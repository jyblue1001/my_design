magic
tech sky130A
timestamp 1738096553
<< error_p >>
rect -1355 332 -1335 335
rect -1355 268 -1352 332
rect -1338 268 -1335 332
rect -1355 265 -1335 268
rect -1135 332 -1115 335
rect -1135 268 -1132 332
rect -1118 268 -1115 332
rect -1135 265 -1115 268
rect -915 332 -895 335
rect -915 268 -912 332
rect -898 268 -895 332
rect -915 265 -895 268
rect -695 332 -675 335
rect -695 268 -692 332
rect -678 268 -675 332
rect -695 265 -675 268
rect -365 332 -345 335
rect -365 268 -362 332
rect -348 268 -345 332
rect -365 265 -345 268
rect -145 332 -125 335
rect -145 268 -142 332
rect -128 268 -125 332
rect -145 265 -125 268
rect 75 332 95 335
rect 75 268 78 332
rect 92 268 95 332
rect 75 265 95 268
rect 295 332 315 335
rect 295 268 298 332
rect 312 268 315 332
rect 295 265 315 268
rect -1355 82 -1335 85
rect -1355 18 -1352 82
rect -1338 18 -1335 82
rect -1355 15 -1335 18
rect -1135 82 -1115 85
rect -1135 18 -1132 82
rect -1118 18 -1115 82
rect -1135 15 -1115 18
rect -695 82 -675 85
rect -695 18 -692 82
rect -678 18 -675 82
rect -695 15 -675 18
rect -475 82 -455 85
rect -475 18 -472 82
rect -458 18 -455 82
rect -475 15 -455 18
rect 75 82 95 85
rect 75 18 78 82
rect 92 18 95 82
rect 75 15 95 18
rect 295 82 315 85
rect 295 18 298 82
rect 312 18 315 82
rect 295 15 315 18
<< nmos >>
rect -2995 200 -2980 400
rect -2845 200 -2830 400
rect -2695 200 -2680 400
rect -2545 200 -2530 400
rect -2395 200 -2380 400
rect -2245 200 -2230 400
rect -2095 200 -2080 400
rect -1945 200 -1930 400
rect -1795 200 -1780 400
rect -1430 250 -1370 350
rect -1320 250 -1260 350
rect -1210 250 -1150 350
rect -1100 250 -1040 350
rect -990 250 -930 350
rect -880 250 -820 350
rect -770 250 -710 350
rect -660 250 -600 350
rect -440 250 -380 350
rect -330 250 -270 350
rect -220 250 -160 350
rect -110 250 -50 350
rect 0 250 60 350
rect 110 250 170 350
rect 220 250 280 350
rect 330 250 390 350
rect -2995 0 -2980 100
rect -2845 0 -2830 100
rect -2695 0 -2680 100
rect -2545 0 -2530 100
rect -2395 0 -2380 100
rect -2245 0 -2230 100
rect -2095 0 -2080 100
rect -1945 0 -1930 100
rect -1795 0 -1780 100
rect -1430 0 -1370 100
rect -1320 0 -1260 100
rect -1210 0 -1150 100
rect -1100 0 -1040 100
rect -770 0 -710 100
rect -660 0 -600 100
rect -550 0 -490 100
rect -440 0 -380 100
rect 0 0 60 100
rect 110 0 170 100
rect 220 0 280 100
rect 330 0 390 100
rect -495 -1300 -480 -1100
rect -345 -1300 -330 -1100
rect -195 -1300 -180 -1100
rect -45 -1300 -30 -1100
rect -495 -1500 -480 -1400
rect -345 -1500 -330 -1400
rect -195 -1500 -180 -1400
rect -45 -1500 -30 -1400
rect 205 -1500 220 -1300
rect -495 -1800 -480 -1600
rect -345 -1800 -330 -1600
rect -195 -1800 -180 -1600
rect -45 -1800 -30 -1600
rect 205 -1700 220 -1600
rect -495 -2000 -480 -1900
rect -345 -2000 -330 -1900
rect -195 -2000 -180 -1900
rect -45 -2000 -30 -1900
<< ndiff >>
rect -3045 385 -2995 400
rect -3045 215 -3030 385
rect -3010 215 -2995 385
rect -3045 200 -2995 215
rect -2980 385 -2930 400
rect -2980 215 -2965 385
rect -2945 215 -2930 385
rect -2980 200 -2930 215
rect -2895 385 -2845 400
rect -2895 215 -2880 385
rect -2860 215 -2845 385
rect -2895 200 -2845 215
rect -2830 385 -2780 400
rect -2830 215 -2815 385
rect -2795 215 -2780 385
rect -2830 200 -2780 215
rect -2745 385 -2695 400
rect -2745 215 -2730 385
rect -2710 215 -2695 385
rect -2745 200 -2695 215
rect -2680 385 -2630 400
rect -2680 215 -2665 385
rect -2645 215 -2630 385
rect -2680 200 -2630 215
rect -2595 385 -2545 400
rect -2595 215 -2580 385
rect -2560 215 -2545 385
rect -2595 200 -2545 215
rect -2530 385 -2480 400
rect -2530 215 -2515 385
rect -2495 215 -2480 385
rect -2530 200 -2480 215
rect -2445 385 -2395 400
rect -2445 215 -2430 385
rect -2410 215 -2395 385
rect -2445 200 -2395 215
rect -2380 385 -2330 400
rect -2380 215 -2365 385
rect -2345 215 -2330 385
rect -2380 200 -2330 215
rect -2295 385 -2245 400
rect -2295 215 -2280 385
rect -2260 215 -2245 385
rect -2295 200 -2245 215
rect -2230 385 -2180 400
rect -2230 215 -2215 385
rect -2195 215 -2180 385
rect -2230 200 -2180 215
rect -2145 385 -2095 400
rect -2145 215 -2130 385
rect -2110 215 -2095 385
rect -2145 200 -2095 215
rect -2080 385 -2030 400
rect -2080 215 -2065 385
rect -2045 215 -2030 385
rect -2080 200 -2030 215
rect -1995 385 -1945 400
rect -1995 215 -1980 385
rect -1960 215 -1945 385
rect -1995 200 -1945 215
rect -1930 385 -1880 400
rect -1930 215 -1915 385
rect -1895 215 -1880 385
rect -1930 200 -1880 215
rect -1845 385 -1795 400
rect -1845 215 -1830 385
rect -1810 215 -1795 385
rect -1845 200 -1795 215
rect -1780 385 -1730 400
rect -1780 215 -1765 385
rect -1745 215 -1730 385
rect -1480 335 -1430 350
rect -1480 265 -1465 335
rect -1445 265 -1430 335
rect -1480 250 -1430 265
rect -1370 335 -1320 350
rect -1370 265 -1355 335
rect -1335 265 -1320 335
rect -1370 250 -1320 265
rect -1260 335 -1210 350
rect -1260 265 -1245 335
rect -1225 265 -1210 335
rect -1260 250 -1210 265
rect -1150 335 -1100 350
rect -1150 265 -1135 335
rect -1115 265 -1100 335
rect -1150 250 -1100 265
rect -1040 335 -990 350
rect -1040 265 -1025 335
rect -1005 265 -990 335
rect -1040 250 -990 265
rect -930 335 -880 350
rect -930 265 -915 335
rect -895 265 -880 335
rect -930 250 -880 265
rect -820 335 -770 350
rect -820 265 -805 335
rect -785 265 -770 335
rect -820 250 -770 265
rect -710 335 -660 350
rect -710 265 -695 335
rect -675 265 -660 335
rect -710 250 -660 265
rect -600 335 -550 350
rect -600 265 -585 335
rect -565 265 -550 335
rect -600 250 -550 265
rect -490 335 -440 350
rect -490 265 -475 335
rect -455 265 -440 335
rect -490 250 -440 265
rect -380 335 -330 350
rect -380 265 -365 335
rect -345 265 -330 335
rect -380 250 -330 265
rect -270 335 -220 350
rect -270 265 -255 335
rect -235 265 -220 335
rect -270 250 -220 265
rect -160 335 -110 350
rect -160 265 -145 335
rect -125 265 -110 335
rect -160 250 -110 265
rect -50 335 0 350
rect -50 265 -35 335
rect -15 265 0 335
rect -50 250 0 265
rect 60 335 110 350
rect 60 265 75 335
rect 95 265 110 335
rect 60 250 110 265
rect 170 335 220 350
rect 170 265 185 335
rect 205 265 220 335
rect 170 250 220 265
rect 280 335 330 350
rect 280 265 295 335
rect 315 265 330 335
rect 280 250 330 265
rect 390 335 440 350
rect 390 265 405 335
rect 425 265 440 335
rect 390 250 440 265
rect -1780 200 -1730 215
rect -3045 85 -2995 100
rect -3045 15 -3030 85
rect -3010 15 -2995 85
rect -3045 0 -2995 15
rect -2980 85 -2930 100
rect -2980 15 -2965 85
rect -2945 15 -2930 85
rect -2980 0 -2930 15
rect -2895 85 -2845 100
rect -2895 15 -2880 85
rect -2860 15 -2845 85
rect -2895 0 -2845 15
rect -2830 85 -2780 100
rect -2830 15 -2815 85
rect -2795 15 -2780 85
rect -2830 0 -2780 15
rect -2745 85 -2695 100
rect -2745 15 -2730 85
rect -2710 15 -2695 85
rect -2745 0 -2695 15
rect -2680 85 -2630 100
rect -2680 15 -2665 85
rect -2645 15 -2630 85
rect -2680 0 -2630 15
rect -2595 85 -2545 100
rect -2595 15 -2580 85
rect -2560 15 -2545 85
rect -2595 0 -2545 15
rect -2530 85 -2480 100
rect -2530 15 -2515 85
rect -2495 15 -2480 85
rect -2530 0 -2480 15
rect -2445 85 -2395 100
rect -2445 15 -2430 85
rect -2410 15 -2395 85
rect -2445 0 -2395 15
rect -2380 85 -2330 100
rect -2380 15 -2365 85
rect -2345 15 -2330 85
rect -2380 0 -2330 15
rect -2295 85 -2245 100
rect -2295 15 -2280 85
rect -2260 15 -2245 85
rect -2295 0 -2245 15
rect -2230 85 -2180 100
rect -2230 15 -2215 85
rect -2195 15 -2180 85
rect -2230 0 -2180 15
rect -2145 85 -2095 100
rect -2145 15 -2130 85
rect -2110 15 -2095 85
rect -2145 0 -2095 15
rect -2080 85 -2030 100
rect -2080 15 -2065 85
rect -2045 15 -2030 85
rect -2080 0 -2030 15
rect -1995 85 -1945 100
rect -1995 15 -1980 85
rect -1960 15 -1945 85
rect -1995 0 -1945 15
rect -1930 85 -1880 100
rect -1930 15 -1915 85
rect -1895 15 -1880 85
rect -1930 0 -1880 15
rect -1845 85 -1795 100
rect -1845 15 -1830 85
rect -1810 15 -1795 85
rect -1845 0 -1795 15
rect -1780 85 -1730 100
rect -1780 15 -1765 85
rect -1745 15 -1730 85
rect -1780 0 -1730 15
rect -1480 85 -1430 100
rect -1480 15 -1465 85
rect -1445 15 -1430 85
rect -1480 0 -1430 15
rect -1370 85 -1320 100
rect -1370 15 -1355 85
rect -1335 15 -1320 85
rect -1370 0 -1320 15
rect -1260 85 -1210 100
rect -1260 15 -1245 85
rect -1225 15 -1210 85
rect -1260 0 -1210 15
rect -1150 85 -1100 100
rect -1150 15 -1135 85
rect -1115 15 -1100 85
rect -1150 0 -1100 15
rect -1040 85 -990 100
rect -1040 15 -1025 85
rect -1005 15 -990 85
rect -1040 0 -990 15
rect -820 85 -770 100
rect -820 15 -805 85
rect -785 15 -770 85
rect -820 0 -770 15
rect -710 85 -660 100
rect -710 15 -695 85
rect -675 15 -660 85
rect -710 0 -660 15
rect -600 85 -550 100
rect -600 15 -585 85
rect -565 15 -550 85
rect -600 0 -550 15
rect -490 85 -440 100
rect -490 15 -475 85
rect -455 15 -440 85
rect -490 0 -440 15
rect -380 85 -330 100
rect -380 15 -365 85
rect -345 15 -330 85
rect -380 0 -330 15
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 60 85 110 100
rect 60 15 75 85
rect 95 15 110 85
rect 60 0 110 15
rect 170 85 220 100
rect 170 15 185 85
rect 205 15 220 85
rect 170 0 220 15
rect 280 85 330 100
rect 280 15 295 85
rect 315 15 330 85
rect 280 0 330 15
rect 390 85 440 100
rect 390 15 405 85
rect 425 15 440 85
rect 390 0 440 15
rect -545 -1115 -495 -1100
rect -545 -1285 -530 -1115
rect -510 -1285 -495 -1115
rect -545 -1300 -495 -1285
rect -480 -1115 -430 -1100
rect -480 -1285 -465 -1115
rect -445 -1285 -430 -1115
rect -480 -1300 -430 -1285
rect -395 -1115 -345 -1100
rect -395 -1285 -380 -1115
rect -360 -1285 -345 -1115
rect -395 -1300 -345 -1285
rect -330 -1115 -280 -1100
rect -330 -1285 -315 -1115
rect -295 -1285 -280 -1115
rect -330 -1300 -280 -1285
rect -245 -1115 -195 -1100
rect -245 -1285 -230 -1115
rect -210 -1285 -195 -1115
rect -245 -1300 -195 -1285
rect -180 -1115 -130 -1100
rect -180 -1285 -165 -1115
rect -145 -1285 -130 -1115
rect -180 -1300 -130 -1285
rect -95 -1115 -45 -1100
rect -95 -1285 -80 -1115
rect -60 -1285 -45 -1115
rect -95 -1300 -45 -1285
rect -30 -1115 20 -1100
rect -30 -1285 -15 -1115
rect 5 -1285 20 -1115
rect -30 -1300 20 -1285
rect 155 -1315 205 -1300
rect -545 -1415 -495 -1400
rect -545 -1485 -530 -1415
rect -510 -1485 -495 -1415
rect -545 -1500 -495 -1485
rect -480 -1415 -430 -1400
rect -480 -1485 -465 -1415
rect -445 -1485 -430 -1415
rect -480 -1500 -430 -1485
rect -395 -1415 -345 -1400
rect -395 -1485 -380 -1415
rect -360 -1485 -345 -1415
rect -395 -1500 -345 -1485
rect -330 -1415 -280 -1400
rect -330 -1485 -315 -1415
rect -295 -1485 -280 -1415
rect -330 -1500 -280 -1485
rect -245 -1415 -195 -1400
rect -245 -1485 -230 -1415
rect -210 -1485 -195 -1415
rect -245 -1500 -195 -1485
rect -180 -1415 -130 -1400
rect -180 -1485 -165 -1415
rect -145 -1485 -130 -1415
rect -180 -1500 -130 -1485
rect -95 -1415 -45 -1400
rect -95 -1485 -80 -1415
rect -60 -1485 -45 -1415
rect -95 -1500 -45 -1485
rect -30 -1415 20 -1400
rect -30 -1485 -15 -1415
rect 5 -1485 20 -1415
rect -30 -1500 20 -1485
rect 155 -1485 170 -1315
rect 190 -1485 205 -1315
rect 155 -1500 205 -1485
rect 220 -1315 270 -1300
rect 220 -1485 235 -1315
rect 255 -1485 270 -1315
rect 220 -1500 270 -1485
rect -545 -1615 -495 -1600
rect -545 -1785 -530 -1615
rect -510 -1785 -495 -1615
rect -545 -1800 -495 -1785
rect -480 -1615 -430 -1600
rect -480 -1785 -465 -1615
rect -445 -1785 -430 -1615
rect -480 -1800 -430 -1785
rect -395 -1615 -345 -1600
rect -395 -1785 -380 -1615
rect -360 -1785 -345 -1615
rect -395 -1800 -345 -1785
rect -330 -1615 -280 -1600
rect -330 -1785 -315 -1615
rect -295 -1785 -280 -1615
rect -330 -1800 -280 -1785
rect -245 -1615 -195 -1600
rect -245 -1785 -230 -1615
rect -210 -1785 -195 -1615
rect -245 -1800 -195 -1785
rect -180 -1615 -130 -1600
rect -180 -1785 -165 -1615
rect -145 -1785 -130 -1615
rect -180 -1800 -130 -1785
rect -95 -1615 -45 -1600
rect -95 -1785 -80 -1615
rect -60 -1785 -45 -1615
rect -95 -1800 -45 -1785
rect -30 -1615 20 -1600
rect -30 -1785 -15 -1615
rect 5 -1785 20 -1615
rect 155 -1615 205 -1600
rect 155 -1685 170 -1615
rect 190 -1685 205 -1615
rect 155 -1700 205 -1685
rect 220 -1615 270 -1600
rect 220 -1685 235 -1615
rect 255 -1685 270 -1615
rect 220 -1700 270 -1685
rect -30 -1800 20 -1785
rect -545 -1915 -495 -1900
rect -545 -1985 -530 -1915
rect -510 -1985 -495 -1915
rect -545 -2000 -495 -1985
rect -480 -1915 -430 -1900
rect -480 -1985 -465 -1915
rect -445 -1985 -430 -1915
rect -480 -2000 -430 -1985
rect -395 -1915 -345 -1900
rect -395 -1985 -380 -1915
rect -360 -1985 -345 -1915
rect -395 -2000 -345 -1985
rect -330 -1915 -280 -1900
rect -330 -1985 -315 -1915
rect -295 -1985 -280 -1915
rect -330 -2000 -280 -1985
rect -245 -1915 -195 -1900
rect -245 -1985 -230 -1915
rect -210 -1985 -195 -1915
rect -245 -2000 -195 -1985
rect -180 -1915 -130 -1900
rect -180 -1985 -165 -1915
rect -145 -1985 -130 -1915
rect -180 -2000 -130 -1985
rect -95 -1915 -45 -1900
rect -95 -1985 -80 -1915
rect -60 -1985 -45 -1915
rect -95 -2000 -45 -1985
rect -30 -1915 20 -1900
rect -30 -1985 -15 -1915
rect 5 -1985 20 -1915
rect -30 -2000 20 -1985
<< ndiffc >>
rect -3030 215 -3010 385
rect -2965 215 -2945 385
rect -2880 215 -2860 385
rect -2815 215 -2795 385
rect -2730 215 -2710 385
rect -2665 215 -2645 385
rect -2580 215 -2560 385
rect -2515 215 -2495 385
rect -2430 215 -2410 385
rect -2365 215 -2345 385
rect -2280 215 -2260 385
rect -2215 215 -2195 385
rect -2130 215 -2110 385
rect -2065 215 -2045 385
rect -1980 215 -1960 385
rect -1915 215 -1895 385
rect -1830 215 -1810 385
rect -1765 215 -1745 385
rect -1465 265 -1445 335
rect -1355 265 -1335 335
rect -1245 265 -1225 335
rect -1135 265 -1115 335
rect -1025 265 -1005 335
rect -915 265 -895 335
rect -805 265 -785 335
rect -695 265 -675 335
rect -585 265 -565 335
rect -475 265 -455 335
rect -365 265 -345 335
rect -255 265 -235 335
rect -145 265 -125 335
rect -35 265 -15 335
rect 75 265 95 335
rect 185 265 205 335
rect 295 265 315 335
rect 405 265 425 335
rect -3030 15 -3010 85
rect -2965 15 -2945 85
rect -2880 15 -2860 85
rect -2815 15 -2795 85
rect -2730 15 -2710 85
rect -2665 15 -2645 85
rect -2580 15 -2560 85
rect -2515 15 -2495 85
rect -2430 15 -2410 85
rect -2365 15 -2345 85
rect -2280 15 -2260 85
rect -2215 15 -2195 85
rect -2130 15 -2110 85
rect -2065 15 -2045 85
rect -1980 15 -1960 85
rect -1915 15 -1895 85
rect -1830 15 -1810 85
rect -1765 15 -1745 85
rect -1465 15 -1445 85
rect -1355 15 -1335 85
rect -1245 15 -1225 85
rect -1135 15 -1115 85
rect -1025 15 -1005 85
rect -805 15 -785 85
rect -695 15 -675 85
rect -585 15 -565 85
rect -475 15 -455 85
rect -365 15 -345 85
rect -35 15 -15 85
rect 75 15 95 85
rect 185 15 205 85
rect 295 15 315 85
rect 405 15 425 85
rect -530 -1285 -510 -1115
rect -465 -1285 -445 -1115
rect -380 -1285 -360 -1115
rect -315 -1285 -295 -1115
rect -230 -1285 -210 -1115
rect -165 -1285 -145 -1115
rect -80 -1285 -60 -1115
rect -15 -1285 5 -1115
rect -530 -1485 -510 -1415
rect -465 -1485 -445 -1415
rect -380 -1485 -360 -1415
rect -315 -1485 -295 -1415
rect -230 -1485 -210 -1415
rect -165 -1485 -145 -1415
rect -80 -1485 -60 -1415
rect -15 -1485 5 -1415
rect 170 -1485 190 -1315
rect 235 -1485 255 -1315
rect -530 -1785 -510 -1615
rect -465 -1785 -445 -1615
rect -380 -1785 -360 -1615
rect -315 -1785 -295 -1615
rect -230 -1785 -210 -1615
rect -165 -1785 -145 -1615
rect -80 -1785 -60 -1615
rect -15 -1785 5 -1615
rect 170 -1685 190 -1615
rect 235 -1685 255 -1615
rect -530 -1985 -510 -1915
rect -465 -1985 -445 -1915
rect -380 -1985 -360 -1915
rect -315 -1985 -295 -1915
rect -230 -1985 -210 -1915
rect -165 -1985 -145 -1915
rect -80 -1985 -60 -1915
rect -15 -1985 5 -1915
<< poly >>
rect -2845 480 -1780 495
rect -2845 455 -2830 480
rect -1795 455 -1780 480
rect -2870 445 -2830 455
rect -2870 425 -2860 445
rect -2840 425 -2830 445
rect -2870 415 -2830 425
rect -2560 445 -2520 455
rect -2560 425 -2550 445
rect -2530 425 -2520 445
rect -2560 415 -2520 425
rect -1795 445 -1755 455
rect -1795 425 -1785 445
rect -1765 425 -1755 445
rect -1795 415 -1755 425
rect -2995 400 -2980 415
rect -2845 400 -2830 415
rect -2695 400 -2680 415
rect -2545 400 -2530 415
rect -2395 400 -2380 415
rect -2245 400 -2230 415
rect -2095 400 -2080 415
rect -1945 400 -1930 415
rect -1795 400 -1780 415
rect -1430 350 -1370 365
rect -1320 350 -1260 365
rect -1210 350 -1150 365
rect -1100 350 -1040 365
rect -990 350 -930 365
rect -880 350 -820 365
rect -770 350 -710 365
rect -660 350 -600 365
rect -440 350 -380 365
rect -330 350 -270 365
rect -220 350 -160 365
rect -110 350 -50 365
rect 0 350 60 365
rect 110 350 170 365
rect 220 350 280 365
rect 330 350 390 365
rect -1430 240 -1370 250
rect -1320 240 -1260 250
rect -1210 240 -1150 250
rect -1100 240 -1040 250
rect -990 240 -930 250
rect -880 240 -820 250
rect -770 240 -710 250
rect -660 240 -600 250
rect -1430 225 -600 240
rect -440 240 -380 250
rect -330 240 -270 250
rect -220 240 -160 250
rect -110 240 -50 250
rect 0 240 60 250
rect 110 240 170 250
rect 220 240 280 250
rect 330 240 390 250
rect -440 225 390 240
rect -2995 155 -2980 200
rect -2845 170 -2830 200
rect -2695 170 -2680 200
rect -2545 185 -2530 200
rect -3060 140 -2980 155
rect -2995 100 -2980 140
rect -2870 160 -2830 170
rect -2870 140 -2860 160
rect -2840 140 -2830 160
rect -2870 130 -2830 140
rect -2720 160 -2680 170
rect -2720 140 -2710 160
rect -2690 140 -2680 160
rect -2395 155 -2380 200
rect -2245 185 -2230 200
rect -2095 185 -2080 200
rect -1945 185 -1930 200
rect -1795 185 -1780 200
rect -2095 170 -1855 185
rect -2720 130 -2680 140
rect -2845 100 -2830 130
rect -2695 125 -2680 130
rect -2470 140 -2380 155
rect -2695 110 -2530 125
rect -2695 100 -2680 110
rect -2545 100 -2530 110
rect -2995 -15 -2980 0
rect -2845 -15 -2830 0
rect -2695 -15 -2680 0
rect -2545 -15 -2530 0
rect -2470 -40 -2455 140
rect -2395 100 -2380 140
rect -2120 160 -2080 170
rect -2120 140 -2110 160
rect -2090 140 -2080 160
rect -2120 130 -2080 140
rect -2245 100 -2230 115
rect -2095 100 -2080 130
rect -1870 125 -1855 170
rect -1690 180 15 195
rect -1690 160 -1675 180
rect -1715 150 -1675 160
rect -1715 130 -1705 150
rect -1685 130 -1675 150
rect -1945 100 -1930 115
rect -1870 110 -1780 125
rect -1715 120 -1675 130
rect -1475 145 -1435 155
rect -1475 125 -1465 145
rect -1445 125 -1435 145
rect -1255 145 -1215 155
rect -1255 125 -1245 145
rect -1225 125 -1215 145
rect -1035 145 -995 155
rect -1035 125 -1025 145
rect -1005 125 -995 145
rect 0 125 15 180
rect -1475 115 -380 125
rect -1465 110 -380 115
rect -1795 100 -1780 110
rect -1430 100 -1370 110
rect -1320 100 -1260 110
rect -1210 100 -1150 110
rect -1100 100 -1040 110
rect -770 100 -710 110
rect -660 100 -600 110
rect -550 100 -490 110
rect -440 100 -380 110
rect 0 110 390 125
rect 0 100 60 110
rect 110 100 170 110
rect 220 100 280 110
rect 330 100 390 110
rect -2395 -15 -2380 0
rect -2245 -15 -2230 0
rect -2095 -15 -2080 0
rect -1945 -15 -1930 0
rect -1795 -15 -1780 0
rect -1430 -15 -1370 0
rect -1320 -15 -1260 0
rect -1210 -15 -1150 0
rect -1100 -15 -1040 0
rect -770 -15 -710 0
rect -660 -15 -600 0
rect -550 -15 -490 0
rect -440 -15 -380 0
rect 0 -15 60 0
rect 110 -15 170 0
rect 220 -15 280 0
rect 330 -15 390 0
rect -3060 -55 -2455 -40
rect -1970 -25 -1930 -15
rect -1970 -45 -1960 -25
rect -1940 -45 -1930 -25
rect -1970 -55 -1930 -45
rect -495 -1100 -480 -1085
rect -345 -1100 -330 -1085
rect -195 -1100 -180 -1085
rect -45 -1090 220 -1075
rect -45 -1100 -30 -1090
rect 205 -1300 220 -1090
rect -495 -1345 -480 -1300
rect -345 -1330 -330 -1300
rect -195 -1330 -180 -1300
rect -45 -1315 -30 -1300
rect -560 -1360 -480 -1345
rect -495 -1400 -480 -1360
rect -370 -1340 -330 -1330
rect -370 -1360 -360 -1340
rect -340 -1360 -330 -1340
rect -370 -1370 -330 -1360
rect -220 -1340 -180 -1330
rect -220 -1360 -210 -1340
rect -190 -1360 -180 -1340
rect -70 -1325 -30 -1315
rect -70 -1345 -60 -1325
rect -40 -1345 -30 -1325
rect -70 -1355 -30 -1345
rect -220 -1370 -180 -1360
rect -345 -1400 -330 -1370
rect -195 -1400 -180 -1370
rect -45 -1400 -30 -1385
rect -495 -1515 -480 -1500
rect -345 -1515 -330 -1500
rect -195 -1515 -180 -1500
rect -45 -1515 -30 -1500
rect 205 -1515 220 -1500
rect -495 -1600 -480 -1585
rect -345 -1600 -330 -1585
rect -195 -1600 -180 -1585
rect -45 -1600 -30 -1585
rect 205 -1600 220 -1585
rect -495 -1845 -480 -1800
rect -345 -1830 -330 -1800
rect -195 -1830 -180 -1800
rect -45 -1815 -30 -1800
rect -560 -1860 -480 -1845
rect -495 -1900 -480 -1860
rect -220 -1840 -180 -1830
rect -220 -1860 -210 -1840
rect -190 -1860 -180 -1840
rect -220 -1870 -180 -1860
rect -345 -1900 -330 -1870
rect -195 -1900 -180 -1870
rect -70 -1855 -30 -1845
rect -70 -1875 -60 -1855
rect -40 -1875 -30 -1855
rect -70 -1885 -30 -1875
rect -45 -1900 -30 -1885
rect -495 -2015 -480 -2000
rect -345 -2015 -330 -2000
rect -195 -2015 -180 -2000
rect -45 -2010 -30 -2000
rect 205 -2010 220 -1700
rect -45 -2025 220 -2010
<< polycont >>
rect -2860 425 -2840 445
rect -2550 425 -2530 445
rect -1785 425 -1765 445
rect -2860 140 -2840 160
rect -2710 140 -2690 160
rect -2110 140 -2090 160
rect -1705 130 -1685 150
rect -1465 125 -1445 145
rect -1245 125 -1225 145
rect -1025 125 -1005 145
rect -1960 -45 -1940 -25
rect -360 -1360 -340 -1340
rect -210 -1360 -190 -1340
rect -60 -1345 -40 -1325
rect -210 -1860 -190 -1840
rect -60 -1875 -40 -1855
<< locali >>
rect -2805 475 -1820 495
rect -2870 445 -2830 455
rect -2870 425 -2860 445
rect -2840 425 -2830 445
rect -2870 415 -2830 425
rect -2805 395 -2785 475
rect -2560 445 -2520 455
rect -2560 435 -2550 445
rect -2665 425 -2550 435
rect -2530 425 -2520 445
rect -2665 415 -2520 425
rect -2665 395 -2645 415
rect -1840 395 -1820 475
rect -1795 445 -1755 455
rect -1795 425 -1785 445
rect -1765 425 -1755 445
rect -1795 415 -1755 425
rect -3040 385 -3000 395
rect -3040 215 -3030 385
rect -3010 215 -3000 385
rect -3040 205 -3000 215
rect -2975 385 -2935 395
rect -2975 215 -2965 385
rect -2945 215 -2935 385
rect -2975 205 -2935 215
rect -2890 385 -2850 395
rect -2890 215 -2880 385
rect -2860 215 -2850 385
rect -2890 205 -2850 215
rect -2825 385 -2785 395
rect -2825 215 -2815 385
rect -2795 215 -2785 385
rect -2825 205 -2785 215
rect -2740 385 -2700 395
rect -2740 215 -2730 385
rect -2710 215 -2700 385
rect -2740 205 -2700 215
rect -2675 385 -2635 395
rect -2675 215 -2665 385
rect -2645 215 -2635 385
rect -2675 205 -2635 215
rect -2590 385 -2550 395
rect -2590 215 -2580 385
rect -2560 215 -2550 385
rect -2590 205 -2550 215
rect -2525 385 -2485 395
rect -2525 215 -2515 385
rect -2495 215 -2485 385
rect -2525 205 -2485 215
rect -2440 385 -2400 395
rect -2440 215 -2430 385
rect -2410 215 -2400 385
rect -2440 205 -2400 215
rect -2375 385 -2335 395
rect -2375 215 -2365 385
rect -2345 215 -2335 385
rect -2375 205 -2335 215
rect -2290 385 -2250 395
rect -2290 215 -2280 385
rect -2260 215 -2250 385
rect -2290 205 -2250 215
rect -2225 385 -2185 395
rect -2225 215 -2215 385
rect -2195 215 -2185 385
rect -2225 205 -2185 215
rect -2140 385 -2100 395
rect -2140 215 -2130 385
rect -2110 215 -2100 385
rect -2140 205 -2100 215
rect -2075 385 -2035 395
rect -2075 215 -2065 385
rect -2045 215 -2035 385
rect -2075 205 -2035 215
rect -1990 385 -1950 395
rect -1990 215 -1980 385
rect -1960 215 -1950 385
rect -1990 205 -1950 215
rect -1925 385 -1885 395
rect -1925 215 -1915 385
rect -1895 215 -1885 385
rect -1925 205 -1885 215
rect -1840 385 -1800 395
rect -1840 215 -1830 385
rect -1810 215 -1800 385
rect -1840 205 -1800 215
rect -1775 385 -1735 395
rect -1775 215 -1765 385
rect -1745 215 -1735 385
rect -1465 365 -565 385
rect -1465 345 -1445 365
rect -1355 345 -1335 365
rect -1245 345 -1225 365
rect -1135 345 -1115 365
rect -1025 345 -1005 365
rect -915 345 -895 365
rect -805 345 -785 365
rect -695 345 -675 365
rect -585 345 -565 365
rect -475 365 425 385
rect -475 345 -455 365
rect -365 345 -345 365
rect -255 345 -235 365
rect -145 345 -125 365
rect -35 345 -15 365
rect 75 345 95 365
rect 185 345 205 365
rect 295 345 315 365
rect 405 345 425 365
rect -1475 335 -1435 345
rect -1475 265 -1465 335
rect -1445 265 -1435 335
rect -1475 255 -1435 265
rect -1365 335 -1325 345
rect -1365 265 -1355 335
rect -1335 265 -1325 335
rect -1365 255 -1325 265
rect -1255 335 -1215 345
rect -1255 265 -1245 335
rect -1225 265 -1215 335
rect -1255 255 -1215 265
rect -1145 335 -1105 345
rect -1145 265 -1135 335
rect -1115 265 -1105 335
rect -1145 255 -1105 265
rect -1035 335 -995 345
rect -1035 265 -1025 335
rect -1005 265 -995 335
rect -1035 255 -995 265
rect -925 335 -885 345
rect -925 265 -915 335
rect -895 265 -885 335
rect -925 255 -885 265
rect -815 335 -775 345
rect -815 265 -805 335
rect -785 265 -775 335
rect -815 255 -775 265
rect -705 335 -665 345
rect -705 265 -695 335
rect -675 265 -665 335
rect -705 255 -665 265
rect -595 335 -555 345
rect -595 265 -585 335
rect -565 265 -555 335
rect -595 255 -555 265
rect -485 335 -445 345
rect -485 265 -475 335
rect -455 265 -445 335
rect -485 255 -445 265
rect -375 335 -335 345
rect -375 265 -365 335
rect -345 265 -335 335
rect -375 255 -335 265
rect -265 335 -225 345
rect -265 265 -255 335
rect -235 265 -225 335
rect -265 255 -225 265
rect -155 335 -115 345
rect -155 265 -145 335
rect -125 265 -115 335
rect -155 255 -115 265
rect -45 335 -5 345
rect -45 265 -35 335
rect -15 265 -5 335
rect -45 255 -5 265
rect 65 335 105 345
rect 65 265 75 335
rect 95 265 105 335
rect 65 255 105 265
rect 175 335 215 345
rect 175 265 185 335
rect 205 265 215 335
rect 175 255 215 265
rect 285 335 325 345
rect 285 265 295 335
rect 315 265 325 335
rect 285 255 325 265
rect 395 335 435 345
rect 395 265 405 335
rect 425 265 435 335
rect 395 255 435 265
rect -1775 205 -1735 215
rect -2955 160 -2935 205
rect -2870 160 -2830 170
rect -2955 140 -2860 160
rect -2840 140 -2830 160
rect -2955 95 -2935 140
rect -2870 130 -2830 140
rect -2805 160 -2785 205
rect -2720 160 -2680 170
rect -2805 140 -2710 160
rect -2690 140 -2680 160
rect -2805 95 -2785 140
rect -2720 130 -2680 140
rect -2655 95 -2635 205
rect -2580 95 -2560 205
rect -2515 95 -2495 205
rect -2355 160 -2335 205
rect -2280 160 -2260 205
rect -2355 140 -2260 160
rect -2355 95 -2335 140
rect -2280 95 -2260 140
rect -2215 160 -2195 205
rect -2120 160 -2080 170
rect -2215 140 -2110 160
rect -2090 140 -2080 160
rect -2215 95 -2195 140
rect -2120 130 -2080 140
rect -2055 95 -2035 205
rect -1980 95 -1960 205
rect -1915 95 -1895 205
rect -1715 150 -1675 160
rect -1715 130 -1705 150
rect -1685 130 -1675 150
rect -1715 120 -1675 130
rect -1475 145 -1435 155
rect -1475 125 -1465 145
rect -1445 125 -1435 145
rect -1475 115 -1435 125
rect -1255 145 -1215 155
rect -1255 125 -1245 145
rect -1225 125 -1215 145
rect -1255 115 -1215 125
rect -1035 145 -995 155
rect -1035 125 -1025 145
rect -1005 125 -995 145
rect -1035 115 -995 125
rect -1465 95 -1445 115
rect -1245 95 -1225 115
rect -1025 95 -1005 115
rect -585 95 -565 255
rect 405 95 425 255
rect -3040 85 -3000 95
rect -3040 15 -3030 85
rect -3010 15 -3000 85
rect -3040 5 -3000 15
rect -2975 85 -2935 95
rect -2975 15 -2965 85
rect -2945 15 -2935 85
rect -2975 5 -2935 15
rect -2890 85 -2850 95
rect -2890 15 -2880 85
rect -2860 15 -2850 85
rect -2890 5 -2850 15
rect -2825 85 -2785 95
rect -2825 15 -2815 85
rect -2795 15 -2785 85
rect -2825 5 -2785 15
rect -2740 85 -2700 95
rect -2740 15 -2730 85
rect -2710 15 -2700 85
rect -2740 5 -2700 15
rect -2675 85 -2635 95
rect -2675 15 -2665 85
rect -2645 15 -2635 85
rect -2675 5 -2635 15
rect -2590 85 -2550 95
rect -2590 15 -2580 85
rect -2560 15 -2550 85
rect -2590 5 -2550 15
rect -2525 85 -2485 95
rect -2525 15 -2515 85
rect -2495 15 -2485 85
rect -2525 5 -2485 15
rect -2440 85 -2400 95
rect -2440 15 -2430 85
rect -2410 15 -2400 85
rect -2440 5 -2400 15
rect -2375 85 -2335 95
rect -2375 15 -2365 85
rect -2345 15 -2335 85
rect -2375 5 -2335 15
rect -2290 85 -2250 95
rect -2290 15 -2280 85
rect -2260 15 -2250 85
rect -2290 5 -2250 15
rect -2225 85 -2185 95
rect -2225 15 -2215 85
rect -2195 15 -2185 85
rect -2225 5 -2185 15
rect -2140 85 -2100 95
rect -2140 15 -2130 85
rect -2110 15 -2100 85
rect -2140 5 -2100 15
rect -2075 85 -2035 95
rect -2075 15 -2065 85
rect -2045 15 -2035 85
rect -2075 5 -2035 15
rect -1990 85 -1950 95
rect -1990 15 -1980 85
rect -1960 15 -1950 85
rect -1990 5 -1950 15
rect -1925 85 -1885 95
rect -1925 15 -1915 85
rect -1895 25 -1885 85
rect -1840 85 -1800 95
rect -1840 25 -1830 85
rect -1895 15 -1830 25
rect -1810 15 -1800 85
rect -1925 5 -1800 15
rect -1775 85 -1735 95
rect -1775 15 -1765 85
rect -1745 15 -1735 85
rect -1775 5 -1735 15
rect -1475 85 -1435 95
rect -1475 15 -1465 85
rect -1445 15 -1435 85
rect -1475 5 -1435 15
rect -1365 85 -1325 95
rect -1365 15 -1355 85
rect -1335 15 -1325 85
rect -1365 5 -1325 15
rect -1255 85 -1215 95
rect -1255 15 -1245 85
rect -1225 15 -1215 85
rect -1255 5 -1215 15
rect -1145 85 -1105 95
rect -1145 15 -1135 85
rect -1115 15 -1105 85
rect -1145 5 -1105 15
rect -1035 85 -995 95
rect -1035 15 -1025 85
rect -1005 15 -995 85
rect -1035 5 -995 15
rect -815 85 -775 95
rect -815 15 -805 85
rect -785 15 -775 85
rect -815 5 -775 15
rect -705 85 -665 95
rect -705 15 -695 85
rect -675 15 -665 85
rect -705 5 -665 15
rect -595 85 -555 95
rect -595 15 -585 85
rect -565 15 -555 85
rect -595 5 -555 15
rect -485 85 -445 95
rect -485 15 -475 85
rect -455 15 -445 85
rect -485 5 -445 15
rect -375 85 -335 95
rect -375 15 -365 85
rect -345 15 -335 85
rect -375 5 -335 15
rect -45 85 -5 95
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 5 -5 15
rect 65 85 105 95
rect 65 15 75 85
rect 95 15 105 85
rect 65 5 105 15
rect 175 85 215 95
rect 175 15 185 85
rect 205 15 215 85
rect 175 5 215 15
rect 285 85 325 95
rect 285 15 295 85
rect 315 15 325 85
rect 285 5 325 15
rect 395 85 435 95
rect 395 15 405 85
rect 425 15 435 85
rect 395 5 435 15
rect -2055 -15 -2035 5
rect -1465 -15 -1445 5
rect -1355 -15 -1335 5
rect -1245 -15 -1225 5
rect -1135 -15 -1115 5
rect -1025 -15 -1005 5
rect -2055 -25 -1930 -15
rect -2055 -35 -1960 -25
rect -1970 -45 -1960 -35
rect -1940 -45 -1930 -25
rect -1465 -35 -1005 -15
rect -805 -15 -785 5
rect -695 -15 -675 5
rect -585 -15 -565 5
rect -475 -15 -455 5
rect -365 -15 -345 5
rect -805 -35 -345 -15
rect -35 -15 -15 5
rect 75 -15 95 5
rect 185 -15 205 5
rect 295 -15 315 5
rect 405 -15 425 5
rect -35 -35 425 -15
rect -1970 -55 -1930 -45
rect -540 -1115 -500 -1105
rect -540 -1285 -530 -1115
rect -510 -1285 -500 -1115
rect -540 -1295 -500 -1285
rect -475 -1115 -435 -1105
rect -475 -1285 -465 -1115
rect -445 -1285 -435 -1115
rect -475 -1295 -435 -1285
rect -390 -1115 -350 -1105
rect -390 -1285 -380 -1115
rect -360 -1285 -350 -1115
rect -390 -1295 -350 -1285
rect -325 -1115 -285 -1105
rect -325 -1285 -315 -1115
rect -295 -1285 -285 -1115
rect -325 -1295 -285 -1285
rect -240 -1115 -200 -1105
rect -240 -1285 -230 -1115
rect -210 -1285 -200 -1115
rect -240 -1295 -200 -1285
rect -175 -1115 -135 -1105
rect -175 -1285 -165 -1115
rect -145 -1285 -135 -1115
rect -175 -1295 -135 -1285
rect -90 -1115 -50 -1105
rect -90 -1285 -80 -1115
rect -60 -1285 -50 -1115
rect -90 -1295 -50 -1285
rect -25 -1115 15 -1105
rect -25 -1285 -15 -1115
rect 5 -1285 15 -1115
rect -25 -1295 15 -1285
rect -455 -1340 -435 -1295
rect -370 -1340 -330 -1330
rect -455 -1360 -360 -1340
rect -340 -1360 -330 -1340
rect -455 -1405 -435 -1360
rect -370 -1370 -330 -1360
rect -305 -1340 -285 -1295
rect -155 -1315 -135 -1295
rect -5 -1315 15 -1295
rect 160 -1315 200 -1305
rect -155 -1325 -30 -1315
rect -220 -1340 -180 -1330
rect -305 -1360 -210 -1340
rect -190 -1360 -180 -1340
rect -305 -1405 -285 -1360
rect -220 -1370 -180 -1360
rect -155 -1335 -60 -1325
rect -155 -1405 -135 -1335
rect -70 -1345 -60 -1335
rect -40 -1345 -30 -1325
rect -70 -1355 -30 -1345
rect -5 -1335 170 -1315
rect -5 -1405 15 -1335
rect -540 -1415 -500 -1405
rect -540 -1485 -530 -1415
rect -510 -1485 -500 -1415
rect -540 -1495 -500 -1485
rect -475 -1415 -435 -1405
rect -475 -1485 -465 -1415
rect -445 -1485 -435 -1415
rect -475 -1495 -435 -1485
rect -390 -1415 -350 -1405
rect -390 -1485 -380 -1415
rect -360 -1485 -350 -1415
rect -390 -1495 -350 -1485
rect -325 -1415 -285 -1405
rect -325 -1485 -315 -1415
rect -295 -1485 -285 -1415
rect -325 -1495 -285 -1485
rect -240 -1415 -200 -1405
rect -240 -1485 -230 -1415
rect -210 -1485 -200 -1415
rect -240 -1495 -200 -1485
rect -175 -1415 -135 -1405
rect -175 -1485 -165 -1415
rect -145 -1485 -135 -1415
rect -175 -1495 -135 -1485
rect -90 -1415 -50 -1405
rect -90 -1485 -80 -1415
rect -60 -1485 -50 -1415
rect -90 -1495 -50 -1485
rect -25 -1415 15 -1405
rect -25 -1485 -15 -1415
rect 5 -1485 15 -1415
rect -25 -1495 15 -1485
rect 160 -1485 170 -1335
rect 190 -1485 200 -1315
rect 160 -1495 200 -1485
rect 225 -1315 265 -1305
rect 225 -1485 235 -1315
rect 255 -1485 265 -1315
rect 225 -1495 265 -1485
rect -540 -1615 -500 -1605
rect -540 -1785 -530 -1615
rect -510 -1785 -500 -1615
rect -540 -1795 -500 -1785
rect -475 -1615 -435 -1605
rect -475 -1785 -465 -1615
rect -445 -1785 -435 -1615
rect -475 -1795 -435 -1785
rect -390 -1615 -350 -1605
rect -390 -1785 -380 -1615
rect -360 -1785 -350 -1615
rect -390 -1795 -350 -1785
rect -325 -1615 -285 -1605
rect -325 -1785 -315 -1615
rect -295 -1785 -285 -1615
rect -325 -1795 -285 -1785
rect -240 -1615 -200 -1605
rect -240 -1785 -230 -1615
rect -210 -1785 -200 -1615
rect -240 -1795 -200 -1785
rect -175 -1615 -135 -1605
rect -175 -1785 -165 -1615
rect -145 -1785 -135 -1615
rect -175 -1795 -135 -1785
rect -90 -1615 -50 -1605
rect -90 -1785 -80 -1615
rect -60 -1785 -50 -1615
rect -90 -1795 -50 -1785
rect -25 -1615 15 -1605
rect -25 -1785 -15 -1615
rect 5 -1785 15 -1615
rect 160 -1615 200 -1605
rect 160 -1685 170 -1615
rect 190 -1685 200 -1615
rect 160 -1695 200 -1685
rect 225 -1615 265 -1605
rect 225 -1685 235 -1615
rect 255 -1685 265 -1615
rect 225 -1695 265 -1685
rect -25 -1795 15 -1785
rect -455 -1840 -435 -1795
rect -380 -1840 -360 -1795
rect -455 -1860 -360 -1840
rect -455 -1905 -435 -1860
rect -380 -1905 -360 -1860
rect -315 -1840 -295 -1795
rect -220 -1840 -180 -1830
rect -315 -1860 -210 -1840
rect -190 -1860 -180 -1840
rect -315 -1905 -295 -1860
rect -220 -1870 -180 -1860
rect -155 -1855 -135 -1795
rect -5 -1835 15 -1795
rect 170 -1835 190 -1695
rect -70 -1855 -30 -1845
rect -155 -1875 -60 -1855
rect -40 -1875 -30 -1855
rect -155 -1905 -135 -1875
rect -70 -1885 -30 -1875
rect -5 -1860 190 -1835
rect -5 -1905 15 -1860
rect -540 -1915 -500 -1905
rect -540 -1985 -530 -1915
rect -510 -1985 -500 -1915
rect -540 -1995 -500 -1985
rect -475 -1915 -435 -1905
rect -475 -1985 -465 -1915
rect -445 -1985 -435 -1915
rect -475 -1995 -435 -1985
rect -390 -1915 -350 -1905
rect -390 -1985 -380 -1915
rect -360 -1985 -350 -1915
rect -390 -1995 -350 -1985
rect -325 -1915 -285 -1905
rect -325 -1985 -315 -1915
rect -295 -1985 -285 -1915
rect -325 -1995 -285 -1985
rect -240 -1915 -200 -1905
rect -240 -1985 -230 -1915
rect -210 -1985 -200 -1915
rect -240 -1995 -200 -1985
rect -175 -1915 -135 -1905
rect -175 -1985 -165 -1915
rect -145 -1985 -135 -1915
rect -175 -1995 -135 -1985
rect -90 -1915 -50 -1905
rect -90 -1985 -80 -1915
rect -60 -1985 -50 -1915
rect -90 -1995 -50 -1985
rect -25 -1915 15 -1905
rect -25 -1985 -15 -1915
rect 5 -1985 15 -1915
rect -25 -1995 15 -1985
<< viali >>
rect -1355 265 -1335 335
rect -1135 265 -1115 335
rect -915 265 -895 335
rect -695 265 -675 335
rect -365 265 -345 335
rect -145 265 -125 335
rect 75 265 95 335
rect 295 265 315 335
rect -1355 15 -1335 85
rect -1135 15 -1115 85
rect -695 15 -675 85
rect -475 15 -455 85
rect 75 15 95 85
rect 295 15 315 85
<< end >>
