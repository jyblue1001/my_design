* PEX produced on Sun Jun 29 09:46:22 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_4.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_4 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 a_n8798_9160.t1 a_n7190_9280.t1 GNDA.t138 sky130_fd_pr__res_xhigh_po_0p35 l=6
X1 VDDA.t429 ref_volt_cur_gen_dummy_magic_0.V_mir2.t17 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t10 VDDA.t428 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X2 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA.t324 GNDA.t326 GNDA.t325 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X3 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t11 ref_volt_cur_gen_dummy_magic_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VDDA.t350 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 VDDA.t349 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X8 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t11 ref_volt_cur_gen_dummy_magic_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_0.V_err_gate.t12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDDA.t458 ref_volt_cur_gen_dummy_magic_0.V_mir1.t14 ref_volt_cur_gen_dummy_magic_0.V_mir1.t15 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X13 GNDA.t32 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X14 two_stage_opamp_dummy_magic_0.X.t13 GNDA.t321 GNDA.t323 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X15 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 VDDA.t58 two_stage_opamp_dummy_magic_0.X.t26 VOUT-.t5 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X19 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_0.Y.t25 VDDA.t89 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X20 VDDA.t220 VDDA.t217 VDDA.t219 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X21 ref_volt_cur_gen_dummy_magic_0.V_TOP.t14 VDDA.t309 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t352 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X23 ref_volt_cur_gen_dummy_magic_0.V_p_2.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 ref_volt_cur_gen_dummy_magic_0.V_mir2.t2 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X24 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 GNDA.t238 GNDA.t319 ref_volt_cur_gen_dummy_magic_0.Vbe2.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X26 VDDA.t27 ref_volt_cur_gen_dummy_magic_0.V_TOP.t15 ref_volt_cur_gen_dummy_magic_0.START_UP.t5 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X27 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5750_2946.t0 GNDA.t51 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X28 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VDDA.t377 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X32 ref_volt_cur_gen_dummy_magic_0.V_p_1.t7 ref_volt_cur_gen_dummy_magic_0.Vin+.t6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t7 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X33 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X34 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VDDA.t460 ref_volt_cur_gen_dummy_magic_0.V_TOP.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X37 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 GNDA.t119 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X39 GNDA.t229 GNDA.t320 ref_volt_cur_gen_dummy_magic_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X40 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t12 ref_volt_cur_gen_dummy_magic_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VDDA.t80 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.VD3.t8 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X43 VDDA.t216 VDDA.t214 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X44 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 two_stage_opamp_dummy_magic_0.Y.t15 GNDA.t316 GNDA.t318 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X47 two_stage_opamp_dummy_magic_0.Y.t12 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD1.t11 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X48 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t379 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X51 VOUT-.t6 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X52 two_stage_opamp_dummy_magic_0.V_p.t3 two_stage_opamp_dummy_magic_0.Vb1.t0 two_stage_opamp_dummy_magic_0.Vb1.t1 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.3
X53 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X54 VDDA.t441 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t12 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t9 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X55 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t13 ref_volt_cur_gen_dummy_magic_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 VDDA.t474 two_stage_opamp_dummy_magic_0.Vb3.t17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 VDDA.t473 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X58 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t5 GNDA.t164 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X59 two_stage_opamp_dummy_magic_0.VD1.t14 VIN-.t0 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X60 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X64 VDDA.t231 ref_volt_cur_gen_dummy_magic_0.V_TOP.t17 ref_volt_cur_gen_dummy_magic_0.Vin+.t4 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X65 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 GNDA.t133 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X68 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 GNDA.t176 ref_volt_cur_gen_dummy_magic_0.START_UP_NFET1.t1 ref_volt_cur_gen_dummy_magic_0.START_UP_NFET1.t0 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X70 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t1 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X71 VDDA.t71 two_stage_opamp_dummy_magic_0.Vb3.t18 two_stage_opamp_dummy_magic_0.VD3.t7 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X72 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 two_stage_opamp_dummy_magic_0.X.t16 two_stage_opamp_dummy_magic_0.Vb2.t9 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X74 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t13 ref_volt_cur_gen_dummy_magic_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 GNDA.t47 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 VOUT+.t1 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X77 GNDA.t208 two_stage_opamp_dummy_magic_0.X.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X78 GNDA.t64 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X79 VDDA.t439 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t14 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t8 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X80 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t313 GNDA.t315 GNDA.t314 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X81 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 GNDA.t312 GNDA.t310 two_stage_opamp_dummy_magic_0.VD1.t18 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X83 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t14 ref_volt_cur_gen_dummy_magic_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT+.t14 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t272 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X89 GNDA.t309 GNDA.t307 GNDA.t309 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X90 GNDA.t306 GNDA.t304 two_stage_opamp_dummy_magic_0.VD1.t17 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X91 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t211 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.5
X92 VDDA.t50 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X93 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 ref_volt_cur_gen_dummy_magic_0.V_TOP.t18 VDDA.t331 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 GNDA.t303 GNDA.t301 VOUT+.t18 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X96 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_0.X.t29 VDDA.t375 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X97 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t15 ref_volt_cur_gen_dummy_magic_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.Vb2.t10 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X99 a_5230_5852.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA.t150 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X100 GNDA.t300 GNDA.t298 two_stage_opamp_dummy_magic_0.X.t12 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X101 GNDA.t297 GNDA.t295 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA.t296 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X102 GNDA.t124 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t2 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t3 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X103 ref_volt_cur_gen_dummy_magic_0.V_TOP.t19 VDDA.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X105 VOUT-.t16 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X106 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t4 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t3 ref_volt_cur_gen_dummy_magic_0.V_p_2.t5 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X112 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 VDDA.t210 VDDA.t208 two_stage_opamp_dummy_magic_0.Vb1.t3 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X115 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t7 ref_volt_cur_gen_dummy_magic_0.V_mir2.t18 VDDA.t427 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X117 VDDA.t207 VDDA.t205 two_stage_opamp_dummy_magic_0.VD3.t11 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X118 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t6 GNDA.t170 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X119 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 ref_volt_cur_gen_dummy_magic_0.V_TOP.t20 VDDA.t285 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 GNDA.t137 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X122 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t16 ref_volt_cur_gen_dummy_magic_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VDDA.t382 two_stage_opamp_dummy_magic_0.X.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X125 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X126 ref_volt_cur_gen_dummy_magic_0.V_mir1.t13 ref_volt_cur_gen_dummy_magic_0.V_mir1.t12 VDDA.t445 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X127 GNDA.t220 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X128 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 GNDA.t294 GNDA.t292 two_stage_opamp_dummy_magic_0.Y.t14 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X130 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t17 ref_volt_cur_gen_dummy_magic_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 GNDA.t125 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X132 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 ref_volt_cur_gen_dummy_magic_0.V_TOP.t21 VDDA.t468 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 GNDA.t66 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X135 GNDA.t126 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 VDDA.t255 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X136 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X137 ref_volt_cur_gen_dummy_magic_0.Vin+.t3 ref_volt_cur_gen_dummy_magic_0.V_TOP.t22 VDDA.t260 VDDA.t259 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X138 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 two_stage_opamp_dummy_magic_0.V_p.t33 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X141 ref_volt_cur_gen_dummy_magic_0.V_mir2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 ref_volt_cur_gen_dummy_magic_0.V_p_2.t9 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X142 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t12 VDDA.t346 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X144 VOUT-.t7 a_5750_2946.t1 GNDA.t71 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X145 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t6 ref_volt_cur_gen_dummy_magic_0.Vin+.t7 ref_volt_cur_gen_dummy_magic_0.V_p_1.t6 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X148 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t18 ref_volt_cur_gen_dummy_magic_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t13 two_stage_opamp_dummy_magic_0.Y.t29 VDDA.t284 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X150 two_stage_opamp_dummy_magic_0.V_p.t20 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X151 two_stage_opamp_dummy_magic_0.V_p.t32 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X152 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VDDA.t248 ref_volt_cur_gen_dummy_magic_0.V_mir1.t17 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t8 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X155 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X156 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VDDA.t201 VDDA.t199 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X158 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 a_n9700_9790.t1 GNDA.t149 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X162 VOUT+.t17 GNDA.t289 GNDA.t291 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X163 a_14520_5852.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X164 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t14 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X165 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t7 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t15 VDDA.t437 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X166 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 two_stage_opamp_dummy_magic_0.VD2.t3 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t6 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X169 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t16 ref_volt_cur_gen_dummy_magic_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 VOUT-.t3 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X173 VOUT-.t4 two_stage_opamp_dummy_magic_0.X.t35 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X174 VDDA.t65 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X175 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 VOUT-.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X178 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t17 ref_volt_cur_gen_dummy_magic_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t4 GNDA.t70 sky130_fd_pr__res_high_po_1p41 l=1.41
X180 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 GNDA.t43 two_stage_opamp_dummy_magic_0.Y.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X182 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.Vb3.t20 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X184 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.X.t17 two_stage_opamp_dummy_magic_0.VD3.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X186 two_stage_opamp_dummy_magic_0.err_amp_out.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X187 VDDA.t204 VDDA.t202 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.5
X188 VDDA.t9 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X189 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t18 ref_volt_cur_gen_dummy_magic_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 GNDA.t238 GNDA.t288 ref_volt_cur_gen_dummy_magic_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X191 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 ref_volt_cur_gen_dummy_magic_0.START_UP_NFET1.t0 ref_volt_cur_gen_dummy_magic_0.START_UP.t0 ref_volt_cur_gen_dummy_magic_0.START_UP.t1 GNDA.t355 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X193 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t1 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t4 ref_volt_cur_gen_dummy_magic_0.V_p_2.t2 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X194 two_stage_opamp_dummy_magic_0.VD1.t10 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X195 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t19 VDDA.t435 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X198 VDDA.t198 VDDA.t196 two_stage_opamp_dummy_magic_0.V_err_p.t4 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X199 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 GNDA.t158 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X203 two_stage_opamp_dummy_magic_0.err_amp_out.t11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X204 GNDA.t1 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X205 GNDA.t174 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X206 VDDA.t42 ref_volt_cur_gen_dummy_magic_0.V_mir1.t10 ref_volt_cur_gen_dummy_magic_0.V_mir1.t11 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t20 ref_volt_cur_gen_dummy_magic_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_0.V_p.t31 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t335 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X214 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 two_stage_opamp_dummy_magic_0.V_p.t18 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA.t24 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X216 VDDA.t299 two_stage_opamp_dummy_magic_0.Vb3.t21 two_stage_opamp_dummy_magic_0.VD4.t15 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X217 VOUT+.t12 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X218 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X219 two_stage_opamp_dummy_magic_0.Vb3.t9 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t9 GNDA.t218 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X220 two_stage_opamp_dummy_magic_0.V_p.t38 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t344 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X221 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA.t285 GNDA.t287 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X222 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t19 ref_volt_cur_gen_dummy_magic_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 ref_volt_cur_gen_dummy_magic_0.V_TOP.t23 VDDA.t463 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t1 VDDA.t193 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X226 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t12 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X227 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X228 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VDDA.t348 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X233 two_stage_opamp_dummy_magic_0.VD2.t20 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t22 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X234 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 ref_volt_cur_gen_dummy_magic_0.V_p_2.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 ref_volt_cur_gen_dummy_magic_0.V_mir2.t0 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X236 GNDA.t284 GNDA.t282 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X237 ref_volt_cur_gen_dummy_magic_0.cap_res1.t20 ref_volt_cur_gen_dummy_magic_0.V_TOP.t13 GNDA.t127 sky130_fd_pr__res_high_po_0p35 l=2.05
X238 VOUT-.t14 two_stage_opamp_dummy_magic_0.X.t38 VDDA.t301 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X239 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VDDA.t16 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X241 VDDA.t308 ref_volt_cur_gen_dummy_magic_0.V_mir1.t8 ref_volt_cur_gen_dummy_magic_0.V_mir1.t9 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X242 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t190 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X248 GNDA.t86 two_stage_opamp_dummy_magic_0.Y.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X249 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VDDA.t189 VDDA.t187 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.5
X251 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.VD4.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 GNDA.t87 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X253 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t343 GNDA.t342 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X256 VDDA.t447 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t20 ref_volt_cur_gen_dummy_magic_0.V_TOP.t12 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X257 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA.t198 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X258 VDDA.t302 two_stage_opamp_dummy_magic_0.X.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X259 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 VDDA.t305 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X261 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t21 ref_volt_cur_gen_dummy_magic_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 VDDA.t450 ref_volt_cur_gen_dummy_magic_0.V_TOP.t24 ref_volt_cur_gen_dummy_magic_0.Vin-.t6 VDDA.t449 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X264 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 two_stage_opamp_dummy_magic_0.VD1.t9 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t8 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X266 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VDDA.t8 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t11 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X268 VDDA.t325 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t324 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X269 GNDA.t115 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X270 ref_volt_cur_gen_dummy_magic_0.V_p_2.t3 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t5 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t2 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X271 GNDA.t26 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X272 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X273 GNDA.t117 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 VOUT-.t12 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X274 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t3 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X275 two_stage_opamp_dummy_magic_0.V_p.t4 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t12 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X276 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 GNDA.t196 two_stage_opamp_dummy_magic_0.err_amp_out.t12 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X278 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t14 VDDA.t341 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X282 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VDDA.t24 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.VD3.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X284 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t9 ref_volt_cur_gen_dummy_magic_0.V_mir1.t18 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X286 VOUT+.t11 two_stage_opamp_dummy_magic_0.Y.t36 VDDA.t295 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X287 two_stage_opamp_dummy_magic_0.V_p.t30 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t19 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X288 two_stage_opamp_dummy_magic_0.V_p.t16 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA.t60 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X289 VOUT+.t10 two_stage_opamp_dummy_magic_0.Y.t37 VDDA.t297 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X290 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t16 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X291 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 GNDA.t21 a_n9700_9790.t0 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X294 ref_volt_cur_gen_dummy_magic_0.V_p_2.t1 VDDA.t475 GNDA.t333 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X295 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t21 ref_volt_cur_gen_dummy_magic_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 a_14640_5852.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA.t14 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X297 VDDA.t425 ref_volt_cur_gen_dummy_magic_0.V_mir2.t7 ref_volt_cur_gen_dummy_magic_0.V_mir2.t8 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X298 ref_volt_cur_gen_dummy_magic_0.V_TOP.t6 VDDA.t476 GNDA.t334 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X299 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_0.Vb3.t5 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t11 GNDA.t167 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X303 GNDA.t246 GNDA.t281 ref_volt_cur_gen_dummy_magic_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X304 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t6 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X305 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t5 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X306 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t33 two_stage_opamp_dummy_magic_0.VD4.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X307 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VDDA.t268 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X310 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 ref_volt_cur_gen_dummy_magic_0.START_UP.t4 ref_volt_cur_gen_dummy_magic_0.V_TOP.t25 VDDA.t472 VDDA.t471 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X314 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_0.VD4.t17 VDDA.t184 VDDA.t186 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X318 ref_volt_cur_gen_dummy_magic_0.V_TOP.t26 VDDA.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X320 GNDA.t49 VDDA.t181 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X321 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X322 ref_volt_cur_gen_dummy_magic_0.V_p_2.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 ref_volt_cur_gen_dummy_magic_0.V_mir2.t1 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X323 VDDA.t423 ref_volt_cur_gen_dummy_magic_0.V_mir2.t15 ref_volt_cur_gen_dummy_magic_0.V_mir2.t16 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X324 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VDDA.t306 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X328 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 two_stage_opamp_dummy_magic_0.Vb2.t6 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t12 GNDA.t35 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X330 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA.t278 GNDA.t280 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X331 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 two_stage_opamp_dummy_magic_0.VD1.t8 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.Y.t24 GNDA.t350 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X333 VDDA.t44 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X334 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 GNDA.t62 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_p_mir.t1 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X336 ref_volt_cur_gen_dummy_magic_0.V_TOP.t1 ref_volt_cur_gen_dummy_magic_0.START_UP.t6 ref_volt_cur_gen_dummy_magic_0.Vin-.t2 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X337 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X338 ref_volt_cur_gen_dummy_magic_0.V_mir1.t7 ref_volt_cur_gen_dummy_magic_0.V_mir1.t6 VDDA.t454 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X339 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 GNDA.t152 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X343 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X344 two_stage_opamp_dummy_magic_0.V_p.t2 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X345 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t15 VDDA.t343 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X347 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 ref_volt_cur_gen_dummy_magic_0.V_p_1.t10 ref_volt_cur_gen_dummy_magic_0.Vin-.t8 ref_volt_cur_gen_dummy_magic_0.V_mir1.t16 GNDA.t352 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X349 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.Vb3.t23 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X350 two_stage_opamp_dummy_magic_0.Vb2.t2 two_stage_opamp_dummy_magic_0.Vb2.t1 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X351 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.Y.t18 two_stage_opamp_dummy_magic_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X352 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t22 ref_volt_cur_gen_dummy_magic_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 GNDA.t238 GNDA.t237 ref_volt_cur_gen_dummy_magic_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X354 VOUT+.t4 VDDA.t178 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X355 two_stage_opamp_dummy_magic_0.V_p.t24 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X356 ref_volt_cur_gen_dummy_magic_0.V_TOP.t27 VDDA.t330 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 two_stage_opamp_dummy_magic_0.V_p.t14 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t154 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X358 two_stage_opamp_dummy_magic_0.Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t21 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t23 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t22 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.24 ps=2 w=0.6 l=0.2
X359 GNDA.t229 GNDA.t233 ref_volt_cur_gen_dummy_magic_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X360 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 VDDA.t175 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.32 ps=2.4 w=0.8 l=0.2
X361 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t16 VDDA.t393 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X362 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t5 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t22 VDDA.t433 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X363 two_stage_opamp_dummy_magic_0.Vb2.t5 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t13 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X364 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 ref_volt_cur_gen_dummy_magic_0.cap_res2.t0 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t3 GNDA.t127 sky130_fd_pr__res_high_po_0p35 l=2.05
X367 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 ref_volt_cur_gen_dummy_magic_0.V_TOP.t28 VDDA.t328 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 ref_volt_cur_gen_dummy_magic_0.V_mir2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 ref_volt_cur_gen_dummy_magic_0.V_p_2.t6 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X370 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VDDA.t174 VDDA.t172 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X372 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t10 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X373 two_stage_opamp_dummy_magic_0.VD2.t11 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t14 GNDA.t327 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X374 ref_volt_cur_gen_dummy_magic_0.V_mir1.t5 ref_volt_cur_gen_dummy_magic_0.V_mir1.t4 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X375 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VDDA.t269 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X378 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t169 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.5
X380 VDDA.t280 two_stage_opamp_dummy_magic_0.Y.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X381 VDDA.t421 ref_volt_cur_gen_dummy_magic_0.V_mir2.t19 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t9 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X382 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t250 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X384 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.Y.t4 GNDA.t142 sky130_fd_pr__res_high_po_1p41 l=1.41
X385 two_stage_opamp_dummy_magic_0.VD4.t29 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Y.t19 two_stage_opamp_dummy_magic_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X386 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 VDDA.t166 VDDA.t168 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X387 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t23 ref_volt_cur_gen_dummy_magic_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 two_stage_opamp_dummy_magic_0.V_err_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X390 ref_volt_cur_gen_dummy_magic_0.V_mir1.t3 ref_volt_cur_gen_dummy_magic_0.Vin-.t9 ref_volt_cur_gen_dummy_magic_0.V_p_1.t9 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X391 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.VD3.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X393 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA.t348 GNDA.t347 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X395 two_stage_opamp_dummy_magic_0.Vb3.t8 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t14 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X396 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t4 GNDA.t275 GNDA.t277 GNDA.t276 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X397 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 ref_volt_cur_gen_dummy_magic_0.V_TOP.t29 VDDA.t312 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t24 ref_volt_cur_gen_dummy_magic_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VDDA.t456 ref_volt_cur_gen_dummy_magic_0.V_TOP.t30 ref_volt_cur_gen_dummy_magic_0.Vin-.t5 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X402 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t229 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X403 two_stage_opamp_dummy_magic_0.VD1.t7 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t5 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X404 VDDA.t2 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X405 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X406 two_stage_opamp_dummy_magic_0.VD1.t6 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X407 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VDDA.t165 VDDA.t163 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t0 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X411 two_stage_opamp_dummy_magic_0.Vb1.t5 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t17 VDDA.t395 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X412 GNDA.t274 GNDA.t271 GNDA.t273 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X413 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 two_stage_opamp_dummy_magic_0.V_err_p.t19 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X414 GNDA.t187 VDDA.t121 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X415 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t25 ref_volt_cur_gen_dummy_magic_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 two_stage_opamp_dummy_magic_0.V_p.t28 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t16 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X418 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VDDA.t337 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t336 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X422 VDDA.t4 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t8 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X423 VDDA.t162 VDDA.t160 GNDA.t48 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X424 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 a_14640_5852.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t161 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X427 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t23 ref_volt_cur_gen_dummy_magic_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 GNDA.t189 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X429 ref_volt_cur_gen_dummy_magic_0.V_mir2.t14 ref_volt_cur_gen_dummy_magic_0.V_mir2.t13 VDDA.t419 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X430 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VOUT+.t2 a_14240_2946.t0 GNDA.t54 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X432 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t26 ref_volt_cur_gen_dummy_magic_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VDDA.t314 ref_volt_cur_gen_dummy_magic_0.V_TOP.t31 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X436 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X438 VDDA.t159 VDDA.t157 ref_volt_cur_gen_dummy_magic_0.V_TOP.t5 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X439 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VDDA.t339 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X441 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t7 VDDA.t452 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X444 VDDA.t156 VDDA.t154 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t0 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X445 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X446 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_0.X.t42 GNDA.t186 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X447 VOUT-.t10 VDDA.t151 VDDA.t153 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X448 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t4 ref_volt_cur_gen_dummy_magic_0.Vin+.t8 ref_volt_cur_gen_dummy_magic_0.V_p_1.t5 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X449 VDDA.t405 GNDA.t268 GNDA.t270 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X450 VDDA.t88 two_stage_opamp_dummy_magic_0.Vb3.t26 two_stage_opamp_dummy_magic_0.VD4.t12 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X451 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 ref_volt_cur_gen_dummy_magic_0.V_TOP.t32 VDDA.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 GNDA.t102 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X455 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 ref_volt_cur_gen_dummy_magic_0.V_mir2.t12 ref_volt_cur_gen_dummy_magic_0.V_mir2.t11 VDDA.t417 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X457 VDDA.t150 VDDA.t148 VOUT+.t3 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X458 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X460 ref_volt_cur_gen_dummy_magic_0.V_TOP.t4 VDDA.t145 VDDA.t147 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X461 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 ref_volt_cur_gen_dummy_magic_0.V_TOP.t33 VDDA.t358 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA.t265 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X465 VOUT+.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t39 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X466 GNDA.t238 GNDA.t264 ref_volt_cur_gen_dummy_magic_0.Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X467 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 GNDA.t229 GNDA.t228 ref_volt_cur_gen_dummy_magic_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X471 two_stage_opamp_dummy_magic_0.V_err_gate.t9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X472 VDDA.t222 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t24 ref_volt_cur_gen_dummy_magic_0.V_TOP.t11 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X473 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VDDA.t321 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X475 VDDA.t367 two_stage_opamp_dummy_magic_0.X.t43 VOUT-.t15 VDDA.t366 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X476 ref_volt_cur_gen_dummy_magic_0.V_mir1.t0 ref_volt_cur_gen_dummy_magic_0.Vin-.t10 ref_volt_cur_gen_dummy_magic_0.V_p_1.t0 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X477 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t142 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X478 VDDA.t242 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD4.t11 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X479 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X483 two_stage_opamp_dummy_magic_0.V_p.t37 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t341 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X484 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t25 ref_volt_cur_gen_dummy_magic_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.Vb3.t28 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X486 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT+.t16 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t110 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X488 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.VD3.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X489 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_0.Y.t41 GNDA.t136 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X492 ref_volt_cur_gen_dummy_magic_0.V_TOP.t34 VDDA.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t27 ref_volt_cur_gen_dummy_magic_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 ref_volt_cur_gen_dummy_magic_0.Vin-.t4 ref_volt_cur_gen_dummy_magic_0.V_TOP.t35 VDDA.t462 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X496 VDDA.t333 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X497 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t1 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t21 VDDA.t335 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X498 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VDDA.t399 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t26 ref_volt_cur_gen_dummy_magic_0.V_TOP.t10 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X500 VDDA.t304 two_stage_opamp_dummy_magic_0.Vb3.t29 two_stage_opamp_dummy_magic_0.VD4.t10 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X501 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 GNDA.t331 VDDA.t477 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t2 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X503 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 two_stage_opamp_dummy_magic_0.V_p.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA.t205 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X505 two_stage_opamp_dummy_magic_0.V_p.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA.t207 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X506 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_0.X.t44 GNDA.t122 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X507 two_stage_opamp_dummy_magic_0.VD2.t4 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.X.t8 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X508 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb3.t30 VDDA.t386 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X509 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t18 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t19 sky130_fd_pr__pfet_01v8 ad=0.24 pd=2 as=0.12 ps=1 w=0.6 l=0.2
X510 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t5 ref_volt_cur_gen_dummy_magic_0.V_mir2.t20 VDDA.t415 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X511 VDDA.t141 VDDA.t139 GNDA.t67 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X512 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t22 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X514 GNDA.t332 VDDA.t478 ref_volt_cur_gen_dummy_magic_0.V_p_1.t1 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X515 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 two_stage_opamp_dummy_magic_0.VD1.t15 VIN-.t6 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X517 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 ref_volt_cur_gen_dummy_magic_0.V_p_1.t4 ref_volt_cur_gen_dummy_magic_0.Vin+.t9 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t3 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X523 GNDA.t73 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X524 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 a_5230_5852.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X526 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t19 two_stage_opamp_dummy_magic_0.VD3.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X527 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t28 ref_volt_cur_gen_dummy_magic_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 GNDA.t82 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X529 VDDA.t226 two_stage_opamp_dummy_magic_0.Y.t42 VOUT+.t9 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X530 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 ref_volt_cur_gen_dummy_magic_0.V_TOP.t36 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X531 two_stage_opamp_dummy_magic_0.VD1.t21 VIN-.t7 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA.t346 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X532 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t23 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X534 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t24 VDDA.t317 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X538 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VDDA.t288 two_stage_opamp_dummy_magic_0.Vb3.t31 two_stage_opamp_dummy_magic_0.VD4.t9 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X541 VDDA.t404 GNDA.t261 GNDA.t263 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X542 two_stage_opamp_dummy_magic_0.Y.t20 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X543 VDDA.t413 ref_volt_cur_gen_dummy_magic_0.V_mir2.t5 ref_volt_cur_gen_dummy_magic_0.V_mir2.t6 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X544 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X545 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t29 ref_volt_cur_gen_dummy_magic_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VDDA.t253 two_stage_opamp_dummy_magic_0.X.t45 VOUT-.t13 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X548 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 VDDA.t138 VDDA.t136 VOUT-.t9 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X550 two_stage_opamp_dummy_magic_0.V_err_gate.t13 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t17 GNDA.t354 GNDA.t353 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X551 GNDA.t260 GNDA.t258 VDDA.t403 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X552 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 ref_volt_cur_gen_dummy_magic_0.V_TOP.t3 VDDA.t133 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X555 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 a_14520_5852.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t13 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X558 VDDA.t411 ref_volt_cur_gen_dummy_magic_0.V_mir2.t21 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t8 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X559 VDDA.t362 ref_volt_cur_gen_dummy_magic_0.V_mir1.t19 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t10 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X560 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_2946.t1 GNDA.t96 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X563 ref_volt_cur_gen_dummy_magic_0.Vin-.t3 ref_volt_cur_gen_dummy_magic_0.V_TOP.t37 VDDA.t465 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X564 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_0.Y.t43 GNDA.t88 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X565 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 GNDA.t257 GNDA.t255 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X569 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.VD3.t30 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.VD3.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X570 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.X.t46 VDDA.t363 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X571 ref_volt_cur_gen_dummy_magic_0.V_TOP.t9 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t27 VDDA.t401 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X572 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 two_stage_opamp_dummy_magic_0.Y.t11 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X575 ref_volt_cur_gen_dummy_magic_0.V_p_2.t0 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t0 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X576 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 ref_volt_cur_gen_dummy_magic_0.V_p_1.t2 ref_volt_cur_gen_dummy_magic_0.Vin-.t11 ref_volt_cur_gen_dummy_magic_0.V_mir1.t1 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X578 GNDA.t9 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 VOUT-.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X579 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X581 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t28 ref_volt_cur_gen_dummy_magic_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t11 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X584 two_stage_opamp_dummy_magic_0.VD4.t8 two_stage_opamp_dummy_magic_0.Vb3.t32 VDDA.t373 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X585 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 two_stage_opamp_dummy_magic_0.VD2.t6 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.X.t9 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X587 two_stage_opamp_dummy_magic_0.V_p.t10 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X588 VDDA.t132 VDDA.t130 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X589 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_0.X.t47 GNDA.t185 VDDA.t364 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X590 VDDA.t384 two_stage_opamp_dummy_magic_0.Vb3.t33 two_stage_opamp_dummy_magic_0.VD3.t15 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X591 GNDA.t98 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 VOUT+.t15 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X592 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 ref_volt_cur_gen_dummy_magic_0.V_TOP.t38 VDDA.t329 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VDDA.t319 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 VDDA.t318 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X595 GNDA.t78 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X596 VDDA.t292 two_stage_opamp_dummy_magic_0.Y.t44 VOUT+.t8 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X597 GNDA.t222 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X598 GNDA.t232 GNDA.t230 VOUT-.t18 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X599 two_stage_opamp_dummy_magic_0.VD2.t21 VIN+.t7 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA.t360 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X600 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 ref_volt_cur_gen_dummy_magic_0.V_TOP.t8 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t29 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X602 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 ref_volt_cur_gen_dummy_magic_0.V_TOP.t39 VDDA.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 VDDA.t103 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.5
X606 two_stage_opamp_dummy_magic_0.V_err_gate.t3 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X607 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 ref_volt_cur_gen_dummy_magic_0.V_p_1.t3 ref_volt_cur_gen_dummy_magic_0.Vin+.t10 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X609 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X612 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 VDDA.t39 two_stage_opamp_dummy_magic_0.X.t48 VOUT-.t2 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X615 VDDA.t101 two_stage_opamp_dummy_magic_0.Vb3.t34 two_stage_opamp_dummy_magic_0.VD3.t9 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X616 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 two_stage_opamp_dummy_magic_0.Y.t45 VDDA.t293 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X617 VDDA.t467 ref_volt_cur_gen_dummy_magic_0.V_TOP.t40 ref_volt_cur_gen_dummy_magic_0.Vin+.t2 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X618 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X619 ref_volt_cur_gen_dummy_magic_0.V_TOP.t41 VDDA.t315 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t30 ref_volt_cur_gen_dummy_magic_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 VDDA.t105 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t27 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X622 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t46 GNDA.t129 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X624 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t130 VDDA.t267 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X627 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 ref_volt_cur_gen_dummy_magic_0.V_TOP.t7 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t30 VDDA.t397 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X629 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.Vb3.t35 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X630 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 GNDA.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X632 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t40 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X633 GNDA.t254 GNDA.t252 VDDA.t402 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X634 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t31 ref_volt_cur_gen_dummy_magic_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X636 two_stage_opamp_dummy_magic_0.Vb1.t2 VDDA.t127 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X637 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 VDDA.t431 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t32 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t4 VDDA.t430 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X640 two_stage_opamp_dummy_magic_0.Y.t16 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t4 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X641 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t31 ref_volt_cur_gen_dummy_magic_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X645 two_stage_opamp_dummy_magic_0.V_p.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X646 two_stage_opamp_dummy_magic_0.V_err_p.t15 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X647 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_0.X.t50 GNDA.t76 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X648 two_stage_opamp_dummy_magic_0.VD2.t18 VIN+.t8 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA.t340 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X649 GNDA.t251 GNDA.t249 GNDA.t251 GNDA.t250 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X650 a_5350_5852.t0 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t160 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X651 two_stage_opamp_dummy_magic_0.X.t20 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X652 GNDA.t248 GNDA.t247 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X653 VDDA.t258 ref_volt_cur_gen_dummy_magic_0.V_TOP.t42 ref_volt_cur_gen_dummy_magic_0.START_UP.t3 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X654 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t33 ref_volt_cur_gen_dummy_magic_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t1 ref_volt_cur_gen_dummy_magic_0.V_mir1.t20 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X656 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 VDDA.t75 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t28 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t1 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X659 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t32 ref_volt_cur_gen_dummy_magic_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 two_stage_opamp_dummy_magic_0.VD3.t10 VDDA.t124 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X662 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 VDDA.t277 two_stage_opamp_dummy_magic_0.Y.t48 VOUT+.t7 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X664 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 two_stage_opamp_dummy_magic_0.VD2.t16 VIN+.t9 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA.t338 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X667 a_n8798_9040.t0 a_n7190_9400.t0 GNDA.t95 sky130_fd_pr__res_xhigh_po_0p35 l=6
X668 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.Vb3.t36 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X669 VDDA.t279 two_stage_opamp_dummy_magic_0.Y.t49 VOUT+.t6 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X670 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 GNDA.t357 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA.t356 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X672 a_n8798_9040.t1 ref_volt_cur_gen_dummy_magic_0.Vin+.t5 GNDA.t138 sky130_fd_pr__res_xhigh_po_0p35 l=6
X673 GNDA.t246 GNDA.t245 ref_volt_cur_gen_dummy_magic_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X674 ref_volt_cur_gen_dummy_magic_0.V_mir2.t10 ref_volt_cur_gen_dummy_magic_0.V_mir2.t9 VDDA.t409 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X675 GNDA.t12 a_n9760_9260.t0 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=6
X676 VOUT-.t17 GNDA.t242 GNDA.t244 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X677 ref_volt_cur_gen_dummy_magic_0.V_TOP.t43 VDDA.t256 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 two_stage_opamp_dummy_magic_0.V_err_gate.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X679 two_stage_opamp_dummy_magic_0.X.t15 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X680 ref_volt_cur_gen_dummy_magic_0.V_TOP.t44 VDDA.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 VDDA.t97 two_stage_opamp_dummy_magic_0.X.t51 VOUT-.t8 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X682 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 two_stage_opamp_dummy_magic_0.Y.t50 VDDA.t289 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X683 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t2 ref_volt_cur_gen_dummy_magic_0.V_mir1.t21 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X685 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t33 ref_volt_cur_gen_dummy_magic_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t19 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X688 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 VOUT-.t11 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X691 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 VDDA.t244 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X693 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_0.Y.t51 GNDA.t140 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X694 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 ref_volt_cur_gen_dummy_magic_0.V_TOP.t45 VDDA.t451 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.VD4.t0 two_stage_opamp_dummy_magic_0.Y.t9 two_stage_opamp_dummy_magic_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X697 GNDA.t172 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X698 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t3 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t7 ref_volt_cur_gen_dummy_magic_0.V_p_2.t4 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X699 GNDA.t200 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X700 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2.t32 two_stage_opamp_dummy_magic_0.Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X702 ref_volt_cur_gen_dummy_magic_0.V_mir1.t2 ref_volt_cur_gen_dummy_magic_0.Vin-.t12 ref_volt_cur_gen_dummy_magic_0.V_p_1.t8 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X703 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t354 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X704 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t34 ref_volt_cur_gen_dummy_magic_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 VDDA.t99 two_stage_opamp_dummy_magic_0.Vb3.t37 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X706 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 two_stage_opamp_dummy_magic_0.Y.t6 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t3 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X708 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 two_stage_opamp_dummy_magic_0.V_err_p.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X710 ref_volt_cur_gen_dummy_magic_0.Vin+.t1 ref_volt_cur_gen_dummy_magic_0.V_TOP.t46 VDDA.t262 VDDA.t261 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X711 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.Vb3.t38 VDDA.t443 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X712 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 ref_volt_cur_gen_dummy_magic_0.V_TOP.t47 VDDA.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 ref_volt_cur_gen_dummy_magic_0.Vin-.t1 ref_volt_cur_gen_dummy_magic_0.START_UP.t7 ref_volt_cur_gen_dummy_magic_0.V_TOP.t0 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X715 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X716 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t29 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X717 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t35 ref_volt_cur_gen_dummy_magic_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 two_stage_opamp_dummy_magic_0.V_p.t6 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t359 GNDA.t358 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X719 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t8 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X720 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA.t239 GNDA.t241 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X721 two_stage_opamp_dummy_magic_0.V_p_mir.t2 VIN-.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t349 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X722 two_stage_opamp_dummy_magic_0.VD1.t13 VIN-.t9 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X723 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 GNDA.t106 a_n7190_9400.t1 GNDA.t105 sky130_fd_pr__res_xhigh_po_0p35 l=6
X728 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t34 ref_volt_cur_gen_dummy_magic_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VDDA.t94 ref_volt_cur_gen_dummy_magic_0.V_mir1.t22 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t5 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X732 VDDA.t120 VDDA.t118 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.4 as=0.16 ps=1.2 w=0.8 l=0.2
X733 VDDA.t274 two_stage_opamp_dummy_magic_0.Y.t52 VOUT+.t5 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X734 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 a_n8798_9160.t0 ref_volt_cur_gen_dummy_magic_0.Vin-.t0 GNDA.t138 sky130_fd_pr__res_xhigh_po_0p35 l=6
X736 two_stage_opamp_dummy_magic_0.VD1.t1 VIN-.t10 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X737 GNDA.t56 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X738 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t2 a_n9760_9260.t1 GNDA.t108 sky130_fd_pr__res_xhigh_po_0p35 l=6
X739 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 ref_volt_cur_gen_dummy_magic_0.V_TOP.t48 VDDA.t264 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X742 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 ref_volt_cur_gen_dummy_magic_0.START_UP.t2 ref_volt_cur_gen_dummy_magic_0.V_TOP.t49 VDDA.t470 VDDA.t469 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X745 two_stage_opamp_dummy_magic_0.V_err_gate.t1 VDDA.t115 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X746 two_stage_opamp_dummy_magic_0.V_err_gate.t0 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X747 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t36 ref_volt_cur_gen_dummy_magic_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.Vb3.t39 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X749 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X750 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t0 VDDA.t112 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X751 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.Vb2.t33 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X752 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_0.Y.t53 VDDA.t275 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X754 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_0.Y.t54 VDDA.t265 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X757 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t6 ref_volt_cur_gen_dummy_magic_0.V_mir2.t22 VDDA.t407 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X761 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VDDA.t238 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t5 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X766 ref_volt_cur_gen_dummy_magic_0.Vbe2.t0 ref_volt_cur_gen_dummy_magic_0.Vin+.t0 GNDA.t104 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X767 GNDA.t193 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X768 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t35 ref_volt_cur_gen_dummy_magic_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 GNDA.t94 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X771 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X773 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_0.X.t53 VDDA.t355 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X775 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t36 ref_volt_cur_gen_dummy_magic_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X778 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t240 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X779 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.Vb2.t34 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X780 GNDA.t75 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X781 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 a_5350_5852.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t351 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X783 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 two_stage_opamp_dummy_magic_0.V_p_mir.t0 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t58 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X787 VDDA.t111 VDDA.t109 ref_volt_cur_gen_dummy_magic_0.V_TOP.t2 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X788 two_stage_opamp_dummy_magic_0.V_err_p.t21 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t7 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X789 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t177 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X790 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA.t234 GNDA.t236 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X792 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 GNDA.t182 a_n7190_9280.t0 GNDA.t181 sky130_fd_pr__res_xhigh_po_0p35 l=6
X794 two_stage_opamp_dummy_magic_0.VD2.t17 VIN+.t10 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X795 two_stage_opamp_dummy_magic_0.Vb2.t3 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t23 GNDA.t224 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X796 GNDA.t227 GNDA.t225 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X797 VDDA.t108 VDDA.t106 two_stage_opamp_dummy_magic_0.VD4.t16 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X798 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 a_n8798_9160.t0 a_n8798_9160.t1 258.591
R1 a_n7190_9280.t0 a_n7190_9280.t1 376.99
R2 GNDA.n1549 GNDA.n1548 59084.7
R3 GNDA.n570 GNDA.n569 41670.6
R4 GNDA.n567 GNDA.n566 41670.6
R5 GNDA.n726 GNDA.n725 41223.8
R6 GNDA.n724 GNDA.n549 32661.5
R7 GNDA.n720 GNDA.n549 32661.5
R8 GNDA.n569 GNDA.n564 30739.1
R9 GNDA.n567 GNDA.n564 30739.1
R10 GNDA.n1546 GNDA.n813 29808.3
R11 GNDA.n569 GNDA.n568 29723.7
R12 GNDA.n719 GNDA.n585 28430.8
R13 GNDA.n725 GNDA.n563 28430.8
R14 GNDA.n723 GNDA.n722 28372.4
R15 GNDA.n722 GNDA.n721 27462.1
R16 GNDA.n1547 GNDA.n1546 26648.4
R17 GNDA.n813 GNDA.n487 26086.2
R18 GNDA.n568 GNDA.n567 25662.2
R19 GNDA.n570 GNDA.n565 25113.6
R20 GNDA.n566 GNDA.n565 24015.7
R21 GNDA.n1548 GNDA.n487 22164.5
R22 GNDA.n1547 GNDA.n812 20494.1
R23 GNDA.n1550 GNDA.n1549 20492.6
R24 GNDA.n764 GNDA.n549 19630.8
R25 GNDA.n722 GNDA.n549 19630.8
R26 GNDA.n721 GNDA.n720 14782.8
R27 GNDA.n724 GNDA.n723 14773.1
R28 GNDA.n820 GNDA.n815 12361.8
R29 GNDA.n819 GNDA.n815 12312.5
R30 GNDA.n2467 GNDA.n2466 12175.2
R31 GNDA.n1544 GNDA.n820 11918.5
R32 GNDA.n1544 GNDA.n819 11869.2
R33 GNDA.n1548 GNDA.n1547 11169.2
R34 GNDA.n1550 GNDA.n487 11132.4
R35 GNDA.n765 GNDA.n547 10835
R36 GNDA.n765 GNDA.n548 10835
R37 GNDA.n763 GNDA.n547 10835
R38 GNDA.n763 GNDA.n548 10835
R39 GNDA.n1546 GNDA.n1545 10371.4
R40 GNDA.n719 GNDA.n718 10371.4
R41 GNDA.n722 GNDA.n564 9476.92
R42 GNDA.n729 GNDA.n527 9308.25
R43 GNDA.n769 GNDA.n527 9308.25
R44 GNDA.n729 GNDA.n528 9308.25
R45 GNDA.n769 GNDA.n528 9308.25
R46 GNDA.n711 GNDA.n586 9259
R47 GNDA.n711 GNDA.n589 8914.25
R48 GNDA.n497 GNDA.n488 8911.86
R49 GNDA.n1551 GNDA.n466 8878.67
R50 GNDA.n568 GNDA.n565 8677.78
R51 GNDA.n1561 GNDA.n478 8175.5
R52 GNDA.n705 GNDA.n586 8175.5
R53 GNDA.n1565 GNDA.n478 8126.25
R54 GNDA.n854 GNDA.n852 7880
R55 GNDA.n1535 GNDA.n852 7880
R56 GNDA.n1493 GNDA.n1485 7880
R57 GNDA.n1493 GNDA.n1486 7880
R58 GNDA.n855 GNDA.n854 7830.75
R59 GNDA.n1535 GNDA.n855 7830.75
R60 GNDA.n1485 GNDA.n1476 7830.75
R61 GNDA.n1486 GNDA.n1476 7830.75
R62 GNDA.n705 GNDA.n589 7830.75
R63 GNDA.n1561 GNDA.n479 7732.25
R64 GNDA.n716 GNDA.n511 7732.25
R65 GNDA.n798 GNDA.n511 7732.25
R66 GNDA.n716 GNDA.n512 7732.25
R67 GNDA.n798 GNDA.n512 7732.25
R68 GNDA.n655 GNDA.n595 7732.25
R69 GNDA.n655 GNDA.n596 7732.25
R70 GNDA.n657 GNDA.n595 7732.25
R71 GNDA.n657 GNDA.n596 7732.25
R72 GNDA.n1565 GNDA.n479 7683
R73 GNDA.n1553 GNDA.n484 6845.75
R74 GNDA.n1553 GNDA.n485 6845.75
R75 GNDA.n1558 GNDA.n484 6796.5
R76 GNDA.n1558 GNDA.n485 6796.5
R77 GNDA.n1932 GNDA.n467 6698
R78 GNDA.n1936 GNDA.n467 6698
R79 GNDA.n1932 GNDA.n468 6648.75
R80 GNDA.n1936 GNDA.n468 6648.75
R81 GNDA.n1468 GNDA.n816 6254.75
R82 GNDA.n1525 GNDA.n816 6254.75
R83 GNDA.n1468 GNDA.n818 6254.75
R84 GNDA.n1525 GNDA.n818 6254.75
R85 GNDA.n648 GNDA.n601 6057.75
R86 GNDA.n648 GNDA.n603 6057.75
R87 GNDA.n649 GNDA.n601 6057.75
R88 GNDA.n649 GNDA.n603 6057.75
R89 GNDA.n803 GNDA.n506 6057.75
R90 GNDA.n804 GNDA.n506 6057.75
R91 GNDA.n804 GNDA.n509 6057.75
R92 GNDA.n803 GNDA.n509 6057.75
R93 GNDA.n1393 GNDA.n1278 5502.84
R94 GNDA.n1464 GNDA.n1459 5368.25
R95 GNDA.n1532 GNDA.n1459 5368.25
R96 GNDA.n1464 GNDA.n1460 5368.25
R97 GNDA.n1532 GNDA.n1460 5368.25
R98 GNDA.n1481 GNDA.n1472 5368.25
R99 GNDA.n1504 GNDA.n1472 5368.25
R100 GNDA.n1481 GNDA.n1473 5368.25
R101 GNDA.n1504 GNDA.n1473 5368.25
R102 GNDA.n576 GNDA.n489 5338.7
R103 GNDA.n632 GNDA.n609 5338.7
R104 GNDA.n576 GNDA.n490 5319
R105 GNDA.n632 GNDA.n610 5319
R106 GNDA.n810 GNDA.n489 5289.45
R107 GNDA.n627 GNDA.n609 5289.45
R108 GNDA.n810 GNDA.n490 5269.75
R109 GNDA.n627 GNDA.n610 5269.75
R110 GNDA.n584 GNDA.n572 5171.25
R111 GNDA.n639 GNDA.n604 5171.25
R112 GNDA.n580 GNDA.n572 5122
R113 GNDA.n635 GNDA.n604 5122
R114 GNDA.n1521 GNDA.n1512 4974.25
R115 GNDA.n1521 GNDA.n1516 4974.25
R116 GNDA.n584 GNDA.n573 4944.7
R117 GNDA.n639 GNDA.n605 4944.7
R118 GNDA.n741 GNDA.n550 4925
R119 GNDA.n755 GNDA.n550 4925
R120 GNDA.n580 GNDA.n573 4895.45
R121 GNDA.n635 GNDA.n605 4895.45
R122 GNDA.n723 GNDA.n563 4826.13
R123 GNDA.n721 GNDA.n571 4816.22
R124 GNDA.n741 GNDA.n551 4728
R125 GNDA.n755 GNDA.n551 4728
R126 GNDA.n1401 GNDA.n475 4678.75
R127 GNDA.n1405 GNDA.n475 4629.5
R128 GNDA.n1401 GNDA.n477 4629.5
R129 GNDA.n1731 GNDA.n1729 4580.25
R130 GNDA.n1731 GNDA.n1730 4580.25
R131 GNDA.n1405 GNDA.n477 4580.25
R132 GNDA.n1738 GNDA.n1737 4580.25
R133 GNDA.n1737 GNDA.n1736 4580.25
R134 GNDA.n1512 GNDA.n1510 4531
R135 GNDA.n1516 GNDA.n1510 4531
R136 GNDA.n1742 GNDA.n1729 4481.75
R137 GNDA.n1742 GNDA.n1730 4481.75
R138 GNDA.n1738 GNDA.n1728 4481.75
R139 GNDA.n1736 GNDA.n1728 4481.75
R140 GNDA.n1551 GNDA.n1550 4377.76
R141 GNDA.n1242 GNDA.n813 4091.78
R142 GNDA.n1938 GNDA.n1937 3691.95
R143 GNDA.n732 GNDA.n557 3595.25
R144 GNDA.n738 GNDA.n557 3595.25
R145 GNDA.n732 GNDA.n558 3250.5
R146 GNDA.n738 GNDA.n558 3250.5
R147 GNDA.n1939 GNDA.n1938 3225.54
R148 GNDA.n773 GNDA.n525 3053.5
R149 GNDA.n773 GNDA.n526 3004.25
R150 GNDA.n1937 GNDA.n466 2978.29
R151 GNDA.n774 GNDA.n525 2955
R152 GNDA.n725 GNDA.n724 2933.33
R153 GNDA.n720 GNDA.n719 2933.33
R154 GNDA.n774 GNDA.n526 2905.75
R155 GNDA.n571 GNDA.n488 2582.96
R156 GNDA.n1549 GNDA.n488 2582.96
R157 GNDA.n1497 GNDA.n1474 2371.15
R158 GNDA.n1500 GNDA.n1474 2371.15
R159 GNDA.n494 GNDA.n493 2326.02
R160 GNDA.n498 GNDA.n493 2326.02
R161 GNDA.n623 GNDA.n614 2326.02
R162 GNDA.n616 GNDA.n614 2326.02
R163 GNDA.n626 GNDA.n624 2310.78
R164 GNDA.n1482 GNDA.n812 2121.65
R165 GNDA.n812 GNDA.n811 1469.8
R166 GNDA.n1475 GNDA.n1474 1301.55
R167 GNDA.n1400 GNDA.n1399 1285.24
R168 GNDA.n1552 GNDA.n1551 1242.27
R169 GNDA.n1900 GNDA.n1709 1214.72
R170 GNDA.n1900 GNDA.n1710 1214.72
R171 GNDA.n1858 GNDA.n1710 1214.72
R172 GNDA.n1866 GNDA.n1858 1214.72
R173 GNDA.n1866 GNDA.n1865 1214.72
R174 GNDA.n1881 GNDA.n1849 1214.72
R175 GNDA.n1881 GNDA.n1845 1214.72
R176 GNDA.n1888 GNDA.n1845 1214.72
R177 GNDA.n1888 GNDA.n410 1214.72
R178 GNDA.n2131 GNDA.n410 1214.72
R179 GNDA.n496 GNDA.n494 1164.49
R180 GNDA.n495 GNDA.n493 1114.8
R181 GNDA.n619 GNDA.n614 1114.8
R182 GNDA.n497 GNDA.t70 965.764
R183 GNDA.n1966 GNDA.n1965 949.682
R184 GNDA.n2497 GNDA.t238 949.682
R185 GNDA.n1393 GNDA.t229 875.452
R186 GNDA.n1849 GNDA.t229 823.313
R187 GNDA.n1542 GNDA.n1541 803.201
R188 GNDA.n1541 GNDA.n821 800
R189 GNDA.n1543 GNDA.n1542 774.4
R190 GNDA.n1543 GNDA.n821 771.201
R191 GNDA.n645 GNDA.t268 734.418
R192 GNDA.n643 GNDA.t258 734.418
R193 GNDA.n504 GNDA.t261 734.418
R194 GNDA.n800 GNDA.t252 734.418
R195 GNDA.n762 GNDA.n761 704
R196 GNDA.n762 GNDA.n521 697.601
R197 GNDA.n591 GNDA.t271 682.201
R198 GNDA.n2514 GNDA.n2513 669.307
R199 GNDA.n702 GNDA.t307 666.134
R200 GNDA.n566 GNDA.n563 624.324
R201 GNDA.n571 GNDA.n570 624.324
R202 GNDA.n1981 GNDA.n1966 623.755
R203 GNDA.n2491 GNDA.t238 623.755
R204 GNDA.n622 GNDA.n615 617.601
R205 GNDA.n499 GNDA.n492 617.601
R206 GNDA.n710 GNDA.n590 601.601
R207 GNDA.n768 GNDA.n767 598.4
R208 GNDA.n767 GNDA.n538 598.4
R209 GNDA.n1453 GNDA.n862 588.271
R210 GNDA.n1191 GNDA.n970 588.271
R211 GNDA.n2494 GNDA.n15 585
R212 GNDA.n205 GNDA.n14 585
R213 GNDA.n2372 GNDA.n2368 585
R214 GNDA.n2373 GNDA.n204 585
R215 GNDA.n2374 GNDA.n203 585
R216 GNDA.n2363 GNDA.n200 585
R217 GNDA.n2379 GNDA.n199 585
R218 GNDA.n2380 GNDA.n198 585
R219 GNDA.n2381 GNDA.n197 585
R220 GNDA.n2360 GNDA.n195 585
R221 GNDA.n2359 GNDA.n192 585
R222 GNDA.n2389 GNDA.n2388 585
R223 GNDA.n2392 GNDA.n2391 585
R224 GNDA.n2391 GNDA.n46 585
R225 GNDA.n2495 GNDA.n2494 585
R226 GNDA.n2370 GNDA.n14 585
R227 GNDA.n2372 GNDA.n2371 585
R228 GNDA.n2373 GNDA.n202 585
R229 GNDA.n2375 GNDA.n2374 585
R230 GNDA.n2377 GNDA.n200 585
R231 GNDA.n2379 GNDA.n2378 585
R232 GNDA.n2380 GNDA.n196 585
R233 GNDA.n2382 GNDA.n2381 585
R234 GNDA.n2384 GNDA.n195 585
R235 GNDA.n2385 GNDA.n192 585
R236 GNDA.n2388 GNDA.n2387 585
R237 GNDA.n2127 GNDA.n2126 585
R238 GNDA.n2014 GNDA.n2008 585
R239 GNDA.n2122 GNDA.n2121 585
R240 GNDA.n2016 GNDA.n2013 585
R241 GNDA.n2044 GNDA.n2043 585
R242 GNDA.n2048 GNDA.n2047 585
R243 GNDA.n2046 GNDA.n2037 585
R244 GNDA.n2055 GNDA.n2054 585
R245 GNDA.n2057 GNDA.n2056 585
R246 GNDA.n2062 GNDA.n2059 585
R247 GNDA.n2064 GNDA.n2063 585
R248 GNDA.n2060 GNDA.n193 585
R249 GNDA.n2324 GNDA.n69 585
R250 GNDA.n2318 GNDA.n364 585
R251 GNDA.n2320 GNDA.n2319 585
R252 GNDA.n2317 GNDA.n369 585
R253 GNDA.n2316 GNDA.n2315 585
R254 GNDA.n2314 GNDA.n2313 585
R255 GNDA.n2312 GNDA.n2311 585
R256 GNDA.n2310 GNDA.n2309 585
R257 GNDA.n2308 GNDA.n2307 585
R258 GNDA.n2306 GNDA.n2305 585
R259 GNDA.n2304 GNDA.n2303 585
R260 GNDA.n2302 GNDA.n2301 585
R261 GNDA.n2268 GNDA.n2267 585
R262 GNDA.n2265 GNDA.n388 585
R263 GNDA.n2158 GNDA.n2157 585
R264 GNDA.n2186 GNDA.n2185 585
R265 GNDA.n2188 GNDA.n2187 585
R266 GNDA.n2193 GNDA.n2192 585
R267 GNDA.n2195 GNDA.n2194 585
R268 GNDA.n2200 GNDA.n2199 585
R269 GNDA.n2202 GNDA.n2201 585
R270 GNDA.n2256 GNDA.n2204 585
R271 GNDA.n2258 GNDA.n2257 585
R272 GNDA.n2254 GNDA.n346 585
R273 GNDA.n2132 GNDA.n409 585
R274 GNDA.n2132 GNDA.n2131 585
R275 GNDA.n1885 GNDA.n408 585
R276 GNDA.n410 GNDA.n408 585
R277 GNDA.n1887 GNDA.n1886 585
R278 GNDA.n1888 GNDA.n1887 585
R279 GNDA.n1884 GNDA.n1846 585
R280 GNDA.n1846 GNDA.n1845 585
R281 GNDA.n1883 GNDA.n1882 585
R282 GNDA.n1882 GNDA.n1881 585
R283 GNDA.n1848 GNDA.n1847 585
R284 GNDA.n1849 GNDA.n1848 585
R285 GNDA.n1864 GNDA.n1863 585
R286 GNDA.n1865 GNDA.n1864 585
R287 GNDA.n1862 GNDA.n1859 585
R288 GNDA.n1866 GNDA.n1859 585
R289 GNDA.n1861 GNDA.n1860 585
R290 GNDA.n1860 GNDA.n1858 585
R291 GNDA.n1708 GNDA.n1707 585
R292 GNDA.n1710 GNDA.n1708 585
R293 GNDA.n1902 GNDA.n1901 585
R294 GNDA.n1901 GNDA.n1900 585
R295 GNDA.n1903 GNDA.n1706 585
R296 GNDA.n1709 GNDA.n1706 585
R297 GNDA.n1769 GNDA.n1711 585
R298 GNDA.n1711 GNDA.n1709 585
R299 GNDA.n1899 GNDA.n1898 585
R300 GNDA.n1900 GNDA.n1899 585
R301 GNDA.n1771 GNDA.n1712 585
R302 GNDA.n1712 GNDA.n1710 585
R303 GNDA.n1856 GNDA.n1855 585
R304 GNDA.n1858 GNDA.n1856 585
R305 GNDA.n1868 GNDA.n1867 585
R306 GNDA.n1867 GNDA.n1866 585
R307 GNDA.n1857 GNDA.n1851 585
R308 GNDA.n1865 GNDA.n1857 585
R309 GNDA.n1873 GNDA.n1850 585
R310 GNDA.n1850 GNDA.n1849 585
R311 GNDA.n1880 GNDA.n1879 585
R312 GNDA.n1881 GNDA.n1880 585
R313 GNDA.n1875 GNDA.n1844 585
R314 GNDA.n1845 GNDA.n1844 585
R315 GNDA.n1890 GNDA.n1889 585
R316 GNDA.n1889 GNDA.n1888 585
R317 GNDA.n1891 GNDA.n411 585
R318 GNDA.n411 GNDA.n410 585
R319 GNDA.n2130 GNDA.n2129 585
R320 GNDA.n2131 GNDA.n2130 585
R321 GNDA.n1154 GNDA.n969 585
R322 GNDA.n1152 GNDA.n1151 585
R323 GNDA.n973 GNDA.n971 585
R324 GNDA.n1054 GNDA.n1052 585
R325 GNDA.n1061 GNDA.n1060 585
R326 GNDA.n1063 GNDA.n1050 585
R327 GNDA.n1066 GNDA.n1065 585
R328 GNDA.n1048 GNDA.n1047 585
R329 GNDA.n1073 GNDA.n1072 585
R330 GNDA.n1075 GNDA.n995 585
R331 GNDA.n1144 GNDA.n1143 585
R332 GNDA.n1141 GNDA.n1140 585
R333 GNDA.n1703 GNDA.n1702 585
R334 GNDA.n1907 GNDA.n1703 585
R335 GNDA.n1910 GNDA.n1909 585
R336 GNDA.n1909 GNDA.n1908 585
R337 GNDA.n1911 GNDA.n1700 585
R338 GNDA.n1704 GNDA.n1700 585
R339 GNDA.n1913 GNDA.n1912 585
R340 GNDA.n1914 GNDA.n1913 585
R341 GNDA.n1701 GNDA.n1698 585
R342 GNDA.n1915 GNDA.n1698 585
R343 GNDA.n1918 GNDA.n1917 585
R344 GNDA.n1917 GNDA.n1916 585
R345 GNDA.n1919 GNDA.n1696 585
R346 GNDA.n1696 GNDA.n1695 585
R347 GNDA.n1921 GNDA.n1920 585
R348 GNDA.n1922 GNDA.n1921 585
R349 GNDA.n1697 GNDA.n1693 585
R350 GNDA.n1923 GNDA.n1693 585
R351 GNDA.n1925 GNDA.n1694 585
R352 GNDA.n1925 GNDA.n1924 585
R353 GNDA.n1926 GNDA.n1568 585
R354 GNDA.n1929 GNDA.n1928 585
R355 GNDA.n1691 GNDA.n1690 585
R356 GNDA.n1690 GNDA.n1567 585
R357 GNDA.n1905 GNDA.n1904 585
R358 GNDA.n1906 GNDA.n1905 585
R359 GNDA.n1727 GNDA.n1726 585
R360 GNDA.n1727 GNDA.n465 585
R361 GNDA.n1746 GNDA.n1745 585
R362 GNDA.n1745 GNDA.n1744 585
R363 GNDA.n1747 GNDA.n1724 585
R364 GNDA.n1724 GNDA.n1723 585
R365 GNDA.n1749 GNDA.n1748 585
R366 GNDA.n1750 GNDA.n1749 585
R367 GNDA.n1725 GNDA.n1722 585
R368 GNDA.n1751 GNDA.n1722 585
R369 GNDA.n1754 GNDA.n1753 585
R370 GNDA.n1753 GNDA.n1752 585
R371 GNDA.n1755 GNDA.n1720 585
R372 GNDA.n1720 GNDA.n1719 585
R373 GNDA.n1757 GNDA.n1756 585
R374 GNDA.n1758 GNDA.n1757 585
R375 GNDA.n1721 GNDA.n1716 585
R376 GNDA.n1759 GNDA.n1716 585
R377 GNDA.n1761 GNDA.n1717 585
R378 GNDA.n1761 GNDA.n1760 585
R379 GNDA.n1762 GNDA.n1715 585
R380 GNDA.n1765 GNDA.n1764 585
R381 GNDA.n1768 GNDA.n1767 585
R382 GNDA.n1767 GNDA.n1766 585
R383 GNDA.n2133 GNDA.n371 585
R384 GNDA.n425 GNDA.n406 585
R385 GNDA.n2138 GNDA.n405 585
R386 GNDA.n2139 GNDA.n404 585
R387 GNDA.n2140 GNDA.n403 585
R388 GNDA.n422 GNDA.n400 585
R389 GNDA.n2145 GNDA.n399 585
R390 GNDA.n2146 GNDA.n398 585
R391 GNDA.n2147 GNDA.n397 585
R392 GNDA.n419 GNDA.n395 585
R393 GNDA.n418 GNDA.n392 585
R394 GNDA.n2154 GNDA.n391 585
R395 GNDA.n380 GNDA.n374 585
R396 GNDA.n2299 GNDA.n374 585
R397 GNDA.n2300 GNDA.n372 585
R398 GNDA.n2300 GNDA.n2299 585
R399 GNDA.n1984 GNDA.n451 585
R400 GNDA.n449 GNDA.n446 585
R401 GNDA.n1989 GNDA.n445 585
R402 GNDA.n1990 GNDA.n443 585
R403 GNDA.n1991 GNDA.n442 585
R404 GNDA.n440 GNDA.n437 585
R405 GNDA.n1996 GNDA.n436 585
R406 GNDA.n1997 GNDA.n434 585
R407 GNDA.n1998 GNDA.n433 585
R408 GNDA.n429 GNDA.n428 585
R409 GNDA.n2004 GNDA.n2003 585
R410 GNDA.n2006 GNDA.n415 585
R411 GNDA.n414 GNDA.n373 585
R412 GNDA.n2299 GNDA.n373 585
R413 GNDA.n2134 GNDA.n2133 585
R414 GNDA.n2136 GNDA.n406 585
R415 GNDA.n2138 GNDA.n2137 585
R416 GNDA.n2139 GNDA.n402 585
R417 GNDA.n2141 GNDA.n2140 585
R418 GNDA.n2143 GNDA.n400 585
R419 GNDA.n2145 GNDA.n2144 585
R420 GNDA.n2146 GNDA.n396 585
R421 GNDA.n2148 GNDA.n2147 585
R422 GNDA.n2150 GNDA.n395 585
R423 GNDA.n2151 GNDA.n392 585
R424 GNDA.n2154 GNDA.n2153 585
R425 GNDA.n1985 GNDA.n1984 585
R426 GNDA.n1987 GNDA.n446 585
R427 GNDA.n1989 GNDA.n1988 585
R428 GNDA.n1990 GNDA.n439 585
R429 GNDA.n1992 GNDA.n1991 585
R430 GNDA.n1994 GNDA.n437 585
R431 GNDA.n1996 GNDA.n1995 585
R432 GNDA.n1997 GNDA.n431 585
R433 GNDA.n1999 GNDA.n1998 585
R434 GNDA.n2001 GNDA.n429 585
R435 GNDA.n2003 GNDA.n2002 585
R436 GNDA.n415 GNDA.n412 585
R437 GNDA.n1689 GNDA.n1688 585
R438 GNDA.n1577 GNDA.n1571 585
R439 GNDA.n1684 GNDA.n1683 585
R440 GNDA.n1579 GNDA.n1576 585
R441 GNDA.n1607 GNDA.n1606 585
R442 GNDA.n1611 GNDA.n1610 585
R443 GNDA.n1609 GNDA.n1600 585
R444 GNDA.n1618 GNDA.n1617 585
R445 GNDA.n1620 GNDA.n1619 585
R446 GNDA.n1624 GNDA.n1622 585
R447 GNDA.n1626 GNDA.n1625 585
R448 GNDA.n393 GNDA.n390 585
R449 GNDA.n1432 GNDA.n379 585
R450 GNDA.n1426 GNDA.n1233 585
R451 GNDA.n1428 GNDA.n1427 585
R452 GNDA.n1425 GNDA.n1238 585
R453 GNDA.n1424 GNDA.n1423 585
R454 GNDA.n1422 GNDA.n1421 585
R455 GNDA.n1420 GNDA.n1419 585
R456 GNDA.n1418 GNDA.n1417 585
R457 GNDA.n1416 GNDA.n1415 585
R458 GNDA.n1414 GNDA.n1413 585
R459 GNDA.n1412 GNDA.n1411 585
R460 GNDA.n1410 GNDA.n1409 585
R461 GNDA.n1252 GNDA.n1240 585
R462 GNDA.n1241 GNDA.n1240 585
R463 GNDA.n1254 GNDA.n1253 585
R464 GNDA.n1255 GNDA.n1254 585
R465 GNDA.n1258 GNDA.n1257 585
R466 GNDA.n1257 GNDA.n1256 585
R467 GNDA.n1259 GNDA.n1251 585
R468 GNDA.n1251 GNDA.n1250 585
R469 GNDA.n1261 GNDA.n1260 585
R470 GNDA.n1262 GNDA.n1261 585
R471 GNDA.n1249 GNDA.n1248 585
R472 GNDA.n1263 GNDA.n1249 585
R473 GNDA.n1266 GNDA.n1265 585
R474 GNDA.n1265 GNDA.n1264 585
R475 GNDA.n1267 GNDA.n1247 585
R476 GNDA.n1247 GNDA.n476 585
R477 GNDA.n1269 GNDA.n1268 585
R478 GNDA.n1269 GNDA.n474 585
R479 GNDA.n1270 GNDA.n1245 585
R480 GNDA.n1271 GNDA.n1270 585
R481 GNDA.n1408 GNDA.n1239 585
R482 GNDA.n1408 GNDA.n1407 585
R483 GNDA.n1273 GNDA.n1272 585
R484 GNDA.n1246 GNDA.n1243 585
R485 GNDA.n1398 GNDA.n1397 585
R486 GNDA.n1399 GNDA.n1398 585
R487 GNDA.n1396 GNDA.n1395 585
R488 GNDA.n1280 GNDA.n1277 585
R489 GNDA.n1391 GNDA.n1390 585
R490 GNDA.n1282 GNDA.n1279 585
R491 GNDA.n1313 GNDA.n1312 585
R492 GNDA.n1314 GNDA.n1313 585
R493 GNDA.n1317 GNDA.n1316 585
R494 GNDA.n1316 GNDA.n1315 585
R495 GNDA.n1318 GNDA.n1305 585
R496 GNDA.n1305 GNDA.n1304 585
R497 GNDA.n1327 GNDA.n1326 585
R498 GNDA.n1328 GNDA.n1327 585
R499 GNDA.n1307 GNDA.n1303 585
R500 GNDA.n1329 GNDA.n1303 585
R501 GNDA.n1332 GNDA.n1331 585
R502 GNDA.n1331 GNDA.n1330 585
R503 GNDA.n1333 GNDA.n858 585
R504 GNDA.n858 GNDA.n857 585
R505 GNDA.n1455 GNDA.n1454 585
R506 GNDA.n1456 GNDA.n1455 585
R507 GNDA.n1206 GNDA.n861 585
R508 GNDA.n1204 GNDA.n1203 585
R509 GNDA.n865 GNDA.n863 585
R510 GNDA.n946 GNDA.n944 585
R511 GNDA.n953 GNDA.n952 585
R512 GNDA.n955 GNDA.n942 585
R513 GNDA.n958 GNDA.n957 585
R514 GNDA.n940 GNDA.n939 585
R515 GNDA.n965 GNDA.n964 585
R516 GNDA.n967 GNDA.n887 585
R517 GNDA.n1196 GNDA.n1195 585
R518 GNDA.n1193 GNDA.n1192 585
R519 GNDA.n378 GNDA.n376 585
R520 GNDA.n1231 GNDA.n1230 585
R521 GNDA.n1437 GNDA.n1228 585
R522 GNDA.n1438 GNDA.n1226 585
R523 GNDA.n1439 GNDA.n1225 585
R524 GNDA.n1223 GNDA.n1220 585
R525 GNDA.n1444 GNDA.n1219 585
R526 GNDA.n1445 GNDA.n1217 585
R527 GNDA.n1446 GNDA.n1216 585
R528 GNDA.n1214 GNDA.n1211 585
R529 GNDA.n1451 GNDA.n1210 585
R530 GNDA.n1452 GNDA.n1208 585
R531 GNDA.n862 GNDA.n856 585
R532 GNDA.n2298 GNDA.n2297 585
R533 GNDA.n2299 GNDA.n2298 585
R534 GNDA.n1433 GNDA.n378 585
R535 GNDA.n1435 GNDA.n1231 585
R536 GNDA.n1437 GNDA.n1436 585
R537 GNDA.n1438 GNDA.n1222 585
R538 GNDA.n1440 GNDA.n1439 585
R539 GNDA.n1442 GNDA.n1220 585
R540 GNDA.n1444 GNDA.n1443 585
R541 GNDA.n1445 GNDA.n1213 585
R542 GNDA.n1447 GNDA.n1446 585
R543 GNDA.n1449 GNDA.n1211 585
R544 GNDA.n1451 GNDA.n1450 585
R545 GNDA.n1452 GNDA.n859 585
R546 GNDA.n2354 GNDA.n2353 585
R547 GNDA.n2278 GNDA.n223 585
R548 GNDA.n2280 GNDA.n2279 585
R549 GNDA.n2281 GNDA.n2276 585
R550 GNDA.n2283 GNDA.n2282 585
R551 GNDA.n2285 GNDA.n2274 585
R552 GNDA.n2287 GNDA.n2286 585
R553 GNDA.n2288 GNDA.n2273 585
R554 GNDA.n2290 GNDA.n2289 585
R555 GNDA.n2292 GNDA.n381 585
R556 GNDA.n2294 GNDA.n2293 585
R557 GNDA.n2295 GNDA.n377 585
R558 GNDA.n1116 GNDA.n1088 585
R559 GNDA.n1114 GNDA.n1113 585
R560 GNDA.n1112 GNDA.n1089 585
R561 GNDA.n1111 GNDA.n1110 585
R562 GNDA.n1108 GNDA.n1090 585
R563 GNDA.n1106 GNDA.n1105 585
R564 GNDA.n1104 GNDA.n1091 585
R565 GNDA.n1103 GNDA.n1102 585
R566 GNDA.n1100 GNDA.n1092 585
R567 GNDA.n1098 GNDA.n1097 585
R568 GNDA.n1096 GNDA.n1095 585
R569 GNDA.n1093 GNDA.n224 585
R570 GNDA.n2357 GNDA.n2356 585
R571 GNDA.n219 GNDA.n217 585
R572 GNDA.n1175 GNDA.n1171 585
R573 GNDA.n1176 GNDA.n1170 585
R574 GNDA.n1177 GNDA.n1169 585
R575 GNDA.n1166 GNDA.n1165 585
R576 GNDA.n1182 GNDA.n1164 585
R577 GNDA.n1183 GNDA.n1163 585
R578 GNDA.n1184 GNDA.n1162 585
R579 GNDA.n1159 GNDA.n1158 585
R580 GNDA.n1189 GNDA.n1157 585
R581 GNDA.n1190 GNDA.n1156 585
R582 GNDA.n970 GNDA.n856 585
R583 GNDA.n220 GNDA.n218 585
R584 GNDA.n218 GNDA.n46 585
R585 GNDA.n2356 GNDA.n2355 585
R586 GNDA.n1173 GNDA.n219 585
R587 GNDA.n1175 GNDA.n1174 585
R588 GNDA.n1176 GNDA.n1168 585
R589 GNDA.n1178 GNDA.n1177 585
R590 GNDA.n1180 GNDA.n1166 585
R591 GNDA.n1182 GNDA.n1181 585
R592 GNDA.n1183 GNDA.n1161 585
R593 GNDA.n1185 GNDA.n1184 585
R594 GNDA.n1187 GNDA.n1159 585
R595 GNDA.n1189 GNDA.n1188 585
R596 GNDA.n1190 GNDA.n968 585
R597 GNDA.n2326 GNDA.n2325 585
R598 GNDA.n362 GNDA.n361 585
R599 GNDA.n2331 GNDA.n360 585
R600 GNDA.n2332 GNDA.n359 585
R601 GNDA.n2333 GNDA.n358 585
R602 GNDA.n355 GNDA.n354 585
R603 GNDA.n2338 GNDA.n353 585
R604 GNDA.n2339 GNDA.n352 585
R605 GNDA.n2340 GNDA.n351 585
R606 GNDA.n349 GNDA.n348 585
R607 GNDA.n347 GNDA.n345 585
R608 GNDA.n2348 GNDA.n2347 585
R609 GNDA.n2351 GNDA.n2350 585
R610 GNDA.n2350 GNDA.n46 585
R611 GNDA.n70 GNDA.n68 585
R612 GNDA.n68 GNDA.n46 585
R613 GNDA.n2327 GNDA.n2326 585
R614 GNDA.n2329 GNDA.n362 585
R615 GNDA.n2331 GNDA.n2330 585
R616 GNDA.n2332 GNDA.n357 585
R617 GNDA.n2334 GNDA.n2333 585
R618 GNDA.n2336 GNDA.n355 585
R619 GNDA.n2338 GNDA.n2337 585
R620 GNDA.n2339 GNDA.n350 585
R621 GNDA.n2341 GNDA.n2340 585
R622 GNDA.n2343 GNDA.n349 585
R623 GNDA.n2344 GNDA.n345 585
R624 GNDA.n2347 GNDA.n2346 585
R625 GNDA.n344 GNDA.n343 585
R626 GNDA.n341 GNDA.n340 585
R627 GNDA.n339 GNDA.n338 585
R628 GNDA.n257 GNDA.n230 585
R629 GNDA.n261 GNDA.n260 585
R630 GNDA.n263 GNDA.n256 585
R631 GNDA.n266 GNDA.n265 585
R632 GNDA.n252 GNDA.n251 585
R633 GNDA.n276 GNDA.n275 585
R634 GNDA.n278 GNDA.n249 585
R635 GNDA.n281 GNDA.n280 585
R636 GNDA.n52 GNDA.n50 585
R637 GNDA.n2417 GNDA.n2416 585
R638 GNDA.n2415 GNDA.n2414 585
R639 GNDA.n2413 GNDA.n63 585
R640 GNDA.n2411 GNDA.n2410 585
R641 GNDA.n2409 GNDA.n64 585
R642 GNDA.n2408 GNDA.n2407 585
R643 GNDA.n2405 GNDA.n65 585
R644 GNDA.n2403 GNDA.n2402 585
R645 GNDA.n2401 GNDA.n66 585
R646 GNDA.n2400 GNDA.n2399 585
R647 GNDA.n2397 GNDA.n67 585
R648 GNDA.n2395 GNDA.n2394 585
R649 GNDA.n190 GNDA.n189 585
R650 GNDA.n187 GNDA.n186 585
R651 GNDA.n185 GNDA.n184 585
R652 GNDA.n103 GNDA.n76 585
R653 GNDA.n107 GNDA.n106 585
R654 GNDA.n109 GNDA.n102 585
R655 GNDA.n112 GNDA.n111 585
R656 GNDA.n98 GNDA.n97 585
R657 GNDA.n122 GNDA.n121 585
R658 GNDA.n124 GNDA.n95 585
R659 GNDA.n127 GNDA.n126 585
R660 GNDA.n41 GNDA.n40 585
R661 GNDA.n1117 GNDA.n1087 585
R662 GNDA.n1117 GNDA.n48 585
R663 GNDA.n1120 GNDA.n1119 585
R664 GNDA.n1119 GNDA.n1118 585
R665 GNDA.n1121 GNDA.n1085 585
R666 GNDA.n1085 GNDA.n1084 585
R667 GNDA.n1123 GNDA.n1122 585
R668 GNDA.n1124 GNDA.n1123 585
R669 GNDA.n1086 GNDA.n1083 585
R670 GNDA.n1125 GNDA.n1083 585
R671 GNDA.n1127 GNDA.n1082 585
R672 GNDA.n1127 GNDA.n1126 585
R673 GNDA.n1130 GNDA.n1129 585
R674 GNDA.n1129 GNDA.n1128 585
R675 GNDA.n1131 GNDA.n1081 585
R676 GNDA.n1081 GNDA.n1080 585
R677 GNDA.n1133 GNDA.n1132 585
R678 GNDA.n1134 GNDA.n1133 585
R679 GNDA.n1078 GNDA.n1077 585
R680 GNDA.n1135 GNDA.n1078 585
R681 GNDA.n1137 GNDA.n1136 585
R682 GNDA.n1079 GNDA.n1076 585
R683 GNDA.n2418 GNDA.n61 585
R684 GNDA.n2418 GNDA.n43 585
R685 GNDA.n2421 GNDA.n2420 585
R686 GNDA.n2420 GNDA.n2419 585
R687 GNDA.n2422 GNDA.n60 585
R688 GNDA.n60 GNDA.n59 585
R689 GNDA.n2424 GNDA.n2423 585
R690 GNDA.n2425 GNDA.n2424 585
R691 GNDA.n58 GNDA.n57 585
R692 GNDA.n2426 GNDA.n58 585
R693 GNDA.n2429 GNDA.n2428 585
R694 GNDA.n2428 GNDA.n2427 585
R695 GNDA.n2430 GNDA.n56 585
R696 GNDA.n56 GNDA.n55 585
R697 GNDA.n2432 GNDA.n2431 585
R698 GNDA.n2433 GNDA.n2432 585
R699 GNDA.n54 GNDA.n53 585
R700 GNDA.n2434 GNDA.n54 585
R701 GNDA.n2437 GNDA.n2436 585
R702 GNDA.n2436 GNDA.n2435 585
R703 GNDA.n51 GNDA.n49 585
R704 GNDA.n2441 GNDA.n2440 585
R705 GNDA.n30 GNDA.n29 585
R706 GNDA.n2466 GNDA.n30 585
R707 GNDA.n2464 GNDA.n2463 585
R708 GNDA.n2465 GNDA.n2464 585
R709 GNDA.n2462 GNDA.n32 585
R710 GNDA.n32 GNDA.n31 585
R711 GNDA.n2461 GNDA.n2460 585
R712 GNDA.n2460 GNDA.n2459 585
R713 GNDA.n34 GNDA.n33 585
R714 GNDA.n2458 GNDA.n34 585
R715 GNDA.n2456 GNDA.n2455 585
R716 GNDA.n2457 GNDA.n2456 585
R717 GNDA.n2454 GNDA.n35 585
R718 GNDA.n2450 GNDA.n35 585
R719 GNDA.n2453 GNDA.n2452 585
R720 GNDA.n2452 GNDA.n2451 585
R721 GNDA.n37 GNDA.n36 585
R722 GNDA.n2449 GNDA.n37 585
R723 GNDA.n2447 GNDA.n2446 585
R724 GNDA.n2448 GNDA.n2447 585
R725 GNDA.n39 GNDA.n38 585
R726 GNDA.n2443 GNDA.n2442 585
R727 GNDA.n2493 GNDA.n2492 585
R728 GNDA.n2492 GNDA.n2491 585
R729 GNDA.n2469 GNDA.n2468 585
R730 GNDA.n2468 GNDA.n2467 585
R731 GNDA.n2470 GNDA.n28 585
R732 GNDA.n28 GNDA.n27 585
R733 GNDA.n2472 GNDA.n2471 585
R734 GNDA.n2473 GNDA.n2472 585
R735 GNDA.n25 GNDA.n24 585
R736 GNDA.n2474 GNDA.n25 585
R737 GNDA.n2477 GNDA.n2476 585
R738 GNDA.n2476 GNDA.n2475 585
R739 GNDA.n2478 GNDA.n23 585
R740 GNDA.n26 GNDA.n23 585
R741 GNDA.n2480 GNDA.n2479 585
R742 GNDA.n2481 GNDA.n2480 585
R743 GNDA.n22 GNDA.n21 585
R744 GNDA.n2482 GNDA.n22 585
R745 GNDA.n2485 GNDA.n2484 585
R746 GNDA.n2484 GNDA.n2483 585
R747 GNDA.n2486 GNDA.n19 585
R748 GNDA.n19 GNDA.n18 585
R749 GNDA.n2488 GNDA.n2487 585
R750 GNDA.n2489 GNDA.n2488 585
R751 GNDA.n20 GNDA.n17 585
R752 GNDA.n2490 GNDA.n17 585
R753 GNDA.n4 GNDA.n3 585
R754 GNDA.n2511 GNDA.n2510 585
R755 GNDA.n2512 GNDA.n2511 585
R756 GNDA.n1983 GNDA.n1982 585
R757 GNDA.n1982 GNDA.n1981 585
R758 GNDA.n2496 GNDA.n12 585
R759 GNDA.n2497 GNDA.n2496 585
R760 GNDA.n2500 GNDA.n2499 585
R761 GNDA.n2499 GNDA.n2498 585
R762 GNDA.n2501 GNDA.n11 585
R763 GNDA.n11 GNDA.n10 585
R764 GNDA.n2503 GNDA.n2502 585
R765 GNDA.n2504 GNDA.n2503 585
R766 GNDA.n9 GNDA.n7 585
R767 GNDA.n2505 GNDA.n9 585
R768 GNDA.n2508 GNDA.n2507 585
R769 GNDA.n2507 GNDA.n2506 585
R770 GNDA.n8 GNDA.n6 585
R771 GNDA.n8 GNDA.n5 585
R772 GNDA.n1971 GNDA.n1970 585
R773 GNDA.n1972 GNDA.n1971 585
R774 GNDA.n1975 GNDA.n1974 585
R775 GNDA.n1974 GNDA.n1973 585
R776 GNDA.n1976 GNDA.n1968 585
R777 GNDA.n1968 GNDA.n1967 585
R778 GNDA.n1978 GNDA.n1977 585
R779 GNDA.n1979 GNDA.n1978 585
R780 GNDA.n1969 GNDA.n453 585
R781 GNDA.n1980 GNDA.n453 585
R782 GNDA.n464 GNDA.n463 585
R783 GNDA.n1939 GNDA.n464 585
R784 GNDA.n1961 GNDA.n448 585
R785 GNDA.n1965 GNDA.n448 585
R786 GNDA.n1963 GNDA.n1962 585
R787 GNDA.n1964 GNDA.n1963 585
R788 GNDA.n1960 GNDA.n455 585
R789 GNDA.n455 GNDA.n454 585
R790 GNDA.n1959 GNDA.n1958 585
R791 GNDA.n1958 GNDA.n1957 585
R792 GNDA.n457 GNDA.n456 585
R793 GNDA.n1956 GNDA.n457 585
R794 GNDA.n1954 GNDA.n1953 585
R795 GNDA.n1955 GNDA.n1954 585
R796 GNDA.n1952 GNDA.n458 585
R797 GNDA.n1948 GNDA.n458 585
R798 GNDA.n1951 GNDA.n1950 585
R799 GNDA.n1950 GNDA.n1949 585
R800 GNDA.n460 GNDA.n459 585
R801 GNDA.n1947 GNDA.n460 585
R802 GNDA.n1945 GNDA.n1944 585
R803 GNDA.n1946 GNDA.n1945 585
R804 GNDA.n1943 GNDA.n462 585
R805 GNDA.n462 GNDA.n461 585
R806 GNDA.n1942 GNDA.n1941 585
R807 GNDA.n1941 GNDA.n1940 585
R808 GNDA.n597 GNDA.t301 535.191
R809 GNDA.n513 GNDA.t242 535.191
R810 GNDA.n516 GNDA.t230 535.191
R811 GNDA.n652 GNDA.t289 535.191
R812 GNDA.n1563 GNDA.n1562 531.201
R813 GNDA.n706 GNDA.n590 531.201
R814 GNDA.n1564 GNDA.n1563 528
R815 GNDA.n1709 GNDA.n1705 512.884
R816 GNDA.n1537 GNDA.n851 512
R817 GNDA.n1537 GNDA.n1536 512
R818 GNDA.n1492 GNDA.n1487 512
R819 GNDA.n1492 GNDA.n1489 512
R820 GNDA.n853 GNDA.n851 508.8
R821 GNDA.n1536 GNDA.n853 508.8
R822 GNDA.n1488 GNDA.n1487 508.8
R823 GNDA.n1489 GNDA.n1488 508.8
R824 GNDA.n1940 GNDA.n1939 505.748
R825 GNDA.n1940 GNDA.n461 505.748
R826 GNDA.n1946 GNDA.n461 505.748
R827 GNDA.n1947 GNDA.n1946 505.748
R828 GNDA.n1949 GNDA.n1947 505.748
R829 GNDA.n1949 GNDA.n1948 505.748
R830 GNDA.n1956 GNDA.n1955 505.748
R831 GNDA.n1957 GNDA.n1956 505.748
R832 GNDA.n1957 GNDA.n454 505.748
R833 GNDA.n1964 GNDA.n454 505.748
R834 GNDA.n1965 GNDA.n1964 505.748
R835 GNDA.n1981 GNDA.n1980 505.748
R836 GNDA.n1980 GNDA.n1979 505.748
R837 GNDA.n1979 GNDA.n1967 505.748
R838 GNDA.n1973 GNDA.n1967 505.748
R839 GNDA.n1973 GNDA.n1972 505.748
R840 GNDA.n1972 GNDA.n5 505.748
R841 GNDA.n2506 GNDA.n2505 505.748
R842 GNDA.n2505 GNDA.n2504 505.748
R843 GNDA.n2504 GNDA.n10 505.748
R844 GNDA.n2498 GNDA.n10 505.748
R845 GNDA.n2498 GNDA.n2497 505.748
R846 GNDA.n2491 GNDA.n2490 505.748
R847 GNDA.n2490 GNDA.n2489 505.748
R848 GNDA.n2489 GNDA.n18 505.748
R849 GNDA.n2483 GNDA.n18 505.748
R850 GNDA.n2483 GNDA.n2482 505.748
R851 GNDA.n2482 GNDA.n2481 505.748
R852 GNDA.n2475 GNDA.n26 505.748
R853 GNDA.n2475 GNDA.n2474 505.748
R854 GNDA.n2474 GNDA.n2473 505.748
R855 GNDA.n2473 GNDA.n27 505.748
R856 GNDA.n2467 GNDA.n27 505.748
R857 GNDA.n1562 GNDA.n481 499.2
R858 GNDA.n796 GNDA.n519 496
R859 GNDA.n658 GNDA.n594 496
R860 GNDA.n529 GNDA.t321 493.418
R861 GNDA.n533 GNDA.t298 493.418
R862 GNDA.n532 GNDA.t316 493.418
R863 GNDA.n531 GNDA.t292 493.418
R864 GNDA.n543 GNDA.t324 493.418
R865 GNDA.n542 GNDA.t304 493.418
R866 GNDA.n541 GNDA.t285 493.418
R867 GNDA.n539 GNDA.t247 493.418
R868 GNDA.n758 GNDA.t234 493.418
R869 GNDA.n757 GNDA.t310 493.418
R870 GNDA.n797 GNDA.n796 489.601
R871 GNDA.n658 GNDA.n593 489.601
R872 GNDA.n1564 GNDA.n472 486.401
R873 GNDA.n1400 GNDA.n1242 467.039
R874 GNDA.n812 GNDA.n488 466.103
R875 GNDA.n1554 GNDA.n486 444.8
R876 GNDA.n1555 GNDA.n1554 444.8
R877 GNDA.n1498 GNDA.n1497 444.695
R878 GNDA.n1557 GNDA.n486 441.601
R879 GNDA.n560 GNDA.t239 441.2
R880 GNDA.n1556 GNDA.n1555 438.401
R881 GNDA.n1935 GNDA.n469 435.2
R882 GNDA.n709 GNDA.n708 428.8
R883 GNDA.n1935 GNDA.n1934 425.601
R884 GNDA.n561 GNDA.t249 425.134
R885 GNDA.n537 GNDA.n536 422.401
R886 GNDA.n534 GNDA.n530 422.401
R887 GNDA.n545 GNDA.n544 422.401
R888 GNDA.n760 GNDA.n759 422.401
R889 GNDA.n1933 GNDA.n471 422.401
R890 GNDA.n1934 GNDA.n1933 419.2
R891 GNDA.n1533 GNDA.n1458 408.661
R892 GNDA.n1506 GNDA.n1465 406.401
R893 GNDA.n1526 GNDA.n1465 406.401
R894 GNDA.n1865 GNDA.t229 391.411
R895 GNDA.n650 GNDA.n600 387.2
R896 GNDA.n805 GNDA.n507 387.2
R897 GNDA.n650 GNDA.n599 380.8
R898 GNDA.n806 GNDA.n805 380.8
R899 GNDA.n1498 GNDA.n1475 377.149
R900 GNDA.n708 GNDA.n707 355.2
R901 GNDA.n1399 GNDA.n1243 354.67
R902 GNDA.n1766 GNDA.n1765 354.67
R903 GNDA.n1315 GNDA.n1314 352.627
R904 GNDA.n1328 GNDA.n1304 352.627
R905 GNDA.n1329 GNDA.n1328 352.627
R906 GNDA.n1330 GNDA.n1329 352.627
R907 GNDA.n1330 GNDA.n857 352.627
R908 GNDA.n1456 GNDA.n857 352.627
R909 GNDA.n1527 GNDA.n1461 348.8
R910 GNDA.n1531 GNDA.n1461 348.8
R911 GNDA.n1480 GNDA.n1469 348.8
R912 GNDA.n1505 GNDA.n1469 348.8
R913 GNDA.n631 GNDA.n611 346.88
R914 GNDA.n503 GNDA.n502 346.88
R915 GNDA.n1955 GNDA.t229 342.784
R916 GNDA.n2506 GNDA.t238 342.784
R917 GNDA.n26 GNDA.t238 342.784
R918 GNDA.n629 GNDA.n628 342.401
R919 GNDA.n809 GNDA.n808 342.401
R920 GNDA.n1407 GNDA.n1241 337.111
R921 GNDA.n1907 GNDA.n1906 337.111
R922 GNDA.n636 GNDA.n607 332.8
R923 GNDA.n581 GNDA.n574 332.8
R924 GNDA.n552 GNDA.t265 332.75
R925 GNDA.n554 GNDA.t255 332.75
R926 GNDA.t238 GNDA.n47 172.876
R927 GNDA.n44 GNDA.t238 172.876
R928 GNDA.n42 GNDA.t238 172.615
R929 GNDA.t238 GNDA.n45 172.615
R930 GNDA.n1520 GNDA.n1519 323.2
R931 GNDA.n638 GNDA.n637 321.281
R932 GNDA.n583 GNDA.n582 321.281
R933 GNDA.n637 GNDA.n636 318.08
R934 GNDA.n582 GNDA.n581 318.08
R935 GNDA.n628 GNDA.n612 318.08
R936 GNDA.n809 GNDA.n501 318.08
R937 GNDA.n1520 GNDA.n1517 316.8
R938 GNDA.n1272 GNDA.n1243 316.043
R939 GNDA.n1272 GNDA.n1271 316.043
R940 GNDA.n1271 GNDA.n474 316.043
R941 GNDA.n1264 GNDA.n476 316.043
R942 GNDA.n1263 GNDA.n1262 316.043
R943 GNDA.n1262 GNDA.n1250 316.043
R944 GNDA.n1256 GNDA.n1250 316.043
R945 GNDA.n1256 GNDA.n1255 316.043
R946 GNDA.n1255 GNDA.n1241 316.043
R947 GNDA.n1929 GNDA.n1568 316.043
R948 GNDA.n1924 GNDA.n1568 316.043
R949 GNDA.n1924 GNDA.n1923 316.043
R950 GNDA.n1923 GNDA.n1922 316.043
R951 GNDA.n1922 GNDA.n1695 316.043
R952 GNDA.n1916 GNDA.n1915 316.043
R953 GNDA.n1915 GNDA.n1914 316.043
R954 GNDA.n1908 GNDA.n1704 316.043
R955 GNDA.n1908 GNDA.n1907 316.043
R956 GNDA.n1765 GNDA.n1715 316.043
R957 GNDA.n1760 GNDA.n1759 316.043
R958 GNDA.n1759 GNDA.n1758 316.043
R959 GNDA.n1758 GNDA.n1719 316.043
R960 GNDA.n1752 GNDA.n1751 316.043
R961 GNDA.n1751 GNDA.n1750 316.043
R962 GNDA.n1750 GNDA.n1723 316.043
R963 GNDA.n1744 GNDA.n1723 316.043
R964 GNDA.n519 GNDA.n518 310.401
R965 GNDA.n653 GNDA.n594 310.401
R966 GNDA.n1906 GNDA.n1705 305.507
R967 GNDA.n1402 GNDA.n480 304
R968 GNDA.n797 GNDA.n514 304
R969 GNDA.n598 GNDA.n593 304
R970 GNDA.n1458 GNDA.n856 303.363
R971 GNDA.n1567 GNDA.t229 301.995
R972 GNDA.n1766 GNDA.n1705 301.995
R973 GNDA.n1404 GNDA.n480 300.8
R974 GNDA.n1403 GNDA.n1402 300.8
R975 GNDA.n607 GNDA.n606 300.8
R976 GNDA.n754 GNDA.n753 300.8
R977 GNDA.n753 GNDA.n742 300.8
R978 GNDA.n574 GNDA.n515 300.8
R979 GNDA.n1404 GNDA.n1403 297.601
R980 GNDA.n1732 GNDA.n470 297.601
R981 GNDA.n1740 GNDA.n1732 297.601
R982 GNDA.n1739 GNDA.n1733 297.601
R983 GNDA.n1735 GNDA.n1733 297.601
R984 GNDA.n620 GNDA.n615 296
R985 GNDA.n492 GNDA.n491 296
R986 GNDA.n1519 GNDA.n1518 294.401
R987 GNDA.n1467 GNDA.t282 292.584
R988 GNDA.n1466 GNDA.t275 292.584
R989 GNDA.n1462 GNDA.t313 292.584
R990 GNDA.n1463 GNDA.t295 292.584
R991 GNDA.n1477 GNDA.t225 292.584
R992 GNDA.n1470 GNDA.t278 292.584
R993 GNDA.n481 GNDA.n479 292.5
R994 GNDA.n479 GNDA.n473 292.5
R995 GNDA.n1563 GNDA.n478 292.5
R996 GNDA.n478 GNDA.n473 292.5
R997 GNDA.n1562 GNDA.n1561 292.5
R998 GNDA.n1561 GNDA.n1560 292.5
R999 GNDA.n1558 GNDA.n1557 292.5
R1000 GNDA.n1559 GNDA.n1558 292.5
R1001 GNDA.n486 GNDA.n484 292.5
R1002 GNDA.n484 GNDA.n482 292.5
R1003 GNDA.n1554 GNDA.n1553 292.5
R1004 GNDA.n1553 GNDA.n1552 292.5
R1005 GNDA.n526 GNDA.n524 292.5
R1006 GNDA.n771 GNDA.n526 292.5
R1007 GNDA.n775 GNDA.n774 292.5
R1008 GNDA.n774 GNDA.t162 292.5
R1009 GNDA.n525 GNDA.n523 292.5
R1010 GNDA.n587 GNDA.n525 292.5
R1011 GNDA.n773 GNDA.n772 292.5
R1012 GNDA.t162 GNDA.n773 292.5
R1013 GNDA.n738 GNDA.n737 292.5
R1014 GNDA.n739 GNDA.n738 292.5
R1015 GNDA.n735 GNDA.n558 292.5
R1016 GNDA.n728 GNDA.n558 292.5
R1017 GNDA.n733 GNDA.n732 292.5
R1018 GNDA.n732 GNDA.n731 292.5
R1019 GNDA.n559 GNDA.n557 292.5
R1020 GNDA.n728 GNDA.n557 292.5
R1021 GNDA.n711 GNDA.n710 292.5
R1022 GNDA.n712 GNDA.n711 292.5
R1023 GNDA.n708 GNDA.n589 292.5
R1024 GNDA.n589 GNDA.n588 292.5
R1025 GNDA.n706 GNDA.n705 292.5
R1026 GNDA.n705 GNDA.n704 292.5
R1027 GNDA.n590 GNDA.n586 292.5
R1028 GNDA.n588 GNDA.n586 292.5
R1029 GNDA.n548 GNDA.n521 292.5
R1030 GNDA.n713 GNDA.n548 292.5
R1031 GNDA.n763 GNDA.n762 292.5
R1032 GNDA.n764 GNDA.n763 292.5
R1033 GNDA.n761 GNDA.n547 292.5
R1034 GNDA.n727 GNDA.n547 292.5
R1035 GNDA.n766 GNDA.n765 292.5
R1036 GNDA.n765 GNDA.n764 292.5
R1037 GNDA.n769 GNDA.n768 292.5
R1038 GNDA.n770 GNDA.n769 292.5
R1039 GNDA.n767 GNDA.n528 292.5
R1040 GNDA.n764 GNDA.n528 292.5
R1041 GNDA.n729 GNDA.n538 292.5
R1042 GNDA.n730 GNDA.n729 292.5
R1043 GNDA.n535 GNDA.n527 292.5
R1044 GNDA.n764 GNDA.n527 292.5
R1045 GNDA.n755 GNDA.n754 292.5
R1046 GNDA.n756 GNDA.n755 292.5
R1047 GNDA.n555 GNDA.n550 292.5
R1048 GNDA.n703 GNDA.n550 292.5
R1049 GNDA.n742 GNDA.n741 292.5
R1050 GNDA.n741 GNDA.n740 292.5
R1051 GNDA.n753 GNDA.n551 292.5
R1052 GNDA.n703 GNDA.n551 292.5
R1053 GNDA.n611 GNDA.n609 292.5
R1054 GNDA.n613 GNDA.n609 292.5
R1055 GNDA.n620 GNDA.n619 292.5
R1056 GNDA.n619 GNDA.n618 292.5
R1057 GNDA.n639 GNDA.n638 292.5
R1058 GNDA.n640 GNDA.n639 292.5
R1059 GNDA.n637 GNDA.n605 292.5
R1060 GNDA.n608 GNDA.n605 292.5
R1061 GNDA.n636 GNDA.n635 292.5
R1062 GNDA.n635 GNDA.n634 292.5
R1063 GNDA.n607 GNDA.n604 292.5
R1064 GNDA.n608 GNDA.n604 292.5
R1065 GNDA.n596 GNDA.n594 292.5
R1066 GNDA.n596 GNDA.n562 292.5
R1067 GNDA.n658 GNDA.n657 292.5
R1068 GNDA.n657 GNDA.n656 292.5
R1069 GNDA.n595 GNDA.n593 292.5
R1070 GNDA.n642 GNDA.n595 292.5
R1071 GNDA.n655 GNDA.n654 292.5
R1072 GNDA.n656 GNDA.n655 292.5
R1073 GNDA.n603 GNDA.n600 292.5
R1074 GNDA.n603 GNDA.n602 292.5
R1075 GNDA.n650 GNDA.n649 292.5
R1076 GNDA.n649 GNDA.t46 292.5
R1077 GNDA.n601 GNDA.n599 292.5
R1078 GNDA.n641 GNDA.n601 292.5
R1079 GNDA.n648 GNDA.n647 292.5
R1080 GNDA.t46 GNDA.n648 292.5
R1081 GNDA.n632 GNDA.n631 292.5
R1082 GNDA.n633 GNDA.n632 292.5
R1083 GNDA.n629 GNDA.n610 292.5
R1084 GNDA.n625 GNDA.n610 292.5
R1085 GNDA.n628 GNDA.n627 292.5
R1086 GNDA.n627 GNDA.n626 292.5
R1087 GNDA.n584 GNDA.n583 292.5
R1088 GNDA.n585 GNDA.n584 292.5
R1089 GNDA.n798 GNDA.n797 292.5
R1090 GNDA.n799 GNDA.n798 292.5
R1091 GNDA.n796 GNDA.n512 292.5
R1092 GNDA.n714 GNDA.n512 292.5
R1093 GNDA.n716 GNDA.n519 292.5
R1094 GNDA.n717 GNDA.n716 292.5
R1095 GNDA.n517 GNDA.n511 292.5
R1096 GNDA.n714 GNDA.n511 292.5
R1097 GNDA.n803 GNDA.n802 292.5
R1098 GNDA.t89 GNDA.n803 292.5
R1099 GNDA.n509 GNDA.n507 292.5
R1100 GNDA.n715 GNDA.n509 292.5
R1101 GNDA.n805 GNDA.n804 292.5
R1102 GNDA.n804 GNDA.t89 292.5
R1103 GNDA.n806 GNDA.n506 292.5
R1104 GNDA.n510 GNDA.n506 292.5
R1105 GNDA.n495 GNDA.n491 292.5
R1106 GNDA.n496 GNDA.n495 292.5
R1107 GNDA.n581 GNDA.n580 292.5
R1108 GNDA.n580 GNDA.n579 292.5
R1109 GNDA.n582 GNDA.n573 292.5
R1110 GNDA.n575 GNDA.n573 292.5
R1111 GNDA.n574 GNDA.n572 292.5
R1112 GNDA.n575 GNDA.n572 292.5
R1113 GNDA.n1505 GNDA.n1504 292.5
R1114 GNDA.n1504 GNDA.n1503 292.5
R1115 GNDA.n1478 GNDA.n1473 292.5
R1116 GNDA.n1495 GNDA.n1473 292.5
R1117 GNDA.n1481 GNDA.n1480 292.5
R1118 GNDA.n1482 GNDA.n1481 292.5
R1119 GNDA.n1472 GNDA.n1469 292.5
R1120 GNDA.n1495 GNDA.n1472 292.5
R1121 GNDA.n1526 GNDA.n1525 292.5
R1122 GNDA.n1525 GNDA.n1524 292.5
R1123 GNDA.n1508 GNDA.n818 292.5
R1124 GNDA.n1545 GNDA.n818 292.5
R1125 GNDA.n1506 GNDA.n1468 292.5
R1126 GNDA.n1502 GNDA.n1468 292.5
R1127 GNDA.n1465 GNDA.n816 292.5
R1128 GNDA.n1545 GNDA.n816 292.5
R1129 GNDA.n1532 GNDA.n1531 292.5
R1130 GNDA.n1533 GNDA.n1532 292.5
R1131 GNDA.n1529 GNDA.n1460 292.5
R1132 GNDA.n1513 GNDA.n1460 292.5
R1133 GNDA.n1527 GNDA.n1464 292.5
R1134 GNDA.n1523 GNDA.n1464 292.5
R1135 GNDA.n1461 GNDA.n1459 292.5
R1136 GNDA.n1513 GNDA.n1459 292.5
R1137 GNDA.n1542 GNDA.n820 292.5
R1138 GNDA.n1514 GNDA.n820 292.5
R1139 GNDA.n1544 GNDA.n1543 292.5
R1140 GNDA.n1545 GNDA.n1544 292.5
R1141 GNDA.n821 GNDA.n819 292.5
R1142 GNDA.n1483 GNDA.n819 292.5
R1143 GNDA.n1541 GNDA.n815 292.5
R1144 GNDA.n1545 GNDA.n815 292.5
R1145 GNDA.n1489 GNDA.n1486 292.5
R1146 GNDA.n1486 GNDA.n814 292.5
R1147 GNDA.n1493 GNDA.n1492 292.5
R1148 GNDA.n1494 GNDA.n1493 292.5
R1149 GNDA.n1487 GNDA.n1485 292.5
R1150 GNDA.n1485 GNDA.n1484 292.5
R1151 GNDA.n1488 GNDA.n1476 292.5
R1152 GNDA.n1494 GNDA.n1476 292.5
R1153 GNDA.n1536 GNDA.n1535 292.5
R1154 GNDA.n1535 GNDA.n1534 292.5
R1155 GNDA.n1537 GNDA.n852 292.5
R1156 GNDA.n1522 GNDA.n852 292.5
R1157 GNDA.n854 GNDA.n851 292.5
R1158 GNDA.n854 GNDA.n817 292.5
R1159 GNDA.n855 GNDA.n853 292.5
R1160 GNDA.n1522 GNDA.n855 292.5
R1161 GNDA.n810 GNDA.n809 292.5
R1162 GNDA.n811 GNDA.n810 292.5
R1163 GNDA.n808 GNDA.n490 292.5
R1164 GNDA.n578 GNDA.n490 292.5
R1165 GNDA.n576 GNDA.n503 292.5
R1166 GNDA.n577 GNDA.n576 292.5
R1167 GNDA.n502 GNDA.n489 292.5
R1168 GNDA.n578 GNDA.n489 292.5
R1169 GNDA.n1500 GNDA.n1499 292.5
R1170 GNDA.n1501 GNDA.n1500 292.5
R1171 GNDA.n1497 GNDA.n1496 292.5
R1172 GNDA.n1494 GNDA.n1475 292.5
R1173 GNDA.n1519 GNDA.n1516 292.5
R1174 GNDA.n1516 GNDA.n1515 292.5
R1175 GNDA.n1518 GNDA.n1510 292.5
R1176 GNDA.n1522 GNDA.n1510 292.5
R1177 GNDA.n1517 GNDA.n1512 292.5
R1178 GNDA.n1512 GNDA.n1511 292.5
R1179 GNDA.n1521 GNDA.n1520 292.5
R1180 GNDA.n1522 GNDA.n1521 292.5
R1181 GNDA.n1734 GNDA.n1728 292.5
R1182 GNDA.n1743 GNDA.n1728 292.5
R1183 GNDA.n1736 GNDA.n1735 292.5
R1184 GNDA.n1736 GNDA.n1718 292.5
R1185 GNDA.n1737 GNDA.n1733 292.5
R1186 GNDA.n1737 GNDA.n1699 292.5
R1187 GNDA.n1739 GNDA.n1738 292.5
R1188 GNDA.n1738 GNDA.n1718 292.5
R1189 GNDA.n1405 GNDA.n1404 292.5
R1190 GNDA.n1406 GNDA.n1405 292.5
R1191 GNDA.n1403 GNDA.n477 292.5
R1192 GNDA.n1566 GNDA.n477 292.5
R1193 GNDA.n1402 GNDA.n1401 292.5
R1194 GNDA.n1401 GNDA.n1400 292.5
R1195 GNDA.n480 GNDA.n475 292.5
R1196 GNDA.n1566 GNDA.n475 292.5
R1197 GNDA.n1742 GNDA.n1741 292.5
R1198 GNDA.n1743 GNDA.n1742 292.5
R1199 GNDA.n1740 GNDA.n1730 292.5
R1200 GNDA.n1730 GNDA.n1718 292.5
R1201 GNDA.n1732 GNDA.n1731 292.5
R1202 GNDA.n1731 GNDA.n1699 292.5
R1203 GNDA.n1729 GNDA.n470 292.5
R1204 GNDA.n1729 GNDA.n1718 292.5
R1205 GNDA.n1565 GNDA.n1564 292.5
R1206 GNDA.n1566 GNDA.n1565 292.5
R1207 GNDA.n1555 GNDA.n485 292.5
R1208 GNDA.n485 GNDA.n466 292.5
R1209 GNDA.n1936 GNDA.n1935 292.5
R1210 GNDA.n1937 GNDA.n1936 292.5
R1211 GNDA.n469 GNDA.n467 292.5
R1212 GNDA.n483 GNDA.n467 292.5
R1213 GNDA.n1933 GNDA.n1932 292.5
R1214 GNDA.n1932 GNDA.n1931 292.5
R1215 GNDA.n1934 GNDA.n468 292.5
R1216 GNDA.n1718 GNDA.n468 292.5
R1217 GNDA.n1741 GNDA.n470 291.2
R1218 GNDA.n1741 GNDA.n1740 291.2
R1219 GNDA.n1739 GNDA.n1734 291.2
R1220 GNDA.n1735 GNDA.n1734 291.2
R1221 GNDA.n1518 GNDA.n1517 288
R1222 GNDA.n1508 GNDA.n1507 288
R1223 GNDA.n1509 GNDA.n1508 288
R1224 GNDA.n1704 GNDA.n1699 270.392
R1225 GNDA.n552 GNDA.t267 258.601
R1226 GNDA.n554 GNDA.t257 258.601
R1227 GNDA.n301 GNDA.n242 258.334
R1228 GNDA.n921 GNDA.n876 258.334
R1229 GNDA.n1353 GNDA.n1295 258.334
R1230 GNDA.n2084 GNDA.n2029 258.334
R1231 GNDA.n147 GNDA.n88 258.334
R1232 GNDA.n1824 GNDA.n1782 258.334
R1233 GNDA.n2237 GNDA.n2169 258.334
R1234 GNDA.n1646 GNDA.n1592 258.334
R1235 GNDA.n1029 GNDA.n984 258.334
R1236 GNDA.n2440 GNDA.n50 257.466
R1237 GNDA.n1193 GNDA.n968 257.466
R1238 GNDA.n2130 GNDA.n412 257.466
R1239 GNDA.n2153 GNDA.n393 257.466
R1240 GNDA.n2387 GNDA.n193 257.466
R1241 GNDA.n2443 GNDA.n41 257.466
R1242 GNDA.n2346 GNDA.n346 257.466
R1243 GNDA.n1141 GNDA.n1076 257.466
R1244 GNDA.n1455 GNDA.n859 257.466
R1245 GNDA.n1139 GNDA.n1138 254.442
R1246 GNDA.n2366 GNDA.n2365 254.34
R1247 GNDA.n2367 GNDA.n2366 254.34
R1248 GNDA.n2366 GNDA.n2364 254.34
R1249 GNDA.n2366 GNDA.n2362 254.34
R1250 GNDA.n2366 GNDA.n2361 254.34
R1251 GNDA.n2366 GNDA.n191 254.34
R1252 GNDA.n194 GNDA.n13 254.34
R1253 GNDA.n2369 GNDA.n194 254.34
R1254 GNDA.n2376 GNDA.n194 254.34
R1255 GNDA.n201 GNDA.n194 254.34
R1256 GNDA.n2383 GNDA.n194 254.34
R1257 GNDA.n2386 GNDA.n194 254.34
R1258 GNDA.n2125 GNDA.n2124 254.34
R1259 GNDA.n2124 GNDA.n2123 254.34
R1260 GNDA.n2124 GNDA.n2012 254.34
R1261 GNDA.n2124 GNDA.n2011 254.34
R1262 GNDA.n2124 GNDA.n2010 254.34
R1263 GNDA.n2124 GNDA.n2009 254.34
R1264 GNDA.n2323 GNDA.n2322 254.34
R1265 GNDA.n2322 GNDA.n2321 254.34
R1266 GNDA.n2322 GNDA.n368 254.34
R1267 GNDA.n2322 GNDA.n367 254.34
R1268 GNDA.n2322 GNDA.n366 254.34
R1269 GNDA.n2322 GNDA.n365 254.34
R1270 GNDA.n2270 GNDA.n2269 254.34
R1271 GNDA.n2270 GNDA.n387 254.34
R1272 GNDA.n2270 GNDA.n386 254.34
R1273 GNDA.n2270 GNDA.n385 254.34
R1274 GNDA.n2270 GNDA.n384 254.34
R1275 GNDA.n2270 GNDA.n383 254.34
R1276 GNDA.n1153 GNDA.n856 254.34
R1277 GNDA.n1051 GNDA.n856 254.34
R1278 GNDA.n1062 GNDA.n856 254.34
R1279 GNDA.n1064 GNDA.n856 254.34
R1280 GNDA.n1074 GNDA.n856 254.34
R1281 GNDA.n1142 GNDA.n856 254.34
R1282 GNDA.n1927 GNDA.n1692 254.34
R1283 GNDA.n1763 GNDA.n1713 254.34
R1284 GNDA.n427 GNDA.n426 254.34
R1285 GNDA.n427 GNDA.n424 254.34
R1286 GNDA.n427 GNDA.n423 254.34
R1287 GNDA.n427 GNDA.n421 254.34
R1288 GNDA.n427 GNDA.n420 254.34
R1289 GNDA.n427 GNDA.n417 254.34
R1290 GNDA.n450 GNDA.n427 254.34
R1291 GNDA.n444 GNDA.n427 254.34
R1292 GNDA.n441 GNDA.n427 254.34
R1293 GNDA.n435 GNDA.n427 254.34
R1294 GNDA.n432 GNDA.n427 254.34
R1295 GNDA.n2005 GNDA.n427 254.34
R1296 GNDA.n2135 GNDA.n394 254.34
R1297 GNDA.n407 GNDA.n394 254.34
R1298 GNDA.n2142 GNDA.n394 254.34
R1299 GNDA.n401 GNDA.n394 254.34
R1300 GNDA.n2149 GNDA.n394 254.34
R1301 GNDA.n2152 GNDA.n394 254.34
R1302 GNDA.n1986 GNDA.n394 254.34
R1303 GNDA.n447 GNDA.n394 254.34
R1304 GNDA.n1993 GNDA.n394 254.34
R1305 GNDA.n438 GNDA.n394 254.34
R1306 GNDA.n2000 GNDA.n394 254.34
R1307 GNDA.n430 GNDA.n394 254.34
R1308 GNDA.n1687 GNDA.n1686 254.34
R1309 GNDA.n1686 GNDA.n1685 254.34
R1310 GNDA.n1686 GNDA.n1575 254.34
R1311 GNDA.n1686 GNDA.n1574 254.34
R1312 GNDA.n1686 GNDA.n1573 254.34
R1313 GNDA.n1686 GNDA.n1572 254.34
R1314 GNDA.n1431 GNDA.n1430 254.34
R1315 GNDA.n1430 GNDA.n1429 254.34
R1316 GNDA.n1430 GNDA.n1237 254.34
R1317 GNDA.n1430 GNDA.n1236 254.34
R1318 GNDA.n1430 GNDA.n1235 254.34
R1319 GNDA.n1430 GNDA.n1234 254.34
R1320 GNDA.n1275 GNDA.n1274 254.34
R1321 GNDA.n1394 GNDA.n1393 254.34
R1322 GNDA.n1393 GNDA.n1392 254.34
R1323 GNDA.n1205 GNDA.n856 254.34
R1324 GNDA.n943 GNDA.n856 254.34
R1325 GNDA.n954 GNDA.n856 254.34
R1326 GNDA.n956 GNDA.n856 254.34
R1327 GNDA.n966 GNDA.n856 254.34
R1328 GNDA.n1194 GNDA.n856 254.34
R1329 GNDA.n1229 GNDA.n427 254.34
R1330 GNDA.n1227 GNDA.n427 254.34
R1331 GNDA.n1224 GNDA.n427 254.34
R1332 GNDA.n1218 GNDA.n427 254.34
R1333 GNDA.n1215 GNDA.n427 254.34
R1334 GNDA.n1209 GNDA.n427 254.34
R1335 GNDA.n1434 GNDA.n394 254.34
R1336 GNDA.n1232 GNDA.n394 254.34
R1337 GNDA.n1441 GNDA.n394 254.34
R1338 GNDA.n1221 GNDA.n394 254.34
R1339 GNDA.n1448 GNDA.n394 254.34
R1340 GNDA.n1212 GNDA.n394 254.34
R1341 GNDA.n2272 GNDA.n222 254.34
R1342 GNDA.n2277 GNDA.n2272 254.34
R1343 GNDA.n2284 GNDA.n2272 254.34
R1344 GNDA.n2275 GNDA.n2272 254.34
R1345 GNDA.n2291 GNDA.n2272 254.34
R1346 GNDA.n2272 GNDA.n382 254.34
R1347 GNDA.n1115 GNDA.n42 254.34
R1348 GNDA.n1109 GNDA.n42 254.34
R1349 GNDA.n1107 GNDA.n42 254.34
R1350 GNDA.n1101 GNDA.n42 254.34
R1351 GNDA.n1099 GNDA.n42 254.34
R1352 GNDA.n1094 GNDA.n42 254.34
R1353 GNDA.n2366 GNDA.n2358 254.34
R1354 GNDA.n2366 GNDA.n216 254.34
R1355 GNDA.n2366 GNDA.n215 254.34
R1356 GNDA.n2366 GNDA.n214 254.34
R1357 GNDA.n2366 GNDA.n213 254.34
R1358 GNDA.n2366 GNDA.n212 254.34
R1359 GNDA.n221 GNDA.n194 254.34
R1360 GNDA.n1172 GNDA.n194 254.34
R1361 GNDA.n1179 GNDA.n194 254.34
R1362 GNDA.n1167 GNDA.n194 254.34
R1363 GNDA.n1186 GNDA.n194 254.34
R1364 GNDA.n1160 GNDA.n194 254.34
R1365 GNDA.n2366 GNDA.n211 254.34
R1366 GNDA.n2366 GNDA.n210 254.34
R1367 GNDA.n2366 GNDA.n209 254.34
R1368 GNDA.n2366 GNDA.n208 254.34
R1369 GNDA.n2366 GNDA.n207 254.34
R1370 GNDA.n2366 GNDA.n206 254.34
R1371 GNDA.n2328 GNDA.n194 254.34
R1372 GNDA.n363 GNDA.n194 254.34
R1373 GNDA.n2335 GNDA.n194 254.34
R1374 GNDA.n356 GNDA.n194 254.34
R1375 GNDA.n2342 GNDA.n194 254.34
R1376 GNDA.n2345 GNDA.n194 254.34
R1377 GNDA.n226 GNDA.n47 254.34
R1378 GNDA.n229 GNDA.n47 254.34
R1379 GNDA.n262 GNDA.n47 254.34
R1380 GNDA.n264 GNDA.n47 254.34
R1381 GNDA.n277 GNDA.n47 254.34
R1382 GNDA.n279 GNDA.n47 254.34
R1383 GNDA.n62 GNDA.n45 254.34
R1384 GNDA.n2412 GNDA.n45 254.34
R1385 GNDA.n2406 GNDA.n45 254.34
R1386 GNDA.n2404 GNDA.n45 254.34
R1387 GNDA.n2398 GNDA.n45 254.34
R1388 GNDA.n2396 GNDA.n45 254.34
R1389 GNDA.n72 GNDA.n44 254.34
R1390 GNDA.n75 GNDA.n44 254.34
R1391 GNDA.n108 GNDA.n44 254.34
R1392 GNDA.n110 GNDA.n44 254.34
R1393 GNDA.n123 GNDA.n44 254.34
R1394 GNDA.n125 GNDA.n44 254.34
R1395 GNDA.n2439 GNDA.n2438 254.34
R1396 GNDA.n2445 GNDA.n2444 254.34
R1397 GNDA.n2418 GNDA.n2417 251.614
R1398 GNDA.n2355 GNDA.n2354 251.614
R1399 GNDA.n1985 GNDA.n448 251.614
R1400 GNDA.n2134 GNDA.n2132 251.614
R1401 GNDA.n2496 GNDA.n2495 251.614
R1402 GNDA.n2468 GNDA.n30 251.614
R1403 GNDA.n2327 GNDA.n2324 251.614
R1404 GNDA.n1117 GNDA.n1116 251.614
R1405 GNDA.n1433 GNDA.n1432 251.614
R1406 GNDA.n2513 GNDA.n2512 250.349
R1407 GNDA.n1304 GNDA.t229 239.004
R1408 GNDA.n622 GNDA.n621 238.4
R1409 GNDA.n500 GNDA.n499 238.4
R1410 GNDA.n733 GNDA.n559 233.601
R1411 GNDA.n737 GNDA.n559 233.601
R1412 GNDA.n748 GNDA.n746 227.096
R1413 GNDA.n745 GNDA.n743 227.096
R1414 GNDA.n748 GNDA.n747 226.534
R1415 GNDA.n745 GNDA.n744 226.534
R1416 GNDA.n597 GNDA.t303 224.525
R1417 GNDA.n513 GNDA.t244 224.525
R1418 GNDA.n516 GNDA.t232 224.525
R1419 GNDA.n652 GNDA.t291 224.525
R1420 GNDA.n1530 GNDA.n1529 224
R1421 GNDA.n1529 GNDA.n1528 224
R1422 GNDA.n1479 GNDA.n1478 224
R1423 GNDA.n1478 GNDA.n1471 224
R1424 GNDA.n751 GNDA.n750 222.034
R1425 GNDA.n1930 GNDA.n1567 221.23
R1426 GNDA.n556 GNDA.n555 211.201
R1427 GNDA.n555 GNDA.n553 211.201
R1428 GNDA.n647 GNDA.n644 211.201
R1429 GNDA.n647 GNDA.n646 211.201
R1430 GNDA.n630 GNDA.n629 211.201
R1431 GNDA.n802 GNDA.n801 211.201
R1432 GNDA.n802 GNDA.n505 211.201
R1433 GNDA.n808 GNDA.n807 211.201
R1434 GNDA.n779 GNDA.n777 206.052
R1435 GNDA.n664 GNDA.n662 206.052
R1436 GNDA.n787 GNDA.n786 205.488
R1437 GNDA.n785 GNDA.n784 205.488
R1438 GNDA.n783 GNDA.n782 205.488
R1439 GNDA.n781 GNDA.n780 205.488
R1440 GNDA.n779 GNDA.n778 205.488
R1441 GNDA.n672 GNDA.n671 205.488
R1442 GNDA.n670 GNDA.n669 205.488
R1443 GNDA.n668 GNDA.n667 205.488
R1444 GNDA.n666 GNDA.n665 205.488
R1445 GNDA.n664 GNDA.n663 205.488
R1446 GNDA.n1407 GNDA.n1406 200.161
R1447 GNDA.t11 GNDA.n1715 200.161
R1448 GNDA.n1743 GNDA.n465 200.161
R1449 GNDA.n772 GNDA.n523 198.4
R1450 GNDA.n2511 GNDA.n4 197
R1451 GNDA.n772 GNDA.n524 195.201
R1452 GNDA.n2349 GNDA.n2348 195.049
R1453 GNDA.n1208 GNDA.n1207 195.049
R1454 GNDA.n1764 GNDA.n1714 195.049
R1455 GNDA.n1928 GNDA.n1569 195.049
R1456 GNDA.n2007 GNDA.n2006 195.049
R1457 GNDA.n2390 GNDA.n2389 195.049
R1458 GNDA.n391 GNDA.n389 195.049
R1459 GNDA.n1156 GNDA.n1155 195.049
R1460 GNDA.n1246 GNDA.n1244 195.049
R1461 GNDA.n616 GNDA.n615 195
R1462 GNDA.n617 GNDA.n616 195
R1463 GNDA.n623 GNDA.n622 195
R1464 GNDA.n624 GNDA.n623 195
R1465 GNDA.n499 GNDA.n498 195
R1466 GNDA.n498 GNDA.n497 195
R1467 GNDA.n494 GNDA.n492 195
R1468 GNDA.n518 GNDA.n517 192
R1469 GNDA.n654 GNDA.n653 192
R1470 GNDA.t238 GNDA.n2441 190.773
R1471 GNDA.n2442 GNDA.t238 190.773
R1472 GNDA.n2325 GNDA.n68 187.249
R1473 GNDA.n2298 GNDA.n376 187.249
R1474 GNDA.n1727 GNDA.n464 187.249
R1475 GNDA.n1905 GNDA.n1703 187.249
R1476 GNDA.n1982 GNDA.n451 187.249
R1477 GNDA.n2492 GNDA.n15 187.249
R1478 GNDA.n2300 GNDA.n371 187.249
R1479 GNDA.n2357 GNDA.n218 187.249
R1480 GNDA.n1408 GNDA.n1240 187.249
R1481 GNDA.t238 GNDA.n48 186.691
R1482 GNDA.t238 GNDA.n43 186.691
R1483 GNDA.n775 GNDA.n523 185.601
R1484 GNDA.n299 GNDA.n242 185
R1485 GNDA.n242 GNDA.t281 185
R1486 GNDA.n298 GNDA.n297 185
R1487 GNDA.n295 GNDA.n243 185
R1488 GNDA.n294 GNDA.n244 185
R1489 GNDA.n292 GNDA.n291 185
R1490 GNDA.n290 GNDA.n245 185
R1491 GNDA.n289 GNDA.n288 185
R1492 GNDA.n286 GNDA.n246 185
R1493 GNDA.n286 GNDA.t281 185
R1494 GNDA.n285 GNDA.n247 185
R1495 GNDA.n301 GNDA.n300 185
R1496 GNDA.n303 GNDA.n240 185
R1497 GNDA.n305 GNDA.n304 185
R1498 GNDA.n306 GNDA.n239 185
R1499 GNDA.n308 GNDA.n307 185
R1500 GNDA.n310 GNDA.n237 185
R1501 GNDA.n312 GNDA.n311 185
R1502 GNDA.n313 GNDA.n236 185
R1503 GNDA.n315 GNDA.n314 185
R1504 GNDA.n317 GNDA.n235 185
R1505 GNDA.n320 GNDA.n319 185
R1506 GNDA.n321 GNDA.n234 185
R1507 GNDA.n323 GNDA.n322 185
R1508 GNDA.n325 GNDA.n233 185
R1509 GNDA.n328 GNDA.n327 185
R1510 GNDA.n329 GNDA.n232 185
R1511 GNDA.n331 GNDA.n330 185
R1512 GNDA.n333 GNDA.n227 185
R1513 GNDA.n923 GNDA.n876 185
R1514 GNDA.t237 GNDA.n876 185
R1515 GNDA.n925 GNDA.n924 185
R1516 GNDA.n927 GNDA.n926 185
R1517 GNDA.n929 GNDA.n928 185
R1518 GNDA.n931 GNDA.n930 185
R1519 GNDA.n933 GNDA.n932 185
R1520 GNDA.n935 GNDA.n934 185
R1521 GNDA.n936 GNDA.n881 185
R1522 GNDA.t237 GNDA.n881 185
R1523 GNDA.n937 GNDA.n885 185
R1524 GNDA.n922 GNDA.n921 185
R1525 GNDA.n920 GNDA.n919 185
R1526 GNDA.n918 GNDA.n917 185
R1527 GNDA.n916 GNDA.n915 185
R1528 GNDA.n914 GNDA.n913 185
R1529 GNDA.n912 GNDA.n911 185
R1530 GNDA.n910 GNDA.n909 185
R1531 GNDA.n908 GNDA.n907 185
R1532 GNDA.n906 GNDA.n905 185
R1533 GNDA.n904 GNDA.n903 185
R1534 GNDA.n902 GNDA.n901 185
R1535 GNDA.n900 GNDA.n899 185
R1536 GNDA.n898 GNDA.n897 185
R1537 GNDA.n896 GNDA.n895 185
R1538 GNDA.n894 GNDA.n893 185
R1539 GNDA.n892 GNDA.n891 185
R1540 GNDA.n890 GNDA.n889 185
R1541 GNDA.n888 GNDA.n866 185
R1542 GNDA.n1351 GNDA.n1295 185
R1543 GNDA.n1295 GNDA.t233 185
R1544 GNDA.n1350 GNDA.n1349 185
R1545 GNDA.n1347 GNDA.n1296 185
R1546 GNDA.n1346 GNDA.n1297 185
R1547 GNDA.n1344 GNDA.n1343 185
R1548 GNDA.n1342 GNDA.n1298 185
R1549 GNDA.n1341 GNDA.n1340 185
R1550 GNDA.n1338 GNDA.n1299 185
R1551 GNDA.n1338 GNDA.t233 185
R1552 GNDA.n1337 GNDA.n1300 185
R1553 GNDA.n1353 GNDA.n1352 185
R1554 GNDA.n1355 GNDA.n1293 185
R1555 GNDA.n1357 GNDA.n1356 185
R1556 GNDA.n1358 GNDA.n1292 185
R1557 GNDA.n1360 GNDA.n1359 185
R1558 GNDA.n1362 GNDA.n1290 185
R1559 GNDA.n1364 GNDA.n1363 185
R1560 GNDA.n1365 GNDA.n1289 185
R1561 GNDA.n1367 GNDA.n1366 185
R1562 GNDA.n1369 GNDA.n1288 185
R1563 GNDA.n1371 GNDA.n1370 185
R1564 GNDA.n1373 GNDA.n1372 185
R1565 GNDA.n1376 GNDA.n1375 185
R1566 GNDA.n1377 GNDA.n1286 185
R1567 GNDA.n1379 GNDA.n1378 185
R1568 GNDA.n1381 GNDA.n1285 185
R1569 GNDA.n1383 GNDA.n1382 185
R1570 GNDA.n1385 GNDA.n1384 185
R1571 GNDA.n2082 GNDA.n2029 185
R1572 GNDA.n2029 GNDA.t319 185
R1573 GNDA.n2081 GNDA.n2080 185
R1574 GNDA.n2078 GNDA.n2030 185
R1575 GNDA.n2077 GNDA.n2031 185
R1576 GNDA.n2075 GNDA.n2074 185
R1577 GNDA.n2073 GNDA.n2032 185
R1578 GNDA.n2072 GNDA.n2071 185
R1579 GNDA.n2069 GNDA.n2033 185
R1580 GNDA.n2069 GNDA.t319 185
R1581 GNDA.n2068 GNDA.n2034 185
R1582 GNDA.n2084 GNDA.n2083 185
R1583 GNDA.n2086 GNDA.n2027 185
R1584 GNDA.n2088 GNDA.n2087 185
R1585 GNDA.n2089 GNDA.n2026 185
R1586 GNDA.n2091 GNDA.n2090 185
R1587 GNDA.n2093 GNDA.n2024 185
R1588 GNDA.n2095 GNDA.n2094 185
R1589 GNDA.n2096 GNDA.n2023 185
R1590 GNDA.n2098 GNDA.n2097 185
R1591 GNDA.n2100 GNDA.n2022 185
R1592 GNDA.n2102 GNDA.n2101 185
R1593 GNDA.n2104 GNDA.n2103 185
R1594 GNDA.n2107 GNDA.n2106 185
R1595 GNDA.n2108 GNDA.n2020 185
R1596 GNDA.n2110 GNDA.n2109 185
R1597 GNDA.n2112 GNDA.n2019 185
R1598 GNDA.n2114 GNDA.n2113 185
R1599 GNDA.n2116 GNDA.n2115 185
R1600 GNDA.n145 GNDA.n88 185
R1601 GNDA.n88 GNDA.t245 185
R1602 GNDA.n144 GNDA.n143 185
R1603 GNDA.n141 GNDA.n89 185
R1604 GNDA.n140 GNDA.n90 185
R1605 GNDA.n138 GNDA.n137 185
R1606 GNDA.n136 GNDA.n91 185
R1607 GNDA.n135 GNDA.n134 185
R1608 GNDA.n132 GNDA.n92 185
R1609 GNDA.n132 GNDA.t245 185
R1610 GNDA.n131 GNDA.n93 185
R1611 GNDA.n147 GNDA.n146 185
R1612 GNDA.n149 GNDA.n86 185
R1613 GNDA.n151 GNDA.n150 185
R1614 GNDA.n152 GNDA.n85 185
R1615 GNDA.n154 GNDA.n153 185
R1616 GNDA.n156 GNDA.n83 185
R1617 GNDA.n158 GNDA.n157 185
R1618 GNDA.n159 GNDA.n82 185
R1619 GNDA.n161 GNDA.n160 185
R1620 GNDA.n163 GNDA.n81 185
R1621 GNDA.n166 GNDA.n165 185
R1622 GNDA.n167 GNDA.n80 185
R1623 GNDA.n169 GNDA.n168 185
R1624 GNDA.n171 GNDA.n79 185
R1625 GNDA.n174 GNDA.n173 185
R1626 GNDA.n175 GNDA.n78 185
R1627 GNDA.n177 GNDA.n176 185
R1628 GNDA.n179 GNDA.n73 185
R1629 GNDA.n180 GNDA.n74 185
R1630 GNDA.n183 GNDA.n182 185
R1631 GNDA.n104 GNDA.n77 185
R1632 GNDA.n105 GNDA.n101 185
R1633 GNDA.n114 GNDA.n113 185
R1634 GNDA.n116 GNDA.n99 185
R1635 GNDA.n119 GNDA.n118 185
R1636 GNDA.n120 GNDA.n94 185
R1637 GNDA.n129 GNDA.n128 185
R1638 GNDA.n1826 GNDA.n1782 185
R1639 GNDA.t320 GNDA.n1782 185
R1640 GNDA.n1828 GNDA.n1827 185
R1641 GNDA.n1830 GNDA.n1829 185
R1642 GNDA.n1832 GNDA.n1831 185
R1643 GNDA.n1834 GNDA.n1833 185
R1644 GNDA.n1836 GNDA.n1835 185
R1645 GNDA.n1838 GNDA.n1837 185
R1646 GNDA.n1839 GNDA.n1787 185
R1647 GNDA.t320 GNDA.n1787 185
R1648 GNDA.n1841 GNDA.n1840 185
R1649 GNDA.n1825 GNDA.n1824 185
R1650 GNDA.n1823 GNDA.n1822 185
R1651 GNDA.n1821 GNDA.n1820 185
R1652 GNDA.n1819 GNDA.n1818 185
R1653 GNDA.n1817 GNDA.n1816 185
R1654 GNDA.n1815 GNDA.n1814 185
R1655 GNDA.n1813 GNDA.n1812 185
R1656 GNDA.n1811 GNDA.n1810 185
R1657 GNDA.n1809 GNDA.n1808 185
R1658 GNDA.n1807 GNDA.n1806 185
R1659 GNDA.n1805 GNDA.n1804 185
R1660 GNDA.n1803 GNDA.n1802 185
R1661 GNDA.n1801 GNDA.n1800 185
R1662 GNDA.n1799 GNDA.n1798 185
R1663 GNDA.n1797 GNDA.n1796 185
R1664 GNDA.n1795 GNDA.n1794 185
R1665 GNDA.n1793 GNDA.n1792 185
R1666 GNDA.n1791 GNDA.n1772 185
R1667 GNDA.n1897 GNDA.n1896 185
R1668 GNDA.n1854 GNDA.n1773 185
R1669 GNDA.n1853 GNDA.n1852 185
R1670 GNDA.n1870 GNDA.n1869 185
R1671 GNDA.n1872 GNDA.n1871 185
R1672 GNDA.n1876 GNDA.n1874 185
R1673 GNDA.n1878 GNDA.n1877 185
R1674 GNDA.n1843 GNDA.n1842 185
R1675 GNDA.n1893 GNDA.n1892 185
R1676 GNDA.n2117 GNDA.n2015 185
R1677 GNDA.n2120 GNDA.n2119 185
R1678 GNDA.n2042 GNDA.n2017 185
R1679 GNDA.n2045 GNDA.n2041 185
R1680 GNDA.n2050 GNDA.n2049 185
R1681 GNDA.n2053 GNDA.n2052 185
R1682 GNDA.n2039 GNDA.n2036 185
R1683 GNDA.n2058 GNDA.n2035 185
R1684 GNDA.n2066 GNDA.n2065 185
R1685 GNDA.n2239 GNDA.n2169 185
R1686 GNDA.t264 GNDA.n2169 185
R1687 GNDA.n2241 GNDA.n2240 185
R1688 GNDA.n2243 GNDA.n2242 185
R1689 GNDA.n2245 GNDA.n2244 185
R1690 GNDA.n2247 GNDA.n2246 185
R1691 GNDA.n2249 GNDA.n2248 185
R1692 GNDA.n2251 GNDA.n2250 185
R1693 GNDA.n2252 GNDA.n2174 185
R1694 GNDA.t264 GNDA.n2174 185
R1695 GNDA.n2253 GNDA.n2178 185
R1696 GNDA.n2238 GNDA.n2237 185
R1697 GNDA.n2236 GNDA.n2235 185
R1698 GNDA.n2234 GNDA.n2233 185
R1699 GNDA.n2232 GNDA.n2231 185
R1700 GNDA.n2230 GNDA.n2229 185
R1701 GNDA.n2228 GNDA.n2227 185
R1702 GNDA.n2226 GNDA.n2225 185
R1703 GNDA.n2224 GNDA.n2223 185
R1704 GNDA.n2222 GNDA.n2221 185
R1705 GNDA.n2220 GNDA.n2219 185
R1706 GNDA.n2218 GNDA.n2217 185
R1707 GNDA.n2216 GNDA.n2215 185
R1708 GNDA.n2214 GNDA.n2213 185
R1709 GNDA.n2212 GNDA.n2211 185
R1710 GNDA.n2210 GNDA.n2209 185
R1711 GNDA.n2208 GNDA.n2207 185
R1712 GNDA.n2206 GNDA.n2205 185
R1713 GNDA.n2159 GNDA.n2156 185
R1714 GNDA.n1644 GNDA.n1592 185
R1715 GNDA.n1592 GNDA.t228 185
R1716 GNDA.n1643 GNDA.n1642 185
R1717 GNDA.n1640 GNDA.n1593 185
R1718 GNDA.n1639 GNDA.n1594 185
R1719 GNDA.n1637 GNDA.n1636 185
R1720 GNDA.n1635 GNDA.n1595 185
R1721 GNDA.n1634 GNDA.n1633 185
R1722 GNDA.n1631 GNDA.n1596 185
R1723 GNDA.n1631 GNDA.t228 185
R1724 GNDA.n1630 GNDA.n1597 185
R1725 GNDA.n1646 GNDA.n1645 185
R1726 GNDA.n1648 GNDA.n1590 185
R1727 GNDA.n1650 GNDA.n1649 185
R1728 GNDA.n1651 GNDA.n1589 185
R1729 GNDA.n1653 GNDA.n1652 185
R1730 GNDA.n1655 GNDA.n1587 185
R1731 GNDA.n1657 GNDA.n1656 185
R1732 GNDA.n1658 GNDA.n1586 185
R1733 GNDA.n1660 GNDA.n1659 185
R1734 GNDA.n1662 GNDA.n1585 185
R1735 GNDA.n1664 GNDA.n1663 185
R1736 GNDA.n1666 GNDA.n1665 185
R1737 GNDA.n1669 GNDA.n1668 185
R1738 GNDA.n1670 GNDA.n1583 185
R1739 GNDA.n1672 GNDA.n1671 185
R1740 GNDA.n1674 GNDA.n1582 185
R1741 GNDA.n1676 GNDA.n1675 185
R1742 GNDA.n1678 GNDA.n1677 185
R1743 GNDA.n1679 GNDA.n1578 185
R1744 GNDA.n1682 GNDA.n1681 185
R1745 GNDA.n1605 GNDA.n1580 185
R1746 GNDA.n1608 GNDA.n1604 185
R1747 GNDA.n1613 GNDA.n1612 185
R1748 GNDA.n1616 GNDA.n1615 185
R1749 GNDA.n1602 GNDA.n1599 185
R1750 GNDA.n1621 GNDA.n1598 185
R1751 GNDA.n1628 GNDA.n1627 185
R1752 GNDA.n2264 GNDA.n2263 185
R1753 GNDA.n2184 GNDA.n2160 185
R1754 GNDA.n2183 GNDA.n2182 185
R1755 GNDA.n2191 GNDA.n2190 185
R1756 GNDA.n2189 GNDA.n2181 185
R1757 GNDA.n2198 GNDA.n2197 185
R1758 GNDA.n2196 GNDA.n2180 185
R1759 GNDA.n2203 GNDA.n2179 185
R1760 GNDA.n2260 GNDA.n2259 185
R1761 GNDA.n1031 GNDA.n984 185
R1762 GNDA.t288 GNDA.n984 185
R1763 GNDA.n1033 GNDA.n1032 185
R1764 GNDA.n1035 GNDA.n1034 185
R1765 GNDA.n1037 GNDA.n1036 185
R1766 GNDA.n1039 GNDA.n1038 185
R1767 GNDA.n1041 GNDA.n1040 185
R1768 GNDA.n1043 GNDA.n1042 185
R1769 GNDA.n1044 GNDA.n989 185
R1770 GNDA.t288 GNDA.n989 185
R1771 GNDA.n1045 GNDA.n993 185
R1772 GNDA.n1030 GNDA.n1029 185
R1773 GNDA.n1028 GNDA.n1027 185
R1774 GNDA.n1026 GNDA.n1025 185
R1775 GNDA.n1024 GNDA.n1023 185
R1776 GNDA.n1022 GNDA.n1021 185
R1777 GNDA.n1020 GNDA.n1019 185
R1778 GNDA.n1018 GNDA.n1017 185
R1779 GNDA.n1016 GNDA.n1015 185
R1780 GNDA.n1014 GNDA.n1013 185
R1781 GNDA.n1012 GNDA.n1011 185
R1782 GNDA.n1010 GNDA.n1009 185
R1783 GNDA.n1008 GNDA.n1007 185
R1784 GNDA.n1006 GNDA.n1005 185
R1785 GNDA.n1004 GNDA.n1003 185
R1786 GNDA.n1002 GNDA.n1001 185
R1787 GNDA.n1000 GNDA.n999 185
R1788 GNDA.n998 GNDA.n997 185
R1789 GNDA.n996 GNDA.n974 185
R1790 GNDA.n1150 GNDA.n1149 185
R1791 GNDA.n1053 GNDA.n975 185
R1792 GNDA.n1056 GNDA.n1055 185
R1793 GNDA.n1059 GNDA.n1058 185
R1794 GNDA.n1057 GNDA.n1049 185
R1795 GNDA.n1068 GNDA.n1067 185
R1796 GNDA.n1070 GNDA.n1069 185
R1797 GNDA.n1071 GNDA.n994 185
R1798 GNDA.n1146 GNDA.n1145 185
R1799 GNDA.n1386 GNDA.n1281 185
R1800 GNDA.n1389 GNDA.n1388 185
R1801 GNDA.n1311 GNDA.n1283 185
R1802 GNDA.n1310 GNDA.n1309 185
R1803 GNDA.n1320 GNDA.n1319 185
R1804 GNDA.n1322 GNDA.n1306 185
R1805 GNDA.n1325 GNDA.n1324 185
R1806 GNDA.n1302 GNDA.n1301 185
R1807 GNDA.n1335 GNDA.n1334 185
R1808 GNDA.n1202 GNDA.n1201 185
R1809 GNDA.n945 GNDA.n867 185
R1810 GNDA.n948 GNDA.n947 185
R1811 GNDA.n951 GNDA.n950 185
R1812 GNDA.n949 GNDA.n941 185
R1813 GNDA.n960 GNDA.n959 185
R1814 GNDA.n962 GNDA.n961 185
R1815 GNDA.n963 GNDA.n886 185
R1816 GNDA.n1198 GNDA.n1197 185
R1817 GNDA.n334 GNDA.n228 185
R1818 GNDA.n337 GNDA.n336 185
R1819 GNDA.n258 GNDA.n231 185
R1820 GNDA.n259 GNDA.n255 185
R1821 GNDA.n268 GNDA.n267 185
R1822 GNDA.n270 GNDA.n253 185
R1823 GNDA.n273 GNDA.n272 185
R1824 GNDA.n274 GNDA.n248 185
R1825 GNDA.n283 GNDA.n282 185
R1826 GNDA.n775 GNDA.n524 182.4
R1827 GNDA.n646 GNDA.n600 182.4
R1828 GNDA.n801 GNDA.n507 182.4
R1829 GNDA.n718 GNDA.n713 179.363
R1830 GNDA.n644 GNDA.n599 176
R1831 GNDA.n806 GNDA.n505 176
R1832 GNDA.n2399 GNDA.n2397 175.546
R1833 GNDA.n2403 GNDA.n66 175.546
R1834 GNDA.n2407 GNDA.n2405 175.546
R1835 GNDA.n2411 GNDA.n64 175.546
R1836 GNDA.n2414 GNDA.n2413 175.546
R1837 GNDA.n2436 GNDA.n51 175.546
R1838 GNDA.n2436 GNDA.n54 175.546
R1839 GNDA.n2432 GNDA.n54 175.546
R1840 GNDA.n2432 GNDA.n56 175.546
R1841 GNDA.n2428 GNDA.n56 175.546
R1842 GNDA.n2428 GNDA.n58 175.546
R1843 GNDA.n2424 GNDA.n58 175.546
R1844 GNDA.n2424 GNDA.n60 175.546
R1845 GNDA.n2420 GNDA.n60 175.546
R1846 GNDA.n2420 GNDA.n2418 175.546
R1847 GNDA.n340 GNDA.n339 175.546
R1848 GNDA.n261 GNDA.n257 175.546
R1849 GNDA.n265 GNDA.n263 175.546
R1850 GNDA.n276 GNDA.n251 175.546
R1851 GNDA.n280 GNDA.n278 175.546
R1852 GNDA.n348 GNDA.n347 175.546
R1853 GNDA.n352 GNDA.n351 175.546
R1854 GNDA.n354 GNDA.n353 175.546
R1855 GNDA.n359 GNDA.n358 175.546
R1856 GNDA.n361 GNDA.n360 175.546
R1857 GNDA.n1214 GNDA.n1210 175.546
R1858 GNDA.n1217 GNDA.n1216 175.546
R1859 GNDA.n1223 GNDA.n1219 175.546
R1860 GNDA.n1226 GNDA.n1225 175.546
R1861 GNDA.n1230 GNDA.n1228 175.546
R1862 GNDA.n2293 GNDA.n2292 175.546
R1863 GNDA.n2290 GNDA.n2273 175.546
R1864 GNDA.n2286 GNDA.n2285 175.546
R1865 GNDA.n2283 GNDA.n2276 175.546
R1866 GNDA.n2279 GNDA.n2278 175.546
R1867 GNDA.n1188 GNDA.n1187 175.546
R1868 GNDA.n1185 GNDA.n1161 175.546
R1869 GNDA.n1181 GNDA.n1180 175.546
R1870 GNDA.n1178 GNDA.n1168 175.546
R1871 GNDA.n1174 GNDA.n1173 175.546
R1872 GNDA.n1204 GNDA.n863 175.546
R1873 GNDA.n953 GNDA.n944 175.546
R1874 GNDA.n957 GNDA.n955 175.546
R1875 GNDA.n965 GNDA.n939 175.546
R1876 GNDA.n1195 GNDA.n967 175.546
R1877 GNDA.n1762 GNDA.n1761 175.546
R1878 GNDA.n1761 GNDA.n1716 175.546
R1879 GNDA.n1757 GNDA.n1716 175.546
R1880 GNDA.n1757 GNDA.n1720 175.546
R1881 GNDA.n1753 GNDA.n1720 175.546
R1882 GNDA.n1753 GNDA.n1722 175.546
R1883 GNDA.n1749 GNDA.n1722 175.546
R1884 GNDA.n1749 GNDA.n1724 175.546
R1885 GNDA.n1745 GNDA.n1724 175.546
R1886 GNDA.n1745 GNDA.n1727 175.546
R1887 GNDA.n1941 GNDA.n462 175.546
R1888 GNDA.n1945 GNDA.n462 175.546
R1889 GNDA.n1945 GNDA.n460 175.546
R1890 GNDA.n1950 GNDA.n460 175.546
R1891 GNDA.n1950 GNDA.n458 175.546
R1892 GNDA.n1954 GNDA.n458 175.546
R1893 GNDA.n1954 GNDA.n457 175.546
R1894 GNDA.n1958 GNDA.n457 175.546
R1895 GNDA.n1958 GNDA.n455 175.546
R1896 GNDA.n1963 GNDA.n455 175.546
R1897 GNDA.n1963 GNDA.n448 175.546
R1898 GNDA.n2002 GNDA.n2001 175.546
R1899 GNDA.n1999 GNDA.n431 175.546
R1900 GNDA.n1995 GNDA.n1994 175.546
R1901 GNDA.n1992 GNDA.n439 175.546
R1902 GNDA.n1988 GNDA.n1987 175.546
R1903 GNDA.n1899 GNDA.n1711 175.546
R1904 GNDA.n1899 GNDA.n1712 175.546
R1905 GNDA.n1856 GNDA.n1712 175.546
R1906 GNDA.n1867 GNDA.n1856 175.546
R1907 GNDA.n1867 GNDA.n1857 175.546
R1908 GNDA.n1857 GNDA.n1850 175.546
R1909 GNDA.n1880 GNDA.n1850 175.546
R1910 GNDA.n1880 GNDA.n1844 175.546
R1911 GNDA.n1889 GNDA.n1844 175.546
R1912 GNDA.n1889 GNDA.n411 175.546
R1913 GNDA.n2130 GNDA.n411 175.546
R1914 GNDA.n1926 GNDA.n1925 175.546
R1915 GNDA.n1925 GNDA.n1693 175.546
R1916 GNDA.n1921 GNDA.n1693 175.546
R1917 GNDA.n1921 GNDA.n1696 175.546
R1918 GNDA.n1917 GNDA.n1696 175.546
R1919 GNDA.n1917 GNDA.n1698 175.546
R1920 GNDA.n1913 GNDA.n1698 175.546
R1921 GNDA.n1913 GNDA.n1700 175.546
R1922 GNDA.n1909 GNDA.n1700 175.546
R1923 GNDA.n1909 GNDA.n1703 175.546
R1924 GNDA.n1684 GNDA.n1571 175.546
R1925 GNDA.n1606 GNDA.n1576 175.546
R1926 GNDA.n1610 GNDA.n1609 175.546
R1927 GNDA.n1619 GNDA.n1618 175.546
R1928 GNDA.n1625 GNDA.n1624 175.546
R1929 GNDA.n2151 GNDA.n2150 175.546
R1930 GNDA.n2148 GNDA.n396 175.546
R1931 GNDA.n2144 GNDA.n2143 175.546
R1932 GNDA.n2141 GNDA.n402 175.546
R1933 GNDA.n2137 GNDA.n2136 175.546
R1934 GNDA.n1901 GNDA.n1706 175.546
R1935 GNDA.n1901 GNDA.n1708 175.546
R1936 GNDA.n1860 GNDA.n1708 175.546
R1937 GNDA.n1860 GNDA.n1859 175.546
R1938 GNDA.n1864 GNDA.n1859 175.546
R1939 GNDA.n1864 GNDA.n1848 175.546
R1940 GNDA.n1882 GNDA.n1848 175.546
R1941 GNDA.n1882 GNDA.n1846 175.546
R1942 GNDA.n1887 GNDA.n1846 175.546
R1943 GNDA.n1887 GNDA.n408 175.546
R1944 GNDA.n2132 GNDA.n408 175.546
R1945 GNDA.n2122 GNDA.n2008 175.546
R1946 GNDA.n2043 GNDA.n2013 175.546
R1947 GNDA.n2047 GNDA.n2046 175.546
R1948 GNDA.n2056 GNDA.n2055 175.546
R1949 GNDA.n2063 GNDA.n2062 175.546
R1950 GNDA.n2004 GNDA.n428 175.546
R1951 GNDA.n434 GNDA.n433 175.546
R1952 GNDA.n440 GNDA.n436 175.546
R1953 GNDA.n443 GNDA.n442 175.546
R1954 GNDA.n449 GNDA.n445 175.546
R1955 GNDA.n1978 GNDA.n453 175.546
R1956 GNDA.n1978 GNDA.n1968 175.546
R1957 GNDA.n1974 GNDA.n1968 175.546
R1958 GNDA.n1974 GNDA.n1971 175.546
R1959 GNDA.n1971 GNDA.n8 175.546
R1960 GNDA.n2507 GNDA.n8 175.546
R1961 GNDA.n2507 GNDA.n9 175.546
R1962 GNDA.n2503 GNDA.n9 175.546
R1963 GNDA.n2503 GNDA.n11 175.546
R1964 GNDA.n2499 GNDA.n11 175.546
R1965 GNDA.n2499 GNDA.n2496 175.546
R1966 GNDA.n2385 GNDA.n2384 175.546
R1967 GNDA.n2382 GNDA.n196 175.546
R1968 GNDA.n2378 GNDA.n2377 175.546
R1969 GNDA.n2375 GNDA.n202 175.546
R1970 GNDA.n2371 GNDA.n2370 175.546
R1971 GNDA.n2488 GNDA.n17 175.546
R1972 GNDA.n2488 GNDA.n19 175.546
R1973 GNDA.n2484 GNDA.n19 175.546
R1974 GNDA.n2484 GNDA.n22 175.546
R1975 GNDA.n2480 GNDA.n22 175.546
R1976 GNDA.n2480 GNDA.n23 175.546
R1977 GNDA.n2476 GNDA.n23 175.546
R1978 GNDA.n2476 GNDA.n25 175.546
R1979 GNDA.n2472 GNDA.n25 175.546
R1980 GNDA.n2472 GNDA.n28 175.546
R1981 GNDA.n2468 GNDA.n28 175.546
R1982 GNDA.n2447 GNDA.n39 175.546
R1983 GNDA.n2447 GNDA.n37 175.546
R1984 GNDA.n2452 GNDA.n37 175.546
R1985 GNDA.n2452 GNDA.n35 175.546
R1986 GNDA.n2456 GNDA.n35 175.546
R1987 GNDA.n2456 GNDA.n34 175.546
R1988 GNDA.n2460 GNDA.n34 175.546
R1989 GNDA.n2460 GNDA.n32 175.546
R1990 GNDA.n2464 GNDA.n32 175.546
R1991 GNDA.n2464 GNDA.n30 175.546
R1992 GNDA.n186 GNDA.n185 175.546
R1993 GNDA.n107 GNDA.n103 175.546
R1994 GNDA.n111 GNDA.n109 175.546
R1995 GNDA.n122 GNDA.n97 175.546
R1996 GNDA.n126 GNDA.n124 175.546
R1997 GNDA.n2360 GNDA.n2359 175.546
R1998 GNDA.n198 GNDA.n197 175.546
R1999 GNDA.n2363 GNDA.n199 175.546
R2000 GNDA.n204 GNDA.n203 175.546
R2001 GNDA.n2368 GNDA.n205 175.546
R2002 GNDA.n419 GNDA.n418 175.546
R2003 GNDA.n398 GNDA.n397 175.546
R2004 GNDA.n422 GNDA.n399 175.546
R2005 GNDA.n404 GNDA.n403 175.546
R2006 GNDA.n425 GNDA.n405 175.546
R2007 GNDA.n2305 GNDA.n2304 175.546
R2008 GNDA.n2309 GNDA.n2308 175.546
R2009 GNDA.n2313 GNDA.n2312 175.546
R2010 GNDA.n2315 GNDA.n369 175.546
R2011 GNDA.n2320 GNDA.n364 175.546
R2012 GNDA.n2344 GNDA.n2343 175.546
R2013 GNDA.n2341 GNDA.n350 175.546
R2014 GNDA.n2337 GNDA.n2336 175.546
R2015 GNDA.n2334 GNDA.n357 175.546
R2016 GNDA.n2330 GNDA.n2329 175.546
R2017 GNDA.n2157 GNDA.n388 175.546
R2018 GNDA.n2187 GNDA.n2186 175.546
R2019 GNDA.n2194 GNDA.n2193 175.546
R2020 GNDA.n2201 GNDA.n2200 175.546
R2021 GNDA.n2257 GNDA.n2256 175.546
R2022 GNDA.n1158 GNDA.n1157 175.546
R2023 GNDA.n1163 GNDA.n1162 175.546
R2024 GNDA.n1165 GNDA.n1164 175.546
R2025 GNDA.n1170 GNDA.n1169 175.546
R2026 GNDA.n1171 GNDA.n217 175.546
R2027 GNDA.n1098 GNDA.n1095 175.546
R2028 GNDA.n1102 GNDA.n1100 175.546
R2029 GNDA.n1106 GNDA.n1091 175.546
R2030 GNDA.n1110 GNDA.n1108 175.546
R2031 GNDA.n1114 GNDA.n1089 175.546
R2032 GNDA.n1137 GNDA.n1078 175.546
R2033 GNDA.n1133 GNDA.n1078 175.546
R2034 GNDA.n1133 GNDA.n1081 175.546
R2035 GNDA.n1129 GNDA.n1081 175.546
R2036 GNDA.n1129 GNDA.n1127 175.546
R2037 GNDA.n1127 GNDA.n1083 175.546
R2038 GNDA.n1123 GNDA.n1083 175.546
R2039 GNDA.n1123 GNDA.n1085 175.546
R2040 GNDA.n1119 GNDA.n1085 175.546
R2041 GNDA.n1119 GNDA.n1117 175.546
R2042 GNDA.n1152 GNDA.n971 175.546
R2043 GNDA.n1061 GNDA.n1052 175.546
R2044 GNDA.n1065 GNDA.n1063 175.546
R2045 GNDA.n1073 GNDA.n1047 175.546
R2046 GNDA.n1143 GNDA.n1075 175.546
R2047 GNDA.n1273 GNDA.n1270 175.546
R2048 GNDA.n1270 GNDA.n1269 175.546
R2049 GNDA.n1269 GNDA.n1247 175.546
R2050 GNDA.n1265 GNDA.n1247 175.546
R2051 GNDA.n1265 GNDA.n1249 175.546
R2052 GNDA.n1261 GNDA.n1249 175.546
R2053 GNDA.n1261 GNDA.n1251 175.546
R2054 GNDA.n1257 GNDA.n1251 175.546
R2055 GNDA.n1257 GNDA.n1254 175.546
R2056 GNDA.n1254 GNDA.n1240 175.546
R2057 GNDA.n1391 GNDA.n1277 175.546
R2058 GNDA.n1313 GNDA.n1279 175.546
R2059 GNDA.n1316 GNDA.n1313 175.546
R2060 GNDA.n1316 GNDA.n1305 175.546
R2061 GNDA.n1327 GNDA.n1305 175.546
R2062 GNDA.n1327 GNDA.n1303 175.546
R2063 GNDA.n1331 GNDA.n1303 175.546
R2064 GNDA.n1331 GNDA.n858 175.546
R2065 GNDA.n1455 GNDA.n858 175.546
R2066 GNDA.n1450 GNDA.n1449 175.546
R2067 GNDA.n1447 GNDA.n1213 175.546
R2068 GNDA.n1443 GNDA.n1442 175.546
R2069 GNDA.n1440 GNDA.n1222 175.546
R2070 GNDA.n1436 GNDA.n1435 175.546
R2071 GNDA.n1413 GNDA.n1412 175.546
R2072 GNDA.n1417 GNDA.n1416 175.546
R2073 GNDA.n1421 GNDA.n1420 175.546
R2074 GNDA.n1423 GNDA.n1238 175.546
R2075 GNDA.n1428 GNDA.n1233 175.546
R2076 GNDA.n2271 GNDA.n2270 173.881
R2077 GNDA.n2124 GNDA.t238 172.876
R2078 GNDA.n1686 GNDA.t229 172.876
R2079 GNDA.n2322 GNDA.t238 172.615
R2080 GNDA.n1430 GNDA.t229 172.615
R2081 GNDA.n718 GNDA.n717 171.817
R2082 GNDA.n2272 GNDA.n2271 171.624
R2083 GNDA.n1278 GNDA.n1242 170.543
R2084 GNDA.t229 GNDA.n1263 165.044
R2085 GNDA.n1916 GNDA.t229 165.044
R2086 GNDA.n1752 GNDA.t229 165.044
R2087 GNDA.n713 GNDA.n712 164.906
R2088 GNDA.n334 GNDA.n333 163.333
R2089 GNDA.n1201 GNDA.n866 163.333
R2090 GNDA.n1386 GNDA.n1385 163.333
R2091 GNDA.n2117 GNDA.n2116 163.333
R2092 GNDA.n180 GNDA.n179 163.333
R2093 GNDA.n1896 GNDA.n1772 163.333
R2094 GNDA.n2263 GNDA.n2159 163.333
R2095 GNDA.n1679 GNDA.n1678 163.333
R2096 GNDA.n1149 GNDA.n974 163.333
R2097 GNDA.n1948 GNDA.t229 162.964
R2098 GNDA.n2481 GNDA.t238 162.964
R2099 GNDA.t251 GNDA.n561 162.857
R2100 GNDA.n560 GNDA.t241 162.857
R2101 GNDA.n1467 GNDA.t284 160.725
R2102 GNDA.n1466 GNDA.t277 160.725
R2103 GNDA.n1462 GNDA.t315 160.725
R2104 GNDA.n1463 GNDA.t297 160.725
R2105 GNDA.n1477 GNDA.t227 160.725
R2106 GNDA.n1470 GNDA.t280 160.725
R2107 GNDA.n768 GNDA.n530 160
R2108 GNDA.n538 GNDA.n537 160
R2109 GNDA.n761 GNDA.n760 160
R2110 GNDA.n824 GNDA.t21 157.555
R2111 GNDA.n823 GNDA.t12 157.555
R2112 GNDA.n734 GNDA.n733 156.8
R2113 GNDA.n544 GNDA.n521 153.601
R2114 GNDA.n707 GNDA.n706 153.601
R2115 GNDA.n514 GNDA.n508 153.601
R2116 GNDA.n651 GNDA.n598 153.601
R2117 GNDA.n847 GNDA.t176 153.294
R2118 GNDA.n645 GNDA.t270 152.994
R2119 GNDA.n643 GNDA.t260 152.994
R2120 GNDA.n504 GNDA.t263 152.994
R2121 GNDA.n800 GNDA.t254 152.994
R2122 GNDA.n1264 GNDA.t229 150.999
R2123 GNDA.t229 GNDA.n1695 150.999
R2124 GNDA.t229 GNDA.n1719 150.999
R2125 GNDA.n710 GNDA.n709 150.4
R2126 GNDA.n737 GNDA.n736 150.4
R2127 GNDA.n336 GNDA.n231 150
R2128 GNDA.n268 GNDA.n255 150
R2129 GNDA.n272 GNDA.n270 150
R2130 GNDA.n283 GNDA.n248 150
R2131 GNDA.n331 GNDA.n232 150
R2132 GNDA.n327 GNDA.n325 150
R2133 GNDA.n323 GNDA.n234 150
R2134 GNDA.n319 GNDA.n317 150
R2135 GNDA.n315 GNDA.n236 150
R2136 GNDA.n311 GNDA.n310 150
R2137 GNDA.n308 GNDA.n239 150
R2138 GNDA.n304 GNDA.n303 150
R2139 GNDA.n286 GNDA.n285 150
R2140 GNDA.n288 GNDA.n286 150
R2141 GNDA.n292 GNDA.n245 150
R2142 GNDA.n295 GNDA.n294 150
R2143 GNDA.n297 GNDA.n242 150
R2144 GNDA.n947 GNDA.n867 150
R2145 GNDA.n950 GNDA.n949 150
R2146 GNDA.n961 GNDA.n960 150
R2147 GNDA.n1198 GNDA.n886 150
R2148 GNDA.n891 GNDA.n890 150
R2149 GNDA.n895 GNDA.n894 150
R2150 GNDA.n899 GNDA.n898 150
R2151 GNDA.n903 GNDA.n902 150
R2152 GNDA.n907 GNDA.n906 150
R2153 GNDA.n911 GNDA.n910 150
R2154 GNDA.n915 GNDA.n914 150
R2155 GNDA.n919 GNDA.n918 150
R2156 GNDA.n885 GNDA.n881 150
R2157 GNDA.n934 GNDA.n881 150
R2158 GNDA.n932 GNDA.n931 150
R2159 GNDA.n928 GNDA.n927 150
R2160 GNDA.n924 GNDA.n876 150
R2161 GNDA.n1388 GNDA.n1283 150
R2162 GNDA.n1320 GNDA.n1309 150
R2163 GNDA.n1324 GNDA.n1322 150
R2164 GNDA.n1335 GNDA.n1301 150
R2165 GNDA.n1382 GNDA.n1381 150
R2166 GNDA.n1379 GNDA.n1286 150
R2167 GNDA.n1375 GNDA.n1373 150
R2168 GNDA.n1370 GNDA.n1369 150
R2169 GNDA.n1367 GNDA.n1289 150
R2170 GNDA.n1363 GNDA.n1362 150
R2171 GNDA.n1360 GNDA.n1292 150
R2172 GNDA.n1356 GNDA.n1355 150
R2173 GNDA.n1338 GNDA.n1337 150
R2174 GNDA.n1340 GNDA.n1338 150
R2175 GNDA.n1344 GNDA.n1298 150
R2176 GNDA.n1347 GNDA.n1346 150
R2177 GNDA.n1349 GNDA.n1295 150
R2178 GNDA.n2119 GNDA.n2017 150
R2179 GNDA.n2050 GNDA.n2041 150
R2180 GNDA.n2052 GNDA.n2039 150
R2181 GNDA.n2066 GNDA.n2035 150
R2182 GNDA.n2113 GNDA.n2112 150
R2183 GNDA.n2110 GNDA.n2020 150
R2184 GNDA.n2106 GNDA.n2104 150
R2185 GNDA.n2101 GNDA.n2100 150
R2186 GNDA.n2098 GNDA.n2023 150
R2187 GNDA.n2094 GNDA.n2093 150
R2188 GNDA.n2091 GNDA.n2026 150
R2189 GNDA.n2087 GNDA.n2086 150
R2190 GNDA.n2069 GNDA.n2068 150
R2191 GNDA.n2071 GNDA.n2069 150
R2192 GNDA.n2075 GNDA.n2032 150
R2193 GNDA.n2078 GNDA.n2077 150
R2194 GNDA.n2080 GNDA.n2029 150
R2195 GNDA.n182 GNDA.n77 150
R2196 GNDA.n114 GNDA.n101 150
R2197 GNDA.n118 GNDA.n116 150
R2198 GNDA.n129 GNDA.n94 150
R2199 GNDA.n177 GNDA.n78 150
R2200 GNDA.n173 GNDA.n171 150
R2201 GNDA.n169 GNDA.n80 150
R2202 GNDA.n165 GNDA.n163 150
R2203 GNDA.n161 GNDA.n82 150
R2204 GNDA.n157 GNDA.n156 150
R2205 GNDA.n154 GNDA.n85 150
R2206 GNDA.n150 GNDA.n149 150
R2207 GNDA.n132 GNDA.n131 150
R2208 GNDA.n134 GNDA.n132 150
R2209 GNDA.n138 GNDA.n91 150
R2210 GNDA.n141 GNDA.n140 150
R2211 GNDA.n143 GNDA.n88 150
R2212 GNDA.n1852 GNDA.n1773 150
R2213 GNDA.n1871 GNDA.n1870 150
R2214 GNDA.n1877 GNDA.n1876 150
R2215 GNDA.n1893 GNDA.n1842 150
R2216 GNDA.n1794 GNDA.n1793 150
R2217 GNDA.n1798 GNDA.n1797 150
R2218 GNDA.n1802 GNDA.n1801 150
R2219 GNDA.n1806 GNDA.n1805 150
R2220 GNDA.n1810 GNDA.n1809 150
R2221 GNDA.n1814 GNDA.n1813 150
R2222 GNDA.n1818 GNDA.n1817 150
R2223 GNDA.n1822 GNDA.n1821 150
R2224 GNDA.n1841 GNDA.n1787 150
R2225 GNDA.n1837 GNDA.n1787 150
R2226 GNDA.n1835 GNDA.n1834 150
R2227 GNDA.n1831 GNDA.n1830 150
R2228 GNDA.n1827 GNDA.n1782 150
R2229 GNDA.n2182 GNDA.n2160 150
R2230 GNDA.n2190 GNDA.n2189 150
R2231 GNDA.n2197 GNDA.n2196 150
R2232 GNDA.n2260 GNDA.n2179 150
R2233 GNDA.n2207 GNDA.n2206 150
R2234 GNDA.n2211 GNDA.n2210 150
R2235 GNDA.n2215 GNDA.n2214 150
R2236 GNDA.n2219 GNDA.n2218 150
R2237 GNDA.n2223 GNDA.n2222 150
R2238 GNDA.n2227 GNDA.n2226 150
R2239 GNDA.n2231 GNDA.n2230 150
R2240 GNDA.n2235 GNDA.n2234 150
R2241 GNDA.n2178 GNDA.n2174 150
R2242 GNDA.n2250 GNDA.n2174 150
R2243 GNDA.n2248 GNDA.n2247 150
R2244 GNDA.n2244 GNDA.n2243 150
R2245 GNDA.n2240 GNDA.n2169 150
R2246 GNDA.n1681 GNDA.n1580 150
R2247 GNDA.n1613 GNDA.n1604 150
R2248 GNDA.n1615 GNDA.n1602 150
R2249 GNDA.n1628 GNDA.n1598 150
R2250 GNDA.n1675 GNDA.n1674 150
R2251 GNDA.n1672 GNDA.n1583 150
R2252 GNDA.n1668 GNDA.n1666 150
R2253 GNDA.n1663 GNDA.n1662 150
R2254 GNDA.n1660 GNDA.n1586 150
R2255 GNDA.n1656 GNDA.n1655 150
R2256 GNDA.n1653 GNDA.n1589 150
R2257 GNDA.n1649 GNDA.n1648 150
R2258 GNDA.n1631 GNDA.n1630 150
R2259 GNDA.n1633 GNDA.n1631 150
R2260 GNDA.n1637 GNDA.n1595 150
R2261 GNDA.n1640 GNDA.n1639 150
R2262 GNDA.n1642 GNDA.n1592 150
R2263 GNDA.n1055 GNDA.n975 150
R2264 GNDA.n1058 GNDA.n1057 150
R2265 GNDA.n1069 GNDA.n1068 150
R2266 GNDA.n1146 GNDA.n994 150
R2267 GNDA.n999 GNDA.n998 150
R2268 GNDA.n1003 GNDA.n1002 150
R2269 GNDA.n1007 GNDA.n1006 150
R2270 GNDA.n1011 GNDA.n1010 150
R2271 GNDA.n1015 GNDA.n1014 150
R2272 GNDA.n1019 GNDA.n1018 150
R2273 GNDA.n1023 GNDA.n1022 150
R2274 GNDA.n1027 GNDA.n1026 150
R2275 GNDA.n993 GNDA.n989 150
R2276 GNDA.n1042 GNDA.n989 150
R2277 GNDA.n1040 GNDA.n1039 150
R2278 GNDA.n1036 GNDA.n1035 150
R2279 GNDA.n1032 GNDA.n984 150
R2280 GNDA.n1499 GNDA.n1498 149.181
R2281 GNDA.n825 GNDA.t106 148.906
R2282 GNDA.n825 GNDA.t182 148.653
R2283 GNDA.n618 GNDA.n617 148.38
R2284 GNDA.n617 GNDA.n563 148.38
R2285 GNDA.n1552 GNDA.t149 141.583
R2286 GNDA.t138 GNDA.t104 140.464
R2287 GNDA.n829 GNDA.n827 140.077
R2288 GNDA.n845 GNDA.n844 139.077
R2289 GNDA.n843 GNDA.n842 139.077
R2290 GNDA.n841 GNDA.n840 139.077
R2291 GNDA.n839 GNDA.n838 139.077
R2292 GNDA.n837 GNDA.n836 139.077
R2293 GNDA.n835 GNDA.n834 139.077
R2294 GNDA.n833 GNDA.n832 139.077
R2295 GNDA.n831 GNDA.n830 139.077
R2296 GNDA.n829 GNDA.n828 139.077
R2297 GNDA.n677 GNDA.n676 139.077
R2298 GNDA.t20 GNDA.t181 137.016
R2299 GNDA.n1930 GNDA.n1929 133.44
R2300 GNDA.t226 GNDA.n1482 131.625
R2301 GNDA.t314 GNDA.n1533 131.625
R2302 GNDA.n602 GNDA.t269 130.731
R2303 GNDA.n715 GNDA.t253 130.731
R2304 GNDA.n727 GNDA.n726 127.249
R2305 GNDA.n2395 GNDA.n68 126.782
R2306 GNDA.n2298 GNDA.n377 126.782
R2307 GNDA.n1941 GNDA.n464 126.782
R2308 GNDA.n1905 GNDA.n1706 126.782
R2309 GNDA.n1982 GNDA.n453 126.782
R2310 GNDA.n2492 GNDA.n17 126.782
R2311 GNDA.n2301 GNDA.n2300 126.782
R2312 GNDA.n1093 GNDA.n218 126.782
R2313 GNDA.n1409 GNDA.n1408 126.782
R2314 GNDA.n2349 GNDA.n344 124.832
R2315 GNDA.n1207 GNDA.n1206 124.832
R2316 GNDA.n1714 GNDA.n1711 124.832
R2317 GNDA.n1688 GNDA.n1569 124.832
R2318 GNDA.n2126 GNDA.n2007 124.832
R2319 GNDA.n2390 GNDA.n190 124.832
R2320 GNDA.n2268 GNDA.n389 124.832
R2321 GNDA.n1155 GNDA.n1154 124.832
R2322 GNDA.n1395 GNDA.n1244 124.832
R2323 GNDA.n631 GNDA.n630 121.6
R2324 GNDA.n807 GNDA.n503 121.6
R2325 GNDA.n642 GNDA.n641 119.525
R2326 GNDA.n799 GNDA.n510 119.525
R2327 GNDA.n1531 GNDA.n1530 118.4
R2328 GNDA.n1528 GNDA.n1527 118.4
R2329 GNDA.n1526 GNDA.n1509 118.4
R2330 GNDA.n1507 GNDA.n1506 118.4
R2331 GNDA.n1480 GNDA.n1479 118.4
R2332 GNDA.n1505 GNDA.n1471 118.4
R2333 GNDA.n1744 GNDA.n1743 115.882
R2334 GNDA.n626 GNDA.t13 115.79
R2335 GNDA.n640 GNDA.t54 115.79
R2336 GNDA.n529 GNDA.t323 113.974
R2337 GNDA.n533 GNDA.t300 113.974
R2338 GNDA.n532 GNDA.t318 113.974
R2339 GNDA.n531 GNDA.t294 113.974
R2340 GNDA.n543 GNDA.t326 113.974
R2341 GNDA.n542 GNDA.t306 113.974
R2342 GNDA.n541 GNDA.t287 113.974
R2343 GNDA.n539 GNDA.t248 113.974
R2344 GNDA.n758 GNDA.t236 113.974
R2345 GNDA.n757 GNDA.t312 113.974
R2346 GNDA.n1315 GNDA.t229 113.624
R2347 GNDA.t173 GNDA.t166 112.822
R2348 GNDA.t199 GNDA.t223 112.822
R2349 GNDA.t223 GNDA.t114 112.822
R2350 GNDA.t101 GNDA.t36 112.822
R2351 GNDA.t353 GNDA.t101 112.822
R2352 GNDA.t219 GNDA.t217 112.822
R2353 GNDA.n2512 GNDA.t238 112.388
R2354 GNDA.n634 GNDA.n633 112.055
R2355 GNDA.t105 GNDA.t95 109.612
R2356 GNDA.n754 GNDA.n553 108.8
R2357 GNDA.n742 GNDA.n556 108.8
R2358 GNDA.t169 GNDA.n1483 106.553
R2359 GNDA.n1406 GNDA.t229 105.347
R2360 GNDA.n2366 GNDA.n0 14.555
R2361 GNDA.n731 GNDA.t311 101.194
R2362 GNDA.n1514 GNDA.t72 100.285
R2363 GNDA.n1966 GNDA.n394 99.6276
R2364 GNDA.n700 GNDA.n699 99.0842
R2365 GNDA.n698 GNDA.n697 99.0842
R2366 GNDA.n696 GNDA.n695 99.0842
R2367 GNDA.n694 GNDA.n693 99.0842
R2368 GNDA.n692 GNDA.n691 99.0842
R2369 GNDA.n690 GNDA.n689 99.0842
R2370 GNDA.n688 GNDA.n687 99.0842
R2371 GNDA.n686 GNDA.n685 99.0842
R2372 GNDA.n684 GNDA.n683 99.0842
R2373 GNDA.n682 GNDA.n681 99.0842
R2374 GNDA.n680 GNDA.n679 99.0842
R2375 GNDA.n585 GNDA.t71 97.1515
R2376 GNDA.n811 GNDA.t44 97.1515
R2377 GNDA.n795 GNDA.n794 95.101
R2378 GNDA.n659 GNDA.n592 95.101
R2379 GNDA.n702 GNDA.t309 94.8842
R2380 GNDA.n591 GNDA.t274 94.8842
R2381 GNDA.t138 GNDA.n474 94.813
R2382 GNDA.n661 GNDA.n660 94.601
R2383 GNDA.n793 GNDA.n792 94.601
R2384 GNDA.n579 GNDA.n577 94.0176
R2385 GNDA.n1136 GNDA.n1079 91.8159
R2386 GNDA.n1136 GNDA.n1135 91.8159
R2387 GNDA.n1135 GNDA.n1134 91.8159
R2388 GNDA.n1134 GNDA.n1080 91.8159
R2389 GNDA.n1128 GNDA.n1080 91.8159
R2390 GNDA.n1126 GNDA.n1125 91.8159
R2391 GNDA.n1125 GNDA.n1124 91.8159
R2392 GNDA.n1124 GNDA.n1084 91.8159
R2393 GNDA.n1118 GNDA.n1084 91.8159
R2394 GNDA.n1118 GNDA.n48 91.8159
R2395 GNDA.n2441 GNDA.n49 91.8159
R2396 GNDA.n2435 GNDA.n49 91.8159
R2397 GNDA.n2435 GNDA.n2434 91.8159
R2398 GNDA.n2434 GNDA.n2433 91.8159
R2399 GNDA.n2433 GNDA.n55 91.8159
R2400 GNDA.n2427 GNDA.n2426 91.8159
R2401 GNDA.n2426 GNDA.n2425 91.8159
R2402 GNDA.n2425 GNDA.n59 91.8159
R2403 GNDA.n2419 GNDA.n59 91.8159
R2404 GNDA.n2419 GNDA.n43 91.8159
R2405 GNDA.n2442 GNDA.n38 91.8159
R2406 GNDA.n2448 GNDA.n38 91.8159
R2407 GNDA.n2449 GNDA.n2448 91.8159
R2408 GNDA.n2451 GNDA.n2449 91.8159
R2409 GNDA.n2451 GNDA.n2450 91.8159
R2410 GNDA.n2458 GNDA.n2457 91.8159
R2411 GNDA.n2459 GNDA.n2458 91.8159
R2412 GNDA.n2459 GNDA.n31 91.8159
R2413 GNDA.n2465 GNDA.n31 91.8159
R2414 GNDA.n2466 GNDA.n2465 91.8159
R2415 GNDA.n1559 GNDA.n483 91.3437
R2416 GNDA.n624 GNDA.n613 91.3105
R2417 GNDA.n731 GNDA.n727 89.9494
R2418 GNDA.t13 GNDA.t161 89.644
R2419 GNDA.t14 GNDA.t15 89.644
R2420 GNDA.n1484 GNDA.t226 87.7498
R2421 GNDA.n1534 GNDA.t314 87.7498
R2422 GNDA.n1538 GNDA.n850 85.2842
R2423 GNDA.n1491 GNDA.n1490 85.2842
R2424 GNDA.n2513 GNDA.n4 84.306
R2425 GNDA.n1457 GNDA.n394 83.2184
R2426 GNDA.t42 GNDA.t259 82.1737
R2427 GNDA.t4 GNDA.t141 82.1737
R2428 GNDA.t131 GNDA.t139 82.1737
R2429 GNDA.t132 GNDA.t134 82.1737
R2430 GNDA.t178 GNDA.t146 82.1737
R2431 GNDA.t184 GNDA.t0 82.1737
R2432 GNDA.t19 GNDA.t144 82.1737
R2433 GNDA.t209 GNDA.t262 82.1737
R2434 GNDA.n2131 GNDA.t229 80.9821
R2435 GNDA.t290 GNDA.t69 78.4385
R2436 GNDA.t231 GNDA.t145 78.4385
R2437 GNDA.n2271 GNDA.t238 76.3879
R2438 GNDA.n2397 GNDA.n2396 76.3222
R2439 GNDA.n2398 GNDA.n66 76.3222
R2440 GNDA.n2405 GNDA.n2404 76.3222
R2441 GNDA.n2406 GNDA.n64 76.3222
R2442 GNDA.n2413 GNDA.n2412 76.3222
R2443 GNDA.n2417 GNDA.n62 76.3222
R2444 GNDA.n2440 GNDA.n2439 76.3222
R2445 GNDA.n344 GNDA.n226 76.3222
R2446 GNDA.n339 GNDA.n229 76.3222
R2447 GNDA.n262 GNDA.n261 76.3222
R2448 GNDA.n265 GNDA.n264 76.3222
R2449 GNDA.n277 GNDA.n276 76.3222
R2450 GNDA.n280 GNDA.n279 76.3222
R2451 GNDA.n2348 GNDA.n206 76.3222
R2452 GNDA.n348 GNDA.n207 76.3222
R2453 GNDA.n352 GNDA.n208 76.3222
R2454 GNDA.n354 GNDA.n209 76.3222
R2455 GNDA.n359 GNDA.n210 76.3222
R2456 GNDA.n2325 GNDA.n211 76.3222
R2457 GNDA.n1210 GNDA.n1209 76.3222
R2458 GNDA.n1216 GNDA.n1215 76.3222
R2459 GNDA.n1219 GNDA.n1218 76.3222
R2460 GNDA.n1225 GNDA.n1224 76.3222
R2461 GNDA.n1228 GNDA.n1227 76.3222
R2462 GNDA.n1229 GNDA.n376 76.3222
R2463 GNDA.n2293 GNDA.n382 76.3222
R2464 GNDA.n2291 GNDA.n2290 76.3222
R2465 GNDA.n2286 GNDA.n2275 76.3222
R2466 GNDA.n2284 GNDA.n2283 76.3222
R2467 GNDA.n2279 GNDA.n2277 76.3222
R2468 GNDA.n2354 GNDA.n222 76.3222
R2469 GNDA.n1188 GNDA.n1160 76.3222
R2470 GNDA.n1186 GNDA.n1185 76.3222
R2471 GNDA.n1181 GNDA.n1167 76.3222
R2472 GNDA.n1179 GNDA.n1178 76.3222
R2473 GNDA.n1174 GNDA.n1172 76.3222
R2474 GNDA.n2355 GNDA.n221 76.3222
R2475 GNDA.n1206 GNDA.n1205 76.3222
R2476 GNDA.n943 GNDA.n863 76.3222
R2477 GNDA.n954 GNDA.n953 76.3222
R2478 GNDA.n957 GNDA.n956 76.3222
R2479 GNDA.n966 GNDA.n965 76.3222
R2480 GNDA.n1195 GNDA.n1194 76.3222
R2481 GNDA.n1763 GNDA.n1762 76.3222
R2482 GNDA.n2002 GNDA.n430 76.3222
R2483 GNDA.n2000 GNDA.n1999 76.3222
R2484 GNDA.n1995 GNDA.n438 76.3222
R2485 GNDA.n1993 GNDA.n1992 76.3222
R2486 GNDA.n1988 GNDA.n447 76.3222
R2487 GNDA.n1986 GNDA.n1985 76.3222
R2488 GNDA.n1927 GNDA.n1926 76.3222
R2489 GNDA.n1688 GNDA.n1687 76.3222
R2490 GNDA.n1685 GNDA.n1684 76.3222
R2491 GNDA.n1606 GNDA.n1575 76.3222
R2492 GNDA.n1609 GNDA.n1574 76.3222
R2493 GNDA.n1619 GNDA.n1573 76.3222
R2494 GNDA.n1625 GNDA.n1572 76.3222
R2495 GNDA.n2152 GNDA.n2151 76.3222
R2496 GNDA.n2149 GNDA.n2148 76.3222
R2497 GNDA.n2144 GNDA.n401 76.3222
R2498 GNDA.n2142 GNDA.n2141 76.3222
R2499 GNDA.n2137 GNDA.n407 76.3222
R2500 GNDA.n2135 GNDA.n2134 76.3222
R2501 GNDA.n2126 GNDA.n2125 76.3222
R2502 GNDA.n2123 GNDA.n2122 76.3222
R2503 GNDA.n2043 GNDA.n2012 76.3222
R2504 GNDA.n2046 GNDA.n2011 76.3222
R2505 GNDA.n2056 GNDA.n2010 76.3222
R2506 GNDA.n2063 GNDA.n2009 76.3222
R2507 GNDA.n2005 GNDA.n2004 76.3222
R2508 GNDA.n433 GNDA.n432 76.3222
R2509 GNDA.n436 GNDA.n435 76.3222
R2510 GNDA.n442 GNDA.n441 76.3222
R2511 GNDA.n445 GNDA.n444 76.3222
R2512 GNDA.n451 GNDA.n450 76.3222
R2513 GNDA.n2386 GNDA.n2385 76.3222
R2514 GNDA.n2383 GNDA.n2382 76.3222
R2515 GNDA.n2378 GNDA.n201 76.3222
R2516 GNDA.n2376 GNDA.n2375 76.3222
R2517 GNDA.n2371 GNDA.n2369 76.3222
R2518 GNDA.n2495 GNDA.n13 76.3222
R2519 GNDA.n2444 GNDA.n39 76.3222
R2520 GNDA.n190 GNDA.n72 76.3222
R2521 GNDA.n185 GNDA.n75 76.3222
R2522 GNDA.n108 GNDA.n107 76.3222
R2523 GNDA.n111 GNDA.n110 76.3222
R2524 GNDA.n123 GNDA.n122 76.3222
R2525 GNDA.n126 GNDA.n125 76.3222
R2526 GNDA.n2389 GNDA.n191 76.3222
R2527 GNDA.n2361 GNDA.n2360 76.3222
R2528 GNDA.n2362 GNDA.n198 76.3222
R2529 GNDA.n2364 GNDA.n2363 76.3222
R2530 GNDA.n2367 GNDA.n204 76.3222
R2531 GNDA.n2365 GNDA.n205 76.3222
R2532 GNDA.n2365 GNDA.n15 76.3222
R2533 GNDA.n2368 GNDA.n2367 76.3222
R2534 GNDA.n2364 GNDA.n203 76.3222
R2535 GNDA.n2362 GNDA.n199 76.3222
R2536 GNDA.n2361 GNDA.n197 76.3222
R2537 GNDA.n2359 GNDA.n191 76.3222
R2538 GNDA.n2370 GNDA.n13 76.3222
R2539 GNDA.n2369 GNDA.n202 76.3222
R2540 GNDA.n2377 GNDA.n2376 76.3222
R2541 GNDA.n201 GNDA.n196 76.3222
R2542 GNDA.n2384 GNDA.n2383 76.3222
R2543 GNDA.n2387 GNDA.n2386 76.3222
R2544 GNDA.n2125 GNDA.n2008 76.3222
R2545 GNDA.n2123 GNDA.n2013 76.3222
R2546 GNDA.n2047 GNDA.n2012 76.3222
R2547 GNDA.n2055 GNDA.n2011 76.3222
R2548 GNDA.n2062 GNDA.n2010 76.3222
R2549 GNDA.n2009 GNDA.n193 76.3222
R2550 GNDA.n418 GNDA.n417 76.3222
R2551 GNDA.n420 GNDA.n397 76.3222
R2552 GNDA.n421 GNDA.n399 76.3222
R2553 GNDA.n423 GNDA.n403 76.3222
R2554 GNDA.n424 GNDA.n405 76.3222
R2555 GNDA.n426 GNDA.n371 76.3222
R2556 GNDA.n2301 GNDA.n365 76.3222
R2557 GNDA.n2305 GNDA.n366 76.3222
R2558 GNDA.n2309 GNDA.n367 76.3222
R2559 GNDA.n2313 GNDA.n368 76.3222
R2560 GNDA.n2321 GNDA.n369 76.3222
R2561 GNDA.n2323 GNDA.n364 76.3222
R2562 GNDA.n2324 GNDA.n2323 76.3222
R2563 GNDA.n2321 GNDA.n2320 76.3222
R2564 GNDA.n2315 GNDA.n368 76.3222
R2565 GNDA.n2312 GNDA.n367 76.3222
R2566 GNDA.n2308 GNDA.n366 76.3222
R2567 GNDA.n2304 GNDA.n365 76.3222
R2568 GNDA.n2345 GNDA.n2344 76.3222
R2569 GNDA.n2342 GNDA.n2341 76.3222
R2570 GNDA.n2337 GNDA.n356 76.3222
R2571 GNDA.n2335 GNDA.n2334 76.3222
R2572 GNDA.n2330 GNDA.n363 76.3222
R2573 GNDA.n2328 GNDA.n2327 76.3222
R2574 GNDA.n2269 GNDA.n388 76.3222
R2575 GNDA.n2186 GNDA.n387 76.3222
R2576 GNDA.n2193 GNDA.n386 76.3222
R2577 GNDA.n2200 GNDA.n385 76.3222
R2578 GNDA.n2256 GNDA.n384 76.3222
R2579 GNDA.n383 GNDA.n346 76.3222
R2580 GNDA.n2269 GNDA.n2268 76.3222
R2581 GNDA.n2157 GNDA.n387 76.3222
R2582 GNDA.n2187 GNDA.n386 76.3222
R2583 GNDA.n2194 GNDA.n385 76.3222
R2584 GNDA.n2201 GNDA.n384 76.3222
R2585 GNDA.n2257 GNDA.n383 76.3222
R2586 GNDA.n1156 GNDA.n212 76.3222
R2587 GNDA.n1158 GNDA.n213 76.3222
R2588 GNDA.n1163 GNDA.n214 76.3222
R2589 GNDA.n1165 GNDA.n215 76.3222
R2590 GNDA.n1170 GNDA.n216 76.3222
R2591 GNDA.n2358 GNDA.n217 76.3222
R2592 GNDA.n1094 GNDA.n1093 76.3222
R2593 GNDA.n1099 GNDA.n1098 76.3222
R2594 GNDA.n1102 GNDA.n1101 76.3222
R2595 GNDA.n1107 GNDA.n1106 76.3222
R2596 GNDA.n1110 GNDA.n1109 76.3222
R2597 GNDA.n1115 GNDA.n1114 76.3222
R2598 GNDA.n1138 GNDA.n1137 76.3222
R2599 GNDA.n1154 GNDA.n1153 76.3222
R2600 GNDA.n1051 GNDA.n971 76.3222
R2601 GNDA.n1062 GNDA.n1061 76.3222
R2602 GNDA.n1065 GNDA.n1064 76.3222
R2603 GNDA.n1074 GNDA.n1073 76.3222
R2604 GNDA.n1143 GNDA.n1142 76.3222
R2605 GNDA.n1153 GNDA.n1152 76.3222
R2606 GNDA.n1052 GNDA.n1051 76.3222
R2607 GNDA.n1063 GNDA.n1062 76.3222
R2608 GNDA.n1064 GNDA.n1047 76.3222
R2609 GNDA.n1075 GNDA.n1074 76.3222
R2610 GNDA.n1142 GNDA.n1141 76.3222
R2611 GNDA.n1928 GNDA.n1927 76.3222
R2612 GNDA.n1764 GNDA.n1763 76.3222
R2613 GNDA.n426 GNDA.n425 76.3222
R2614 GNDA.n424 GNDA.n404 76.3222
R2615 GNDA.n423 GNDA.n422 76.3222
R2616 GNDA.n421 GNDA.n398 76.3222
R2617 GNDA.n420 GNDA.n419 76.3222
R2618 GNDA.n417 GNDA.n391 76.3222
R2619 GNDA.n450 GNDA.n449 76.3222
R2620 GNDA.n444 GNDA.n443 76.3222
R2621 GNDA.n441 GNDA.n440 76.3222
R2622 GNDA.n435 GNDA.n434 76.3222
R2623 GNDA.n432 GNDA.n428 76.3222
R2624 GNDA.n2006 GNDA.n2005 76.3222
R2625 GNDA.n2136 GNDA.n2135 76.3222
R2626 GNDA.n407 GNDA.n402 76.3222
R2627 GNDA.n2143 GNDA.n2142 76.3222
R2628 GNDA.n401 GNDA.n396 76.3222
R2629 GNDA.n2150 GNDA.n2149 76.3222
R2630 GNDA.n2153 GNDA.n2152 76.3222
R2631 GNDA.n1987 GNDA.n1986 76.3222
R2632 GNDA.n447 GNDA.n439 76.3222
R2633 GNDA.n1994 GNDA.n1993 76.3222
R2634 GNDA.n438 GNDA.n431 76.3222
R2635 GNDA.n2001 GNDA.n2000 76.3222
R2636 GNDA.n430 GNDA.n412 76.3222
R2637 GNDA.n1687 GNDA.n1571 76.3222
R2638 GNDA.n1685 GNDA.n1576 76.3222
R2639 GNDA.n1610 GNDA.n1575 76.3222
R2640 GNDA.n1618 GNDA.n1574 76.3222
R2641 GNDA.n1624 GNDA.n1573 76.3222
R2642 GNDA.n1572 GNDA.n393 76.3222
R2643 GNDA.n1274 GNDA.n1273 76.3222
R2644 GNDA.n1395 GNDA.n1394 76.3222
R2645 GNDA.n1392 GNDA.n1391 76.3222
R2646 GNDA.n1450 GNDA.n1212 76.3222
R2647 GNDA.n1448 GNDA.n1447 76.3222
R2648 GNDA.n1443 GNDA.n1221 76.3222
R2649 GNDA.n1441 GNDA.n1440 76.3222
R2650 GNDA.n1436 GNDA.n1232 76.3222
R2651 GNDA.n1434 GNDA.n1433 76.3222
R2652 GNDA.n1409 GNDA.n1234 76.3222
R2653 GNDA.n1413 GNDA.n1235 76.3222
R2654 GNDA.n1417 GNDA.n1236 76.3222
R2655 GNDA.n1421 GNDA.n1237 76.3222
R2656 GNDA.n1429 GNDA.n1238 76.3222
R2657 GNDA.n1431 GNDA.n1233 76.3222
R2658 GNDA.n1432 GNDA.n1431 76.3222
R2659 GNDA.n1429 GNDA.n1428 76.3222
R2660 GNDA.n1423 GNDA.n1237 76.3222
R2661 GNDA.n1420 GNDA.n1236 76.3222
R2662 GNDA.n1416 GNDA.n1235 76.3222
R2663 GNDA.n1412 GNDA.n1234 76.3222
R2664 GNDA.n1274 GNDA.n1246 76.3222
R2665 GNDA.n1394 GNDA.n1277 76.3222
R2666 GNDA.n1392 GNDA.n1279 76.3222
R2667 GNDA.n1205 GNDA.n1204 76.3222
R2668 GNDA.n944 GNDA.n943 76.3222
R2669 GNDA.n955 GNDA.n954 76.3222
R2670 GNDA.n956 GNDA.n939 76.3222
R2671 GNDA.n967 GNDA.n966 76.3222
R2672 GNDA.n1194 GNDA.n1193 76.3222
R2673 GNDA.n1230 GNDA.n1229 76.3222
R2674 GNDA.n1227 GNDA.n1226 76.3222
R2675 GNDA.n1224 GNDA.n1223 76.3222
R2676 GNDA.n1218 GNDA.n1217 76.3222
R2677 GNDA.n1215 GNDA.n1214 76.3222
R2678 GNDA.n1209 GNDA.n1208 76.3222
R2679 GNDA.n1435 GNDA.n1434 76.3222
R2680 GNDA.n1232 GNDA.n1222 76.3222
R2681 GNDA.n1442 GNDA.n1441 76.3222
R2682 GNDA.n1221 GNDA.n1213 76.3222
R2683 GNDA.n1449 GNDA.n1448 76.3222
R2684 GNDA.n1212 GNDA.n859 76.3222
R2685 GNDA.n2278 GNDA.n222 76.3222
R2686 GNDA.n2277 GNDA.n2276 76.3222
R2687 GNDA.n2285 GNDA.n2284 76.3222
R2688 GNDA.n2275 GNDA.n2273 76.3222
R2689 GNDA.n2292 GNDA.n2291 76.3222
R2690 GNDA.n382 GNDA.n377 76.3222
R2691 GNDA.n1116 GNDA.n1115 76.3222
R2692 GNDA.n1109 GNDA.n1089 76.3222
R2693 GNDA.n1108 GNDA.n1107 76.3222
R2694 GNDA.n1101 GNDA.n1091 76.3222
R2695 GNDA.n1100 GNDA.n1099 76.3222
R2696 GNDA.n1095 GNDA.n1094 76.3222
R2697 GNDA.n2358 GNDA.n2357 76.3222
R2698 GNDA.n1171 GNDA.n216 76.3222
R2699 GNDA.n1169 GNDA.n215 76.3222
R2700 GNDA.n1164 GNDA.n214 76.3222
R2701 GNDA.n1162 GNDA.n213 76.3222
R2702 GNDA.n1157 GNDA.n212 76.3222
R2703 GNDA.n1173 GNDA.n221 76.3222
R2704 GNDA.n1172 GNDA.n1168 76.3222
R2705 GNDA.n1180 GNDA.n1179 76.3222
R2706 GNDA.n1167 GNDA.n1161 76.3222
R2707 GNDA.n1187 GNDA.n1186 76.3222
R2708 GNDA.n1160 GNDA.n968 76.3222
R2709 GNDA.n361 GNDA.n211 76.3222
R2710 GNDA.n360 GNDA.n210 76.3222
R2711 GNDA.n358 GNDA.n209 76.3222
R2712 GNDA.n353 GNDA.n208 76.3222
R2713 GNDA.n351 GNDA.n207 76.3222
R2714 GNDA.n347 GNDA.n206 76.3222
R2715 GNDA.n2329 GNDA.n2328 76.3222
R2716 GNDA.n363 GNDA.n357 76.3222
R2717 GNDA.n2336 GNDA.n2335 76.3222
R2718 GNDA.n356 GNDA.n350 76.3222
R2719 GNDA.n2343 GNDA.n2342 76.3222
R2720 GNDA.n2346 GNDA.n2345 76.3222
R2721 GNDA.n340 GNDA.n226 76.3222
R2722 GNDA.n257 GNDA.n229 76.3222
R2723 GNDA.n263 GNDA.n262 76.3222
R2724 GNDA.n264 GNDA.n251 76.3222
R2725 GNDA.n278 GNDA.n277 76.3222
R2726 GNDA.n279 GNDA.n50 76.3222
R2727 GNDA.n2414 GNDA.n62 76.3222
R2728 GNDA.n2412 GNDA.n2411 76.3222
R2729 GNDA.n2407 GNDA.n2406 76.3222
R2730 GNDA.n2404 GNDA.n2403 76.3222
R2731 GNDA.n2399 GNDA.n2398 76.3222
R2732 GNDA.n2396 GNDA.n2395 76.3222
R2733 GNDA.n186 GNDA.n72 76.3222
R2734 GNDA.n103 GNDA.n75 76.3222
R2735 GNDA.n109 GNDA.n108 76.3222
R2736 GNDA.n110 GNDA.n97 76.3222
R2737 GNDA.n124 GNDA.n123 76.3222
R2738 GNDA.n125 GNDA.n41 76.3222
R2739 GNDA.n1138 GNDA.n1076 76.3222
R2740 GNDA.n2439 GNDA.n51 76.3222
R2741 GNDA.n2444 GNDA.n2443 76.3222
R2742 GNDA.t150 GNDA.t351 75.2142
R2743 GNDA.t160 GNDA.t44 75.2142
R2744 GNDA.t27 GNDA.t31 75.2142
R2745 GNDA.t107 GNDA.t100 75.2142
R2746 GNDA.t41 GNDA.t45 75.2142
R2747 GNDA.t40 GNDA.t352 75.2142
R2748 GNDA.n284 GNDA.n283 74.5978
R2749 GNDA.n285 GNDA.n284 74.5978
R2750 GNDA.n1199 GNDA.n1198 74.5978
R2751 GNDA.n1199 GNDA.n885 74.5978
R2752 GNDA.n1336 GNDA.n1335 74.5978
R2753 GNDA.n1337 GNDA.n1336 74.5978
R2754 GNDA.n2067 GNDA.n2066 74.5978
R2755 GNDA.n2068 GNDA.n2067 74.5978
R2756 GNDA.n130 GNDA.n129 74.5978
R2757 GNDA.n131 GNDA.n130 74.5978
R2758 GNDA.n1894 GNDA.n1893 74.5978
R2759 GNDA.n1894 GNDA.n1841 74.5978
R2760 GNDA.n2261 GNDA.n2260 74.5978
R2761 GNDA.n2261 GNDA.n2178 74.5978
R2762 GNDA.n1629 GNDA.n1628 74.5978
R2763 GNDA.n1630 GNDA.n1629 74.5978
R2764 GNDA.n1147 GNDA.n1146 74.5978
R2765 GNDA.n1147 GNDA.n993 74.5978
R2766 GNDA.t302 GNDA.t42 70.9682
R2767 GNDA.t69 GNDA.t97 70.9682
R2768 GNDA.t145 GNDA.t2 70.9682
R2769 GNDA.t243 GNDA.t209 70.9682
R2770 GNDA.n1938 GNDA.n465 70.2319
R2771 GNDA.n317 GNDA.n316 69.3109
R2772 GNDA.n316 GNDA.n315 69.3109
R2773 GNDA.n903 GNDA.n875 69.3109
R2774 GNDA.n906 GNDA.n875 69.3109
R2775 GNDA.n1369 GNDA.n1368 69.3109
R2776 GNDA.n1368 GNDA.n1367 69.3109
R2777 GNDA.n2100 GNDA.n2099 69.3109
R2778 GNDA.n2099 GNDA.n2098 69.3109
R2779 GNDA.n163 GNDA.n162 69.3109
R2780 GNDA.n162 GNDA.n161 69.3109
R2781 GNDA.n1806 GNDA.n1781 69.3109
R2782 GNDA.n1809 GNDA.n1781 69.3109
R2783 GNDA.n2219 GNDA.n2168 69.3109
R2784 GNDA.n2222 GNDA.n2168 69.3109
R2785 GNDA.n1662 GNDA.n1661 69.3109
R2786 GNDA.n1661 GNDA.n1660 69.3109
R2787 GNDA.n1011 GNDA.n983 69.3109
R2788 GNDA.n1014 GNDA.n983 69.3109
R2789 GNDA.n296 GNDA.t281 65.8183
R2790 GNDA.n293 GNDA.t281 65.8183
R2791 GNDA.n287 GNDA.t281 65.8183
R2792 GNDA.n302 GNDA.t281 65.8183
R2793 GNDA.n241 GNDA.t281 65.8183
R2794 GNDA.n309 GNDA.t281 65.8183
R2795 GNDA.n238 GNDA.t281 65.8183
R2796 GNDA.n318 GNDA.t281 65.8183
R2797 GNDA.n324 GNDA.t281 65.8183
R2798 GNDA.n326 GNDA.t281 65.8183
R2799 GNDA.n332 GNDA.t281 65.8183
R2800 GNDA.t237 GNDA.n874 65.8183
R2801 GNDA.t237 GNDA.n872 65.8183
R2802 GNDA.t237 GNDA.n870 65.8183
R2803 GNDA.t237 GNDA.n877 65.8183
R2804 GNDA.t237 GNDA.n878 65.8183
R2805 GNDA.t237 GNDA.n879 65.8183
R2806 GNDA.t237 GNDA.n880 65.8183
R2807 GNDA.t237 GNDA.n873 65.8183
R2808 GNDA.t237 GNDA.n871 65.8183
R2809 GNDA.t237 GNDA.n869 65.8183
R2810 GNDA.t237 GNDA.n868 65.8183
R2811 GNDA.n1348 GNDA.t233 65.8183
R2812 GNDA.n1345 GNDA.t233 65.8183
R2813 GNDA.n1339 GNDA.t233 65.8183
R2814 GNDA.n1354 GNDA.t233 65.8183
R2815 GNDA.n1294 GNDA.t233 65.8183
R2816 GNDA.n1361 GNDA.t233 65.8183
R2817 GNDA.n1291 GNDA.t233 65.8183
R2818 GNDA.n1287 GNDA.t233 65.8183
R2819 GNDA.n1374 GNDA.t233 65.8183
R2820 GNDA.n1380 GNDA.t233 65.8183
R2821 GNDA.n1284 GNDA.t233 65.8183
R2822 GNDA.n2079 GNDA.t319 65.8183
R2823 GNDA.n2076 GNDA.t319 65.8183
R2824 GNDA.n2070 GNDA.t319 65.8183
R2825 GNDA.n2085 GNDA.t319 65.8183
R2826 GNDA.n2028 GNDA.t319 65.8183
R2827 GNDA.n2092 GNDA.t319 65.8183
R2828 GNDA.n2025 GNDA.t319 65.8183
R2829 GNDA.n2021 GNDA.t319 65.8183
R2830 GNDA.n2105 GNDA.t319 65.8183
R2831 GNDA.n2111 GNDA.t319 65.8183
R2832 GNDA.n2018 GNDA.t319 65.8183
R2833 GNDA.n142 GNDA.t245 65.8183
R2834 GNDA.n139 GNDA.t245 65.8183
R2835 GNDA.n133 GNDA.t245 65.8183
R2836 GNDA.n148 GNDA.t245 65.8183
R2837 GNDA.n87 GNDA.t245 65.8183
R2838 GNDA.n155 GNDA.t245 65.8183
R2839 GNDA.n84 GNDA.t245 65.8183
R2840 GNDA.n164 GNDA.t245 65.8183
R2841 GNDA.n170 GNDA.t245 65.8183
R2842 GNDA.n172 GNDA.t245 65.8183
R2843 GNDA.n178 GNDA.t245 65.8183
R2844 GNDA.n181 GNDA.t245 65.8183
R2845 GNDA.n100 GNDA.t245 65.8183
R2846 GNDA.n115 GNDA.t245 65.8183
R2847 GNDA.n117 GNDA.t245 65.8183
R2848 GNDA.t320 GNDA.n1780 65.8183
R2849 GNDA.t320 GNDA.n1778 65.8183
R2850 GNDA.t320 GNDA.n1776 65.8183
R2851 GNDA.t320 GNDA.n1783 65.8183
R2852 GNDA.t320 GNDA.n1784 65.8183
R2853 GNDA.t320 GNDA.n1785 65.8183
R2854 GNDA.t320 GNDA.n1786 65.8183
R2855 GNDA.t320 GNDA.n1779 65.8183
R2856 GNDA.t320 GNDA.n1777 65.8183
R2857 GNDA.t320 GNDA.n1775 65.8183
R2858 GNDA.t320 GNDA.n1774 65.8183
R2859 GNDA.n1895 GNDA.t320 65.8183
R2860 GNDA.t320 GNDA.n1788 65.8183
R2861 GNDA.t320 GNDA.n1789 65.8183
R2862 GNDA.t320 GNDA.n1790 65.8183
R2863 GNDA.n2118 GNDA.t319 65.8183
R2864 GNDA.n2040 GNDA.t319 65.8183
R2865 GNDA.n2051 GNDA.t319 65.8183
R2866 GNDA.n2038 GNDA.t319 65.8183
R2867 GNDA.t264 GNDA.n2167 65.8183
R2868 GNDA.t264 GNDA.n2165 65.8183
R2869 GNDA.t264 GNDA.n2163 65.8183
R2870 GNDA.t264 GNDA.n2170 65.8183
R2871 GNDA.t264 GNDA.n2171 65.8183
R2872 GNDA.t264 GNDA.n2172 65.8183
R2873 GNDA.t264 GNDA.n2173 65.8183
R2874 GNDA.t264 GNDA.n2166 65.8183
R2875 GNDA.t264 GNDA.n2164 65.8183
R2876 GNDA.t264 GNDA.n2162 65.8183
R2877 GNDA.t264 GNDA.n2161 65.8183
R2878 GNDA.n1641 GNDA.t228 65.8183
R2879 GNDA.n1638 GNDA.t228 65.8183
R2880 GNDA.n1632 GNDA.t228 65.8183
R2881 GNDA.n1647 GNDA.t228 65.8183
R2882 GNDA.n1591 GNDA.t228 65.8183
R2883 GNDA.n1654 GNDA.t228 65.8183
R2884 GNDA.n1588 GNDA.t228 65.8183
R2885 GNDA.n1584 GNDA.t228 65.8183
R2886 GNDA.n1667 GNDA.t228 65.8183
R2887 GNDA.n1673 GNDA.t228 65.8183
R2888 GNDA.n1581 GNDA.t228 65.8183
R2889 GNDA.n1680 GNDA.t228 65.8183
R2890 GNDA.n1603 GNDA.t228 65.8183
R2891 GNDA.n1614 GNDA.t228 65.8183
R2892 GNDA.n1601 GNDA.t228 65.8183
R2893 GNDA.n2262 GNDA.t264 65.8183
R2894 GNDA.t264 GNDA.n2175 65.8183
R2895 GNDA.t264 GNDA.n2176 65.8183
R2896 GNDA.t264 GNDA.n2177 65.8183
R2897 GNDA.t288 GNDA.n982 65.8183
R2898 GNDA.t288 GNDA.n980 65.8183
R2899 GNDA.t288 GNDA.n978 65.8183
R2900 GNDA.t288 GNDA.n985 65.8183
R2901 GNDA.t288 GNDA.n986 65.8183
R2902 GNDA.t288 GNDA.n987 65.8183
R2903 GNDA.t288 GNDA.n988 65.8183
R2904 GNDA.t288 GNDA.n981 65.8183
R2905 GNDA.t288 GNDA.n979 65.8183
R2906 GNDA.t288 GNDA.n977 65.8183
R2907 GNDA.t288 GNDA.n976 65.8183
R2908 GNDA.n1148 GNDA.t288 65.8183
R2909 GNDA.t288 GNDA.n990 65.8183
R2910 GNDA.t288 GNDA.n991 65.8183
R2911 GNDA.t288 GNDA.n992 65.8183
R2912 GNDA.n1387 GNDA.t233 65.8183
R2913 GNDA.n1308 GNDA.t233 65.8183
R2914 GNDA.n1321 GNDA.t233 65.8183
R2915 GNDA.n1323 GNDA.t233 65.8183
R2916 GNDA.n1200 GNDA.t237 65.8183
R2917 GNDA.t237 GNDA.n882 65.8183
R2918 GNDA.t237 GNDA.n883 65.8183
R2919 GNDA.t237 GNDA.n884 65.8183
R2920 GNDA.n335 GNDA.t281 65.8183
R2921 GNDA.n254 GNDA.t281 65.8183
R2922 GNDA.n269 GNDA.t281 65.8183
R2923 GNDA.n271 GNDA.t281 65.8183
R2924 GNDA.n766 GNDA.n546 64.0005
R2925 GNDA.n766 GNDA.n540 64.0005
R2926 GNDA.t183 GNDA.t120 62.6786
R2927 GNDA.t22 GNDA.t279 62.6786
R2928 GNDA.t91 GNDA.t296 62.6786
R2929 GNDA.t10 GNDA.t192 62.6786
R2930 GNDA.t238 GNDA.n0 32.9056
R2931 GNDA.n736 GNDA.n735 60.8005
R2932 GNDA.t52 GNDA.t272 59.9664
R2933 GNDA.n1566 GNDA.n476 59.6972
R2934 GNDA.n1760 GNDA.n1718 59.6972
R2935 GNDA.t149 GNDA.n482 59.3736
R2936 GNDA.n316 GNDA.t281 57.8461
R2937 GNDA.t237 GNDA.n875 57.8461
R2938 GNDA.n1368 GNDA.t233 57.8461
R2939 GNDA.n2099 GNDA.t319 57.8461
R2940 GNDA.n162 GNDA.t245 57.8461
R2941 GNDA.t320 GNDA.n1781 57.8461
R2942 GNDA.t264 GNDA.n2168 57.8461
R2943 GNDA.n1661 GNDA.t228 57.8461
R2944 GNDA.t288 GNDA.n983 57.8461
R2945 GNDA.t142 GNDA.n613 56.4986
R2946 GNDA.n1495 GNDA.t221 56.4108
R2947 GNDA.t283 GNDA.t28 56.4108
R2948 GNDA.t28 GNDA.t34 56.4108
R2949 GNDA.t34 GNDA.n1501 56.4108
R2950 GNDA.n1501 GNDA.t199 56.4108
R2951 GNDA.n1511 GNDA.t353 56.4108
R2952 GNDA.n1511 GNDA.t123 56.4108
R2953 GNDA.t123 GNDA.t191 56.4108
R2954 GNDA.t191 GNDA.t276 56.4108
R2955 GNDA.n1513 GNDA.t163 56.4108
R2956 GNDA.t109 GNDA.t4 56.0277
R2957 GNDA.t134 GNDA.t38 56.0277
R2958 GNDA.t146 GNDA.t8 56.0277
R2959 GNDA.t116 GNDA.t19 56.0277
R2960 GNDA.n130 GNDA.t245 55.2026
R2961 GNDA.t320 GNDA.n1894 55.2026
R2962 GNDA.n2067 GNDA.t319 55.2026
R2963 GNDA.n1629 GNDA.t228 55.2026
R2964 GNDA.t264 GNDA.n2261 55.2026
R2965 GNDA.t288 GNDA.n1147 55.2026
R2966 GNDA.n1336 GNDA.t233 55.2026
R2967 GNDA.t237 GNDA.n1199 55.2026
R2968 GNDA.n284 GNDA.t281 55.2026
R2969 GNDA.n735 GNDA.n734 54.4005
R2970 GNDA.n335 GNDA.n334 53.3664
R2971 GNDA.n254 GNDA.n231 53.3664
R2972 GNDA.n269 GNDA.n268 53.3664
R2973 GNDA.n272 GNDA.n271 53.3664
R2974 GNDA.n333 GNDA.n332 53.3664
R2975 GNDA.n326 GNDA.n232 53.3664
R2976 GNDA.n325 GNDA.n324 53.3664
R2977 GNDA.n318 GNDA.n234 53.3664
R2978 GNDA.n311 GNDA.n238 53.3664
R2979 GNDA.n309 GNDA.n308 53.3664
R2980 GNDA.n304 GNDA.n241 53.3664
R2981 GNDA.n302 GNDA.n301 53.3664
R2982 GNDA.n288 GNDA.n287 53.3664
R2983 GNDA.n293 GNDA.n292 53.3664
R2984 GNDA.n296 GNDA.n295 53.3664
R2985 GNDA.n297 GNDA.n296 53.3664
R2986 GNDA.n294 GNDA.n293 53.3664
R2987 GNDA.n287 GNDA.n245 53.3664
R2988 GNDA.n303 GNDA.n302 53.3664
R2989 GNDA.n241 GNDA.n239 53.3664
R2990 GNDA.n310 GNDA.n309 53.3664
R2991 GNDA.n238 GNDA.n236 53.3664
R2992 GNDA.n319 GNDA.n318 53.3664
R2993 GNDA.n324 GNDA.n323 53.3664
R2994 GNDA.n327 GNDA.n326 53.3664
R2995 GNDA.n332 GNDA.n331 53.3664
R2996 GNDA.n1201 GNDA.n1200 53.3664
R2997 GNDA.n947 GNDA.n882 53.3664
R2998 GNDA.n949 GNDA.n883 53.3664
R2999 GNDA.n961 GNDA.n884 53.3664
R3000 GNDA.n868 GNDA.n866 53.3664
R3001 GNDA.n891 GNDA.n869 53.3664
R3002 GNDA.n895 GNDA.n871 53.3664
R3003 GNDA.n899 GNDA.n873 53.3664
R3004 GNDA.n910 GNDA.n880 53.3664
R3005 GNDA.n914 GNDA.n879 53.3664
R3006 GNDA.n918 GNDA.n878 53.3664
R3007 GNDA.n921 GNDA.n877 53.3664
R3008 GNDA.n934 GNDA.n870 53.3664
R3009 GNDA.n931 GNDA.n872 53.3664
R3010 GNDA.n927 GNDA.n874 53.3664
R3011 GNDA.n924 GNDA.n874 53.3664
R3012 GNDA.n928 GNDA.n872 53.3664
R3013 GNDA.n932 GNDA.n870 53.3664
R3014 GNDA.n919 GNDA.n877 53.3664
R3015 GNDA.n915 GNDA.n878 53.3664
R3016 GNDA.n911 GNDA.n879 53.3664
R3017 GNDA.n907 GNDA.n880 53.3664
R3018 GNDA.n902 GNDA.n873 53.3664
R3019 GNDA.n898 GNDA.n871 53.3664
R3020 GNDA.n894 GNDA.n869 53.3664
R3021 GNDA.n890 GNDA.n868 53.3664
R3022 GNDA.n1387 GNDA.n1386 53.3664
R3023 GNDA.n1308 GNDA.n1283 53.3664
R3024 GNDA.n1321 GNDA.n1320 53.3664
R3025 GNDA.n1324 GNDA.n1323 53.3664
R3026 GNDA.n1385 GNDA.n1284 53.3664
R3027 GNDA.n1381 GNDA.n1380 53.3664
R3028 GNDA.n1374 GNDA.n1286 53.3664
R3029 GNDA.n1373 GNDA.n1287 53.3664
R3030 GNDA.n1363 GNDA.n1291 53.3664
R3031 GNDA.n1361 GNDA.n1360 53.3664
R3032 GNDA.n1356 GNDA.n1294 53.3664
R3033 GNDA.n1354 GNDA.n1353 53.3664
R3034 GNDA.n1340 GNDA.n1339 53.3664
R3035 GNDA.n1345 GNDA.n1344 53.3664
R3036 GNDA.n1348 GNDA.n1347 53.3664
R3037 GNDA.n1349 GNDA.n1348 53.3664
R3038 GNDA.n1346 GNDA.n1345 53.3664
R3039 GNDA.n1339 GNDA.n1298 53.3664
R3040 GNDA.n1355 GNDA.n1354 53.3664
R3041 GNDA.n1294 GNDA.n1292 53.3664
R3042 GNDA.n1362 GNDA.n1361 53.3664
R3043 GNDA.n1291 GNDA.n1289 53.3664
R3044 GNDA.n1370 GNDA.n1287 53.3664
R3045 GNDA.n1375 GNDA.n1374 53.3664
R3046 GNDA.n1380 GNDA.n1379 53.3664
R3047 GNDA.n1382 GNDA.n1284 53.3664
R3048 GNDA.n2118 GNDA.n2117 53.3664
R3049 GNDA.n2040 GNDA.n2017 53.3664
R3050 GNDA.n2051 GNDA.n2050 53.3664
R3051 GNDA.n2039 GNDA.n2038 53.3664
R3052 GNDA.n2116 GNDA.n2018 53.3664
R3053 GNDA.n2112 GNDA.n2111 53.3664
R3054 GNDA.n2105 GNDA.n2020 53.3664
R3055 GNDA.n2104 GNDA.n2021 53.3664
R3056 GNDA.n2094 GNDA.n2025 53.3664
R3057 GNDA.n2092 GNDA.n2091 53.3664
R3058 GNDA.n2087 GNDA.n2028 53.3664
R3059 GNDA.n2085 GNDA.n2084 53.3664
R3060 GNDA.n2071 GNDA.n2070 53.3664
R3061 GNDA.n2076 GNDA.n2075 53.3664
R3062 GNDA.n2079 GNDA.n2078 53.3664
R3063 GNDA.n2080 GNDA.n2079 53.3664
R3064 GNDA.n2077 GNDA.n2076 53.3664
R3065 GNDA.n2070 GNDA.n2032 53.3664
R3066 GNDA.n2086 GNDA.n2085 53.3664
R3067 GNDA.n2028 GNDA.n2026 53.3664
R3068 GNDA.n2093 GNDA.n2092 53.3664
R3069 GNDA.n2025 GNDA.n2023 53.3664
R3070 GNDA.n2101 GNDA.n2021 53.3664
R3071 GNDA.n2106 GNDA.n2105 53.3664
R3072 GNDA.n2111 GNDA.n2110 53.3664
R3073 GNDA.n2113 GNDA.n2018 53.3664
R3074 GNDA.n181 GNDA.n180 53.3664
R3075 GNDA.n100 GNDA.n77 53.3664
R3076 GNDA.n115 GNDA.n114 53.3664
R3077 GNDA.n118 GNDA.n117 53.3664
R3078 GNDA.n179 GNDA.n178 53.3664
R3079 GNDA.n172 GNDA.n78 53.3664
R3080 GNDA.n171 GNDA.n170 53.3664
R3081 GNDA.n164 GNDA.n80 53.3664
R3082 GNDA.n157 GNDA.n84 53.3664
R3083 GNDA.n155 GNDA.n154 53.3664
R3084 GNDA.n150 GNDA.n87 53.3664
R3085 GNDA.n148 GNDA.n147 53.3664
R3086 GNDA.n134 GNDA.n133 53.3664
R3087 GNDA.n139 GNDA.n138 53.3664
R3088 GNDA.n142 GNDA.n141 53.3664
R3089 GNDA.n143 GNDA.n142 53.3664
R3090 GNDA.n140 GNDA.n139 53.3664
R3091 GNDA.n133 GNDA.n91 53.3664
R3092 GNDA.n149 GNDA.n148 53.3664
R3093 GNDA.n87 GNDA.n85 53.3664
R3094 GNDA.n156 GNDA.n155 53.3664
R3095 GNDA.n84 GNDA.n82 53.3664
R3096 GNDA.n165 GNDA.n164 53.3664
R3097 GNDA.n170 GNDA.n169 53.3664
R3098 GNDA.n173 GNDA.n172 53.3664
R3099 GNDA.n178 GNDA.n177 53.3664
R3100 GNDA.n182 GNDA.n181 53.3664
R3101 GNDA.n101 GNDA.n100 53.3664
R3102 GNDA.n116 GNDA.n115 53.3664
R3103 GNDA.n117 GNDA.n94 53.3664
R3104 GNDA.n1896 GNDA.n1895 53.3664
R3105 GNDA.n1852 GNDA.n1788 53.3664
R3106 GNDA.n1871 GNDA.n1789 53.3664
R3107 GNDA.n1877 GNDA.n1790 53.3664
R3108 GNDA.n1774 GNDA.n1772 53.3664
R3109 GNDA.n1794 GNDA.n1775 53.3664
R3110 GNDA.n1798 GNDA.n1777 53.3664
R3111 GNDA.n1802 GNDA.n1779 53.3664
R3112 GNDA.n1813 GNDA.n1786 53.3664
R3113 GNDA.n1817 GNDA.n1785 53.3664
R3114 GNDA.n1821 GNDA.n1784 53.3664
R3115 GNDA.n1824 GNDA.n1783 53.3664
R3116 GNDA.n1837 GNDA.n1776 53.3664
R3117 GNDA.n1834 GNDA.n1778 53.3664
R3118 GNDA.n1830 GNDA.n1780 53.3664
R3119 GNDA.n1827 GNDA.n1780 53.3664
R3120 GNDA.n1831 GNDA.n1778 53.3664
R3121 GNDA.n1835 GNDA.n1776 53.3664
R3122 GNDA.n1822 GNDA.n1783 53.3664
R3123 GNDA.n1818 GNDA.n1784 53.3664
R3124 GNDA.n1814 GNDA.n1785 53.3664
R3125 GNDA.n1810 GNDA.n1786 53.3664
R3126 GNDA.n1805 GNDA.n1779 53.3664
R3127 GNDA.n1801 GNDA.n1777 53.3664
R3128 GNDA.n1797 GNDA.n1775 53.3664
R3129 GNDA.n1793 GNDA.n1774 53.3664
R3130 GNDA.n1895 GNDA.n1773 53.3664
R3131 GNDA.n1870 GNDA.n1788 53.3664
R3132 GNDA.n1876 GNDA.n1789 53.3664
R3133 GNDA.n1842 GNDA.n1790 53.3664
R3134 GNDA.n2119 GNDA.n2118 53.3664
R3135 GNDA.n2041 GNDA.n2040 53.3664
R3136 GNDA.n2052 GNDA.n2051 53.3664
R3137 GNDA.n2038 GNDA.n2035 53.3664
R3138 GNDA.n2263 GNDA.n2262 53.3664
R3139 GNDA.n2182 GNDA.n2175 53.3664
R3140 GNDA.n2189 GNDA.n2176 53.3664
R3141 GNDA.n2196 GNDA.n2177 53.3664
R3142 GNDA.n2161 GNDA.n2159 53.3664
R3143 GNDA.n2207 GNDA.n2162 53.3664
R3144 GNDA.n2211 GNDA.n2164 53.3664
R3145 GNDA.n2215 GNDA.n2166 53.3664
R3146 GNDA.n2226 GNDA.n2173 53.3664
R3147 GNDA.n2230 GNDA.n2172 53.3664
R3148 GNDA.n2234 GNDA.n2171 53.3664
R3149 GNDA.n2237 GNDA.n2170 53.3664
R3150 GNDA.n2250 GNDA.n2163 53.3664
R3151 GNDA.n2247 GNDA.n2165 53.3664
R3152 GNDA.n2243 GNDA.n2167 53.3664
R3153 GNDA.n2240 GNDA.n2167 53.3664
R3154 GNDA.n2244 GNDA.n2165 53.3664
R3155 GNDA.n2248 GNDA.n2163 53.3664
R3156 GNDA.n2235 GNDA.n2170 53.3664
R3157 GNDA.n2231 GNDA.n2171 53.3664
R3158 GNDA.n2227 GNDA.n2172 53.3664
R3159 GNDA.n2223 GNDA.n2173 53.3664
R3160 GNDA.n2218 GNDA.n2166 53.3664
R3161 GNDA.n2214 GNDA.n2164 53.3664
R3162 GNDA.n2210 GNDA.n2162 53.3664
R3163 GNDA.n2206 GNDA.n2161 53.3664
R3164 GNDA.n1680 GNDA.n1679 53.3664
R3165 GNDA.n1603 GNDA.n1580 53.3664
R3166 GNDA.n1614 GNDA.n1613 53.3664
R3167 GNDA.n1602 GNDA.n1601 53.3664
R3168 GNDA.n1678 GNDA.n1581 53.3664
R3169 GNDA.n1674 GNDA.n1673 53.3664
R3170 GNDA.n1667 GNDA.n1583 53.3664
R3171 GNDA.n1666 GNDA.n1584 53.3664
R3172 GNDA.n1656 GNDA.n1588 53.3664
R3173 GNDA.n1654 GNDA.n1653 53.3664
R3174 GNDA.n1649 GNDA.n1591 53.3664
R3175 GNDA.n1647 GNDA.n1646 53.3664
R3176 GNDA.n1633 GNDA.n1632 53.3664
R3177 GNDA.n1638 GNDA.n1637 53.3664
R3178 GNDA.n1641 GNDA.n1640 53.3664
R3179 GNDA.n1642 GNDA.n1641 53.3664
R3180 GNDA.n1639 GNDA.n1638 53.3664
R3181 GNDA.n1632 GNDA.n1595 53.3664
R3182 GNDA.n1648 GNDA.n1647 53.3664
R3183 GNDA.n1591 GNDA.n1589 53.3664
R3184 GNDA.n1655 GNDA.n1654 53.3664
R3185 GNDA.n1588 GNDA.n1586 53.3664
R3186 GNDA.n1663 GNDA.n1584 53.3664
R3187 GNDA.n1668 GNDA.n1667 53.3664
R3188 GNDA.n1673 GNDA.n1672 53.3664
R3189 GNDA.n1675 GNDA.n1581 53.3664
R3190 GNDA.n1681 GNDA.n1680 53.3664
R3191 GNDA.n1604 GNDA.n1603 53.3664
R3192 GNDA.n1615 GNDA.n1614 53.3664
R3193 GNDA.n1601 GNDA.n1598 53.3664
R3194 GNDA.n2262 GNDA.n2160 53.3664
R3195 GNDA.n2190 GNDA.n2175 53.3664
R3196 GNDA.n2197 GNDA.n2176 53.3664
R3197 GNDA.n2179 GNDA.n2177 53.3664
R3198 GNDA.n1149 GNDA.n1148 53.3664
R3199 GNDA.n1055 GNDA.n990 53.3664
R3200 GNDA.n1057 GNDA.n991 53.3664
R3201 GNDA.n1069 GNDA.n992 53.3664
R3202 GNDA.n976 GNDA.n974 53.3664
R3203 GNDA.n999 GNDA.n977 53.3664
R3204 GNDA.n1003 GNDA.n979 53.3664
R3205 GNDA.n1007 GNDA.n981 53.3664
R3206 GNDA.n1018 GNDA.n988 53.3664
R3207 GNDA.n1022 GNDA.n987 53.3664
R3208 GNDA.n1026 GNDA.n986 53.3664
R3209 GNDA.n1029 GNDA.n985 53.3664
R3210 GNDA.n1042 GNDA.n978 53.3664
R3211 GNDA.n1039 GNDA.n980 53.3664
R3212 GNDA.n1035 GNDA.n982 53.3664
R3213 GNDA.n1032 GNDA.n982 53.3664
R3214 GNDA.n1036 GNDA.n980 53.3664
R3215 GNDA.n1040 GNDA.n978 53.3664
R3216 GNDA.n1027 GNDA.n985 53.3664
R3217 GNDA.n1023 GNDA.n986 53.3664
R3218 GNDA.n1019 GNDA.n987 53.3664
R3219 GNDA.n1015 GNDA.n988 53.3664
R3220 GNDA.n1010 GNDA.n981 53.3664
R3221 GNDA.n1006 GNDA.n979 53.3664
R3222 GNDA.n1002 GNDA.n977 53.3664
R3223 GNDA.n998 GNDA.n976 53.3664
R3224 GNDA.n1148 GNDA.n975 53.3664
R3225 GNDA.n1058 GNDA.n990 53.3664
R3226 GNDA.n1068 GNDA.n991 53.3664
R3227 GNDA.n994 GNDA.n992 53.3664
R3228 GNDA.n1388 GNDA.n1387 53.3664
R3229 GNDA.n1309 GNDA.n1308 53.3664
R3230 GNDA.n1322 GNDA.n1321 53.3664
R3231 GNDA.n1323 GNDA.n1301 53.3664
R3232 GNDA.n1200 GNDA.n867 53.3664
R3233 GNDA.n950 GNDA.n882 53.3664
R3234 GNDA.n960 GNDA.n883 53.3664
R3235 GNDA.n886 GNDA.n884 53.3664
R3236 GNDA.n336 GNDA.n335 53.3664
R3237 GNDA.n255 GNDA.n254 53.3664
R3238 GNDA.n270 GNDA.n269 53.3664
R3239 GNDA.n271 GNDA.n248 53.3664
R3240 GNDA.t68 GNDA.t347 52.4707
R3241 GNDA.t147 GNDA.t118 52.4707
R3242 GNDA.t317 GNDA.t266 52.4707
R3243 GNDA.n546 GNDA.n545 51.2005
R3244 GNDA.n759 GNDA.n540 51.2005
R3245 GNDA.n1457 GNDA.n1456 50.9355
R3246 GNDA.n2512 GNDA.n5 50.5752
R3247 GNDA.n1496 GNDA.t166 50.1429
R3248 GNDA.t221 GNDA.t183 50.1429
R3249 GNDA.t74 GNDA.t22 50.1429
R3250 GNDA.t215 GNDA.t91 50.1429
R3251 GNDA.t163 GNDA.t10 50.1429
R3252 GNDA.n1515 GNDA.t219 50.1429
R3253 GNDA.n625 GNDA.t14 48.5574
R3254 GNDA.n608 GNDA.t54 48.5574
R3255 GNDA.n656 GNDA.t135 48.5574
R3256 GNDA.t179 GNDA.n714 48.5574
R3257 GNDA.n856 GNDA.t238 48.2626
R3258 GNDA.n750 GNDA.t343 48.0005
R3259 GNDA.n750 GNDA.t172 48.0005
R3260 GNDA.n747 GNDA.t113 48.0005
R3261 GNDA.n747 GNDA.t94 48.0005
R3262 GNDA.n746 GNDA.t348 48.0005
R3263 GNDA.n746 GNDA.t119 48.0005
R3264 GNDA.n744 GNDA.t198 48.0005
R3265 GNDA.n744 GNDA.t189 48.0005
R3266 GNDA.n743 GNDA.t213 48.0005
R3267 GNDA.n743 GNDA.t6 48.0005
R3268 GNDA.n1126 GNDA.t238 47.9486
R3269 GNDA.n2427 GNDA.t238 47.9486
R3270 GNDA.n2457 GNDA.t238 47.9486
R3271 GNDA.n194 GNDA.t238 47.6748
R3272 GNDA.n1560 GNDA.n482 45.6721
R3273 GNDA.n1914 GNDA.n1699 45.6509
R3274 GNDA.t111 GNDA.t65 44.9749
R3275 GNDA.t214 GNDA.t83 44.9749
R3276 GNDA.t329 GNDA.t79 44.9749
R3277 GNDA.t143 GNDA.t25 44.9749
R3278 GNDA.t211 GNDA.t358 44.9749
R3279 GNDA.t201 GNDA.t151 44.9749
R3280 GNDA.t50 GNDA.t206 44.9749
R3281 GNDA.t327 GNDA.t61 44.9749
R3282 GNDA.n641 GNDA.n640 44.8222
R3283 GNDA.n585 GNDA.n510 44.8222
R3284 GNDA.n621 GNDA.n620 44.8005
R3285 GNDA.n500 GNDA.n491 44.8005
R3286 GNDA.n1503 GNDA.t29 43.8751
R3287 GNDA.n1523 GNDA.t159 43.8751
R3288 GNDA.n1128 GNDA.t238 43.8679
R3289 GNDA.t238 GNDA.n55 43.8679
R3290 GNDA.n2450 GNDA.t238 43.8679
R3291 GNDA.n1314 GNDA.n1278 43.0993
R3292 GNDA.n730 GNDA.t194 41.2271
R3293 GNDA.n764 GNDA.t349 41.2271
R3294 GNDA.n588 GNDA.t204 41.2271
R3295 GNDA.t180 GNDA.n770 41.2271
R3296 GNDA.n770 GNDA.t325 41.2271
R3297 GNDA.t108 GNDA.n473 41.1049
R3298 GNDA.t161 GNDA.n625 41.0871
R3299 GNDA.t96 GNDA.n608 41.0871
R3300 GNDA.t46 GNDA.t131 41.0871
R3301 GNDA.t46 GNDA.t128 41.0871
R3302 GNDA.t89 GNDA.t210 41.0871
R3303 GNDA.t89 GNDA.t184 41.0871
R3304 GNDA.n575 GNDA.t71 40.7412
R3305 GNDA.t351 GNDA.n578 40.7412
R3306 GNDA.t165 GNDA.n1494 37.6073
R3307 GNDA.n1494 GNDA.t29 37.6073
R3308 GNDA.n1502 GNDA.t107 37.6073
R3309 GNDA.n1545 GNDA.n814 37.6073
R3310 GNDA.n1545 GNDA.n817 37.6073
R3311 GNDA.n1524 GNDA.t45 37.6073
R3312 GNDA.t159 GNDA.n1522 37.6073
R3313 GNDA.n1522 GNDA.t99 37.6073
R3314 GNDA.t311 GNDA.t250 37.4792
R3315 GNDA.t337 GNDA.t240 37.4792
R3316 GNDA.t339 GNDA.t256 37.4792
R3317 GNDA.t5 GNDA.t190 37.4792
R3318 GNDA.t340 GNDA.t188 37.4792
R3319 GNDA.t85 GNDA.t342 37.4792
R3320 GNDA.t103 GNDA.t171 37.4792
R3321 GNDA.t53 GNDA.t112 37.4792
R3322 GNDA.t235 GNDA.t93 37.4792
R3323 GNDA.t18 GNDA.t63 37.4792
R3324 GNDA.t204 GNDA.t111 37.4792
R3325 GNDA.n788 GNDA.n787 36.9067
R3326 GNDA.n673 GNDA.n672 36.6567
R3327 GNDA.t51 GNDA.n575 34.4734
R3328 GNDA.n578 GNDA.t160 34.4734
R3329 GNDA.t194 GNDA.n728 33.7313
R3330 GNDA.n740 GNDA.t195 33.7313
R3331 GNDA.n739 GNDA.t212 33.7313
R3332 GNDA.n704 GNDA.t197 33.7313
R3333 GNDA.t153 GNDA.n756 33.7313
R3334 GNDA.t322 GNDA.n771 33.7313
R3335 GNDA.n656 GNDA.t128 33.6168
R3336 GNDA.n714 GNDA.t210 33.6168
R3337 GNDA.n375 GNDA.t238 31.6472
R3338 GNDA.n1718 GNDA.t127 31.6047
R3339 GNDA.n1503 GNDA.t30 31.3395
R3340 GNDA.t92 GNDA.n1523 31.3395
R3341 GNDA.t240 GNDA.t293 29.9835
R3342 GNDA.t256 GNDA.t33 29.9835
R3343 GNDA.t17 GNDA.t212 29.9835
R3344 GNDA.t203 GNDA.t5 29.9835
R3345 GNDA.t197 GNDA.t7 29.9835
R3346 GNDA.t286 GNDA.t299 29.9835
R3347 GNDA.n602 GNDA.n562 29.8817
R3348 GNDA.n717 GNDA.n715 29.8817
R3349 GNDA.n630 GNDA.n599 28.413
R3350 GNDA.n807 GNDA.n806 28.413
R3351 GNDA.n1933 GNDA.n472 28.1318
R3352 GNDA.n606 GNDA.n593 28.038
R3353 GNDA.n797 GNDA.n515 28.038
R3354 GNDA.n1527 GNDA.n1526 27.8193
R3355 GNDA.n1506 GNDA.n1505 27.8193
R3356 GNDA.n300 GNDA.n299 27.5561
R3357 GNDA.n923 GNDA.n922 27.5561
R3358 GNDA.n1352 GNDA.n1351 27.5561
R3359 GNDA.n2083 GNDA.n2082 27.5561
R3360 GNDA.n146 GNDA.n145 27.5561
R3361 GNDA.n1826 GNDA.n1825 27.5561
R3362 GNDA.n2239 GNDA.n2238 27.5561
R3363 GNDA.n1645 GNDA.n1644 27.5561
R3364 GNDA.n1031 GNDA.n1030 27.5561
R3365 GNDA.n1931 GNDA.n1930 27.4034
R3366 GNDA.n0 GNDA.n46 8.60107
R3367 GNDA.n764 GNDA.t55 26.2356
R3368 GNDA.n587 GNDA.t157 26.2356
R3369 GNDA.n712 GNDA.t325 26.2356
R3370 GNDA.t139 GNDA.t109 26.1465
R3371 GNDA.t38 GNDA.t135 26.1465
R3372 GNDA.t8 GNDA.t179 26.1465
R3373 GNDA.t0 GNDA.t116 26.1465
R3374 GNDA.n517 GNDA.n508 25.6005
R3375 GNDA.n654 GNDA.n651 25.6005
R3376 GNDA.n1484 GNDA.t169 25.0717
R3377 GNDA.t31 GNDA.t74 25.0717
R3378 GNDA.t30 GNDA.t175 25.0717
R3379 GNDA.t355 GNDA.t92 25.0717
R3380 GNDA.t352 GNDA.t215 25.0717
R3381 GNDA.n1534 GNDA.t72 25.0717
R3382 GNDA.t127 GNDA.t11 24.5815
R3383 GNDA.n1079 GNDA.t238 24.4846
R3384 GNDA.n844 GNDA.t170 24.0005
R3385 GNDA.n844 GNDA.t174 24.0005
R3386 GNDA.n842 GNDA.t167 24.0005
R3387 GNDA.n842 GNDA.t222 24.0005
R3388 GNDA.n840 GNDA.t121 24.0005
R3389 GNDA.n840 GNDA.t75 24.0005
R3390 GNDA.n838 GNDA.t35 24.0005
R3391 GNDA.n838 GNDA.t200 24.0005
R3392 GNDA.n836 GNDA.t224 24.0005
R3393 GNDA.n836 GNDA.t115 24.0005
R3394 GNDA.n834 GNDA.t37 24.0005
R3395 GNDA.n834 GNDA.t102 24.0005
R3396 GNDA.n832 GNDA.t354 24.0005
R3397 GNDA.n832 GNDA.t124 24.0005
R3398 GNDA.n830 GNDA.t216 24.0005
R3399 GNDA.n830 GNDA.t193 24.0005
R3400 GNDA.n828 GNDA.t164 24.0005
R3401 GNDA.n828 GNDA.t220 24.0005
R3402 GNDA.n827 GNDA.t218 24.0005
R3403 GNDA.n827 GNDA.t73 24.0005
R3404 GNDA.n676 GNDA.t251 24.0005
R3405 GNDA.n676 GNDA.t196 24.0005
R3406 GNDA.n314 GNDA.n235 23.6449
R3407 GNDA.n905 GNDA.n904 23.6449
R3408 GNDA.n1366 GNDA.n1288 23.6449
R3409 GNDA.n2097 GNDA.n2022 23.6449
R3410 GNDA.n160 GNDA.n81 23.6449
R3411 GNDA.n1808 GNDA.n1807 23.6449
R3412 GNDA.n2221 GNDA.n2220 23.6449
R3413 GNDA.n1659 GNDA.n1585 23.6449
R3414 GNDA.n1013 GNDA.n1012 23.6449
R3415 GNDA.n1458 GNDA.n1457 23.509
R3416 GNDA.n790 GNDA.n521 23.488
R3417 GNDA.t65 GNDA.t305 22.4877
R3418 GNDA.t83 GNDA.t346 22.4877
R3419 GNDA.t157 GNDA.t336 22.4877
R3420 GNDA.t79 GNDA.t360 22.4877
R3421 GNDA.t25 GNDA.t344 22.4877
R3422 GNDA.t358 GNDA.t16 22.4877
R3423 GNDA.t151 GNDA.t335 22.4877
R3424 GNDA.t206 GNDA.t338 22.4877
R3425 GNDA.t61 GNDA.t328 22.4877
R3426 GNDA.t57 GNDA.t52 22.4877
R3427 GNDA.t272 GNDA.t180 22.4877
R3428 GNDA.n638 GNDA.n606 22.4005
R3429 GNDA.n536 GNDA.n535 22.4005
R3430 GNDA.n535 GNDA.n534 22.4005
R3431 GNDA.n707 GNDA.n702 22.4005
R3432 GNDA.n709 GNDA.n591 22.4005
R3433 GNDA.n734 GNDA.n561 22.4005
R3434 GNDA.n736 GNDA.n560 22.4005
R3435 GNDA.n583 GNDA.n515 22.4005
R3436 GNDA.n1934 GNDA.n2 21.4917
R3437 GNDA.n1507 GNDA.n1467 21.3338
R3438 GNDA.n1509 GNDA.n1466 21.3338
R3439 GNDA.n1530 GNDA.n1462 21.3338
R3440 GNDA.n1528 GNDA.n1463 21.3338
R3441 GNDA.n1479 GNDA.n1477 21.3338
R3442 GNDA.n1471 GNDA.n1470 21.3338
R3443 GNDA.n598 GNDA.n597 21.3338
R3444 GNDA.n530 GNDA.n529 21.3338
R3445 GNDA.n534 GNDA.n533 21.3338
R3446 GNDA.n536 GNDA.n532 21.3338
R3447 GNDA.n537 GNDA.n531 21.3338
R3448 GNDA.n544 GNDA.n543 21.3338
R3449 GNDA.n545 GNDA.n542 21.3338
R3450 GNDA.n546 GNDA.n541 21.3338
R3451 GNDA.n540 GNDA.n539 21.3338
R3452 GNDA.n759 GNDA.n758 21.3338
R3453 GNDA.n760 GNDA.n757 21.3338
R3454 GNDA.n553 GNDA.n552 21.3338
R3455 GNDA.n556 GNDA.n554 21.3338
R3456 GNDA.n514 GNDA.n513 21.3338
R3457 GNDA.n518 GNDA.n516 21.3338
R3458 GNDA.n653 GNDA.n652 21.3338
R3459 GNDA.n646 GNDA.n645 21.3338
R3460 GNDA.n644 GNDA.n643 21.3338
R3461 GNDA.n505 GNDA.n504 21.3338
R3462 GNDA.n801 GNDA.n800 21.3338
R3463 GNDA.t104 GNDA.n1566 21.0699
R3464 GNDA.n789 GNDA 20.281
R3465 GNDA.n621 GNDA.n612 20.2755
R3466 GNDA.n501 GNDA.n500 20.2755
R3467 GNDA.n826 GNDA.n825 19.7404
R3468 GNDA.n786 GNDA.t177 19.7005
R3469 GNDA.n786 GNDA.t187 19.7005
R3470 GNDA.n784 GNDA.t122 19.7005
R3471 GNDA.n784 GNDA.t125 19.7005
R3472 GNDA.n782 GNDA.t186 19.7005
R3473 GNDA.n782 GNDA.t208 19.7005
R3474 GNDA.n780 GNDA.t76 19.7005
R3475 GNDA.n780 GNDA.t32 19.7005
R3476 GNDA.n778 GNDA.t185 19.7005
R3477 GNDA.n778 GNDA.t1 19.7005
R3478 GNDA.n777 GNDA.t67 19.7005
R3479 GNDA.n777 GNDA.t126 19.7005
R3480 GNDA.n671 GNDA.t48 19.7005
R3481 GNDA.n671 GNDA.t133 19.7005
R3482 GNDA.n669 GNDA.t136 19.7005
R3483 GNDA.n669 GNDA.t137 19.7005
R3484 GNDA.n667 GNDA.t88 19.7005
R3485 GNDA.n667 GNDA.t43 19.7005
R3486 GNDA.n665 GNDA.t130 19.7005
R3487 GNDA.n665 GNDA.t87 19.7005
R3488 GNDA.n663 GNDA.t129 19.7005
R3489 GNDA.n663 GNDA.t86 19.7005
R3490 GNDA.n662 GNDA.t140 19.7005
R3491 GNDA.n662 GNDA.t49 19.7005
R3492 GNDA.n767 GNDA.n766 19.288
R3493 GNDA.n1934 GNDA.n470 19.2005
R3494 GNDA.n1564 GNDA.n480 19.2005
R3495 GNDA.n1740 GNDA.n1739 19.2005
R3496 GNDA.n1538 GNDA.n1537 19.2005
R3497 GNDA.n1492 GNDA.n1491 19.2005
R3498 GNDA.n1556 GNDA.n471 19.2005
R3499 GNDA.n805 GNDA.n508 19.1005
R3500 GNDA.n651 GNDA.n650 19.1005
R3501 GNDA.t100 GNDA.t283 18.8039
R3502 GNDA.t114 GNDA.n814 18.8039
R3503 GNDA.t36 GNDA.n817 18.8039
R3504 GNDA.t276 GNDA.t41 18.8039
R3505 GNDA.t345 GNDA.n587 18.7399
R3506 GNDA.n848 GNDA.n826 18.4413
R3507 GNDA.n1480 GNDA.n1 18.3355
R3508 GNDA.t95 GNDA.t108 18.2691
R3509 GNDA.n1931 GNDA.n473 18.2691
R3510 GNDA.t11 GNDA.t138 18.2691
R3511 GNDA.n1539 GNDA.n1538 17.613
R3512 GNDA.n2515 GNDA.n2514 17.4917
R3513 GNDA.n2469 GNDA.n29 17.0672
R3514 GNDA.n1088 GNDA.n1087 17.0672
R3515 GNDA.n2416 GNDA.n61 17.0672
R3516 GNDA.n2510 GNDA.n2509 16.9605
R3517 GNDA.n247 GNDA.n246 16.0005
R3518 GNDA.n289 GNDA.n246 16.0005
R3519 GNDA.n290 GNDA.n289 16.0005
R3520 GNDA.n291 GNDA.n290 16.0005
R3521 GNDA.n291 GNDA.n244 16.0005
R3522 GNDA.n244 GNDA.n243 16.0005
R3523 GNDA.n298 GNDA.n243 16.0005
R3524 GNDA.n299 GNDA.n298 16.0005
R3525 GNDA.n314 GNDA.n313 16.0005
R3526 GNDA.n313 GNDA.n312 16.0005
R3527 GNDA.n312 GNDA.n237 16.0005
R3528 GNDA.n307 GNDA.n237 16.0005
R3529 GNDA.n307 GNDA.n306 16.0005
R3530 GNDA.n306 GNDA.n305 16.0005
R3531 GNDA.n305 GNDA.n240 16.0005
R3532 GNDA.n300 GNDA.n240 16.0005
R3533 GNDA.n330 GNDA.n227 16.0005
R3534 GNDA.n330 GNDA.n329 16.0005
R3535 GNDA.n329 GNDA.n328 16.0005
R3536 GNDA.n328 GNDA.n233 16.0005
R3537 GNDA.n322 GNDA.n233 16.0005
R3538 GNDA.n321 GNDA.n320 16.0005
R3539 GNDA.n320 GNDA.n235 16.0005
R3540 GNDA.n937 GNDA.n936 16.0005
R3541 GNDA.n936 GNDA.n935 16.0005
R3542 GNDA.n935 GNDA.n933 16.0005
R3543 GNDA.n933 GNDA.n930 16.0005
R3544 GNDA.n930 GNDA.n929 16.0005
R3545 GNDA.n929 GNDA.n926 16.0005
R3546 GNDA.n926 GNDA.n925 16.0005
R3547 GNDA.n925 GNDA.n923 16.0005
R3548 GNDA.n908 GNDA.n905 16.0005
R3549 GNDA.n909 GNDA.n908 16.0005
R3550 GNDA.n912 GNDA.n909 16.0005
R3551 GNDA.n913 GNDA.n912 16.0005
R3552 GNDA.n916 GNDA.n913 16.0005
R3553 GNDA.n917 GNDA.n916 16.0005
R3554 GNDA.n920 GNDA.n917 16.0005
R3555 GNDA.n922 GNDA.n920 16.0005
R3556 GNDA.n889 GNDA.n888 16.0005
R3557 GNDA.n892 GNDA.n889 16.0005
R3558 GNDA.n893 GNDA.n892 16.0005
R3559 GNDA.n896 GNDA.n893 16.0005
R3560 GNDA.n897 GNDA.n896 16.0005
R3561 GNDA.n901 GNDA.n900 16.0005
R3562 GNDA.n904 GNDA.n901 16.0005
R3563 GNDA.n1300 GNDA.n1299 16.0005
R3564 GNDA.n1341 GNDA.n1299 16.0005
R3565 GNDA.n1342 GNDA.n1341 16.0005
R3566 GNDA.n1343 GNDA.n1342 16.0005
R3567 GNDA.n1343 GNDA.n1297 16.0005
R3568 GNDA.n1297 GNDA.n1296 16.0005
R3569 GNDA.n1350 GNDA.n1296 16.0005
R3570 GNDA.n1351 GNDA.n1350 16.0005
R3571 GNDA.n1366 GNDA.n1365 16.0005
R3572 GNDA.n1365 GNDA.n1364 16.0005
R3573 GNDA.n1364 GNDA.n1290 16.0005
R3574 GNDA.n1359 GNDA.n1290 16.0005
R3575 GNDA.n1359 GNDA.n1358 16.0005
R3576 GNDA.n1358 GNDA.n1357 16.0005
R3577 GNDA.n1357 GNDA.n1293 16.0005
R3578 GNDA.n1352 GNDA.n1293 16.0005
R3579 GNDA.n1384 GNDA.n1383 16.0005
R3580 GNDA.n1383 GNDA.n1285 16.0005
R3581 GNDA.n1378 GNDA.n1285 16.0005
R3582 GNDA.n1378 GNDA.n1377 16.0005
R3583 GNDA.n1377 GNDA.n1376 16.0005
R3584 GNDA.n1372 GNDA.n1371 16.0005
R3585 GNDA.n1371 GNDA.n1288 16.0005
R3586 GNDA.n2034 GNDA.n2033 16.0005
R3587 GNDA.n2072 GNDA.n2033 16.0005
R3588 GNDA.n2073 GNDA.n2072 16.0005
R3589 GNDA.n2074 GNDA.n2073 16.0005
R3590 GNDA.n2074 GNDA.n2031 16.0005
R3591 GNDA.n2031 GNDA.n2030 16.0005
R3592 GNDA.n2081 GNDA.n2030 16.0005
R3593 GNDA.n2082 GNDA.n2081 16.0005
R3594 GNDA.n2097 GNDA.n2096 16.0005
R3595 GNDA.n2096 GNDA.n2095 16.0005
R3596 GNDA.n2095 GNDA.n2024 16.0005
R3597 GNDA.n2090 GNDA.n2024 16.0005
R3598 GNDA.n2090 GNDA.n2089 16.0005
R3599 GNDA.n2089 GNDA.n2088 16.0005
R3600 GNDA.n2088 GNDA.n2027 16.0005
R3601 GNDA.n2083 GNDA.n2027 16.0005
R3602 GNDA.n2115 GNDA.n2114 16.0005
R3603 GNDA.n2114 GNDA.n2019 16.0005
R3604 GNDA.n2109 GNDA.n2019 16.0005
R3605 GNDA.n2109 GNDA.n2108 16.0005
R3606 GNDA.n2108 GNDA.n2107 16.0005
R3607 GNDA.n2103 GNDA.n2102 16.0005
R3608 GNDA.n2102 GNDA.n2022 16.0005
R3609 GNDA.n93 GNDA.n92 16.0005
R3610 GNDA.n135 GNDA.n92 16.0005
R3611 GNDA.n136 GNDA.n135 16.0005
R3612 GNDA.n137 GNDA.n136 16.0005
R3613 GNDA.n137 GNDA.n90 16.0005
R3614 GNDA.n90 GNDA.n89 16.0005
R3615 GNDA.n144 GNDA.n89 16.0005
R3616 GNDA.n145 GNDA.n144 16.0005
R3617 GNDA.n160 GNDA.n159 16.0005
R3618 GNDA.n159 GNDA.n158 16.0005
R3619 GNDA.n158 GNDA.n83 16.0005
R3620 GNDA.n153 GNDA.n83 16.0005
R3621 GNDA.n153 GNDA.n152 16.0005
R3622 GNDA.n152 GNDA.n151 16.0005
R3623 GNDA.n151 GNDA.n86 16.0005
R3624 GNDA.n146 GNDA.n86 16.0005
R3625 GNDA.n176 GNDA.n73 16.0005
R3626 GNDA.n176 GNDA.n175 16.0005
R3627 GNDA.n175 GNDA.n174 16.0005
R3628 GNDA.n174 GNDA.n79 16.0005
R3629 GNDA.n168 GNDA.n79 16.0005
R3630 GNDA.n167 GNDA.n166 16.0005
R3631 GNDA.n166 GNDA.n81 16.0005
R3632 GNDA.n2510 GNDA.n3 16.0005
R3633 GNDA.n2514 GNDA.n3 16.0005
R3634 GNDA.n1840 GNDA.n1839 16.0005
R3635 GNDA.n1839 GNDA.n1838 16.0005
R3636 GNDA.n1838 GNDA.n1836 16.0005
R3637 GNDA.n1836 GNDA.n1833 16.0005
R3638 GNDA.n1833 GNDA.n1832 16.0005
R3639 GNDA.n1832 GNDA.n1829 16.0005
R3640 GNDA.n1829 GNDA.n1828 16.0005
R3641 GNDA.n1828 GNDA.n1826 16.0005
R3642 GNDA.n1811 GNDA.n1808 16.0005
R3643 GNDA.n1812 GNDA.n1811 16.0005
R3644 GNDA.n1815 GNDA.n1812 16.0005
R3645 GNDA.n1816 GNDA.n1815 16.0005
R3646 GNDA.n1819 GNDA.n1816 16.0005
R3647 GNDA.n1820 GNDA.n1819 16.0005
R3648 GNDA.n1823 GNDA.n1820 16.0005
R3649 GNDA.n1825 GNDA.n1823 16.0005
R3650 GNDA.n1792 GNDA.n1791 16.0005
R3651 GNDA.n1795 GNDA.n1792 16.0005
R3652 GNDA.n1796 GNDA.n1795 16.0005
R3653 GNDA.n1799 GNDA.n1796 16.0005
R3654 GNDA.n1800 GNDA.n1799 16.0005
R3655 GNDA.n1804 GNDA.n1803 16.0005
R3656 GNDA.n1807 GNDA.n1804 16.0005
R3657 GNDA.n2253 GNDA.n2252 16.0005
R3658 GNDA.n2252 GNDA.n2251 16.0005
R3659 GNDA.n2251 GNDA.n2249 16.0005
R3660 GNDA.n2249 GNDA.n2246 16.0005
R3661 GNDA.n2246 GNDA.n2245 16.0005
R3662 GNDA.n2245 GNDA.n2242 16.0005
R3663 GNDA.n2242 GNDA.n2241 16.0005
R3664 GNDA.n2241 GNDA.n2239 16.0005
R3665 GNDA.n2224 GNDA.n2221 16.0005
R3666 GNDA.n2225 GNDA.n2224 16.0005
R3667 GNDA.n2228 GNDA.n2225 16.0005
R3668 GNDA.n2229 GNDA.n2228 16.0005
R3669 GNDA.n2232 GNDA.n2229 16.0005
R3670 GNDA.n2233 GNDA.n2232 16.0005
R3671 GNDA.n2236 GNDA.n2233 16.0005
R3672 GNDA.n2238 GNDA.n2236 16.0005
R3673 GNDA.n2205 GNDA.n2156 16.0005
R3674 GNDA.n2208 GNDA.n2205 16.0005
R3675 GNDA.n2209 GNDA.n2208 16.0005
R3676 GNDA.n2212 GNDA.n2209 16.0005
R3677 GNDA.n2213 GNDA.n2212 16.0005
R3678 GNDA.n2217 GNDA.n2216 16.0005
R3679 GNDA.n2220 GNDA.n2217 16.0005
R3680 GNDA.n1597 GNDA.n1596 16.0005
R3681 GNDA.n1634 GNDA.n1596 16.0005
R3682 GNDA.n1635 GNDA.n1634 16.0005
R3683 GNDA.n1636 GNDA.n1635 16.0005
R3684 GNDA.n1636 GNDA.n1594 16.0005
R3685 GNDA.n1594 GNDA.n1593 16.0005
R3686 GNDA.n1643 GNDA.n1593 16.0005
R3687 GNDA.n1644 GNDA.n1643 16.0005
R3688 GNDA.n1659 GNDA.n1658 16.0005
R3689 GNDA.n1658 GNDA.n1657 16.0005
R3690 GNDA.n1657 GNDA.n1587 16.0005
R3691 GNDA.n1652 GNDA.n1587 16.0005
R3692 GNDA.n1652 GNDA.n1651 16.0005
R3693 GNDA.n1651 GNDA.n1650 16.0005
R3694 GNDA.n1650 GNDA.n1590 16.0005
R3695 GNDA.n1645 GNDA.n1590 16.0005
R3696 GNDA.n1677 GNDA.n1676 16.0005
R3697 GNDA.n1676 GNDA.n1582 16.0005
R3698 GNDA.n1671 GNDA.n1582 16.0005
R3699 GNDA.n1671 GNDA.n1670 16.0005
R3700 GNDA.n1670 GNDA.n1669 16.0005
R3701 GNDA.n1665 GNDA.n1664 16.0005
R3702 GNDA.n1664 GNDA.n1585 16.0005
R3703 GNDA.n1045 GNDA.n1044 16.0005
R3704 GNDA.n1044 GNDA.n1043 16.0005
R3705 GNDA.n1043 GNDA.n1041 16.0005
R3706 GNDA.n1041 GNDA.n1038 16.0005
R3707 GNDA.n1038 GNDA.n1037 16.0005
R3708 GNDA.n1037 GNDA.n1034 16.0005
R3709 GNDA.n1034 GNDA.n1033 16.0005
R3710 GNDA.n1033 GNDA.n1031 16.0005
R3711 GNDA.n1016 GNDA.n1013 16.0005
R3712 GNDA.n1017 GNDA.n1016 16.0005
R3713 GNDA.n1020 GNDA.n1017 16.0005
R3714 GNDA.n1021 GNDA.n1020 16.0005
R3715 GNDA.n1024 GNDA.n1021 16.0005
R3716 GNDA.n1025 GNDA.n1024 16.0005
R3717 GNDA.n1028 GNDA.n1025 16.0005
R3718 GNDA.n1030 GNDA.n1028 16.0005
R3719 GNDA.n997 GNDA.n996 16.0005
R3720 GNDA.n1000 GNDA.n997 16.0005
R3721 GNDA.n1001 GNDA.n1000 16.0005
R3722 GNDA.n1004 GNDA.n1001 16.0005
R3723 GNDA.n1005 GNDA.n1004 16.0005
R3724 GNDA.n1009 GNDA.n1008 16.0005
R3725 GNDA.n1012 GNDA.n1009 16.0005
R3726 GNDA.n2296 GNDA.n380 15.5383
R3727 GNDA.n2393 GNDA.n2392 15.5383
R3728 GNDA.n414 GNDA.n370 15.5383
R3729 GNDA.n2352 GNDA.n2351 15.5383
R3730 GNDA.n1517 GNDA.n822 15.363
R3731 GNDA.n1499 GNDA.n822 15.363
R3732 GNDA.t293 GNDA.t339 14.992
R3733 GNDA.t33 GNDA.t202 14.992
R3734 GNDA.t190 GNDA.t17 14.992
R3735 GNDA.t341 GNDA.t203 14.992
R3736 GNDA.t7 GNDA.t340 14.992
R3737 GNDA.t188 GNDA.t308 14.992
R3738 GNDA.t308 GNDA.t330 14.992
R3739 GNDA.t330 GNDA.t85 14.992
R3740 GNDA.t342 GNDA.t81 14.992
R3741 GNDA.t81 GNDA.t168 14.992
R3742 GNDA.t171 GNDA.t155 14.992
R3743 GNDA.t155 GNDA.t148 14.992
R3744 GNDA.t148 GNDA.t53 14.992
R3745 GNDA.t112 GNDA.t77 14.992
R3746 GNDA.t77 GNDA.t350 14.992
R3747 GNDA.t350 GNDA.t235 14.992
R3748 GNDA.t93 GNDA.t23 14.992
R3749 GNDA.t23 GNDA.t68 14.992
R3750 GNDA.t347 GNDA.t356 14.992
R3751 GNDA.t356 GNDA.t147 14.992
R3752 GNDA.t118 GNDA.t59 14.992
R3753 GNDA.t59 GNDA.t317 14.992
R3754 GNDA.t266 GNDA.t55 14.992
R3755 GNDA.t349 GNDA.t153 14.992
R3756 GNDA.t63 GNDA.t286 14.992
R3757 GNDA.t305 GNDA.t214 14.992
R3758 GNDA.t346 GNDA.t345 14.992
R3759 GNDA.t336 GNDA.t329 14.992
R3760 GNDA.t360 GNDA.t143 14.992
R3761 GNDA.t344 GNDA.t211 14.992
R3762 GNDA.t335 GNDA.t50 14.992
R3763 GNDA.t338 GNDA.t327 14.992
R3764 GNDA.t328 GNDA.t322 14.992
R3765 GNDA.n726 GNDA.n562 14.9411
R3766 GNDA.n796 GNDA.n795 14.0505
R3767 GNDA.n659 GNDA.n658 14.0505
R3768 GNDA.n776 GNDA.n775 14.0193
R3769 GNDA.n427 GNDA.n375 13.9984
R3770 GNDA.n1491 GNDA.n849 13.8005
R3771 GNDA.n591 GNDA.n520 13.8005
R3772 GNDA.n702 GNDA.n701 13.8005
R3773 GNDA.n678 GNDA.n560 13.8005
R3774 GNDA.n675 GNDA.n561 13.8005
R3775 GNDA.n483 GNDA.t105 13.702
R3776 GNDA.n2516 GNDA.n2515 13.4945
R3777 GNDA GNDA.n321 12.9783
R3778 GNDA.n900 GNDA 12.9783
R3779 GNDA.n1372 GNDA 12.9783
R3780 GNDA.n2103 GNDA 12.9783
R3781 GNDA GNDA.n167 12.9783
R3782 GNDA.n1803 GNDA 12.9783
R3783 GNDA.n2216 GNDA 12.9783
R3784 GNDA.n1665 GNDA 12.9783
R3785 GNDA.n1008 GNDA 12.9783
R3786 GNDA.n612 GNDA.n611 12.8005
R3787 GNDA.n502 GNDA.n501 12.8005
R3788 GNDA.t120 GNDA.t27 12.5361
R3789 GNDA.t279 GNDA.t165 12.5361
R3790 GNDA.t175 GNDA.n1502 12.5361
R3791 GNDA.n1524 GNDA.t355 12.5361
R3792 GNDA.t296 GNDA.t99 12.5361
R3793 GNDA.t192 GNDA.t40 12.5361
R3794 GNDA.t217 GNDA.n1514 12.5361
R3795 GNDA.n1726 GNDA.n463 12.4126
R3796 GNDA.n1904 GNDA.n1702 12.4126
R3797 GNDA.n1252 GNDA.n1239 12.4126
R3798 GNDA.n2446 GNDA.n36 11.6369
R3799 GNDA.n2453 GNDA.n36 11.6369
R3800 GNDA.n2454 GNDA.n2453 11.6369
R3801 GNDA.n2455 GNDA.n2454 11.6369
R3802 GNDA.n2455 GNDA.n33 11.6369
R3803 GNDA.n2461 GNDA.n33 11.6369
R3804 GNDA.n2462 GNDA.n2461 11.6369
R3805 GNDA.n2463 GNDA.n2462 11.6369
R3806 GNDA.n2463 GNDA.n29 11.6369
R3807 GNDA.n1721 GNDA.n1717 11.6369
R3808 GNDA.n1756 GNDA.n1721 11.6369
R3809 GNDA.n1756 GNDA.n1755 11.6369
R3810 GNDA.n1755 GNDA.n1754 11.6369
R3811 GNDA.n1748 GNDA.n1725 11.6369
R3812 GNDA.n1748 GNDA.n1747 11.6369
R3813 GNDA.n1747 GNDA.n1746 11.6369
R3814 GNDA.n1746 GNDA.n1726 11.6369
R3815 GNDA.n1943 GNDA.n1942 11.6369
R3816 GNDA.n1944 GNDA.n1943 11.6369
R3817 GNDA.n1944 GNDA.n459 11.6369
R3818 GNDA.n1951 GNDA.n459 11.6369
R3819 GNDA.n1952 GNDA.n1951 11.6369
R3820 GNDA.n1953 GNDA.n1952 11.6369
R3821 GNDA.n1953 GNDA.n456 11.6369
R3822 GNDA.n1959 GNDA.n456 11.6369
R3823 GNDA.n1960 GNDA.n1959 11.6369
R3824 GNDA.n1962 GNDA.n1960 11.6369
R3825 GNDA.n1962 GNDA.n1961 11.6369
R3826 GNDA.n1977 GNDA.n1969 11.6369
R3827 GNDA.n1977 GNDA.n1976 11.6369
R3828 GNDA.n1976 GNDA.n1975 11.6369
R3829 GNDA.n1975 GNDA.n1970 11.6369
R3830 GNDA.n1970 GNDA.n6 11.6369
R3831 GNDA.n2508 GNDA.n7 11.6369
R3832 GNDA.n2502 GNDA.n7 11.6369
R3833 GNDA.n2502 GNDA.n2501 11.6369
R3834 GNDA.n2501 GNDA.n2500 11.6369
R3835 GNDA.n2500 GNDA.n12 11.6369
R3836 GNDA.n2487 GNDA.n20 11.6369
R3837 GNDA.n2487 GNDA.n2486 11.6369
R3838 GNDA.n2486 GNDA.n2485 11.6369
R3839 GNDA.n2485 GNDA.n21 11.6369
R3840 GNDA.n2479 GNDA.n21 11.6369
R3841 GNDA.n2479 GNDA.n2478 11.6369
R3842 GNDA.n2478 GNDA.n2477 11.6369
R3843 GNDA.n2477 GNDA.n24 11.6369
R3844 GNDA.n2471 GNDA.n24 11.6369
R3845 GNDA.n2471 GNDA.n2470 11.6369
R3846 GNDA.n2470 GNDA.n2469 11.6369
R3847 GNDA.n2303 GNDA.n2302 11.6369
R3848 GNDA.n2306 GNDA.n2303 11.6369
R3849 GNDA.n2307 GNDA.n2306 11.6369
R3850 GNDA.n2310 GNDA.n2307 11.6369
R3851 GNDA.n2311 GNDA.n2310 11.6369
R3852 GNDA.n2314 GNDA.n2311 11.6369
R3853 GNDA.n2316 GNDA.n2314 11.6369
R3854 GNDA.n2317 GNDA.n2316 11.6369
R3855 GNDA.n2319 GNDA.n2317 11.6369
R3856 GNDA.n2319 GNDA.n2318 11.6369
R3857 GNDA.n2318 GNDA.n69 11.6369
R3858 GNDA.n1697 GNDA.n1694 11.6369
R3859 GNDA.n1920 GNDA.n1697 11.6369
R3860 GNDA.n1920 GNDA.n1919 11.6369
R3861 GNDA.n1919 GNDA.n1918 11.6369
R3862 GNDA.n1912 GNDA.n1701 11.6369
R3863 GNDA.n1912 GNDA.n1911 11.6369
R3864 GNDA.n1911 GNDA.n1910 11.6369
R3865 GNDA.n1910 GNDA.n1702 11.6369
R3866 GNDA.n1903 GNDA.n1902 11.6369
R3867 GNDA.n1902 GNDA.n1707 11.6369
R3868 GNDA.n1861 GNDA.n1707 11.6369
R3869 GNDA.n1862 GNDA.n1861 11.6369
R3870 GNDA.n1863 GNDA.n1862 11.6369
R3871 GNDA.n1863 GNDA.n1847 11.6369
R3872 GNDA.n1883 GNDA.n1847 11.6369
R3873 GNDA.n1884 GNDA.n1883 11.6369
R3874 GNDA.n1886 GNDA.n1884 11.6369
R3875 GNDA.n1886 GNDA.n1885 11.6369
R3876 GNDA.n1885 GNDA.n409 11.6369
R3877 GNDA.n1132 GNDA.n1077 11.6369
R3878 GNDA.n1132 GNDA.n1131 11.6369
R3879 GNDA.n1131 GNDA.n1130 11.6369
R3880 GNDA.n1130 GNDA.n1082 11.6369
R3881 GNDA.n1086 GNDA.n1082 11.6369
R3882 GNDA.n1122 GNDA.n1086 11.6369
R3883 GNDA.n1122 GNDA.n1121 11.6369
R3884 GNDA.n1121 GNDA.n1120 11.6369
R3885 GNDA.n1120 GNDA.n1087 11.6369
R3886 GNDA.n1411 GNDA.n1410 11.6369
R3887 GNDA.n1414 GNDA.n1411 11.6369
R3888 GNDA.n1415 GNDA.n1414 11.6369
R3889 GNDA.n1418 GNDA.n1415 11.6369
R3890 GNDA.n1419 GNDA.n1418 11.6369
R3891 GNDA.n1422 GNDA.n1419 11.6369
R3892 GNDA.n1424 GNDA.n1422 11.6369
R3893 GNDA.n1425 GNDA.n1424 11.6369
R3894 GNDA.n1427 GNDA.n1425 11.6369
R3895 GNDA.n1427 GNDA.n1426 11.6369
R3896 GNDA.n1426 GNDA.n379 11.6369
R3897 GNDA.n1268 GNDA.n1245 11.6369
R3898 GNDA.n1268 GNDA.n1267 11.6369
R3899 GNDA.n1267 GNDA.n1266 11.6369
R3900 GNDA.n1266 GNDA.n1248 11.6369
R3901 GNDA.n1260 GNDA.n1259 11.6369
R3902 GNDA.n1259 GNDA.n1258 11.6369
R3903 GNDA.n1258 GNDA.n1253 11.6369
R3904 GNDA.n1253 GNDA.n1252 11.6369
R3905 GNDA.n2295 GNDA.n2294 11.6369
R3906 GNDA.n2294 GNDA.n381 11.6369
R3907 GNDA.n2289 GNDA.n381 11.6369
R3908 GNDA.n2289 GNDA.n2288 11.6369
R3909 GNDA.n2288 GNDA.n2287 11.6369
R3910 GNDA.n2287 GNDA.n2274 11.6369
R3911 GNDA.n2282 GNDA.n2274 11.6369
R3912 GNDA.n2282 GNDA.n2281 11.6369
R3913 GNDA.n2281 GNDA.n2280 11.6369
R3914 GNDA.n2280 GNDA.n223 11.6369
R3915 GNDA.n2353 GNDA.n223 11.6369
R3916 GNDA.n1096 GNDA.n224 11.6369
R3917 GNDA.n1097 GNDA.n1096 11.6369
R3918 GNDA.n1097 GNDA.n1092 11.6369
R3919 GNDA.n1103 GNDA.n1092 11.6369
R3920 GNDA.n1104 GNDA.n1103 11.6369
R3921 GNDA.n1105 GNDA.n1104 11.6369
R3922 GNDA.n1105 GNDA.n1090 11.6369
R3923 GNDA.n1111 GNDA.n1090 11.6369
R3924 GNDA.n1112 GNDA.n1111 11.6369
R3925 GNDA.n1113 GNDA.n1112 11.6369
R3926 GNDA.n1113 GNDA.n1088 11.6369
R3927 GNDA.n2437 GNDA.n53 11.6369
R3928 GNDA.n2431 GNDA.n53 11.6369
R3929 GNDA.n2431 GNDA.n2430 11.6369
R3930 GNDA.n2430 GNDA.n2429 11.6369
R3931 GNDA.n2429 GNDA.n57 11.6369
R3932 GNDA.n2423 GNDA.n57 11.6369
R3933 GNDA.n2423 GNDA.n2422 11.6369
R3934 GNDA.n2422 GNDA.n2421 11.6369
R3935 GNDA.n2421 GNDA.n61 11.6369
R3936 GNDA.n2394 GNDA.n67 11.6369
R3937 GNDA.n2400 GNDA.n67 11.6369
R3938 GNDA.n2401 GNDA.n2400 11.6369
R3939 GNDA.n2402 GNDA.n2401 11.6369
R3940 GNDA.n2402 GNDA.n65 11.6369
R3941 GNDA.n2408 GNDA.n65 11.6369
R3942 GNDA.n2409 GNDA.n2408 11.6369
R3943 GNDA.n2410 GNDA.n2409 11.6369
R3944 GNDA.n2410 GNDA.n63 11.6369
R3945 GNDA.n2415 GNDA.n63 11.6369
R3946 GNDA.n2416 GNDA.n2415 11.6369
R3947 GNDA.n674 GNDA.n673 11.6255
R3948 GNDA.n1717 GNDA.n1713 11.3514
R3949 GNDA.n1694 GNDA.n1692 11.3514
R3950 GNDA.n1275 GNDA.n1245 11.3514
R3951 GNDA.n2446 GNDA.n2445 11.249
R3952 GNDA.n1139 GNDA.n1077 11.249
R3953 GNDA.n2438 GNDA.n2437 11.249
R3954 GNDA.n740 GNDA.t337 11.2441
R3955 GNDA.t168 GNDA.n703 11.2441
R3956 GNDA.t162 GNDA.t201 11.2441
R3957 GNDA.n771 GNDA.t57 11.2441
R3958 GNDA.t259 GNDA.n642 11.2059
R3959 GNDA.t141 GNDA.t302 11.2059
R3960 GNDA.t97 GNDA.t132 11.2059
R3961 GNDA.t2 GNDA.t178 11.2059
R3962 GNDA.t144 GNDA.t243 11.2059
R3963 GNDA.t262 GNDA.n799 11.2059
R3964 GNDA.n2509 GNDA.n2508 10.4732
R3965 GNDA.n1725 GNDA 10.3439
R3966 GNDA.n1701 GNDA 10.3439
R3967 GNDA.n1260 GNDA 10.3439
R3968 GNDA.n1541 GNDA.n1540 9.78488
R3969 GNDA.n850 GNDA.t334 9.6005
R3970 GNDA.n850 GNDA.t332 9.6005
R3971 GNDA.n1490 GNDA.t333 9.6005
R3972 GNDA.n1490 GNDA.t331 9.6005
R3973 GNDA.n699 GNDA.t309 9.6005
R3974 GNDA.n699 GNDA.t82 9.6005
R3975 GNDA.n697 GNDA.t156 9.6005
R3976 GNDA.n697 GNDA.t78 9.6005
R3977 GNDA.n695 GNDA.t24 9.6005
R3978 GNDA.n695 GNDA.t357 9.6005
R3979 GNDA.n693 GNDA.t60 9.6005
R3980 GNDA.n693 GNDA.t56 9.6005
R3981 GNDA.n691 GNDA.t154 9.6005
R3982 GNDA.n691 GNDA.t64 9.6005
R3983 GNDA.n689 GNDA.t205 9.6005
R3984 GNDA.n689 GNDA.t66 9.6005
R3985 GNDA.n687 GNDA.t84 9.6005
R3986 GNDA.n687 GNDA.t158 9.6005
R3987 GNDA.n685 GNDA.t80 9.6005
R3988 GNDA.n685 GNDA.t26 9.6005
R3989 GNDA.n683 GNDA.t359 9.6005
R3990 GNDA.n683 GNDA.t152 9.6005
R3991 GNDA.n681 GNDA.t207 9.6005
R3992 GNDA.n681 GNDA.t62 9.6005
R3993 GNDA.n679 GNDA.t58 9.6005
R3994 GNDA.n679 GNDA.t273 9.6005
R3995 GNDA.n849 GNDA.n848 9.37925
R3996 GNDA.n753 GNDA.n752 9.3005
R3997 GNDA.n2299 GNDA.n375 8.98697
R3998 GNDA.n1942 GNDA.n463 8.79242
R3999 GNDA.n1904 GNDA.n1903 8.79242
R4000 GNDA.n1410 GNDA.n1239 8.79242
R4001 GNDA.n1969 GNDA.n452 8.53383
R4002 GNDA.n20 GNDA.n16 8.53383
R4003 GNDA.n2302 GNDA.n370 8.53383
R4004 GNDA.n2296 GNDA.n2295 8.53383
R4005 GNDA.n2352 GNDA.n224 8.53383
R4006 GNDA.n2394 GNDA.n2393 8.53383
R4007 GNDA.n250 GNDA.n247 8.35606
R4008 GNDA.n938 GNDA.n937 8.35606
R4009 GNDA.n1300 GNDA.n860 8.35606
R4010 GNDA.n2061 GNDA.n2034 8.35606
R4011 GNDA.n96 GNDA.n93 8.35606
R4012 GNDA.n1840 GNDA.n413 8.35606
R4013 GNDA.n2255 GNDA.n2253 8.35606
R4014 GNDA.n1623 GNDA.n1597 8.35606
R4015 GNDA.n1046 GNDA.n1045 8.35606
R4016 GNDA.n1457 GNDA.t229 8.20508
R4017 GNDA.n1966 GNDA.t238 8.20508
R4018 GNDA.n1540 GNDA.n822 7.71925
R4019 GNDA.n471 GNDA.n469 6.4005
R4020 GNDA.n1483 GNDA.t173 6.26831
R4021 GNDA.n1496 GNDA.n1495 6.26831
R4022 GNDA.n1515 GNDA.n1513 6.26831
R4023 GNDA.n846 GNDA.n845 6.0355
R4024 GNDA GNDA.n2516 5.86508
R4025 GNDA.n776 GNDA.n522 5.03175
R4026 GNDA.n673 GNDA.n522 4.90675
R4027 GNDA.n752 GNDA.n522 4.7505
R4028 GNDA.n1769 GNDA.n1768 4.6085
R4029 GNDA.n1691 GNDA.n1689 4.6085
R4030 GNDA.n1397 GNDA.n1396 4.6085
R4031 GNDA.n1560 GNDA.t20 4.56766
R4032 GNDA.t181 GNDA.n1559 4.56766
R4033 GNDA.n1930 GNDA.t138 4.56766
R4034 GNDA.n1984 GNDA.n1983 4.55161
R4035 GNDA.n2494 GNDA.n2493 4.55161
R4036 GNDA.n2133 GNDA.n372 4.55161
R4037 GNDA.n2297 GNDA.n378 4.55161
R4038 GNDA.n2356 GNDA.n220 4.55161
R4039 GNDA.n2326 GNDA.n70 4.55161
R4040 GNDA.n1540 GNDA.n1539 4.5005
R4041 GNDA.n751 GNDA.n749 4.5005
R4042 GNDA.n789 GNDA.n788 4.5005
R4043 GNDA.n791 GNDA.n790 4.5005
R4044 GNDA.n1961 GNDA.n452 4.39646
R4045 GNDA.n16 GNDA.n12 4.39646
R4046 GNDA.n2393 GNDA.n69 4.39646
R4047 GNDA.n409 GNDA.n370 4.39646
R4048 GNDA.n2296 GNDA.n379 4.39646
R4049 GNDA.n2353 GNDA.n2352 4.39646
R4050 GNDA.n2445 GNDA.n40 4.3013
R4051 GNDA.n2438 GNDA.n52 4.3013
R4052 GNDA.n2003 GNDA.n415 4.26717
R4053 GNDA.n2003 GNDA.n429 4.26717
R4054 GNDA.n1998 GNDA.n429 4.26717
R4055 GNDA.n1998 GNDA.n1997 4.26717
R4056 GNDA.n1997 GNDA.n1996 4.26717
R4057 GNDA.n1996 GNDA.n437 4.26717
R4058 GNDA.n1991 GNDA.n1990 4.26717
R4059 GNDA.n1990 GNDA.n1989 4.26717
R4060 GNDA.n1989 GNDA.n446 4.26717
R4061 GNDA.n1984 GNDA.n446 4.26717
R4062 GNDA.n2388 GNDA.n192 4.26717
R4063 GNDA.n195 GNDA.n192 4.26717
R4064 GNDA.n2381 GNDA.n195 4.26717
R4065 GNDA.n2381 GNDA.n2380 4.26717
R4066 GNDA.n2380 GNDA.n2379 4.26717
R4067 GNDA.n2379 GNDA.n200 4.26717
R4068 GNDA.n2374 GNDA.n2373 4.26717
R4069 GNDA.n2373 GNDA.n2372 4.26717
R4070 GNDA.n2372 GNDA.n14 4.26717
R4071 GNDA.n2494 GNDA.n14 4.26717
R4072 GNDA.n2154 GNDA.n392 4.26717
R4073 GNDA.n395 GNDA.n392 4.26717
R4074 GNDA.n2147 GNDA.n395 4.26717
R4075 GNDA.n2147 GNDA.n2146 4.26717
R4076 GNDA.n2146 GNDA.n2145 4.26717
R4077 GNDA.n2145 GNDA.n400 4.26717
R4078 GNDA.n2140 GNDA.n2139 4.26717
R4079 GNDA.n2139 GNDA.n2138 4.26717
R4080 GNDA.n2138 GNDA.n406 4.26717
R4081 GNDA.n2133 GNDA.n406 4.26717
R4082 GNDA.n1452 GNDA.n1451 4.26717
R4083 GNDA.n1451 GNDA.n1211 4.26717
R4084 GNDA.n1446 GNDA.n1211 4.26717
R4085 GNDA.n1446 GNDA.n1445 4.26717
R4086 GNDA.n1445 GNDA.n1444 4.26717
R4087 GNDA.n1444 GNDA.n1220 4.26717
R4088 GNDA.n1439 GNDA.n1438 4.26717
R4089 GNDA.n1438 GNDA.n1437 4.26717
R4090 GNDA.n1437 GNDA.n1231 4.26717
R4091 GNDA.n1231 GNDA.n378 4.26717
R4092 GNDA.n1190 GNDA.n1189 4.26717
R4093 GNDA.n1189 GNDA.n1159 4.26717
R4094 GNDA.n1184 GNDA.n1159 4.26717
R4095 GNDA.n1184 GNDA.n1183 4.26717
R4096 GNDA.n1183 GNDA.n1182 4.26717
R4097 GNDA.n1182 GNDA.n1166 4.26717
R4098 GNDA.n1177 GNDA.n1176 4.26717
R4099 GNDA.n1176 GNDA.n1175 4.26717
R4100 GNDA.n1175 GNDA.n219 4.26717
R4101 GNDA.n2356 GNDA.n219 4.26717
R4102 GNDA.n2347 GNDA.n345 4.26717
R4103 GNDA.n349 GNDA.n345 4.26717
R4104 GNDA.n2340 GNDA.n349 4.26717
R4105 GNDA.n2340 GNDA.n2339 4.26717
R4106 GNDA.n2339 GNDA.n2338 4.26717
R4107 GNDA.n2338 GNDA.n355 4.26717
R4108 GNDA.n2333 GNDA.n2332 4.26717
R4109 GNDA.n2332 GNDA.n2331 4.26717
R4110 GNDA.n2331 GNDA.n362 4.26717
R4111 GNDA.n2326 GNDA.n362 4.26717
R4112 GNDA.n1140 GNDA.n1139 4.1989
R4113 GNDA.n1539 GNDA.n849 3.813
R4114 GNDA.n1991 GNDA 3.79309
R4115 GNDA.n2374 GNDA 3.79309
R4116 GNDA.n2140 GNDA 3.79309
R4117 GNDA.n1439 GNDA 3.79309
R4118 GNDA.n1177 GNDA 3.79309
R4119 GNDA.n2333 GNDA 3.79309
R4120 GNDA.t250 GNDA.n730 3.74837
R4121 GNDA.n728 GNDA.t195 3.74837
R4122 GNDA.t202 GNDA.n739 3.74837
R4123 GNDA.n704 GNDA.t341 3.74837
R4124 GNDA.n703 GNDA.t103 3.74837
R4125 GNDA.n756 GNDA.t299 3.74837
R4126 GNDA.n588 GNDA.t18 3.74837
R4127 GNDA.t162 GNDA.t16 3.74837
R4128 GNDA.n634 GNDA.t15 3.73564
R4129 GNDA.n633 GNDA.t96 3.73564
R4130 GNDA.t269 GNDA.t290 3.73564
R4131 GNDA.t253 GNDA.t231 3.73564
R4132 GNDA.t70 GNDA.n496 3.72931
R4133 GNDA.n788 GNDA.n776 3.6255
R4134 GNDA.n184 GNDA.n74 3.5845
R4135 GNDA.n183 GNDA.n76 3.5845
R4136 GNDA.n106 GNDA.n104 3.5845
R4137 GNDA.n105 GNDA.n102 3.5845
R4138 GNDA.n113 GNDA.n112 3.5845
R4139 GNDA.n99 GNDA.n98 3.5845
R4140 GNDA.n121 GNDA.n119 3.5845
R4141 GNDA.n120 GNDA.n95 3.5845
R4142 GNDA.n128 GNDA.n127 3.5845
R4143 GNDA.n1897 GNDA.n1771 3.5845
R4144 GNDA.n1855 GNDA.n1854 3.5845
R4145 GNDA.n1868 GNDA.n1853 3.5845
R4146 GNDA.n1869 GNDA.n1851 3.5845
R4147 GNDA.n1873 GNDA.n1872 3.5845
R4148 GNDA.n1879 GNDA.n1874 3.5845
R4149 GNDA.n1878 GNDA.n1875 3.5845
R4150 GNDA.n1890 GNDA.n1843 3.5845
R4151 GNDA.n1892 GNDA.n1891 3.5845
R4152 GNDA.n2121 GNDA.n2015 3.5845
R4153 GNDA.n2120 GNDA.n2016 3.5845
R4154 GNDA.n2044 GNDA.n2042 3.5845
R4155 GNDA.n2048 GNDA.n2045 3.5845
R4156 GNDA.n2049 GNDA.n2037 3.5845
R4157 GNDA.n2054 GNDA.n2053 3.5845
R4158 GNDA.n2057 GNDA.n2036 3.5845
R4159 GNDA.n2059 GNDA.n2058 3.5845
R4160 GNDA.n2065 GNDA.n2064 3.5845
R4161 GNDA.n1683 GNDA.n1578 3.5845
R4162 GNDA.n1682 GNDA.n1579 3.5845
R4163 GNDA.n1607 GNDA.n1605 3.5845
R4164 GNDA.n1611 GNDA.n1608 3.5845
R4165 GNDA.n1612 GNDA.n1600 3.5845
R4166 GNDA.n1617 GNDA.n1616 3.5845
R4167 GNDA.n1620 GNDA.n1599 3.5845
R4168 GNDA.n1622 GNDA.n1621 3.5845
R4169 GNDA.n1627 GNDA.n1626 3.5845
R4170 GNDA.n2264 GNDA.n2158 3.5845
R4171 GNDA.n2185 GNDA.n2184 3.5845
R4172 GNDA.n2188 GNDA.n2183 3.5845
R4173 GNDA.n2192 GNDA.n2191 3.5845
R4174 GNDA.n2195 GNDA.n2181 3.5845
R4175 GNDA.n2199 GNDA.n2198 3.5845
R4176 GNDA.n2202 GNDA.n2180 3.5845
R4177 GNDA.n2204 GNDA.n2203 3.5845
R4178 GNDA.n2259 GNDA.n2258 3.5845
R4179 GNDA.n1150 GNDA.n973 3.5845
R4180 GNDA.n1054 GNDA.n1053 3.5845
R4181 GNDA.n1060 GNDA.n1056 3.5845
R4182 GNDA.n1059 GNDA.n1050 3.5845
R4183 GNDA.n1066 GNDA.n1049 3.5845
R4184 GNDA.n1067 GNDA.n1048 3.5845
R4185 GNDA.n1072 GNDA.n1070 3.5845
R4186 GNDA.n1071 GNDA.n995 3.5845
R4187 GNDA.n1145 GNDA.n1144 3.5845
R4188 GNDA.n1390 GNDA.n1281 3.5845
R4189 GNDA.n1389 GNDA.n1282 3.5845
R4190 GNDA.n1312 GNDA.n1311 3.5845
R4191 GNDA.n1317 GNDA.n1310 3.5845
R4192 GNDA.n1319 GNDA.n1318 3.5845
R4193 GNDA.n1326 GNDA.n1306 3.5845
R4194 GNDA.n1325 GNDA.n1307 3.5845
R4195 GNDA.n1332 GNDA.n1302 3.5845
R4196 GNDA.n1334 GNDA.n1333 3.5845
R4197 GNDA.n1202 GNDA.n865 3.5845
R4198 GNDA.n946 GNDA.n945 3.5845
R4199 GNDA.n952 GNDA.n948 3.5845
R4200 GNDA.n951 GNDA.n942 3.5845
R4201 GNDA.n958 GNDA.n941 3.5845
R4202 GNDA.n959 GNDA.n940 3.5845
R4203 GNDA.n964 GNDA.n962 3.5845
R4204 GNDA.n963 GNDA.n887 3.5845
R4205 GNDA.n1197 GNDA.n1196 3.5845
R4206 GNDA.n338 GNDA.n228 3.5845
R4207 GNDA.n337 GNDA.n230 3.5845
R4208 GNDA.n260 GNDA.n258 3.5845
R4209 GNDA.n259 GNDA.n256 3.5845
R4210 GNDA.n267 GNDA.n266 3.5845
R4211 GNDA.n253 GNDA.n252 3.5845
R4212 GNDA.n275 GNDA.n273 3.5845
R4213 GNDA.n274 GNDA.n249 3.5845
R4214 GNDA.n282 GNDA.n281 3.5845
R4215 GNDA.n660 GNDA.t39 3.42907
R4216 GNDA.n660 GNDA.t98 3.42907
R4217 GNDA.n792 GNDA.t3 3.42907
R4218 GNDA.n792 GNDA.t9 3.42907
R4219 GNDA.n794 GNDA.t90 3.42907
R4220 GNDA.n794 GNDA.t117 3.42907
R4221 GNDA.n592 GNDA.t110 3.42907
R4222 GNDA.n592 GNDA.t47 3.42907
R4223 GNDA.n189 GNDA.n71 3.3797
R4224 GNDA.n96 GNDA.n40 3.3797
R4225 GNDA.n2129 GNDA.n413 3.3797
R4226 GNDA.n2128 GNDA.n2127 3.3797
R4227 GNDA.n2061 GNDA.n2060 3.3797
R4228 GNDA.n1623 GNDA.n390 3.3797
R4229 GNDA.n2267 GNDA.n2155 3.3797
R4230 GNDA.n2255 GNDA.n2254 3.3797
R4231 GNDA.n1191 GNDA.n969 3.3797
R4232 GNDA.n1140 GNDA.n1046 3.3797
R4233 GNDA.n1454 GNDA.n860 3.3797
R4234 GNDA.n1453 GNDA.n861 3.3797
R4235 GNDA.n1192 GNDA.n938 3.3797
R4236 GNDA.n343 GNDA.n225 3.3797
R4237 GNDA.n250 GNDA.n52 3.3797
R4238 GNDA.n2128 GNDA.n414 3.27161
R4239 GNDA.n2392 GNDA.n71 3.27161
R4240 GNDA.n2155 GNDA.n380 3.27161
R4241 GNDA.n2351 GNDA.n225 3.27161
R4242 GNDA.n833 GNDA.n831 3.21925
R4243 GNDA.n841 GNDA.n839 3.21925
R4244 GNDA.n1557 GNDA.n1556 3.2005
R4245 GNDA.n481 GNDA.n472 3.2005
R4246 GNDA.n577 GNDA.t51 3.1344
R4247 GNDA.n579 GNDA.t150 3.1344
R4248 GNDA.n322 GNDA 3.02272
R4249 GNDA.n897 GNDA 3.02272
R4250 GNDA.n1376 GNDA 3.02272
R4251 GNDA.n2107 GNDA 3.02272
R4252 GNDA.n168 GNDA 3.02272
R4253 GNDA.n1800 GNDA 3.02272
R4254 GNDA.n2213 GNDA 3.02272
R4255 GNDA.n1669 GNDA 3.02272
R4256 GNDA.n1005 GNDA 3.02272
R4257 GNDA.n188 GNDA.n187 2.8677
R4258 GNDA.n1898 GNDA.n1770 2.8677
R4259 GNDA.n2014 GNDA.n416 2.8677
R4260 GNDA.n1577 GNDA.n1570 2.8677
R4261 GNDA.n2266 GNDA.n2265 2.8677
R4262 GNDA.n1151 GNDA.n972 2.8677
R4263 GNDA.n1280 GNDA.n1276 2.8677
R4264 GNDA.n1203 GNDA.n864 2.8677
R4265 GNDA.n342 GNDA.n341 2.8677
R4266 GNDA.n790 GNDA.n789 2.5005
R4267 GNDA.n342 GNDA.n227 2.31161
R4268 GNDA.n888 GNDA.n864 2.31161
R4269 GNDA.n1384 GNDA.n1276 2.31161
R4270 GNDA.n2115 GNDA.n416 2.31161
R4271 GNDA.n188 GNDA.n73 2.31161
R4272 GNDA.n1791 GNDA.n1770 2.31161
R4273 GNDA.n2266 GNDA.n2156 2.31161
R4274 GNDA.n1677 GNDA.n1570 2.31161
R4275 GNDA.n996 GNDA.n972 2.31161
R4276 GNDA.n793 GNDA.n791 2.063
R4277 GNDA.n2350 GNDA.n2349 1.951
R4278 GNDA.n1207 GNDA.n862 1.951
R4279 GNDA.n1767 GNDA.n1714 1.951
R4280 GNDA.n1690 GNDA.n1569 1.951
R4281 GNDA.n2007 GNDA.n373 1.951
R4282 GNDA.n2391 GNDA.n2390 1.951
R4283 GNDA.n389 GNDA.n374 1.951
R4284 GNDA.n1155 GNDA.n970 1.951
R4285 GNDA.n1398 GNDA.n1244 1.951
R4286 GNDA.n674 GNDA.n661 1.813
R4287 GNDA.n791 GNDA.n520 1.78175
R4288 GNDA.n675 GNDA.n674 1.78175
R4289 GNDA.n189 GNDA.n188 1.7413
R4290 GNDA.n1770 GNDA.n1769 1.7413
R4291 GNDA.n2129 GNDA.n2128 1.7413
R4292 GNDA.n2127 GNDA.n416 1.7413
R4293 GNDA.n2060 GNDA.n71 1.7413
R4294 GNDA.n1689 GNDA.n1570 1.7413
R4295 GNDA.n2155 GNDA.n390 1.7413
R4296 GNDA.n2267 GNDA.n2266 1.7413
R4297 GNDA.n2254 GNDA.n225 1.7413
R4298 GNDA.n972 GNDA.n969 1.7413
R4299 GNDA.n1396 GNDA.n1276 1.7413
R4300 GNDA.n1454 GNDA.n1453 1.7413
R4301 GNDA.n864 GNDA.n861 1.7413
R4302 GNDA.n1192 GNDA.n1191 1.7413
R4303 GNDA.n343 GNDA.n342 1.7413
R4304 GNDA.n2515 GNDA.n2 1.73362
R4305 GNDA.n2128 GNDA.n415 1.51754
R4306 GNDA.n2388 GNDA.n71 1.51754
R4307 GNDA.n2155 GNDA.n2154 1.51754
R4308 GNDA.n1453 GNDA.n1452 1.51754
R4309 GNDA.n1191 GNDA.n1190 1.51754
R4310 GNDA.n2347 GNDA.n225 1.51754
R4311 GNDA.n1754 GNDA 1.29343
R4312 GNDA.n1918 GNDA 1.29343
R4313 GNDA GNDA.n1248 1.29343
R4314 GNDA.n127 GNDA.n96 1.2293
R4315 GNDA.n1891 GNDA.n413 1.2293
R4316 GNDA.n2064 GNDA.n2061 1.2293
R4317 GNDA.n1626 GNDA.n1623 1.2293
R4318 GNDA.n2258 GNDA.n2255 1.2293
R4319 GNDA.n1144 GNDA.n1046 1.2293
R4320 GNDA.n1333 GNDA.n860 1.2293
R4321 GNDA.n1196 GNDA.n938 1.2293
R4322 GNDA.n281 GNDA.n250 1.2293
R4323 GNDA.n701 GNDA.n678 1.21925
R4324 GNDA.n1768 GNDA.n1713 1.1781
R4325 GNDA.n1692 GNDA.n1691 1.1781
R4326 GNDA.n1397 GNDA.n1275 1.1781
R4327 GNDA.n2509 GNDA.n6 1.16414
R4328 GNDA.n187 GNDA.n74 1.0245
R4329 GNDA.n184 GNDA.n183 1.0245
R4330 GNDA.n104 GNDA.n76 1.0245
R4331 GNDA.n106 GNDA.n105 1.0245
R4332 GNDA.n113 GNDA.n102 1.0245
R4333 GNDA.n112 GNDA.n99 1.0245
R4334 GNDA.n119 GNDA.n98 1.0245
R4335 GNDA.n121 GNDA.n120 1.0245
R4336 GNDA.n128 GNDA.n95 1.0245
R4337 GNDA.n1898 GNDA.n1897 1.0245
R4338 GNDA.n1854 GNDA.n1771 1.0245
R4339 GNDA.n1855 GNDA.n1853 1.0245
R4340 GNDA.n1869 GNDA.n1868 1.0245
R4341 GNDA.n1872 GNDA.n1851 1.0245
R4342 GNDA.n1874 GNDA.n1873 1.0245
R4343 GNDA.n1879 GNDA.n1878 1.0245
R4344 GNDA.n1875 GNDA.n1843 1.0245
R4345 GNDA.n1892 GNDA.n1890 1.0245
R4346 GNDA.n2015 GNDA.n2014 1.0245
R4347 GNDA.n2121 GNDA.n2120 1.0245
R4348 GNDA.n2042 GNDA.n2016 1.0245
R4349 GNDA.n2045 GNDA.n2044 1.0245
R4350 GNDA.n2049 GNDA.n2048 1.0245
R4351 GNDA.n2053 GNDA.n2037 1.0245
R4352 GNDA.n2054 GNDA.n2036 1.0245
R4353 GNDA.n2058 GNDA.n2057 1.0245
R4354 GNDA.n2065 GNDA.n2059 1.0245
R4355 GNDA.n1578 GNDA.n1577 1.0245
R4356 GNDA.n1683 GNDA.n1682 1.0245
R4357 GNDA.n1605 GNDA.n1579 1.0245
R4358 GNDA.n1608 GNDA.n1607 1.0245
R4359 GNDA.n1612 GNDA.n1611 1.0245
R4360 GNDA.n1616 GNDA.n1600 1.0245
R4361 GNDA.n1617 GNDA.n1599 1.0245
R4362 GNDA.n1621 GNDA.n1620 1.0245
R4363 GNDA.n1627 GNDA.n1622 1.0245
R4364 GNDA.n2265 GNDA.n2264 1.0245
R4365 GNDA.n2184 GNDA.n2158 1.0245
R4366 GNDA.n2185 GNDA.n2183 1.0245
R4367 GNDA.n2191 GNDA.n2188 1.0245
R4368 GNDA.n2192 GNDA.n2181 1.0245
R4369 GNDA.n2198 GNDA.n2195 1.0245
R4370 GNDA.n2199 GNDA.n2180 1.0245
R4371 GNDA.n2203 GNDA.n2202 1.0245
R4372 GNDA.n2259 GNDA.n2204 1.0245
R4373 GNDA.n1151 GNDA.n1150 1.0245
R4374 GNDA.n1053 GNDA.n973 1.0245
R4375 GNDA.n1056 GNDA.n1054 1.0245
R4376 GNDA.n1060 GNDA.n1059 1.0245
R4377 GNDA.n1050 GNDA.n1049 1.0245
R4378 GNDA.n1067 GNDA.n1066 1.0245
R4379 GNDA.n1070 GNDA.n1048 1.0245
R4380 GNDA.n1072 GNDA.n1071 1.0245
R4381 GNDA.n1145 GNDA.n995 1.0245
R4382 GNDA.n1281 GNDA.n1280 1.0245
R4383 GNDA.n1390 GNDA.n1389 1.0245
R4384 GNDA.n1311 GNDA.n1282 1.0245
R4385 GNDA.n1312 GNDA.n1310 1.0245
R4386 GNDA.n1319 GNDA.n1317 1.0245
R4387 GNDA.n1318 GNDA.n1306 1.0245
R4388 GNDA.n1326 GNDA.n1325 1.0245
R4389 GNDA.n1307 GNDA.n1302 1.0245
R4390 GNDA.n1334 GNDA.n1332 1.0245
R4391 GNDA.n1203 GNDA.n1202 1.0245
R4392 GNDA.n945 GNDA.n865 1.0245
R4393 GNDA.n948 GNDA.n946 1.0245
R4394 GNDA.n952 GNDA.n951 1.0245
R4395 GNDA.n942 GNDA.n941 1.0245
R4396 GNDA.n959 GNDA.n958 1.0245
R4397 GNDA.n962 GNDA.n940 1.0245
R4398 GNDA.n964 GNDA.n963 1.0245
R4399 GNDA.n1197 GNDA.n887 1.0245
R4400 GNDA.n341 GNDA.n228 1.0245
R4401 GNDA.n338 GNDA.n337 1.0245
R4402 GNDA.n258 GNDA.n230 1.0245
R4403 GNDA.n260 GNDA.n259 1.0245
R4404 GNDA.n267 GNDA.n256 1.0245
R4405 GNDA.n266 GNDA.n253 1.0245
R4406 GNDA.n273 GNDA.n252 1.0245
R4407 GNDA.n275 GNDA.n274 1.0245
R4408 GNDA.n282 GNDA.n249 1.0245
R4409 GNDA.n831 GNDA.n829 1.0005
R4410 GNDA.n835 GNDA.n833 1.0005
R4411 GNDA.n837 GNDA.n835 1.0005
R4412 GNDA.n839 GNDA.n837 1.0005
R4413 GNDA.n843 GNDA.n841 1.0005
R4414 GNDA.n845 GNDA.n843 1.0005
R4415 GNDA.n678 GNDA.n677 0.6255
R4416 GNDA.n618 GNDA.t142 0.571187
R4417 GNDA.n781 GNDA.n779 0.563
R4418 GNDA.n783 GNDA.n781 0.563
R4419 GNDA.n785 GNDA.n783 0.563
R4420 GNDA.n787 GNDA.n785 0.563
R4421 GNDA.n749 GNDA.n748 0.563
R4422 GNDA.n749 GNDA.n745 0.563
R4423 GNDA.n666 GNDA.n664 0.563
R4424 GNDA.n668 GNDA.n666 0.563
R4425 GNDA.n670 GNDA.n668 0.563
R4426 GNDA.n672 GNDA.n670 0.563
R4427 GNDA.n682 GNDA.n680 0.563
R4428 GNDA.n684 GNDA.n682 0.563
R4429 GNDA.n686 GNDA.n684 0.563
R4430 GNDA.n688 GNDA.n686 0.563
R4431 GNDA.n690 GNDA.n688 0.563
R4432 GNDA.n692 GNDA.n690 0.563
R4433 GNDA.n694 GNDA.n692 0.563
R4434 GNDA.n696 GNDA.n694 0.563
R4435 GNDA.n698 GNDA.n696 0.563
R4436 GNDA.n700 GNDA.n698 0.563
R4437 GNDA.n795 GNDA.n793 0.5005
R4438 GNDA.n661 GNDA.n659 0.5005
R4439 GNDA GNDA.n437 0.474574
R4440 GNDA GNDA.n200 0.474574
R4441 GNDA GNDA.n400 0.474574
R4442 GNDA GNDA.n1220 0.474574
R4443 GNDA GNDA.n1166 0.474574
R4444 GNDA GNDA.n355 0.474574
R4445 GNDA.n826 GNDA.n824 0.4705
R4446 GNDA.n824 GNDA.n823 0.311875
R4447 GNDA.n680 GNDA.n520 0.28175
R4448 GNDA.n848 GNDA.n847 0.276625
R4449 GNDA.n2516 GNDA.n1 0.276625
R4450 GNDA.n752 GNDA.n751 0.2505
R4451 GNDA.n701 GNDA.n700 0.2505
R4452 GNDA.n677 GNDA.n675 0.2505
R4453 GNDA.n847 GNDA.n846 0.22375
R4454 GNDA.n846 GNDA.n1 0.100375
R4455 GNDA.n1983 GNDA.n452 0.0953148
R4456 GNDA.n2493 GNDA.n16 0.0953148
R4457 GNDA.n372 GNDA.n370 0.0953148
R4458 GNDA.n2297 GNDA.n2296 0.0953148
R4459 GNDA.n2352 GNDA.n220 0.0953148
R4460 GNDA.n2393 GNDA.n70 0.0953148
R4461 GNDA.n823 GNDA.n2 0.076875
R4462 ref_volt_cur_gen_dummy_magic_0.V_mir2.n5 ref_volt_cur_gen_dummy_magic_0.V_mir2.n1 325.473
R4463 ref_volt_cur_gen_dummy_magic_0.V_mir2.n10 ref_volt_cur_gen_dummy_magic_0.V_mir2.n6 325.471
R4464 ref_volt_cur_gen_dummy_magic_0.V_mir2.n19 ref_volt_cur_gen_dummy_magic_0.V_mir2.n18 325.471
R4465 ref_volt_cur_gen_dummy_magic_0.V_mir2.n15 ref_volt_cur_gen_dummy_magic_0.V_mir2.t18 310.488
R4466 ref_volt_cur_gen_dummy_magic_0.V_mir2.n7 ref_volt_cur_gen_dummy_magic_0.V_mir2.t22 310.488
R4467 ref_volt_cur_gen_dummy_magic_0.V_mir2.n2 ref_volt_cur_gen_dummy_magic_0.V_mir2.t20 310.488
R4468 ref_volt_cur_gen_dummy_magic_0.V_mir2.n13 ref_volt_cur_gen_dummy_magic_0.V_mir2.t1 278.312
R4469 ref_volt_cur_gen_dummy_magic_0.V_mir2.n13 ref_volt_cur_gen_dummy_magic_0.V_mir2.n12 228.939
R4470 ref_volt_cur_gen_dummy_magic_0.V_mir2.n0 ref_volt_cur_gen_dummy_magic_0.V_mir2.n11 224.439
R4471 ref_volt_cur_gen_dummy_magic_0.V_mir2.n17 ref_volt_cur_gen_dummy_magic_0.V_mir2.t5 184.097
R4472 ref_volt_cur_gen_dummy_magic_0.V_mir2.n9 ref_volt_cur_gen_dummy_magic_0.V_mir2.t7 184.097
R4473 ref_volt_cur_gen_dummy_magic_0.V_mir2.n4 ref_volt_cur_gen_dummy_magic_0.V_mir2.t15 184.097
R4474 ref_volt_cur_gen_dummy_magic_0.V_mir2.n16 ref_volt_cur_gen_dummy_magic_0.V_mir2.n15 167.094
R4475 ref_volt_cur_gen_dummy_magic_0.V_mir2.n8 ref_volt_cur_gen_dummy_magic_0.V_mir2.n7 167.094
R4476 ref_volt_cur_gen_dummy_magic_0.V_mir2.n3 ref_volt_cur_gen_dummy_magic_0.V_mir2.n2 167.094
R4477 ref_volt_cur_gen_dummy_magic_0.V_mir2.n10 ref_volt_cur_gen_dummy_magic_0.V_mir2.n9 152
R4478 ref_volt_cur_gen_dummy_magic_0.V_mir2.n5 ref_volt_cur_gen_dummy_magic_0.V_mir2.n4 152
R4479 ref_volt_cur_gen_dummy_magic_0.V_mir2.n18 ref_volt_cur_gen_dummy_magic_0.V_mir2.n17 152
R4480 ref_volt_cur_gen_dummy_magic_0.V_mir2.n15 ref_volt_cur_gen_dummy_magic_0.V_mir2.t17 120.501
R4481 ref_volt_cur_gen_dummy_magic_0.V_mir2.n16 ref_volt_cur_gen_dummy_magic_0.V_mir2.t9 120.501
R4482 ref_volt_cur_gen_dummy_magic_0.V_mir2.n7 ref_volt_cur_gen_dummy_magic_0.V_mir2.t21 120.501
R4483 ref_volt_cur_gen_dummy_magic_0.V_mir2.n8 ref_volt_cur_gen_dummy_magic_0.V_mir2.t13 120.501
R4484 ref_volt_cur_gen_dummy_magic_0.V_mir2.n2 ref_volt_cur_gen_dummy_magic_0.V_mir2.t19 120.501
R4485 ref_volt_cur_gen_dummy_magic_0.V_mir2.n3 ref_volt_cur_gen_dummy_magic_0.V_mir2.t11 120.501
R4486 ref_volt_cur_gen_dummy_magic_0.V_mir2.n12 ref_volt_cur_gen_dummy_magic_0.V_mir2.t2 48.0005
R4487 ref_volt_cur_gen_dummy_magic_0.V_mir2.n12 ref_volt_cur_gen_dummy_magic_0.V_mir2.t3 48.0005
R4488 ref_volt_cur_gen_dummy_magic_0.V_mir2.n11 ref_volt_cur_gen_dummy_magic_0.V_mir2.t0 48.0005
R4489 ref_volt_cur_gen_dummy_magic_0.V_mir2.n11 ref_volt_cur_gen_dummy_magic_0.V_mir2.t4 48.0005
R4490 ref_volt_cur_gen_dummy_magic_0.V_mir2.n17 ref_volt_cur_gen_dummy_magic_0.V_mir2.n16 40.7027
R4491 ref_volt_cur_gen_dummy_magic_0.V_mir2.n9 ref_volt_cur_gen_dummy_magic_0.V_mir2.n8 40.7027
R4492 ref_volt_cur_gen_dummy_magic_0.V_mir2.n4 ref_volt_cur_gen_dummy_magic_0.V_mir2.n3 40.7027
R4493 ref_volt_cur_gen_dummy_magic_0.V_mir2.n6 ref_volt_cur_gen_dummy_magic_0.V_mir2.t8 39.4005
R4494 ref_volt_cur_gen_dummy_magic_0.V_mir2.n6 ref_volt_cur_gen_dummy_magic_0.V_mir2.t14 39.4005
R4495 ref_volt_cur_gen_dummy_magic_0.V_mir2.n1 ref_volt_cur_gen_dummy_magic_0.V_mir2.t16 39.4005
R4496 ref_volt_cur_gen_dummy_magic_0.V_mir2.n1 ref_volt_cur_gen_dummy_magic_0.V_mir2.t12 39.4005
R4497 ref_volt_cur_gen_dummy_magic_0.V_mir2.t6 ref_volt_cur_gen_dummy_magic_0.V_mir2.n19 39.4005
R4498 ref_volt_cur_gen_dummy_magic_0.V_mir2.n19 ref_volt_cur_gen_dummy_magic_0.V_mir2.t10 39.4005
R4499 ref_volt_cur_gen_dummy_magic_0.V_mir2.n14 ref_volt_cur_gen_dummy_magic_0.V_mir2.n5 15.8005
R4500 ref_volt_cur_gen_dummy_magic_0.V_mir2.n18 ref_volt_cur_gen_dummy_magic_0.V_mir2.n14 15.8005
R4501 ref_volt_cur_gen_dummy_magic_0.V_mir2.n0 ref_volt_cur_gen_dummy_magic_0.V_mir2.n10 9.3005
R4502 ref_volt_cur_gen_dummy_magic_0.V_mir2.n0 ref_volt_cur_gen_dummy_magic_0.V_mir2.n13 5.8755
R4503 ref_volt_cur_gen_dummy_magic_0.V_mir2.n14 ref_volt_cur_gen_dummy_magic_0.V_mir2.n0 5.28175
R4504 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t32 354.854
R4505 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t22 346.8
R4506 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n11 339.522
R4507 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n4 339.522
R4508 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n6 335.022
R4509 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n8 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t4 275.909
R4510 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n8 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n7 227.909
R4511 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n9 222.034
R4512 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n10 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t19 184.097
R4513 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n10 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t14 184.097
R4514 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n5 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t15 184.097
R4515 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n5 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t12 184.097
R4516 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n10 166.05
R4517 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n5 166.05
R4518 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 58.0259
R4519 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n9 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t0 48.0005
R4520 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n9 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t3 48.0005
R4521 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n7 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t2 48.0005
R4522 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n7 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t1 48.0005
R4523 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t8 39.4005
R4524 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t6 39.4005
R4525 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n4 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t10 39.4005
R4526 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n4 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t7 39.4005
R4527 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n11 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t9 39.4005
R4528 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n11 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t5 39.4005
R4529 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n0 5.6255
R4530 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n3 5.28175
R4531 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t11 4.8295
R4532 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t28 4.8295
R4533 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t18 4.8295
R4534 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t34 4.8295
R4535 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t36 4.8295
R4536 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t27 4.8295
R4537 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t21 4.8295
R4538 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n8 4.5005
R4539 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t20 4.5005
R4540 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t26 4.5005
R4541 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t33 4.5005
R4542 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t25 4.5005
R4543 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t31 4.5005
R4544 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t13 4.5005
R4545 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t17 4.5005
R4546 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t24 4.5005
R4547 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t30 4.5005
R4548 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t29 4.5005
R4549 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t35 4.5005
R4550 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t16 4.5005
R4551 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t23 4.5005
R4552 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 3.8075
R4553 VDDA.n348 VDDA.n344 6600
R4554 VDDA.n348 VDDA.n345 6600
R4555 VDDA.n350 VDDA.n344 6570
R4556 VDDA.n350 VDDA.n345 6570
R4557 VDDA.n434 VDDA.n381 4710
R4558 VDDA.n434 VDDA.n382 4710
R4559 VDDA.n432 VDDA.n381 4710
R4560 VDDA.n432 VDDA.n382 4710
R4561 VDDA.n410 VDDA.n403 4710
R4562 VDDA.n412 VDDA.n403 4710
R4563 VDDA.n410 VDDA.n409 4710
R4564 VDDA.n412 VDDA.n409 4710
R4565 VDDA.n141 VDDA.n137 4605
R4566 VDDA.n141 VDDA.n138 4605
R4567 VDDA.n42 VDDA.n28 4605
R4568 VDDA.n44 VDDA.n28 4605
R4569 VDDA.n206 VDDA.n182 4590
R4570 VDDA.n208 VDDA.n182 4590
R4571 VDDA.n208 VDDA.n183 4590
R4572 VDDA.n206 VDDA.n183 4590
R4573 VDDA.n143 VDDA.n137 4575
R4574 VDDA.n143 VDDA.n138 4575
R4575 VDDA.n42 VDDA.n29 4575
R4576 VDDA.n44 VDDA.n29 4575
R4577 VDDA.n282 VDDA.n275 4500
R4578 VDDA.n284 VDDA.n275 4500
R4579 VDDA.n282 VDDA.n276 4350
R4580 VDDA.n284 VDDA.n276 4350
R4581 VDDA.n101 VDDA.n94 4020
R4582 VDDA.n103 VDDA.n94 4020
R4583 VDDA.n101 VDDA.n100 4020
R4584 VDDA.n103 VDDA.n100 4020
R4585 VDDA.n77 VDDA.n70 4020
R4586 VDDA.n79 VDDA.n70 4020
R4587 VDDA.n77 VDDA.n76 4020
R4588 VDDA.n79 VDDA.n76 4020
R4589 VDDA.n121 VDDA.n114 3390
R4590 VDDA.n123 VDDA.n114 3390
R4591 VDDA.n121 VDDA.n120 3390
R4592 VDDA.n123 VDDA.n120 3390
R4593 VDDA.n21 VDDA.n14 3390
R4594 VDDA.n23 VDDA.n14 3390
R4595 VDDA.n21 VDDA.n20 3390
R4596 VDDA.n23 VDDA.n20 3390
R4597 VDDA.n305 VDDA.n299 3180
R4598 VDDA.n305 VDDA.n300 3180
R4599 VDDA.n303 VDDA.n299 3180
R4600 VDDA.n303 VDDA.n300 3180
R4601 VDDA.n266 VDDA.n260 3180
R4602 VDDA.n266 VDDA.n261 3180
R4603 VDDA.n264 VDDA.n260 3180
R4604 VDDA.n264 VDDA.n261 3180
R4605 VDDA.n230 VDDA.n221 3060
R4606 VDDA.n230 VDDA.n222 2970
R4607 VDDA.n163 VDDA.n157 2940
R4608 VDDA.n165 VDDA.n157 2940
R4609 VDDA.n165 VDDA.n162 2940
R4610 VDDA.n163 VDDA.n162 2940
R4611 VDDA.n171 VDDA.n152 2940
R4612 VDDA.n173 VDDA.n152 2940
R4613 VDDA.n173 VDDA.n170 2940
R4614 VDDA.n171 VDDA.n170 2940
R4615 VDDA.n232 VDDA.n221 2820
R4616 VDDA.n232 VDDA.n222 2730
R4617 VDDA.n363 VDDA.n358 2190
R4618 VDDA.n365 VDDA.n358 2190
R4619 VDDA.n363 VDDA.n361 2190
R4620 VDDA.n365 VDDA.n361 2190
R4621 VDDA.n335 VDDA.n330 1770
R4622 VDDA.n337 VDDA.n330 1770
R4623 VDDA.n335 VDDA.n333 1770
R4624 VDDA.n337 VDDA.n333 1770
R4625 VDDA.n135 VDDA.t151 1216.42
R4626 VDDA.n146 VDDA.t136 1216.42
R4627 VDDA.n39 VDDA.t148 1216.42
R4628 VDDA.n47 VDDA.t178 1216.42
R4629 VDDA.n347 VDDA.n346 704
R4630 VDDA.n347 VDDA.n313 704
R4631 VDDA.n159 VDDA.t132 689.4
R4632 VDDA.n158 VDDA.t144 689.4
R4633 VDDA.n154 VDDA.t216 689.4
R4634 VDDA.n153 VDDA.t117 689.4
R4635 VDDA.n218 VDDA.t201 675.274
R4636 VDDA.n219 VDDA.t220 675.274
R4637 VDDA.n202 VDDA.t198 663.801
R4638 VDDA.n212 VDDA.t192 663.801
R4639 VDDA.n97 VDDA.t205 660.109
R4640 VDDA.n95 VDDA.t124 660.109
R4641 VDDA.n73 VDDA.t106 660.109
R4642 VDDA.n71 VDDA.t184 660.109
R4643 VDDA.n223 VDDA.t120 634.25
R4644 VDDA.n238 VDDA.t177 634.25
R4645 VDDA.n216 VDDA.n215 632.933
R4646 VDDA.n225 VDDA.n224 632.933
R4647 VDDA.n241 VDDA.n240 631.227
R4648 VDDA.n179 VDDA.n178 626.534
R4649 VDDA.n185 VDDA.n184 626.534
R4650 VDDA.n187 VDDA.n186 626.534
R4651 VDDA.n189 VDDA.n188 626.534
R4652 VDDA.n191 VDDA.n190 626.534
R4653 VDDA.n193 VDDA.n192 626.534
R4654 VDDA.n195 VDDA.n194 626.534
R4655 VDDA.n197 VDDA.n196 626.534
R4656 VDDA.n199 VDDA.n198 626.534
R4657 VDDA.n201 VDDA.n200 626.534
R4658 VDDA.n117 VDDA.t139 573.75
R4659 VDDA.n115 VDDA.t121 573.75
R4660 VDDA.n17 VDDA.t160 573.75
R4661 VDDA.n15 VDDA.t181 573.75
R4662 VDDA.n352 VDDA.n351 518.4
R4663 VDDA.n351 VDDA.n343 518.4
R4664 VDDA.n414 VDDA.n413 496
R4665 VDDA.n414 VDDA.n402 496
R4666 VDDA.n140 VDDA.n112 491.2
R4667 VDDA.n140 VDDA.n139 491.2
R4668 VDDA.n45 VDDA.n27 491.2
R4669 VDDA.n41 VDDA.n27 491.2
R4670 VDDA.n205 VDDA.n181 489.601
R4671 VDDA.n209 VDDA.n181 489.601
R4672 VDDA.n285 VDDA.n274 464
R4673 VDDA.n281 VDDA.n274 464
R4674 VDDA.n105 VDDA.n104 428.8
R4675 VDDA.n105 VDDA.n93 428.8
R4676 VDDA.n81 VDDA.n80 428.8
R4677 VDDA.n81 VDDA.n69 428.8
R4678 VDDA.n328 VDDA.t109 413.084
R4679 VDDA.n331 VDDA.t133 413.084
R4680 VDDA.n287 VDDA.t114 403.051
R4681 VDDA.n279 VDDA.t165 403.051
R4682 VDDA.t209 VDDA.n363 394.774
R4683 VDDA.n365 VDDA.t128 394.774
R4684 VDDA.t200 VDDA.t176 392.065
R4685 VDDA.t197 VDDA.n206 389.375
R4686 VDDA.n208 VDDA.t191 389.375
R4687 VDDA.t215 VDDA.n170 389.375
R4688 VDDA.t116 VDDA.n152 389.375
R4689 VDDA.n356 VDDA.t210 389.185
R4690 VDDA.n359 VDDA.t129 389.185
R4691 VDDA.n204 VDDA.n180 387.2
R4692 VDDA.n210 VDDA.n180 387.2
R4693 VDDA.n328 VDDA.t111 384.918
R4694 VDDA.n331 VDDA.t135 384.918
R4695 VDDA.n383 VDDA.t156 384.918
R4696 VDDA.n385 VDDA.t195 384.918
R4697 VDDA.n406 VDDA.t159 384.918
R4698 VDDA.n404 VDDA.t147 384.918
R4699 VDDA.t131 VDDA.n162 384.168
R4700 VDDA.t143 VDDA.n157 384.168
R4701 VDDA.n431 VDDA.n384 384
R4702 VDDA.n431 VDDA.n430 384
R4703 VDDA.n408 VDDA.n407 384
R4704 VDDA.n408 VDDA.n405 384
R4705 VDDA.t164 VDDA.n282 369.584
R4706 VDDA.n284 VDDA.t113 369.584
R4707 VDDA.t119 VDDA.n230 363.93
R4708 VDDA.n232 VDDA.t218 363.93
R4709 VDDA.n342 VDDA.t166 360.868
R4710 VDDA.n353 VDDA.t172 360.868
R4711 VDDA.n383 VDDA.t154 358.858
R4712 VDDA.n385 VDDA.t193 358.858
R4713 VDDA.n406 VDDA.t157 358.858
R4714 VDDA.n404 VDDA.t145 358.858
R4715 VDDA.n272 VDDA.n271 355.272
R4716 VDDA.n278 VDDA.n277 355.272
R4717 VDDA.n289 VDDA.n288 355.272
R4718 VDDA.n291 VDDA.n290 355.272
R4719 VDDA.n125 VDDA.n124 355.2
R4720 VDDA.n125 VDDA.n113 355.2
R4721 VDDA.n25 VDDA.n24 355.2
R4722 VDDA.n25 VDDA.n13 355.2
R4723 VDDA.t155 VDDA.n381 351.591
R4724 VDDA.t194 VDDA.n382 351.591
R4725 VDDA.t158 VDDA.n410 351.591
R4726 VDDA.n412 VDDA.t146 351.591
R4727 VDDA.n294 VDDA.n293 350.772
R4728 VDDA.n280 VDDA.n273 345.601
R4729 VDDA.n286 VDDA.n273 345.601
R4730 VDDA.t110 VDDA.n335 344.394
R4731 VDDA.n337 VDDA.t134 344.394
R4732 VDDA.n397 VDDA.n395 342.301
R4733 VDDA.n425 VDDA.n424 341.676
R4734 VDDA.n423 VDDA.n422 341.676
R4735 VDDA.n421 VDDA.n420 341.676
R4736 VDDA.n419 VDDA.n418 341.676
R4737 VDDA.n401 VDDA.n400 341.676
R4738 VDDA.n399 VDDA.n398 341.676
R4739 VDDA.n397 VDDA.n396 341.676
R4740 VDDA.n302 VDDA.n301 339.2
R4741 VDDA.n302 VDDA.n250 339.2
R4742 VDDA.n263 VDDA.n262 339.2
R4743 VDDA.n263 VDDA.n255 339.2
R4744 VDDA.n393 VDDA.n392 337.176
R4745 VDDA.n390 VDDA.n388 337.176
R4746 VDDA.n379 VDDA.n378 337.176
R4747 VDDA.n436 VDDA.n377 337.176
R4748 VDDA.n439 VDDA.n438 337.176
R4749 VDDA.n443 VDDA.n442 337.176
R4750 VDDA.n446 VDDA.n445 337.176
R4751 VDDA.n449 VDDA.n373 337.176
R4752 VDDA.n427 VDDA.n387 337.176
R4753 VDDA.n416 VDDA.n415 337.176
R4754 VDDA.n297 VDDA.t211 336.767
R4755 VDDA.n308 VDDA.t202 336.767
R4756 VDDA.n258 VDDA.t169 336.767
R4757 VDDA.n269 VDDA.t187 336.767
R4758 VDDA.n369 VDDA.n355 335.022
R4759 VDDA.n227 VDDA.t118 334.759
R4760 VDDA.n237 VDDA.t175 334.759
R4761 VDDA.n203 VDDA.t196 332.75
R4762 VDDA.n211 VDDA.t190 332.75
R4763 VDDA.n159 VDDA.t130 332.75
R4764 VDDA.n158 VDDA.t142 332.75
R4765 VDDA.n154 VDDA.t214 332.75
R4766 VDDA.n153 VDDA.t115 332.75
R4767 VDDA.t118 VDDA.n226 326.726
R4768 VDDA.n229 VDDA.n220 326.401
R4769 VDDA.n218 VDDA.t199 314.274
R4770 VDDA.n219 VDDA.t217 314.274
R4771 VDDA.n161 VDDA.n156 313.601
R4772 VDDA.n168 VDDA.n156 307.2
R4773 VDDA.n176 VDDA.n151 307.2
R4774 VDDA.n169 VDDA.n151 307.2
R4775 VDDA.n233 VDDA.n220 300.8
R4776 VDDA.t140 VDDA.n121 285.815
R4777 VDDA.n123 VDDA.t122 285.815
R4778 VDDA.t161 VDDA.n21 285.815
R4779 VDDA.n23 VDDA.t182 285.815
R4780 VDDA.t173 VDDA.n344 278.95
R4781 VDDA.t167 VDDA.n345 278.95
R4782 VDDA.n117 VDDA.t141 277.916
R4783 VDDA.n115 VDDA.t123 277.916
R4784 VDDA.n17 VDDA.t162 277.916
R4785 VDDA.n15 VDDA.t183 277.916
R4786 VDDA.n145 VDDA.n112 276.8
R4787 VDDA.n139 VDDA.n136 276.8
R4788 VDDA.n46 VDDA.n45 276.8
R4789 VDDA.n41 VDDA.n40 276.8
R4790 VDDA.n356 VDDA.t208 274.509
R4791 VDDA.n359 VDDA.t127 274.509
R4792 VDDA.n353 VDDA.t174 270.705
R4793 VDDA.n342 VDDA.t168 270.705
R4794 VDDA.n279 VDDA.t163 264.668
R4795 VDDA.n287 VDDA.t112 264.668
R4796 VDDA.t394 VDDA.t209 259.091
R4797 VDDA.t128 VDDA.t332 259.091
R4798 VDDA.t206 VDDA.n101 239.915
R4799 VDDA.n103 VDDA.t125 239.915
R4800 VDDA.t107 VDDA.n77 239.915
R4801 VDDA.n79 VDDA.t185 239.915
R4802 VDDA.t334 VDDA.t164 237.5
R4803 VDDA.t318 VDDA.t334 237.5
R4804 VDDA.t345 VDDA.t318 237.5
R4805 VDDA.t347 VDDA.t345 237.5
R4806 VDDA.t316 VDDA.t347 237.5
R4807 VDDA.t76 VDDA.t104 237.5
R4808 VDDA.t349 VDDA.t76 237.5
R4809 VDDA.t392 VDDA.t349 237.5
R4810 VDDA.t74 VDDA.t392 237.5
R4811 VDDA.t113 VDDA.t74 237.5
R4812 VDDA.t203 VDDA.n299 234.242
R4813 VDDA.t212 VDDA.n300 234.242
R4814 VDDA.n366 VDDA.n360 233.601
R4815 VDDA.n362 VDDA.n360 233.601
R4816 VDDA.t188 VDDA.n260 232.1
R4817 VDDA.t170 VDDA.n261 232.1
R4818 VDDA.n99 VDDA.n98 230.4
R4819 VDDA.n99 VDDA.n96 230.4
R4820 VDDA.n75 VDDA.n74 230.4
R4821 VDDA.n75 VDDA.n72 230.4
R4822 VDDA.n166 VDDA.n160 211.201
R4823 VDDA.n167 VDDA.n166 211.201
R4824 VDDA.n175 VDDA.n174 211.201
R4825 VDDA.n119 VDDA.n118 211.201
R4826 VDDA.n119 VDDA.n116 211.201
R4827 VDDA.n19 VDDA.n18 211.201
R4828 VDDA.n19 VDDA.n16 211.201
R4829 VDDA.n228 VDDA.n217 208
R4830 VDDA.n145 VDDA.n144 204.8
R4831 VDDA.n144 VDDA.n136 204.8
R4832 VDDA.n40 VDDA.n26 204.8
R4833 VDDA.n46 VDDA.n26 204.8
R4834 VDDA.n174 VDDA.n155 202.971
R4835 VDDA.n104 VDDA.n96 198.4
R4836 VDDA.n98 VDDA.n93 198.4
R4837 VDDA.n80 VDDA.n72 198.4
R4838 VDDA.n74 VDDA.n69 198.4
R4839 VDDA.n338 VDDA.n332 188.8
R4840 VDDA.n334 VDDA.n332 188.8
R4841 VDDA.n429 VDDA.n428 188.8
R4842 VDDA.n448 VDDA.n374 188.8
R4843 VDDA.t322 VDDA.t197 186.607
R4844 VDDA.t324 VDDA.t322 186.607
R4845 VDDA.t19 VDDA.t324 186.607
R4846 VDDA.t7 VDDA.t19 186.607
R4847 VDDA.t245 VDDA.t7 186.607
R4848 VDDA.t43 VDDA.t245 186.607
R4849 VDDA.t239 VDDA.t43 186.607
R4850 VDDA.t1 VDDA.t239 186.607
R4851 VDDA.t378 VDDA.t1 186.607
R4852 VDDA.t320 VDDA.t378 186.607
R4853 VDDA.t3 VDDA.t5 186.607
R4854 VDDA.t47 VDDA.t3 186.607
R4855 VDDA.t243 VDDA.t47 186.607
R4856 VDDA.t326 VDDA.t243 186.607
R4857 VDDA.t237 VDDA.t326 186.607
R4858 VDDA.t45 VDDA.t237 186.607
R4859 VDDA.t376 VDDA.t45 186.607
R4860 VDDA.t21 VDDA.t376 186.607
R4861 VDDA.t49 VDDA.t21 186.607
R4862 VDDA.t191 VDDA.t49 186.607
R4863 VDDA.t235 VDDA.t215 186.607
R4864 VDDA.t344 VDDA.t235 186.607
R4865 VDDA.t31 VDDA.t344 186.607
R4866 VDDA.t55 VDDA.t31 186.607
R4867 VDDA.t78 VDDA.t55 186.607
R4868 VDDA.t452 VDDA.t232 186.607
R4869 VDDA.t232 VDDA.t391 186.607
R4870 VDDA.t391 VDDA.t236 186.607
R4871 VDDA.t236 VDDA.t389 186.607
R4872 VDDA.t389 VDDA.t116 186.607
R4873 VDDA.n308 VDDA.t204 183.661
R4874 VDDA.n297 VDDA.t213 183.661
R4875 VDDA.n269 VDDA.t189 183.661
R4876 VDDA.n258 VDDA.t171 183.661
R4877 VDDA.t390 VDDA.t131 183.333
R4878 VDDA.t286 VDDA.t390 183.333
R4879 VDDA.t13 VDDA.t286 183.333
R4880 VDDA.t233 VDDA.t13 183.333
R4881 VDDA.t61 VDDA.t233 183.333
R4882 VDDA.t67 VDDA.t63 183.333
R4883 VDDA.t63 VDDA.t234 183.333
R4884 VDDA.t234 VDDA.t56 183.333
R4885 VDDA.t56 VDDA.t448 183.333
R4886 VDDA.t448 VDDA.t143 183.333
R4887 VDDA.n346 VDDA.n343 182.4
R4888 VDDA.n352 VDDA.n313 182.4
R4889 VDDA.n249 VDDA.n248 181.701
R4890 VDDA.n252 VDDA.n251 181.701
R4891 VDDA.n254 VDDA.n253 181.701
R4892 VDDA.n257 VDDA.n256 181.701
R4893 VDDA.t249 VDDA.t119 180.952
R4894 VDDA.t473 VDDA.t249 180.952
R4895 VDDA.t385 VDDA.t473 180.952
R4896 VDDA.t98 VDDA.t385 180.952
R4897 VDDA.t17 VDDA.t200 180.952
R4898 VDDA.t218 VDDA.t17 180.952
R4899 VDDA.t340 VDDA.t203 178.125
R4900 VDDA.t336 VDDA.t340 178.125
R4901 VDDA.t83 VDDA.t102 178.125
R4902 VDDA.t102 VDDA.t212 178.125
R4903 VDDA.n134 VDDA.t153 178.124
R4904 VDDA.n147 VDDA.t138 178.124
R4905 VDDA.n38 VDDA.t150 178.124
R4906 VDDA.n48 VDDA.t180 178.124
R4907 VDDA.t342 VDDA.t188 176.29
R4908 VDDA.t338 VDDA.t342 176.29
R4909 VDDA.t85 VDDA.t351 176.29
R4910 VDDA.t351 VDDA.t170 176.29
R4911 VDDA.n307 VDDA.n306 172.8
R4912 VDDA.n306 VDDA.n298 172.8
R4913 VDDA.n268 VDDA.n267 172.8
R4914 VDDA.n267 VDDA.n259 172.8
R4915 VDDA.t432 VDDA.t155 172.727
R4916 VDDA.t412 VDDA.t432 172.727
R4917 VDDA.t408 VDDA.t412 172.727
R4918 VDDA.t428 VDDA.t408 172.727
R4919 VDDA.t426 VDDA.t428 172.727
R4920 VDDA.t440 VDDA.t426 172.727
R4921 VDDA.t436 VDDA.t440 172.727
R4922 VDDA.t424 VDDA.t436 172.727
R4923 VDDA.t418 VDDA.t424 172.727
R4924 VDDA.t410 VDDA.t406 172.727
R4925 VDDA.t406 VDDA.t438 172.727
R4926 VDDA.t438 VDDA.t434 172.727
R4927 VDDA.t434 VDDA.t422 172.727
R4928 VDDA.t422 VDDA.t416 172.727
R4929 VDDA.t416 VDDA.t420 172.727
R4930 VDDA.t420 VDDA.t414 172.727
R4931 VDDA.t414 VDDA.t430 172.727
R4932 VDDA.t430 VDDA.t194 172.727
R4933 VDDA.t400 VDDA.t158 172.727
R4934 VDDA.t247 VDDA.t400 172.727
R4935 VDDA.t359 VDDA.t247 172.727
R4936 VDDA.t41 VDDA.t359 172.727
R4937 VDDA.t453 VDDA.t41 172.727
R4938 VDDA.t221 VDDA.t453 172.727
R4939 VDDA.t370 VDDA.t221 172.727
R4940 VDDA.t93 VDDA.t370 172.727
R4941 VDDA.t34 VDDA.t93 172.727
R4942 VDDA.t368 VDDA.t307 172.727
R4943 VDDA.t398 VDDA.t368 172.727
R4944 VDDA.t396 VDDA.t398 172.727
R4945 VDDA.t361 VDDA.t396 172.727
R4946 VDDA.t36 VDDA.t361 172.727
R4947 VDDA.t457 VDDA.t36 172.727
R4948 VDDA.t444 VDDA.t457 172.727
R4949 VDDA.t446 VDDA.t444 172.727
R4950 VDDA.t146 VDDA.t446 172.727
R4951 VDDA.n312 VDDA.n311 168.435
R4952 VDDA.n315 VDDA.n314 168.435
R4953 VDDA.n317 VDDA.n316 168.435
R4954 VDDA.n319 VDDA.n318 168.435
R4955 VDDA.n321 VDDA.n320 168.435
R4956 VDDA.n323 VDDA.n322 168.435
R4957 VDDA.n325 VDDA.n324 168.435
R4958 VDDA.n327 VDDA.n326 168.435
R4959 VDDA.n301 VDDA.n298 166.4
R4960 VDDA.n307 VDDA.n250 166.4
R4961 VDDA.n262 VDDA.n259 166.4
R4962 VDDA.n268 VDDA.n255 166.4
R4963 VDDA.n231 VDDA.t98 165.874
R4964 VDDA.t137 VDDA.n137 161.817
R4965 VDDA.t152 VDDA.n138 161.817
R4966 VDDA.t149 VDDA.n42 161.817
R4967 VDDA.n44 VDDA.t179 161.817
R4968 VDDA.n91 VDDA.n89 160.428
R4969 VDDA.n88 VDDA.n86 160.428
R4970 VDDA.n67 VDDA.n65 160.428
R4971 VDDA.n64 VDDA.n62 160.428
R4972 VDDA.t263 VDDA.t173 159.814
R4973 VDDA.t26 VDDA.t263 159.814
R4974 VDDA.t471 VDDA.t26 159.814
R4975 VDDA.t455 VDDA.t471 159.814
R4976 VDDA.t461 VDDA.t455 159.814
R4977 VDDA.t230 VDDA.t461 159.814
R4978 VDDA.t259 VDDA.t230 159.814
R4979 VDDA.t313 VDDA.t259 159.814
R4980 VDDA.t310 VDDA.t466 159.814
R4981 VDDA.t466 VDDA.t261 159.814
R4982 VDDA.t261 VDDA.t449 159.814
R4983 VDDA.t449 VDDA.t464 159.814
R4984 VDDA.t464 VDDA.t257 159.814
R4985 VDDA.t257 VDDA.t469 159.814
R4986 VDDA.t469 VDDA.t459 159.814
R4987 VDDA.t459 VDDA.t167 159.814
R4988 VDDA.n91 VDDA.n90 159.803
R4989 VDDA.n88 VDDA.n87 159.803
R4990 VDDA.n67 VDDA.n66 159.803
R4991 VDDA.n64 VDDA.n63 159.803
R4992 VDDA.t82 VDDA.t110 158.333
R4993 VDDA.t134 VDDA.t64 158.333
R4994 VDDA.n97 VDDA.t207 155.125
R4995 VDDA.n95 VDDA.t126 155.125
R4996 VDDA.n73 VDDA.t108 155.125
R4997 VDDA.n71 VDDA.t186 155.125
R4998 VDDA.n134 VDDA.n133 151.882
R4999 VDDA.n38 VDDA.n37 151.882
R5000 VDDA.n148 VDDA.n147 151.321
R5001 VDDA.n49 VDDA.n48 151.321
R5002 VDDA.n124 VDDA.n116 150.4
R5003 VDDA.n118 VDDA.n113 150.4
R5004 VDDA.n24 VDDA.n16 150.4
R5005 VDDA.n18 VDDA.n13 150.4
R5006 VDDA.n107 VDDA.n106 146.002
R5007 VDDA.n83 VDDA.n82 146.002
R5008 VDDA.n111 VDDA.n110 145.429
R5009 VDDA.n127 VDDA.n126 145.429
R5010 VDDA.n129 VDDA.n128 145.429
R5011 VDDA.n131 VDDA.n130 145.429
R5012 VDDA.n133 VDDA.n132 145.429
R5013 VDDA.n12 VDDA.n11 145.429
R5014 VDDA.n31 VDDA.n30 145.429
R5015 VDDA.n33 VDDA.n32 145.429
R5016 VDDA.n35 VDDA.n34 145.429
R5017 VDDA.n37 VDDA.n36 145.429
R5018 VDDA.n147 VDDA.n146 135.387
R5019 VDDA.n135 VDDA.n134 135.387
R5020 VDDA.n48 VDDA.n47 135.387
R5021 VDDA.n39 VDDA.n38 135.387
R5022 VDDA.n286 VDDA.n285 134.4
R5023 VDDA.n281 VDDA.n280 134.4
R5024 VDDA.n364 VDDA.t394 129.546
R5025 VDDA.t332 VDDA.n364 129.546
R5026 VDDA.t255 VDDA.t140 121.513
R5027 VDDA.t364 VDDA.t255 121.513
R5028 VDDA.t10 VDDA.t364 121.513
R5029 VDDA.t95 VDDA.t10 121.513
R5030 VDDA.t62 VDDA.t95 121.513
R5031 VDDA.t374 VDDA.t365 121.513
R5032 VDDA.t251 VDDA.t374 121.513
R5033 VDDA.t254 VDDA.t251 121.513
R5034 VDDA.t353 VDDA.t254 121.513
R5035 VDDA.t122 VDDA.t353 121.513
R5036 VDDA.t270 VDDA.t161 121.513
R5037 VDDA.t281 VDDA.t270 121.513
R5038 VDDA.t282 VDDA.t281 121.513
R5039 VDDA.t227 VDDA.t282 121.513
R5040 VDDA.t66 VDDA.t227 121.513
R5041 VDDA.t224 VDDA.t267 121.513
R5042 VDDA.t266 VDDA.t224 121.513
R5043 VDDA.t223 VDDA.t266 121.513
R5044 VDDA.t290 VDDA.t223 121.513
R5045 VDDA.t182 VDDA.t290 121.513
R5046 VDDA.n283 VDDA.t316 118.751
R5047 VDDA.t104 VDDA.n283 118.751
R5048 VDDA.n367 VDDA.n366 118.4
R5049 VDDA.n362 VDDA.n357 118.4
R5050 VDDA.n339 VDDA.n338 118.4
R5051 VDDA.n334 VDDA.n329 118.4
R5052 VDDA.n430 VDDA.n429 118.4
R5053 VDDA.n384 VDDA.n374 118.4
R5054 VDDA.n413 VDDA.n405 118.4
R5055 VDDA.n407 VDDA.n402 118.4
R5056 VDDA.n235 VDDA.n234 115.201
R5057 VDDA.n229 VDDA.n228 108.8
R5058 VDDA.n234 VDDA.n233 108.8
R5059 VDDA.n368 VDDA.n367 107.52
R5060 VDDA.n368 VDDA.n357 107.52
R5061 VDDA.n205 VDDA.n204 102.4
R5062 VDDA.n210 VDDA.n209 102.4
R5063 VDDA.n161 VDDA.n160 102.4
R5064 VDDA.t68 VDDA.t206 98.2764
R5065 VDDA.t70 VDDA.t68 98.2764
R5066 VDDA.t32 VDDA.t70 98.2764
R5067 VDDA.t100 VDDA.t32 98.2764
R5068 VDDA.t387 VDDA.t100 98.2764
R5069 VDDA.t356 VDDA.t23 98.2764
R5070 VDDA.t79 VDDA.t356 98.2764
R5071 VDDA.t442 VDDA.t79 98.2764
R5072 VDDA.t383 VDDA.t442 98.2764
R5073 VDDA.t125 VDDA.t383 98.2764
R5074 VDDA.t90 VDDA.t107 98.2764
R5075 VDDA.t287 VDDA.t90 98.2764
R5076 VDDA.t228 VDDA.t287 98.2764
R5077 VDDA.t241 VDDA.t228 98.2764
R5078 VDDA.t11 VDDA.t241 98.2764
R5079 VDDA.t72 VDDA.t298 98.2764
R5080 VDDA.t303 VDDA.t72 98.2764
R5081 VDDA.t372 VDDA.t303 98.2764
R5082 VDDA.t87 VDDA.t372 98.2764
R5083 VDDA.t185 VDDA.t87 98.2764
R5084 VDDA.n52 VDDA.n50 97.4034
R5085 VDDA.n2 VDDA.n0 97.4034
R5086 VDDA.n60 VDDA.n59 96.8409
R5087 VDDA.n58 VDDA.n57 96.8409
R5088 VDDA.n56 VDDA.n55 96.8409
R5089 VDDA.n54 VDDA.n53 96.8409
R5090 VDDA.n52 VDDA.n51 96.8409
R5091 VDDA.n10 VDDA.n9 96.8409
R5092 VDDA.n8 VDDA.n7 96.8409
R5093 VDDA.n6 VDDA.n5 96.8409
R5094 VDDA.n4 VDDA.n3 96.8409
R5095 VDDA.n2 VDDA.n1 96.8409
R5096 VDDA.n168 VDDA.n167 96.0005
R5097 VDDA.n169 VDDA.n155 96.0005
R5098 VDDA.n176 VDDA.n175 96.0005
R5099 VDDA.n207 VDDA.t320 93.3041
R5100 VDDA.t5 VDDA.n207 93.3041
R5101 VDDA.n172 VDDA.t78 93.3041
R5102 VDDA.n172 VDDA.t452 93.3041
R5103 VDDA.n230 VDDA.n229 92.5005
R5104 VDDA.n221 VDDA.n220 92.5005
R5105 VDDA.n231 VDDA.n221 92.5005
R5106 VDDA.n233 VDDA.n232 92.5005
R5107 VDDA.n222 VDDA.n217 92.5005
R5108 VDDA.n231 VDDA.n222 92.5005
R5109 VDDA.n206 VDDA.n205 92.5005
R5110 VDDA.n182 VDDA.n181 92.5005
R5111 VDDA.n207 VDDA.n182 92.5005
R5112 VDDA.n209 VDDA.n208 92.5005
R5113 VDDA.n183 VDDA.n180 92.5005
R5114 VDDA.n207 VDDA.n183 92.5005
R5115 VDDA.n163 VDDA.n156 92.5005
R5116 VDDA.n164 VDDA.n163 92.5005
R5117 VDDA.n162 VDDA.n161 92.5005
R5118 VDDA.n166 VDDA.n165 92.5005
R5119 VDDA.n165 VDDA.n164 92.5005
R5120 VDDA.n168 VDDA.n157 92.5005
R5121 VDDA.n171 VDDA.n151 92.5005
R5122 VDDA.n172 VDDA.n171 92.5005
R5123 VDDA.n170 VDDA.n169 92.5005
R5124 VDDA.n174 VDDA.n173 92.5005
R5125 VDDA.n173 VDDA.n172 92.5005
R5126 VDDA.n176 VDDA.n152 92.5005
R5127 VDDA.n124 VDDA.n123 92.5005
R5128 VDDA.n120 VDDA.n119 92.5005
R5129 VDDA.n122 VDDA.n120 92.5005
R5130 VDDA.n121 VDDA.n113 92.5005
R5131 VDDA.n125 VDDA.n114 92.5005
R5132 VDDA.n122 VDDA.n114 92.5005
R5133 VDDA.n144 VDDA.n143 92.5005
R5134 VDDA.n143 VDDA.n142 92.5005
R5135 VDDA.n141 VDDA.n140 92.5005
R5136 VDDA.n142 VDDA.n141 92.5005
R5137 VDDA.n104 VDDA.n103 92.5005
R5138 VDDA.n100 VDDA.n99 92.5005
R5139 VDDA.n102 VDDA.n100 92.5005
R5140 VDDA.n101 VDDA.n93 92.5005
R5141 VDDA.n105 VDDA.n94 92.5005
R5142 VDDA.n102 VDDA.n94 92.5005
R5143 VDDA.n80 VDDA.n79 92.5005
R5144 VDDA.n76 VDDA.n75 92.5005
R5145 VDDA.n78 VDDA.n76 92.5005
R5146 VDDA.n77 VDDA.n69 92.5005
R5147 VDDA.n81 VDDA.n70 92.5005
R5148 VDDA.n78 VDDA.n70 92.5005
R5149 VDDA.n24 VDDA.n23 92.5005
R5150 VDDA.n20 VDDA.n19 92.5005
R5151 VDDA.n22 VDDA.n20 92.5005
R5152 VDDA.n21 VDDA.n13 92.5005
R5153 VDDA.n25 VDDA.n14 92.5005
R5154 VDDA.n22 VDDA.n14 92.5005
R5155 VDDA.n29 VDDA.n26 92.5005
R5156 VDDA.n43 VDDA.n29 92.5005
R5157 VDDA.n28 VDDA.n27 92.5005
R5158 VDDA.n43 VDDA.n28 92.5005
R5159 VDDA.n303 VDDA.n302 92.5005
R5160 VDDA.n304 VDDA.n303 92.5005
R5161 VDDA.n306 VDDA.n305 92.5005
R5162 VDDA.n305 VDDA.n304 92.5005
R5163 VDDA.n285 VDDA.n284 92.5005
R5164 VDDA.n276 VDDA.n274 92.5005
R5165 VDDA.n283 VDDA.n276 92.5005
R5166 VDDA.n282 VDDA.n281 92.5005
R5167 VDDA.n275 VDDA.n273 92.5005
R5168 VDDA.n283 VDDA.n275 92.5005
R5169 VDDA.n264 VDDA.n263 92.5005
R5170 VDDA.n265 VDDA.n264 92.5005
R5171 VDDA.n267 VDDA.n266 92.5005
R5172 VDDA.n266 VDDA.n265 92.5005
R5173 VDDA.n366 VDDA.n365 92.5005
R5174 VDDA.n363 VDDA.n362 92.5005
R5175 VDDA.n346 VDDA.n345 92.5005
R5176 VDDA.n348 VDDA.n347 92.5005
R5177 VDDA.n349 VDDA.n348 92.5005
R5178 VDDA.n344 VDDA.n313 92.5005
R5179 VDDA.n351 VDDA.n350 92.5005
R5180 VDDA.n350 VDDA.n349 92.5005
R5181 VDDA.n338 VDDA.n337 92.5005
R5182 VDDA.n333 VDDA.n332 92.5005
R5183 VDDA.n336 VDDA.n333 92.5005
R5184 VDDA.n335 VDDA.n334 92.5005
R5185 VDDA.n340 VDDA.n330 92.5005
R5186 VDDA.n336 VDDA.n330 92.5005
R5187 VDDA.n429 VDDA.n382 92.5005
R5188 VDDA.n432 VDDA.n431 92.5005
R5189 VDDA.n433 VDDA.n432 92.5005
R5190 VDDA.n381 VDDA.n374 92.5005
R5191 VDDA.n435 VDDA.n434 92.5005
R5192 VDDA.n434 VDDA.n433 92.5005
R5193 VDDA.n413 VDDA.n412 92.5005
R5194 VDDA.n409 VDDA.n408 92.5005
R5195 VDDA.n411 VDDA.n409 92.5005
R5196 VDDA.n410 VDDA.n402 92.5005
R5197 VDDA.n414 VDDA.n403 92.5005
R5198 VDDA.n411 VDDA.n403 92.5005
R5199 VDDA.n164 VDDA.t61 91.6672
R5200 VDDA.n164 VDDA.t67 91.6672
R5201 VDDA.n304 VDDA.t336 89.063
R5202 VDDA.n304 VDDA.t83 89.063
R5203 VDDA.n265 VDDA.t338 88.1448
R5204 VDDA.n265 VDDA.t85 88.1448
R5205 VDDA.n433 VDDA.t418 86.3641
R5206 VDDA.n433 VDDA.t410 86.3641
R5207 VDDA.n411 VDDA.t34 86.3641
R5208 VDDA.t307 VDDA.n411 86.3641
R5209 VDDA.n349 VDDA.t313 79.907
R5210 VDDA.n349 VDDA.t310 79.907
R5211 VDDA.n336 VDDA.t82 79.1672
R5212 VDDA.t64 VDDA.n336 79.1672
R5213 VDDA.n178 VDDA.t22 78.8005
R5214 VDDA.n178 VDDA.t50 78.8005
R5215 VDDA.n184 VDDA.t46 78.8005
R5216 VDDA.n184 VDDA.t377 78.8005
R5217 VDDA.n186 VDDA.t327 78.8005
R5218 VDDA.n186 VDDA.t238 78.8005
R5219 VDDA.n188 VDDA.t48 78.8005
R5220 VDDA.n188 VDDA.t244 78.8005
R5221 VDDA.n190 VDDA.t6 78.8005
R5222 VDDA.n190 VDDA.t4 78.8005
R5223 VDDA.n192 VDDA.t379 78.8005
R5224 VDDA.n192 VDDA.t321 78.8005
R5225 VDDA.n194 VDDA.t240 78.8005
R5226 VDDA.n194 VDDA.t2 78.8005
R5227 VDDA.n196 VDDA.t246 78.8005
R5228 VDDA.n196 VDDA.t44 78.8005
R5229 VDDA.n198 VDDA.t20 78.8005
R5230 VDDA.n198 VDDA.t8 78.8005
R5231 VDDA.n200 VDDA.t323 78.8005
R5232 VDDA.n200 VDDA.t325 78.8005
R5233 VDDA.n340 VDDA.n339 64.0005
R5234 VDDA.n340 VDDA.n329 64.0005
R5235 VDDA.n448 VDDA.n447 64.0005
R5236 VDDA.n447 VDDA.n444 64.0005
R5237 VDDA.n444 VDDA.n375 64.0005
R5238 VDDA.n435 VDDA.n375 64.0005
R5239 VDDA.n435 VDDA.n380 64.0005
R5240 VDDA.n389 VDDA.n380 64.0005
R5241 VDDA.n389 VDDA.n386 64.0005
R5242 VDDA.n428 VDDA.n386 64.0005
R5243 VDDA.t53 VDDA.t137 62.9523
R5244 VDDA.t38 VDDA.t53 62.9523
R5245 VDDA.t300 VDDA.t38 62.9523
R5246 VDDA.t96 VDDA.t300 62.9523
R5247 VDDA.t59 VDDA.t96 62.9523
R5248 VDDA.t366 VDDA.t380 62.9523
R5249 VDDA.t380 VDDA.t252 62.9523
R5250 VDDA.t252 VDDA.t51 62.9523
R5251 VDDA.t51 VDDA.t57 62.9523
R5252 VDDA.t57 VDDA.t152 62.9523
R5253 VDDA.t271 VDDA.t149 62.9523
R5254 VDDA.t225 VDDA.t271 62.9523
R5255 VDDA.t283 VDDA.t225 62.9523
R5256 VDDA.t291 VDDA.t283 62.9523
R5257 VDDA.t14 VDDA.t291 62.9523
R5258 VDDA.t296 VDDA.t278 62.9523
R5259 VDDA.t276 VDDA.t296 62.9523
R5260 VDDA.t294 VDDA.t276 62.9523
R5261 VDDA.t273 VDDA.t294 62.9523
R5262 VDDA.t179 VDDA.t273 62.9523
R5263 VDDA.n240 VDDA.t18 62.5402
R5264 VDDA.n240 VDDA.t219 62.5402
R5265 VDDA.n137 VDDA.n112 61.6672
R5266 VDDA.n139 VDDA.n138 61.6672
R5267 VDDA.n45 VDDA.n44 61.6672
R5268 VDDA.n42 VDDA.n41 61.6672
R5269 VDDA.n122 VDDA.t62 60.7563
R5270 VDDA.t365 VDDA.n122 60.7563
R5271 VDDA.n22 VDDA.t66 60.7563
R5272 VDDA.t267 VDDA.n22 60.7563
R5273 VDDA.n452 VDDA.t476 59.5681
R5274 VDDA.n453 VDDA.t477 59.5681
R5275 VDDA.n452 VDDA.t478 51.8887
R5276 VDDA.n215 VDDA.t386 49.2505
R5277 VDDA.n215 VDDA.t99 49.2505
R5278 VDDA.n224 VDDA.t250 49.2505
R5279 VDDA.n224 VDDA.t474 49.2505
R5280 VDDA.n102 VDDA.t387 49.1384
R5281 VDDA.t23 VDDA.n102 49.1384
R5282 VDDA.n78 VDDA.t11 49.1384
R5283 VDDA.t298 VDDA.n78 49.1384
R5284 VDDA.n454 VDDA.t475 48.9557
R5285 VDDA.n239 VDDA.n238 47.9338
R5286 VDDA.n361 VDDA.n360 46.2505
R5287 VDDA.n364 VDDA.n361 46.2505
R5288 VDDA.n368 VDDA.n358 46.2505
R5289 VDDA.n364 VDDA.n358 46.2505
R5290 VDDA.n236 VDDA.n235 44.8005
R5291 VDDA.n202 VDDA.n201 42.0963
R5292 VDDA.n213 VDDA.n212 41.5338
R5293 VDDA.n293 VDDA.t317 39.4005
R5294 VDDA.n293 VDDA.t105 39.4005
R5295 VDDA.n271 VDDA.t346 39.4005
R5296 VDDA.n271 VDDA.t348 39.4005
R5297 VDDA.n277 VDDA.t335 39.4005
R5298 VDDA.n277 VDDA.t319 39.4005
R5299 VDDA.n288 VDDA.t393 39.4005
R5300 VDDA.n288 VDDA.t75 39.4005
R5301 VDDA.n290 VDDA.t77 39.4005
R5302 VDDA.n290 VDDA.t350 39.4005
R5303 VDDA.n355 VDDA.t395 39.4005
R5304 VDDA.n355 VDDA.t333 39.4005
R5305 VDDA.n392 VDDA.t417 39.4005
R5306 VDDA.n392 VDDA.t421 39.4005
R5307 VDDA.n388 VDDA.t435 39.4005
R5308 VDDA.n388 VDDA.t423 39.4005
R5309 VDDA.n378 VDDA.t407 39.4005
R5310 VDDA.n378 VDDA.t439 39.4005
R5311 VDDA.n377 VDDA.t419 39.4005
R5312 VDDA.n377 VDDA.t411 39.4005
R5313 VDDA.n438 VDDA.t437 39.4005
R5314 VDDA.n438 VDDA.t425 39.4005
R5315 VDDA.n442 VDDA.t427 39.4005
R5316 VDDA.n442 VDDA.t441 39.4005
R5317 VDDA.n445 VDDA.t409 39.4005
R5318 VDDA.n445 VDDA.t429 39.4005
R5319 VDDA.n373 VDDA.t433 39.4005
R5320 VDDA.n373 VDDA.t413 39.4005
R5321 VDDA.n387 VDDA.t415 39.4005
R5322 VDDA.n387 VDDA.t431 39.4005
R5323 VDDA.n424 VDDA.t401 39.4005
R5324 VDDA.n424 VDDA.t248 39.4005
R5325 VDDA.n422 VDDA.t360 39.4005
R5326 VDDA.n422 VDDA.t42 39.4005
R5327 VDDA.n420 VDDA.t454 39.4005
R5328 VDDA.n420 VDDA.t222 39.4005
R5329 VDDA.n418 VDDA.t371 39.4005
R5330 VDDA.n418 VDDA.t94 39.4005
R5331 VDDA.n415 VDDA.t35 39.4005
R5332 VDDA.n415 VDDA.t308 39.4005
R5333 VDDA.n400 VDDA.t369 39.4005
R5334 VDDA.n400 VDDA.t399 39.4005
R5335 VDDA.n398 VDDA.t397 39.4005
R5336 VDDA.n398 VDDA.t362 39.4005
R5337 VDDA.n396 VDDA.t37 39.4005
R5338 VDDA.n396 VDDA.t458 39.4005
R5339 VDDA.n395 VDDA.t445 39.4005
R5340 VDDA.n395 VDDA.t447 39.4005
R5341 VDDA.n226 VDDA.n223 34.1338
R5342 VDDA.n238 VDDA.n237 32.0005
R5343 VDDA.n227 VDDA.n223 32.0005
R5344 VDDA.n142 VDDA.t59 31.4764
R5345 VDDA.n142 VDDA.t366 31.4764
R5346 VDDA.n43 VDDA.t14 31.4764
R5347 VDDA.t278 VDDA.n43 31.4764
R5348 VDDA.n169 VDDA.n168 28.663
R5349 VDDA.n456 VDDA.n455 28.3925
R5350 VDDA.n301 VDDA.n300 26.4291
R5351 VDDA.n299 VDDA.n250 26.4291
R5352 VDDA.n262 VDDA.n261 26.4291
R5353 VDDA.n260 VDDA.n255 26.4291
R5354 VDDA.n212 VDDA.n211 25.6005
R5355 VDDA.n203 VDDA.n202 25.6005
R5356 VDDA.n237 VDDA.n236 24.5338
R5357 VDDA.n235 VDDA.n218 24.5338
R5358 VDDA.n234 VDDA.n219 24.5338
R5359 VDDA.n228 VDDA.n227 24.5338
R5360 VDDA.n236 VDDA.n217 22.4005
R5361 VDDA VDDA.n242 22.2202
R5362 VDDA.n211 VDDA.n210 21.3338
R5363 VDDA.n204 VDDA.n203 21.3338
R5364 VDDA.n160 VDDA.n159 21.3338
R5365 VDDA.n167 VDDA.n158 21.3338
R5366 VDDA.n155 VDDA.n154 21.3338
R5367 VDDA.n175 VDDA.n153 21.3338
R5368 VDDA.n118 VDDA.n117 21.3338
R5369 VDDA.n116 VDDA.n115 21.3338
R5370 VDDA.n146 VDDA.n145 21.3338
R5371 VDDA.n136 VDDA.n135 21.3338
R5372 VDDA.n98 VDDA.n97 21.3338
R5373 VDDA.n96 VDDA.n95 21.3338
R5374 VDDA.n74 VDDA.n73 21.3338
R5375 VDDA.n72 VDDA.n71 21.3338
R5376 VDDA.n18 VDDA.n17 21.3338
R5377 VDDA.n16 VDDA.n15 21.3338
R5378 VDDA.n47 VDDA.n46 21.3338
R5379 VDDA.n40 VDDA.n39 21.3338
R5380 VDDA.n357 VDDA.n356 21.3338
R5381 VDDA.n367 VDDA.n359 21.3338
R5382 VDDA.n329 VDDA.n328 21.3338
R5383 VDDA.n339 VDDA.n331 21.3338
R5384 VDDA.n384 VDDA.n383 21.3338
R5385 VDDA.n430 VDDA.n385 21.3338
R5386 VDDA.n407 VDDA.n406 21.3338
R5387 VDDA.n405 VDDA.n404 21.3338
R5388 VDDA.n61 VDDA.n60 21.1567
R5389 VDDA.n177 VDDA.n176 19.5505
R5390 VDDA.n144 VDDA.n125 19.538
R5391 VDDA.n26 VDDA.n25 19.538
R5392 VDDA.n107 VDDA.n105 19.2005
R5393 VDDA.n83 VDDA.n81 19.2005
R5394 VDDA.n308 VDDA.n307 19.2005
R5395 VDDA.n298 VDDA.n297 19.2005
R5396 VDDA.n287 VDDA.n286 19.2005
R5397 VDDA.n280 VDDA.n279 19.2005
R5398 VDDA.n269 VDDA.n268 19.2005
R5399 VDDA.n259 VDDA.n258 19.2005
R5400 VDDA.n353 VDDA.n352 19.2005
R5401 VDDA.n343 VDDA.n342 19.2005
R5402 VDDA.n150 VDDA.n10 16.8443
R5403 VDDA.n341 VDDA.n340 16.363
R5404 VDDA.n248 VDDA.t341 15.7605
R5405 VDDA.n248 VDDA.t337 15.7605
R5406 VDDA.n251 VDDA.t84 15.7605
R5407 VDDA.n251 VDDA.t103 15.7605
R5408 VDDA.n253 VDDA.t343 15.7605
R5409 VDDA.n253 VDDA.t339 15.7605
R5410 VDDA.n256 VDDA.t86 15.7605
R5411 VDDA.n256 VDDA.t352 15.7605
R5412 VDDA.t176 VDDA.n231 15.0799
R5413 VDDA.n247 VDDA.t463 15.0181
R5414 VDDA.n289 VDDA.n287 14.8005
R5415 VDDA.n279 VDDA.n278 14.8005
R5416 VDDA.n258 VDDA.n257 14.8005
R5417 VDDA.n226 VDDA.n225 14.4255
R5418 VDDA.n297 VDDA.n296 13.8005
R5419 VDDA.n270 VDDA.n269 13.8005
R5420 VDDA.n309 VDDA.n308 13.8005
R5421 VDDA.n342 VDDA.n341 13.8005
R5422 VDDA.n354 VDDA.n353 13.8005
R5423 VDDA.n311 VDDA.t264 13.1338
R5424 VDDA.n311 VDDA.t27 13.1338
R5425 VDDA.n314 VDDA.t472 13.1338
R5426 VDDA.n314 VDDA.t456 13.1338
R5427 VDDA.n316 VDDA.t462 13.1338
R5428 VDDA.n316 VDDA.t231 13.1338
R5429 VDDA.n318 VDDA.t260 13.1338
R5430 VDDA.n318 VDDA.t314 13.1338
R5431 VDDA.n320 VDDA.t311 13.1338
R5432 VDDA.n320 VDDA.t467 13.1338
R5433 VDDA.n322 VDDA.t262 13.1338
R5434 VDDA.n322 VDDA.t450 13.1338
R5435 VDDA.n324 VDDA.t465 13.1338
R5436 VDDA.n324 VDDA.t258 13.1338
R5437 VDDA.n326 VDDA.t470 13.1338
R5438 VDDA.n326 VDDA.t460 13.1338
R5439 VDDA.n106 VDDA.t388 11.2576
R5440 VDDA.n106 VDDA.t24 11.2576
R5441 VDDA.n90 VDDA.t357 11.2576
R5442 VDDA.n90 VDDA.t80 11.2576
R5443 VDDA.n89 VDDA.t443 11.2576
R5444 VDDA.n89 VDDA.t384 11.2576
R5445 VDDA.n87 VDDA.t33 11.2576
R5446 VDDA.n87 VDDA.t101 11.2576
R5447 VDDA.n86 VDDA.t69 11.2576
R5448 VDDA.n86 VDDA.t71 11.2576
R5449 VDDA.n82 VDDA.t12 11.2576
R5450 VDDA.n82 VDDA.t299 11.2576
R5451 VDDA.n66 VDDA.t73 11.2576
R5452 VDDA.n66 VDDA.t304 11.2576
R5453 VDDA.n65 VDDA.t373 11.2576
R5454 VDDA.n65 VDDA.t88 11.2576
R5455 VDDA.n63 VDDA.t229 11.2576
R5456 VDDA.n63 VDDA.t242 11.2576
R5457 VDDA.n62 VDDA.t91 11.2576
R5458 VDDA.n62 VDDA.t288 11.2576
R5459 VDDA.n108 VDDA.n107 9.3005
R5460 VDDA.n84 VDDA.n83 9.3005
R5461 VDDA.n369 VDDA.n368 9.3005
R5462 VDDA.n449 VDDA.n448 9.3005
R5463 VDDA.n447 VDDA.n446 9.3005
R5464 VDDA.n444 VDDA.n443 9.3005
R5465 VDDA.n439 VDDA.n375 9.3005
R5466 VDDA.n436 VDDA.n435 9.3005
R5467 VDDA.n380 VDDA.n379 9.3005
R5468 VDDA.n390 VDDA.n389 9.3005
R5469 VDDA.n393 VDDA.n386 9.3005
R5470 VDDA.n428 VDDA.n427 9.3005
R5471 VDDA.n416 VDDA.n414 9.3005
R5472 VDDA.n455 VDDA.n454 8.03219
R5473 VDDA.n59 VDDA.t89 8.0005
R5474 VDDA.n59 VDDA.t405 8.0005
R5475 VDDA.n57 VDDA.t275 8.0005
R5476 VDDA.n57 VDDA.t269 8.0005
R5477 VDDA.n55 VDDA.t265 8.0005
R5478 VDDA.n55 VDDA.t280 8.0005
R5479 VDDA.n53 VDDA.t289 8.0005
R5480 VDDA.n53 VDDA.t268 8.0005
R5481 VDDA.n51 VDDA.t293 8.0005
R5482 VDDA.n51 VDDA.t16 8.0005
R5483 VDDA.n50 VDDA.t403 8.0005
R5484 VDDA.n50 VDDA.t65 8.0005
R5485 VDDA.n9 VDDA.t402 8.0005
R5486 VDDA.n9 VDDA.t305 8.0005
R5487 VDDA.n7 VDDA.t354 8.0005
R5488 VDDA.n7 VDDA.t306 8.0005
R5489 VDDA.n5 VDDA.t355 8.0005
R5490 VDDA.n5 VDDA.t382 8.0005
R5491 VDDA.n3 VDDA.t363 8.0005
R5492 VDDA.n3 VDDA.t9 8.0005
R5493 VDDA.n1 VDDA.t40 8.0005
R5494 VDDA.n1 VDDA.t302 8.0005
R5495 VDDA.n0 VDDA.t375 8.0005
R5496 VDDA.n0 VDDA.t404 8.0005
R5497 VDDA.n214 VDDA.n213 7.438
R5498 VDDA.n242 VDDA.n241 7.03175
R5499 VDDA.n110 VDDA.t54 6.56717
R5500 VDDA.n110 VDDA.t39 6.56717
R5501 VDDA.n126 VDDA.t301 6.56717
R5502 VDDA.n126 VDDA.t97 6.56717
R5503 VDDA.n128 VDDA.t60 6.56717
R5504 VDDA.n128 VDDA.t367 6.56717
R5505 VDDA.n130 VDDA.t381 6.56717
R5506 VDDA.n130 VDDA.t253 6.56717
R5507 VDDA.n132 VDDA.t52 6.56717
R5508 VDDA.n132 VDDA.t58 6.56717
R5509 VDDA.n11 VDDA.t295 6.56717
R5510 VDDA.n11 VDDA.t274 6.56717
R5511 VDDA.n30 VDDA.t297 6.56717
R5512 VDDA.n30 VDDA.t277 6.56717
R5513 VDDA.n32 VDDA.t15 6.56717
R5514 VDDA.n32 VDDA.t279 6.56717
R5515 VDDA.n34 VDDA.t284 6.56717
R5516 VDDA.n34 VDDA.t292 6.56717
R5517 VDDA.n36 VDDA.t272 6.56717
R5518 VDDA.n36 VDDA.t226 6.56717
R5519 VDDA.n109 VDDA.n85 6.313
R5520 VDDA.n451 VDDA.n450 6.098
R5521 VDDA.n371 VDDA.n370 5.69621
R5522 VDDA.n295 VDDA.n270 5.188
R5523 VDDA.n296 VDDA.n295 5.188
R5524 VDDA.n456 VDDA.n247 5.16125
R5525 VDDA.n310 VDDA.n309 5.1605
R5526 VDDA.n295 VDDA.n294 5.15675
R5527 VDDA.n109 VDDA.n108 5.063
R5528 VDDA.n85 VDDA.n84 5.063
R5529 VDDA.n370 VDDA.n369 4.50831
R5530 VDDA.n108 VDDA.n92 4.5005
R5531 VDDA.n84 VDDA.n68 4.5005
R5532 VDDA.n150 VDDA.n149 4.5005
R5533 VDDA.n294 VDDA.n292 4.5005
R5534 VDDA.n417 VDDA.n416 4.5005
R5535 VDDA.n427 VDDA.n426 4.5005
R5536 VDDA.n394 VDDA.n393 4.5005
R5537 VDDA.n391 VDDA.n390 4.5005
R5538 VDDA.n379 VDDA.n376 4.5005
R5539 VDDA.n437 VDDA.n436 4.5005
R5540 VDDA.n440 VDDA.n439 4.5005
R5541 VDDA.n443 VDDA.n441 4.5005
R5542 VDDA.n446 VDDA.n372 4.5005
R5543 VDDA.n450 VDDA.n449 4.5005
R5544 VDDA.n453 VDDA.n452 4.12334
R5545 VDDA.n85 VDDA.n61 3.688
R5546 VDDA.n149 VDDA.n109 3.5005
R5547 VDDA.n426 VDDA.n425 3.3755
R5548 VDDA.n454 VDDA.n453 2.93377
R5549 VDDA.n370 VDDA.n354 2.91121
R5550 VDDA.n214 VDDA.n177 2.813
R5551 VDDA.n242 VDDA.n214 2.563
R5552 VDDA.n177 VDDA.n150 1.46925
R5553 VDDA.n241 VDDA.n239 1.063
R5554 VDDA.n292 VDDA.n291 1.0005
R5555 VDDA.n291 VDDA.n289 1.0005
R5556 VDDA.n278 VDDA.n272 1.0005
R5557 VDDA.n292 VDDA.n272 1.0005
R5558 VDDA.n257 VDDA.n254 1.0005
R5559 VDDA.n270 VDDA.n254 1.0005
R5560 VDDA.n296 VDDA.n252 1.0005
R5561 VDDA.n252 VDDA.n249 1.0005
R5562 VDDA.n309 VDDA.n249 1.0005
R5563 VDDA.n341 VDDA.n327 1.0005
R5564 VDDA.n327 VDDA.n325 1.0005
R5565 VDDA.n325 VDDA.n323 1.0005
R5566 VDDA.n323 VDDA.n321 1.0005
R5567 VDDA.n321 VDDA.n319 1.0005
R5568 VDDA.n319 VDDA.n317 1.0005
R5569 VDDA.n317 VDDA.n315 1.0005
R5570 VDDA.n315 VDDA.n312 1.0005
R5571 VDDA.n354 VDDA.n312 1.0005
R5572 VDDA.n149 VDDA.n148 0.938
R5573 VDDA.n455 VDDA.n451 0.840625
R5574 VDDA.n61 VDDA.n49 0.7505
R5575 VDDA.n451 VDDA.n371 0.74075
R5576 VDDA.n371 VDDA.n310 0.723125
R5577 VDDA.n225 VDDA.n216 0.6255
R5578 VDDA.n239 VDDA.n216 0.6255
R5579 VDDA.n92 VDDA.n91 0.6255
R5580 VDDA.n92 VDDA.n88 0.6255
R5581 VDDA.n68 VDDA.n67 0.6255
R5582 VDDA.n68 VDDA.n64 0.6255
R5583 VDDA.n399 VDDA.n397 0.6255
R5584 VDDA.n401 VDDA.n399 0.6255
R5585 VDDA.n417 VDDA.n401 0.6255
R5586 VDDA.n419 VDDA.n417 0.6255
R5587 VDDA.n421 VDDA.n419 0.6255
R5588 VDDA.n423 VDDA.n421 0.6255
R5589 VDDA.n425 VDDA.n423 0.6255
R5590 VDDA.n426 VDDA.n394 0.6255
R5591 VDDA.n394 VDDA.n391 0.6255
R5592 VDDA.n391 VDDA.n376 0.6255
R5593 VDDA.n437 VDDA.n376 0.6255
R5594 VDDA.n440 VDDA.n437 0.6255
R5595 VDDA.n441 VDDA.n440 0.6255
R5596 VDDA.n441 VDDA.n372 0.6255
R5597 VDDA.n450 VDDA.n372 0.6255
R5598 VDDA.n201 VDDA.n199 0.563
R5599 VDDA.n199 VDDA.n197 0.563
R5600 VDDA.n197 VDDA.n195 0.563
R5601 VDDA.n195 VDDA.n193 0.563
R5602 VDDA.n193 VDDA.n191 0.563
R5603 VDDA.n191 VDDA.n189 0.563
R5604 VDDA.n189 VDDA.n187 0.563
R5605 VDDA.n187 VDDA.n185 0.563
R5606 VDDA.n185 VDDA.n179 0.563
R5607 VDDA.n213 VDDA.n179 0.563
R5608 VDDA.n133 VDDA.n131 0.563
R5609 VDDA.n131 VDDA.n129 0.563
R5610 VDDA.n129 VDDA.n127 0.563
R5611 VDDA.n127 VDDA.n111 0.563
R5612 VDDA.n148 VDDA.n111 0.563
R5613 VDDA.n54 VDDA.n52 0.563
R5614 VDDA.n56 VDDA.n54 0.563
R5615 VDDA.n58 VDDA.n56 0.563
R5616 VDDA.n60 VDDA.n58 0.563
R5617 VDDA.n37 VDDA.n35 0.563
R5618 VDDA.n35 VDDA.n33 0.563
R5619 VDDA.n33 VDDA.n31 0.563
R5620 VDDA.n31 VDDA.n12 0.563
R5621 VDDA.n49 VDDA.n12 0.563
R5622 VDDA.n4 VDDA.n2 0.563
R5623 VDDA.n6 VDDA.n4 0.563
R5624 VDDA.n8 VDDA.n6 0.563
R5625 VDDA.n10 VDDA.n8 0.563
R5626 VDDA.n310 VDDA.n247 0.253125
R5627 VDDA.t0 VDDA.t256 0.1603
R5628 VDDA.t330 VDDA.t468 0.1603
R5629 VDDA.t81 VDDA.t331 0.1603
R5630 VDDA.t329 VDDA.t328 0.1603
R5631 VDDA.t28 VDDA.t30 0.1603
R5632 VDDA.t309 VDDA.t92 0.1603
R5633 VDDA.t29 VDDA.t285 0.1603
R5634 VDDA.t315 VDDA.t312 0.1603
R5635 VDDA.n244 VDDA.t25 0.159278
R5636 VDDA.n245 VDDA.t451 0.159278
R5637 VDDA.n246 VDDA.t358 0.159278
R5638 VDDA.n246 VDDA.t0 0.1368
R5639 VDDA.n246 VDDA.t330 0.1368
R5640 VDDA.n245 VDDA.t81 0.1368
R5641 VDDA.n245 VDDA.t329 0.1368
R5642 VDDA.n244 VDDA.t28 0.1368
R5643 VDDA.n244 VDDA.t309 0.1368
R5644 VDDA.n243 VDDA.t29 0.1368
R5645 VDDA.n243 VDDA.t315 0.1368
R5646 VDDA VDDA.n456 0.024
R5647 VDDA.t25 VDDA.n243 0.00152174
R5648 VDDA.t451 VDDA.n244 0.00152174
R5649 VDDA.t358 VDDA.n245 0.00152174
R5650 VDDA.t463 VDDA.n246 0.00152174
R5651 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 114.719
R5652 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5653 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5654 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 114.156
R5655 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5656 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5657 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5658 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5659 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5660 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5661 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5662 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5663 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5664 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5665 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5666 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5667 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5668 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5669 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5670 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5671 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5672 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5673 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5674 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5675 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5676 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5677 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5678 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5679 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5680 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5681 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5682 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5683 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5684 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5685 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5686 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5687 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5688 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5689 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5690 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5691 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n8 0.563
R5692 VOUT-.n14 VOUT-.n6 145.989
R5693 VOUT-.n9 VOUT-.n7 145.989
R5694 VOUT-.n13 VOUT-.n12 145.427
R5695 VOUT-.n11 VOUT-.n10 145.427
R5696 VOUT-.n9 VOUT-.n8 145.427
R5697 VOUT-.n16 VOUT-.n15 140.927
R5698 VOUT-.n5 VOUT-.t7 113.192
R5699 VOUT-.n2 VOUT-.n0 95.7303
R5700 VOUT-.n4 VOUT-.n3 94.6053
R5701 VOUT-.n2 VOUT-.n1 94.6053
R5702 VOUT-.n100 VOUT-.n16 20.5943
R5703 VOUT-.n100 VOUT-.n99 11.7059
R5704 VOUT- VOUT-.n100 7.813
R5705 VOUT-.n15 VOUT-.t2 6.56717
R5706 VOUT-.n15 VOUT-.t14 6.56717
R5707 VOUT-.n12 VOUT-.t8 6.56717
R5708 VOUT-.n12 VOUT-.t6 6.56717
R5709 VOUT-.n10 VOUT-.t15 6.56717
R5710 VOUT-.n10 VOUT-.t16 6.56717
R5711 VOUT-.n8 VOUT-.t13 6.56717
R5712 VOUT-.n8 VOUT-.t3 6.56717
R5713 VOUT-.n7 VOUT-.t5 6.56717
R5714 VOUT-.n7 VOUT-.t10 6.56717
R5715 VOUT-.n6 VOUT-.t9 6.56717
R5716 VOUT-.n6 VOUT-.t4 6.56717
R5717 VOUT-.n46 VOUT-.t83 4.8295
R5718 VOUT-.n48 VOUT-.t90 4.8295
R5719 VOUT-.n51 VOUT-.t128 4.8295
R5720 VOUT-.n54 VOUT-.t26 4.8295
R5721 VOUT-.n57 VOUT-.t74 4.8295
R5722 VOUT-.n70 VOUT-.t39 4.8295
R5723 VOUT-.n72 VOUT-.t34 4.8295
R5724 VOUT-.n73 VOUT-.t136 4.8295
R5725 VOUT-.n75 VOUT-.t68 4.8295
R5726 VOUT-.n76 VOUT-.t36 4.8295
R5727 VOUT-.n78 VOUT-.t94 4.8295
R5728 VOUT-.n79 VOUT-.t64 4.8295
R5729 VOUT-.n81 VOUT-.t54 4.8295
R5730 VOUT-.n82 VOUT-.t29 4.8295
R5731 VOUT-.n84 VOUT-.t89 4.8295
R5732 VOUT-.n85 VOUT-.t57 4.8295
R5733 VOUT-.n87 VOUT-.t48 4.8295
R5734 VOUT-.n88 VOUT-.t20 4.8295
R5735 VOUT-.n90 VOUT-.t148 4.8295
R5736 VOUT-.n91 VOUT-.t121 4.8295
R5737 VOUT-.n93 VOUT-.t43 4.8295
R5738 VOUT-.n94 VOUT-.t152 4.8295
R5739 VOUT-.n17 VOUT-.t107 4.8295
R5740 VOUT-.n29 VOUT-.t28 4.8295
R5741 VOUT-.n31 VOUT-.t24 4.8295
R5742 VOUT-.n32 VOUT-.t129 4.8295
R5743 VOUT-.n34 VOUT-.t59 4.8295
R5744 VOUT-.n35 VOUT-.t32 4.8295
R5745 VOUT-.n37 VOUT-.t99 4.8295
R5746 VOUT-.n38 VOUT-.t69 4.8295
R5747 VOUT-.n40 VOUT-.t67 4.8295
R5748 VOUT-.n41 VOUT-.t35 4.8295
R5749 VOUT-.n43 VOUT-.t104 4.8295
R5750 VOUT-.n44 VOUT-.t76 4.8295
R5751 VOUT-.n96 VOUT-.t115 4.8295
R5752 VOUT-.n69 VOUT-.t132 4.806
R5753 VOUT-.n68 VOUT-.t114 4.806
R5754 VOUT-.n67 VOUT-.t146 4.806
R5755 VOUT-.n66 VOUT-.t45 4.806
R5756 VOUT-.n65 VOUT-.t85 4.806
R5757 VOUT-.n64 VOUT-.t63 4.806
R5758 VOUT-.n63 VOUT-.t101 4.806
R5759 VOUT-.n62 VOUT-.t134 4.806
R5760 VOUT-.n61 VOUT-.t119 4.806
R5761 VOUT-.n60 VOUT-.t155 4.806
R5762 VOUT-.n28 VOUT-.t47 4.806
R5763 VOUT-.n27 VOUT-.t91 4.806
R5764 VOUT-.n26 VOUT-.t41 4.806
R5765 VOUT-.n25 VOUT-.t130 4.806
R5766 VOUT-.n24 VOUT-.t82 4.806
R5767 VOUT-.n23 VOUT-.t124 4.806
R5768 VOUT-.n22 VOUT-.t72 4.806
R5769 VOUT-.n21 VOUT-.t23 4.806
R5770 VOUT-.n20 VOUT-.t62 4.806
R5771 VOUT-.n19 VOUT-.t150 4.806
R5772 VOUT-.n47 VOUT-.t95 4.5005
R5773 VOUT-.n46 VOUT-.t56 4.5005
R5774 VOUT-.n48 VOUT-.t131 4.5005
R5775 VOUT-.n49 VOUT-.t103 4.5005
R5776 VOUT-.n50 VOUT-.t71 4.5005
R5777 VOUT-.n51 VOUT-.t31 4.5005
R5778 VOUT-.n52 VOUT-.t138 4.5005
R5779 VOUT-.n53 VOUT-.t106 4.5005
R5780 VOUT-.n54 VOUT-.t60 4.5005
R5781 VOUT-.n55 VOUT-.t40 4.5005
R5782 VOUT-.n56 VOUT-.t143 4.5005
R5783 VOUT-.n57 VOUT-.t113 4.5005
R5784 VOUT-.n58 VOUT-.t21 4.5005
R5785 VOUT-.n59 VOUT-.t125 4.5005
R5786 VOUT-.n60 VOUT-.t118 4.5005
R5787 VOUT-.n61 VOUT-.t80 4.5005
R5788 VOUT-.n62 VOUT-.t96 4.5005
R5789 VOUT-.n63 VOUT-.t61 4.5005
R5790 VOUT-.n64 VOUT-.t27 4.5005
R5791 VOUT-.n65 VOUT-.t44 4.5005
R5792 VOUT-.n66 VOUT-.t144 4.5005
R5793 VOUT-.n67 VOUT-.t111 4.5005
R5794 VOUT-.n68 VOUT-.t75 4.5005
R5795 VOUT-.n69 VOUT-.t92 4.5005
R5796 VOUT-.n71 VOUT-.t55 4.5005
R5797 VOUT-.n70 VOUT-.t19 4.5005
R5798 VOUT-.n72 VOUT-.t51 4.5005
R5799 VOUT-.n74 VOUT-.t156 4.5005
R5800 VOUT-.n73 VOUT-.t120 4.5005
R5801 VOUT-.n75 VOUT-.t87 4.5005
R5802 VOUT-.n77 VOUT-.t49 4.5005
R5803 VOUT-.n76 VOUT-.t151 4.5005
R5804 VOUT-.n78 VOUT-.t42 4.5005
R5805 VOUT-.n80 VOUT-.t145 4.5005
R5806 VOUT-.n79 VOUT-.t117 4.5005
R5807 VOUT-.n81 VOUT-.t141 4.5005
R5808 VOUT-.n83 VOUT-.t110 4.5005
R5809 VOUT-.n82 VOUT-.t79 4.5005
R5810 VOUT-.n84 VOUT-.t38 4.5005
R5811 VOUT-.n86 VOUT-.t139 4.5005
R5812 VOUT-.n85 VOUT-.t108 4.5005
R5813 VOUT-.n87 VOUT-.t135 4.5005
R5814 VOUT-.n89 VOUT-.t102 4.5005
R5815 VOUT-.n88 VOUT-.t70 4.5005
R5816 VOUT-.n90 VOUT-.t98 4.5005
R5817 VOUT-.n92 VOUT-.t66 4.5005
R5818 VOUT-.n91 VOUT-.t33 4.5005
R5819 VOUT-.n93 VOUT-.t133 4.5005
R5820 VOUT-.n95 VOUT-.t97 4.5005
R5821 VOUT-.n94 VOUT-.t65 4.5005
R5822 VOUT-.n18 VOUT-.t100 4.5005
R5823 VOUT-.n17 VOUT-.t149 4.5005
R5824 VOUT-.n19 VOUT-.t86 4.5005
R5825 VOUT-.n20 VOUT-.t50 4.5005
R5826 VOUT-.n21 VOUT-.t137 4.5005
R5827 VOUT-.n22 VOUT-.t105 4.5005
R5828 VOUT-.n23 VOUT-.t73 4.5005
R5829 VOUT-.n24 VOUT-.t25 4.5005
R5830 VOUT-.n25 VOUT-.t127 4.5005
R5831 VOUT-.n26 VOUT-.t88 4.5005
R5832 VOUT-.n27 VOUT-.t53 4.5005
R5833 VOUT-.n28 VOUT-.t140 4.5005
R5834 VOUT-.n30 VOUT-.t109 4.5005
R5835 VOUT-.n29 VOUT-.t78 4.5005
R5836 VOUT-.n31 VOUT-.t112 4.5005
R5837 VOUT-.n33 VOUT-.t77 4.5005
R5838 VOUT-.n32 VOUT-.t37 4.5005
R5839 VOUT-.n34 VOUT-.t147 4.5005
R5840 VOUT-.n36 VOUT-.t116 4.5005
R5841 VOUT-.n35 VOUT-.t81 4.5005
R5842 VOUT-.n37 VOUT-.t46 4.5005
R5843 VOUT-.n39 VOUT-.t153 4.5005
R5844 VOUT-.n38 VOUT-.t122 4.5005
R5845 VOUT-.n40 VOUT-.t154 4.5005
R5846 VOUT-.n42 VOUT-.t123 4.5005
R5847 VOUT-.n41 VOUT-.t84 4.5005
R5848 VOUT-.n43 VOUT-.t52 4.5005
R5849 VOUT-.n45 VOUT-.t22 4.5005
R5850 VOUT-.n44 VOUT-.t126 4.5005
R5851 VOUT-.n99 VOUT-.t142 4.5005
R5852 VOUT-.n98 VOUT-.t93 4.5005
R5853 VOUT-.n97 VOUT-.t58 4.5005
R5854 VOUT-.n96 VOUT-.t30 4.5005
R5855 VOUT-.n16 VOUT-.n14 4.5005
R5856 VOUT-.n3 VOUT-.t12 3.42907
R5857 VOUT-.n3 VOUT-.t17 3.42907
R5858 VOUT-.n1 VOUT-.t1 3.42907
R5859 VOUT-.n1 VOUT-.t11 3.42907
R5860 VOUT-.n0 VOUT-.t18 3.42907
R5861 VOUT-.n0 VOUT-.t0 3.42907
R5862 VOUT- VOUT-.n5 2.84425
R5863 VOUT-.n5 VOUT-.n4 2.03175
R5864 VOUT-.n4 VOUT-.n2 1.1255
R5865 VOUT-.n11 VOUT-.n9 0.563
R5866 VOUT-.n13 VOUT-.n11 0.563
R5867 VOUT-.n14 VOUT-.n13 0.563
R5868 VOUT-.n47 VOUT-.n46 0.3295
R5869 VOUT-.n50 VOUT-.n49 0.3295
R5870 VOUT-.n49 VOUT-.n48 0.3295
R5871 VOUT-.n53 VOUT-.n52 0.3295
R5872 VOUT-.n52 VOUT-.n51 0.3295
R5873 VOUT-.n56 VOUT-.n55 0.3295
R5874 VOUT-.n55 VOUT-.n54 0.3295
R5875 VOUT-.n59 VOUT-.n58 0.3295
R5876 VOUT-.n58 VOUT-.n57 0.3295
R5877 VOUT-.n61 VOUT-.n60 0.3295
R5878 VOUT-.n62 VOUT-.n61 0.3295
R5879 VOUT-.n63 VOUT-.n62 0.3295
R5880 VOUT-.n64 VOUT-.n63 0.3295
R5881 VOUT-.n65 VOUT-.n64 0.3295
R5882 VOUT-.n66 VOUT-.n65 0.3295
R5883 VOUT-.n67 VOUT-.n66 0.3295
R5884 VOUT-.n68 VOUT-.n67 0.3295
R5885 VOUT-.n69 VOUT-.n68 0.3295
R5886 VOUT-.n71 VOUT-.n69 0.3295
R5887 VOUT-.n71 VOUT-.n70 0.3295
R5888 VOUT-.n74 VOUT-.n72 0.3295
R5889 VOUT-.n74 VOUT-.n73 0.3295
R5890 VOUT-.n77 VOUT-.n75 0.3295
R5891 VOUT-.n77 VOUT-.n76 0.3295
R5892 VOUT-.n80 VOUT-.n78 0.3295
R5893 VOUT-.n80 VOUT-.n79 0.3295
R5894 VOUT-.n83 VOUT-.n81 0.3295
R5895 VOUT-.n83 VOUT-.n82 0.3295
R5896 VOUT-.n86 VOUT-.n84 0.3295
R5897 VOUT-.n86 VOUT-.n85 0.3295
R5898 VOUT-.n89 VOUT-.n87 0.3295
R5899 VOUT-.n89 VOUT-.n88 0.3295
R5900 VOUT-.n92 VOUT-.n90 0.3295
R5901 VOUT-.n92 VOUT-.n91 0.3295
R5902 VOUT-.n95 VOUT-.n93 0.3295
R5903 VOUT-.n95 VOUT-.n94 0.3295
R5904 VOUT-.n18 VOUT-.n17 0.3295
R5905 VOUT-.n20 VOUT-.n19 0.3295
R5906 VOUT-.n21 VOUT-.n20 0.3295
R5907 VOUT-.n22 VOUT-.n21 0.3295
R5908 VOUT-.n23 VOUT-.n22 0.3295
R5909 VOUT-.n24 VOUT-.n23 0.3295
R5910 VOUT-.n25 VOUT-.n24 0.3295
R5911 VOUT-.n26 VOUT-.n25 0.3295
R5912 VOUT-.n27 VOUT-.n26 0.3295
R5913 VOUT-.n28 VOUT-.n27 0.3295
R5914 VOUT-.n30 VOUT-.n28 0.3295
R5915 VOUT-.n30 VOUT-.n29 0.3295
R5916 VOUT-.n33 VOUT-.n31 0.3295
R5917 VOUT-.n33 VOUT-.n32 0.3295
R5918 VOUT-.n36 VOUT-.n34 0.3295
R5919 VOUT-.n36 VOUT-.n35 0.3295
R5920 VOUT-.n39 VOUT-.n37 0.3295
R5921 VOUT-.n39 VOUT-.n38 0.3295
R5922 VOUT-.n42 VOUT-.n40 0.3295
R5923 VOUT-.n42 VOUT-.n41 0.3295
R5924 VOUT-.n45 VOUT-.n43 0.3295
R5925 VOUT-.n45 VOUT-.n44 0.3295
R5926 VOUT-.n99 VOUT-.n98 0.3295
R5927 VOUT-.n98 VOUT-.n97 0.3295
R5928 VOUT-.n97 VOUT-.n96 0.3295
R5929 VOUT-.n67 VOUT-.n50 0.306
R5930 VOUT-.n66 VOUT-.n53 0.306
R5931 VOUT-.n65 VOUT-.n56 0.306
R5932 VOUT-.n64 VOUT-.n59 0.306
R5933 VOUT-.n71 VOUT-.n47 0.2825
R5934 VOUT-.n74 VOUT-.n71 0.2825
R5935 VOUT-.n77 VOUT-.n74 0.2825
R5936 VOUT-.n80 VOUT-.n77 0.2825
R5937 VOUT-.n83 VOUT-.n80 0.2825
R5938 VOUT-.n86 VOUT-.n83 0.2825
R5939 VOUT-.n89 VOUT-.n86 0.2825
R5940 VOUT-.n92 VOUT-.n89 0.2825
R5941 VOUT-.n95 VOUT-.n92 0.2825
R5942 VOUT-.n30 VOUT-.n18 0.2825
R5943 VOUT-.n33 VOUT-.n30 0.2825
R5944 VOUT-.n36 VOUT-.n33 0.2825
R5945 VOUT-.n39 VOUT-.n36 0.2825
R5946 VOUT-.n42 VOUT-.n39 0.2825
R5947 VOUT-.n45 VOUT-.n42 0.2825
R5948 VOUT-.n97 VOUT-.n45 0.2825
R5949 VOUT-.n97 VOUT-.n95 0.2825
R5950 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.083
R5951 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1603
R5952 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1603
R5953 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R5954 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R5955 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R5956 two_stage_opamp_dummy_magic_0.cap_res_X.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R5957 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R5958 two_stage_opamp_dummy_magic_0.cap_res_X.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1603
R5959 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R5960 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.1603
R5961 two_stage_opamp_dummy_magic_0.cap_res_X.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1603
R5962 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1603
R5963 two_stage_opamp_dummy_magic_0.cap_res_X.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R5964 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1603
R5965 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R5966 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1603
R5967 two_stage_opamp_dummy_magic_0.cap_res_X.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1603
R5968 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R5969 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1603
R5970 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1603
R5971 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R5972 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R5973 two_stage_opamp_dummy_magic_0.cap_res_X.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R5974 two_stage_opamp_dummy_magic_0.cap_res_X.t3 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R5975 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R5976 two_stage_opamp_dummy_magic_0.cap_res_X.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R5977 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R5978 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R5979 two_stage_opamp_dummy_magic_0.cap_res_X.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1603
R5980 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1603
R5981 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R5982 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.1603
R5983 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R5984 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R5985 two_stage_opamp_dummy_magic_0.cap_res_X.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R5986 two_stage_opamp_dummy_magic_0.cap_res_X.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.1603
R5987 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.1603
R5988 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1603
R5989 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R5990 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R5991 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1603
R5992 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R5993 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.1603
R5994 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R5995 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1603
R5996 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R5997 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R5998 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1603
R5999 two_stage_opamp_dummy_magic_0.cap_res_X.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R6000 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R6001 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R6002 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R6003 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1603
R6004 two_stage_opamp_dummy_magic_0.cap_res_X.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R6005 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R6006 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R6007 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R6008 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.1603
R6009 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.159278
R6010 two_stage_opamp_dummy_magic_0.cap_res_X.t48 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R6011 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R6012 two_stage_opamp_dummy_magic_0.cap_res_X.t41 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R6013 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R6014 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R6015 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R6016 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R6017 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R6018 two_stage_opamp_dummy_magic_0.cap_res_X.t91 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R6019 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R6020 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.159278
R6021 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.159278
R6022 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.159278
R6023 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.159278
R6024 two_stage_opamp_dummy_magic_0.cap_res_X.t1 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.159278
R6025 two_stage_opamp_dummy_magic_0.cap_res_X.t102 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.159278
R6026 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.159278
R6027 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.159278
R6028 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.159278
R6029 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.159278
R6030 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.159278
R6031 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.159278
R6032 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.159278
R6033 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.159278
R6034 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.159278
R6035 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.159278
R6036 two_stage_opamp_dummy_magic_0.cap_res_X.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.137822
R6037 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1368
R6038 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.1368
R6039 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.1368
R6040 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1368
R6041 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.1368
R6042 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1368
R6043 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1368
R6044 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R6045 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R6046 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1368
R6047 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R6048 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1368
R6049 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R6050 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R6051 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1368
R6052 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1368
R6053 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R6054 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R6055 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.1368
R6056 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R6057 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R6058 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1368
R6059 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1368
R6060 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1368
R6061 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1368
R6062 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R6063 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1368
R6064 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1368
R6065 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1368
R6066 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R6067 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R6068 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.118
R6069 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.114322
R6070 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R6071 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R6072 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R6073 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.1133
R6074 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.1133
R6075 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.1133
R6076 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.1133
R6077 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.1133
R6078 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.1133
R6079 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R6080 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R6081 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R6082 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R6083 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R6084 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R6085 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R6086 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R6087 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R6088 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R6089 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.00152174
R6090 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.00152174
R6091 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.00152174
R6092 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.00152174
R6093 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R6094 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R6095 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.00152174
R6096 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.00152174
R6097 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R6098 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.00152174
R6099 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.00152174
R6100 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R6101 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.00152174
R6102 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R6103 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.00152174
R6104 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.00152174
R6105 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R6106 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R6107 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.00152174
R6108 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.00152174
R6109 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R6110 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R6111 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R6112 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.00152174
R6113 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R6114 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.00152174
R6115 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.00152174
R6116 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R6117 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R6118 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.00152174
R6119 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.00152174
R6120 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.00152174
R6121 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R6122 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R6123 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.00152174
R6124 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R6125 ref_volt_cur_gen_dummy_magic_0.cap_res2.t0 ref_volt_cur_gen_dummy_magic_0.cap_res2.t18 188.963
R6126 ref_volt_cur_gen_dummy_magic_0.cap_res2.t13 ref_volt_cur_gen_dummy_magic_0.cap_res2.t14 0.1603
R6127 ref_volt_cur_gen_dummy_magic_0.cap_res2.t2 ref_volt_cur_gen_dummy_magic_0.cap_res2.t7 0.1603
R6128 ref_volt_cur_gen_dummy_magic_0.cap_res2.t6 ref_volt_cur_gen_dummy_magic_0.cap_res2.t9 0.1603
R6129 ref_volt_cur_gen_dummy_magic_0.cap_res2.t17 ref_volt_cur_gen_dummy_magic_0.cap_res2.t1 0.1603
R6130 ref_volt_cur_gen_dummy_magic_0.cap_res2.t19 ref_volt_cur_gen_dummy_magic_0.cap_res2.t3 0.1603
R6131 ref_volt_cur_gen_dummy_magic_0.cap_res2.t11 ref_volt_cur_gen_dummy_magic_0.cap_res2.t16 0.1603
R6132 ref_volt_cur_gen_dummy_magic_0.cap_res2.t4 ref_volt_cur_gen_dummy_magic_0.cap_res2.t8 0.1603
R6133 ref_volt_cur_gen_dummy_magic_0.cap_res2.t15 ref_volt_cur_gen_dummy_magic_0.cap_res2.t20 0.1603
R6134 ref_volt_cur_gen_dummy_magic_0.cap_res2.n1 ref_volt_cur_gen_dummy_magic_0.cap_res2.t10 0.159278
R6135 ref_volt_cur_gen_dummy_magic_0.cap_res2.n2 ref_volt_cur_gen_dummy_magic_0.cap_res2.t5 0.159278
R6136 ref_volt_cur_gen_dummy_magic_0.cap_res2.n3 ref_volt_cur_gen_dummy_magic_0.cap_res2.t12 0.159278
R6137 ref_volt_cur_gen_dummy_magic_0.cap_res2.n3 ref_volt_cur_gen_dummy_magic_0.cap_res2.t13 0.1368
R6138 ref_volt_cur_gen_dummy_magic_0.cap_res2.n3 ref_volt_cur_gen_dummy_magic_0.cap_res2.t2 0.1368
R6139 ref_volt_cur_gen_dummy_magic_0.cap_res2.n2 ref_volt_cur_gen_dummy_magic_0.cap_res2.t6 0.1368
R6140 ref_volt_cur_gen_dummy_magic_0.cap_res2.n2 ref_volt_cur_gen_dummy_magic_0.cap_res2.t17 0.1368
R6141 ref_volt_cur_gen_dummy_magic_0.cap_res2.n1 ref_volt_cur_gen_dummy_magic_0.cap_res2.t19 0.1368
R6142 ref_volt_cur_gen_dummy_magic_0.cap_res2.n1 ref_volt_cur_gen_dummy_magic_0.cap_res2.t11 0.1368
R6143 ref_volt_cur_gen_dummy_magic_0.cap_res2.n0 ref_volt_cur_gen_dummy_magic_0.cap_res2.t4 0.1368
R6144 ref_volt_cur_gen_dummy_magic_0.cap_res2.n0 ref_volt_cur_gen_dummy_magic_0.cap_res2.t15 0.1368
R6145 ref_volt_cur_gen_dummy_magic_0.cap_res2.t10 ref_volt_cur_gen_dummy_magic_0.cap_res2.n0 0.00152174
R6146 ref_volt_cur_gen_dummy_magic_0.cap_res2.t5 ref_volt_cur_gen_dummy_magic_0.cap_res2.n1 0.00152174
R6147 ref_volt_cur_gen_dummy_magic_0.cap_res2.t12 ref_volt_cur_gen_dummy_magic_0.cap_res2.n2 0.00152174
R6148 ref_volt_cur_gen_dummy_magic_0.cap_res2.t18 ref_volt_cur_gen_dummy_magic_0.cap_res2.n3 0.00152174
R6149 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n5 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t11 345.433
R6150 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n4 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t15 345.433
R6151 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n2 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t26 345.433
R6152 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n1 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t14 345.433
R6153 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n23 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n21 341.397
R6154 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n25 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n24 339.272
R6155 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n23 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n22 339.272
R6156 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n28 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n27 334.772
R6157 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n8 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t21 273.134
R6158 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n11 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t28 273.134
R6159 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n9 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n8 224.934
R6160 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n10 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n9 224.934
R6161 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n16 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n15 224.934
R6162 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n12 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n11 224.934
R6163 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n13 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n12 224.934
R6164 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n18 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n17 217.919
R6165 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n14 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n7 217.919
R6166 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t3 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n29 194.895
R6167 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n7 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n6 172.363
R6168 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n20 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n0 169.832
R6169 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n19 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n3 168.863
R6170 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n5 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t23 120.501
R6171 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n4 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t19 120.501
R6172 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n2 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t22 120.501
R6173 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n1 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t18 120.501
R6174 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n0 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t20 117.823
R6175 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n0 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t17 117.823
R6176 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n26 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t2 100.635
R6177 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n6 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n5 69.6227
R6178 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n6 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n4 69.6227
R6179 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n3 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n2 69.6227
R6180 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n3 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n1 69.6227
R6181 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n8 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t25 48.2005
R6182 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n9 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t12 48.2005
R6183 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n10 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t13 48.2005
R6184 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n17 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n10 48.2005
R6185 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n16 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t24 48.2005
R6186 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n17 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n16 48.2005
R6187 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n15 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t27 48.2005
R6188 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n11 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t16 48.2005
R6189 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n12 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t10 48.2005
R6190 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n13 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t29 48.2005
R6191 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n14 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n13 48.2005
R6192 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n15 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n14 48.2005
R6193 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n27 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t4 39.4005
R6194 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n27 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t1 39.4005
R6195 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n24 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t8 39.4005
R6196 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n24 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t6 39.4005
R6197 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n22 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t9 39.4005
R6198 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n22 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t7 39.4005
R6199 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n21 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t0 39.4005
R6200 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n21 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t5 39.4005
R6201 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n20 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n19 26.938
R6202 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n29 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n28 5.15675
R6203 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n28 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n26 4.5005
R6204 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n29 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n20 4.188
R6205 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n19 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n18 3.3755
R6206 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n25 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n23 2.1255
R6207 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n26 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n25 2.1255
R6208 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n18 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n7 1.0005
R6209 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 610.534
R6210 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 610.534
R6211 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R6212 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R6213 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R6214 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R6215 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R6216 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R6217 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R6218 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R6219 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R6220 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R6221 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 433.8
R6222 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R6223 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R6224 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R6225 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R6226 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R6227 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R6228 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 433.8
R6229 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 340.272
R6230 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 339.272
R6231 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R6232 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 334.772
R6233 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 221.293
R6234 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 176.733
R6235 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 176.733
R6236 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R6237 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R6238 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R6239 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R6240 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R6241 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R6242 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R6243 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 176.733
R6244 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R6245 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R6246 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R6247 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R6248 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R6249 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R6250 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 118.45
R6251 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 76.5943
R6252 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 64.5799
R6253 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 56.2338
R6254 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 56.2338
R6255 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 53.2453
R6256 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R6257 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R6258 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R6259 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R6260 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R6261 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 39.4005
R6262 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R6263 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R6264 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R6265 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R6266 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R6267 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 16.0005
R6268 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 5.5005
R6269 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 1.0005
R6270 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t27 355.293
R6271 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t20 346.8
R6272 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n10 339.522
R6273 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n8 339.522
R6274 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n12 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n4 335.022
R6275 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t0 275.909
R6276 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n6 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n5 227.909
R6277 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n4 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n7 222.034
R6278 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n11 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t30 184.097
R6279 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n11 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t26 184.097
R6280 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n9 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t29 184.097
R6281 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n9 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t24 184.097
R6282 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n11 166.05
R6283 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n9 166.05
R6284 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n7 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t7 48.0005
R6285 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n7 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t6 48.0005
R6286 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n5 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t3 48.0005
R6287 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n5 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t4 48.0005
R6288 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n10 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t10 39.4005
R6289 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n10 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t2 39.4005
R6290 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n8 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t8 39.4005
R6291 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n8 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t9 39.4005
R6292 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n12 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t5 39.4005
R6293 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n12 39.4005
R6294 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n0 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 32.0499
R6295 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n4 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n1 5.28175
R6296 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n1 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n0 5.188
R6297 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t36 4.8295
R6298 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t15 4.8295
R6299 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t17 4.8295
R6300 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t21 4.8295
R6301 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t35 4.8295
R6302 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t13 4.8295
R6303 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t31 4.8295
R6304 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t18 4.5005
R6305 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t12 4.5005
R6306 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t33 4.5005
R6307 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t22 4.5005
R6308 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t19 4.5005
R6309 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t14 4.5005
R6310 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t16 4.5005
R6311 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t11 4.5005
R6312 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t32 4.5005
R6313 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t25 4.5005
R6314 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t34 4.5005
R6315 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t28 4.5005
R6316 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t23 4.5005
R6317 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n4 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n6 4.5005
R6318 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 3.8075
R6319 ref_volt_cur_gen_dummy_magic_0.cap_res1.t20 ref_volt_cur_gen_dummy_magic_0.cap_res1.t6 179.073
R6320 ref_volt_cur_gen_dummy_magic_0.cap_res1.t8 ref_volt_cur_gen_dummy_magic_0.cap_res1.t5 0.1603
R6321 ref_volt_cur_gen_dummy_magic_0.cap_res1.t2 ref_volt_cur_gen_dummy_magic_0.cap_res1.t7 0.1603
R6322 ref_volt_cur_gen_dummy_magic_0.cap_res1.t4 ref_volt_cur_gen_dummy_magic_0.cap_res1.t17 0.1603
R6323 ref_volt_cur_gen_dummy_magic_0.cap_res1.t14 ref_volt_cur_gen_dummy_magic_0.cap_res1.t1 0.1603
R6324 ref_volt_cur_gen_dummy_magic_0.cap_res1.t16 ref_volt_cur_gen_dummy_magic_0.cap_res1.t10 0.1603
R6325 ref_volt_cur_gen_dummy_magic_0.cap_res1.t9 ref_volt_cur_gen_dummy_magic_0.cap_res1.t13 0.1603
R6326 ref_volt_cur_gen_dummy_magic_0.cap_res1.t3 ref_volt_cur_gen_dummy_magic_0.cap_res1.t15 0.1603
R6327 ref_volt_cur_gen_dummy_magic_0.cap_res1.t12 ref_volt_cur_gen_dummy_magic_0.cap_res1.t0 0.1603
R6328 ref_volt_cur_gen_dummy_magic_0.cap_res1.n1 ref_volt_cur_gen_dummy_magic_0.cap_res1.t18 0.159278
R6329 ref_volt_cur_gen_dummy_magic_0.cap_res1.n2 ref_volt_cur_gen_dummy_magic_0.cap_res1.t11 0.159278
R6330 ref_volt_cur_gen_dummy_magic_0.cap_res1.n3 ref_volt_cur_gen_dummy_magic_0.cap_res1.t19 0.159278
R6331 ref_volt_cur_gen_dummy_magic_0.cap_res1.n3 ref_volt_cur_gen_dummy_magic_0.cap_res1.t8 0.1368
R6332 ref_volt_cur_gen_dummy_magic_0.cap_res1.n3 ref_volt_cur_gen_dummy_magic_0.cap_res1.t2 0.1368
R6333 ref_volt_cur_gen_dummy_magic_0.cap_res1.n2 ref_volt_cur_gen_dummy_magic_0.cap_res1.t4 0.1368
R6334 ref_volt_cur_gen_dummy_magic_0.cap_res1.n2 ref_volt_cur_gen_dummy_magic_0.cap_res1.t14 0.1368
R6335 ref_volt_cur_gen_dummy_magic_0.cap_res1.n1 ref_volt_cur_gen_dummy_magic_0.cap_res1.t16 0.1368
R6336 ref_volt_cur_gen_dummy_magic_0.cap_res1.n1 ref_volt_cur_gen_dummy_magic_0.cap_res1.t9 0.1368
R6337 ref_volt_cur_gen_dummy_magic_0.cap_res1.n0 ref_volt_cur_gen_dummy_magic_0.cap_res1.t3 0.1368
R6338 ref_volt_cur_gen_dummy_magic_0.cap_res1.n0 ref_volt_cur_gen_dummy_magic_0.cap_res1.t12 0.1368
R6339 ref_volt_cur_gen_dummy_magic_0.cap_res1.t18 ref_volt_cur_gen_dummy_magic_0.cap_res1.n0 0.00152174
R6340 ref_volt_cur_gen_dummy_magic_0.cap_res1.t11 ref_volt_cur_gen_dummy_magic_0.cap_res1.n1 0.00152174
R6341 ref_volt_cur_gen_dummy_magic_0.cap_res1.t19 ref_volt_cur_gen_dummy_magic_0.cap_res1.n2 0.00152174
R6342 ref_volt_cur_gen_dummy_magic_0.cap_res1.t6 ref_volt_cur_gen_dummy_magic_0.cap_res1.n3 0.00152174
R6343 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 688.859
R6344 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 514.134
R6345 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 323.491
R6346 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 322.692
R6347 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6348 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6349 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 270.591
R6350 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 270.591
R6351 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 233.374
R6352 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 233.374
R6353 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 233.374
R6354 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 233.374
R6355 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 208.838
R6356 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 197.964
R6357 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 174.726
R6358 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6359 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 174.726
R6360 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 174.726
R6361 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 169.215
R6362 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 169.215
R6363 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 169.215
R6364 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 129.24
R6365 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 129.24
R6366 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6367 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6368 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 128.534
R6369 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 128.534
R6370 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 16.8443
R6371 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6372 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 13.1338
R6373 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6374 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6375 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6376 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6377 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 4.3755
R6378 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 4.3755
R6379 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 3.688
R6380 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 3.2505
R6381 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 3.1255
R6382 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 1.2755
R6383 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 1.2755
R6384 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 0.8005
R6385 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 632.186
R6386 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 630.264
R6387 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6388 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6389 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 628.003
R6390 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 628.003
R6391 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 626.753
R6392 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 626.753
R6393 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 625.756
R6394 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 622.231
R6395 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6396 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6397 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6398 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6399 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6400 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6401 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6402 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6403 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6404 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6405 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6406 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6407 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6408 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6409 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6410 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6411 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6412 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6413 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6414 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6415 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 7.94147
R6416 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 6.188
R6417 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 630.857
R6418 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 626.784
R6419 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n28 626.784
R6420 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n29 626.784
R6421 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n5 626.784
R6422 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.n25 585
R6423 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6424 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6425 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 176.733
R6426 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6427 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6428 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6429 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6430 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6431 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6432 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6433 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6434 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6435 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6436 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6437 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6438 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6439 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6440 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.n20 176.733
R6441 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n24 162.214
R6442 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n3 136.702
R6443 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6444 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6445 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6446 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6447 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6448 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6449 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6450 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6451 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6452 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6453 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6454 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6455 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6456 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6457 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6458 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6459 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6460 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6461 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6462 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6463 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6464 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R6465 two_stage_opamp_dummy_magic_0.V_err_gate.n29 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R6466 two_stage_opamp_dummy_magic_0.V_err_gate.n29 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6467 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R6468 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6469 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6470 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6471 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6472 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6473 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n2 67.6186
R6474 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n23 49.8072
R6475 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n21 49.8072
R6476 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 41.7838
R6477 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6478 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t4 24.0005
R6479 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t13 24.0005
R6480 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 1.1255
R6481 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n1 1.11856
R6482 ref_volt_cur_gen_dummy_magic_0.V_mir1.n20 ref_volt_cur_gen_dummy_magic_0.V_mir1.n19 325.473
R6483 ref_volt_cur_gen_dummy_magic_0.V_mir1.n9 ref_volt_cur_gen_dummy_magic_0.V_mir1.n5 325.471
R6484 ref_volt_cur_gen_dummy_magic_0.V_mir1.n4 ref_volt_cur_gen_dummy_magic_0.V_mir1.n0 325.471
R6485 ref_volt_cur_gen_dummy_magic_0.V_mir1.n16 ref_volt_cur_gen_dummy_magic_0.V_mir1.t19 310.488
R6486 ref_volt_cur_gen_dummy_magic_0.V_mir1.n6 ref_volt_cur_gen_dummy_magic_0.V_mir1.t22 310.488
R6487 ref_volt_cur_gen_dummy_magic_0.V_mir1.n1 ref_volt_cur_gen_dummy_magic_0.V_mir1.t17 310.488
R6488 ref_volt_cur_gen_dummy_magic_0.V_mir1.n12 ref_volt_cur_gen_dummy_magic_0.V_mir1.t3 278.312
R6489 ref_volt_cur_gen_dummy_magic_0.V_mir1.n12 ref_volt_cur_gen_dummy_magic_0.V_mir1.n11 228.939
R6490 ref_volt_cur_gen_dummy_magic_0.V_mir1.n13 ref_volt_cur_gen_dummy_magic_0.V_mir1.n10 224.439
R6491 ref_volt_cur_gen_dummy_magic_0.V_mir1.n18 ref_volt_cur_gen_dummy_magic_0.V_mir1.t12 184.097
R6492 ref_volt_cur_gen_dummy_magic_0.V_mir1.n8 ref_volt_cur_gen_dummy_magic_0.V_mir1.t4 184.097
R6493 ref_volt_cur_gen_dummy_magic_0.V_mir1.n3 ref_volt_cur_gen_dummy_magic_0.V_mir1.t6 184.097
R6494 ref_volt_cur_gen_dummy_magic_0.V_mir1.n17 ref_volt_cur_gen_dummy_magic_0.V_mir1.n16 167.094
R6495 ref_volt_cur_gen_dummy_magic_0.V_mir1.n7 ref_volt_cur_gen_dummy_magic_0.V_mir1.n6 167.094
R6496 ref_volt_cur_gen_dummy_magic_0.V_mir1.n2 ref_volt_cur_gen_dummy_magic_0.V_mir1.n1 167.094
R6497 ref_volt_cur_gen_dummy_magic_0.V_mir1.n9 ref_volt_cur_gen_dummy_magic_0.V_mir1.n8 152
R6498 ref_volt_cur_gen_dummy_magic_0.V_mir1.n4 ref_volt_cur_gen_dummy_magic_0.V_mir1.n3 152
R6499 ref_volt_cur_gen_dummy_magic_0.V_mir1.n19 ref_volt_cur_gen_dummy_magic_0.V_mir1.n18 152
R6500 ref_volt_cur_gen_dummy_magic_0.V_mir1.n16 ref_volt_cur_gen_dummy_magic_0.V_mir1.t21 120.501
R6501 ref_volt_cur_gen_dummy_magic_0.V_mir1.n17 ref_volt_cur_gen_dummy_magic_0.V_mir1.t14 120.501
R6502 ref_volt_cur_gen_dummy_magic_0.V_mir1.n6 ref_volt_cur_gen_dummy_magic_0.V_mir1.t20 120.501
R6503 ref_volt_cur_gen_dummy_magic_0.V_mir1.n7 ref_volt_cur_gen_dummy_magic_0.V_mir1.t8 120.501
R6504 ref_volt_cur_gen_dummy_magic_0.V_mir1.n1 ref_volt_cur_gen_dummy_magic_0.V_mir1.t18 120.501
R6505 ref_volt_cur_gen_dummy_magic_0.V_mir1.n2 ref_volt_cur_gen_dummy_magic_0.V_mir1.t10 120.501
R6506 ref_volt_cur_gen_dummy_magic_0.V_mir1.n11 ref_volt_cur_gen_dummy_magic_0.V_mir1.t1 48.0005
R6507 ref_volt_cur_gen_dummy_magic_0.V_mir1.n11 ref_volt_cur_gen_dummy_magic_0.V_mir1.t2 48.0005
R6508 ref_volt_cur_gen_dummy_magic_0.V_mir1.n10 ref_volt_cur_gen_dummy_magic_0.V_mir1.t16 48.0005
R6509 ref_volt_cur_gen_dummy_magic_0.V_mir1.n10 ref_volt_cur_gen_dummy_magic_0.V_mir1.t0 48.0005
R6510 ref_volt_cur_gen_dummy_magic_0.V_mir1.n18 ref_volt_cur_gen_dummy_magic_0.V_mir1.n17 40.7027
R6511 ref_volt_cur_gen_dummy_magic_0.V_mir1.n8 ref_volt_cur_gen_dummy_magic_0.V_mir1.n7 40.7027
R6512 ref_volt_cur_gen_dummy_magic_0.V_mir1.n3 ref_volt_cur_gen_dummy_magic_0.V_mir1.n2 40.7027
R6513 ref_volt_cur_gen_dummy_magic_0.V_mir1.n5 ref_volt_cur_gen_dummy_magic_0.V_mir1.t9 39.4005
R6514 ref_volt_cur_gen_dummy_magic_0.V_mir1.n5 ref_volt_cur_gen_dummy_magic_0.V_mir1.t5 39.4005
R6515 ref_volt_cur_gen_dummy_magic_0.V_mir1.n0 ref_volt_cur_gen_dummy_magic_0.V_mir1.t11 39.4005
R6516 ref_volt_cur_gen_dummy_magic_0.V_mir1.n0 ref_volt_cur_gen_dummy_magic_0.V_mir1.t7 39.4005
R6517 ref_volt_cur_gen_dummy_magic_0.V_mir1.t15 ref_volt_cur_gen_dummy_magic_0.V_mir1.n20 39.4005
R6518 ref_volt_cur_gen_dummy_magic_0.V_mir1.n20 ref_volt_cur_gen_dummy_magic_0.V_mir1.t13 39.4005
R6519 ref_volt_cur_gen_dummy_magic_0.V_mir1.n15 ref_volt_cur_gen_dummy_magic_0.V_mir1.n4 15.8005
R6520 ref_volt_cur_gen_dummy_magic_0.V_mir1.n19 ref_volt_cur_gen_dummy_magic_0.V_mir1.n15 15.8005
R6521 ref_volt_cur_gen_dummy_magic_0.V_mir1.n14 ref_volt_cur_gen_dummy_magic_0.V_mir1.n9 9.3005
R6522 ref_volt_cur_gen_dummy_magic_0.V_mir1.n13 ref_volt_cur_gen_dummy_magic_0.V_mir1.n12 5.8755
R6523 ref_volt_cur_gen_dummy_magic_0.V_mir1.n15 ref_volt_cur_gen_dummy_magic_0.V_mir1.n14 4.5005
R6524 ref_volt_cur_gen_dummy_magic_0.V_mir1.n14 ref_volt_cur_gen_dummy_magic_0.V_mir1.n13 0.78175
R6525 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t26 1172.87
R6526 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t35 1172.87
R6527 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.t45 996.134
R6528 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t34 996.134
R6529 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t48 996.134
R6530 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t38 996.134
R6531 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t51 996.134
R6532 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t27 996.134
R6533 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t43 996.134
R6534 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t30 996.134
R6535 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t29 690.867
R6536 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t40 690.867
R6537 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t54 530.201
R6538 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t33 530.201
R6539 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t39 514.134
R6540 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t49 514.134
R6541 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t36 514.134
R6542 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t46 514.134
R6543 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t31 514.134
R6544 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 514.134
R6545 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t41 514.134
R6546 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t52 514.134
R6547 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6548 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.t50 353.467
R6549 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t25 353.467
R6550 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t42 353.467
R6551 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t28 353.467
R6552 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t44 353.467
R6553 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t32 353.467
R6554 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t47 353.467
R6555 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 176.733
R6556 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R6557 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R6558 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R6559 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R6560 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.n47 176.733
R6561 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 176.733
R6562 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 176.733
R6563 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 176.733
R6564 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R6565 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6566 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6567 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 176.733
R6568 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6569 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R6570 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6571 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6572 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6573 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 166.436
R6574 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n31 161.875
R6575 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n40 161.686
R6576 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n0 160.427
R6577 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 159.802
R6578 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 159.802
R6579 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 159.802
R6580 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n1 159.802
R6581 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 155.302
R6582 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n13 114.689
R6583 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n12 114.689
R6584 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 114.126
R6585 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 114.126
R6586 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 114.126
R6587 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n11 109.626
R6588 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 51.9494
R6589 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R6590 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 51.9494
R6591 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n23 51.9494
R6592 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R6593 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n32 51.9494
R6594 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.X.n52 49.3036
R6595 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t22 16.0005
R6596 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R6597 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t8 16.0005
R6598 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t10 16.0005
R6599 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t9 16.0005
R6600 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R6601 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R6602 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t13 16.0005
R6603 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t12 16.0005
R6604 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t2 16.0005
R6605 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t6 16.0005
R6606 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t11 16.0005
R6607 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n42 15.7193
R6608 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t21 11.2576
R6609 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t18 11.2576
R6610 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t24 11.2576
R6611 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t20 11.2576
R6612 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t19 11.2576
R6613 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R6614 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t17 11.2576
R6615 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t16 11.2576
R6616 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t23 11.2576
R6617 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R6618 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R6619 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R6620 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n22 10.188
R6621 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 6.188
R6622 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n8 5.1255
R6623 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n20 4.5005
R6624 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 0.6255
R6625 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.6255
R6626 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.6255
R6627 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n15 0.563
R6628 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n17 0.563
R6629 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 0.563
R6630 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n10 0.5005
R6631 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 0.438
R6632 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 206.052
R6633 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 205.488
R6634 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 205.488
R6635 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 205.488
R6636 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 205.488
R6637 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 182.701
R6638 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 181.701
R6639 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 121.222
R6640 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 104.106
R6641 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 97.5005
R6642 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 85.2005
R6643 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 44.0317
R6644 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 19.7005
R6645 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R6646 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 19.7005
R6647 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R6648 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 19.7005
R6649 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R6650 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R6651 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R6652 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R6653 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R6654 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 15.7605
R6655 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 15.7605
R6656 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 15.7605
R6657 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 15.7605
R6658 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 15.7605
R6659 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 15.7605
R6660 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 6.09425
R6661 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 0.563
R6662 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 0.563
R6663 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 0.563
R6664 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t52 1172.87
R6665 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t27 1172.87
R6666 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t44 996.134
R6667 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6668 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t49 996.134
R6669 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t37 996.134
R6670 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R6671 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t36 996.134
R6672 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t42 996.134
R6673 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.t29 996.134
R6674 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t25 690.867
R6675 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t30 690.867
R6676 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t51 530.201
R6677 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t26 530.201
R6678 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t39 514.134
R6679 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t53 514.134
R6680 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t40 514.134
R6681 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R6682 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t38 514.134
R6683 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t50 514.134
R6684 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R6685 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 514.134
R6686 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t34 353.467
R6687 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R6688 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t28 353.467
R6689 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t43 353.467
R6690 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t31 353.467
R6691 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R6692 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t35 353.467
R6693 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t46 353.467
R6694 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R6695 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R6696 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R6697 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R6698 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R6699 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 176.733
R6700 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R6701 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6702 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6703 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6704 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R6705 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R6706 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R6707 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R6708 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R6709 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R6710 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R6711 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R6712 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 166.375
R6713 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.875
R6714 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.686
R6715 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n0 160.427
R6716 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n7 159.802
R6717 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 159.802
R6718 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 159.802
R6719 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n1 159.802
R6720 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 155.302
R6721 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 114.689
R6722 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n12 114.689
R6723 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 114.126
R6724 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n15 114.126
R6725 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 114.126
R6726 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n11 109.626
R6727 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R6728 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n42 51.9494
R6729 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R6730 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n28 51.9494
R6731 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R6732 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n37 51.9494
R6733 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t4 49.2412
R6734 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R6735 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R6736 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t8 16.0005
R6737 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R6738 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t0 16.0005
R6739 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t16 16.0005
R6740 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R6741 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t12 16.0005
R6742 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t14 16.0005
R6743 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t2 16.0005
R6744 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t24 16.0005
R6745 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t3 16.0005
R6746 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 15.6567
R6747 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t18 11.2576
R6748 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t7 11.2576
R6749 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t10 11.2576
R6750 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t23 11.2576
R6751 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t17 11.2576
R6752 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t20 11.2576
R6753 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t19 11.2576
R6754 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t22 11.2576
R6755 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t13 11.2576
R6756 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t21 11.2576
R6757 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t9 11.2576
R6758 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t11 11.2576
R6759 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n51 10.313
R6760 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n40 6.063
R6761 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n8 5.1255
R6762 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 4.5005
R6763 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n2 0.6255
R6764 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n4 0.6255
R6765 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n6 0.6255
R6766 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n14 0.563
R6767 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n16 0.563
R6768 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n18 0.563
R6769 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n10 0.5005
R6770 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n21 0.438
R6771 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 145.702
R6772 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 134.577
R6773 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 108.66
R6774 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 97.4009
R6775 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 96.8384
R6776 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 96.8384
R6777 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 96.8384
R6778 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 96.8384
R6779 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 73.063
R6780 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R6781 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 24.0005
R6782 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 24.0005
R6783 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 24.0005
R6784 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 18.4067
R6785 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R6786 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R6787 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R6788 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 8.0005
R6789 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R6790 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 8.0005
R6791 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R6792 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 8.0005
R6793 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R6794 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R6795 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 2.71925
R6796 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 0.563
R6797 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 0.563
R6798 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.563
R6799 ref_volt_cur_gen_dummy_magic_0.V_TOP.n0 ref_volt_cur_gen_dummy_magic_0.V_TOP.t16 369.534
R6800 ref_volt_cur_gen_dummy_magic_0.V_TOP.n10 ref_volt_cur_gen_dummy_magic_0.V_TOP.n8 339.959
R6801 ref_volt_cur_gen_dummy_magic_0.V_TOP.n7 ref_volt_cur_gen_dummy_magic_0.V_TOP.n6 339.272
R6802 ref_volt_cur_gen_dummy_magic_0.V_TOP.n15 ref_volt_cur_gen_dummy_magic_0.V_TOP.n14 339.272
R6803 ref_volt_cur_gen_dummy_magic_0.V_TOP.n17 ref_volt_cur_gen_dummy_magic_0.V_TOP.n16 339.272
R6804 ref_volt_cur_gen_dummy_magic_0.V_TOP.n10 ref_volt_cur_gen_dummy_magic_0.V_TOP.n9 339.272
R6805 ref_volt_cur_gen_dummy_magic_0.V_TOP.n12 ref_volt_cur_gen_dummy_magic_0.V_TOP.n11 334.772
R6806 ref_volt_cur_gen_dummy_magic_0.V_TOP.n1 ref_volt_cur_gen_dummy_magic_0.V_TOP.n0 224.934
R6807 ref_volt_cur_gen_dummy_magic_0.V_TOP.n2 ref_volt_cur_gen_dummy_magic_0.V_TOP.n1 224.934
R6808 ref_volt_cur_gen_dummy_magic_0.V_TOP.n3 ref_volt_cur_gen_dummy_magic_0.V_TOP.n2 224.934
R6809 ref_volt_cur_gen_dummy_magic_0.V_TOP.n4 ref_volt_cur_gen_dummy_magic_0.V_TOP.n3 224.934
R6810 ref_volt_cur_gen_dummy_magic_0.V_TOP.n5 ref_volt_cur_gen_dummy_magic_0.V_TOP.n4 224.934
R6811 ref_volt_cur_gen_dummy_magic_0.V_TOP.n27 ref_volt_cur_gen_dummy_magic_0.V_TOP.n26 224.934
R6812 ref_volt_cur_gen_dummy_magic_0.V_TOP.n26 ref_volt_cur_gen_dummy_magic_0.V_TOP.n25 224.934
R6813 ref_volt_cur_gen_dummy_magic_0.V_TOP.n25 ref_volt_cur_gen_dummy_magic_0.V_TOP.n24 224.934
R6814 ref_volt_cur_gen_dummy_magic_0.V_TOP.n24 ref_volt_cur_gen_dummy_magic_0.V_TOP.n23 224.934
R6815 ref_volt_cur_gen_dummy_magic_0.V_TOP.n23 ref_volt_cur_gen_dummy_magic_0.V_TOP.n22 224.934
R6816 ref_volt_cur_gen_dummy_magic_0.V_TOP.n22 ref_volt_cur_gen_dummy_magic_0.V_TOP.n21 224.934
R6817 ref_volt_cur_gen_dummy_magic_0.V_TOP.n21 ref_volt_cur_gen_dummy_magic_0.V_TOP.n20 224.934
R6818 ref_volt_cur_gen_dummy_magic_0.V_TOP ref_volt_cur_gen_dummy_magic_0.V_TOP.t48 214.222
R6819 ref_volt_cur_gen_dummy_magic_0.V_TOP ref_volt_cur_gen_dummy_magic_0.V_TOP.n40 204.002
R6820 ref_volt_cur_gen_dummy_magic_0.V_TOP.n7 ref_volt_cur_gen_dummy_magic_0.V_TOP.t13 176.114
R6821 ref_volt_cur_gen_dummy_magic_0.V_TOP.n19 ref_volt_cur_gen_dummy_magic_0.V_TOP.n18 163.175
R6822 ref_volt_cur_gen_dummy_magic_0.V_TOP.n0 ref_volt_cur_gen_dummy_magic_0.V_TOP.t49 144.601
R6823 ref_volt_cur_gen_dummy_magic_0.V_TOP.n1 ref_volt_cur_gen_dummy_magic_0.V_TOP.t42 144.601
R6824 ref_volt_cur_gen_dummy_magic_0.V_TOP.n2 ref_volt_cur_gen_dummy_magic_0.V_TOP.t37 144.601
R6825 ref_volt_cur_gen_dummy_magic_0.V_TOP.n3 ref_volt_cur_gen_dummy_magic_0.V_TOP.t24 144.601
R6826 ref_volt_cur_gen_dummy_magic_0.V_TOP.n4 ref_volt_cur_gen_dummy_magic_0.V_TOP.t46 144.601
R6827 ref_volt_cur_gen_dummy_magic_0.V_TOP.n5 ref_volt_cur_gen_dummy_magic_0.V_TOP.t40 144.601
R6828 ref_volt_cur_gen_dummy_magic_0.V_TOP.n27 ref_volt_cur_gen_dummy_magic_0.V_TOP.t15 144.601
R6829 ref_volt_cur_gen_dummy_magic_0.V_TOP.n26 ref_volt_cur_gen_dummy_magic_0.V_TOP.t25 144.601
R6830 ref_volt_cur_gen_dummy_magic_0.V_TOP.n25 ref_volt_cur_gen_dummy_magic_0.V_TOP.t30 144.601
R6831 ref_volt_cur_gen_dummy_magic_0.V_TOP.n24 ref_volt_cur_gen_dummy_magic_0.V_TOP.t35 144.601
R6832 ref_volt_cur_gen_dummy_magic_0.V_TOP.n23 ref_volt_cur_gen_dummy_magic_0.V_TOP.t17 144.601
R6833 ref_volt_cur_gen_dummy_magic_0.V_TOP.n22 ref_volt_cur_gen_dummy_magic_0.V_TOP.t22 144.601
R6834 ref_volt_cur_gen_dummy_magic_0.V_TOP.n21 ref_volt_cur_gen_dummy_magic_0.V_TOP.t31 144.601
R6835 ref_volt_cur_gen_dummy_magic_0.V_TOP.n20 ref_volt_cur_gen_dummy_magic_0.V_TOP.t36 144.601
R6836 ref_volt_cur_gen_dummy_magic_0.V_TOP.n18 ref_volt_cur_gen_dummy_magic_0.V_TOP.t6 95.447
R6837 ref_volt_cur_gen_dummy_magic_0.V_TOP.n19 ref_volt_cur_gen_dummy_magic_0.V_TOP.n5 69.6227
R6838 ref_volt_cur_gen_dummy_magic_0.V_TOP ref_volt_cur_gen_dummy_magic_0.V_TOP.n27 69.6227
R6839 ref_volt_cur_gen_dummy_magic_0.V_TOP.n20 ref_volt_cur_gen_dummy_magic_0.V_TOP.n19 69.6227
R6840 ref_volt_cur_gen_dummy_magic_0.V_TOP.n6 ref_volt_cur_gen_dummy_magic_0.V_TOP.t12 39.4005
R6841 ref_volt_cur_gen_dummy_magic_0.V_TOP.n6 ref_volt_cur_gen_dummy_magic_0.V_TOP.t4 39.4005
R6842 ref_volt_cur_gen_dummy_magic_0.V_TOP.n11 ref_volt_cur_gen_dummy_magic_0.V_TOP.t10 39.4005
R6843 ref_volt_cur_gen_dummy_magic_0.V_TOP.n11 ref_volt_cur_gen_dummy_magic_0.V_TOP.t7 39.4005
R6844 ref_volt_cur_gen_dummy_magic_0.V_TOP.n9 ref_volt_cur_gen_dummy_magic_0.V_TOP.t2 39.4005
R6845 ref_volt_cur_gen_dummy_magic_0.V_TOP.n9 ref_volt_cur_gen_dummy_magic_0.V_TOP.t1 39.4005
R6846 ref_volt_cur_gen_dummy_magic_0.V_TOP.n8 ref_volt_cur_gen_dummy_magic_0.V_TOP.t0 39.4005
R6847 ref_volt_cur_gen_dummy_magic_0.V_TOP.n8 ref_volt_cur_gen_dummy_magic_0.V_TOP.t3 39.4005
R6848 ref_volt_cur_gen_dummy_magic_0.V_TOP.n14 ref_volt_cur_gen_dummy_magic_0.V_TOP.t11 39.4005
R6849 ref_volt_cur_gen_dummy_magic_0.V_TOP.n14 ref_volt_cur_gen_dummy_magic_0.V_TOP.t8 39.4005
R6850 ref_volt_cur_gen_dummy_magic_0.V_TOP.n16 ref_volt_cur_gen_dummy_magic_0.V_TOP.t5 39.4005
R6851 ref_volt_cur_gen_dummy_magic_0.V_TOP.n16 ref_volt_cur_gen_dummy_magic_0.V_TOP.t9 39.4005
R6852 ref_volt_cur_gen_dummy_magic_0.V_TOP.n12 ref_volt_cur_gen_dummy_magic_0.V_TOP.n10 8.313
R6853 ref_volt_cur_gen_dummy_magic_0.V_TOP.n18 ref_volt_cur_gen_dummy_magic_0.V_TOP.n17 5.188
R6854 ref_volt_cur_gen_dummy_magic_0.V_TOP.n28 ref_volt_cur_gen_dummy_magic_0.V_TOP.t29 4.8295
R6855 ref_volt_cur_gen_dummy_magic_0.V_TOP.n29 ref_volt_cur_gen_dummy_magic_0.V_TOP.t20 4.8295
R6856 ref_volt_cur_gen_dummy_magic_0.V_TOP.n31 ref_volt_cur_gen_dummy_magic_0.V_TOP.t39 4.8295
R6857 ref_volt_cur_gen_dummy_magic_0.V_TOP.n32 ref_volt_cur_gen_dummy_magic_0.V_TOP.t26 4.8295
R6858 ref_volt_cur_gen_dummy_magic_0.V_TOP.n34 ref_volt_cur_gen_dummy_magic_0.V_TOP.t28 4.8295
R6859 ref_volt_cur_gen_dummy_magic_0.V_TOP.n35 ref_volt_cur_gen_dummy_magic_0.V_TOP.t18 4.8295
R6860 ref_volt_cur_gen_dummy_magic_0.V_TOP.n37 ref_volt_cur_gen_dummy_magic_0.V_TOP.t43 4.8295
R6861 ref_volt_cur_gen_dummy_magic_0.V_TOP.n28 ref_volt_cur_gen_dummy_magic_0.V_TOP.t41 4.5005
R6862 ref_volt_cur_gen_dummy_magic_0.V_TOP.n30 ref_volt_cur_gen_dummy_magic_0.V_TOP.t34 4.5005
R6863 ref_volt_cur_gen_dummy_magic_0.V_TOP.n29 ref_volt_cur_gen_dummy_magic_0.V_TOP.t47 4.5005
R6864 ref_volt_cur_gen_dummy_magic_0.V_TOP.n31 ref_volt_cur_gen_dummy_magic_0.V_TOP.t14 4.5005
R6865 ref_volt_cur_gen_dummy_magic_0.V_TOP.n33 ref_volt_cur_gen_dummy_magic_0.V_TOP.t45 4.5005
R6866 ref_volt_cur_gen_dummy_magic_0.V_TOP.n32 ref_volt_cur_gen_dummy_magic_0.V_TOP.t19 4.5005
R6867 ref_volt_cur_gen_dummy_magic_0.V_TOP.n34 ref_volt_cur_gen_dummy_magic_0.V_TOP.t38 4.5005
R6868 ref_volt_cur_gen_dummy_magic_0.V_TOP.n36 ref_volt_cur_gen_dummy_magic_0.V_TOP.t33 4.5005
R6869 ref_volt_cur_gen_dummy_magic_0.V_TOP.n35 ref_volt_cur_gen_dummy_magic_0.V_TOP.t44 4.5005
R6870 ref_volt_cur_gen_dummy_magic_0.V_TOP.n40 ref_volt_cur_gen_dummy_magic_0.V_TOP.t21 4.5005
R6871 ref_volt_cur_gen_dummy_magic_0.V_TOP.n39 ref_volt_cur_gen_dummy_magic_0.V_TOP.t27 4.5005
R6872 ref_volt_cur_gen_dummy_magic_0.V_TOP.n38 ref_volt_cur_gen_dummy_magic_0.V_TOP.t23 4.5005
R6873 ref_volt_cur_gen_dummy_magic_0.V_TOP.n37 ref_volt_cur_gen_dummy_magic_0.V_TOP.t32 4.5005
R6874 ref_volt_cur_gen_dummy_magic_0.V_TOP.n13 ref_volt_cur_gen_dummy_magic_0.V_TOP.n12 4.5005
R6875 ref_volt_cur_gen_dummy_magic_0.V_TOP.n17 ref_volt_cur_gen_dummy_magic_0.V_TOP.n15 2.1255
R6876 ref_volt_cur_gen_dummy_magic_0.V_TOP.n15 ref_volt_cur_gen_dummy_magic_0.V_TOP.n13 2.1255
R6877 ref_volt_cur_gen_dummy_magic_0.V_TOP.n13 ref_volt_cur_gen_dummy_magic_0.V_TOP.n7 2.1255
R6878 ref_volt_cur_gen_dummy_magic_0.V_TOP.n30 ref_volt_cur_gen_dummy_magic_0.V_TOP.n28 0.3295
R6879 ref_volt_cur_gen_dummy_magic_0.V_TOP.n30 ref_volt_cur_gen_dummy_magic_0.V_TOP.n29 0.3295
R6880 ref_volt_cur_gen_dummy_magic_0.V_TOP.n33 ref_volt_cur_gen_dummy_magic_0.V_TOP.n31 0.3295
R6881 ref_volt_cur_gen_dummy_magic_0.V_TOP.n33 ref_volt_cur_gen_dummy_magic_0.V_TOP.n32 0.3295
R6882 ref_volt_cur_gen_dummy_magic_0.V_TOP.n36 ref_volt_cur_gen_dummy_magic_0.V_TOP.n34 0.3295
R6883 ref_volt_cur_gen_dummy_magic_0.V_TOP.n36 ref_volt_cur_gen_dummy_magic_0.V_TOP.n35 0.3295
R6884 ref_volt_cur_gen_dummy_magic_0.V_TOP.n40 ref_volt_cur_gen_dummy_magic_0.V_TOP.n39 0.3295
R6885 ref_volt_cur_gen_dummy_magic_0.V_TOP.n39 ref_volt_cur_gen_dummy_magic_0.V_TOP.n38 0.3295
R6886 ref_volt_cur_gen_dummy_magic_0.V_TOP.n38 ref_volt_cur_gen_dummy_magic_0.V_TOP.n37 0.3295
R6887 ref_volt_cur_gen_dummy_magic_0.V_TOP.n33 ref_volt_cur_gen_dummy_magic_0.V_TOP.n30 0.2825
R6888 ref_volt_cur_gen_dummy_magic_0.V_TOP.n36 ref_volt_cur_gen_dummy_magic_0.V_TOP.n33 0.2825
R6889 ref_volt_cur_gen_dummy_magic_0.V_TOP.n38 ref_volt_cur_gen_dummy_magic_0.V_TOP.n36 0.2825
R6890 ref_volt_cur_gen_dummy_magic_0.V_p_2.n1 ref_volt_cur_gen_dummy_magic_0.V_p_2.n5 229.562
R6891 ref_volt_cur_gen_dummy_magic_0.V_p_2.n1 ref_volt_cur_gen_dummy_magic_0.V_p_2.n4 228.939
R6892 ref_volt_cur_gen_dummy_magic_0.V_p_2.n0 ref_volt_cur_gen_dummy_magic_0.V_p_2.n3 228.939
R6893 ref_volt_cur_gen_dummy_magic_0.V_p_2.n0 ref_volt_cur_gen_dummy_magic_0.V_p_2.n2 228.939
R6894 ref_volt_cur_gen_dummy_magic_0.V_p_2.n6 ref_volt_cur_gen_dummy_magic_0.V_p_2.n1 228.938
R6895 ref_volt_cur_gen_dummy_magic_0.V_p_2.n0 ref_volt_cur_gen_dummy_magic_0.V_p_2.t1 98.2282
R6896 ref_volt_cur_gen_dummy_magic_0.V_p_2.n5 ref_volt_cur_gen_dummy_magic_0.V_p_2.t2 48.0005
R6897 ref_volt_cur_gen_dummy_magic_0.V_p_2.n5 ref_volt_cur_gen_dummy_magic_0.V_p_2.t7 48.0005
R6898 ref_volt_cur_gen_dummy_magic_0.V_p_2.n4 ref_volt_cur_gen_dummy_magic_0.V_p_2.t4 48.0005
R6899 ref_volt_cur_gen_dummy_magic_0.V_p_2.n4 ref_volt_cur_gen_dummy_magic_0.V_p_2.t10 48.0005
R6900 ref_volt_cur_gen_dummy_magic_0.V_p_2.n3 ref_volt_cur_gen_dummy_magic_0.V_p_2.t6 48.0005
R6901 ref_volt_cur_gen_dummy_magic_0.V_p_2.n3 ref_volt_cur_gen_dummy_magic_0.V_p_2.t0 48.0005
R6902 ref_volt_cur_gen_dummy_magic_0.V_p_2.n2 ref_volt_cur_gen_dummy_magic_0.V_p_2.t5 48.0005
R6903 ref_volt_cur_gen_dummy_magic_0.V_p_2.n2 ref_volt_cur_gen_dummy_magic_0.V_p_2.t8 48.0005
R6904 ref_volt_cur_gen_dummy_magic_0.V_p_2.t9 ref_volt_cur_gen_dummy_magic_0.V_p_2.n6 48.0005
R6905 ref_volt_cur_gen_dummy_magic_0.V_p_2.n6 ref_volt_cur_gen_dummy_magic_0.V_p_2.t3 48.0005
R6906 ref_volt_cur_gen_dummy_magic_0.V_p_2.n1 ref_volt_cur_gen_dummy_magic_0.V_p_2.n0 1.8755
R6907 VOUT+.n2 VOUT+.n0 145.989
R6908 VOUT+.n8 VOUT+.n7 145.989
R6909 VOUT+.n6 VOUT+.n5 145.427
R6910 VOUT+.n4 VOUT+.n3 145.427
R6911 VOUT+.n2 VOUT+.n1 145.427
R6912 VOUT+.n10 VOUT+.n9 140.927
R6913 VOUT+.n100 VOUT+.t2 113.192
R6914 VOUT+.n97 VOUT+.n95 95.7303
R6915 VOUT+.n99 VOUT+.n98 94.6053
R6916 VOUT+.n97 VOUT+.n96 94.6053
R6917 VOUT+.n94 VOUT+.n10 20.5943
R6918 VOUT+.n94 VOUT+.n93 11.7059
R6919 VOUT+ VOUT+.n94 7.813
R6920 VOUT+.n9 VOUT+.t7 6.56717
R6921 VOUT+.n9 VOUT+.t11 6.56717
R6922 VOUT+.n7 VOUT+.t5 6.56717
R6923 VOUT+.n7 VOUT+.t4 6.56717
R6924 VOUT+.n5 VOUT+.t6 6.56717
R6925 VOUT+.n5 VOUT+.t10 6.56717
R6926 VOUT+.n3 VOUT+.t8 6.56717
R6927 VOUT+.n3 VOUT+.t12 6.56717
R6928 VOUT+.n1 VOUT+.t9 6.56717
R6929 VOUT+.n1 VOUT+.t13 6.56717
R6930 VOUT+.n0 VOUT+.t3 6.56717
R6931 VOUT+.n0 VOUT+.t14 6.56717
R6932 VOUT+.n40 VOUT+.t108 4.8295
R6933 VOUT+.n52 VOUT+.t25 4.8295
R6934 VOUT+.n49 VOUT+.t76 4.8295
R6935 VOUT+.n46 VOUT+.t113 4.8295
R6936 VOUT+.n43 VOUT+.t145 4.8295
R6937 VOUT+.n42 VOUT+.t68 4.8295
R6938 VOUT+.n66 VOUT+.t28 4.8295
R6939 VOUT+.n67 VOUT+.t77 4.8295
R6940 VOUT+.n69 VOUT+.t63 4.8295
R6941 VOUT+.n70 VOUT+.t111 4.8295
R6942 VOUT+.n72 VOUT+.t114 4.8295
R6943 VOUT+.n73 VOUT+.t99 4.8295
R6944 VOUT+.n75 VOUT+.t74 4.8295
R6945 VOUT+.n76 VOUT+.t56 4.8295
R6946 VOUT+.n78 VOUT+.t109 4.8295
R6947 VOUT+.n79 VOUT+.t92 4.8295
R6948 VOUT+.n81 VOUT+.t69 4.8295
R6949 VOUT+.n82 VOUT+.t53 4.8295
R6950 VOUT+.n84 VOUT+.t30 4.8295
R6951 VOUT+.n85 VOUT+.t153 4.8295
R6952 VOUT+.n87 VOUT+.t64 4.8295
R6953 VOUT+.n88 VOUT+.t47 4.8295
R6954 VOUT+.n11 VOUT+.t117 4.8295
R6955 VOUT+.n13 VOUT+.t72 4.8295
R6956 VOUT+.n25 VOUT+.t38 4.8295
R6957 VOUT+.n26 VOUT+.t20 4.8295
R6958 VOUT+.n28 VOUT+.t80 4.8295
R6959 VOUT+.n29 VOUT+.t61 4.8295
R6960 VOUT+.n31 VOUT+.t121 4.8295
R6961 VOUT+.n32 VOUT+.t104 4.8295
R6962 VOUT+.n34 VOUT+.t85 4.8295
R6963 VOUT+.n35 VOUT+.t67 4.8295
R6964 VOUT+.n37 VOUT+.t123 4.8295
R6965 VOUT+.n38 VOUT+.t107 4.8295
R6966 VOUT+.n90 VOUT+.t22 4.8295
R6967 VOUT+.n55 VOUT+.t33 4.806
R6968 VOUT+.n56 VOUT+.t150 4.806
R6969 VOUT+.n57 VOUT+.t51 4.806
R6970 VOUT+.n58 VOUT+.t88 4.806
R6971 VOUT+.n59 VOUT+.t125 4.806
R6972 VOUT+.n60 VOUT+.t105 4.806
R6973 VOUT+.n61 VOUT+.t140 4.806
R6974 VOUT+.n62 VOUT+.t37 4.806
R6975 VOUT+.n63 VOUT+.t156 4.806
R6976 VOUT+.n64 VOUT+.t54 4.806
R6977 VOUT+.n14 VOUT+.t73 4.806
R6978 VOUT+.n15 VOUT+.t116 4.806
R6979 VOUT+.n16 VOUT+.t65 4.806
R6980 VOUT+.n17 VOUT+.t154 4.806
R6981 VOUT+.n18 VOUT+.t106 4.806
R6982 VOUT+.n19 VOUT+.t143 4.806
R6983 VOUT+.n20 VOUT+.t96 4.806
R6984 VOUT+.n21 VOUT+.t43 4.806
R6985 VOUT+.n22 VOUT+.t87 4.806
R6986 VOUT+.n23 VOUT+.t35 4.806
R6987 VOUT+.n40 VOUT+.t70 4.5005
R6988 VOUT+.n41 VOUT+.t91 4.5005
R6989 VOUT+.n52 VOUT+.t66 4.5005
R6990 VOUT+.n53 VOUT+.t81 4.5005
R6991 VOUT+.n54 VOUT+.t44 4.5005
R6992 VOUT+.n49 VOUT+.t118 4.5005
R6993 VOUT+.n50 VOUT+.t57 4.5005
R6994 VOUT+.n51 VOUT+.t21 4.5005
R6995 VOUT+.n46 VOUT+.t151 4.5005
R6996 VOUT+.n47 VOUT+.t98 4.5005
R6997 VOUT+.n48 VOUT+.t60 4.5005
R6998 VOUT+.n43 VOUT+.t45 4.5005
R6999 VOUT+.n44 VOUT+.t136 4.5005
R7000 VOUT+.n45 VOUT+.t101 4.5005
R7001 VOUT+.n42 VOUT+.t31 4.5005
R7002 VOUT+.n65 VOUT+.t52 4.5005
R7003 VOUT+.n64 VOUT+.t155 4.5005
R7004 VOUT+.n63 VOUT+.t119 4.5005
R7005 VOUT+.n62 VOUT+.t139 4.5005
R7006 VOUT+.n61 VOUT+.t102 4.5005
R7007 VOUT+.n60 VOUT+.t62 4.5005
R7008 VOUT+.n59 VOUT+.t86 4.5005
R7009 VOUT+.n58 VOUT+.t46 4.5005
R7010 VOUT+.n57 VOUT+.t147 4.5005
R7011 VOUT+.n56 VOUT+.t110 4.5005
R7012 VOUT+.n55 VOUT+.t134 4.5005
R7013 VOUT+.n66 VOUT+.t130 4.5005
R7014 VOUT+.n68 VOUT+.t152 4.5005
R7015 VOUT+.n67 VOUT+.t115 4.5005
R7016 VOUT+.n69 VOUT+.t23 4.5005
R7017 VOUT+.n71 VOUT+.t48 4.5005
R7018 VOUT+.n70 VOUT+.t148 4.5005
R7019 VOUT+.n72 VOUT+.t79 4.5005
R7020 VOUT+.n74 VOUT+.t27 4.5005
R7021 VOUT+.n73 VOUT+.t132 4.5005
R7022 VOUT+.n75 VOUT+.t40 4.5005
R7023 VOUT+.n77 VOUT+.t128 4.5005
R7024 VOUT+.n76 VOUT+.t93 4.5005
R7025 VOUT+.n78 VOUT+.t71 4.5005
R7026 VOUT+.n80 VOUT+.t19 4.5005
R7027 VOUT+.n79 VOUT+.t126 4.5005
R7028 VOUT+.n81 VOUT+.t34 4.5005
R7029 VOUT+.n83 VOUT+.t122 4.5005
R7030 VOUT+.n82 VOUT+.t89 4.5005
R7031 VOUT+.n84 VOUT+.t135 4.5005
R7032 VOUT+.n86 VOUT+.t83 4.5005
R7033 VOUT+.n85 VOUT+.t49 4.5005
R7034 VOUT+.n87 VOUT+.t29 4.5005
R7035 VOUT+.n89 VOUT+.t120 4.5005
R7036 VOUT+.n88 VOUT+.t82 4.5005
R7037 VOUT+.n11 VOUT+.t26 4.5005
R7038 VOUT+.n12 VOUT+.t124 4.5005
R7039 VOUT+.n13 VOUT+.t39 4.5005
R7040 VOUT+.n24 VOUT+.t127 4.5005
R7041 VOUT+.n23 VOUT+.t95 4.5005
R7042 VOUT+.n22 VOUT+.t55 4.5005
R7043 VOUT+.n21 VOUT+.t144 4.5005
R7044 VOUT+.n20 VOUT+.t112 4.5005
R7045 VOUT+.n19 VOUT+.t75 4.5005
R7046 VOUT+.n18 VOUT+.t24 4.5005
R7047 VOUT+.n17 VOUT+.t131 4.5005
R7048 VOUT+.n16 VOUT+.t97 4.5005
R7049 VOUT+.n15 VOUT+.t59 4.5005
R7050 VOUT+.n14 VOUT+.t149 4.5005
R7051 VOUT+.n25 VOUT+.t142 4.5005
R7052 VOUT+.n27 VOUT+.t94 4.5005
R7053 VOUT+.n26 VOUT+.t58 4.5005
R7054 VOUT+.n28 VOUT+.t42 4.5005
R7055 VOUT+.n30 VOUT+.t133 4.5005
R7056 VOUT+.n29 VOUT+.t100 4.5005
R7057 VOUT+.n31 VOUT+.t84 4.5005
R7058 VOUT+.n33 VOUT+.t32 4.5005
R7059 VOUT+.n32 VOUT+.t137 4.5005
R7060 VOUT+.n34 VOUT+.t50 4.5005
R7061 VOUT+.n36 VOUT+.t138 4.5005
R7062 VOUT+.n35 VOUT+.t103 4.5005
R7063 VOUT+.n37 VOUT+.t90 4.5005
R7064 VOUT+.n39 VOUT+.t36 4.5005
R7065 VOUT+.n38 VOUT+.t141 4.5005
R7066 VOUT+.n90 VOUT+.t129 4.5005
R7067 VOUT+.n91 VOUT+.t78 4.5005
R7068 VOUT+.n92 VOUT+.t41 4.5005
R7069 VOUT+.n93 VOUT+.t146 4.5005
R7070 VOUT+.n10 VOUT+.n8 4.5005
R7071 VOUT+.n98 VOUT+.t18 3.42907
R7072 VOUT+.n98 VOUT+.t16 3.42907
R7073 VOUT+.n96 VOUT+.t1 3.42907
R7074 VOUT+.n96 VOUT+.t0 3.42907
R7075 VOUT+.n95 VOUT+.t15 3.42907
R7076 VOUT+.n95 VOUT+.t17 3.42907
R7077 VOUT+ VOUT+.n100 2.84425
R7078 VOUT+.n100 VOUT+.n99 2.03175
R7079 VOUT+.n99 VOUT+.n97 1.1255
R7080 VOUT+.n4 VOUT+.n2 0.563
R7081 VOUT+.n6 VOUT+.n4 0.563
R7082 VOUT+.n8 VOUT+.n6 0.563
R7083 VOUT+.n41 VOUT+.n40 0.3295
R7084 VOUT+.n54 VOUT+.n53 0.3295
R7085 VOUT+.n53 VOUT+.n52 0.3295
R7086 VOUT+.n51 VOUT+.n50 0.3295
R7087 VOUT+.n50 VOUT+.n49 0.3295
R7088 VOUT+.n48 VOUT+.n47 0.3295
R7089 VOUT+.n47 VOUT+.n46 0.3295
R7090 VOUT+.n45 VOUT+.n44 0.3295
R7091 VOUT+.n44 VOUT+.n43 0.3295
R7092 VOUT+.n65 VOUT+.n42 0.3295
R7093 VOUT+.n65 VOUT+.n64 0.3295
R7094 VOUT+.n64 VOUT+.n63 0.3295
R7095 VOUT+.n63 VOUT+.n62 0.3295
R7096 VOUT+.n62 VOUT+.n61 0.3295
R7097 VOUT+.n61 VOUT+.n60 0.3295
R7098 VOUT+.n60 VOUT+.n59 0.3295
R7099 VOUT+.n59 VOUT+.n58 0.3295
R7100 VOUT+.n58 VOUT+.n57 0.3295
R7101 VOUT+.n57 VOUT+.n56 0.3295
R7102 VOUT+.n56 VOUT+.n55 0.3295
R7103 VOUT+.n68 VOUT+.n66 0.3295
R7104 VOUT+.n68 VOUT+.n67 0.3295
R7105 VOUT+.n71 VOUT+.n69 0.3295
R7106 VOUT+.n71 VOUT+.n70 0.3295
R7107 VOUT+.n74 VOUT+.n72 0.3295
R7108 VOUT+.n74 VOUT+.n73 0.3295
R7109 VOUT+.n77 VOUT+.n75 0.3295
R7110 VOUT+.n77 VOUT+.n76 0.3295
R7111 VOUT+.n80 VOUT+.n78 0.3295
R7112 VOUT+.n80 VOUT+.n79 0.3295
R7113 VOUT+.n83 VOUT+.n81 0.3295
R7114 VOUT+.n83 VOUT+.n82 0.3295
R7115 VOUT+.n86 VOUT+.n84 0.3295
R7116 VOUT+.n86 VOUT+.n85 0.3295
R7117 VOUT+.n89 VOUT+.n87 0.3295
R7118 VOUT+.n89 VOUT+.n88 0.3295
R7119 VOUT+.n12 VOUT+.n11 0.3295
R7120 VOUT+.n24 VOUT+.n13 0.3295
R7121 VOUT+.n24 VOUT+.n23 0.3295
R7122 VOUT+.n23 VOUT+.n22 0.3295
R7123 VOUT+.n22 VOUT+.n21 0.3295
R7124 VOUT+.n21 VOUT+.n20 0.3295
R7125 VOUT+.n20 VOUT+.n19 0.3295
R7126 VOUT+.n19 VOUT+.n18 0.3295
R7127 VOUT+.n18 VOUT+.n17 0.3295
R7128 VOUT+.n17 VOUT+.n16 0.3295
R7129 VOUT+.n16 VOUT+.n15 0.3295
R7130 VOUT+.n15 VOUT+.n14 0.3295
R7131 VOUT+.n27 VOUT+.n25 0.3295
R7132 VOUT+.n27 VOUT+.n26 0.3295
R7133 VOUT+.n30 VOUT+.n28 0.3295
R7134 VOUT+.n30 VOUT+.n29 0.3295
R7135 VOUT+.n33 VOUT+.n31 0.3295
R7136 VOUT+.n33 VOUT+.n32 0.3295
R7137 VOUT+.n36 VOUT+.n34 0.3295
R7138 VOUT+.n36 VOUT+.n35 0.3295
R7139 VOUT+.n39 VOUT+.n37 0.3295
R7140 VOUT+.n39 VOUT+.n38 0.3295
R7141 VOUT+.n91 VOUT+.n90 0.3295
R7142 VOUT+.n92 VOUT+.n91 0.3295
R7143 VOUT+.n93 VOUT+.n92 0.3295
R7144 VOUT+.n59 VOUT+.n54 0.306
R7145 VOUT+.n60 VOUT+.n51 0.306
R7146 VOUT+.n61 VOUT+.n48 0.306
R7147 VOUT+.n62 VOUT+.n45 0.306
R7148 VOUT+.n65 VOUT+.n41 0.2825
R7149 VOUT+.n68 VOUT+.n65 0.2825
R7150 VOUT+.n71 VOUT+.n68 0.2825
R7151 VOUT+.n74 VOUT+.n71 0.2825
R7152 VOUT+.n77 VOUT+.n74 0.2825
R7153 VOUT+.n80 VOUT+.n77 0.2825
R7154 VOUT+.n83 VOUT+.n80 0.2825
R7155 VOUT+.n86 VOUT+.n83 0.2825
R7156 VOUT+.n89 VOUT+.n86 0.2825
R7157 VOUT+.n24 VOUT+.n12 0.2825
R7158 VOUT+.n27 VOUT+.n24 0.2825
R7159 VOUT+.n30 VOUT+.n27 0.2825
R7160 VOUT+.n33 VOUT+.n30 0.2825
R7161 VOUT+.n36 VOUT+.n33 0.2825
R7162 VOUT+.n39 VOUT+.n36 0.2825
R7163 VOUT+.n91 VOUT+.n39 0.2825
R7164 VOUT+.n91 VOUT+.n89 0.2825
R7165 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 49.2006
R7166 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1603
R7167 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R7168 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1603
R7169 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.1603
R7170 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R7171 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.1603
R7172 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1603
R7173 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R7174 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R7175 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R7176 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.1603
R7177 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R7178 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.1603
R7179 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R7180 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1603
R7181 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1603
R7182 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1603
R7183 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.1603
R7184 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.1603
R7185 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1603
R7186 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.1603
R7187 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R7188 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1603
R7189 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1603
R7190 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1603
R7191 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R7192 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.1603
R7193 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1603
R7194 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R7195 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.1603
R7196 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R7197 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1603
R7198 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R7199 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1603
R7200 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R7201 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R7202 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R7203 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1603
R7204 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R7205 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R7206 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R7207 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.1603
R7208 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R7209 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R7210 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.1603
R7211 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R7212 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.1603
R7213 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R7214 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R7215 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R7216 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1603
R7217 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.1603
R7218 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1603
R7219 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R7220 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.1603
R7221 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.1603
R7222 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1603
R7223 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1603
R7224 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.159278
R7225 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.159278
R7226 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.159278
R7227 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.159278
R7228 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.159278
R7229 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.159278
R7230 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.159278
R7231 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.159278
R7232 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.159278
R7233 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.159278
R7234 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.159278
R7235 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.159278
R7236 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.159278
R7237 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R7238 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R7239 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R7240 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7241 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7242 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7243 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7244 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7245 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7246 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7247 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.159278
R7248 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 0.159278
R7249 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.159278
R7250 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.159278
R7251 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.137822
R7252 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.1368
R7253 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1368
R7254 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1368
R7255 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1368
R7256 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1368
R7257 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.1368
R7258 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1368
R7259 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.1368
R7260 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1368
R7261 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1368
R7262 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1368
R7263 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.1368
R7264 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1368
R7265 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.1368
R7266 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1368
R7267 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.1368
R7268 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1368
R7269 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1368
R7270 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1368
R7271 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R7272 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1368
R7273 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1368
R7274 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.1368
R7275 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.1368
R7276 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1368
R7277 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1368
R7278 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1368
R7279 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1368
R7280 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1368
R7281 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7282 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.1368
R7283 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.114322
R7284 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.1133
R7285 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.1133
R7286 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7287 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7288 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7289 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7290 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7291 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7292 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7293 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7294 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7295 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7296 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7297 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7298 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.1133
R7299 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.1133
R7300 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.1133
R7301 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.1133
R7302 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R7303 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.00152174
R7304 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R7305 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.00152174
R7306 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.00152174
R7307 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.00152174
R7308 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.00152174
R7309 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.00152174
R7310 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.00152174
R7311 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.00152174
R7312 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.00152174
R7313 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.00152174
R7314 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R7315 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.00152174
R7316 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.00152174
R7317 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.00152174
R7318 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.00152174
R7319 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R7320 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.00152174
R7321 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.00152174
R7322 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.00152174
R7323 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R7324 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.00152174
R7325 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.00152174
R7326 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.00152174
R7327 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.00152174
R7328 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.00152174
R7329 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.00152174
R7330 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.00152174
R7331 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.00152174
R7332 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.00152174
R7333 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.00152174
R7334 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.00152174
R7335 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.00152174
R7336 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R7337 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.00152174
R7338 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R7339 ref_volt_cur_gen_dummy_magic_0.Vbe2.n102 ref_volt_cur_gen_dummy_magic_0.Vbe2.t0 162.458
R7340 ref_volt_cur_gen_dummy_magic_0.Vbe2.n117 ref_volt_cur_gen_dummy_magic_0.Vbe2.n116 83.5719
R7341 ref_volt_cur_gen_dummy_magic_0.Vbe2.n115 ref_volt_cur_gen_dummy_magic_0.Vbe2.n9 83.5719
R7342 ref_volt_cur_gen_dummy_magic_0.Vbe2.n114 ref_volt_cur_gen_dummy_magic_0.Vbe2.n113 83.5719
R7343 ref_volt_cur_gen_dummy_magic_0.Vbe2.n105 ref_volt_cur_gen_dummy_magic_0.Vbe2.n12 83.5719
R7344 ref_volt_cur_gen_dummy_magic_0.Vbe2.n97 ref_volt_cur_gen_dummy_magic_0.Vbe2.n13 83.5719
R7345 ref_volt_cur_gen_dummy_magic_0.Vbe2.n99 ref_volt_cur_gen_dummy_magic_0.Vbe2.n98 83.5719
R7346 ref_volt_cur_gen_dummy_magic_0.Vbe2.n91 ref_volt_cur_gen_dummy_magic_0.Vbe2.n17 83.5719
R7347 ref_volt_cur_gen_dummy_magic_0.Vbe2.n81 ref_volt_cur_gen_dummy_magic_0.Vbe2.n80 83.5719
R7348 ref_volt_cur_gen_dummy_magic_0.Vbe2.n79 ref_volt_cur_gen_dummy_magic_0.Vbe2.n78 83.5719
R7349 ref_volt_cur_gen_dummy_magic_0.Vbe2.n77 ref_volt_cur_gen_dummy_magic_0.Vbe2.n76 83.5719
R7350 ref_volt_cur_gen_dummy_magic_0.Vbe2.n38 ref_volt_cur_gen_dummy_magic_0.Vbe2.n37 83.5719
R7351 ref_volt_cur_gen_dummy_magic_0.Vbe2.n36 ref_volt_cur_gen_dummy_magic_0.Vbe2.n34 83.5719
R7352 ref_volt_cur_gen_dummy_magic_0.Vbe2.n44 ref_volt_cur_gen_dummy_magic_0.Vbe2.n33 83.5719
R7353 ref_volt_cur_gen_dummy_magic_0.Vbe2.n52 ref_volt_cur_gen_dummy_magic_0.Vbe2.n51 83.5719
R7354 ref_volt_cur_gen_dummy_magic_0.Vbe2.n31 ref_volt_cur_gen_dummy_magic_0.Vbe2.n29 83.5719
R7355 ref_volt_cur_gen_dummy_magic_0.Vbe2.n57 ref_volt_cur_gen_dummy_magic_0.Vbe2.n28 83.5719
R7356 ref_volt_cur_gen_dummy_magic_0.Vbe2.n65 ref_volt_cur_gen_dummy_magic_0.Vbe2.n64 83.5719
R7357 ref_volt_cur_gen_dummy_magic_0.Vbe2.n130 ref_volt_cur_gen_dummy_magic_0.Vbe2.n0 83.5719
R7358 ref_volt_cur_gen_dummy_magic_0.Vbe2.n132 ref_volt_cur_gen_dummy_magic_0.Vbe2.n131 83.5719
R7359 ref_volt_cur_gen_dummy_magic_0.Vbe2.n134 ref_volt_cur_gen_dummy_magic_0.Vbe2.n133 83.5719
R7360 ref_volt_cur_gen_dummy_magic_0.Vbe2.n116 ref_volt_cur_gen_dummy_magic_0.Vbe2.n8 73.682
R7361 ref_volt_cur_gen_dummy_magic_0.Vbe2.n37 ref_volt_cur_gen_dummy_magic_0.Vbe2.n35 73.682
R7362 ref_volt_cur_gen_dummy_magic_0.Vbe2.n114 ref_volt_cur_gen_dummy_magic_0.Vbe2.n10 73.3165
R7363 ref_volt_cur_gen_dummy_magic_0.Vbe2.n98 ref_volt_cur_gen_dummy_magic_0.Vbe2.n96 73.3165
R7364 ref_volt_cur_gen_dummy_magic_0.Vbe2.n77 ref_volt_cur_gen_dummy_magic_0.Vbe2.n24 73.3165
R7365 ref_volt_cur_gen_dummy_magic_0.Vbe2.n46 ref_volt_cur_gen_dummy_magic_0.Vbe2.n33 73.3165
R7366 ref_volt_cur_gen_dummy_magic_0.Vbe2.n59 ref_volt_cur_gen_dummy_magic_0.Vbe2.n28 73.3165
R7367 ref_volt_cur_gen_dummy_magic_0.Vbe2.n135 ref_volt_cur_gen_dummy_magic_0.Vbe2.n134 73.3165
R7368 ref_volt_cur_gen_dummy_magic_0.Vbe2.n107 ref_volt_cur_gen_dummy_magic_0.Vbe2.n12 73.19
R7369 ref_volt_cur_gen_dummy_magic_0.Vbe2.n93 ref_volt_cur_gen_dummy_magic_0.Vbe2.n17 73.19
R7370 ref_volt_cur_gen_dummy_magic_0.Vbe2.n82 ref_volt_cur_gen_dummy_magic_0.Vbe2.n81 73.19
R7371 ref_volt_cur_gen_dummy_magic_0.Vbe2.n51 ref_volt_cur_gen_dummy_magic_0.Vbe2.n50 73.19
R7372 ref_volt_cur_gen_dummy_magic_0.Vbe2.n64 ref_volt_cur_gen_dummy_magic_0.Vbe2.n63 73.19
R7373 ref_volt_cur_gen_dummy_magic_0.Vbe2.n130 ref_volt_cur_gen_dummy_magic_0.Vbe2.n4 73.19
R7374 ref_volt_cur_gen_dummy_magic_0.Vbe2.n18 ref_volt_cur_gen_dummy_magic_0.Vbe2.t3 36.6632
R7375 ref_volt_cur_gen_dummy_magic_0.Vbe2.t6 ref_volt_cur_gen_dummy_magic_0.Vbe2.n25 36.6632
R7376 ref_volt_cur_gen_dummy_magic_0.Vbe2.n115 ref_volt_cur_gen_dummy_magic_0.Vbe2.n114 26.074
R7377 ref_volt_cur_gen_dummy_magic_0.Vbe2.n98 ref_volt_cur_gen_dummy_magic_0.Vbe2.n97 26.074
R7378 ref_volt_cur_gen_dummy_magic_0.Vbe2.n79 ref_volt_cur_gen_dummy_magic_0.Vbe2.n77 26.074
R7379 ref_volt_cur_gen_dummy_magic_0.Vbe2.n36 ref_volt_cur_gen_dummy_magic_0.Vbe2.n33 26.074
R7380 ref_volt_cur_gen_dummy_magic_0.Vbe2.n31 ref_volt_cur_gen_dummy_magic_0.Vbe2.n28 26.074
R7381 ref_volt_cur_gen_dummy_magic_0.Vbe2.n134 ref_volt_cur_gen_dummy_magic_0.Vbe2.n132 26.074
R7382 ref_volt_cur_gen_dummy_magic_0.Vbe2.n116 ref_volt_cur_gen_dummy_magic_0.Vbe2.t7 25.7843
R7383 ref_volt_cur_gen_dummy_magic_0.Vbe2.t2 ref_volt_cur_gen_dummy_magic_0.Vbe2.n12 25.7843
R7384 ref_volt_cur_gen_dummy_magic_0.Vbe2.t3 ref_volt_cur_gen_dummy_magic_0.Vbe2.n17 25.7843
R7385 ref_volt_cur_gen_dummy_magic_0.Vbe2.n81 ref_volt_cur_gen_dummy_magic_0.Vbe2.t4 25.7843
R7386 ref_volt_cur_gen_dummy_magic_0.Vbe2.n37 ref_volt_cur_gen_dummy_magic_0.Vbe2.t1 25.7843
R7387 ref_volt_cur_gen_dummy_magic_0.Vbe2.n51 ref_volt_cur_gen_dummy_magic_0.Vbe2.t5 25.7843
R7388 ref_volt_cur_gen_dummy_magic_0.Vbe2.n64 ref_volt_cur_gen_dummy_magic_0.Vbe2.t6 25.7843
R7389 ref_volt_cur_gen_dummy_magic_0.Vbe2.t8 ref_volt_cur_gen_dummy_magic_0.Vbe2.n130 25.7843
R7390 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n3 9.3005
R7391 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 ref_volt_cur_gen_dummy_magic_0.Vbe2.n3 9.3005
R7392 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 ref_volt_cur_gen_dummy_magic_0.Vbe2.n3 9.3005
R7393 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 ref_volt_cur_gen_dummy_magic_0.Vbe2.n3 9.3005
R7394 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n5 9.3005
R7395 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 ref_volt_cur_gen_dummy_magic_0.Vbe2.n5 9.3005
R7396 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 ref_volt_cur_gen_dummy_magic_0.Vbe2.n5 9.3005
R7397 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 ref_volt_cur_gen_dummy_magic_0.Vbe2.n5 9.3005
R7398 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n2 9.3005
R7399 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 ref_volt_cur_gen_dummy_magic_0.Vbe2.n2 9.3005
R7400 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 ref_volt_cur_gen_dummy_magic_0.Vbe2.n2 9.3005
R7401 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 ref_volt_cur_gen_dummy_magic_0.Vbe2.n2 9.3005
R7402 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n6 9.3005
R7403 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 ref_volt_cur_gen_dummy_magic_0.Vbe2.n6 9.3005
R7404 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 ref_volt_cur_gen_dummy_magic_0.Vbe2.n6 9.3005
R7405 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 ref_volt_cur_gen_dummy_magic_0.Vbe2.n6 9.3005
R7406 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 9.3005
R7407 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 9.3005
R7408 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 9.3005
R7409 ref_volt_cur_gen_dummy_magic_0.Vbe2.n123 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 9.3005
R7410 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 9.3005
R7411 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 9.3005
R7412 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 9.3005
R7413 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 9.3005
R7414 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 ref_volt_cur_gen_dummy_magic_0.Vbe2.n123 9.3005
R7415 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 9.3005
R7416 ref_volt_cur_gen_dummy_magic_0.Vbe2.n71 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 9.3005
R7417 ref_volt_cur_gen_dummy_magic_0.Vbe2.n71 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 9.3005
R7418 ref_volt_cur_gen_dummy_magic_0.Vbe2.n71 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 9.3005
R7419 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 ref_volt_cur_gen_dummy_magic_0.Vbe2.n71 9.3005
R7420 ref_volt_cur_gen_dummy_magic_0.Vbe2.n73 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 9.3005
R7421 ref_volt_cur_gen_dummy_magic_0.Vbe2.n73 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 9.3005
R7422 ref_volt_cur_gen_dummy_magic_0.Vbe2.n73 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 9.3005
R7423 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 ref_volt_cur_gen_dummy_magic_0.Vbe2.n73 9.3005
R7424 ref_volt_cur_gen_dummy_magic_0.Vbe2.n70 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 9.3005
R7425 ref_volt_cur_gen_dummy_magic_0.Vbe2.n70 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 9.3005
R7426 ref_volt_cur_gen_dummy_magic_0.Vbe2.n70 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 9.3005
R7427 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 ref_volt_cur_gen_dummy_magic_0.Vbe2.n70 9.3005
R7428 ref_volt_cur_gen_dummy_magic_0.Vbe2.n85 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 9.3005
R7429 ref_volt_cur_gen_dummy_magic_0.Vbe2.n85 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 9.3005
R7430 ref_volt_cur_gen_dummy_magic_0.Vbe2.n85 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 9.3005
R7431 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 ref_volt_cur_gen_dummy_magic_0.Vbe2.n85 9.3005
R7432 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 9.3005
R7433 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 9.3005
R7434 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 9.3005
R7435 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 ref_volt_cur_gen_dummy_magic_0.Vbe2.n19 9.3005
R7436 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 9.3005
R7437 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 9.3005
R7438 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 9.3005
R7439 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 9.3005
R7440 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 ref_volt_cur_gen_dummy_magic_0.Vbe2.n19 9.3005
R7441 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 9.3005
R7442 ref_volt_cur_gen_dummy_magic_0.Vbe2.n123 ref_volt_cur_gen_dummy_magic_0.Vbe2.n121 4.64654
R7443 ref_volt_cur_gen_dummy_magic_0.Vbe2.n127 ref_volt_cur_gen_dummy_magic_0.Vbe2.n126 4.64654
R7444 ref_volt_cur_gen_dummy_magic_0.Vbe2.n123 ref_volt_cur_gen_dummy_magic_0.Vbe2.n122 4.64654
R7445 ref_volt_cur_gen_dummy_magic_0.Vbe2.n127 ref_volt_cur_gen_dummy_magic_0.Vbe2.n125 4.64654
R7446 ref_volt_cur_gen_dummy_magic_0.Vbe2.n128 ref_volt_cur_gen_dummy_magic_0.Vbe2.n127 4.64654
R7447 ref_volt_cur_gen_dummy_magic_0.Vbe2.n72 ref_volt_cur_gen_dummy_magic_0.Vbe2.n19 4.64654
R7448 ref_volt_cur_gen_dummy_magic_0.Vbe2.n83 ref_volt_cur_gen_dummy_magic_0.Vbe2.n75 4.64654
R7449 ref_volt_cur_gen_dummy_magic_0.Vbe2.n74 ref_volt_cur_gen_dummy_magic_0.Vbe2.n19 4.64654
R7450 ref_volt_cur_gen_dummy_magic_0.Vbe2.n84 ref_volt_cur_gen_dummy_magic_0.Vbe2.n83 4.64654
R7451 ref_volt_cur_gen_dummy_magic_0.Vbe2.n83 ref_volt_cur_gen_dummy_magic_0.Vbe2.n21 4.64654
R7452 ref_volt_cur_gen_dummy_magic_0.Vbe2.n108 ref_volt_cur_gen_dummy_magic_0.Vbe2.n107 2.36206
R7453 ref_volt_cur_gen_dummy_magic_0.Vbe2.n94 ref_volt_cur_gen_dummy_magic_0.Vbe2.n93 2.36206
R7454 ref_volt_cur_gen_dummy_magic_0.Vbe2.n50 ref_volt_cur_gen_dummy_magic_0.Vbe2.n48 2.36206
R7455 ref_volt_cur_gen_dummy_magic_0.Vbe2.n63 ref_volt_cur_gen_dummy_magic_0.Vbe2.n61 2.36206
R7456 ref_volt_cur_gen_dummy_magic_0.Vbe2.n109 ref_volt_cur_gen_dummy_magic_0.Vbe2.n10 2.19742
R7457 ref_volt_cur_gen_dummy_magic_0.Vbe2.n96 ref_volt_cur_gen_dummy_magic_0.Vbe2.n95 2.19742
R7458 ref_volt_cur_gen_dummy_magic_0.Vbe2.n47 ref_volt_cur_gen_dummy_magic_0.Vbe2.n46 2.19742
R7459 ref_volt_cur_gen_dummy_magic_0.Vbe2.n60 ref_volt_cur_gen_dummy_magic_0.Vbe2.n59 2.19742
R7460 ref_volt_cur_gen_dummy_magic_0.Vbe2.n90 ref_volt_cur_gen_dummy_magic_0.Vbe2.n18 1.80777
R7461 ref_volt_cur_gen_dummy_magic_0.Vbe2.n66 ref_volt_cur_gen_dummy_magic_0.Vbe2.n25 1.80777
R7462 ref_volt_cur_gen_dummy_magic_0.Vbe2.n62 ref_volt_cur_gen_dummy_magic_0.Vbe2.n26 1.5505
R7463 ref_volt_cur_gen_dummy_magic_0.Vbe2.n67 ref_volt_cur_gen_dummy_magic_0.Vbe2.n66 1.5505
R7464 ref_volt_cur_gen_dummy_magic_0.Vbe2.n49 ref_volt_cur_gen_dummy_magic_0.Vbe2.n30 1.5505
R7465 ref_volt_cur_gen_dummy_magic_0.Vbe2.n54 ref_volt_cur_gen_dummy_magic_0.Vbe2.n53 1.5505
R7466 ref_volt_cur_gen_dummy_magic_0.Vbe2.n56 ref_volt_cur_gen_dummy_magic_0.Vbe2.n55 1.5505
R7467 ref_volt_cur_gen_dummy_magic_0.Vbe2.n58 ref_volt_cur_gen_dummy_magic_0.Vbe2.n27 1.5505
R7468 ref_volt_cur_gen_dummy_magic_0.Vbe2.n40 ref_volt_cur_gen_dummy_magic_0.Vbe2.n39 1.5505
R7469 ref_volt_cur_gen_dummy_magic_0.Vbe2.n43 ref_volt_cur_gen_dummy_magic_0.Vbe2.n42 1.5505
R7470 ref_volt_cur_gen_dummy_magic_0.Vbe2.n45 ref_volt_cur_gen_dummy_magic_0.Vbe2.n32 1.5505
R7471 ref_volt_cur_gen_dummy_magic_0.Vbe2.n92 ref_volt_cur_gen_dummy_magic_0.Vbe2.n16 1.5505
R7472 ref_volt_cur_gen_dummy_magic_0.Vbe2.n90 ref_volt_cur_gen_dummy_magic_0.Vbe2.n89 1.5505
R7473 ref_volt_cur_gen_dummy_magic_0.Vbe2.n106 ref_volt_cur_gen_dummy_magic_0.Vbe2.n11 1.5505
R7474 ref_volt_cur_gen_dummy_magic_0.Vbe2.n104 ref_volt_cur_gen_dummy_magic_0.Vbe2.n103 1.5505
R7475 ref_volt_cur_gen_dummy_magic_0.Vbe2.n101 ref_volt_cur_gen_dummy_magic_0.Vbe2.n100 1.5505
R7476 ref_volt_cur_gen_dummy_magic_0.Vbe2.n15 ref_volt_cur_gen_dummy_magic_0.Vbe2.n14 1.5505
R7477 ref_volt_cur_gen_dummy_magic_0.Vbe2.n119 ref_volt_cur_gen_dummy_magic_0.Vbe2.n118 1.5505
R7478 ref_volt_cur_gen_dummy_magic_0.Vbe2.n112 ref_volt_cur_gen_dummy_magic_0.Vbe2.n7 1.5505
R7479 ref_volt_cur_gen_dummy_magic_0.Vbe2.n111 ref_volt_cur_gen_dummy_magic_0.Vbe2.n110 1.5505
R7480 ref_volt_cur_gen_dummy_magic_0.Vbe2.n111 ref_volt_cur_gen_dummy_magic_0.Vbe2.n10 1.19225
R7481 ref_volt_cur_gen_dummy_magic_0.Vbe2.n96 ref_volt_cur_gen_dummy_magic_0.Vbe2.n15 1.19225
R7482 ref_volt_cur_gen_dummy_magic_0.Vbe2.n24 ref_volt_cur_gen_dummy_magic_0.Vbe2.n19 1.19225
R7483 ref_volt_cur_gen_dummy_magic_0.Vbe2.n46 ref_volt_cur_gen_dummy_magic_0.Vbe2.n45 1.19225
R7484 ref_volt_cur_gen_dummy_magic_0.Vbe2.n59 ref_volt_cur_gen_dummy_magic_0.Vbe2.n58 1.19225
R7485 ref_volt_cur_gen_dummy_magic_0.Vbe2.n135 ref_volt_cur_gen_dummy_magic_0.Vbe2.n123 1.19225
R7486 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n8 1.07742
R7487 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n35 1.07742
R7488 ref_volt_cur_gen_dummy_magic_0.Vbe2.n118 ref_volt_cur_gen_dummy_magic_0.Vbe2.n9 1.07024
R7489 ref_volt_cur_gen_dummy_magic_0.Vbe2.n104 ref_volt_cur_gen_dummy_magic_0.Vbe2.n13 1.07024
R7490 ref_volt_cur_gen_dummy_magic_0.Vbe2.n78 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 1.07024
R7491 ref_volt_cur_gen_dummy_magic_0.Vbe2.n39 ref_volt_cur_gen_dummy_magic_0.Vbe2.n34 1.07024
R7492 ref_volt_cur_gen_dummy_magic_0.Vbe2.n53 ref_volt_cur_gen_dummy_magic_0.Vbe2.n29 1.07024
R7493 ref_volt_cur_gen_dummy_magic_0.Vbe2.n131 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 1.07024
R7494 ref_volt_cur_gen_dummy_magic_0.Vbe2.n68 ref_volt_cur_gen_dummy_magic_0.Vbe2.n25 1.04793
R7495 ref_volt_cur_gen_dummy_magic_0.Vbe2.n88 ref_volt_cur_gen_dummy_magic_0.Vbe2.n18 1.04793
R7496 ref_volt_cur_gen_dummy_magic_0.Vbe2.n107 ref_volt_cur_gen_dummy_magic_0.Vbe2.n106 1.0237
R7497 ref_volt_cur_gen_dummy_magic_0.Vbe2.n93 ref_volt_cur_gen_dummy_magic_0.Vbe2.n92 1.0237
R7498 ref_volt_cur_gen_dummy_magic_0.Vbe2.n82 ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 1.0237
R7499 ref_volt_cur_gen_dummy_magic_0.Vbe2.n50 ref_volt_cur_gen_dummy_magic_0.Vbe2.n49 1.0237
R7500 ref_volt_cur_gen_dummy_magic_0.Vbe2.n63 ref_volt_cur_gen_dummy_magic_0.Vbe2.n62 1.0237
R7501 ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 ref_volt_cur_gen_dummy_magic_0.Vbe2.n4 1.0237
R7502 ref_volt_cur_gen_dummy_magic_0.Vbe2.n113 ref_volt_cur_gen_dummy_magic_0.Vbe2.n111 0.959578
R7503 ref_volt_cur_gen_dummy_magic_0.Vbe2.n99 ref_volt_cur_gen_dummy_magic_0.Vbe2.n15 0.959578
R7504 ref_volt_cur_gen_dummy_magic_0.Vbe2.n76 ref_volt_cur_gen_dummy_magic_0.Vbe2.n19 0.959578
R7505 ref_volt_cur_gen_dummy_magic_0.Vbe2.n45 ref_volt_cur_gen_dummy_magic_0.Vbe2.n44 0.959578
R7506 ref_volt_cur_gen_dummy_magic_0.Vbe2.n58 ref_volt_cur_gen_dummy_magic_0.Vbe2.n57 0.959578
R7507 ref_volt_cur_gen_dummy_magic_0.Vbe2.n133 ref_volt_cur_gen_dummy_magic_0.Vbe2.n123 0.959578
R7508 ref_volt_cur_gen_dummy_magic_0.Vbe2.n113 ref_volt_cur_gen_dummy_magic_0.Vbe2.n112 0.885803
R7509 ref_volt_cur_gen_dummy_magic_0.Vbe2.n100 ref_volt_cur_gen_dummy_magic_0.Vbe2.n99 0.885803
R7510 ref_volt_cur_gen_dummy_magic_0.Vbe2.n76 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 0.885803
R7511 ref_volt_cur_gen_dummy_magic_0.Vbe2.n44 ref_volt_cur_gen_dummy_magic_0.Vbe2.n43 0.885803
R7512 ref_volt_cur_gen_dummy_magic_0.Vbe2.n57 ref_volt_cur_gen_dummy_magic_0.Vbe2.n56 0.885803
R7513 ref_volt_cur_gen_dummy_magic_0.Vbe2.n133 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 0.885803
R7514 ref_volt_cur_gen_dummy_magic_0.Vbe2.n83 ref_volt_cur_gen_dummy_magic_0.Vbe2.n82 0.812055
R7515 ref_volt_cur_gen_dummy_magic_0.Vbe2.n127 ref_volt_cur_gen_dummy_magic_0.Vbe2.n4 0.812055
R7516 ref_volt_cur_gen_dummy_magic_0.Vbe2.n112 ref_volt_cur_gen_dummy_magic_0.Vbe2.n9 0.77514
R7517 ref_volt_cur_gen_dummy_magic_0.Vbe2.n100 ref_volt_cur_gen_dummy_magic_0.Vbe2.n13 0.77514
R7518 ref_volt_cur_gen_dummy_magic_0.Vbe2.n78 ref_volt_cur_gen_dummy_magic_0.Vbe2.n23 0.77514
R7519 ref_volt_cur_gen_dummy_magic_0.Vbe2.n43 ref_volt_cur_gen_dummy_magic_0.Vbe2.n34 0.77514
R7520 ref_volt_cur_gen_dummy_magic_0.Vbe2.n56 ref_volt_cur_gen_dummy_magic_0.Vbe2.n29 0.77514
R7521 ref_volt_cur_gen_dummy_magic_0.Vbe2.n131 ref_volt_cur_gen_dummy_magic_0.Vbe2.n129 0.77514
R7522 ref_volt_cur_gen_dummy_magic_0.Vbe2.n40 ref_volt_cur_gen_dummy_magic_0.Vbe2.n35 0.763532
R7523 ref_volt_cur_gen_dummy_magic_0.Vbe2.n119 ref_volt_cur_gen_dummy_magic_0.Vbe2.n8 0.763532
R7524 ref_volt_cur_gen_dummy_magic_0.Vbe2.n106 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16.Emitter 0.756696
R7525 ref_volt_cur_gen_dummy_magic_0.Vbe2.n92 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11.Emitter 0.756696
R7526 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n22 0.756696
R7527 ref_volt_cur_gen_dummy_magic_0.Vbe2.n49 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15.Emitter 0.756696
R7528 ref_volt_cur_gen_dummy_magic_0.Vbe2.n62 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10.Emitter 0.756696
R7529 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n138 0.756696
R7530 ref_volt_cur_gen_dummy_magic_0.Vbe2.n86 ref_volt_cur_gen_dummy_magic_0.Vbe2.n24 0.647417
R7531 ref_volt_cur_gen_dummy_magic_0.Vbe2.n136 ref_volt_cur_gen_dummy_magic_0.Vbe2.n135 0.647417
R7532 ref_volt_cur_gen_dummy_magic_0.Vbe2.n118 ref_volt_cur_gen_dummy_magic_0.Vbe2.n117 0.590702
R7533 ref_volt_cur_gen_dummy_magic_0.Vbe2.n105 ref_volt_cur_gen_dummy_magic_0.Vbe2.n104 0.590702
R7534 ref_volt_cur_gen_dummy_magic_0.Vbe2.n91 ref_volt_cur_gen_dummy_magic_0.Vbe2.n90 0.590702
R7535 ref_volt_cur_gen_dummy_magic_0.Vbe2.n80 ref_volt_cur_gen_dummy_magic_0.Vbe2.n20 0.590702
R7536 ref_volt_cur_gen_dummy_magic_0.Vbe2.n39 ref_volt_cur_gen_dummy_magic_0.Vbe2.n38 0.590702
R7537 ref_volt_cur_gen_dummy_magic_0.Vbe2.n53 ref_volt_cur_gen_dummy_magic_0.Vbe2.n52 0.590702
R7538 ref_volt_cur_gen_dummy_magic_0.Vbe2.n66 ref_volt_cur_gen_dummy_magic_0.Vbe2.n65 0.590702
R7539 ref_volt_cur_gen_dummy_magic_0.Vbe2.n124 ref_volt_cur_gen_dummy_magic_0.Vbe2.n0 0.590702
R7540 ref_volt_cur_gen_dummy_magic_0.Vbe2.n117 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14.Emitter 0.498483
R7541 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n105 0.498483
R7542 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n91 0.498483
R7543 ref_volt_cur_gen_dummy_magic_0.Vbe2.n80 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9.Emitter 0.498483
R7544 ref_volt_cur_gen_dummy_magic_0.Vbe2.n38 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12.Emitter 0.498483
R7545 ref_volt_cur_gen_dummy_magic_0.Vbe2.n52 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15.Emitter 0.498483
R7546 ref_volt_cur_gen_dummy_magic_0.Vbe2.n65 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10.Emitter 0.498483
R7547 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13.Emitter ref_volt_cur_gen_dummy_magic_0.Vbe2.n0 0.498483
R7548 ref_volt_cur_gen_dummy_magic_0.Vbe2.t7 ref_volt_cur_gen_dummy_magic_0.Vbe2.n115 0.290206
R7549 ref_volt_cur_gen_dummy_magic_0.Vbe2.n97 ref_volt_cur_gen_dummy_magic_0.Vbe2.t2 0.290206
R7550 ref_volt_cur_gen_dummy_magic_0.Vbe2.t4 ref_volt_cur_gen_dummy_magic_0.Vbe2.n79 0.290206
R7551 ref_volt_cur_gen_dummy_magic_0.Vbe2.t1 ref_volt_cur_gen_dummy_magic_0.Vbe2.n36 0.290206
R7552 ref_volt_cur_gen_dummy_magic_0.Vbe2.t5 ref_volt_cur_gen_dummy_magic_0.Vbe2.n31 0.290206
R7553 ref_volt_cur_gen_dummy_magic_0.Vbe2.n132 ref_volt_cur_gen_dummy_magic_0.Vbe2.t8 0.290206
R7554 ref_volt_cur_gen_dummy_magic_0.Vbe2.n61 ref_volt_cur_gen_dummy_magic_0.Vbe2.n60 0.154071
R7555 ref_volt_cur_gen_dummy_magic_0.Vbe2.n48 ref_volt_cur_gen_dummy_magic_0.Vbe2.n47 0.154071
R7556 ref_volt_cur_gen_dummy_magic_0.Vbe2.n95 ref_volt_cur_gen_dummy_magic_0.Vbe2.n94 0.154071
R7557 ref_volt_cur_gen_dummy_magic_0.Vbe2.n109 ref_volt_cur_gen_dummy_magic_0.Vbe2.n108 0.154071
R7558 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 ref_volt_cur_gen_dummy_magic_0.Vbe2.n120 0.137464
R7559 ref_volt_cur_gen_dummy_magic_0.Vbe2.n88 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 0.137464
R7560 ref_volt_cur_gen_dummy_magic_0.Vbe2.n41 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 0.134964
R7561 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 ref_volt_cur_gen_dummy_magic_0.Vbe2.n68 0.134964
R7562 ref_volt_cur_gen_dummy_magic_0.Vbe2.n67 ref_volt_cur_gen_dummy_magic_0.Vbe2.n26 0.0183571
R7563 ref_volt_cur_gen_dummy_magic_0.Vbe2.n61 ref_volt_cur_gen_dummy_magic_0.Vbe2.n26 0.0183571
R7564 ref_volt_cur_gen_dummy_magic_0.Vbe2.n60 ref_volt_cur_gen_dummy_magic_0.Vbe2.n27 0.0183571
R7565 ref_volt_cur_gen_dummy_magic_0.Vbe2.n55 ref_volt_cur_gen_dummy_magic_0.Vbe2.n27 0.0183571
R7566 ref_volt_cur_gen_dummy_magic_0.Vbe2.n55 ref_volt_cur_gen_dummy_magic_0.Vbe2.n54 0.0183571
R7567 ref_volt_cur_gen_dummy_magic_0.Vbe2.n54 ref_volt_cur_gen_dummy_magic_0.Vbe2.n30 0.0183571
R7568 ref_volt_cur_gen_dummy_magic_0.Vbe2.n48 ref_volt_cur_gen_dummy_magic_0.Vbe2.n30 0.0183571
R7569 ref_volt_cur_gen_dummy_magic_0.Vbe2.n47 ref_volt_cur_gen_dummy_magic_0.Vbe2.n32 0.0183571
R7570 ref_volt_cur_gen_dummy_magic_0.Vbe2.n42 ref_volt_cur_gen_dummy_magic_0.Vbe2.n32 0.0183571
R7571 ref_volt_cur_gen_dummy_magic_0.Vbe2.n89 ref_volt_cur_gen_dummy_magic_0.Vbe2.n16 0.0183571
R7572 ref_volt_cur_gen_dummy_magic_0.Vbe2.n94 ref_volt_cur_gen_dummy_magic_0.Vbe2.n16 0.0183571
R7573 ref_volt_cur_gen_dummy_magic_0.Vbe2.n95 ref_volt_cur_gen_dummy_magic_0.Vbe2.n14 0.0183571
R7574 ref_volt_cur_gen_dummy_magic_0.Vbe2.n101 ref_volt_cur_gen_dummy_magic_0.Vbe2.n14 0.0183571
R7575 ref_volt_cur_gen_dummy_magic_0.Vbe2.n103 ref_volt_cur_gen_dummy_magic_0.Vbe2.n11 0.0183571
R7576 ref_volt_cur_gen_dummy_magic_0.Vbe2.n108 ref_volt_cur_gen_dummy_magic_0.Vbe2.n11 0.0183571
R7577 ref_volt_cur_gen_dummy_magic_0.Vbe2.n110 ref_volt_cur_gen_dummy_magic_0.Vbe2.n109 0.0183571
R7578 ref_volt_cur_gen_dummy_magic_0.Vbe2.n110 ref_volt_cur_gen_dummy_magic_0.Vbe2.n7 0.0183571
R7579 ref_volt_cur_gen_dummy_magic_0.Vbe2.n68 ref_volt_cur_gen_dummy_magic_0.Vbe2.n67 0.0106786
R7580 ref_volt_cur_gen_dummy_magic_0.Vbe2.n41 ref_volt_cur_gen_dummy_magic_0.Vbe2.n40 0.0106786
R7581 ref_volt_cur_gen_dummy_magic_0.Vbe2.n89 ref_volt_cur_gen_dummy_magic_0.Vbe2.n88 0.0106786
R7582 ref_volt_cur_gen_dummy_magic_0.Vbe2.n120 ref_volt_cur_gen_dummy_magic_0.Vbe2.n119 0.0106786
R7583 ref_volt_cur_gen_dummy_magic_0.Vbe2.n102 ref_volt_cur_gen_dummy_magic_0.Vbe2.n101 0.00996429
R7584 ref_volt_cur_gen_dummy_magic_0.Vbe2.n137 ref_volt_cur_gen_dummy_magic_0.Vbe2.n128 0.00992001
R7585 ref_volt_cur_gen_dummy_magic_0.Vbe2.n121 ref_volt_cur_gen_dummy_magic_0.Vbe2.n5 0.00992001
R7586 ref_volt_cur_gen_dummy_magic_0.Vbe2.n126 ref_volt_cur_gen_dummy_magic_0.Vbe2.n2 0.00992001
R7587 ref_volt_cur_gen_dummy_magic_0.Vbe2.n122 ref_volt_cur_gen_dummy_magic_0.Vbe2.n6 0.00992001
R7588 ref_volt_cur_gen_dummy_magic_0.Vbe2.n125 ref_volt_cur_gen_dummy_magic_0.Vbe2.n1 0.00992001
R7589 ref_volt_cur_gen_dummy_magic_0.Vbe2.n128 ref_volt_cur_gen_dummy_magic_0.Vbe2.n3 0.00992001
R7590 ref_volt_cur_gen_dummy_magic_0.Vbe2.n121 ref_volt_cur_gen_dummy_magic_0.Vbe2.n3 0.00992001
R7591 ref_volt_cur_gen_dummy_magic_0.Vbe2.n126 ref_volt_cur_gen_dummy_magic_0.Vbe2.n5 0.00992001
R7592 ref_volt_cur_gen_dummy_magic_0.Vbe2.n122 ref_volt_cur_gen_dummy_magic_0.Vbe2.n2 0.00992001
R7593 ref_volt_cur_gen_dummy_magic_0.Vbe2.n125 ref_volt_cur_gen_dummy_magic_0.Vbe2.n6 0.00992001
R7594 ref_volt_cur_gen_dummy_magic_0.Vbe2.n87 ref_volt_cur_gen_dummy_magic_0.Vbe2.n21 0.00992001
R7595 ref_volt_cur_gen_dummy_magic_0.Vbe2.n73 ref_volt_cur_gen_dummy_magic_0.Vbe2.n72 0.00992001
R7596 ref_volt_cur_gen_dummy_magic_0.Vbe2.n75 ref_volt_cur_gen_dummy_magic_0.Vbe2.n70 0.00992001
R7597 ref_volt_cur_gen_dummy_magic_0.Vbe2.n85 ref_volt_cur_gen_dummy_magic_0.Vbe2.n74 0.00992001
R7598 ref_volt_cur_gen_dummy_magic_0.Vbe2.n84 ref_volt_cur_gen_dummy_magic_0.Vbe2.n69 0.00992001
R7599 ref_volt_cur_gen_dummy_magic_0.Vbe2.n71 ref_volt_cur_gen_dummy_magic_0.Vbe2.n21 0.00992001
R7600 ref_volt_cur_gen_dummy_magic_0.Vbe2.n72 ref_volt_cur_gen_dummy_magic_0.Vbe2.n71 0.00992001
R7601 ref_volt_cur_gen_dummy_magic_0.Vbe2.n75 ref_volt_cur_gen_dummy_magic_0.Vbe2.n73 0.00992001
R7602 ref_volt_cur_gen_dummy_magic_0.Vbe2.n74 ref_volt_cur_gen_dummy_magic_0.Vbe2.n70 0.00992001
R7603 ref_volt_cur_gen_dummy_magic_0.Vbe2.n85 ref_volt_cur_gen_dummy_magic_0.Vbe2.n84 0.00992001
R7604 ref_volt_cur_gen_dummy_magic_0.Vbe2.n103 ref_volt_cur_gen_dummy_magic_0.Vbe2.n102 0.00889286
R7605 ref_volt_cur_gen_dummy_magic_0.Vbe2.n42 ref_volt_cur_gen_dummy_magic_0.Vbe2.n41 0.00817857
R7606 ref_volt_cur_gen_dummy_magic_0.Vbe2.n120 ref_volt_cur_gen_dummy_magic_0.Vbe2.n7 0.00817857
R7607 ref_volt_cur_gen_dummy_magic_0.START_UP.n1 ref_volt_cur_gen_dummy_magic_0.START_UP.t7 238.322
R7608 ref_volt_cur_gen_dummy_magic_0.START_UP.n1 ref_volt_cur_gen_dummy_magic_0.START_UP.t6 238.322
R7609 ref_volt_cur_gen_dummy_magic_0.START_UP.n5 ref_volt_cur_gen_dummy_magic_0.START_UP.n4 175.558
R7610 ref_volt_cur_gen_dummy_magic_0.START_UP.n4 ref_volt_cur_gen_dummy_magic_0.START_UP.n3 168.935
R7611 ref_volt_cur_gen_dummy_magic_0.START_UP.n2 ref_volt_cur_gen_dummy_magic_0.START_UP.n1 166.925
R7612 ref_volt_cur_gen_dummy_magic_0.START_UP.n0 ref_volt_cur_gen_dummy_magic_0.START_UP.t1 130.001
R7613 ref_volt_cur_gen_dummy_magic_0.START_UP.n0 ref_volt_cur_gen_dummy_magic_0.START_UP.t0 81.7084
R7614 ref_volt_cur_gen_dummy_magic_0.START_UP.n2 ref_volt_cur_gen_dummy_magic_0.START_UP.n0 53.0427
R7615 ref_volt_cur_gen_dummy_magic_0.START_UP.n3 ref_volt_cur_gen_dummy_magic_0.START_UP.t3 13.1338
R7616 ref_volt_cur_gen_dummy_magic_0.START_UP.n3 ref_volt_cur_gen_dummy_magic_0.START_UP.t2 13.1338
R7617 ref_volt_cur_gen_dummy_magic_0.START_UP.t5 ref_volt_cur_gen_dummy_magic_0.START_UP.n5 13.1338
R7618 ref_volt_cur_gen_dummy_magic_0.START_UP.n5 ref_volt_cur_gen_dummy_magic_0.START_UP.t4 13.1338
R7619 ref_volt_cur_gen_dummy_magic_0.START_UP.n4 ref_volt_cur_gen_dummy_magic_0.START_UP.n2 4.21925
R7620 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 525.38
R7621 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 525.38
R7622 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 366.856
R7623 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 366.856
R7624 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7625 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 281.168
R7626 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 281.168
R7627 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 281.168
R7628 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7629 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7630 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7631 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7632 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7633 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7634 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7635 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7636 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 39.5005
R7637 a_5750_2946.t0 a_5750_2946.t1 169.905
R7638 ref_volt_cur_gen_dummy_magic_0.Vin+.n3 ref_volt_cur_gen_dummy_magic_0.Vin+.n2 526.183
R7639 ref_volt_cur_gen_dummy_magic_0.Vin+.n1 ref_volt_cur_gen_dummy_magic_0.Vin+.n0 514.134
R7640 ref_volt_cur_gen_dummy_magic_0.Vin+.n0 ref_volt_cur_gen_dummy_magic_0.Vin+.t9 303.259
R7641 ref_volt_cur_gen_dummy_magic_0.Vin+.n7 ref_volt_cur_gen_dummy_magic_0.Vin+.n3 215.732
R7642 ref_volt_cur_gen_dummy_magic_0.Vin+.n0 ref_volt_cur_gen_dummy_magic_0.Vin+.t8 174.726
R7643 ref_volt_cur_gen_dummy_magic_0.Vin+.n1 ref_volt_cur_gen_dummy_magic_0.Vin+.t6 174.726
R7644 ref_volt_cur_gen_dummy_magic_0.Vin+.n2 ref_volt_cur_gen_dummy_magic_0.Vin+.t7 174.726
R7645 ref_volt_cur_gen_dummy_magic_0.Vin+.n6 ref_volt_cur_gen_dummy_magic_0.Vin+.n4 170.56
R7646 ref_volt_cur_gen_dummy_magic_0.Vin+.n6 ref_volt_cur_gen_dummy_magic_0.Vin+.n5 168.435
R7647 ref_volt_cur_gen_dummy_magic_0.Vin+.t0 ref_volt_cur_gen_dummy_magic_0.Vin+.n8 158.796
R7648 ref_volt_cur_gen_dummy_magic_0.Vin+.n8 ref_volt_cur_gen_dummy_magic_0.Vin+.t5 147.981
R7649 ref_volt_cur_gen_dummy_magic_0.Vin+.n2 ref_volt_cur_gen_dummy_magic_0.Vin+.n1 128.534
R7650 ref_volt_cur_gen_dummy_magic_0.Vin+.n3 ref_volt_cur_gen_dummy_magic_0.Vin+.t10 96.4005
R7651 ref_volt_cur_gen_dummy_magic_0.Vin+.n7 ref_volt_cur_gen_dummy_magic_0.Vin+.n6 13.5005
R7652 ref_volt_cur_gen_dummy_magic_0.Vin+.n5 ref_volt_cur_gen_dummy_magic_0.Vin+.t2 13.1338
R7653 ref_volt_cur_gen_dummy_magic_0.Vin+.n5 ref_volt_cur_gen_dummy_magic_0.Vin+.t1 13.1338
R7654 ref_volt_cur_gen_dummy_magic_0.Vin+.n4 ref_volt_cur_gen_dummy_magic_0.Vin+.t4 13.1338
R7655 ref_volt_cur_gen_dummy_magic_0.Vin+.n4 ref_volt_cur_gen_dummy_magic_0.Vin+.t3 13.1338
R7656 ref_volt_cur_gen_dummy_magic_0.Vin+.n8 ref_volt_cur_gen_dummy_magic_0.Vin+.n7 1.438
R7657 ref_volt_cur_gen_dummy_magic_0.V_p_1.n1 ref_volt_cur_gen_dummy_magic_0.V_p_1.n2 229.562
R7658 ref_volt_cur_gen_dummy_magic_0.V_p_1.n0 ref_volt_cur_gen_dummy_magic_0.V_p_1.n5 228.939
R7659 ref_volt_cur_gen_dummy_magic_0.V_p_1.n0 ref_volt_cur_gen_dummy_magic_0.V_p_1.n4 228.939
R7660 ref_volt_cur_gen_dummy_magic_0.V_p_1.n1 ref_volt_cur_gen_dummy_magic_0.V_p_1.n3 228.939
R7661 ref_volt_cur_gen_dummy_magic_0.V_p_1.n6 ref_volt_cur_gen_dummy_magic_0.V_p_1.n1 228.938
R7662 ref_volt_cur_gen_dummy_magic_0.V_p_1.n0 ref_volt_cur_gen_dummy_magic_0.V_p_1.t1 98.2282
R7663 ref_volt_cur_gen_dummy_magic_0.V_p_1.n5 ref_volt_cur_gen_dummy_magic_0.V_p_1.t6 48.0005
R7664 ref_volt_cur_gen_dummy_magic_0.V_p_1.n5 ref_volt_cur_gen_dummy_magic_0.V_p_1.t10 48.0005
R7665 ref_volt_cur_gen_dummy_magic_0.V_p_1.n4 ref_volt_cur_gen_dummy_magic_0.V_p_1.t0 48.0005
R7666 ref_volt_cur_gen_dummy_magic_0.V_p_1.n4 ref_volt_cur_gen_dummy_magic_0.V_p_1.t3 48.0005
R7667 ref_volt_cur_gen_dummy_magic_0.V_p_1.n3 ref_volt_cur_gen_dummy_magic_0.V_p_1.t5 48.0005
R7668 ref_volt_cur_gen_dummy_magic_0.V_p_1.n3 ref_volt_cur_gen_dummy_magic_0.V_p_1.t2 48.0005
R7669 ref_volt_cur_gen_dummy_magic_0.V_p_1.n2 ref_volt_cur_gen_dummy_magic_0.V_p_1.t9 48.0005
R7670 ref_volt_cur_gen_dummy_magic_0.V_p_1.n2 ref_volt_cur_gen_dummy_magic_0.V_p_1.t4 48.0005
R7671 ref_volt_cur_gen_dummy_magic_0.V_p_1.n6 ref_volt_cur_gen_dummy_magic_0.V_p_1.t8 48.0005
R7672 ref_volt_cur_gen_dummy_magic_0.V_p_1.t7 ref_volt_cur_gen_dummy_magic_0.V_p_1.n6 48.0005
R7673 ref_volt_cur_gen_dummy_magic_0.V_p_1.n1 ref_volt_cur_gen_dummy_magic_0.V_p_1.n0 1.8755
R7674 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7675 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7676 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7677 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7678 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t33 660.109
R7679 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t30 660.109
R7680 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n14 428.8
R7681 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n15 428.8
R7682 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.n16 239.915
R7683 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.VD3.n17 239.915
R7684 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n19 230.4
R7685 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n21 230.4
R7686 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n14 198.4
R7687 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n15 198.4
R7688 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n11 160.428
R7689 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 160.427
R7690 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 160.427
R7691 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 160.053
R7692 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 159.803
R7693 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 159.803
R7694 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 159.802
R7695 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n3 159.802
R7696 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 159.802
R7697 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 155.302
R7698 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t32 155.125
R7699 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t35 155.125
R7700 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n27 146.002
R7701 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.VD3.t34 98.2764
R7702 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.t21 98.2764
R7703 two_stage_opamp_dummy_magic_0.VD3.t26 two_stage_opamp_dummy_magic_0.VD3.t36 98.2764
R7704 two_stage_opamp_dummy_magic_0.VD3.t23 two_stage_opamp_dummy_magic_0.VD3.t26 98.2764
R7705 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.VD3.t23 98.2764
R7706 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.t17 98.2764
R7707 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t28 98.2764
R7708 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.VD3.t12 98.2764
R7709 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t3 98.2764
R7710 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t31 98.2764
R7711 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.n14 92.5005
R7712 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n25 92.5005
R7713 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 92.5005
R7714 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 92.5005
R7715 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 92.5005
R7716 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.n23 92.5005
R7717 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t1 49.1384
R7718 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t19 49.1384
R7719 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 21.3338
R7720 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 21.3338
R7721 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n26 19.2005
R7722 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n28 13.8005
R7723 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t18 11.2576
R7724 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R7725 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t8 11.2576
R7726 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R7727 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R7728 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t10 11.2576
R7729 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t0 11.2576
R7730 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t14 11.2576
R7731 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R7732 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t16 11.2576
R7733 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R7734 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R7735 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R7736 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t6 11.2576
R7737 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R7738 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t4 11.2576
R7739 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R7740 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R7741 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R7742 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R7743 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t2 11.2576
R7744 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R7745 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n33 5.40675
R7746 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n8 4.5005
R7747 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n10 0.78175
R7748 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R7749 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R7750 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n6 0.6255
R7751 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n29 0.6255
R7752 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n13 0.6255
R7753 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n31 0.2505
R7754 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 628.034
R7755 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 626.784
R7756 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 626.784
R7757 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 289.2
R7758 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 289.2
R7759 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 228.252
R7760 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 212.733
R7761 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 212.733
R7762 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 176.733
R7763 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 176.733
R7764 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R7765 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 176.733
R7766 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 176.733
R7767 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 152
R7768 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 152
R7769 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R7770 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R7771 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 112.468
R7772 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 112.468
R7773 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R7774 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R7775 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 112.468
R7776 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 112.468
R7777 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 78.8005
R7778 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R7779 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R7780 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R7781 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 78.8005
R7782 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R7783 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 48.0005
R7784 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 48.0005
R7785 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R7786 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R7787 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 48.0005
R7788 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 48.0005
R7789 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 45.5227
R7790 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 45.5227
R7791 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 45.5227
R7792 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R7793 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 33.8443
R7794 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 14.2693
R7795 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 14.2693
R7796 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 1.2505
R7797 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 1.2505
R7798 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.n4 629.293
R7799 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.n7 628.668
R7800 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.n6 628.668
R7801 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.n5 628.668
R7802 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t33 611.739
R7803 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t20 611.739
R7804 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t26 611.739
R7805 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t36 611.739
R7806 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t38 421.75
R7807 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R7808 two_stage_opamp_dummy_magic_0.Vb3.n27 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R7809 two_stage_opamp_dummy_magic_0.Vb3.n28 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R7810 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R7811 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t39 421.75
R7812 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.t34 421.75
R7813 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R7814 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t32 421.75
R7815 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t29 421.75
R7816 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t35 421.75
R7817 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R7818 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t31 421.75
R7819 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t25 421.75
R7820 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R7821 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R7822 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t37 286.389
R7823 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t24 286.389
R7824 two_stage_opamp_dummy_magic_0.Vb3.n30 two_stage_opamp_dummy_magic_0.Vb3.n20 172.436
R7825 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 167.094
R7826 two_stage_opamp_dummy_magic_0.Vb3.n27 two_stage_opamp_dummy_magic_0.Vb3.n26 167.094
R7827 two_stage_opamp_dummy_magic_0.Vb3.n28 two_stage_opamp_dummy_magic_0.Vb3.n27 167.094
R7828 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 167.094
R7829 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 167.094
R7830 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 167.094
R7831 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R7832 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.n17 167.094
R7833 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R7834 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 167.094
R7835 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n13 167.094
R7836 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R7837 two_stage_opamp_dummy_magic_0.Vb3.n30 two_stage_opamp_dummy_magic_0.Vb3.n29 166.25
R7838 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 165.8
R7839 two_stage_opamp_dummy_magic_0.Vb3.n34 two_stage_opamp_dummy_magic_0.Vb3.n33 141.421
R7840 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n1 141.421
R7841 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 139.296
R7842 two_stage_opamp_dummy_magic_0.Vb3.n35 two_stage_opamp_dummy_magic_0.Vb3.n34 139.296
R7843 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t30 96.4005
R7844 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t17 96.4005
R7845 two_stage_opamp_dummy_magic_0.Vb3.n32 two_stage_opamp_dummy_magic_0.Vb3.n31 79.2817
R7846 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t3 65.6672
R7847 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t1 65.6672
R7848 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t7 65.6672
R7849 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t13 65.6672
R7850 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t4 65.6672
R7851 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t15 65.6672
R7852 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.t0 65.6672
R7853 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.t14 65.6672
R7854 two_stage_opamp_dummy_magic_0.Vb3.n29 two_stage_opamp_dummy_magic_0.Vb3.n28 47.1294
R7855 two_stage_opamp_dummy_magic_0.Vb3.n29 two_stage_opamp_dummy_magic_0.Vb3.n24 47.1294
R7856 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 47.1294
R7857 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n15 47.1294
R7858 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 38.5605
R7859 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n8 38.5605
R7860 two_stage_opamp_dummy_magic_0.Vb3.n33 two_stage_opamp_dummy_magic_0.Vb3.t10 24.0005
R7861 two_stage_opamp_dummy_magic_0.Vb3.n33 two_stage_opamp_dummy_magic_0.Vb3.t9 24.0005
R7862 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R7863 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t11 24.0005
R7864 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R7865 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R7866 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.Vb3.n35 24.0005
R7867 two_stage_opamp_dummy_magic_0.Vb3.n35 two_stage_opamp_dummy_magic_0.Vb3.t8 24.0005
R7868 two_stage_opamp_dummy_magic_0.Vb3.n31 two_stage_opamp_dummy_magic_0.Vb3.n30 16.5943
R7869 two_stage_opamp_dummy_magic_0.Vb3.n31 two_stage_opamp_dummy_magic_0.Vb3.n11 10.1567
R7870 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n0 4.938
R7871 two_stage_opamp_dummy_magic_0.Vb3.n32 two_stage_opamp_dummy_magic_0.Vb3.n3 4.34425
R7872 two_stage_opamp_dummy_magic_0.Vb3.n34 two_stage_opamp_dummy_magic_0.Vb3.n32 4.34425
R7873 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7874 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7875 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t14 449.868
R7876 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t18 449.868
R7877 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n21 340.397
R7878 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 339.272
R7879 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7880 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7881 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7882 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R7883 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7884 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7885 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7886 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7887 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7888 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7889 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7890 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7891 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R7892 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7893 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7894 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7895 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t1 184.498
R7896 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R7897 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.n15 176.733
R7898 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7899 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 176.733
R7900 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n11 176.733
R7901 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 176.733
R7902 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R7903 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.n6 176.733
R7904 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7905 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 176.733
R7906 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.n2 176.733
R7907 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R7908 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n9 170.269
R7909 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 165.8
R7910 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t0 58.5723
R7911 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 56.2338
R7912 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n13 56.2338
R7913 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 56.2338
R7914 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n4 56.2338
R7915 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n20 53.7505
R7916 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7917 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.t2 39.4005
R7918 two_stage_opamp_dummy_magic_0.Vb1.t3 two_stage_opamp_dummy_magic_0.Vb1.n23 39.4005
R7919 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7920 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 22.3599
R7921 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n0 7.09288
R7922 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n7 114.719
R7923 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7924 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n8 114.156
R7925 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7926 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7927 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7928 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7929 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7930 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7931 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7932 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7933 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7934 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7935 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7936 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7937 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7938 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7939 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7940 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7941 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7942 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7943 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7944 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7945 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7946 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7947 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7948 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7949 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7950 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7951 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7952 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7953 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7954 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7955 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7956 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7957 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7958 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7959 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7960 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7961 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 0.563
R7962 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7963 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7964 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7965 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7966 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7967 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7968 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7969 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7970 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7971 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7972 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7973 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7974 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7975 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7976 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7977 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7978 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7979 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7980 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7981 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7982 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7983 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7984 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7985 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7986 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7987 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7988 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7989 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7990 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7991 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7992 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7993 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7994 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7995 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7996 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7997 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7998 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7999 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.3272
R8000 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R8001 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R8002 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R8003 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R8004 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R8005 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.n0 237.327
R8006 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.t3 202.407
R8007 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n9 118.168
R8008 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.n2 117.831
R8009 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n16 117.269
R8010 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.n14 117.269
R8011 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.n12 117.269
R8012 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n10 117.269
R8013 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.n7 117.269
R8014 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.n5 117.269
R8015 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.n3 117.269
R8016 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.n1 113.136
R8017 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.n29 99.647
R8018 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.n37 99.0857
R8019 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n32 99.0845
R8020 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.n30 99.0845
R8021 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n27 99.0845
R8022 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.n25 99.0845
R8023 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.n23 99.0845
R8024 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.n34 94.5845
R8025 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n20 94.5845
R8026 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t27 24.0005
R8027 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t29 24.0005
R8028 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.t39 16.0005
R8029 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.t32 16.0005
R8030 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t40 16.0005
R8031 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t38 16.0005
R8032 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t0 16.0005
R8033 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t31 16.0005
R8034 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t34 16.0005
R8035 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t30 16.0005
R8036 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.t1 16.0005
R8037 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.t24 16.0005
R8038 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.t36 16.0005
R8039 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.t4 16.0005
R8040 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.t25 16.0005
R8041 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.t37 16.0005
R8042 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t35 16.0005
R8043 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t28 16.0005
R8044 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.t26 16.0005
R8045 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.t33 16.0005
R8046 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t23 16.0005
R8047 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t2 16.0005
R8048 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.t21 9.6005
R8049 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.t10 9.6005
R8050 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.t19 9.6005
R8051 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.t8 9.6005
R8052 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.t17 9.6005
R8053 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.t6 9.6005
R8054 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t15 9.6005
R8055 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t12 9.6005
R8056 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t5 9.6005
R8057 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t14 9.6005
R8058 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.t7 9.6005
R8059 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.t16 9.6005
R8060 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.t9 9.6005
R8061 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.t18 9.6005
R8062 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t11 9.6005
R8063 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t20 9.6005
R8064 two_stage_opamp_dummy_magic_0.V_p.t22 two_stage_opamp_dummy_magic_0.V_p.n38 9.6005
R8065 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.t13 9.6005
R8066 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n35 4.5005
R8067 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.n18 4.5005
R8068 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.n21 4.5005
R8069 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n17 3.65675
R8070 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n19 1.28175
R8071 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n31 0.563
R8072 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n33 0.563
R8073 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n36 0.563
R8074 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.n11 0.563
R8075 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.n13 0.563
R8076 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n15 0.563
R8077 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.n4 0.563
R8078 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.n6 0.563
R8079 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.n22 0.563
R8080 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.n24 0.563
R8081 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n26 0.563
R8082 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n28 0.563
R8083 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n8 0.53175
R8084 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R8085 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R8086 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R8087 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R8088 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R8089 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R8090 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R8091 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.n0 165.8
R8092 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R8093 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R8094 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R8095 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R8096 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R8097 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R8098 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t3 117.591
R8099 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t2 117.591
R8100 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t1 108.424
R8101 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 108.424
R8102 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 42.9559
R8103 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 21.6434
R8104 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n8 17.0005
R8105 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 3.31612
R8106 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 1.26612
R8107 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.2505
R8108 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n4 1.15363
R8109 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 2445
R8110 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2430
R8111 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 2430
R8112 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2415
R8113 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t20 650.668
R8114 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t23 650.668
R8115 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n22 637.288
R8116 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n25 636.663
R8117 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n23 636.663
R8118 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 628.668
R8119 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 628.668
R8120 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n21 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 624.168
R8121 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t22 387.329
R8122 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 356.495
R8123 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t21 310.659
R8124 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t18 310.659
R8125 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 259.2
R8126 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 257.601
R8127 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t19 196.553
R8128 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t14 196.553
R8129 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 196.553
R8130 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 196.553
R8131 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t12 196.553
R8132 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t22 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 196.553
R8133 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 153.601
R8134 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 153.601
R8135 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 107.201
R8136 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 105.6
R8137 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t16 98.2764
R8138 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 98.2764
R8139 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8140 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8141 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 92.5005
R8142 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8143 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 92.5005
R8144 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t15 65.6672
R8145 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 65.6672
R8146 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t17 65.6672
R8147 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t11 65.6672
R8148 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t13 65.6672
R8149 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 65.6672
R8150 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 61.6672
R8151 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 49.2505
R8152 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 49.2505
R8153 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 49.2505
R8154 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 49.2505
R8155 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n22 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 49.2505
R8156 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n22 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 49.2505
R8157 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 44.2922
R8158 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 44.2922
R8159 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 27.7338
R8160 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 27.7338
R8161 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 21.3338
R8162 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 21.3338
R8163 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n21 7.188
R8164 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n21 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n20 4.5005
R8165 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n26 1.688
R8166 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n24 0.6255
R8167 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n19 0.6255
R8168 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 0.6255
R8169 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n19 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n0 392.666
R8170 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n10 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t16 273.134
R8171 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n9 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t14 273.134
R8172 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n7 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t22 273.134
R8173 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n4 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t6 273.134
R8174 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n1 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t12 273.134
R8175 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t2 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n18 273.134
R8176 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n11 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n10 224.934
R8177 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n12 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n11 224.934
R8178 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n5 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n4 224.934
R8179 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n6 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n5 224.934
R8180 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n2 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n1 224.934
R8181 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n3 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n2 224.934
R8182 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n17 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n16 224.934
R8183 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n18 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n17 224.934
R8184 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n19 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t2 200.201
R8185 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n14 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n13 171.582
R8186 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n14 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n8 171.582
R8187 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n15 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n14 166.113
R8188 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n20 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n19 150.876
R8189 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n13 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n12 69.6227
R8190 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n13 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n9 69.6227
R8191 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n8 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n7 69.6227
R8192 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n8 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n6 69.6227
R8193 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n15 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n3 69.6227
R8194 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n16 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n15 69.6227
R8195 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n10 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t9 48.2005
R8196 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n11 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t7 48.2005
R8197 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n12 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t5 48.2005
R8198 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n9 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t21 48.2005
R8199 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n7 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t19 48.2005
R8200 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n4 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t8 48.2005
R8201 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n5 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t11 48.2005
R8202 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n6 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t18 48.2005
R8203 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n1 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t20 48.2005
R8204 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n2 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t23 48.2005
R8205 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n3 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t10 48.2005
R8206 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n16 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t13 48.2005
R8207 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n17 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t15 48.2005
R8208 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n18 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t17 48.2005
R8209 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n0 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t1 39.4005
R8210 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n0 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t0 39.4005
R8211 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t3 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n20 24.0005
R8212 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.n20 ref_volt_cur_gen_dummy_magic_0.NFET_GATE_10uA.t4 24.0005
R8213 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 145.702
R8214 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 134.577
R8215 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 108.66
R8216 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 97.4009
R8217 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 96.8384
R8218 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 96.8384
R8219 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 96.8384
R8220 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 96.8384
R8221 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 48.7817
R8222 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 24.0005
R8223 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 24.0005
R8224 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 24.0005
R8225 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 24.0005
R8226 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 18.4067
R8227 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R8228 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R8229 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R8230 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R8231 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R8232 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R8233 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R8234 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 8.0005
R8235 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R8236 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R8237 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 0.563
R8238 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 0.563
R8239 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.563
R8240 VIN-.n4 VIN-.t8 485.021
R8241 VIN-.n1 VIN-.t6 484.159
R8242 VIN-.n5 VIN-.t7 483.358
R8243 VIN-.n8 VIN-.t10 431.536
R8244 VIN-.n2 VIN-.t9 431.536
R8245 VIN-.n6 VIN-.t1 431.257
R8246 VIN-.n0 VIN-.t0 431.257
R8247 VIN-.n6 VIN-.t2 289.908
R8248 VIN-.n0 VIN-.t5 289.908
R8249 VIN-.n8 VIN-.t4 279.183
R8250 VIN-.n2 VIN-.t3 279.183
R8251 VIN-.n7 VIN-.n6 233.374
R8252 VIN-.n1 VIN-.n0 233.374
R8253 VIN-.n9 VIN-.n8 188.989
R8254 VIN-.n3 VIN-.n2 188.989
R8255 VIN-.n4 VIN-.n3 2.463
R8256 VIN- VIN-.n9 2.03175
R8257 VIN-.n5 VIN-.n4 1.563
R8258 VIN-.n3 VIN-.n1 1.2755
R8259 VIN-.n9 VIN-.n7 1.2755
R8260 VIN-.n7 VIN-.n5 0.8005
R8261 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 206.052
R8262 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 205.488
R8263 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 205.488
R8264 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 205.488
R8265 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 205.488
R8266 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 182.701
R8267 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 181.701
R8268 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 181.701
R8269 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 121.192
R8270 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 57.7817
R8271 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 19.7005
R8272 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R8273 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R8274 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R8275 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R8276 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R8277 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R8278 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R8279 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R8280 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 19.7005
R8281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 15.7605
R8282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 15.7605
R8283 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 15.7605
R8284 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 15.7605
R8285 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 15.7605
R8286 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 15.7605
R8287 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 6.1255
R8288 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 4.438
R8289 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 1.0005
R8290 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R8291 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 0.563
R8292 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 0.563
R8293 ref_volt_cur_gen_dummy_magic_0.START_UP_NFET1.t0 ref_volt_cur_gen_dummy_magic_0.START_UP_NFET1.t1 178.194
R8294 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 621.268
R8295 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t24 611.739
R8296 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t10 611.739
R8297 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t18 611.739
R8298 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t27 611.739
R8299 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R8300 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t33 421.75
R8301 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t9 421.75
R8302 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R8303 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t34 421.75
R8304 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.t31 421.75
R8305 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R8306 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R8307 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R8308 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R8309 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R8310 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R8311 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t22 421.75
R8312 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R8313 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R8314 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R8315 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t1 288.166
R8316 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t12 262.288
R8317 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n6 172.811
R8318 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 169.125
R8319 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n18 169.125
R8320 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n23 167.094
R8321 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 167.094
R8322 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.n25 167.094
R8323 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 167.094
R8324 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 167.094
R8325 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 167.094
R8326 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.n14 167.094
R8327 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R8328 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R8329 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.n10 167.094
R8330 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R8331 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R8332 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R8333 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.n3 167.094
R8334 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R8335 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t32 142.325
R8336 two_stage_opamp_dummy_magic_0.Vb2.n31 two_stage_opamp_dummy_magic_0.Vb2.n0 140.077
R8337 two_stage_opamp_dummy_magic_0.Vb2.n32 two_stage_opamp_dummy_magic_0.Vb2.n31 140.077
R8338 two_stage_opamp_dummy_magic_0.Vb2.n30 two_stage_opamp_dummy_magic_0.Vb2.n1 134.577
R8339 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t30 72.3005
R8340 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t16 72.3005
R8341 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t28 72.3005
R8342 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t14 72.3005
R8343 two_stage_opamp_dummy_magic_0.Vb2.n30 two_stage_opamp_dummy_magic_0.Vb2.n29 69.563
R8344 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t0 62.5402
R8345 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t2 62.5402
R8346 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n26 47.1294
R8347 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n22 47.1294
R8348 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 47.1294
R8349 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n13 47.1294
R8350 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n5 47.1294
R8351 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 37.3443
R8352 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R8353 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R8354 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t8 24.0005
R8355 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R8356 two_stage_opamp_dummy_magic_0.Vb2.t7 two_stage_opamp_dummy_magic_0.Vb2.n32 24.0005
R8357 two_stage_opamp_dummy_magic_0.Vb2.n32 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R8358 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 14.6443
R8359 two_stage_opamp_dummy_magic_0.Vb2.n31 two_stage_opamp_dummy_magic_0.Vb2.n30 4.5005
R8360 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n9 2.09425
R8361 a_5230_5852.t0 a_5230_5852.t1 304.579
R8362 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n3 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n2 526.183
R8363 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n1 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n0 514.134
R8364 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n0 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t4 303.259
R8365 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n5 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n4 287.264
R8366 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n5 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n3 282.522
R8367 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t2 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n5 262.411
R8368 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n0 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t5 174.726
R8369 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n1 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t7 174.726
R8370 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n2 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t6 174.726
R8371 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n2 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n1 128.534
R8372 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n3 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t3 96.4005
R8373 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n4 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t0 39.4005
R8374 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.n4 ref_volt_cur_gen_dummy_magic_0.V_CUR_REF_REG.t1 39.4005
R8375 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8376 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8377 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8378 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8379 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t0 660.109
R8380 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t3 660.109
R8381 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 428.8
R8382 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n0 428.8
R8383 two_stage_opamp_dummy_magic_0.VD4.t1 two_stage_opamp_dummy_magic_0.VD4.n8 239.915
R8384 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t4 239.915
R8385 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 230.4
R8386 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n3 230.4
R8387 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 198.4
R8388 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n0 198.4
R8389 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n28 160.428
R8390 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 160.427
R8391 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n14 160.427
R8392 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n13 160.053
R8393 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n29 159.803
R8394 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.803
R8395 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 159.802
R8396 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 159.802
R8397 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 159.802
R8398 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n23 155.302
R8399 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t2 155.125
R8400 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t5 155.125
R8401 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 146.004
R8402 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t1 98.2764
R8403 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t18 98.2764
R8404 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.VD4.t24 98.2764
R8405 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.VD4.t32 98.2764
R8406 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.VD4.t28 98.2764
R8407 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t36 98.2764
R8408 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t20 98.2764
R8409 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.VD4.t26 98.2764
R8410 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.VD4.t22 98.2764
R8411 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.VD4.t30 98.2764
R8412 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R8413 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.n6 92.5005
R8414 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n7 92.5005
R8415 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n0 92.5005
R8416 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8417 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8418 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t34 49.1384
R8419 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.VD4.n9 49.1384
R8420 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n4 21.3338
R8421 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.n2 21.3338
R8422 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n12 19.2005
R8423 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 13.8005
R8424 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R8425 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R8426 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R8427 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R8428 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t33 11.2576
R8429 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R8430 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R8431 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R8432 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R8433 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t14 11.2576
R8434 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R8435 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8436 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R8437 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R8438 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t12 11.2576
R8439 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R8440 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t16 11.2576
R8441 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R8442 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R8443 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R8444 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t35 11.2576
R8445 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.VD4.n33 11.2576
R8446 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 6.188
R8447 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n22 4.5005
R8448 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 0.6255
R8449 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n17 0.6255
R8450 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n19 0.6255
R8451 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 0.6255
R8452 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n27 0.6255
R8453 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.2505
R8454 VIN+.n9 VIN+.t5 485.127
R8455 VIN+.n4 VIN+.t3 485.127
R8456 VIN+.n3 VIN+.t4 485.127
R8457 VIN+.n7 VIN+.t9 318.656
R8458 VIN+.n7 VIN+.t2 318.656
R8459 VIN+.n5 VIN+.t7 318.656
R8460 VIN+.n5 VIN+.t1 318.656
R8461 VIN+.n1 VIN+.t8 318.656
R8462 VIN+.n1 VIN+.t6 318.656
R8463 VIN+.n0 VIN+.t10 318.656
R8464 VIN+.n0 VIN+.t0 318.656
R8465 VIN+.n2 VIN+.n0 167.05
R8466 VIN+.n8 VIN+.n7 165.8
R8467 VIN+.n6 VIN+.n5 165.8
R8468 VIN+.n2 VIN+.n1 165.8
R8469 VIN+.n6 VIN+.n4 2.34425
R8470 VIN+.n4 VIN+.n3 1.3005
R8471 VIN+.n8 VIN+.n6 1.2505
R8472 VIN+ VIN+.n9 1.213
R8473 VIN+.n3 VIN+.n2 1.15675
R8474 VIN+.n9 VIN+.n8 1.15675
R8475 a_n9700_9790.t0 a_n9700_9790.t1 258.591
R8476 a_14520_5852.t0 a_14520_5852.t1 305.31
R8477 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n6 630.607
R8478 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 627.128
R8479 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n10 627.128
R8480 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t12 410.666
R8481 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 227.784
R8482 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 226.534
R8483 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n3 226.534
R8484 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8485 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t11 78.8005
R8486 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t8 78.8005
R8487 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t10 78.8005
R8488 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t7 78.8005
R8489 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t9 78.8005
R8490 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t2 48.0005
R8491 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t4 48.0005
R8492 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t1 48.0005
R8493 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t3 48.0005
R8494 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R8495 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t5 48.0005
R8496 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n5 21.1255
R8497 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.n4 10.8755
R8498 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n7 1.3755
R8499 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.2505
R8500 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 1.2505
R8501 ref_volt_cur_gen_dummy_magic_0.Vin-.n11 ref_volt_cur_gen_dummy_magic_0.Vin-.t9 688.859
R8502 ref_volt_cur_gen_dummy_magic_0.Vin-.n13 ref_volt_cur_gen_dummy_magic_0.Vin-.n12 514.134
R8503 ref_volt_cur_gen_dummy_magic_0.Vin-.n9 ref_volt_cur_gen_dummy_magic_0.Vin-.n8 345.116
R8504 ref_volt_cur_gen_dummy_magic_0.Vin-.n15 ref_volt_cur_gen_dummy_magic_0.Vin-.n14 214.713
R8505 ref_volt_cur_gen_dummy_magic_0.Vin-.n11 ref_volt_cur_gen_dummy_magic_0.Vin-.t11 174.726
R8506 ref_volt_cur_gen_dummy_magic_0.Vin-.n12 ref_volt_cur_gen_dummy_magic_0.Vin-.t12 174.726
R8507 ref_volt_cur_gen_dummy_magic_0.Vin-.n13 ref_volt_cur_gen_dummy_magic_0.Vin-.t8 174.726
R8508 ref_volt_cur_gen_dummy_magic_0.Vin-.n14 ref_volt_cur_gen_dummy_magic_0.Vin-.t10 174.726
R8509 ref_volt_cur_gen_dummy_magic_0.Vin-.n7 ref_volt_cur_gen_dummy_magic_0.Vin-.n5 173.029
R8510 ref_volt_cur_gen_dummy_magic_0.Vin-.n7 ref_volt_cur_gen_dummy_magic_0.Vin-.n6 168.654
R8511 ref_volt_cur_gen_dummy_magic_0.Vin-.n9 ref_volt_cur_gen_dummy_magic_0.Vin-.t0 162.921
R8512 ref_volt_cur_gen_dummy_magic_0.Vin-.n12 ref_volt_cur_gen_dummy_magic_0.Vin-.n11 128.534
R8513 ref_volt_cur_gen_dummy_magic_0.Vin-.n14 ref_volt_cur_gen_dummy_magic_0.Vin-.n13 128.534
R8514 ref_volt_cur_gen_dummy_magic_0.Vin-.n1 ref_volt_cur_gen_dummy_magic_0.Vin-.n0 83.5719
R8515 ref_volt_cur_gen_dummy_magic_0.Vin-.n22 ref_volt_cur_gen_dummy_magic_0.Vin-.n21 83.5719
R8516 ref_volt_cur_gen_dummy_magic_0.Vin-.n20 ref_volt_cur_gen_dummy_magic_0.Vin-.n19 83.5719
R8517 ref_volt_cur_gen_dummy_magic_0.Vin-.n25 ref_volt_cur_gen_dummy_magic_0.Vin-.n1 73.682
R8518 ref_volt_cur_gen_dummy_magic_0.Vin-.n20 ref_volt_cur_gen_dummy_magic_0.Vin-.n4 73.3165
R8519 ref_volt_cur_gen_dummy_magic_0.Vin-.n8 ref_volt_cur_gen_dummy_magic_0.Vin-.t2 39.4005
R8520 ref_volt_cur_gen_dummy_magic_0.Vin-.n8 ref_volt_cur_gen_dummy_magic_0.Vin-.t1 39.4005
R8521 ref_volt_cur_gen_dummy_magic_0.Vin-.n21 ref_volt_cur_gen_dummy_magic_0.Vin-.n20 26.074
R8522 ref_volt_cur_gen_dummy_magic_0.Vin-.t7 ref_volt_cur_gen_dummy_magic_0.Vin-.n1 25.7843
R8523 ref_volt_cur_gen_dummy_magic_0.Vin-.n16 ref_volt_cur_gen_dummy_magic_0.Vin-.n15 17.526
R8524 ref_volt_cur_gen_dummy_magic_0.Vin-.n6 ref_volt_cur_gen_dummy_magic_0.Vin-.t6 13.1338
R8525 ref_volt_cur_gen_dummy_magic_0.Vin-.n6 ref_volt_cur_gen_dummy_magic_0.Vin-.t3 13.1338
R8526 ref_volt_cur_gen_dummy_magic_0.Vin-.n5 ref_volt_cur_gen_dummy_magic_0.Vin-.t5 13.1338
R8527 ref_volt_cur_gen_dummy_magic_0.Vin-.n5 ref_volt_cur_gen_dummy_magic_0.Vin-.t4 13.1338
R8528 ref_volt_cur_gen_dummy_magic_0.Vin-.n15 ref_volt_cur_gen_dummy_magic_0.Vin-.n10 12.5317
R8529 ref_volt_cur_gen_dummy_magic_0.Vin-.n10 ref_volt_cur_gen_dummy_magic_0.Vin-.n9 6.40675
R8530 ref_volt_cur_gen_dummy_magic_0.Vin-.n10 ref_volt_cur_gen_dummy_magic_0.Vin-.n7 3.8755
R8531 ref_volt_cur_gen_dummy_magic_0.Vin-.n16 ref_volt_cur_gen_dummy_magic_0.Vin-.n4 2.19742
R8532 ref_volt_cur_gen_dummy_magic_0.Vin-.n24 ref_volt_cur_gen_dummy_magic_0.Vin-.n23 1.5505
R8533 ref_volt_cur_gen_dummy_magic_0.Vin-.n3 ref_volt_cur_gen_dummy_magic_0.Vin-.n2 1.5505
R8534 ref_volt_cur_gen_dummy_magic_0.Vin-.n18 ref_volt_cur_gen_dummy_magic_0.Vin-.n17 1.5505
R8535 ref_volt_cur_gen_dummy_magic_0.Vin-.n18 ref_volt_cur_gen_dummy_magic_0.Vin-.n4 1.19225
R8536 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter ref_volt_cur_gen_dummy_magic_0.Vin-.n25 1.07742
R8537 ref_volt_cur_gen_dummy_magic_0.Vin-.n23 ref_volt_cur_gen_dummy_magic_0.Vin-.n22 1.07024
R8538 ref_volt_cur_gen_dummy_magic_0.Vin-.n19 ref_volt_cur_gen_dummy_magic_0.Vin-.n18 0.959578
R8539 ref_volt_cur_gen_dummy_magic_0.Vin-.n19 ref_volt_cur_gen_dummy_magic_0.Vin-.n3 0.885803
R8540 ref_volt_cur_gen_dummy_magic_0.Vin-.n22 ref_volt_cur_gen_dummy_magic_0.Vin-.n3 0.77514
R8541 ref_volt_cur_gen_dummy_magic_0.Vin-.n25 ref_volt_cur_gen_dummy_magic_0.Vin-.n24 0.763532
R8542 ref_volt_cur_gen_dummy_magic_0.Vin-.n23 ref_volt_cur_gen_dummy_magic_0.Vin-.n0 0.590702
R8543 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter ref_volt_cur_gen_dummy_magic_0.Vin-.n0 0.498483
R8544 ref_volt_cur_gen_dummy_magic_0.Vin-.n21 ref_volt_cur_gen_dummy_magic_0.Vin-.t7 0.290206
R8545 ref_volt_cur_gen_dummy_magic_0.Vin-.n17 ref_volt_cur_gen_dummy_magic_0.Vin-.n16 0.0183571
R8546 ref_volt_cur_gen_dummy_magic_0.Vin-.n17 ref_volt_cur_gen_dummy_magic_0.Vin-.n2 0.0183571
R8547 ref_volt_cur_gen_dummy_magic_0.Vin-.n24 ref_volt_cur_gen_dummy_magic_0.Vin-.n2 0.0183571
R8548 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 220.678
R8549 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R8550 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t2 16.0005
R8551 two_stage_opamp_dummy_magic_0.V_p_mir.t1 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R8552 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t0 9.6005
R8553 a_14640_5852.t0 a_14640_5852.t1 169.905
R8554 a_14240_2946.t0 a_14240_2946.t1 169.905
R8555 a_5350_5852.t0 a_5350_5852.t1 169.905
R8556 a_n8798_9040.t0 a_n8798_9040.t1 376.99
R8557 a_n7190_9400.t0 a_n7190_9400.t1 258.591
R8558 a_n9760_9260.t0 a_n9760_9260.t1 258.591
C0 VIN+ two_stage_opamp_dummy_magic_0.VD1 0.057219f
C1 VDDA ref_volt_cur_gen_dummy_magic_0.V_TOP 16.055f
C2 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 ref_volt_cur_gen_dummy_magic_0.V_TOP 1.39829f
C3 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.err_amp_out 0.040365f
C4 VDDA ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 2.81641f
C5 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.err_amp_out 0.017581f
C6 VDDA VOUT- 6.77346f
C7 VDDA two_stage_opamp_dummy_magic_0.V_err_gate 3.58589f
C8 VDDA two_stage_opamp_dummy_magic_0.cap_res_X 0.983966f
C9 VDDA VOUT+ 6.69238f
C10 VOUT- two_stage_opamp_dummy_magic_0.V_err_gate 0.068595f
C11 VOUT- two_stage_opamp_dummy_magic_0.cap_res_X 50.7528f
C12 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.V_err_gate 0.356357f
C13 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.VD1 1.06369f
C14 ref_volt_cur_gen_dummy_magic_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.10577f
C15 VDDA two_stage_opamp_dummy_magic_0.V_err_amp_ref 3.98206f
C16 VOUT- VOUT+ 0.210644f
C17 VOUT+ two_stage_opamp_dummy_magic_0.cap_res_X 0.020189f
C18 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.24899f
C19 VDDA m2_n2790_7140# 0.010446f
C20 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 m2_n2790_7140# 0.075543f
C21 VOUT- two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.068695f
C22 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 4.78237f
C23 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.25369f
C24 VDDA two_stage_opamp_dummy_magic_0.VD3 3.70112f
C25 VDDA two_stage_opamp_dummy_magic_0.Vb2_Vb3 1.65321f
C26 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.VD3 0.01134f
C27 VDDA two_stage_opamp_dummy_magic_0.err_amp_out 1.00936f
C28 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.012774f
C29 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.014914f
C30 VOUT+ two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.03526f
C31 VIN- VIN+ 0.555219f
C32 VDDA two_stage_opamp_dummy_magic_0.Y 4.15025f
C33 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.406563f
C34 ref_volt_cur_gen_dummy_magic_0.V_TOP m2_n4150_7140# 0.012f
C35 VDDA m2_n4150_7140# 0.010446f
C36 VOUT+ two_stage_opamp_dummy_magic_0.Y 2.10995f
C37 VIN- two_stage_opamp_dummy_magic_0.VD1 0.881219f
C38 VIN+ GNDA 2.09054f
C39 VIN- GNDA 2.157042f
C40 VOUT+ GNDA 17.828459f
C41 VOUT- GNDA 17.39849f
C42 VDDA GNDA 0.161808p
C43 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.38775f
C44 two_stage_opamp_dummy_magic_0.Y GNDA 4.961036f
C45 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 32.22025f
C46 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2 GNDA 4.662062f
C47 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 3.001013f
C48 ref_volt_cur_gen_dummy_magic_0.V_TOP GNDA 6.652324f
C49 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 8.904718f
C50 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 8.838531f
C51 two_stage_opamp_dummy_magic_0.VD3 GNDA 6.53628f
C52 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.42123f
C53 ref_volt_cur_gen_dummy_magic_0.Vin-.n0 GNDA 0.048818f
C54 ref_volt_cur_gen_dummy_magic_0.Vin-.n1 GNDA 0.333648f
C55 ref_volt_cur_gen_dummy_magic_0.Vin-.n2 GNDA 0.166915f
C56 ref_volt_cur_gen_dummy_magic_0.Vin-.n3 GNDA 0.074468f
C57 ref_volt_cur_gen_dummy_magic_0.Vin-.n4 GNDA 0.338979f
C58 ref_volt_cur_gen_dummy_magic_0.Vin-.t5 GNDA 0.028614f
C59 ref_volt_cur_gen_dummy_magic_0.Vin-.t4 GNDA 0.028614f
C60 ref_volt_cur_gen_dummy_magic_0.Vin-.n5 GNDA 0.099613f
C61 ref_volt_cur_gen_dummy_magic_0.Vin-.t6 GNDA 0.028614f
C62 ref_volt_cur_gen_dummy_magic_0.Vin-.t3 GNDA 0.028614f
C63 ref_volt_cur_gen_dummy_magic_0.Vin-.n6 GNDA 0.095121f
C64 ref_volt_cur_gen_dummy_magic_0.Vin-.n7 GNDA 0.408067f
C65 ref_volt_cur_gen_dummy_magic_0.Vin-.t0 GNDA 0.098662f
C66 ref_volt_cur_gen_dummy_magic_0.Vin-.n8 GNDA 0.025702f
C67 ref_volt_cur_gen_dummy_magic_0.Vin-.n9 GNDA 0.469862f
C68 ref_volt_cur_gen_dummy_magic_0.Vin-.n10 GNDA 0.222852f
C69 ref_volt_cur_gen_dummy_magic_0.Vin-.t9 GNDA 0.023594f
C70 ref_volt_cur_gen_dummy_magic_0.Vin-.n11 GNDA 0.027673f
C71 ref_volt_cur_gen_dummy_magic_0.Vin-.n12 GNDA 0.022653f
C72 ref_volt_cur_gen_dummy_magic_0.Vin-.n13 GNDA 0.022653f
C73 ref_volt_cur_gen_dummy_magic_0.Vin-.n14 GNDA 0.040466f
C74 ref_volt_cur_gen_dummy_magic_0.Vin-.n15 GNDA 0.524007f
C75 ref_volt_cur_gen_dummy_magic_0.Vin-.n16 GNDA 0.461299f
C76 ref_volt_cur_gen_dummy_magic_0.Vin-.n17 GNDA 0.166915f
C77 ref_volt_cur_gen_dummy_magic_0.Vin-.n18 GNDA 0.10855f
C78 ref_volt_cur_gen_dummy_magic_0.Vin-.n19 GNDA 0.082742f
C79 ref_volt_cur_gen_dummy_magic_0.Vin-.n20 GNDA 0.331333f
C80 ref_volt_cur_gen_dummy_magic_0.Vin-.t7 GNDA 0.072966f
C81 ref_volt_cur_gen_dummy_magic_0.Vin-.n21 GNDA 0.073776f
C82 ref_volt_cur_gen_dummy_magic_0.Vin-.n22 GNDA 0.082742f
C83 ref_volt_cur_gen_dummy_magic_0.Vin-.n23 GNDA 0.074468f
C84 ref_volt_cur_gen_dummy_magic_0.Vin-.n24 GNDA 0.656866f
C85 ref_volt_cur_gen_dummy_magic_0.Vin-.n25 GNDA 0.389111f
C86 ref_volt_cur_gen_dummy_magic_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.086659f
C87 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA 0.013323f
C88 two_stage_opamp_dummy_magic_0.err_amp_out.t3 GNDA 0.013323f
C89 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.038344f
C90 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA 0.013323f
C91 two_stage_opamp_dummy_magic_0.err_amp_out.t4 GNDA 0.013323f
C92 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.037203f
C93 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.462683f
C94 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA 0.013323f
C95 two_stage_opamp_dummy_magic_0.err_amp_out.t5 GNDA 0.013323f
C96 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.037203f
C97 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.493922f
C98 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.059015f
C99 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 1.65781f
C100 two_stage_opamp_dummy_magic_0.err_amp_out.t0 GNDA 0.013323f
C101 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA 0.013323f
C102 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 0.030943f
C103 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.914249f
C104 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA 0.013323f
C105 two_stage_opamp_dummy_magic_0.err_amp_out.t10 GNDA 0.013323f
C106 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.031191f
C107 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.349833f
C108 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA 0.013323f
C109 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA 0.013323f
C110 two_stage_opamp_dummy_magic_0.err_amp_out.n10 GNDA 0.031191f
C111 VIN+.t0 GNDA 0.041803f
C112 VIN+.t10 GNDA 0.041803f
C113 VIN+.n0 GNDA 0.086391f
C114 VIN+.t6 GNDA 0.041803f
C115 VIN+.t8 GNDA 0.041803f
C116 VIN+.n1 GNDA 0.085194f
C117 VIN+.n2 GNDA 0.359761f
C118 VIN+.t4 GNDA 0.058811f
C119 VIN+.n3 GNDA 0.215335f
C120 VIN+.t3 GNDA 0.058811f
C121 VIN+.n4 GNDA 0.262589f
C122 VIN+.t1 GNDA 0.041803f
C123 VIN+.t7 GNDA 0.041803f
C124 VIN+.n5 GNDA 0.085194f
C125 VIN+.n6 GNDA 0.248358f
C126 VIN+.t2 GNDA 0.041803f
C127 VIN+.t9 GNDA 0.041803f
C128 VIN+.n7 GNDA 0.085194f
C129 VIN+.n8 GNDA 0.200956f
C130 VIN+.t5 GNDA 0.058811f
C131 VIN+.n9 GNDA 0.211601f
C132 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.024416f
C133 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.069509f
C134 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.094519f
C135 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.120449f
C136 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.042516f
C137 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.078578f
C138 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.050655f
C139 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.120449f
C140 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.042516f
C141 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.078578f
C142 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.050655f
C143 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.050227f
C144 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.094519f
C145 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.281683f
C146 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.420453f
C147 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.242764f
C148 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.242764f
C149 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.242764f
C150 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.242764f
C151 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.182073f
C152 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.121382f
C153 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.182073f
C154 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.242764f
C155 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.242764f
C156 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.242764f
C157 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.242764f
C158 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.420453f
C159 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.281683f
C160 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.069509f
C161 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.097309f
C162 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.024416f
C163 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.024416f
C164 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.084727f
C165 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.024416f
C166 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.024416f
C167 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.084913f
C168 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.024416f
C169 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.024416f
C170 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.084913f
C171 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.024416f
C172 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.024416f
C173 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.084613f
C174 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.15974f
C175 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.024416f
C176 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.024416f
C177 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.084613f
C178 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.082811f
C179 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.024416f
C180 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.024416f
C181 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.084613f
C182 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.082811f
C183 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.099252f
C184 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.024416f
C185 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.024416f
C186 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.08286f
C187 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.100481f
C188 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.094683f
C189 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.024416f
C190 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.024416f
C191 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.084612f
C192 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.078625f
C193 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.024416f
C194 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.024416f
C195 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.084913f
C196 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.024416f
C197 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.024416f
C198 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.084612f
C199 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.15974f
C200 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.029845f
C201 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.057972f
C202 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.079606f
C203 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.024416f
C204 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.023814f
C205 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.023814f
C206 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.023814f
C207 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.077376f
C208 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.023814f
C209 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.023814f
C210 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.071929f
C211 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.014289f
C212 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.014289f
C213 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.014289f
C214 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.014289f
C215 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.031614f
C216 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.04221f
C217 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.03334f
C218 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.03334f
C219 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.029021f
C220 two_stage_opamp_dummy_magic_0.Vb2.t32 GNDA 0.022707f
C221 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.067799f
C222 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.015003f
C223 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.015003f
C224 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.032578f
C225 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.046595f
C226 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.157984f
C227 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.83403f
C228 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.117881f
C229 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.117881f
C230 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.117881f
C231 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.117881f
C232 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.136033f
C233 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.110444f
C234 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.067871f
C235 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.067871f
C236 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.063552f
C237 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.117881f
C238 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.117881f
C239 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.117881f
C240 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.117881f
C241 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.136033f
C242 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.110444f
C243 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.067871f
C244 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.067871f
C245 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.063552f
C246 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.042509f
C247 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.117881f
C248 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.117881f
C249 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.117881f
C250 two_stage_opamp_dummy_magic_0.Vb2.t34 GNDA 0.117881f
C251 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.136033f
C252 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.110444f
C253 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.067871f
C254 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.067871f
C255 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 0.063552f
C256 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.117881f
C257 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.117881f
C258 two_stage_opamp_dummy_magic_0.Vb2.t33 GNDA 0.117881f
C259 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.117881f
C260 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.136033f
C261 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.110444f
C262 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.067871f
C263 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.067871f
C264 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.063552f
C265 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.042509f
C266 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 1.5622f
C267 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 3.36171f
C268 two_stage_opamp_dummy_magic_0.Vb2.n30 GNDA 2.14572f
C269 two_stage_opamp_dummy_magic_0.Vb2.n31 GNDA 0.488234f
C270 two_stage_opamp_dummy_magic_0.Vb2.n32 GNDA 0.077376f
C271 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.023814f
C272 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.080817f
C273 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.012915f
C274 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.012915f
C275 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.037893f
C276 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.012915f
C277 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.012915f
C278 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.037721f
C279 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.130385f
C280 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.012915f
C281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.012915f
C282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.037721f
C283 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.067538f
C284 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.012915f
C285 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.012915f
C286 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.037721f
C287 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.067538f
C288 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.012915f
C289 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.012915f
C290 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.037721f
C291 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.097494f
C292 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.697459f
C293 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.016144f
C294 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.016144f
C295 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.052448f
C296 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.016144f
C297 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.016144f
C298 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.052068f
C299 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.147331f
C300 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.016144f
C301 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.016144f
C302 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.052068f
C303 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 0.113865f
C304 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S3 GNDA 0.626194f
C305 VIN-.t6 GNDA 0.050642f
C306 VIN-.t5 GNDA 0.033412f
C307 VIN-.t0 GNDA 0.041251f
C308 VIN-.n0 GNDA 0.059274f
C309 VIN-.n1 GNDA 0.280478f
C310 VIN-.t3 GNDA 0.032863f
C311 VIN-.t9 GNDA 0.041265f
C312 VIN-.n2 GNDA 0.064892f
C313 VIN-.n3 GNDA 0.200879f
C314 VIN-.t8 GNDA 0.050078f
C315 VIN-.n4 GNDA 0.236241f
C316 VIN-.t7 GNDA 0.050425f
C317 VIN-.n5 GNDA 0.180621f
C318 VIN-.t2 GNDA 0.033412f
C319 VIN-.t1 GNDA 0.041251f
C320 VIN-.n6 GNDA 0.059274f
C321 VIN-.n7 GNDA 0.149629f
C322 VIN-.t4 GNDA 0.032863f
C323 VIN-.t10 GNDA 0.041265f
C324 VIN-.n8 GNDA 0.064892f
C325 VIN-.n9 GNDA 0.186141f
C326 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.028303f
C327 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.022556f
C328 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.607656f
C329 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.022403f
C330 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.022403f
C331 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.092646f
C332 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.022403f
C333 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.022403f
C334 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.09229f
C335 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.127961f
C336 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.022403f
C337 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.022403f
C338 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.09229f
C339 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.066772f
C340 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.022403f
C341 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.022403f
C342 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.09229f
C343 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.066772f
C344 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.022403f
C345 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.022403f
C346 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.09229f
C347 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.161141f
C348 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.619006f
C349 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.084125f
C350 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.09829f
C351 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.011144f
C352 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.018145f
C353 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.106108f
C354 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.021321f
C355 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.094664f
C356 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.011069f
C357 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.090853f
C358 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.021321f
C359 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.066102f
C360 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.021321f
C361 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.202731f
C362 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.098301f
C363 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.09227f
C364 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.515714f
C365 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 0.773533f
C366 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.325901f
C367 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.09227f
C368 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA 0.024781f
C369 two_stage_opamp_dummy_magic_0.V_p.n0 GNDA 0.049064f
C370 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA 0.014869f
C371 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA 0.014869f
C372 two_stage_opamp_dummy_magic_0.V_p.n1 GNDA 0.050516f
C373 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA 0.014869f
C374 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA 0.014869f
C375 two_stage_opamp_dummy_magic_0.V_p.n2 GNDA 0.053418f
C376 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA 0.014869f
C377 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA 0.014869f
C378 two_stage_opamp_dummy_magic_0.V_p.n3 GNDA 0.053005f
C379 two_stage_opamp_dummy_magic_0.V_p.n4 GNDA 0.179254f
C380 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA 0.014869f
C381 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA 0.014869f
C382 two_stage_opamp_dummy_magic_0.V_p.n5 GNDA 0.053005f
C383 two_stage_opamp_dummy_magic_0.V_p.n6 GNDA 0.093302f
C384 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA 0.014869f
C385 two_stage_opamp_dummy_magic_0.V_p.t4 GNDA 0.014869f
C386 two_stage_opamp_dummy_magic_0.V_p.n7 GNDA 0.053005f
C387 two_stage_opamp_dummy_magic_0.V_p.n8 GNDA 0.092807f
C388 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA 0.014869f
C389 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA 0.014869f
C390 two_stage_opamp_dummy_magic_0.V_p.n9 GNDA 0.053395f
C391 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA 0.014869f
C392 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA 0.014869f
C393 two_stage_opamp_dummy_magic_0.V_p.n10 GNDA 0.053005f
C394 two_stage_opamp_dummy_magic_0.V_p.n11 GNDA 0.177493f
C395 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA 0.014869f
C396 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA 0.014869f
C397 two_stage_opamp_dummy_magic_0.V_p.n12 GNDA 0.053005f
C398 two_stage_opamp_dummy_magic_0.V_p.n13 GNDA 0.093302f
C399 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA 0.014869f
C400 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA 0.014869f
C401 two_stage_opamp_dummy_magic_0.V_p.n14 GNDA 0.053005f
C402 two_stage_opamp_dummy_magic_0.V_p.n15 GNDA 0.093302f
C403 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA 0.014869f
C404 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA 0.014869f
C405 two_stage_opamp_dummy_magic_0.V_p.n16 GNDA 0.053005f
C406 two_stage_opamp_dummy_magic_0.V_p.n17 GNDA 0.142369f
C407 two_stage_opamp_dummy_magic_0.V_p.n18 GNDA 0.078308f
C408 two_stage_opamp_dummy_magic_0.V_p.n19 GNDA 0.0836f
C409 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA 0.024781f
C410 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA 0.024781f
C411 two_stage_opamp_dummy_magic_0.V_p.n20 GNDA 0.095622f
C412 two_stage_opamp_dummy_magic_0.V_p.n21 GNDA 0.079333f
C413 two_stage_opamp_dummy_magic_0.V_p.n22 GNDA 0.16901f
C414 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA 0.024781f
C415 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA 0.024781f
C416 two_stage_opamp_dummy_magic_0.V_p.n23 GNDA 0.098392f
C417 two_stage_opamp_dummy_magic_0.V_p.n24 GNDA 0.087962f
C418 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA 0.024781f
C419 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA 0.024781f
C420 two_stage_opamp_dummy_magic_0.V_p.n25 GNDA 0.098392f
C421 two_stage_opamp_dummy_magic_0.V_p.n26 GNDA 0.087962f
C422 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA 0.024781f
C423 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA 0.024781f
C424 two_stage_opamp_dummy_magic_0.V_p.n27 GNDA 0.098392f
C425 two_stage_opamp_dummy_magic_0.V_p.n28 GNDA 0.087962f
C426 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA 0.024781f
C427 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA 0.024781f
C428 two_stage_opamp_dummy_magic_0.V_p.n29 GNDA 0.098849f
C429 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA 0.024781f
C430 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA 0.024781f
C431 two_stage_opamp_dummy_magic_0.V_p.n30 GNDA 0.098392f
C432 two_stage_opamp_dummy_magic_0.V_p.n31 GNDA 0.168527f
C433 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA 0.024781f
C434 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA 0.024781f
C435 two_stage_opamp_dummy_magic_0.V_p.n32 GNDA 0.098392f
C436 two_stage_opamp_dummy_magic_0.V_p.n33 GNDA 0.087962f
C437 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA 0.086517f
C438 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA 0.024781f
C439 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA 0.024781f
C440 two_stage_opamp_dummy_magic_0.V_p.n34 GNDA 0.095622f
C441 two_stage_opamp_dummy_magic_0.V_p.n35 GNDA 0.572198f
C442 two_stage_opamp_dummy_magic_0.V_p.n36 GNDA 0.029737f
C443 two_stage_opamp_dummy_magic_0.V_p.n37 GNDA 0.087962f
C444 two_stage_opamp_dummy_magic_0.V_p.n38 GNDA 0.098392f
C445 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA 0.024781f
C446 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.02127f
C447 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020358f
C448 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020407f
C449 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021244f
C450 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.021116f
C451 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.299998f
C452 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.021116f
C453 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.156484f
C454 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.021116f
C455 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.190977f
C456 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.153542f
C457 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.133374f
C458 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.242929f
C459 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.02127f
C460 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020976f
C461 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.328367f
C462 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020976f
C463 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.180843f
C464 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.180843f
C465 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020976f
C466 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 1.30141f
C467 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.035528f
C468 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.035528f
C469 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.035528f
C470 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.122118f
C471 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.035528f
C472 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.035528f
C473 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.115851f
C474 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 1.06767f
C475 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.021316f
C476 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.021316f
C477 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.048768f
C478 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.021316f
C479 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.021316f
C480 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.048509f
C481 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.021316f
C482 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.021316f
C483 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.048509f
C484 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.021316f
C485 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.021316f
C486 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.048509f
C487 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.031975f
C488 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.058004f
C489 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.065898f
C490 two_stage_opamp_dummy_magic_0.Vb3.t30 GNDA 0.031975f
C491 two_stage_opamp_dummy_magic_0.Vb3.t37 GNDA 0.058004f
C492 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.065898f
C493 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.064006f
C494 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.801298f
C495 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.175861f
C496 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.175861f
C497 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.175861f
C498 two_stage_opamp_dummy_magic_0.Vb3.t31 GNDA 0.175861f
C499 two_stage_opamp_dummy_magic_0.Vb3.t36 GNDA 0.202942f
C500 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.164767f
C501 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.101253f
C502 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.101253f
C503 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.09481f
C504 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.175861f
C505 two_stage_opamp_dummy_magic_0.Vb3.t35 GNDA 0.175861f
C506 two_stage_opamp_dummy_magic_0.Vb3.t29 GNDA 0.175861f
C507 two_stage_opamp_dummy_magic_0.Vb3.t32 GNDA 0.175861f
C508 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.202942f
C509 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.164767f
C510 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.101253f
C511 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.101253f
C512 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.09481f
C513 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.077892f
C514 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.175861f
C515 two_stage_opamp_dummy_magic_0.Vb3.t34 GNDA 0.175861f
C516 two_stage_opamp_dummy_magic_0.Vb3.t39 GNDA 0.175861f
C517 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.175861f
C518 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.202942f
C519 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.164767f
C520 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.101253f
C521 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 0.101253f
C522 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.09481f
C523 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.175861f
C524 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.175861f
C525 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.175861f
C526 two_stage_opamp_dummy_magic_0.Vb3.t38 GNDA 0.175861f
C527 two_stage_opamp_dummy_magic_0.Vb3.t33 GNDA 0.202942f
C528 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.164767f
C529 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 0.101253f
C530 two_stage_opamp_dummy_magic_0.Vb3.n27 GNDA 0.101253f
C531 two_stage_opamp_dummy_magic_0.Vb3.n28 GNDA 0.09481f
C532 two_stage_opamp_dummy_magic_0.Vb3.n29 GNDA 0.057251f
C533 two_stage_opamp_dummy_magic_0.Vb3.n30 GNDA 1.78968f
C534 two_stage_opamp_dummy_magic_0.Vb3.n31 GNDA 4.75238f
C535 two_stage_opamp_dummy_magic_0.Vb3.n32 GNDA 3.71013f
C536 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.035528f
C537 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.035528f
C538 two_stage_opamp_dummy_magic_0.Vb3.n33 GNDA 0.122118f
C539 two_stage_opamp_dummy_magic_0.Vb3.n34 GNDA 1.06767f
C540 two_stage_opamp_dummy_magic_0.Vb3.n35 GNDA 0.115851f
C541 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.035528f
C542 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA 0.020233f
C543 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA 0.020233f
C544 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 GNDA 0.020233f
C545 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 GNDA 0.047731f
C546 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 GNDA 0.020233f
C547 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA 0.020233f
C548 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 GNDA 0.046922f
C549 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 GNDA 0.884615f
C550 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA 0.020233f
C551 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 GNDA 0.020233f
C552 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 GNDA 0.046922f
C553 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 GNDA 2.10658f
C554 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 GNDA 1.98101f
C555 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA 0.020233f
C556 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA 0.020233f
C557 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 GNDA 0.04777f
C558 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA 0.016692f
C559 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA 0.016692f
C560 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA 0.016692f
C561 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA 0.016692f
C562 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA 0.016692f
C563 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA 0.036166f
C564 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 GNDA 0.051623f
C565 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA 0.020233f
C566 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA 0.020233f
C567 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 GNDA 0.04777f
C568 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 GNDA 0.17992f
C569 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 GNDA 0.05811f
C570 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 GNDA 0.039231f
C571 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 GNDA 0.044006f
C572 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 GNDA 0.044006f
C573 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 GNDA 0.039231f
C574 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA 0.016692f
C575 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 GNDA 0.016692f
C576 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA 0.016692f
C577 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA 0.036166f
C578 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 GNDA 0.056399f
C579 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 GNDA 0.044006f
C580 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 GNDA 0.039231f
C581 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 GNDA 0.05811f
C582 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 GNDA 0.17992f
C583 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 GNDA 0.746838f
C584 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 GNDA 0.061393f
C585 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA 0.020233f
C586 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.03144f
C587 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.03144f
C588 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.10934f
C589 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.03144f
C590 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.03144f
C591 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.108953f
C592 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.205692f
C593 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.03144f
C594 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.03144f
C595 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.108953f
C596 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.106633f
C597 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.03144f
C598 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.03144f
C599 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.108953f
C600 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.106633f
C601 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.03144f
C602 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.03144f
C603 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.10934f
C604 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.127804f
C605 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.03144f
C606 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.03144f
C607 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.106696f
C608 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.089361f
C609 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.03144f
C610 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.03144f
C611 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.10934f
C612 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.03144f
C613 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.03144f
C614 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.108953f
C615 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.205693f
C616 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.089505f
C617 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.089505f
C618 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.362715f
C619 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.362715f
C620 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.541405f
C621 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.3126f
C622 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.3126f
C623 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.3126f
C624 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.3126f
C625 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.23445f
C626 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.155099f
C627 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.054747f
C628 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.101182f
C629 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.065226f
C630 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.155099f
C631 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.054747f
C632 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.101182f
C633 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.065226f
C634 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.064676f
C635 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.12171f
C636 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.541405f
C637 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.3126f
C638 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.3126f
C639 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.3126f
C640 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.3126f
C641 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.23445f
C642 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.1563f
C643 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.12171f
C644 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.125303f
C645 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.03144f
C646 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.03144f
C647 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.102506f
C648 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.074649f
C649 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.038431f
C650 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.03144f
C651 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.03144f
C652 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.108953f
C653 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.101243f
C654 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.03144f
C655 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.03144f
C656 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.1091f
C657 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.116136f
C658 ref_volt_cur_gen_dummy_magic_0.Vin+.t5 GNDA 0.125873f
C659 ref_volt_cur_gen_dummy_magic_0.Vin+.t9 GNDA 0.020459f
C660 ref_volt_cur_gen_dummy_magic_0.Vin+.t8 GNDA 0.013299f
C661 ref_volt_cur_gen_dummy_magic_0.Vin+.n0 GNDA 0.04388f
C662 ref_volt_cur_gen_dummy_magic_0.Vin+.t6 GNDA 0.013299f
C663 ref_volt_cur_gen_dummy_magic_0.Vin+.n1 GNDA 0.034146f
C664 ref_volt_cur_gen_dummy_magic_0.Vin+.t7 GNDA 0.013299f
C665 ref_volt_cur_gen_dummy_magic_0.Vin+.n2 GNDA 0.034607f
C666 ref_volt_cur_gen_dummy_magic_0.Vin+.n3 GNDA 0.074523f
C667 ref_volt_cur_gen_dummy_magic_0.Vin+.t4 GNDA 0.043132f
C668 ref_volt_cur_gen_dummy_magic_0.Vin+.t3 GNDA 0.043132f
C669 ref_volt_cur_gen_dummy_magic_0.Vin+.n4 GNDA 0.144858f
C670 ref_volt_cur_gen_dummy_magic_0.Vin+.t2 GNDA 0.043132f
C671 ref_volt_cur_gen_dummy_magic_0.Vin+.t1 GNDA 0.043132f
C672 ref_volt_cur_gen_dummy_magic_0.Vin+.n5 GNDA 0.142496f
C673 ref_volt_cur_gen_dummy_magic_0.Vin+.n6 GNDA 0.656763f
C674 ref_volt_cur_gen_dummy_magic_0.Vin+.n7 GNDA 0.71769f
C675 ref_volt_cur_gen_dummy_magic_0.Vin+.n8 GNDA 0.446219f
C676 ref_volt_cur_gen_dummy_magic_0.Vin+.t0 GNDA 0.137433f
C677 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.163765f
C678 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.409099f
C679 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.409099f
C680 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.485537f
C681 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.256456f
C682 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.162306f
C683 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.446073f
C684 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.149996f
C685 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.917914f
C686 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.446073f
C687 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.409099f
C688 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.409099f
C689 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.485537f
C690 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.256456f
C691 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.162306f
C692 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.149996f
C693 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.917423f
C694 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.163765f
C695 ref_volt_cur_gen_dummy_magic_0.START_UP.t4 GNDA 0.041701f
C696 ref_volt_cur_gen_dummy_magic_0.START_UP.t0 GNDA 1.6623f
C697 ref_volt_cur_gen_dummy_magic_0.START_UP.t1 GNDA 0.043697f
C698 ref_volt_cur_gen_dummy_magic_0.START_UP.n0 GNDA 1.28651f
C699 ref_volt_cur_gen_dummy_magic_0.START_UP.t6 GNDA 0.01567f
C700 ref_volt_cur_gen_dummy_magic_0.START_UP.t7 GNDA 0.01567f
C701 ref_volt_cur_gen_dummy_magic_0.START_UP.n1 GNDA 0.044238f
C702 ref_volt_cur_gen_dummy_magic_0.START_UP.n2 GNDA 0.853868f
C703 ref_volt_cur_gen_dummy_magic_0.START_UP.t3 GNDA 0.041701f
C704 ref_volt_cur_gen_dummy_magic_0.START_UP.t2 GNDA 0.041701f
C705 ref_volt_cur_gen_dummy_magic_0.START_UP.n3 GNDA 0.139173f
C706 ref_volt_cur_gen_dummy_magic_0.START_UP.n4 GNDA 0.720786f
C707 ref_volt_cur_gen_dummy_magic_0.START_UP.n5 GNDA 0.151283f
C708 ref_volt_cur_gen_dummy_magic_0.START_UP.t5 GNDA 0.041701f
C709 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.345114f
C710 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.346365f
C711 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.345114f
C712 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.34782f
C713 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.378304f
C714 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.345114f
C715 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.346365f
C716 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.345114f
C717 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.346365f
C718 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.345114f
C719 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.346365f
C720 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.345114f
C721 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.346365f
C722 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.345114f
C723 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.346365f
C724 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.345114f
C725 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.346365f
C726 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.345114f
C727 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.346365f
C728 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.345114f
C729 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.346365f
C730 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.345114f
C731 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.346365f
C732 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.345114f
C733 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.346365f
C734 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.345114f
C735 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.346365f
C736 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.345114f
C737 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.346365f
C738 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.345114f
C739 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.346365f
C740 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.345114f
C741 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.346365f
C742 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.345114f
C743 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.346365f
C744 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.345114f
C745 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.346365f
C746 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.345114f
C747 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.346365f
C748 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.345114f
C749 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.346365f
C750 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.345114f
C751 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.346365f
C752 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.345114f
C753 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.346365f
C754 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.345114f
C755 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.346365f
C756 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.345114f
C757 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.346365f
C758 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.345114f
C759 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.346365f
C760 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.345114f
C761 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.346365f
C762 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.345114f
C763 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.346365f
C764 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.345114f
C765 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.346365f
C766 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.345114f
C767 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.346365f
C768 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.345114f
C769 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.346365f
C770 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.345114f
C771 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.346365f
C772 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.345114f
C773 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.362035f
C774 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.345114f
C775 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.185368f
C776 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.198389f
C777 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.345114f
C778 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.185368f
C779 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.196789f
C780 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.345114f
C781 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.185368f
C782 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.196789f
C783 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.345114f
C784 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.185368f
C785 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.196789f
C786 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.345114f
C787 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.185368f
C788 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.196789f
C789 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.345114f
C790 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.185368f
C791 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.196789f
C792 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.345114f
C793 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.185368f
C794 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.196789f
C795 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.345114f
C796 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.185368f
C797 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196789f
C798 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.345114f
C799 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.185368f
C800 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196789f
C801 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.345114f
C802 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.346365f
C803 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.166846f
C804 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.215207f
C805 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.18422f
C806 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.233728f
C807 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.18422f
C808 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.250999f
C809 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.18422f
C810 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.250999f
C811 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.18422f
C812 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.250999f
C813 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.18422f
C814 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.250999f
C815 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.18422f
C816 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.250999f
C817 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.18422f
C818 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.250999f
C819 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.18422f
C820 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250999f
C821 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.18422f
C822 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250999f
C823 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.18422f
C824 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250999f
C825 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.18422f
C826 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250999f
C827 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.18422f
C828 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250999f
C829 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.18422f
C830 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250999f
C831 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.18422f
C832 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250999f
C833 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.18422f
C834 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250999f
C835 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.18422f
C836 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.233728f
C837 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.343967f
C838 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.166846f
C839 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.216458f
C840 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.343967f
C841 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.166846f
C842 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.216458f
C843 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.343967f
C844 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.345114f
C845 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.363635f
C846 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.363635f
C847 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.363635f
C848 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.185368f
C849 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.216458f
C850 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.343967f
C851 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.166846f
C852 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.197936f
C853 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.343967f
C854 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.166846f
C855 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.216458f
C856 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.343967f
C857 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.166846f
C858 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.216458f
C859 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.343967f
C860 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.166846f
C861 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216458f
C862 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.343967f
C863 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.345114f
C864 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.363635f
C865 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.363635f
C866 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.363635f
C867 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.185368f
C868 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216458f
C869 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.343967f
C870 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.345114f
C871 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.363635f
C872 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.363635f
C873 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.363635f
C874 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.185368f
C875 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216458f
C876 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.343967f
C877 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216458f
C878 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.185368f
C879 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.363635f
C880 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.363635f
C881 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.363635f
C882 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.602274f
C883 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.298233f
C884 VOUT+.t3 GNDA 0.043577f
C885 VOUT+.t14 GNDA 0.043577f
C886 VOUT+.n0 GNDA 0.175148f
C887 VOUT+.t9 GNDA 0.043577f
C888 VOUT+.t13 GNDA 0.043577f
C889 VOUT+.n1 GNDA 0.174825f
C890 VOUT+.n2 GNDA 0.172223f
C891 VOUT+.t8 GNDA 0.043577f
C892 VOUT+.t12 GNDA 0.043577f
C893 VOUT+.n3 GNDA 0.174825f
C894 VOUT+.n4 GNDA 0.088815f
C895 VOUT+.t6 GNDA 0.043577f
C896 VOUT+.t10 GNDA 0.043577f
C897 VOUT+.n5 GNDA 0.174825f
C898 VOUT+.n6 GNDA 0.088815f
C899 VOUT+.t5 GNDA 0.043577f
C900 VOUT+.t4 GNDA 0.043577f
C901 VOUT+.n7 GNDA 0.175148f
C902 VOUT+.n8 GNDA 0.105197f
C903 VOUT+.t7 GNDA 0.043577f
C904 VOUT+.t11 GNDA 0.043577f
C905 VOUT+.n9 GNDA 0.172685f
C906 VOUT+.n10 GNDA 0.210763f
C907 VOUT+.t117 GNDA 0.295461f
C908 VOUT+.t26 GNDA 0.290513f
C909 VOUT+.n11 GNDA 0.194779f
C910 VOUT+.t124 GNDA 0.290513f
C911 VOUT+.n12 GNDA 0.127099f
C912 VOUT+.t72 GNDA 0.295461f
C913 VOUT+.t39 GNDA 0.290513f
C914 VOUT+.n13 GNDA 0.194779f
C915 VOUT+.t127 GNDA 0.290513f
C916 VOUT+.t35 GNDA 0.294841f
C917 VOUT+.t87 GNDA 0.294841f
C918 VOUT+.t43 GNDA 0.294841f
C919 VOUT+.t96 GNDA 0.294841f
C920 VOUT+.t143 GNDA 0.294841f
C921 VOUT+.t106 GNDA 0.294841f
C922 VOUT+.t154 GNDA 0.294841f
C923 VOUT+.t65 GNDA 0.294841f
C924 VOUT+.t116 GNDA 0.294841f
C925 VOUT+.t73 GNDA 0.294841f
C926 VOUT+.t149 GNDA 0.290513f
C927 VOUT+.n14 GNDA 0.195399f
C928 VOUT+.t59 GNDA 0.290513f
C929 VOUT+.n15 GNDA 0.24987f
C930 VOUT+.t97 GNDA 0.290513f
C931 VOUT+.n16 GNDA 0.24987f
C932 VOUT+.t131 GNDA 0.290513f
C933 VOUT+.n17 GNDA 0.24987f
C934 VOUT+.t24 GNDA 0.290513f
C935 VOUT+.n18 GNDA 0.24987f
C936 VOUT+.t75 GNDA 0.290513f
C937 VOUT+.n19 GNDA 0.24987f
C938 VOUT+.t112 GNDA 0.290513f
C939 VOUT+.n20 GNDA 0.24987f
C940 VOUT+.t144 GNDA 0.290513f
C941 VOUT+.n21 GNDA 0.24987f
C942 VOUT+.t55 GNDA 0.290513f
C943 VOUT+.n22 GNDA 0.24987f
C944 VOUT+.t95 GNDA 0.290513f
C945 VOUT+.n23 GNDA 0.24987f
C946 VOUT+.n24 GNDA 0.236042f
C947 VOUT+.t38 GNDA 0.295461f
C948 VOUT+.t142 GNDA 0.290513f
C949 VOUT+.n25 GNDA 0.194779f
C950 VOUT+.t94 GNDA 0.290513f
C951 VOUT+.t20 GNDA 0.295461f
C952 VOUT+.t58 GNDA 0.290513f
C953 VOUT+.n26 GNDA 0.194779f
C954 VOUT+.n27 GNDA 0.236042f
C955 VOUT+.t80 GNDA 0.295461f
C956 VOUT+.t42 GNDA 0.290513f
C957 VOUT+.n28 GNDA 0.194779f
C958 VOUT+.t133 GNDA 0.290513f
C959 VOUT+.t61 GNDA 0.295461f
C960 VOUT+.t100 GNDA 0.290513f
C961 VOUT+.n29 GNDA 0.194779f
C962 VOUT+.n30 GNDA 0.236042f
C963 VOUT+.t121 GNDA 0.295461f
C964 VOUT+.t84 GNDA 0.290513f
C965 VOUT+.n31 GNDA 0.194779f
C966 VOUT+.t32 GNDA 0.290513f
C967 VOUT+.t104 GNDA 0.295461f
C968 VOUT+.t137 GNDA 0.290513f
C969 VOUT+.n32 GNDA 0.194779f
C970 VOUT+.n33 GNDA 0.236042f
C971 VOUT+.t85 GNDA 0.295461f
C972 VOUT+.t50 GNDA 0.290513f
C973 VOUT+.n34 GNDA 0.194779f
C974 VOUT+.t138 GNDA 0.290513f
C975 VOUT+.t67 GNDA 0.295461f
C976 VOUT+.t103 GNDA 0.290513f
C977 VOUT+.n35 GNDA 0.194779f
C978 VOUT+.n36 GNDA 0.236042f
C979 VOUT+.t123 GNDA 0.295461f
C980 VOUT+.t90 GNDA 0.290513f
C981 VOUT+.n37 GNDA 0.194779f
C982 VOUT+.t36 GNDA 0.290513f
C983 VOUT+.t107 GNDA 0.295337f
C984 VOUT+.t141 GNDA 0.290513f
C985 VOUT+.n38 GNDA 0.193087f
C986 VOUT+.n39 GNDA 0.236042f
C987 VOUT+.t108 GNDA 0.295461f
C988 VOUT+.t70 GNDA 0.290513f
C989 VOUT+.n40 GNDA 0.194779f
C990 VOUT+.t91 GNDA 0.290513f
C991 VOUT+.n41 GNDA 0.127099f
C992 VOUT+.t68 GNDA 0.295461f
C993 VOUT+.t31 GNDA 0.290513f
C994 VOUT+.n42 GNDA 0.194779f
C995 VOUT+.t52 GNDA 0.290513f
C996 VOUT+.t54 GNDA 0.294841f
C997 VOUT+.t156 GNDA 0.294841f
C998 VOUT+.t145 GNDA 0.295461f
C999 VOUT+.t45 GNDA 0.290513f
C1000 VOUT+.n43 GNDA 0.194779f
C1001 VOUT+.t136 GNDA 0.290513f
C1002 VOUT+.n44 GNDA 0.127099f
C1003 VOUT+.t101 GNDA 0.290513f
C1004 VOUT+.n45 GNDA 0.12256f
C1005 VOUT+.t37 GNDA 0.294841f
C1006 VOUT+.t113 GNDA 0.295461f
C1007 VOUT+.t151 GNDA 0.290513f
C1008 VOUT+.n46 GNDA 0.194779f
C1009 VOUT+.t98 GNDA 0.290513f
C1010 VOUT+.n47 GNDA 0.127099f
C1011 VOUT+.t60 GNDA 0.290513f
C1012 VOUT+.n48 GNDA 0.12256f
C1013 VOUT+.t140 GNDA 0.294841f
C1014 VOUT+.t76 GNDA 0.295461f
C1015 VOUT+.t118 GNDA 0.290513f
C1016 VOUT+.n49 GNDA 0.194779f
C1017 VOUT+.t57 GNDA 0.290513f
C1018 VOUT+.n50 GNDA 0.127099f
C1019 VOUT+.t21 GNDA 0.290513f
C1020 VOUT+.n51 GNDA 0.12256f
C1021 VOUT+.t105 GNDA 0.294841f
C1022 VOUT+.t25 GNDA 0.295461f
C1023 VOUT+.t66 GNDA 0.290513f
C1024 VOUT+.n52 GNDA 0.194779f
C1025 VOUT+.t81 GNDA 0.290513f
C1026 VOUT+.n53 GNDA 0.127099f
C1027 VOUT+.t44 GNDA 0.290513f
C1028 VOUT+.n54 GNDA 0.12256f
C1029 VOUT+.t125 GNDA 0.294841f
C1030 VOUT+.t88 GNDA 0.294841f
C1031 VOUT+.t51 GNDA 0.294841f
C1032 VOUT+.t150 GNDA 0.294841f
C1033 VOUT+.t33 GNDA 0.294841f
C1034 VOUT+.t134 GNDA 0.290513f
C1035 VOUT+.n55 GNDA 0.195399f
C1036 VOUT+.t110 GNDA 0.290513f
C1037 VOUT+.n56 GNDA 0.24987f
C1038 VOUT+.t147 GNDA 0.290513f
C1039 VOUT+.n57 GNDA 0.24987f
C1040 VOUT+.t46 GNDA 0.290513f
C1041 VOUT+.n58 GNDA 0.24987f
C1042 VOUT+.t86 GNDA 0.290513f
C1043 VOUT+.n59 GNDA 0.30888f
C1044 VOUT+.t62 GNDA 0.290513f
C1045 VOUT+.n60 GNDA 0.30888f
C1046 VOUT+.t102 GNDA 0.290513f
C1047 VOUT+.n61 GNDA 0.30888f
C1048 VOUT+.t139 GNDA 0.290513f
C1049 VOUT+.n62 GNDA 0.30888f
C1050 VOUT+.t119 GNDA 0.290513f
C1051 VOUT+.n63 GNDA 0.24987f
C1052 VOUT+.t155 GNDA 0.290513f
C1053 VOUT+.n64 GNDA 0.24987f
C1054 VOUT+.n65 GNDA 0.236042f
C1055 VOUT+.t28 GNDA 0.295461f
C1056 VOUT+.t130 GNDA 0.290513f
C1057 VOUT+.n66 GNDA 0.194779f
C1058 VOUT+.t152 GNDA 0.290513f
C1059 VOUT+.t77 GNDA 0.295461f
C1060 VOUT+.t115 GNDA 0.290513f
C1061 VOUT+.n67 GNDA 0.194779f
C1062 VOUT+.n68 GNDA 0.236042f
C1063 VOUT+.t63 GNDA 0.295461f
C1064 VOUT+.t23 GNDA 0.290513f
C1065 VOUT+.n69 GNDA 0.194779f
C1066 VOUT+.t48 GNDA 0.290513f
C1067 VOUT+.t111 GNDA 0.295461f
C1068 VOUT+.t148 GNDA 0.290513f
C1069 VOUT+.n70 GNDA 0.194779f
C1070 VOUT+.n71 GNDA 0.236042f
C1071 VOUT+.t114 GNDA 0.295461f
C1072 VOUT+.t79 GNDA 0.290513f
C1073 VOUT+.n72 GNDA 0.194779f
C1074 VOUT+.t27 GNDA 0.290513f
C1075 VOUT+.t99 GNDA 0.295461f
C1076 VOUT+.t132 GNDA 0.290513f
C1077 VOUT+.n73 GNDA 0.194779f
C1078 VOUT+.n74 GNDA 0.236042f
C1079 VOUT+.t74 GNDA 0.295461f
C1080 VOUT+.t40 GNDA 0.290513f
C1081 VOUT+.n75 GNDA 0.194779f
C1082 VOUT+.t128 GNDA 0.290513f
C1083 VOUT+.t56 GNDA 0.295461f
C1084 VOUT+.t93 GNDA 0.290513f
C1085 VOUT+.n76 GNDA 0.194779f
C1086 VOUT+.n77 GNDA 0.236042f
C1087 VOUT+.t109 GNDA 0.295461f
C1088 VOUT+.t71 GNDA 0.290513f
C1089 VOUT+.n78 GNDA 0.194779f
C1090 VOUT+.t19 GNDA 0.290513f
C1091 VOUT+.t92 GNDA 0.295461f
C1092 VOUT+.t126 GNDA 0.290513f
C1093 VOUT+.n79 GNDA 0.194779f
C1094 VOUT+.n80 GNDA 0.236042f
C1095 VOUT+.t69 GNDA 0.295461f
C1096 VOUT+.t34 GNDA 0.290513f
C1097 VOUT+.n81 GNDA 0.194779f
C1098 VOUT+.t122 GNDA 0.290513f
C1099 VOUT+.t53 GNDA 0.295461f
C1100 VOUT+.t89 GNDA 0.290513f
C1101 VOUT+.n82 GNDA 0.194779f
C1102 VOUT+.n83 GNDA 0.236042f
C1103 VOUT+.t30 GNDA 0.295461f
C1104 VOUT+.t135 GNDA 0.290513f
C1105 VOUT+.n84 GNDA 0.194779f
C1106 VOUT+.t83 GNDA 0.290513f
C1107 VOUT+.t153 GNDA 0.295461f
C1108 VOUT+.t49 GNDA 0.290513f
C1109 VOUT+.n85 GNDA 0.194779f
C1110 VOUT+.n86 GNDA 0.236042f
C1111 VOUT+.t64 GNDA 0.295461f
C1112 VOUT+.t29 GNDA 0.290513f
C1113 VOUT+.n87 GNDA 0.194779f
C1114 VOUT+.t120 GNDA 0.290513f
C1115 VOUT+.t47 GNDA 0.295461f
C1116 VOUT+.t82 GNDA 0.290513f
C1117 VOUT+.n88 GNDA 0.194779f
C1118 VOUT+.n89 GNDA 0.236042f
C1119 VOUT+.t22 GNDA 0.295461f
C1120 VOUT+.t129 GNDA 0.290513f
C1121 VOUT+.n90 GNDA 0.194779f
C1122 VOUT+.t78 GNDA 0.290513f
C1123 VOUT+.n91 GNDA 0.236042f
C1124 VOUT+.t41 GNDA 0.290513f
C1125 VOUT+.n92 GNDA 0.127099f
C1126 VOUT+.t146 GNDA 0.290513f
C1127 VOUT+.n93 GNDA 0.238016f
C1128 VOUT+.n94 GNDA 0.268648f
C1129 VOUT+.t15 GNDA 0.05084f
C1130 VOUT+.t17 GNDA 0.05084f
C1131 VOUT+.n95 GNDA 0.235187f
C1132 VOUT+.t1 GNDA 0.05084f
C1133 VOUT+.t0 GNDA 0.05084f
C1134 VOUT+.n96 GNDA 0.2344f
C1135 VOUT+.n97 GNDA 0.144847f
C1136 VOUT+.t18 GNDA 0.05084f
C1137 VOUT+.t16 GNDA 0.05084f
C1138 VOUT+.n98 GNDA 0.2344f
C1139 VOUT+.n99 GNDA 0.089159f
C1140 VOUT+.t2 GNDA 0.084056f
C1141 VOUT+.n100 GNDA 0.119121f
C1142 ref_volt_cur_gen_dummy_magic_0.V_TOP.t48 GNDA 0.134378f
C1143 ref_volt_cur_gen_dummy_magic_0.V_TOP.t15 GNDA 0.116612f
C1144 ref_volt_cur_gen_dummy_magic_0.V_TOP.t25 GNDA 0.116612f
C1145 ref_volt_cur_gen_dummy_magic_0.V_TOP.t30 GNDA 0.116612f
C1146 ref_volt_cur_gen_dummy_magic_0.V_TOP.t35 GNDA 0.116612f
C1147 ref_volt_cur_gen_dummy_magic_0.V_TOP.t17 GNDA 0.116612f
C1148 ref_volt_cur_gen_dummy_magic_0.V_TOP.t22 GNDA 0.116612f
C1149 ref_volt_cur_gen_dummy_magic_0.V_TOP.t31 GNDA 0.116612f
C1150 ref_volt_cur_gen_dummy_magic_0.V_TOP.t36 GNDA 0.116612f
C1151 ref_volt_cur_gen_dummy_magic_0.V_TOP.t40 GNDA 0.116612f
C1152 ref_volt_cur_gen_dummy_magic_0.V_TOP.t46 GNDA 0.116612f
C1153 ref_volt_cur_gen_dummy_magic_0.V_TOP.t24 GNDA 0.116612f
C1154 ref_volt_cur_gen_dummy_magic_0.V_TOP.t37 GNDA 0.116612f
C1155 ref_volt_cur_gen_dummy_magic_0.V_TOP.t42 GNDA 0.116612f
C1156 ref_volt_cur_gen_dummy_magic_0.V_TOP.t49 GNDA 0.116612f
C1157 ref_volt_cur_gen_dummy_magic_0.V_TOP.t16 GNDA 0.15244f
C1158 ref_volt_cur_gen_dummy_magic_0.V_TOP.n0 GNDA 0.085226f
C1159 ref_volt_cur_gen_dummy_magic_0.V_TOP.n1 GNDA 0.062193f
C1160 ref_volt_cur_gen_dummy_magic_0.V_TOP.n2 GNDA 0.062193f
C1161 ref_volt_cur_gen_dummy_magic_0.V_TOP.n3 GNDA 0.062193f
C1162 ref_volt_cur_gen_dummy_magic_0.V_TOP.n4 GNDA 0.062193f
C1163 ref_volt_cur_gen_dummy_magic_0.V_TOP.n5 GNDA 0.057996f
C1164 ref_volt_cur_gen_dummy_magic_0.V_TOP.t6 GNDA 0.149962f
C1165 ref_volt_cur_gen_dummy_magic_0.V_TOP.t13 GNDA 0.157893f
C1166 ref_volt_cur_gen_dummy_magic_0.V_TOP.t12 GNDA 0.011106f
C1167 ref_volt_cur_gen_dummy_magic_0.V_TOP.t4 GNDA 0.011106f
C1168 ref_volt_cur_gen_dummy_magic_0.V_TOP.n6 GNDA 0.027652f
C1169 ref_volt_cur_gen_dummy_magic_0.V_TOP.n7 GNDA 0.736743f
C1170 ref_volt_cur_gen_dummy_magic_0.V_TOP.t0 GNDA 0.011106f
C1171 ref_volt_cur_gen_dummy_magic_0.V_TOP.t3 GNDA 0.011106f
C1172 ref_volt_cur_gen_dummy_magic_0.V_TOP.n8 GNDA 0.027839f
C1173 ref_volt_cur_gen_dummy_magic_0.V_TOP.t2 GNDA 0.011106f
C1174 ref_volt_cur_gen_dummy_magic_0.V_TOP.t1 GNDA 0.011106f
C1175 ref_volt_cur_gen_dummy_magic_0.V_TOP.n9 GNDA 0.027652f
C1176 ref_volt_cur_gen_dummy_magic_0.V_TOP.n10 GNDA 0.256267f
C1177 ref_volt_cur_gen_dummy_magic_0.V_TOP.t10 GNDA 0.011106f
C1178 ref_volt_cur_gen_dummy_magic_0.V_TOP.t7 GNDA 0.011106f
C1179 ref_volt_cur_gen_dummy_magic_0.V_TOP.n11 GNDA 0.026785f
C1180 ref_volt_cur_gen_dummy_magic_0.V_TOP.n12 GNDA 0.155669f
C1181 ref_volt_cur_gen_dummy_magic_0.V_TOP.n13 GNDA 0.088847f
C1182 ref_volt_cur_gen_dummy_magic_0.V_TOP.t11 GNDA 0.011106f
C1183 ref_volt_cur_gen_dummy_magic_0.V_TOP.t8 GNDA 0.011106f
C1184 ref_volt_cur_gen_dummy_magic_0.V_TOP.n14 GNDA 0.027652f
C1185 ref_volt_cur_gen_dummy_magic_0.V_TOP.n15 GNDA 0.153374f
C1186 ref_volt_cur_gen_dummy_magic_0.V_TOP.t5 GNDA 0.011106f
C1187 ref_volt_cur_gen_dummy_magic_0.V_TOP.t9 GNDA 0.011106f
C1188 ref_volt_cur_gen_dummy_magic_0.V_TOP.n16 GNDA 0.027652f
C1189 ref_volt_cur_gen_dummy_magic_0.V_TOP.n17 GNDA 0.151915f
C1190 ref_volt_cur_gen_dummy_magic_0.V_TOP.n18 GNDA 0.333935f
C1191 ref_volt_cur_gen_dummy_magic_0.V_TOP.n19 GNDA 0.023499f
C1192 ref_volt_cur_gen_dummy_magic_0.V_TOP.n20 GNDA 0.057996f
C1193 ref_volt_cur_gen_dummy_magic_0.V_TOP.n21 GNDA 0.062193f
C1194 ref_volt_cur_gen_dummy_magic_0.V_TOP.n22 GNDA 0.062193f
C1195 ref_volt_cur_gen_dummy_magic_0.V_TOP.n23 GNDA 0.062193f
C1196 ref_volt_cur_gen_dummy_magic_0.V_TOP.n24 GNDA 0.062193f
C1197 ref_volt_cur_gen_dummy_magic_0.V_TOP.n25 GNDA 0.062193f
C1198 ref_volt_cur_gen_dummy_magic_0.V_TOP.n26 GNDA 0.062193f
C1199 ref_volt_cur_gen_dummy_magic_0.V_TOP.n27 GNDA 0.057996f
C1200 ref_volt_cur_gen_dummy_magic_0.V_TOP.t21 GNDA 0.444236f
C1201 ref_volt_cur_gen_dummy_magic_0.V_TOP.t29 GNDA 0.451802f
C1202 ref_volt_cur_gen_dummy_magic_0.V_TOP.t41 GNDA 0.444236f
C1203 ref_volt_cur_gen_dummy_magic_0.V_TOP.n28 GNDA 0.297846f
C1204 ref_volt_cur_gen_dummy_magic_0.V_TOP.t34 GNDA 0.444236f
C1205 ref_volt_cur_gen_dummy_magic_0.V_TOP.t20 GNDA 0.451802f
C1206 ref_volt_cur_gen_dummy_magic_0.V_TOP.t47 GNDA 0.444236f
C1207 ref_volt_cur_gen_dummy_magic_0.V_TOP.n29 GNDA 0.297846f
C1208 ref_volt_cur_gen_dummy_magic_0.V_TOP.n30 GNDA 0.277647f
C1209 ref_volt_cur_gen_dummy_magic_0.V_TOP.t39 GNDA 0.451802f
C1210 ref_volt_cur_gen_dummy_magic_0.V_TOP.t14 GNDA 0.444236f
C1211 ref_volt_cur_gen_dummy_magic_0.V_TOP.n31 GNDA 0.297846f
C1212 ref_volt_cur_gen_dummy_magic_0.V_TOP.t45 GNDA 0.444236f
C1213 ref_volt_cur_gen_dummy_magic_0.V_TOP.t26 GNDA 0.451802f
C1214 ref_volt_cur_gen_dummy_magic_0.V_TOP.t19 GNDA 0.444236f
C1215 ref_volt_cur_gen_dummy_magic_0.V_TOP.n32 GNDA 0.297846f
C1216 ref_volt_cur_gen_dummy_magic_0.V_TOP.n33 GNDA 0.360942f
C1217 ref_volt_cur_gen_dummy_magic_0.V_TOP.t28 GNDA 0.451802f
C1218 ref_volt_cur_gen_dummy_magic_0.V_TOP.t38 GNDA 0.444236f
C1219 ref_volt_cur_gen_dummy_magic_0.V_TOP.n34 GNDA 0.297846f
C1220 ref_volt_cur_gen_dummy_magic_0.V_TOP.t33 GNDA 0.444236f
C1221 ref_volt_cur_gen_dummy_magic_0.V_TOP.t18 GNDA 0.451802f
C1222 ref_volt_cur_gen_dummy_magic_0.V_TOP.t44 GNDA 0.444236f
C1223 ref_volt_cur_gen_dummy_magic_0.V_TOP.n35 GNDA 0.297846f
C1224 ref_volt_cur_gen_dummy_magic_0.V_TOP.n36 GNDA 0.360942f
C1225 ref_volt_cur_gen_dummy_magic_0.V_TOP.t43 GNDA 0.451802f
C1226 ref_volt_cur_gen_dummy_magic_0.V_TOP.t32 GNDA 0.444236f
C1227 ref_volt_cur_gen_dummy_magic_0.V_TOP.n37 GNDA 0.297846f
C1228 ref_volt_cur_gen_dummy_magic_0.V_TOP.t23 GNDA 0.444236f
C1229 ref_volt_cur_gen_dummy_magic_0.V_TOP.n38 GNDA 0.277647f
C1230 ref_volt_cur_gen_dummy_magic_0.V_TOP.t27 GNDA 0.444236f
C1231 ref_volt_cur_gen_dummy_magic_0.V_TOP.n39 GNDA 0.194353f
C1232 ref_volt_cur_gen_dummy_magic_0.V_TOP.n40 GNDA 0.859259f
C1233 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.020502f
C1234 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.016339f
C1235 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.127301f
C1236 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.06094f
C1237 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.016229f
C1238 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.016229f
C1239 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.067112f
C1240 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.016229f
C1241 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.016229f
C1242 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.066854f
C1243 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.092694f
C1244 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.016229f
C1245 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.016229f
C1246 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.066854f
C1247 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.048369f
C1248 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.016229f
C1249 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.016229f
C1250 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.066854f
C1251 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.048369f
C1252 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.016229f
C1253 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.016229f
C1254 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.066854f
C1255 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.116942f
C1256 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.660581f
C1257 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S4 GNDA 0.589511f
C1258 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.053187f
C1259 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.053187f
C1260 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.184972f
C1261 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.053187f
C1262 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.053187f
C1263 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.184316f
C1264 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.347971f
C1265 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.053187f
C1266 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.053187f
C1267 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.184316f
C1268 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.180392f
C1269 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.053187f
C1270 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.053187f
C1271 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.184316f
C1272 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.180392f
C1273 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.053187f
C1274 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.053187f
C1275 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.184316f
C1276 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.212415f
C1277 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.053187f
C1278 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.053187f
C1279 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.180498f
C1280 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.149147f
C1281 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.022794f
C1282 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.022794f
C1283 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.076959f
C1284 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.022794f
C1285 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.022794f
C1286 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.082252f
C1287 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.022794f
C1288 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.022794f
C1289 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.081534f
C1290 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.302737f
C1291 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.022794f
C1292 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.022794f
C1293 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.081534f
C1294 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.157046f
C1295 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.022794f
C1296 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.022794f
C1297 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.081534f
C1298 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.157046f
C1299 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.022794f
C1300 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.022794f
C1301 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.082252f
C1302 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.191279f
C1303 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.123631f
C1304 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.031912f
C1305 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.031912f
C1306 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.031912f
C1307 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.031912f
C1308 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.031912f
C1309 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.031912f
C1310 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.031912f
C1311 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.03875f
C1312 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.03875f
C1313 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.025074f
C1314 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.025074f
C1315 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.025074f
C1316 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.025074f
C1317 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.025074f
C1318 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.022459f
C1319 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.031912f
C1320 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.03875f
C1321 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.036135f
C1322 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.022101f
C1323 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.049008f
C1324 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.049008f
C1325 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.049008f
C1326 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.049008f
C1327 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.049008f
C1328 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.049008f
C1329 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.049008f
C1330 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.055713f
C1331 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.05028f
C1332 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.030772f
C1333 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.030772f
C1334 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.030772f
C1335 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.030772f
C1336 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.030772f
C1337 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.028157f
C1338 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.049008f
C1339 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.055713f
C1340 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.047665f
C1341 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.022031f
C1342 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.153015f
C1343 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.741299f
C1344 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.100295f
C1345 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.100295f
C1346 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.106821f
C1347 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.084651f
C1348 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.045253f
C1349 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.100295f
C1350 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.100295f
C1351 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.100295f
C1352 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.100295f
C1353 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.100295f
C1354 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.100295f
C1355 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.106821f
C1356 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.084651f
C1357 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.047868f
C1358 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.047868f
C1359 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.047868f
C1360 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.047868f
C1361 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.045253f
C1362 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.024415f
C1363 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 1.03694f
C1364 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.458663f
C1365 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.192021f
C1366 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.030665f
C1367 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.030665f
C1368 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.08997f
C1369 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.030665f
C1370 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.030665f
C1371 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.089561f
C1372 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.309576f
C1373 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.030665f
C1374 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.030665f
C1375 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.089561f
C1376 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.160359f
C1377 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.030665f
C1378 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.030665f
C1379 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.089561f
C1380 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.160359f
C1381 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.030665f
C1382 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.030665f
C1383 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.089561f
C1384 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.230381f
C1385 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 1.29517f
C1386 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.038331f
C1387 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.038331f
C1388 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.124528f
C1389 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.038331f
C1390 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.038331f
C1391 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.123627f
C1392 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.45876f
C1393 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.038331f
C1394 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.038331f
C1395 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.076663f
C1396 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 0.210234f
C1397 ref_volt_cur_gen_dummy_magic_0.V_CMFB_S1 GNDA 1.67347f
C1398 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.041329f
C1399 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.041329f
C1400 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.143735f
C1401 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.041329f
C1402 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.041329f
C1403 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.143225f
C1404 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.270395f
C1405 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.041329f
C1406 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.041329f
C1407 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.143225f
C1408 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.140175f
C1409 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.041329f
C1410 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.041329f
C1411 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.143225f
C1412 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.140175f
C1413 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.041329f
C1414 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.041329f
C1415 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.143225f
C1416 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.165059f
C1417 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.041329f
C1418 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.041329f
C1419 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.140258f
C1420 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.115897f
C1421 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.017712f
C1422 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.017712f
C1423 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.059802f
C1424 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.017712f
C1425 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.017712f
C1426 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.063915f
C1427 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.017712f
C1428 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.017712f
C1429 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.063915f
C1430 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.017712f
C1431 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.017712f
C1432 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.063357f
C1433 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.235245f
C1434 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.017712f
C1435 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.017712f
C1436 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.063357f
C1437 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.122034f
C1438 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.017712f
C1439 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.017712f
C1440 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.063357f
C1441 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.122034f
C1442 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.148636f
C1443 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.096069f
C1444 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.101103f
C1445 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.024798f
C1446 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.030111f
C1447 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.028079f
C1448 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.024798f
C1449 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.024798f
C1450 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.024798f
C1451 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.024798f
C1452 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.024798f
C1453 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.024798f
C1454 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.024798f
C1455 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.030111f
C1456 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.030111f
C1457 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.019484f
C1458 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.019484f
C1459 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.019484f
C1460 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.019484f
C1461 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.019484f
C1462 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.017452f
C1463 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.017174f
C1464 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.038082f
C1465 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.043293f
C1466 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.037039f
C1467 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.038082f
C1468 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.038082f
C1469 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.038082f
C1470 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.038082f
C1471 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.038082f
C1472 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.038082f
C1473 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.038082f
C1474 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.043293f
C1475 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.039071f
C1476 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.023912f
C1477 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.023912f
C1478 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.023912f
C1479 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.023912f
C1480 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.023912f
C1481 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.02188f
C1482 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.01712f
C1483 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.120237f
C1484 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.357276f
C1485 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.077935f
C1486 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.077935f
C1487 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.077935f
C1488 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.077935f
C1489 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.077935f
C1490 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.077935f
C1491 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.083006f
C1492 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.065779f
C1493 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.037196f
C1494 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.037196f
C1495 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.037196f
C1496 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.037196f
C1497 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.035164f
C1498 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.077935f
C1499 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.077935f
C1500 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.083006f
C1501 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.065779f
C1502 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.035164f
C1503 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.019054f
C1504 two_stage_opamp_dummy_magic_0.X.n52 GNDA 0.811703f
C1505 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.576893f
C1506 ref_volt_cur_gen_dummy_magic_0.V_mir1.t11 GNDA 0.03537f
C1507 ref_volt_cur_gen_dummy_magic_0.V_mir1.t7 GNDA 0.03537f
C1508 ref_volt_cur_gen_dummy_magic_0.V_mir1.n0 GNDA 0.08097f
C1509 ref_volt_cur_gen_dummy_magic_0.V_mir1.t10 GNDA 0.042444f
C1510 ref_volt_cur_gen_dummy_magic_0.V_mir1.t18 GNDA 0.042444f
C1511 ref_volt_cur_gen_dummy_magic_0.V_mir1.t17 GNDA 0.06851f
C1512 ref_volt_cur_gen_dummy_magic_0.V_mir1.n1 GNDA 0.076506f
C1513 ref_volt_cur_gen_dummy_magic_0.V_mir1.n2 GNDA 0.052264f
C1514 ref_volt_cur_gen_dummy_magic_0.V_mir1.t6 GNDA 0.053881f
C1515 ref_volt_cur_gen_dummy_magic_0.V_mir1.n3 GNDA 0.081315f
C1516 ref_volt_cur_gen_dummy_magic_0.V_mir1.n4 GNDA 0.201563f
C1517 ref_volt_cur_gen_dummy_magic_0.V_mir1.t9 GNDA 0.03537f
C1518 ref_volt_cur_gen_dummy_magic_0.V_mir1.t5 GNDA 0.03537f
C1519 ref_volt_cur_gen_dummy_magic_0.V_mir1.n5 GNDA 0.08097f
C1520 ref_volt_cur_gen_dummy_magic_0.V_mir1.t8 GNDA 0.042444f
C1521 ref_volt_cur_gen_dummy_magic_0.V_mir1.t20 GNDA 0.042444f
C1522 ref_volt_cur_gen_dummy_magic_0.V_mir1.t22 GNDA 0.06851f
C1523 ref_volt_cur_gen_dummy_magic_0.V_mir1.n6 GNDA 0.076506f
C1524 ref_volt_cur_gen_dummy_magic_0.V_mir1.n7 GNDA 0.052264f
C1525 ref_volt_cur_gen_dummy_magic_0.V_mir1.t4 GNDA 0.053881f
C1526 ref_volt_cur_gen_dummy_magic_0.V_mir1.n8 GNDA 0.081315f
C1527 ref_volt_cur_gen_dummy_magic_0.V_mir1.n9 GNDA 0.156007f
C1528 ref_volt_cur_gen_dummy_magic_0.V_mir1.t16 GNDA 0.017685f
C1529 ref_volt_cur_gen_dummy_magic_0.V_mir1.t0 GNDA 0.017685f
C1530 ref_volt_cur_gen_dummy_magic_0.V_mir1.n10 GNDA 0.046242f
C1531 ref_volt_cur_gen_dummy_magic_0.V_mir1.t3 GNDA 0.075466f
C1532 ref_volt_cur_gen_dummy_magic_0.V_mir1.t1 GNDA 0.017685f
C1533 ref_volt_cur_gen_dummy_magic_0.V_mir1.t2 GNDA 0.017685f
C1534 ref_volt_cur_gen_dummy_magic_0.V_mir1.n11 GNDA 0.050199f
C1535 ref_volt_cur_gen_dummy_magic_0.V_mir1.n12 GNDA 0.827814f
C1536 ref_volt_cur_gen_dummy_magic_0.V_mir1.n13 GNDA 0.268286f
C1537 ref_volt_cur_gen_dummy_magic_0.V_mir1.n14 GNDA 0.09373f
C1538 ref_volt_cur_gen_dummy_magic_0.V_mir1.n15 GNDA 0.699157f
C1539 ref_volt_cur_gen_dummy_magic_0.V_mir1.t14 GNDA 0.042444f
C1540 ref_volt_cur_gen_dummy_magic_0.V_mir1.t21 GNDA 0.042444f
C1541 ref_volt_cur_gen_dummy_magic_0.V_mir1.t19 GNDA 0.06851f
C1542 ref_volt_cur_gen_dummy_magic_0.V_mir1.n16 GNDA 0.076506f
C1543 ref_volt_cur_gen_dummy_magic_0.V_mir1.n17 GNDA 0.052264f
C1544 ref_volt_cur_gen_dummy_magic_0.V_mir1.t12 GNDA 0.053881f
C1545 ref_volt_cur_gen_dummy_magic_0.V_mir1.n18 GNDA 0.081315f
C1546 ref_volt_cur_gen_dummy_magic_0.V_mir1.n19 GNDA 0.203577f
C1547 ref_volt_cur_gen_dummy_magic_0.V_mir1.t13 GNDA 0.03537f
C1548 ref_volt_cur_gen_dummy_magic_0.V_mir1.n20 GNDA 0.08097f
C1549 ref_volt_cur_gen_dummy_magic_0.V_mir1.t15 GNDA 0.03537f
C1550 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 0.802776f
C1551 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 0.777013f
C1552 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 5.29905f
C1553 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.045581f
C1554 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.045581f
C1555 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.143682f
C1556 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.022791f
C1557 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.022791f
C1558 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.052798f
C1559 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.022791f
C1560 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.022791f
C1561 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.052854f
C1562 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.018802f
C1563 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.018802f
C1564 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.018802f
C1565 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.018802f
C1566 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.018802f
C1567 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.018802f
C1568 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.018802f
C1569 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.018802f
C1570 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.018802f
C1571 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.018802f
C1572 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.018802f
C1573 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.018802f
C1574 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.018802f
C1575 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.018802f
C1576 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.018802f
C1577 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.018802f
C1578 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.040738f
C1579 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.063528f
C1580 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.049569f
C1581 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.049569f
C1582 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.049569f
C1583 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.049569f
C1584 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.049569f
C1585 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.049569f
C1586 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.049569f
C1587 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.049569f
C1588 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.049569f
C1589 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.049569f
C1590 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.049569f
C1591 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.049569f
C1592 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.049569f
C1593 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.049569f
C1594 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.042418f
C1595 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.018802f
C1596 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.018802f
C1597 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.040738f
C1598 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.063528f
C1599 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.042418f
C1600 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.06835f
C1601 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.022791f
C1602 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.022791f
C1603 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.045581f
C1604 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.135775f
C1605 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.022791f
C1606 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.022791f
C1607 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.052854f
C1608 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.022791f
C1609 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.022791f
C1610 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.052854f
C1611 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.022791f
C1612 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.022791f
C1613 two_stage_opamp_dummy_magic_0.V_err_gate.n29 GNDA 0.052854f
C1614 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.040476f
C1615 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.012714f
C1616 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.023725f
C1617 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.056644f
C1618 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.354182f
C1619 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.012714f
C1620 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.023725f
C1621 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.056644f
C1622 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.327181f
C1623 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.040089f
C1624 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.318577f
C1625 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.012714f
C1626 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.023725f
C1627 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 0.056644f
C1628 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.197826f
C1629 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.012714f
C1630 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.023725f
C1631 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.056644f
C1632 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.307478f
C1633 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.069261f
C1634 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.025899f
C1635 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 0.081234f
C1636 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.025899f
C1637 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.066497f
C1638 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.025899f
C1639 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.066497f
C1640 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.025899f
C1641 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.102019f
C1642 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.661388f
C1643 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.083997f
C1644 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.083997f
C1645 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.281474f
C1646 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 3.17158f
C1647 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.083997f
C1648 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.083997f
C1649 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.281474f
C1650 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.760085f
C1651 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.083997f
C1652 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.083997f
C1653 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.281474f
C1654 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 1.08667f
C1655 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.945272f
C1656 ref_volt_cur_gen_dummy_magic_0.cap_res1.t7 GNDA 0.412521f
C1657 ref_volt_cur_gen_dummy_magic_0.cap_res1.t2 GNDA 0.414016f
C1658 ref_volt_cur_gen_dummy_magic_0.cap_res1.t5 GNDA 0.412521f
C1659 ref_volt_cur_gen_dummy_magic_0.cap_res1.t8 GNDA 0.414016f
C1660 ref_volt_cur_gen_dummy_magic_0.cap_res1.t1 GNDA 0.412521f
C1661 ref_volt_cur_gen_dummy_magic_0.cap_res1.t14 GNDA 0.414016f
C1662 ref_volt_cur_gen_dummy_magic_0.cap_res1.t17 GNDA 0.412521f
C1663 ref_volt_cur_gen_dummy_magic_0.cap_res1.t4 GNDA 0.414016f
C1664 ref_volt_cur_gen_dummy_magic_0.cap_res1.t13 GNDA 0.412521f
C1665 ref_volt_cur_gen_dummy_magic_0.cap_res1.t9 GNDA 0.414016f
C1666 ref_volt_cur_gen_dummy_magic_0.cap_res1.t10 GNDA 0.412521f
C1667 ref_volt_cur_gen_dummy_magic_0.cap_res1.t16 GNDA 0.414016f
C1668 ref_volt_cur_gen_dummy_magic_0.cap_res1.t0 GNDA 0.412521f
C1669 ref_volt_cur_gen_dummy_magic_0.cap_res1.t12 GNDA 0.414016f
C1670 ref_volt_cur_gen_dummy_magic_0.cap_res1.t15 GNDA 0.412521f
C1671 ref_volt_cur_gen_dummy_magic_0.cap_res1.t3 GNDA 0.414016f
C1672 ref_volt_cur_gen_dummy_magic_0.cap_res1.n0 GNDA 0.276513f
C1673 ref_volt_cur_gen_dummy_magic_0.cap_res1.t18 GNDA 0.220202f
C1674 ref_volt_cur_gen_dummy_magic_0.cap_res1.n1 GNDA 0.300024f
C1675 ref_volt_cur_gen_dummy_magic_0.cap_res1.t11 GNDA 0.220202f
C1676 ref_volt_cur_gen_dummy_magic_0.cap_res1.n2 GNDA 0.300024f
C1677 ref_volt_cur_gen_dummy_magic_0.cap_res1.t19 GNDA 0.220202f
C1678 ref_volt_cur_gen_dummy_magic_0.cap_res1.n3 GNDA 0.300024f
C1679 ref_volt_cur_gen_dummy_magic_0.cap_res1.t6 GNDA 0.644091f
C1680 ref_volt_cur_gen_dummy_magic_0.cap_res1.t20 GNDA 0.106417f
C1681 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n0 GNDA 0.551826f
C1682 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n1 GNDA 0.283818f
C1683 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n2 GNDA 1.41958f
C1684 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n3 GNDA 1.86939f
C1685 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n4 GNDA 0.124721f
C1686 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n5 GNDA 0.012445f
C1687 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t0 GNDA 0.018146f
C1688 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n6 GNDA 0.188238f
C1689 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n7 GNDA 0.01126f
C1690 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t27 GNDA 0.020677f
C1691 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n8 GNDA 0.021718f
C1692 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t24 GNDA 0.013124f
C1693 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t29 GNDA 0.013124f
C1694 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n9 GNDA 0.029197f
C1695 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t25 GNDA 0.344612f
C1696 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t36 GNDA 0.350481f
C1697 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t18 GNDA 0.344612f
C1698 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t12 GNDA 0.344612f
C1699 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t15 GNDA 0.350481f
C1700 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t33 GNDA 0.344612f
C1701 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t17 GNDA 0.350481f
C1702 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t22 GNDA 0.344612f
C1703 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t19 GNDA 0.344612f
C1704 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t21 GNDA 0.350481f
C1705 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t14 GNDA 0.344612f
C1706 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t35 GNDA 0.350481f
C1707 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t16 GNDA 0.344612f
C1708 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t11 GNDA 0.344612f
C1709 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t13 GNDA 0.350481f
C1710 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t32 GNDA 0.344612f
C1711 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t31 GNDA 0.350481f
C1712 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t23 GNDA 0.344612f
C1713 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t28 GNDA 0.344612f
C1714 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t34 GNDA 0.344612f
C1715 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t20 GNDA 0.022513f
C1716 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n10 GNDA 0.021718f
C1717 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t26 GNDA 0.013124f
C1718 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.t30 GNDA 0.013124f
C1719 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n11 GNDA 0.029197f
C1720 ref_volt_cur_gen_dummy_magic_0.1st_Vout_1.n12 GNDA 0.020817f
C1721 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.030518f
C1722 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.030518f
C1723 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.030518f
C1724 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.110443f
C1725 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.020346f
C1726 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.020346f
C1727 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.051185f
C1728 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.020346f
C1729 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.020346f
C1730 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.050658f
C1731 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.386452f
C1732 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.020346f
C1733 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.020346f
C1734 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.050658f
C1735 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.25767f
C1736 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.020346f
C1737 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.020346f
C1738 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.049069f
C1739 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 1.95751f
C1740 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 2.30946f
C1741 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.05417f
C1742 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.05417f
C1743 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.05417f
C1744 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.05417f
C1745 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.05417f
C1746 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.05417f
C1747 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.05417f
C1748 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.063225f
C1749 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.059611f
C1750 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.037385f
C1751 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.037385f
C1752 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.037385f
C1753 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.037385f
C1754 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.037385f
C1755 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.033407f
C1756 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.05417f
C1757 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.05417f
C1758 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.05417f
C1759 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.05417f
C1760 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.05417f
C1761 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.05417f
C1762 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.05417f
C1763 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.05417f
C1764 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.05417f
C1765 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.05417f
C1766 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.05417f
C1767 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.063225f
C1768 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.059611f
C1769 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.037385f
C1770 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.037385f
C1771 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.037385f
C1772 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.037385f
C1773 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.037385f
C1774 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.037385f
C1775 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.037385f
C1776 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.037385f
C1777 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.037385f
C1778 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.033407f
C1779 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.083487f
C1780 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.236591f
C1781 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 0.061037f
C1782 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.030518f
C1783 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t17 GNDA 0.170605f
C1784 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t20 GNDA 0.170605f
C1785 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n0 GNDA 0.175172f
C1786 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t18 GNDA 0.332067f
C1787 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t14 GNDA 0.449269f
C1788 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n1 GNDA 0.239778f
C1789 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t22 GNDA 0.332067f
C1790 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t26 GNDA 0.449269f
C1791 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n2 GNDA 0.239778f
C1792 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n3 GNDA 0.091338f
C1793 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t19 GNDA 0.332067f
C1794 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t15 GNDA 0.449269f
C1795 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n4 GNDA 0.239778f
C1796 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t23 GNDA 0.332067f
C1797 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t11 GNDA 0.449269f
C1798 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n5 GNDA 0.239778f
C1799 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n6 GNDA 0.107586f
C1800 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n7 GNDA 1.37913f
C1801 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t13 GNDA 0.115501f
C1802 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t12 GNDA 0.115501f
C1803 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t25 GNDA 0.115501f
C1804 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t21 GNDA 0.204279f
C1805 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n8 GNDA 0.138375f
C1806 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n9 GNDA 0.119352f
C1807 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n10 GNDA 0.09577f
C1808 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t24 GNDA 0.115501f
C1809 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t27 GNDA 0.115501f
C1810 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t29 GNDA 0.115501f
C1811 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t10 GNDA 0.115501f
C1812 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t16 GNDA 0.115501f
C1813 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t28 GNDA 0.204279f
C1814 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n11 GNDA 0.138375f
C1815 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n12 GNDA 0.119352f
C1816 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n13 GNDA 0.09577f
C1817 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n14 GNDA 0.125716f
C1818 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n15 GNDA 0.09577f
C1819 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n16 GNDA 0.09577f
C1820 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n17 GNDA 0.125716f
C1821 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n18 GNDA 0.587506f
C1822 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n19 GNDA 1.51155f
C1823 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n20 GNDA 1.75217f
C1824 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t0 GNDA 0.0385f
C1825 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t5 GNDA 0.0385f
C1826 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n21 GNDA 0.098404f
C1827 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t9 GNDA 0.0385f
C1828 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t7 GNDA 0.0385f
C1829 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n22 GNDA 0.095862f
C1830 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n23 GNDA 0.937648f
C1831 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t8 GNDA 0.0385f
C1832 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t6 GNDA 0.0385f
C1833 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n24 GNDA 0.095862f
C1834 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n25 GNDA 0.531696f
C1835 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t2 GNDA 0.562397f
C1836 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n26 GNDA 1.08542f
C1837 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t4 GNDA 0.0385f
C1838 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t1 GNDA 0.0385f
C1839 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n27 GNDA 0.092855f
C1840 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n28 GNDA 0.341746f
C1841 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.n29 GNDA 3.68874f
C1842 ref_volt_cur_gen_dummy_magic_0.PFET_GATE_10uA.t3 GNDA 0.748699f
C1843 ref_volt_cur_gen_dummy_magic_0.cap_res2.t7 GNDA 0.401569f
C1844 ref_volt_cur_gen_dummy_magic_0.cap_res2.t2 GNDA 0.403025f
C1845 ref_volt_cur_gen_dummy_magic_0.cap_res2.t14 GNDA 0.401569f
C1846 ref_volt_cur_gen_dummy_magic_0.cap_res2.t13 GNDA 0.403025f
C1847 ref_volt_cur_gen_dummy_magic_0.cap_res2.t1 GNDA 0.401569f
C1848 ref_volt_cur_gen_dummy_magic_0.cap_res2.t17 GNDA 0.403025f
C1849 ref_volt_cur_gen_dummy_magic_0.cap_res2.t9 GNDA 0.401569f
C1850 ref_volt_cur_gen_dummy_magic_0.cap_res2.t6 GNDA 0.403025f
C1851 ref_volt_cur_gen_dummy_magic_0.cap_res2.t16 GNDA 0.401569f
C1852 ref_volt_cur_gen_dummy_magic_0.cap_res2.t11 GNDA 0.403025f
C1853 ref_volt_cur_gen_dummy_magic_0.cap_res2.t3 GNDA 0.401569f
C1854 ref_volt_cur_gen_dummy_magic_0.cap_res2.t19 GNDA 0.403025f
C1855 ref_volt_cur_gen_dummy_magic_0.cap_res2.t20 GNDA 0.401569f
C1856 ref_volt_cur_gen_dummy_magic_0.cap_res2.t15 GNDA 0.403025f
C1857 ref_volt_cur_gen_dummy_magic_0.cap_res2.t8 GNDA 0.401569f
C1858 ref_volt_cur_gen_dummy_magic_0.cap_res2.t4 GNDA 0.403025f
C1859 ref_volt_cur_gen_dummy_magic_0.cap_res2.n0 GNDA 0.269172f
C1860 ref_volt_cur_gen_dummy_magic_0.cap_res2.t10 GNDA 0.214356f
C1861 ref_volt_cur_gen_dummy_magic_0.cap_res2.n1 GNDA 0.292058f
C1862 ref_volt_cur_gen_dummy_magic_0.cap_res2.t5 GNDA 0.214356f
C1863 ref_volt_cur_gen_dummy_magic_0.cap_res2.n2 GNDA 0.292058f
C1864 ref_volt_cur_gen_dummy_magic_0.cap_res2.t12 GNDA 0.214356f
C1865 ref_volt_cur_gen_dummy_magic_0.cap_res2.n3 GNDA 0.292058f
C1866 ref_volt_cur_gen_dummy_magic_0.cap_res2.t18 GNDA 0.840875f
C1867 ref_volt_cur_gen_dummy_magic_0.cap_res2.t0 GNDA 0.133954f
C1868 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.344645f
C1869 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.167175f
C1870 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.198327f
C1871 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.344645f
C1872 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.167175f
C1873 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.216884f
C1874 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.344645f
C1875 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.167175f
C1876 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.216884f
C1877 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.344645f
C1878 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.167175f
C1879 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.216884f
C1880 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344645f
C1881 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.345795f
C1882 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.364353f
C1883 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.364353f
C1884 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.364353f
C1885 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.185733f
C1886 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.216884f
C1887 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344645f
C1888 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.345795f
C1889 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.364353f
C1890 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.364353f
C1891 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.364353f
C1892 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.185733f
C1893 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.216884f
C1894 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345795f
C1895 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.347048f
C1896 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345795f
C1897 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.348506f
C1898 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.37905f
C1899 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.345795f
C1900 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.347048f
C1901 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.345795f
C1902 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.347048f
C1903 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.345795f
C1904 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.347048f
C1905 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.345795f
C1906 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.347048f
C1907 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.345795f
C1908 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.347048f
C1909 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.345795f
C1910 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.347048f
C1911 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.345795f
C1912 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.347048f
C1913 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.345795f
C1914 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.347048f
C1915 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345795f
C1916 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.347048f
C1917 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.345795f
C1918 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.347048f
C1919 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.345795f
C1920 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.347048f
C1921 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.345795f
C1922 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.347048f
C1923 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.345795f
C1924 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.347048f
C1925 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.345795f
C1926 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.347048f
C1927 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.345795f
C1928 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.347048f
C1929 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.345795f
C1930 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.347048f
C1931 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.345795f
C1932 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.347048f
C1933 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.345795f
C1934 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.347048f
C1935 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.345795f
C1936 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.347048f
C1937 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.345795f
C1938 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.347048f
C1939 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.345795f
C1940 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.347048f
C1941 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.345795f
C1942 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.347048f
C1943 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.345795f
C1944 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.347048f
C1945 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.345795f
C1946 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.347048f
C1947 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.345795f
C1948 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.347048f
C1949 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.345795f
C1950 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.347048f
C1951 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.345795f
C1952 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.347048f
C1953 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.345795f
C1954 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.347048f
C1955 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.345795f
C1956 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.362749f
C1957 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.345795f
C1958 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.185733f
C1959 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.198781f
C1960 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.345795f
C1961 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.185733f
C1962 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.197177f
C1963 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.345795f
C1964 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.185733f
C1965 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.197177f
C1966 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.345795f
C1967 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.185733f
C1968 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.197177f
C1969 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.345795f
C1970 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185733f
C1971 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.197177f
C1972 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.345795f
C1973 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.185733f
C1974 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.197177f
C1975 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.345795f
C1976 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.185733f
C1977 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.197177f
C1978 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.345795f
C1979 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.185733f
C1980 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.197177f
C1981 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.345795f
C1982 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185733f
C1983 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.197177f
C1984 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.345795f
C1985 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.347048f
C1986 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.345795f
C1987 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.347048f
C1988 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.167175f
C1989 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.215631f
C1990 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.184584f
C1991 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.234189f
C1992 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.184584f
C1993 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.251494f
C1994 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.184584f
C1995 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.251494f
C1996 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.184584f
C1997 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.251494f
C1998 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.184584f
C1999 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.251494f
C2000 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.184584f
C2001 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.251494f
C2002 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.184584f
C2003 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.251494f
C2004 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.184584f
C2005 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.251494f
C2006 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.184584f
C2007 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.251494f
C2008 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.184584f
C2009 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.251494f
C2010 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.184584f
C2011 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.251494f
C2012 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.184584f
C2013 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.251494f
C2014 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.184584f
C2015 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.251494f
C2016 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.184584f
C2017 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.251494f
C2018 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.184584f
C2019 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.251494f
C2020 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.184584f
C2021 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.234189f
C2022 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.344645f
C2023 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.167175f
C2024 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216884f
C2025 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C2026 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.167175f
C2027 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216884f
C2028 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344645f
C2029 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.345795f
C2030 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.364353f
C2031 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.364353f
C2032 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.364353f
C2033 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185733f
C2034 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216884f
C2035 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.344645f
C2036 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216884f
C2037 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185733f
C2038 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.364353f
C2039 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.364353f
C2040 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.364353f
C2041 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.337351f
C2042 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.298183f
C2043 VOUT-.t18 GNDA 0.049273f
C2044 VOUT-.t0 GNDA 0.049273f
C2045 VOUT-.n0 GNDA 0.227938f
C2046 VOUT-.t1 GNDA 0.049273f
C2047 VOUT-.t11 GNDA 0.049273f
C2048 VOUT-.n1 GNDA 0.227175f
C2049 VOUT-.n2 GNDA 0.140383f
C2050 VOUT-.t12 GNDA 0.049273f
C2051 VOUT-.t17 GNDA 0.049273f
C2052 VOUT-.n3 GNDA 0.227175f
C2053 VOUT-.n4 GNDA 0.086411f
C2054 VOUT-.t7 GNDA 0.081465f
C2055 VOUT-.n5 GNDA 0.11545f
C2056 VOUT-.t9 GNDA 0.042234f
C2057 VOUT-.t4 GNDA 0.042234f
C2058 VOUT-.n6 GNDA 0.16975f
C2059 VOUT-.t5 GNDA 0.042234f
C2060 VOUT-.t10 GNDA 0.042234f
C2061 VOUT-.n7 GNDA 0.169749f
C2062 VOUT-.t13 GNDA 0.042234f
C2063 VOUT-.t3 GNDA 0.042234f
C2064 VOUT-.n8 GNDA 0.169437f
C2065 VOUT-.n9 GNDA 0.166915f
C2066 VOUT-.t15 GNDA 0.042234f
C2067 VOUT-.t16 GNDA 0.042234f
C2068 VOUT-.n10 GNDA 0.169437f
C2069 VOUT-.n11 GNDA 0.086077f
C2070 VOUT-.t8 GNDA 0.042234f
C2071 VOUT-.t6 GNDA 0.042234f
C2072 VOUT-.n12 GNDA 0.169437f
C2073 VOUT-.n13 GNDA 0.086077f
C2074 VOUT-.n14 GNDA 0.101954f
C2075 VOUT-.t2 GNDA 0.042234f
C2076 VOUT-.t14 GNDA 0.042234f
C2077 VOUT-.n15 GNDA 0.167363f
C2078 VOUT-.n16 GNDA 0.205258f
C2079 VOUT-.t100 GNDA 0.281558f
C2080 VOUT-.t107 GNDA 0.286354f
C2081 VOUT-.t149 GNDA 0.281558f
C2082 VOUT-.n17 GNDA 0.188776f
C2083 VOUT-.n18 GNDA 0.123182f
C2084 VOUT-.t47 GNDA 0.285754f
C2085 VOUT-.t91 GNDA 0.285754f
C2086 VOUT-.t41 GNDA 0.285754f
C2087 VOUT-.t130 GNDA 0.285754f
C2088 VOUT-.t82 GNDA 0.285754f
C2089 VOUT-.t124 GNDA 0.285754f
C2090 VOUT-.t72 GNDA 0.285754f
C2091 VOUT-.t23 GNDA 0.285754f
C2092 VOUT-.t62 GNDA 0.285754f
C2093 VOUT-.t150 GNDA 0.285754f
C2094 VOUT-.t86 GNDA 0.281558f
C2095 VOUT-.n19 GNDA 0.189376f
C2096 VOUT-.t50 GNDA 0.281558f
C2097 VOUT-.n20 GNDA 0.242168f
C2098 VOUT-.t137 GNDA 0.281558f
C2099 VOUT-.n21 GNDA 0.242168f
C2100 VOUT-.t105 GNDA 0.281558f
C2101 VOUT-.n22 GNDA 0.242168f
C2102 VOUT-.t73 GNDA 0.281558f
C2103 VOUT-.n23 GNDA 0.242168f
C2104 VOUT-.t25 GNDA 0.281558f
C2105 VOUT-.n24 GNDA 0.242168f
C2106 VOUT-.t127 GNDA 0.281558f
C2107 VOUT-.n25 GNDA 0.242168f
C2108 VOUT-.t88 GNDA 0.281558f
C2109 VOUT-.n26 GNDA 0.242168f
C2110 VOUT-.t53 GNDA 0.281558f
C2111 VOUT-.n27 GNDA 0.242168f
C2112 VOUT-.t140 GNDA 0.281558f
C2113 VOUT-.n28 GNDA 0.242168f
C2114 VOUT-.t109 GNDA 0.281558f
C2115 VOUT-.t28 GNDA 0.286354f
C2116 VOUT-.t78 GNDA 0.281558f
C2117 VOUT-.n29 GNDA 0.188776f
C2118 VOUT-.n30 GNDA 0.228766f
C2119 VOUT-.t24 GNDA 0.286354f
C2120 VOUT-.t112 GNDA 0.281558f
C2121 VOUT-.n31 GNDA 0.188776f
C2122 VOUT-.t77 GNDA 0.281558f
C2123 VOUT-.t129 GNDA 0.286354f
C2124 VOUT-.t37 GNDA 0.281558f
C2125 VOUT-.n32 GNDA 0.188776f
C2126 VOUT-.n33 GNDA 0.228766f
C2127 VOUT-.t59 GNDA 0.286354f
C2128 VOUT-.t147 GNDA 0.281558f
C2129 VOUT-.n34 GNDA 0.188776f
C2130 VOUT-.t116 GNDA 0.281558f
C2131 VOUT-.t32 GNDA 0.286354f
C2132 VOUT-.t81 GNDA 0.281558f
C2133 VOUT-.n35 GNDA 0.188776f
C2134 VOUT-.n36 GNDA 0.228766f
C2135 VOUT-.t99 GNDA 0.286354f
C2136 VOUT-.t46 GNDA 0.281558f
C2137 VOUT-.n37 GNDA 0.188776f
C2138 VOUT-.t153 GNDA 0.281558f
C2139 VOUT-.t69 GNDA 0.286354f
C2140 VOUT-.t122 GNDA 0.281558f
C2141 VOUT-.n38 GNDA 0.188776f
C2142 VOUT-.n39 GNDA 0.228766f
C2143 VOUT-.t67 GNDA 0.286354f
C2144 VOUT-.t154 GNDA 0.281558f
C2145 VOUT-.n40 GNDA 0.188776f
C2146 VOUT-.t123 GNDA 0.281558f
C2147 VOUT-.t35 GNDA 0.286354f
C2148 VOUT-.t84 GNDA 0.281558f
C2149 VOUT-.n41 GNDA 0.188776f
C2150 VOUT-.n42 GNDA 0.228766f
C2151 VOUT-.t104 GNDA 0.286354f
C2152 VOUT-.t52 GNDA 0.281558f
C2153 VOUT-.n43 GNDA 0.188776f
C2154 VOUT-.t22 GNDA 0.281558f
C2155 VOUT-.t76 GNDA 0.286354f
C2156 VOUT-.t126 GNDA 0.281558f
C2157 VOUT-.n44 GNDA 0.188776f
C2158 VOUT-.n45 GNDA 0.228766f
C2159 VOUT-.t95 GNDA 0.281558f
C2160 VOUT-.t83 GNDA 0.286354f
C2161 VOUT-.t56 GNDA 0.281558f
C2162 VOUT-.n46 GNDA 0.188776f
C2163 VOUT-.n47 GNDA 0.123182f
C2164 VOUT-.t132 GNDA 0.285754f
C2165 VOUT-.t114 GNDA 0.285754f
C2166 VOUT-.t90 GNDA 0.286354f
C2167 VOUT-.t131 GNDA 0.281558f
C2168 VOUT-.n48 GNDA 0.188776f
C2169 VOUT-.t103 GNDA 0.281558f
C2170 VOUT-.n49 GNDA 0.123182f
C2171 VOUT-.t71 GNDA 0.281558f
C2172 VOUT-.n50 GNDA 0.118782f
C2173 VOUT-.t146 GNDA 0.285754f
C2174 VOUT-.t128 GNDA 0.286354f
C2175 VOUT-.t31 GNDA 0.281558f
C2176 VOUT-.n51 GNDA 0.188776f
C2177 VOUT-.t138 GNDA 0.281558f
C2178 VOUT-.n52 GNDA 0.123182f
C2179 VOUT-.t106 GNDA 0.281558f
C2180 VOUT-.n53 GNDA 0.118782f
C2181 VOUT-.t45 GNDA 0.285754f
C2182 VOUT-.t26 GNDA 0.286354f
C2183 VOUT-.t60 GNDA 0.281558f
C2184 VOUT-.n54 GNDA 0.188776f
C2185 VOUT-.t40 GNDA 0.281558f
C2186 VOUT-.n55 GNDA 0.123182f
C2187 VOUT-.t143 GNDA 0.281558f
C2188 VOUT-.n56 GNDA 0.118782f
C2189 VOUT-.t85 GNDA 0.285754f
C2190 VOUT-.t74 GNDA 0.286354f
C2191 VOUT-.t113 GNDA 0.281558f
C2192 VOUT-.n57 GNDA 0.188776f
C2193 VOUT-.t21 GNDA 0.281558f
C2194 VOUT-.n58 GNDA 0.123182f
C2195 VOUT-.t125 GNDA 0.281558f
C2196 VOUT-.n59 GNDA 0.118782f
C2197 VOUT-.t63 GNDA 0.285754f
C2198 VOUT-.t101 GNDA 0.285754f
C2199 VOUT-.t134 GNDA 0.285754f
C2200 VOUT-.t119 GNDA 0.285754f
C2201 VOUT-.t155 GNDA 0.285754f
C2202 VOUT-.t118 GNDA 0.281558f
C2203 VOUT-.n60 GNDA 0.189376f
C2204 VOUT-.t80 GNDA 0.281558f
C2205 VOUT-.n61 GNDA 0.242168f
C2206 VOUT-.t96 GNDA 0.281558f
C2207 VOUT-.n62 GNDA 0.242168f
C2208 VOUT-.t61 GNDA 0.281558f
C2209 VOUT-.n63 GNDA 0.242168f
C2210 VOUT-.t27 GNDA 0.281558f
C2211 VOUT-.n64 GNDA 0.29936f
C2212 VOUT-.t44 GNDA 0.281558f
C2213 VOUT-.n65 GNDA 0.29936f
C2214 VOUT-.t144 GNDA 0.281558f
C2215 VOUT-.n66 GNDA 0.29936f
C2216 VOUT-.t111 GNDA 0.281558f
C2217 VOUT-.n67 GNDA 0.29936f
C2218 VOUT-.t75 GNDA 0.281558f
C2219 VOUT-.n68 GNDA 0.242168f
C2220 VOUT-.t92 GNDA 0.281558f
C2221 VOUT-.n69 GNDA 0.242168f
C2222 VOUT-.t55 GNDA 0.281558f
C2223 VOUT-.t39 GNDA 0.286354f
C2224 VOUT-.t19 GNDA 0.281558f
C2225 VOUT-.n70 GNDA 0.188776f
C2226 VOUT-.n71 GNDA 0.228766f
C2227 VOUT-.t34 GNDA 0.286354f
C2228 VOUT-.t51 GNDA 0.281558f
C2229 VOUT-.n72 GNDA 0.188776f
C2230 VOUT-.t156 GNDA 0.281558f
C2231 VOUT-.t136 GNDA 0.286354f
C2232 VOUT-.t120 GNDA 0.281558f
C2233 VOUT-.n73 GNDA 0.188776f
C2234 VOUT-.n74 GNDA 0.228766f
C2235 VOUT-.t68 GNDA 0.286354f
C2236 VOUT-.t87 GNDA 0.281558f
C2237 VOUT-.n75 GNDA 0.188776f
C2238 VOUT-.t49 GNDA 0.281558f
C2239 VOUT-.t36 GNDA 0.286354f
C2240 VOUT-.t151 GNDA 0.281558f
C2241 VOUT-.n76 GNDA 0.188776f
C2242 VOUT-.n77 GNDA 0.228766f
C2243 VOUT-.t94 GNDA 0.286354f
C2244 VOUT-.t42 GNDA 0.281558f
C2245 VOUT-.n78 GNDA 0.188776f
C2246 VOUT-.t145 GNDA 0.281558f
C2247 VOUT-.t64 GNDA 0.286354f
C2248 VOUT-.t117 GNDA 0.281558f
C2249 VOUT-.n79 GNDA 0.188776f
C2250 VOUT-.n80 GNDA 0.228766f
C2251 VOUT-.t54 GNDA 0.286354f
C2252 VOUT-.t141 GNDA 0.281558f
C2253 VOUT-.n81 GNDA 0.188776f
C2254 VOUT-.t110 GNDA 0.281558f
C2255 VOUT-.t29 GNDA 0.286354f
C2256 VOUT-.t79 GNDA 0.281558f
C2257 VOUT-.n82 GNDA 0.188776f
C2258 VOUT-.n83 GNDA 0.228766f
C2259 VOUT-.t89 GNDA 0.286354f
C2260 VOUT-.t38 GNDA 0.281558f
C2261 VOUT-.n84 GNDA 0.188776f
C2262 VOUT-.t139 GNDA 0.281558f
C2263 VOUT-.t57 GNDA 0.286354f
C2264 VOUT-.t108 GNDA 0.281558f
C2265 VOUT-.n85 GNDA 0.188776f
C2266 VOUT-.n86 GNDA 0.228766f
C2267 VOUT-.t48 GNDA 0.286354f
C2268 VOUT-.t135 GNDA 0.281558f
C2269 VOUT-.n87 GNDA 0.188776f
C2270 VOUT-.t102 GNDA 0.281558f
C2271 VOUT-.t20 GNDA 0.286354f
C2272 VOUT-.t70 GNDA 0.281558f
C2273 VOUT-.n88 GNDA 0.188776f
C2274 VOUT-.n89 GNDA 0.228766f
C2275 VOUT-.t148 GNDA 0.286354f
C2276 VOUT-.t98 GNDA 0.281558f
C2277 VOUT-.n90 GNDA 0.188776f
C2278 VOUT-.t66 GNDA 0.281558f
C2279 VOUT-.t121 GNDA 0.286354f
C2280 VOUT-.t33 GNDA 0.281558f
C2281 VOUT-.n91 GNDA 0.188776f
C2282 VOUT-.n92 GNDA 0.228766f
C2283 VOUT-.t43 GNDA 0.286354f
C2284 VOUT-.t133 GNDA 0.281558f
C2285 VOUT-.n93 GNDA 0.188776f
C2286 VOUT-.t97 GNDA 0.281558f
C2287 VOUT-.t152 GNDA 0.286354f
C2288 VOUT-.t65 GNDA 0.281558f
C2289 VOUT-.n94 GNDA 0.188776f
C2290 VOUT-.n95 GNDA 0.228766f
C2291 VOUT-.t115 GNDA 0.286354f
C2292 VOUT-.t30 GNDA 0.281558f
C2293 VOUT-.n96 GNDA 0.188776f
C2294 VOUT-.t58 GNDA 0.281558f
C2295 VOUT-.n97 GNDA 0.228766f
C2296 VOUT-.t93 GNDA 0.281558f
C2297 VOUT-.n98 GNDA 0.123182f
C2298 VOUT-.t142 GNDA 0.281558f
C2299 VOUT-.n99 GNDA 0.23068f
C2300 VOUT-.n100 GNDA 0.259376f
C2301 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2302 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2303 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2304 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2305 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2306 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2307 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2308 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2309 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2310 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2311 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2312 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2313 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2314 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2315 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2316 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2317 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2318 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2319 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2320 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2321 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.04969f
C2322 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.186051f
C2323 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2324 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2325 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.050131f
C2326 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2327 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2328 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2329 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.186051f
C2330 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.027755f
C2331 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2332 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2333 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2334 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2335 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2336 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2337 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2338 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2339 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2340 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2341 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2342 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2343 VDDA.t375 GNDA 0.019589f
C2344 VDDA.t404 GNDA 0.019589f
C2345 VDDA.n0 GNDA 0.08101f
C2346 VDDA.t40 GNDA 0.019589f
C2347 VDDA.t302 GNDA 0.019589f
C2348 VDDA.n1 GNDA 0.080699f
C2349 VDDA.n2 GNDA 0.111885f
C2350 VDDA.t363 GNDA 0.019589f
C2351 VDDA.t9 GNDA 0.019589f
C2352 VDDA.n3 GNDA 0.080699f
C2353 VDDA.n4 GNDA 0.058383f
C2354 VDDA.t355 GNDA 0.019589f
C2355 VDDA.t382 GNDA 0.019589f
C2356 VDDA.n5 GNDA 0.080699f
C2357 VDDA.n6 GNDA 0.058383f
C2358 VDDA.t354 GNDA 0.019589f
C2359 VDDA.t306 GNDA 0.019589f
C2360 VDDA.n7 GNDA 0.080699f
C2361 VDDA.n8 GNDA 0.058383f
C2362 VDDA.t402 GNDA 0.019589f
C2363 VDDA.t305 GNDA 0.019589f
C2364 VDDA.n9 GNDA 0.080699f
C2365 VDDA.n10 GNDA 0.168617f
C2366 VDDA.t295 GNDA 0.039178f
C2367 VDDA.t274 GNDA 0.039178f
C2368 VDDA.n11 GNDA 0.157178f
C2369 VDDA.n12 GNDA 0.079851f
C2370 VDDA.t180 GNDA 0.039028f
C2371 VDDA.n13 GNDA 0.052848f
C2372 VDDA.n14 GNDA 0.074595f
C2373 VDDA.t183 GNDA 0.043345f
C2374 VDDA.t181 GNDA 0.018981f
C2375 VDDA.n15 GNDA 0.068758f
C2376 VDDA.n16 GNDA 0.040477f
C2377 VDDA.t162 GNDA 0.043345f
C2378 VDDA.t160 GNDA 0.018981f
C2379 VDDA.n17 GNDA 0.068758f
C2380 VDDA.n18 GNDA 0.040477f
C2381 VDDA.n19 GNDA 0.043096f
C2382 VDDA.n20 GNDA 0.074595f
C2383 VDDA.n21 GNDA 0.215645f
C2384 VDDA.t161 GNDA 0.267071f
C2385 VDDA.t270 GNDA 0.154428f
C2386 VDDA.t281 GNDA 0.154428f
C2387 VDDA.t282 GNDA 0.154428f
C2388 VDDA.t227 GNDA 0.154428f
C2389 VDDA.t66 GNDA 0.115821f
C2390 VDDA.n22 GNDA 0.077214f
C2391 VDDA.t267 GNDA 0.115821f
C2392 VDDA.t224 GNDA 0.154428f
C2393 VDDA.t266 GNDA 0.154428f
C2394 VDDA.t223 GNDA 0.154428f
C2395 VDDA.t290 GNDA 0.154428f
C2396 VDDA.t182 GNDA 0.267071f
C2397 VDDA.n23 GNDA 0.215645f
C2398 VDDA.n24 GNDA 0.052848f
C2399 VDDA.n25 GNDA 0.100005f
C2400 VDDA.n26 GNDA 0.068439f
C2401 VDDA.n27 GNDA 0.101516f
C2402 VDDA.n28 GNDA 0.101516f
C2403 VDDA.n29 GNDA 0.100854f
C2404 VDDA.t150 GNDA 0.039028f
C2405 VDDA.t297 GNDA 0.039178f
C2406 VDDA.t277 GNDA 0.039178f
C2407 VDDA.n30 GNDA 0.157178f
C2408 VDDA.n31 GNDA 0.079851f
C2409 VDDA.t15 GNDA 0.039178f
C2410 VDDA.t279 GNDA 0.039178f
C2411 VDDA.n32 GNDA 0.157178f
C2412 VDDA.n33 GNDA 0.079851f
C2413 VDDA.t284 GNDA 0.039178f
C2414 VDDA.t292 GNDA 0.039178f
C2415 VDDA.n34 GNDA 0.157178f
C2416 VDDA.n35 GNDA 0.079851f
C2417 VDDA.t272 GNDA 0.039178f
C2418 VDDA.t226 GNDA 0.039178f
C2419 VDDA.n36 GNDA 0.157178f
C2420 VDDA.n37 GNDA 0.167794f
C2421 VDDA.n38 GNDA 0.126688f
C2422 VDDA.t148 GNDA 0.047355f
C2423 VDDA.n39 GNDA 0.090605f
C2424 VDDA.n40 GNDA 0.052934f
C2425 VDDA.n41 GNDA 0.079201f
C2426 VDDA.n42 GNDA 0.348615f
C2427 VDDA.t149 GNDA 0.538472f
C2428 VDDA.t271 GNDA 0.298081f
C2429 VDDA.t225 GNDA 0.298081f
C2430 VDDA.t283 GNDA 0.298081f
C2431 VDDA.t291 GNDA 0.298081f
C2432 VDDA.t14 GNDA 0.223561f
C2433 VDDA.n43 GNDA 0.149041f
C2434 VDDA.t278 GNDA 0.223561f
C2435 VDDA.t296 GNDA 0.298081f
C2436 VDDA.t276 GNDA 0.298081f
C2437 VDDA.t294 GNDA 0.298081f
C2438 VDDA.t273 GNDA 0.298081f
C2439 VDDA.t179 GNDA 0.538472f
C2440 VDDA.n44 GNDA 0.348615f
C2441 VDDA.n45 GNDA 0.079201f
C2442 VDDA.n46 GNDA 0.052934f
C2443 VDDA.t178 GNDA 0.047355f
C2444 VDDA.n47 GNDA 0.090605f
C2445 VDDA.n48 GNDA 0.126361f
C2446 VDDA.n49 GNDA 0.0948f
C2447 VDDA.t403 GNDA 0.019589f
C2448 VDDA.t65 GNDA 0.019589f
C2449 VDDA.n50 GNDA 0.08101f
C2450 VDDA.t293 GNDA 0.019589f
C2451 VDDA.t16 GNDA 0.019589f
C2452 VDDA.n51 GNDA 0.080699f
C2453 VDDA.n52 GNDA 0.111885f
C2454 VDDA.t289 GNDA 0.019589f
C2455 VDDA.t268 GNDA 0.019589f
C2456 VDDA.n53 GNDA 0.080699f
C2457 VDDA.n54 GNDA 0.058383f
C2458 VDDA.t265 GNDA 0.019589f
C2459 VDDA.t280 GNDA 0.019589f
C2460 VDDA.n55 GNDA 0.080699f
C2461 VDDA.n56 GNDA 0.058383f
C2462 VDDA.t275 GNDA 0.019589f
C2463 VDDA.t269 GNDA 0.019589f
C2464 VDDA.n57 GNDA 0.080699f
C2465 VDDA.n58 GNDA 0.058383f
C2466 VDDA.t89 GNDA 0.019589f
C2467 VDDA.t405 GNDA 0.019589f
C2468 VDDA.n59 GNDA 0.080699f
C2469 VDDA.n60 GNDA 0.201709f
C2470 VDDA.n61 GNDA 0.186425f
C2471 VDDA.t91 GNDA 0.022854f
C2472 VDDA.t288 GNDA 0.022854f
C2473 VDDA.n62 GNDA 0.079481f
C2474 VDDA.t229 GNDA 0.022854f
C2475 VDDA.t242 GNDA 0.022854f
C2476 VDDA.n63 GNDA 0.0792f
C2477 VDDA.n64 GNDA 0.149521f
C2478 VDDA.t373 GNDA 0.022854f
C2479 VDDA.t88 GNDA 0.022854f
C2480 VDDA.n65 GNDA 0.079481f
C2481 VDDA.t73 GNDA 0.022854f
C2482 VDDA.t304 GNDA 0.022854f
C2483 VDDA.n66 GNDA 0.0792f
C2484 VDDA.n67 GNDA 0.149521f
C2485 VDDA.n68 GNDA 0.020895f
C2486 VDDA.n69 GNDA 0.065063f
C2487 VDDA.n70 GNDA 0.088473f
C2488 VDDA.t186 GNDA 0.112744f
C2489 VDDA.t184 GNDA 0.039797f
C2490 VDDA.n71 GNDA 0.073551f
C2491 VDDA.n72 GNDA 0.047414f
C2492 VDDA.t108 GNDA 0.112744f
C2493 VDDA.t106 GNDA 0.039797f
C2494 VDDA.n73 GNDA 0.073551f
C2495 VDDA.n74 GNDA 0.047414f
C2496 VDDA.n75 GNDA 0.047014f
C2497 VDDA.n76 GNDA 0.088473f
C2498 VDDA.n77 GNDA 0.263664f
C2499 VDDA.t107 GNDA 0.393556f
C2500 VDDA.t90 GNDA 0.227234f
C2501 VDDA.t287 GNDA 0.227234f
C2502 VDDA.t228 GNDA 0.227234f
C2503 VDDA.t241 GNDA 0.227234f
C2504 VDDA.t11 GNDA 0.170425f
C2505 VDDA.n78 GNDA 0.113617f
C2506 VDDA.t298 GNDA 0.170425f
C2507 VDDA.t72 GNDA 0.227234f
C2508 VDDA.t303 GNDA 0.227234f
C2509 VDDA.t372 GNDA 0.227234f
C2510 VDDA.t87 GNDA 0.227234f
C2511 VDDA.t185 GNDA 0.393556f
C2512 VDDA.n79 GNDA 0.263664f
C2513 VDDA.n80 GNDA 0.065063f
C2514 VDDA.n81 GNDA 0.091085f
C2515 VDDA.t12 GNDA 0.022854f
C2516 VDDA.t299 GNDA 0.022854f
C2517 VDDA.n82 GNDA 0.074514f
C2518 VDDA.n83 GNDA 0.050857f
C2519 VDDA.n84 GNDA 0.028368f
C2520 VDDA.n85 GNDA 0.11398f
C2521 VDDA.t69 GNDA 0.022854f
C2522 VDDA.t71 GNDA 0.022854f
C2523 VDDA.n86 GNDA 0.079481f
C2524 VDDA.t33 GNDA 0.022854f
C2525 VDDA.t101 GNDA 0.022854f
C2526 VDDA.n87 GNDA 0.0792f
C2527 VDDA.n88 GNDA 0.149521f
C2528 VDDA.t443 GNDA 0.022854f
C2529 VDDA.t384 GNDA 0.022854f
C2530 VDDA.n89 GNDA 0.079481f
C2531 VDDA.t357 GNDA 0.022854f
C2532 VDDA.t80 GNDA 0.022854f
C2533 VDDA.n90 GNDA 0.0792f
C2534 VDDA.n91 GNDA 0.149521f
C2535 VDDA.n92 GNDA 0.020895f
C2536 VDDA.n93 GNDA 0.065063f
C2537 VDDA.n94 GNDA 0.088473f
C2538 VDDA.t126 GNDA 0.112744f
C2539 VDDA.t124 GNDA 0.039797f
C2540 VDDA.n95 GNDA 0.073551f
C2541 VDDA.n96 GNDA 0.047414f
C2542 VDDA.t207 GNDA 0.112744f
C2543 VDDA.t205 GNDA 0.039797f
C2544 VDDA.n97 GNDA 0.073551f
C2545 VDDA.n98 GNDA 0.047414f
C2546 VDDA.n99 GNDA 0.047014f
C2547 VDDA.n100 GNDA 0.088473f
C2548 VDDA.n101 GNDA 0.263664f
C2549 VDDA.t206 GNDA 0.393556f
C2550 VDDA.t68 GNDA 0.227234f
C2551 VDDA.t70 GNDA 0.227234f
C2552 VDDA.t32 GNDA 0.227234f
C2553 VDDA.t100 GNDA 0.227234f
C2554 VDDA.t387 GNDA 0.170425f
C2555 VDDA.n102 GNDA 0.113617f
C2556 VDDA.t23 GNDA 0.170425f
C2557 VDDA.t356 GNDA 0.227234f
C2558 VDDA.t79 GNDA 0.227234f
C2559 VDDA.t442 GNDA 0.227234f
C2560 VDDA.t383 GNDA 0.227234f
C2561 VDDA.t125 GNDA 0.393556f
C2562 VDDA.n103 GNDA 0.263664f
C2563 VDDA.n104 GNDA 0.065063f
C2564 VDDA.n105 GNDA 0.091085f
C2565 VDDA.t388 GNDA 0.022854f
C2566 VDDA.t24 GNDA 0.022854f
C2567 VDDA.n106 GNDA 0.074514f
C2568 VDDA.n107 GNDA 0.050857f
C2569 VDDA.n108 GNDA 0.028368f
C2570 VDDA.n109 GNDA 0.112021f
C2571 VDDA.t54 GNDA 0.039178f
C2572 VDDA.t39 GNDA 0.039178f
C2573 VDDA.n110 GNDA 0.157178f
C2574 VDDA.n111 GNDA 0.079851f
C2575 VDDA.t138 GNDA 0.039028f
C2576 VDDA.n112 GNDA 0.079201f
C2577 VDDA.n113 GNDA 0.052848f
C2578 VDDA.n114 GNDA 0.074595f
C2579 VDDA.t123 GNDA 0.043345f
C2580 VDDA.t121 GNDA 0.018981f
C2581 VDDA.n115 GNDA 0.068758f
C2582 VDDA.n116 GNDA 0.040477f
C2583 VDDA.t141 GNDA 0.043345f
C2584 VDDA.t139 GNDA 0.018981f
C2585 VDDA.n117 GNDA 0.068758f
C2586 VDDA.n118 GNDA 0.040477f
C2587 VDDA.n119 GNDA 0.043096f
C2588 VDDA.n120 GNDA 0.074595f
C2589 VDDA.n121 GNDA 0.215645f
C2590 VDDA.t140 GNDA 0.267071f
C2591 VDDA.t255 GNDA 0.154428f
C2592 VDDA.t364 GNDA 0.154428f
C2593 VDDA.t10 GNDA 0.154428f
C2594 VDDA.t95 GNDA 0.154428f
C2595 VDDA.t62 GNDA 0.115821f
C2596 VDDA.n122 GNDA 0.077214f
C2597 VDDA.t365 GNDA 0.115821f
C2598 VDDA.t374 GNDA 0.154428f
C2599 VDDA.t251 GNDA 0.154428f
C2600 VDDA.t254 GNDA 0.154428f
C2601 VDDA.t353 GNDA 0.154428f
C2602 VDDA.t122 GNDA 0.267071f
C2603 VDDA.n123 GNDA 0.215645f
C2604 VDDA.n124 GNDA 0.052848f
C2605 VDDA.n125 GNDA 0.100005f
C2606 VDDA.t153 GNDA 0.039028f
C2607 VDDA.t301 GNDA 0.039178f
C2608 VDDA.t97 GNDA 0.039178f
C2609 VDDA.n126 GNDA 0.157178f
C2610 VDDA.n127 GNDA 0.079851f
C2611 VDDA.t60 GNDA 0.039178f
C2612 VDDA.t367 GNDA 0.039178f
C2613 VDDA.n128 GNDA 0.157178f
C2614 VDDA.n129 GNDA 0.079851f
C2615 VDDA.t381 GNDA 0.039178f
C2616 VDDA.t253 GNDA 0.039178f
C2617 VDDA.n130 GNDA 0.157178f
C2618 VDDA.n131 GNDA 0.079851f
C2619 VDDA.t52 GNDA 0.039178f
C2620 VDDA.t58 GNDA 0.039178f
C2621 VDDA.n132 GNDA 0.157178f
C2622 VDDA.n133 GNDA 0.167794f
C2623 VDDA.n134 GNDA 0.126688f
C2624 VDDA.t151 GNDA 0.047355f
C2625 VDDA.n135 GNDA 0.090605f
C2626 VDDA.n136 GNDA 0.052934f
C2627 VDDA.n137 GNDA 0.348615f
C2628 VDDA.n138 GNDA 0.348615f
C2629 VDDA.t137 GNDA 0.538472f
C2630 VDDA.t53 GNDA 0.298081f
C2631 VDDA.t38 GNDA 0.298081f
C2632 VDDA.t300 GNDA 0.298081f
C2633 VDDA.t96 GNDA 0.298081f
C2634 VDDA.t59 GNDA 0.223561f
C2635 VDDA.n139 GNDA 0.079201f
C2636 VDDA.n140 GNDA 0.101516f
C2637 VDDA.n141 GNDA 0.101516f
C2638 VDDA.t152 GNDA 0.538472f
C2639 VDDA.t57 GNDA 0.298081f
C2640 VDDA.t51 GNDA 0.298081f
C2641 VDDA.t252 GNDA 0.298081f
C2642 VDDA.t380 GNDA 0.298081f
C2643 VDDA.t366 GNDA 0.223561f
C2644 VDDA.n142 GNDA 0.149041f
C2645 VDDA.n143 GNDA 0.100854f
C2646 VDDA.n144 GNDA 0.068439f
C2647 VDDA.n145 GNDA 0.052934f
C2648 VDDA.t136 GNDA 0.047355f
C2649 VDDA.n146 GNDA 0.090605f
C2650 VDDA.n147 GNDA 0.126361f
C2651 VDDA.n148 GNDA 0.096759f
C2652 VDDA.n149 GNDA 0.054197f
C2653 VDDA.n150 GNDA 0.183277f
C2654 VDDA.n151 GNDA 0.063257f
C2655 VDDA.n152 GNDA 0.168876f
C2656 VDDA.t117 GNDA 0.012304f
C2657 VDDA.n153 GNDA 0.02618f
C2658 VDDA.t216 GNDA 0.012304f
C2659 VDDA.n154 GNDA 0.02618f
C2660 VDDA.n155 GNDA 0.038012f
C2661 VDDA.n156 GNDA 0.06389f
C2662 VDDA.n157 GNDA 0.17027f
C2663 VDDA.t144 GNDA 0.012304f
C2664 VDDA.n158 GNDA 0.02618f
C2665 VDDA.t132 GNDA 0.012304f
C2666 VDDA.n159 GNDA 0.02618f
C2667 VDDA.n160 GNDA 0.035424f
C2668 VDDA.n161 GNDA 0.043972f
C2669 VDDA.n162 GNDA 0.17027f
C2670 VDDA.t131 GNDA 0.16564f
C2671 VDDA.t390 GNDA 0.102353f
C2672 VDDA.t286 GNDA 0.102353f
C2673 VDDA.t13 GNDA 0.102353f
C2674 VDDA.t233 GNDA 0.102353f
C2675 VDDA.t61 GNDA 0.076765f
C2676 VDDA.t143 GNDA 0.16564f
C2677 VDDA.t448 GNDA 0.102353f
C2678 VDDA.t56 GNDA 0.102353f
C2679 VDDA.t234 GNDA 0.102353f
C2680 VDDA.t63 GNDA 0.102353f
C2681 VDDA.t67 GNDA 0.076765f
C2682 VDDA.n163 GNDA 0.064524f
C2683 VDDA.n164 GNDA 0.051177f
C2684 VDDA.n165 GNDA 0.064524f
C2685 VDDA.n166 GNDA 0.043096f
C2686 VDDA.n167 GNDA 0.034869f
C2687 VDDA.n168 GNDA 0.081074f
C2688 VDDA.n169 GNDA 0.081074f
C2689 VDDA.n170 GNDA 0.168876f
C2690 VDDA.t215 GNDA 0.1623f
C2691 VDDA.t235 GNDA 0.100558f
C2692 VDDA.t344 GNDA 0.100558f
C2693 VDDA.t31 GNDA 0.100558f
C2694 VDDA.t55 GNDA 0.100558f
C2695 VDDA.t78 GNDA 0.075418f
C2696 VDDA.t116 GNDA 0.1623f
C2697 VDDA.t389 GNDA 0.100558f
C2698 VDDA.t236 GNDA 0.100558f
C2699 VDDA.t391 GNDA 0.100558f
C2700 VDDA.t232 GNDA 0.100558f
C2701 VDDA.t452 GNDA 0.075418f
C2702 VDDA.n171 GNDA 0.064524f
C2703 VDDA.n172 GNDA 0.050279f
C2704 VDDA.n173 GNDA 0.064524f
C2705 VDDA.n174 GNDA 0.042891f
C2706 VDDA.n175 GNDA 0.034869f
C2707 VDDA.n176 GNDA 0.067502f
C2708 VDDA.n177 GNDA 0.090296f
C2709 VDDA.n179 GNDA 0.049996f
C2710 VDDA.n180 GNDA 0.07901f
C2711 VDDA.n181 GNDA 0.100246f
C2712 VDDA.n182 GNDA 0.100246f
C2713 VDDA.n183 GNDA 0.100246f
C2714 VDDA.n185 GNDA 0.049996f
C2715 VDDA.n187 GNDA 0.049996f
C2716 VDDA.n189 GNDA 0.049996f
C2717 VDDA.n191 GNDA 0.049996f
C2718 VDDA.n193 GNDA 0.049996f
C2719 VDDA.n195 GNDA 0.049996f
C2720 VDDA.n197 GNDA 0.049996f
C2721 VDDA.n199 GNDA 0.049996f
C2722 VDDA.n201 GNDA 0.081815f
C2723 VDDA.t198 GNDA 0.011897f
C2724 VDDA.n202 GNDA 0.017664f
C2725 VDDA.n203 GNDA 0.015629f
C2726 VDDA.n204 GNDA 0.05338f
C2727 VDDA.n205 GNDA 0.062025f
C2728 VDDA.n206 GNDA 0.204981f
C2729 VDDA.t197 GNDA 0.1623f
C2730 VDDA.t322 GNDA 0.100558f
C2731 VDDA.t324 GNDA 0.100558f
C2732 VDDA.t19 GNDA 0.100558f
C2733 VDDA.t7 GNDA 0.100558f
C2734 VDDA.t245 GNDA 0.100558f
C2735 VDDA.t43 GNDA 0.100558f
C2736 VDDA.t239 GNDA 0.100558f
C2737 VDDA.t1 GNDA 0.100558f
C2738 VDDA.t378 GNDA 0.100558f
C2739 VDDA.t320 GNDA 0.075418f
C2740 VDDA.n207 GNDA 0.050279f
C2741 VDDA.t5 GNDA 0.075418f
C2742 VDDA.t3 GNDA 0.100558f
C2743 VDDA.t47 GNDA 0.100558f
C2744 VDDA.t243 GNDA 0.100558f
C2745 VDDA.t326 GNDA 0.100558f
C2746 VDDA.t237 GNDA 0.100558f
C2747 VDDA.t45 GNDA 0.100558f
C2748 VDDA.t376 GNDA 0.100558f
C2749 VDDA.t21 GNDA 0.100558f
C2750 VDDA.t49 GNDA 0.100558f
C2751 VDDA.t191 GNDA 0.1623f
C2752 VDDA.n208 GNDA 0.204981f
C2753 VDDA.n209 GNDA 0.062025f
C2754 VDDA.n210 GNDA 0.05338f
C2755 VDDA.n211 GNDA 0.015629f
C2756 VDDA.t192 GNDA 0.011897f
C2757 VDDA.n212 GNDA 0.017233f
C2758 VDDA.n213 GNDA 0.085732f
C2759 VDDA.n214 GNDA 0.079723f
C2760 VDDA.n215 GNDA 0.011843f
C2761 VDDA.n216 GNDA 0.056719f
C2762 VDDA.n217 GNDA 0.023507f
C2763 VDDA.t201 GNDA 0.015799f
C2764 VDDA.t199 GNDA 0.012804f
C2765 VDDA.n218 GNDA 0.029209f
C2766 VDDA.t220 GNDA 0.015799f
C2767 VDDA.t217 GNDA 0.012543f
C2768 VDDA.n219 GNDA 0.029209f
C2769 VDDA.n220 GNDA 0.064659f
C2770 VDDA.n221 GNDA 0.064659f
C2771 VDDA.n222 GNDA 0.062638f
C2772 VDDA.t120 GNDA 0.019678f
C2773 VDDA.n223 GNDA 0.015388f
C2774 VDDA.n224 GNDA 0.011843f
C2775 VDDA.n225 GNDA 0.078447f
C2776 VDDA.n226 GNDA 0.025208f
C2777 VDDA.t118 GNDA 0.022936f
C2778 VDDA.n227 GNDA 0.018366f
C2779 VDDA.n228 GNDA 0.036049f
C2780 VDDA.n229 GNDA 0.045849f
C2781 VDDA.n230 GNDA 0.18268f
C2782 VDDA.t119 GNDA 0.193474f
C2783 VDDA.t249 GNDA 0.123412f
C2784 VDDA.t473 GNDA 0.123412f
C2785 VDDA.t385 GNDA 0.123412f
C2786 VDDA.t98 GNDA 0.118269f
C2787 VDDA.n231 GNDA 0.061706f
C2788 VDDA.t176 GNDA 0.138838f
C2789 VDDA.t200 GNDA 0.195402f
C2790 VDDA.t17 GNDA 0.123412f
C2791 VDDA.t218 GNDA 0.193474f
C2792 VDDA.n232 GNDA 0.177404f
C2793 VDDA.n233 GNDA 0.04321f
C2794 VDDA.n234 GNDA 0.026581f
C2795 VDDA.n235 GNDA 0.019206f
C2796 VDDA.t175 GNDA 0.014339f
C2797 VDDA.n237 GNDA 0.018366f
C2798 VDDA.t177 GNDA 0.019678f
C2799 VDDA.n238 GNDA 0.020138f
C2800 VDDA.n239 GNDA 0.044254f
C2801 VDDA.n241 GNDA 0.101146f
C2802 VDDA.n242 GNDA 0.498827f
C2803 VDDA.t468 GNDA 0.365011f
C2804 VDDA.t330 GNDA 0.366334f
C2805 VDDA.t256 GNDA 0.365011f
C2806 VDDA.t0 GNDA 0.366334f
C2807 VDDA.t328 GNDA 0.365011f
C2808 VDDA.t329 GNDA 0.366334f
C2809 VDDA.t331 GNDA 0.365011f
C2810 VDDA.t81 GNDA 0.366334f
C2811 VDDA.t92 GNDA 0.365011f
C2812 VDDA.t309 GNDA 0.366334f
C2813 VDDA.t30 GNDA 0.365011f
C2814 VDDA.t28 GNDA 0.366334f
C2815 VDDA.t312 GNDA 0.365011f
C2816 VDDA.t315 GNDA 0.366334f
C2817 VDDA.t285 GNDA 0.365011f
C2818 VDDA.t29 GNDA 0.366334f
C2819 VDDA.n243 GNDA 0.244667f
C2820 VDDA.t25 GNDA 0.194841f
C2821 VDDA.n244 GNDA 0.26547f
C2822 VDDA.t451 GNDA 0.194841f
C2823 VDDA.n245 GNDA 0.26547f
C2824 VDDA.t358 GNDA 0.194841f
C2825 VDDA.n246 GNDA 0.26547f
C2826 VDDA.t463 GNDA 0.290742f
C2827 VDDA.n247 GNDA 0.45064f
C2828 VDDA.t341 GNDA 0.016324f
C2829 VDDA.t337 GNDA 0.016324f
C2830 VDDA.n248 GNDA 0.05265f
C2831 VDDA.n249 GNDA 0.079251f
C2832 VDDA.n250 GNDA 0.052699f
C2833 VDDA.t211 GNDA 0.080323f
C2834 VDDA.t213 GNDA 0.076112f
C2835 VDDA.t84 GNDA 0.016324f
C2836 VDDA.t103 GNDA 0.016324f
C2837 VDDA.n251 GNDA 0.05265f
C2838 VDDA.n252 GNDA 0.079251f
C2839 VDDA.t343 GNDA 0.016324f
C2840 VDDA.t339 GNDA 0.016324f
C2841 VDDA.n253 GNDA 0.05265f
C2842 VDDA.n254 GNDA 0.079251f
C2843 VDDA.n255 GNDA 0.052699f
C2844 VDDA.t169 GNDA 0.080323f
C2845 VDDA.t171 GNDA 0.076112f
C2846 VDDA.t86 GNDA 0.016324f
C2847 VDDA.t352 GNDA 0.016324f
C2848 VDDA.n256 GNDA 0.05265f
C2849 VDDA.n257 GNDA 0.104081f
C2850 VDDA.n258 GNDA 0.071107f
C2851 VDDA.n259 GNDA 0.038224f
C2852 VDDA.n260 GNDA 0.302361f
C2853 VDDA.n261 GNDA 0.302361f
C2854 VDDA.t188 GNDA 0.338524f
C2855 VDDA.t342 GNDA 0.285022f
C2856 VDDA.t338 GNDA 0.213766f
C2857 VDDA.n262 GNDA 0.052699f
C2858 VDDA.n263 GNDA 0.070201f
C2859 VDDA.n264 GNDA 0.070201f
C2860 VDDA.t170 GNDA 0.338524f
C2861 VDDA.t351 GNDA 0.285022f
C2862 VDDA.t85 GNDA 0.213766f
C2863 VDDA.n265 GNDA 0.142511f
C2864 VDDA.n266 GNDA 0.070201f
C2865 VDDA.n267 GNDA 0.03526f
C2866 VDDA.n268 GNDA 0.038224f
C2867 VDDA.t189 GNDA 0.076112f
C2868 VDDA.t187 GNDA 0.080323f
C2869 VDDA.n269 GNDA 0.069308f
C2870 VDDA.n270 GNDA 0.079521f
C2871 VDDA.n271 GNDA 0.017285f
C2872 VDDA.n272 GNDA 0.068907f
C2873 VDDA.n273 GNDA 0.070521f
C2874 VDDA.n274 GNDA 0.095131f
C2875 VDDA.n275 GNDA 0.098468f
C2876 VDDA.n276 GNDA 0.095131f
C2877 VDDA.t163 GNDA 0.044973f
C2878 VDDA.t165 GNDA 0.025573f
C2879 VDDA.n277 GNDA 0.017285f
C2880 VDDA.n278 GNDA 0.093738f
C2881 VDDA.n279 GNDA 0.04991f
C2882 VDDA.n280 GNDA 0.052518f
C2883 VDDA.n281 GNDA 0.062507f
C2884 VDDA.n282 GNDA 0.243833f
C2885 VDDA.t164 GNDA 0.277731f
C2886 VDDA.t334 GNDA 0.211563f
C2887 VDDA.t318 GNDA 0.211563f
C2888 VDDA.t345 GNDA 0.211563f
C2889 VDDA.t347 GNDA 0.211563f
C2890 VDDA.t316 GNDA 0.158672f
C2891 VDDA.n283 GNDA 0.105781f
C2892 VDDA.t104 GNDA 0.158672f
C2893 VDDA.t76 GNDA 0.211563f
C2894 VDDA.t349 GNDA 0.211563f
C2895 VDDA.t392 GNDA 0.211563f
C2896 VDDA.t74 GNDA 0.211563f
C2897 VDDA.t113 GNDA 0.277731f
C2898 VDDA.n284 GNDA 0.243833f
C2899 VDDA.n285 GNDA 0.062507f
C2900 VDDA.n286 GNDA 0.052518f
C2901 VDDA.t114 GNDA 0.025573f
C2902 VDDA.t112 GNDA 0.044973f
C2903 VDDA.n287 GNDA 0.04991f
C2904 VDDA.n288 GNDA 0.017285f
C2905 VDDA.n289 GNDA 0.093738f
C2906 VDDA.n290 GNDA 0.017285f
C2907 VDDA.n291 GNDA 0.068907f
C2908 VDDA.n292 GNDA 0.028731f
C2909 VDDA.n293 GNDA 0.01677f
C2910 VDDA.n294 GNDA 0.060204f
C2911 VDDA.n295 GNDA 0.118265f
C2912 VDDA.n296 GNDA 0.079521f
C2913 VDDA.n297 GNDA 0.069308f
C2914 VDDA.n298 GNDA 0.038224f
C2915 VDDA.n299 GNDA 0.300244f
C2916 VDDA.n300 GNDA 0.300244f
C2917 VDDA.t203 GNDA 0.334765f
C2918 VDDA.t340 GNDA 0.282084f
C2919 VDDA.t336 GNDA 0.211563f
C2920 VDDA.n301 GNDA 0.052699f
C2921 VDDA.n302 GNDA 0.070201f
C2922 VDDA.n303 GNDA 0.070201f
C2923 VDDA.t212 GNDA 0.334765f
C2924 VDDA.t102 GNDA 0.282084f
C2925 VDDA.t83 GNDA 0.211563f
C2926 VDDA.n304 GNDA 0.141042f
C2927 VDDA.n305 GNDA 0.070201f
C2928 VDDA.n306 GNDA 0.03526f
C2929 VDDA.n307 GNDA 0.038224f
C2930 VDDA.t204 GNDA 0.076112f
C2931 VDDA.t202 GNDA 0.080323f
C2932 VDDA.n308 GNDA 0.069308f
C2933 VDDA.n309 GNDA 0.061731f
C2934 VDDA.n310 GNDA 0.117694f
C2935 VDDA.t264 GNDA 0.019589f
C2936 VDDA.t27 GNDA 0.019589f
C2937 VDDA.n311 GNDA 0.064716f
C2938 VDDA.n312 GNDA 0.083508f
C2939 VDDA.n313 GNDA 0.091744f
C2940 VDDA.t166 GNDA 0.093409f
C2941 VDDA.t168 GNDA 0.060033f
C2942 VDDA.t472 GNDA 0.019589f
C2943 VDDA.t456 GNDA 0.019589f
C2944 VDDA.n314 GNDA 0.064716f
C2945 VDDA.n315 GNDA 0.083508f
C2946 VDDA.t462 GNDA 0.019589f
C2947 VDDA.t231 GNDA 0.019589f
C2948 VDDA.n316 GNDA 0.064716f
C2949 VDDA.n317 GNDA 0.083508f
C2950 VDDA.t260 GNDA 0.019589f
C2951 VDDA.t314 GNDA 0.019589f
C2952 VDDA.n318 GNDA 0.064716f
C2953 VDDA.n319 GNDA 0.083508f
C2954 VDDA.t311 GNDA 0.019589f
C2955 VDDA.t467 GNDA 0.019589f
C2956 VDDA.n320 GNDA 0.064716f
C2957 VDDA.n321 GNDA 0.083508f
C2958 VDDA.t262 GNDA 0.019589f
C2959 VDDA.t450 GNDA 0.019589f
C2960 VDDA.n322 GNDA 0.064716f
C2961 VDDA.n323 GNDA 0.083508f
C2962 VDDA.t465 GNDA 0.019589f
C2963 VDDA.t258 GNDA 0.019589f
C2964 VDDA.n324 GNDA 0.064716f
C2965 VDDA.n325 GNDA 0.083508f
C2966 VDDA.t470 GNDA 0.019589f
C2967 VDDA.t460 GNDA 0.019589f
C2968 VDDA.n326 GNDA 0.064716f
C2969 VDDA.n327 GNDA 0.083508f
C2970 VDDA.t111 GNDA 0.024529f
C2971 VDDA.t109 GNDA 0.012379f
C2972 VDDA.n328 GNDA 0.038673f
C2973 VDDA.n329 GNDA 0.0223f
C2974 VDDA.n330 GNDA 0.039632f
C2975 VDDA.t135 GNDA 0.024529f
C2976 VDDA.t133 GNDA 0.012379f
C2977 VDDA.n331 GNDA 0.038673f
C2978 VDDA.n332 GNDA 0.039632f
C2979 VDDA.n333 GNDA 0.039632f
C2980 VDDA.n334 GNDA 0.032519f
C2981 VDDA.n335 GNDA 0.164144f
C2982 VDDA.t110 GNDA 0.199107f
C2983 VDDA.t82 GNDA 0.088886f
C2984 VDDA.n336 GNDA 0.059257f
C2985 VDDA.t64 GNDA 0.088886f
C2986 VDDA.t134 GNDA 0.196213f
C2987 VDDA.n337 GNDA 0.156264f
C2988 VDDA.n338 GNDA 0.032519f
C2989 VDDA.n339 GNDA 0.0223f
C2990 VDDA.n340 GNDA 0.031329f
C2991 VDDA.n341 GNDA 0.092202f
C2992 VDDA.n342 GNDA 0.11148f
C2993 VDDA.n343 GNDA 0.075143f
C2994 VDDA.n344 GNDA 0.338033f
C2995 VDDA.n345 GNDA 0.338033f
C2996 VDDA.t173 GNDA 0.436176f
C2997 VDDA.t263 GNDA 0.314406f
C2998 VDDA.t26 GNDA 0.314406f
C2999 VDDA.t471 GNDA 0.314406f
C3000 VDDA.t455 GNDA 0.314406f
C3001 VDDA.t461 GNDA 0.314406f
C3002 VDDA.t230 GNDA 0.314406f
C3003 VDDA.t259 GNDA 0.314406f
C3004 VDDA.t313 GNDA 0.235804f
C3005 VDDA.n346 GNDA 0.091744f
C3006 VDDA.n347 GNDA 0.1442f
C3007 VDDA.n348 GNDA 0.1442f
C3008 VDDA.t167 GNDA 0.436176f
C3009 VDDA.t459 GNDA 0.314406f
C3010 VDDA.t469 GNDA 0.314406f
C3011 VDDA.t257 GNDA 0.314406f
C3012 VDDA.t464 GNDA 0.314406f
C3013 VDDA.t449 GNDA 0.314406f
C3014 VDDA.t261 GNDA 0.314406f
C3015 VDDA.t466 GNDA 0.314406f
C3016 VDDA.t310 GNDA 0.235804f
C3017 VDDA.n349 GNDA 0.157203f
C3018 VDDA.n350 GNDA 0.143537f
C3019 VDDA.n351 GNDA 0.105781f
C3020 VDDA.n352 GNDA 0.075143f
C3021 VDDA.t174 GNDA 0.060033f
C3022 VDDA.t172 GNDA 0.093409f
C3023 VDDA.n353 GNDA 0.11148f
C3024 VDDA.n354 GNDA 0.055743f
C3025 VDDA.n355 GNDA 0.01577f
C3026 VDDA.t210 GNDA 0.024711f
C3027 VDDA.t208 GNDA 0.03882f
C3028 VDDA.n356 GNDA 0.036536f
C3029 VDDA.n357 GNDA 0.026675f
C3030 VDDA.n358 GNDA 0.048561f
C3031 VDDA.t129 GNDA 0.024711f
C3032 VDDA.t127 GNDA 0.03882f
C3033 VDDA.n359 GNDA 0.036536f
C3034 VDDA.n360 GNDA 0.048561f
C3035 VDDA.n361 GNDA 0.048561f
C3036 VDDA.n362 GNDA 0.037196f
C3037 VDDA.n363 GNDA 0.193751f
C3038 VDDA.t209 GNDA 0.254272f
C3039 VDDA.t394 GNDA 0.145449f
C3040 VDDA.n364 GNDA 0.096966f
C3041 VDDA.t332 GNDA 0.145449f
C3042 VDDA.t128 GNDA 0.251747f
C3043 VDDA.n365 GNDA 0.185502f
C3044 VDDA.n366 GNDA 0.037196f
C3045 VDDA.n367 GNDA 0.026675f
C3046 VDDA.n368 GNDA 0.032649f
C3047 VDDA.n369 GNDA 0.043637f
C3048 VDDA.n370 GNDA 0.090849f
C3049 VDDA.n371 GNDA 0.175846f
C3050 VDDA.n372 GNDA 0.020895f
C3051 VDDA.n373 GNDA 0.015815f
C3052 VDDA.n374 GNDA 0.032585f
C3053 VDDA.n375 GNDA 0.020895f
C3054 VDDA.n376 GNDA 0.020895f
C3055 VDDA.n377 GNDA 0.015815f
C3056 VDDA.n378 GNDA 0.015815f
C3057 VDDA.n379 GNDA 0.046217f
C3058 VDDA.n380 GNDA 0.020895f
C3059 VDDA.n381 GNDA 0.223805f
C3060 VDDA.n382 GNDA 0.223805f
C3061 VDDA.t155 GNDA 0.204128f
C3062 VDDA.t432 GNDA 0.129288f
C3063 VDDA.t412 GNDA 0.129288f
C3064 VDDA.t408 GNDA 0.129288f
C3065 VDDA.t428 GNDA 0.129288f
C3066 VDDA.t426 GNDA 0.129288f
C3067 VDDA.t440 GNDA 0.129288f
C3068 VDDA.t436 GNDA 0.129288f
C3069 VDDA.t424 GNDA 0.129288f
C3070 VDDA.t418 GNDA 0.096966f
C3071 VDDA.t156 GNDA 0.024529f
C3072 VDDA.t154 GNDA 0.016163f
C3073 VDDA.n383 GNDA 0.03848f
C3074 VDDA.n384 GNDA 0.054752f
C3075 VDDA.t195 GNDA 0.024529f
C3076 VDDA.t193 GNDA 0.016163f
C3077 VDDA.n385 GNDA 0.03848f
C3078 VDDA.n386 GNDA 0.020895f
C3079 VDDA.n387 GNDA 0.015815f
C3080 VDDA.n388 GNDA 0.015815f
C3081 VDDA.n389 GNDA 0.020895f
C3082 VDDA.n390 GNDA 0.046217f
C3083 VDDA.n391 GNDA 0.020895f
C3084 VDDA.n392 GNDA 0.015815f
C3085 VDDA.n393 GNDA 0.046217f
C3086 VDDA.n394 GNDA 0.020895f
C3087 VDDA.n395 GNDA 0.016536f
C3088 VDDA.n396 GNDA 0.016424f
C3089 VDDA.n397 GNDA 0.127672f
C3090 VDDA.n398 GNDA 0.016424f
C3091 VDDA.n399 GNDA 0.066504f
C3092 VDDA.n400 GNDA 0.016424f
C3093 VDDA.n401 GNDA 0.066504f
C3094 VDDA.n402 GNDA 0.064229f
C3095 VDDA.n403 GNDA 0.102932f
C3096 VDDA.t147 GNDA 0.024529f
C3097 VDDA.t145 GNDA 0.016163f
C3098 VDDA.n404 GNDA 0.03848f
C3099 VDDA.n405 GNDA 0.054752f
C3100 VDDA.t159 GNDA 0.024529f
C3101 VDDA.t157 GNDA 0.016163f
C3102 VDDA.n406 GNDA 0.03848f
C3103 VDDA.n407 GNDA 0.054752f
C3104 VDDA.n408 GNDA 0.078356f
C3105 VDDA.n409 GNDA 0.102932f
C3106 VDDA.n410 GNDA 0.223805f
C3107 VDDA.t158 GNDA 0.204128f
C3108 VDDA.t400 GNDA 0.129288f
C3109 VDDA.t247 GNDA 0.129288f
C3110 VDDA.t359 GNDA 0.129288f
C3111 VDDA.t41 GNDA 0.129288f
C3112 VDDA.t453 GNDA 0.129288f
C3113 VDDA.t221 GNDA 0.129288f
C3114 VDDA.t370 GNDA 0.129288f
C3115 VDDA.t93 GNDA 0.129288f
C3116 VDDA.t34 GNDA 0.096966f
C3117 VDDA.n411 GNDA 0.064644f
C3118 VDDA.t307 GNDA 0.096966f
C3119 VDDA.t368 GNDA 0.129288f
C3120 VDDA.t398 GNDA 0.129288f
C3121 VDDA.t396 GNDA 0.129288f
C3122 VDDA.t361 GNDA 0.129288f
C3123 VDDA.t36 GNDA 0.129288f
C3124 VDDA.t457 GNDA 0.129288f
C3125 VDDA.t444 GNDA 0.129288f
C3126 VDDA.t446 GNDA 0.129288f
C3127 VDDA.t146 GNDA 0.204128f
C3128 VDDA.n412 GNDA 0.223805f
C3129 VDDA.n413 GNDA 0.064229f
C3130 VDDA.n414 GNDA 0.109417f
C3131 VDDA.n415 GNDA 0.015815f
C3132 VDDA.n416 GNDA 0.046217f
C3133 VDDA.n417 GNDA 0.020895f
C3134 VDDA.n418 GNDA 0.016424f
C3135 VDDA.n419 GNDA 0.066504f
C3136 VDDA.n420 GNDA 0.016424f
C3137 VDDA.n421 GNDA 0.066504f
C3138 VDDA.n422 GNDA 0.016424f
C3139 VDDA.n423 GNDA 0.066504f
C3140 VDDA.n424 GNDA 0.016424f
C3141 VDDA.n425 GNDA 0.095234f
C3142 VDDA.n426 GNDA 0.049626f
C3143 VDDA.n427 GNDA 0.046217f
C3144 VDDA.n428 GNDA 0.034115f
C3145 VDDA.n429 GNDA 0.032585f
C3146 VDDA.n430 GNDA 0.054752f
C3147 VDDA.n431 GNDA 0.078356f
C3148 VDDA.n432 GNDA 0.102932f
C3149 VDDA.t194 GNDA 0.204128f
C3150 VDDA.t430 GNDA 0.129288f
C3151 VDDA.t414 GNDA 0.129288f
C3152 VDDA.t420 GNDA 0.129288f
C3153 VDDA.t416 GNDA 0.129288f
C3154 VDDA.t422 GNDA 0.129288f
C3155 VDDA.t434 GNDA 0.129288f
C3156 VDDA.t438 GNDA 0.129288f
C3157 VDDA.t406 GNDA 0.129288f
C3158 VDDA.t410 GNDA 0.096966f
C3159 VDDA.n433 GNDA 0.064644f
C3160 VDDA.n434 GNDA 0.102932f
C3161 VDDA.n435 GNDA 0.020895f
C3162 VDDA.n436 GNDA 0.046217f
C3163 VDDA.n437 GNDA 0.020895f
C3164 VDDA.n438 GNDA 0.015815f
C3165 VDDA.n439 GNDA 0.046217f
C3166 VDDA.n440 GNDA 0.020895f
C3167 VDDA.n441 GNDA 0.020895f
C3168 VDDA.n442 GNDA 0.015815f
C3169 VDDA.n443 GNDA 0.046217f
C3170 VDDA.n444 GNDA 0.020895f
C3171 VDDA.n445 GNDA 0.015815f
C3172 VDDA.n446 GNDA 0.046217f
C3173 VDDA.n447 GNDA 0.020895f
C3174 VDDA.n448 GNDA 0.034115f
C3175 VDDA.n449 GNDA 0.046217f
C3176 VDDA.n450 GNDA 0.063258f
C3177 VDDA.n451 GNDA 0.192054f
C3178 VDDA.t475 GNDA 0.721887f
C3179 VDDA.t478 GNDA 0.737779f
C3180 VDDA.t476 GNDA 0.769393f
C3181 VDDA.n452 GNDA 0.515727f
C3182 VDDA.t477 GNDA 0.769393f
C3183 VDDA.n453 GNDA 0.250385f
C3184 VDDA.n454 GNDA 0.321009f
C3185 VDDA.n455 GNDA 2.60145f
C3186 VDDA.n456 GNDA 3.1197f
C3187 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n0 GNDA 0.849209f
C3188 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n1 GNDA 1.77369f
C3189 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n2 GNDA 2.45745f
C3190 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n3 GNDA 0.155832f
C3191 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t29 GNDA 0.430574f
C3192 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t11 GNDA 0.437907f
C3193 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t20 GNDA 0.430574f
C3194 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t26 GNDA 0.430574f
C3195 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t28 GNDA 0.437907f
C3196 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t33 GNDA 0.430574f
C3197 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t18 GNDA 0.437907f
C3198 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t25 GNDA 0.430574f
C3199 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t31 GNDA 0.430574f
C3200 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t34 GNDA 0.437907f
C3201 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t13 GNDA 0.430574f
C3202 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t36 GNDA 0.437907f
C3203 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t17 GNDA 0.430574f
C3204 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t24 GNDA 0.430574f
C3205 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t27 GNDA 0.437907f
C3206 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t30 GNDA 0.430574f
C3207 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t21 GNDA 0.437907f
C3208 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t23 GNDA 0.430574f
C3209 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t16 GNDA 0.430574f
C3210 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t35 GNDA 0.430574f
C3211 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t22 GNDA 0.028128f
C3212 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t10 GNDA 0.010764f
C3213 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t7 GNDA 0.010764f
C3214 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n4 GNDA 0.027135f
C3215 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t12 GNDA 0.016398f
C3216 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t15 GNDA 0.016398f
C3217 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n5 GNDA 0.036479f
C3218 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t8 GNDA 0.010764f
C3219 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t6 GNDA 0.010764f
C3220 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n6 GNDA 0.02601f
C3221 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t4 GNDA 0.022672f
C3222 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n7 GNDA 0.015549f
C3223 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n8 GNDA 0.235193f
C3224 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n9 GNDA 0.014069f
C3225 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t14 GNDA 0.016398f
C3226 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t19 GNDA 0.016398f
C3227 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n10 GNDA 0.036479f
C3228 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t9 GNDA 0.010764f
C3229 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t5 GNDA 0.010764f
C3230 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.n11 GNDA 0.027135f
C3231 ref_volt_cur_gen_dummy_magic_0.1st_Vout_2.t32 GNDA 0.025738f
C3232 ref_volt_cur_gen_dummy_magic_0.V_mir2.n0 GNDA 0.362016f
C3233 ref_volt_cur_gen_dummy_magic_0.V_mir2.t10 GNDA 0.03537f
C3234 ref_volt_cur_gen_dummy_magic_0.V_mir2.t16 GNDA 0.03537f
C3235 ref_volt_cur_gen_dummy_magic_0.V_mir2.t12 GNDA 0.03537f
C3236 ref_volt_cur_gen_dummy_magic_0.V_mir2.n1 GNDA 0.08097f
C3237 ref_volt_cur_gen_dummy_magic_0.V_mir2.t15 GNDA 0.053881f
C3238 ref_volt_cur_gen_dummy_magic_0.V_mir2.t11 GNDA 0.042444f
C3239 ref_volt_cur_gen_dummy_magic_0.V_mir2.t19 GNDA 0.042444f
C3240 ref_volt_cur_gen_dummy_magic_0.V_mir2.t20 GNDA 0.06851f
C3241 ref_volt_cur_gen_dummy_magic_0.V_mir2.n2 GNDA 0.076506f
C3242 ref_volt_cur_gen_dummy_magic_0.V_mir2.n3 GNDA 0.052264f
C3243 ref_volt_cur_gen_dummy_magic_0.V_mir2.n4 GNDA 0.081315f
C3244 ref_volt_cur_gen_dummy_magic_0.V_mir2.n5 GNDA 0.201563f
C3245 ref_volt_cur_gen_dummy_magic_0.V_mir2.t8 GNDA 0.03537f
C3246 ref_volt_cur_gen_dummy_magic_0.V_mir2.t14 GNDA 0.03537f
C3247 ref_volt_cur_gen_dummy_magic_0.V_mir2.n6 GNDA 0.08097f
C3248 ref_volt_cur_gen_dummy_magic_0.V_mir2.t7 GNDA 0.053881f
C3249 ref_volt_cur_gen_dummy_magic_0.V_mir2.t13 GNDA 0.042444f
C3250 ref_volt_cur_gen_dummy_magic_0.V_mir2.t21 GNDA 0.042444f
C3251 ref_volt_cur_gen_dummy_magic_0.V_mir2.t22 GNDA 0.06851f
C3252 ref_volt_cur_gen_dummy_magic_0.V_mir2.n7 GNDA 0.076506f
C3253 ref_volt_cur_gen_dummy_magic_0.V_mir2.n8 GNDA 0.052264f
C3254 ref_volt_cur_gen_dummy_magic_0.V_mir2.n9 GNDA 0.081315f
C3255 ref_volt_cur_gen_dummy_magic_0.V_mir2.n10 GNDA 0.156007f
C3256 ref_volt_cur_gen_dummy_magic_0.V_mir2.t0 GNDA 0.017685f
C3257 ref_volt_cur_gen_dummy_magic_0.V_mir2.t4 GNDA 0.017685f
C3258 ref_volt_cur_gen_dummy_magic_0.V_mir2.n11 GNDA 0.046242f
C3259 ref_volt_cur_gen_dummy_magic_0.V_mir2.t1 GNDA 0.075466f
C3260 ref_volt_cur_gen_dummy_magic_0.V_mir2.t2 GNDA 0.017685f
C3261 ref_volt_cur_gen_dummy_magic_0.V_mir2.t3 GNDA 0.017685f
C3262 ref_volt_cur_gen_dummy_magic_0.V_mir2.n12 GNDA 0.050199f
C3263 ref_volt_cur_gen_dummy_magic_0.V_mir2.n13 GNDA 0.827814f
C3264 ref_volt_cur_gen_dummy_magic_0.V_mir2.n14 GNDA 0.699157f
C3265 ref_volt_cur_gen_dummy_magic_0.V_mir2.t5 GNDA 0.053881f
C3266 ref_volt_cur_gen_dummy_magic_0.V_mir2.t9 GNDA 0.042444f
C3267 ref_volt_cur_gen_dummy_magic_0.V_mir2.t17 GNDA 0.042444f
C3268 ref_volt_cur_gen_dummy_magic_0.V_mir2.t18 GNDA 0.06851f
C3269 ref_volt_cur_gen_dummy_magic_0.V_mir2.n15 GNDA 0.076506f
C3270 ref_volt_cur_gen_dummy_magic_0.V_mir2.n16 GNDA 0.052264f
C3271 ref_volt_cur_gen_dummy_magic_0.V_mir2.n17 GNDA 0.081315f
C3272 ref_volt_cur_gen_dummy_magic_0.V_mir2.n18 GNDA 0.203577f
C3273 ref_volt_cur_gen_dummy_magic_0.V_mir2.n19 GNDA 0.08097f
C3274 ref_volt_cur_gen_dummy_magic_0.V_mir2.t6 GNDA 0.03537f
.ends

