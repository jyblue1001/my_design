* PEX produced on Mon Feb 17 02:31:17 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from charge_pump_cell_5.ext - technology: sky130A

.subckt charge_pump_magic VDDA GNDA x vout UP_b DOWN I_IN UP_input DOWN_input opamp_out
X0 VDDA.t21 VDDA.t18 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X1 GNDA.t30 GNDA.t28 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X2 UP_input.t0 UP_b.t0 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=8.75
X3 x.t3 I_IN.t4 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X4 GNDA.t27 GNDA.t25 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X5 GNDA.t3 I_IN.t5 x.t2 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X6 VDDA.t17 VDDA.t15 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X7 GNDA.t24 GNDA.t21 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X8 GNDA.t20 GNDA.t18 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X9 vout.t5 DOWN_input.t0 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X10 GNDA.t32 DOWN_input.t1 vout.t4 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X11 x.t5 opamp_out.t0 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X12 GNDA.t17 GNDA.t14 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X13 VDDA.t14 VDDA.t12 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X14 VDDA.t11 VDDA.t8 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X15 VDDA.t7 opamp_out.t1 x.t1 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X16 vout.t3 UP_input.t1 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X17 VDDA.t23 UP_input.t2 vout.t2 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X18 GNDA.t9 I_IN.t2 I_IN.t3 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X19 x.t0 opamp_out.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X20 DOWN_input.t2 DOWN.t0 sky130_fd_pr__cap_mim_m3_1 l=2.6 w=3.35
X21 VDDA.t27 opamp_out.t3 x.t4 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X22 VDDA.t5 UP_input.t3 vout.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X23 I_IN.t1 I_IN.t0 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X24 vout.t0 UP_input.t4 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X25 GNDA.t13 GNDA.t10 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
R0 VDDA.n97 VDDA.n2 585
R1 VDDA.n90 VDDA.n2 585
R2 VDDA.n87 VDDA.n86 585
R3 VDDA.n86 VDDA.n85 585
R4 VDDA.n56 VDDA.n55 585
R5 VDDA.n56 VDDA.n45 585
R6 VDDA.t13 VDDA.t22 360.346
R7 VDDA.t22 VDDA.t24 360.346
R8 VDDA.t24 VDDA.t4 360.346
R9 VDDA.t4 VDDA.t0 360.346
R10 VDDA.t0 VDDA.t19 360.346
R11 VDDA.t6 VDDA.t16 360.346
R12 VDDA.t2 VDDA.t6 360.346
R13 VDDA.t26 VDDA.t2 360.346
R14 VDDA.t28 VDDA.t26 360.346
R15 VDDA.t9 VDDA.t28 360.346
R16 VDDA.n51 VDDA.t13 343.966
R17 VDDA.n89 VDDA.t19 343.966
R18 VDDA.t16 VDDA.n89 343.966
R19 VDDA.n95 VDDA.t9 343.966
R20 VDDA.n84 VDDA.t15 336.329
R21 VDDA.n84 VDDA.t18 336.329
R22 VDDA.n46 VDDA.t12 320.7
R23 VDDA.n98 VDDA.t8 320.7
R24 VDDA.n86 VDDA.n10 291.363
R25 VDDA.n82 VDDA.n8 291.363
R26 VDDA.n83 VDDA.n82 291.363
R27 VDDA.n91 VDDA.n2 290.733
R28 VDDA.n56 VDDA.n44 290.733
R29 VDDA.n97 VDDA.n96 230.308
R30 VDDA.n94 VDDA.n90 230.308
R31 VDDA.n88 VDDA.n87 230.308
R32 VDDA.n85 VDDA.n5 230.308
R33 VDDA.n19 VDDA.n18 196.502
R34 VDDA.n16 VDDA.n15 196.502
R35 VDDA.n81 VDDA.n80 196.502
R36 VDDA.n72 VDDA.n37 196.502
R37 VDDA.n65 VDDA.n40 196.502
R38 VDDA.n58 VDDA.n57 196.502
R39 VDDA.n9 VDDA.n6 185
R40 VDDA.n12 VDDA.n11 185
R41 VDDA.n4 VDDA.n3 185
R42 VDDA.n93 VDDA.n92 185
R43 VDDA.n55 VDDA.n47 185
R44 VDDA.n51 VDDA.n47 185
R45 VDDA.n54 VDDA.n53 185
R46 VDDA.n49 VDDA.n48 185
R47 VDDA.n50 VDDA.n45 185
R48 VDDA.n51 VDDA.n50 185
R49 VDDA.n85 VDDA.n84 166.63
R50 VDDA.n93 VDDA.n4 120.001
R51 VDDA.n11 VDDA.n6 120.001
R52 VDDA.n53 VDDA.n47 120.001
R53 VDDA.n50 VDDA.n49 120.001
R54 VDDA.n89 VDDA.n88 69.8479
R55 VDDA.n89 VDDA.n5 69.8479
R56 VDDA.n96 VDDA.n95 69.8479
R57 VDDA.n95 VDDA.n94 69.8479
R58 VDDA.n52 VDDA.n51 69.8479
R59 VDDA.n88 VDDA.n6 45.3071
R60 VDDA.n11 VDDA.n5 45.3071
R61 VDDA.n96 VDDA.n4 45.3071
R62 VDDA.n94 VDDA.n93 45.3071
R63 VDDA.n53 VDDA.n52 45.3071
R64 VDDA.n52 VDDA.n49 45.3071
R65 VDDA.n87 VDDA.n7 32.2291
R66 VDDA.n24 VDDA.n23 32.0005
R67 VDDA.n23 VDDA.n22 32.0005
R68 VDDA.n30 VDDA.n13 32.0005
R69 VDDA.n30 VDDA.n29 32.0005
R70 VDDA.n29 VDDA.n28 32.0005
R71 VDDA.n79 VDDA.n34 32.0005
R72 VDDA.n74 VDDA.n73 32.0005
R73 VDDA.n67 VDDA.n66 32.0005
R74 VDDA.n67 VDDA.n38 32.0005
R75 VDDA.n71 VDDA.n38 32.0005
R76 VDDA.n60 VDDA.n59 32.0005
R77 VDDA.n60 VDDA.n41 32.0005
R78 VDDA.n64 VDDA.n41 32.0005
R79 VDDA.n99 VDDA.n1 28.8005
R80 VDDA.n24 VDDA.n16 28.8005
R81 VDDA.n80 VDDA.n79 28.8005
R82 VDDA.n18 VDDA.t29 24.6255
R83 VDDA.n18 VDDA.t10 24.6255
R84 VDDA.n15 VDDA.t3 24.6255
R85 VDDA.n15 VDDA.t27 24.6255
R86 VDDA.t17 VDDA.n81 24.6255
R87 VDDA.n81 VDDA.t7 24.6255
R88 VDDA.n37 VDDA.t1 24.6255
R89 VDDA.n37 VDDA.t20 24.6255
R90 VDDA.n40 VDDA.t25 24.6255
R91 VDDA.n40 VDDA.t5 24.6255
R92 VDDA.n57 VDDA.t14 24.6255
R93 VDDA.n57 VDDA.t23 24.6255
R94 VDDA.t14 VDDA.n56 24.6255
R95 VDDA.n2 VDDA.t11 24.6255
R96 VDDA.n82 VDDA.t17 24.6255
R97 VDDA.n86 VDDA.t21 24.6255
R98 VDDA.n46 VDDA.n43 24.361
R99 VDDA.n22 VDDA.n19 22.4005
R100 VDDA.n73 VDDA.n72 22.4005
R101 VDDA.n74 VDDA.n7 22.4005
R102 VDDA.n99 VDDA.n98 17.6005
R103 VDDA.n19 VDDA.n1 16.0005
R104 VDDA.n34 VDDA.n7 16.0005
R105 VDDA.n72 VDDA.n71 16.0005
R106 VDDA.n59 VDDA.n58 16.0005
R107 VDDA.n98 VDDA.n97 15.6449
R108 VDDA.n55 VDDA.n46 15.6449
R109 VDDA.n80 VDDA.n13 9.6005
R110 VDDA.n28 VDDA.n16 9.6005
R111 VDDA.n59 VDDA.n42 9.3005
R112 VDDA.n61 VDDA.n60 9.3005
R113 VDDA.n62 VDDA.n41 9.3005
R114 VDDA.n64 VDDA.n63 9.3005
R115 VDDA.n66 VDDA.n39 9.3005
R116 VDDA.n68 VDDA.n67 9.3005
R117 VDDA.n69 VDDA.n38 9.3005
R118 VDDA.n71 VDDA.n70 9.3005
R119 VDDA.n72 VDDA.n36 9.3005
R120 VDDA.n73 VDDA.n35 9.3005
R121 VDDA.n75 VDDA.n74 9.3005
R122 VDDA.n76 VDDA.n7 9.3005
R123 VDDA.n77 VDDA.n34 9.3005
R124 VDDA.n79 VDDA.n78 9.3005
R125 VDDA.n80 VDDA.n33 9.3005
R126 VDDA.n32 VDDA.n13 9.3005
R127 VDDA.n31 VDDA.n30 9.3005
R128 VDDA.n29 VDDA.n14 9.3005
R129 VDDA.n28 VDDA.n27 9.3005
R130 VDDA.n26 VDDA.n16 9.3005
R131 VDDA.n25 VDDA.n24 9.3005
R132 VDDA.n23 VDDA.n17 9.3005
R133 VDDA.n22 VDDA.n21 9.3005
R134 VDDA.n20 VDDA.n19 9.3005
R135 VDDA.n1 VDDA.n0 9.3005
R136 VDDA.n97 VDDA.n3 7.11161
R137 VDDA.n92 VDDA.n90 7.11161
R138 VDDA.n55 VDDA.n54 7.11161
R139 VDDA.n48 VDDA.n45 7.11161
R140 VDDA.n58 VDDA.n43 6.54033
R141 VDDA.n100 VDDA.n99 5.98166
R142 VDDA.n91 VDDA.n3 3.53508
R143 VDDA.n92 VDDA.n91 3.53508
R144 VDDA.n54 VDDA.n44 3.53508
R145 VDDA.n48 VDDA.n44 3.53508
R146 VDDA.n66 VDDA.n65 3.2005
R147 VDDA.n65 VDDA.n64 3.2005
R148 VDDA.n9 VDDA.n8 2.27782
R149 VDDA.n10 VDDA.n9 2.27782
R150 VDDA.n85 VDDA.n83 2.27782
R151 VDDA.n12 VDDA.n10 2.27782
R152 VDDA.n87 VDDA.n8 2.27782
R153 VDDA.n83 VDDA.n12 2.27782
R154 VDDA.n43 VDDA.n42 0.703395
R155 VDDA VDDA.n100 0.527077
R156 VDDA.n100 VDDA.n0 0.224356
R157 VDDA.n61 VDDA.n42 0.15675
R158 VDDA.n62 VDDA.n61 0.15675
R159 VDDA.n63 VDDA.n62 0.15675
R160 VDDA.n63 VDDA.n39 0.15675
R161 VDDA.n68 VDDA.n39 0.15675
R162 VDDA.n69 VDDA.n68 0.15675
R163 VDDA.n70 VDDA.n69 0.15675
R164 VDDA.n70 VDDA.n36 0.15675
R165 VDDA.n36 VDDA.n35 0.15675
R166 VDDA.n75 VDDA.n35 0.15675
R167 VDDA.n76 VDDA.n75 0.15675
R168 VDDA.n77 VDDA.n76 0.15675
R169 VDDA.n78 VDDA.n77 0.15675
R170 VDDA.n78 VDDA.n33 0.15675
R171 VDDA.n33 VDDA.n32 0.15675
R172 VDDA.n32 VDDA.n31 0.15675
R173 VDDA.n31 VDDA.n14 0.15675
R174 VDDA.n27 VDDA.n14 0.15675
R175 VDDA.n27 VDDA.n26 0.15675
R176 VDDA.n26 VDDA.n25 0.15675
R177 VDDA.n25 VDDA.n17 0.15675
R178 VDDA.n21 VDDA.n17 0.15675
R179 VDDA.n21 VDDA.n20 0.15675
R180 VDDA.n20 VDDA.n0 0.15675
R181 GNDA.n113 GNDA.n107 26375.6
R182 GNDA.t31 GNDA.t19 733.333
R183 GNDA.t4 GNDA.t31 733.333
R184 GNDA.t15 GNDA.t4 733.333
R185 GNDA.t2 GNDA.t26 733.333
R186 GNDA.t0 GNDA.t2 733.333
R187 GNDA.t22 GNDA.t0 733.333
R188 GNDA.t29 GNDA.t8 733.333
R189 GNDA.t8 GNDA.t6 733.333
R190 GNDA.t6 GNDA.t11 733.333
R191 GNDA.n107 GNDA.t19 700
R192 GNDA.n80 GNDA.t15 700
R193 GNDA.n80 GNDA.t26 700
R194 GNDA.n59 GNDA.t22 700
R195 GNDA.n59 GNDA.t29 700
R196 GNDA.n113 GNDA.t11 700
R197 GNDA.n58 GNDA.n57 669.307
R198 GNDA.n61 GNDA.n60 669.307
R199 GNDA.n79 GNDA.n78 669.307
R200 GNDA.n82 GNDA.n81 669.307
R201 GNDA.n106 GNDA.n105 669.307
R202 GNDA.n100 GNDA.n6 669.307
R203 GNDA.n104 GNDA.n7 585
R204 GNDA.n102 GNDA.n101 585
R205 GNDA.n22 GNDA.n18 585
R206 GNDA.n20 GNDA.n17 585
R207 GNDA.n39 GNDA.n35 585
R208 GNDA.n37 GNDA.n34 585
R209 GNDA.n112 GNDA.n111 585
R210 GNDA.n113 GNDA.n112 585
R211 GNDA.n110 GNDA.n108 585
R212 GNDA.n4 GNDA.n2 585
R213 GNDA.n115 GNDA.n114 585
R214 GNDA.n114 GNDA.n113 585
R215 GNDA.n36 GNDA.t28 336.329
R216 GNDA.n36 GNDA.t21 336.329
R217 GNDA.n19 GNDA.t25 336.329
R218 GNDA.n19 GNDA.t14 336.329
R219 GNDA.n116 GNDA.t10 320.7
R220 GNDA.n99 GNDA.t18 320.7
R221 GNDA.n107 GNDA.n106 250.349
R222 GNDA.n107 GNDA.n6 250.349
R223 GNDA.n80 GNDA.n79 250.349
R224 GNDA.n81 GNDA.n80 250.349
R225 GNDA.n59 GNDA.n58 250.349
R226 GNDA.n60 GNDA.n59 250.349
R227 GNDA.n113 GNDA.n5 250.349
R228 GNDA.n35 GNDA.n34 197
R229 GNDA.n18 GNDA.n17 197
R230 GNDA.n101 GNDA.n7 197
R231 GNDA.n112 GNDA.n108 197
R232 GNDA.n114 GNDA.n4 197
R233 GNDA.n57 GNDA.n33 185
R234 GNDA.n61 GNDA.n33 185
R235 GNDA.n78 GNDA.n16 185
R236 GNDA.n82 GNDA.n16 185
R237 GNDA.n105 GNDA.n8 185
R238 GNDA.n100 GNDA.n8 185
R239 GNDA.n111 GNDA.n3 185
R240 GNDA.n115 GNDA.n3 185
R241 GNDA.n57 GNDA.n36 166.63
R242 GNDA.n78 GNDA.n19 166.63
R243 GNDA.n89 GNDA.n88 92.2612
R244 GNDA.n97 GNDA.n96 92.2612
R245 GNDA.n75 GNDA.n74 92.2612
R246 GNDA.n68 GNDA.n28 92.2612
R247 GNDA.n54 GNDA.n53 92.2612
R248 GNDA.n47 GNDA.n46 92.2612
R249 GNDA.n38 GNDA.n33 91.3721
R250 GNDA.n56 GNDA.n55 91.3721
R251 GNDA.n55 GNDA.n32 91.3721
R252 GNDA.n21 GNDA.n16 91.3721
R253 GNDA.n77 GNDA.n76 91.3721
R254 GNDA.n76 GNDA.n15 91.3721
R255 GNDA.n103 GNDA.n8 90.7567
R256 GNDA.n109 GNDA.n3 90.7567
R257 GNDA.n106 GNDA.n7 84.306
R258 GNDA.n101 GNDA.n6 84.306
R259 GNDA.n79 GNDA.n18 84.306
R260 GNDA.n81 GNDA.n17 84.306
R261 GNDA.n58 GNDA.n35 84.306
R262 GNDA.n60 GNDA.n34 84.306
R263 GNDA.n108 GNDA.n5 84.306
R264 GNDA.n5 GNDA.n4 84.306
R265 GNDA.n89 GNDA.n87 32.0005
R266 GNDA.n87 GNDA.n12 32.0005
R267 GNDA.n95 GNDA.n94 32.0005
R268 GNDA.n94 GNDA.n10 32.0005
R269 GNDA.n90 GNDA.n10 32.0005
R270 GNDA.n23 GNDA.n14 32.0005
R271 GNDA.n73 GNDA.n26 32.0005
R272 GNDA.n69 GNDA.n26 32.0005
R273 GNDA.n69 GNDA.n68 32.0005
R274 GNDA.n67 GNDA.n29 32.0005
R275 GNDA.n63 GNDA.n29 32.0005
R276 GNDA.n62 GNDA.n31 32.0005
R277 GNDA.n40 GNDA.n31 32.0005
R278 GNDA.n52 GNDA.n44 32.0005
R279 GNDA.n48 GNDA.n44 32.0005
R280 GNDA.n117 GNDA.n1 32.0005
R281 GNDA.n62 GNDA.n61 29.0291
R282 GNDA.n83 GNDA.n82 29.0291
R283 GNDA.n83 GNDA.n14 25.6005
R284 GNDA.n53 GNDA.n52 25.6005
R285 GNDA.n48 GNDA.n47 25.6005
R286 GNDA.n99 GNDA.n98 20.9665
R287 GNDA.n74 GNDA.n23 19.2005
R288 GNDA.n74 GNDA.n73 19.2005
R289 GNDA.n100 GNDA.n99 15.6449
R290 GNDA.n116 GNDA.n115 15.6449
R291 GNDA.n88 GNDA.t5 15.0005
R292 GNDA.n88 GNDA.t16 15.0005
R293 GNDA.n96 GNDA.t20 15.0005
R294 GNDA.n96 GNDA.t32 15.0005
R295 GNDA.t27 GNDA.n75 15.0005
R296 GNDA.n75 GNDA.t3 15.0005
R297 GNDA.n28 GNDA.t1 15.0005
R298 GNDA.n28 GNDA.t23 15.0005
R299 GNDA.t30 GNDA.n54 15.0005
R300 GNDA.n54 GNDA.t9 15.0005
R301 GNDA.n46 GNDA.t7 15.0005
R302 GNDA.n46 GNDA.t12 15.0005
R303 GNDA.n55 GNDA.t30 15.0005
R304 GNDA.n33 GNDA.t24 15.0005
R305 GNDA.n76 GNDA.t27 15.0005
R306 GNDA.n16 GNDA.t17 15.0005
R307 GNDA.t20 GNDA.n8 15.0005
R308 GNDA.n3 GNDA.t13 15.0005
R309 GNDA.n117 GNDA.n116 14.4005
R310 GNDA.n83 GNDA.n12 12.8005
R311 GNDA.n97 GNDA.n95 12.8005
R312 GNDA.n53 GNDA.n40 12.8005
R313 GNDA.n47 GNDA.n1 12.8005
R314 GNDA.n1 GNDA.n0 9.3005
R315 GNDA.n47 GNDA.n45 9.3005
R316 GNDA.n49 GNDA.n48 9.3005
R317 GNDA.n50 GNDA.n44 9.3005
R318 GNDA.n52 GNDA.n51 9.3005
R319 GNDA.n53 GNDA.n43 9.3005
R320 GNDA.n42 GNDA.n40 9.3005
R321 GNDA.n41 GNDA.n31 9.3005
R322 GNDA.n62 GNDA.n30 9.3005
R323 GNDA.n95 GNDA.n9 9.3005
R324 GNDA.n94 GNDA.n93 9.3005
R325 GNDA.n92 GNDA.n10 9.3005
R326 GNDA.n91 GNDA.n90 9.3005
R327 GNDA.n89 GNDA.n11 9.3005
R328 GNDA.n87 GNDA.n86 9.3005
R329 GNDA.n85 GNDA.n12 9.3005
R330 GNDA.n84 GNDA.n83 9.3005
R331 GNDA.n14 GNDA.n13 9.3005
R332 GNDA.n24 GNDA.n23 9.3005
R333 GNDA.n74 GNDA.n25 9.3005
R334 GNDA.n73 GNDA.n72 9.3005
R335 GNDA.n71 GNDA.n26 9.3005
R336 GNDA.n70 GNDA.n69 9.3005
R337 GNDA.n68 GNDA.n27 9.3005
R338 GNDA.n67 GNDA.n66 9.3005
R339 GNDA.n65 GNDA.n29 9.3005
R340 GNDA.n64 GNDA.n63 9.3005
R341 GNDA.n105 GNDA.n104 7.11161
R342 GNDA.n102 GNDA.n100 7.11161
R343 GNDA.n111 GNDA.n110 7.11161
R344 GNDA.n115 GNDA.n2 7.11161
R345 GNDA.n98 GNDA.n97 6.69883
R346 GNDA.n90 GNDA.n89 6.4005
R347 GNDA.n68 GNDA.n67 6.4005
R348 GNDA.n63 GNDA.n62 6.4005
R349 GNDA.n118 GNDA.n117 5.80512
R350 GNDA.n104 GNDA.n103 3.48951
R351 GNDA.n103 GNDA.n102 3.48951
R352 GNDA.n110 GNDA.n109 3.48951
R353 GNDA.n109 GNDA.n2 3.48951
R354 GNDA.n56 GNDA.n39 2.25882
R355 GNDA.n39 GNDA.n38 2.25882
R356 GNDA.n61 GNDA.n32 2.25882
R357 GNDA.n38 GNDA.n37 2.25882
R358 GNDA.n57 GNDA.n56 2.25882
R359 GNDA.n37 GNDA.n32 2.25882
R360 GNDA.n77 GNDA.n22 2.25882
R361 GNDA.n22 GNDA.n21 2.25882
R362 GNDA.n82 GNDA.n15 2.25882
R363 GNDA.n21 GNDA.n20 2.25882
R364 GNDA.n78 GNDA.n77 2.25882
R365 GNDA.n20 GNDA.n15 2.25882
R366 GNDA.n98 GNDA.n9 0.703977
R367 GNDA GNDA.n118 0.223516
R368 GNDA.n118 GNDA.n0 0.215014
R369 GNDA.n93 GNDA.n9 0.15675
R370 GNDA.n93 GNDA.n92 0.15675
R371 GNDA.n92 GNDA.n91 0.15675
R372 GNDA.n91 GNDA.n11 0.15675
R373 GNDA.n86 GNDA.n11 0.15675
R374 GNDA.n86 GNDA.n85 0.15675
R375 GNDA.n85 GNDA.n84 0.15675
R376 GNDA.n84 GNDA.n13 0.15675
R377 GNDA.n24 GNDA.n13 0.15675
R378 GNDA.n25 GNDA.n24 0.15675
R379 GNDA.n72 GNDA.n25 0.15675
R380 GNDA.n72 GNDA.n71 0.15675
R381 GNDA.n71 GNDA.n70 0.15675
R382 GNDA.n70 GNDA.n27 0.15675
R383 GNDA.n66 GNDA.n27 0.15675
R384 GNDA.n66 GNDA.n65 0.15675
R385 GNDA.n65 GNDA.n64 0.15675
R386 GNDA.n64 GNDA.n30 0.15675
R387 GNDA.n41 GNDA.n30 0.15675
R388 GNDA.n42 GNDA.n41 0.15675
R389 GNDA.n43 GNDA.n42 0.15675
R390 GNDA.n51 GNDA.n43 0.15675
R391 GNDA.n51 GNDA.n50 0.15675
R392 GNDA.n50 GNDA.n49 0.15675
R393 GNDA.n49 GNDA.n45 0.15675
R394 GNDA.n45 GNDA.n0 0.15675
R395 UP_input.n1 UP_input.t4 337.401
R396 UP_input UP_input.t0 326.658
R397 UP_input.n2 UP_input.t4 297.233
R398 UP_input.t2 UP_input.n3 297.233
R399 UP_input.n1 UP_input.n0 257.067
R400 UP_input UP_input.n0 226.942
R401 UP_input.n3 UP_input.n2 216.9
R402 UP_input UP_input.t2 92.3838
R403 UP_input.n2 UP_input.t3 80.3338
R404 UP_input.t3 UP_input.n1 80.3338
R405 UP_input.n3 UP_input.t1 80.3338
R406 UP_input.t1 UP_input.n0 80.3338
R407 UP_b UP_b.t0 12.0836
R408 I_IN.n2 I_IN.n1 1269.42
R409 I_IN.n2 I_IN.t0 275.325
R410 I_IN.n4 I_IN.n3 248.4
R411 I_IN I_IN.n4 214.4
R412 I_IN.n1 I_IN.t5 151.792
R413 I_IN.n3 I_IN.t2 140.583
R414 I_IN.n3 I_IN.t0 140.583
R415 I_IN.n4 I_IN.n0 98.6614
R416 I_IN.t2 I_IN.n2 80.3338
R417 I_IN.n1 I_IN.t4 44.2902
R418 I_IN.n0 I_IN.t3 15.0005
R419 I_IN.n0 I_IN.t1 15.0005
R420 x.n2 x.n1 242.903
R421 x.n2 x.n0 172.502
R422 x.n5 x.n4 105.061
R423 x.n5 x.n2 91.2005
R424 x.n0 x.t1 24.6255
R425 x.n0 x.t0 24.6255
R426 x.n1 x.t4 24.6255
R427 x.n1 x.t5 24.6255
R428 x.n4 x.t2 15.0005
R429 x.n4 x.t3 15.0005
R430 x.n5 x.n3 8.0005
R431 x x.n5 6.4005
R432 DOWN_input DOWN_input.t2 326.658
R433 DOWN_input DOWN_input.t0 307.276
R434 DOWN_input.n1 DOWN_input.t0 265.101
R435 DOWN_input.n1 DOWN_input.n0 172.718
R436 DOWN_input DOWN_input.t1 92.3838
R437 DOWN_input.t1 DOWN_input.n1 80.3338
R438 vout.n2 vout.n1 242.903
R439 vout.n2 vout.n0 172.502
R440 vout vout.n3 98.6614
R441 vout vout.n2 28.6428
R442 vout.n0 vout.t2 24.6255
R443 vout.n0 vout.t3 24.6255
R444 vout.n1 vout.t1 24.6255
R445 vout.n1 vout.t0 24.6255
R446 vout.n3 vout.t4 15.0005
R447 vout.n3 vout.t5 15.0005
R448 opamp_out.n1 opamp_out.t1 297.233
R449 opamp_out.n2 opamp_out.t1 297.233
R450 opamp_out.t0 opamp_out.n3 297.233
R451 opamp_out.n3 opamp_out.n2 216.9
R452 opamp_out.n1 opamp_out.n0 216.9
R453 opamp_out opamp_out.n0 184.768
R454 opamp_out opamp_out.t0 112.468
R455 opamp_out.n2 opamp_out.t2 80.3338
R456 opamp_out.t2 opamp_out.n1 80.3338
R457 opamp_out.n3 opamp_out.t3 80.3338
R458 opamp_out.t3 opamp_out.n0 80.3338
R459 DOWN DOWN.t0 12.0784
C0 UP_b VDDA 0.216714f
C1 opamp_out x 0.402621f
C2 UP_b DOWN 0.043302f
C3 UP_input UP_b 0.207944f
C4 I_IN VDDA 0.091388f
C5 I_IN DOWN 0.011064f
C6 UP_input VDDA 1.17012f
C7 vout VDDA 0.4159f
C8 opamp_out VDDA 0.913816f
C9 x VDDA 0.472127f
C10 DOWN_input DOWN 0.199998f
C11 x I_IN 0.163274f
C12 UP_input DOWN_input 0.110282f
C13 DOWN_input vout 0.305623f
C14 UP_input vout 0.565486f
C15 DOWN GNDA 2.74152f
C16 UP_b GNDA 3.71409f
C17 DOWN_input GNDA 1.43625f
C18 I_IN GNDA 2.77981f
C19 vout GNDA 0.512153f
C20 x GNDA 0.553099f
C21 UP_input GNDA 1.07212f
C22 opamp_out GNDA 0.648776f
C23 VDDA GNDA 7.79453f
.ends

