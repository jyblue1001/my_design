magic
tech sky130A
timestamp 1738230223
<< psubdiff >>
rect 955 1770 1005 1785
rect 955 1750 970 1770
rect 990 1750 1005 1770
rect 955 1735 1005 1750
<< nsubdiff >>
rect 235 840 285 855
rect 235 820 250 840
rect 270 820 285 840
rect 235 805 285 820
<< psubdiffcont >>
rect 970 1750 990 1770
<< nsubdiffcont >>
rect 250 820 270 840
<< poly >>
rect -155 2710 20 2720
rect -155 2690 -145 2710
rect -125 2705 20 2710
rect -125 2690 -115 2705
rect -155 2680 -115 2690
rect -75 2545 -35 2555
rect -75 2525 -65 2545
rect -45 2525 -35 2545
rect -75 2515 -35 2525
rect 90 2545 130 2555
rect 90 2525 100 2545
rect 120 2525 130 2545
rect 90 2515 130 2525
rect -50 1280 -35 2515
rect -50 1265 2925 1280
rect 2910 530 2925 1265
<< polycont >>
rect -145 2690 -125 2710
rect -65 2525 -45 2545
rect 100 2525 120 2545
<< locali >>
rect -155 2710 -115 2720
rect -155 2690 -145 2710
rect -125 2690 -115 2710
rect -155 2680 -115 2690
rect -135 950 -115 2680
rect -75 2545 130 2555
rect -75 2525 -65 2545
rect -45 2530 100 2545
rect -45 2525 -35 2530
rect -75 2515 -35 2525
rect 90 2525 100 2530
rect 120 2525 130 2545
rect 90 2515 130 2525
rect 960 1770 1000 1780
rect 960 1750 970 1770
rect 990 1750 1000 1770
rect 960 1740 1000 1750
rect 2640 1105 2660 2410
rect 2170 1085 2660 1105
rect -135 930 100 950
rect 240 840 280 850
rect 2170 840 2190 1085
rect 240 820 250 840
rect 270 820 280 840
rect 795 820 2190 840
rect 240 810 280 820
<< viali >>
rect 970 1750 990 1770
rect 250 820 270 840
<< metal1 >>
rect 1250 3725 3000 3745
rect 1250 3090 1270 3725
rect 2980 3035 3000 3725
rect 2980 3015 3270 3035
rect 955 1770 1005 1785
rect 955 1750 970 1770
rect 990 1750 1005 1770
rect -400 1725 245 1745
rect 955 1735 1005 1750
rect -400 390 -380 1725
rect 3250 1155 3270 3015
rect 2030 1135 3270 1155
rect -400 370 150 390
use charge_pump_8  charge_pump_8_0
timestamp 1738230159
transform 1 0 1665 0 1 -120
box -1665 120 1245 1275
use opamp_6_6  opamp_6_6_0
timestamp 1738229533
transform 1 0 -725 0 1 2440
box 735 -1145 3385 1090
<< labels >>
flabel metal1 -400 780 -400 780 7 FreeSans 400 0 -200 0 GNDA
flabel metal1 3270 1915 3270 1920 3 FreeSans 400 0 200 0 VDDA
flabel space 100 710 100 710 7 FreeSans 400 0 -200 0 x
flabel poly 2925 540 2925 540 3 FreeSans 400 0 200 0 VOUT
<< end >>
