* PEX produced on Fri Jul 18 10:41:38 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_15.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_15 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t222 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_21_0.Vb3.t4 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_0.V_TOP.t13 VDDA.t431 VDDA.t433 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X2 two_stage_opamp_dummy_magic_21_0.err_amp_out.t7 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t17 GNDA.t130 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 two_stage_opamp_dummy_magic_21_0.V_p_mir.t2 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t12 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X4 GNDA.t10 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t2 VOUT-.t9 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X5 two_stage_opamp_dummy_magic_21_0.VD2.t15 GNDA.t317 GNDA.t318 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X6 VOUT+.t19 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VDDA.t122 bgr_0.V_TOP.t14 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t3 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t14 two_stage_opamp_dummy_magic_21_0.Y.t25 GNDA.t66 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X9 VOUT+.t20 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 VOUT+.t21 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 bgr_0.Vin+.t3 bgr_0.V_TOP.t15 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X12 VDDA.t19 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X13 VOUT+.t22 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VOUT+.t23 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 GNDA.t123 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_21_0.V_source.t26 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X17 two_stage_opamp_dummy_magic_21_0.Y.t3 two_stage_opamp_dummy_magic_21_0.Vb2.t11 two_stage_opamp_dummy_magic_21_0.VD4.t25 two_stage_opamp_dummy_magic_21_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X18 bgr_0.1st_Vout_2.t8 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t4 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X19 VDDA.t144 two_stage_opamp_dummy_magic_21_0.Y.t26 VOUT+.t8 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X20 VOUT+.t24 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VOUT+.t25 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 GNDA.t140 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_21_0.V_source.t25 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X23 a_7460_23988.t1 bgr_0.Vin+.t5 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X24 VDDA.t430 VDDA.t428 VDDA.t430 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X25 two_stage_opamp_dummy_magic_21_0.V_err_p.t11 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_21_0.err_amp_out.t1 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X26 VOUT+.t26 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 two_stage_opamp_dummy_magic_21_0.X.t20 GNDA.t315 GNDA.t316 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X29 VDDA.t427 VDDA.t425 bgr_0.NFET_GATE_10uA.t0 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X30 two_stage_opamp_dummy_magic_21_0.X.t4 two_stage_opamp_dummy_magic_21_0.Vb1.t14 two_stage_opamp_dummy_magic_21_0.VD1.t21 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X31 GNDA.t148 a_6930_22564.t1 GNDA.t113 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X32 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t3 bgr_0.PFET_GATE_10uA.t10 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X33 VDDA.t183 two_stage_opamp_dummy_magic_21_0.X.t25 VOUT-.t4 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X34 VDDA.t64 bgr_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t1 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X35 VOUT-.t19 two_stage_opamp_dummy_magic_21_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VDDA.t212 two_stage_opamp_dummy_magic_21_0.X.t26 VOUT-.t11 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X37 VOUT-.t20 two_stage_opamp_dummy_magic_21_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT-.t21 two_stage_opamp_dummy_magic_21_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT+.t27 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VOUT+.t28 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT+.t29 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 bgr_0.1st_Vout_2.t6 bgr_0.V_mir2.t17 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X44 VDDA.t57 bgr_0.V_TOP.t16 bgr_0.Vin-.t3 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X45 VOUT-.t22 two_stage_opamp_dummy_magic_21_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 bgr_0.1st_Vout_1.t8 bgr_0.Vin+.t6 bgr_0.V_p_1.t10 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X47 two_stage_opamp_dummy_magic_21_0.Y.t19 GNDA.t312 GNDA.t314 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X48 GNDA.t38 VDDA.t469 bgr_0.V_p_2.t10 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X49 VOUT+.t30 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 bgr_0.cap_res2.t0 bgr_0.PFET_GATE_10uA.t0 GNDA.t57 sky130_fd_pr__res_high_po_0p35 l=2.05
X51 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 GNDA.t331 two_stage_opamp_dummy_magic_21_0.X.t27 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t13 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X53 VOUT+.t31 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 VOUT-.t23 two_stage_opamp_dummy_magic_21_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 two_stage_opamp_dummy_magic_21_0.Y.t7 two_stage_opamp_dummy_magic_21_0.Vb2.t12 two_stage_opamp_dummy_magic_21_0.VD4.t23 two_stage_opamp_dummy_magic_21_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X56 VOUT-.t24 two_stage_opamp_dummy_magic_21_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t12 GNDA.t180 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X58 VDDA.t258 bgr_0.1st_Vout_1.t13 bgr_0.V_TOP.t7 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X59 bgr_0.V_TOP.t17 VDDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VOUT-.t25 two_stage_opamp_dummy_magic_21_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_21_0.Y.t27 VDDA.t145 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X62 two_stage_opamp_dummy_magic_21_0.VD1.t2 VIN-.t0 two_stage_opamp_dummy_magic_21_0.V_source.t6 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X63 GNDA.t311 GNDA.t309 bgr_0.NFET_GATE_10uA.t1 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X64 bgr_0.START_UP.t3 bgr_0.V_TOP.t18 VDDA.t435 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X65 VOUT-.t26 two_stage_opamp_dummy_magic_21_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 two_stage_opamp_dummy_magic_21_0.V_err_gate.t11 bgr_0.NFET_GATE_10uA.t6 GNDA.t220 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X67 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t7 bgr_0.V_p_1.t9 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X68 VOUT+.t32 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 VOUT-.t27 two_stage_opamp_dummy_magic_21_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VOUT-.t28 two_stage_opamp_dummy_magic_21_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 VOUT-.t29 two_stage_opamp_dummy_magic_21_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 two_stage_opamp_dummy_magic_21_0.V_source.t24 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t15 GNDA.t142 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X73 two_stage_opamp_dummy_magic_21_0.VD3.t35 two_stage_opamp_dummy_magic_21_0.Vb3.t8 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X74 VOUT+.t33 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 two_stage_opamp_dummy_magic_21_0.VD2.t0 VIN+.t0 two_stage_opamp_dummy_magic_21_0.V_source.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X77 bgr_0.V_TOP.t19 VDDA.t436 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t272 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t16 VDDA.t422 VDDA.t424 VDDA.t423 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X80 VOUT-.t30 two_stage_opamp_dummy_magic_21_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t2 bgr_0.PFET_GATE_10uA.t12 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X82 VDDA.t126 bgr_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t3 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X83 two_stage_opamp_dummy_magic_21_0.Vb2_2.t8 two_stage_opamp_dummy_magic_21_0.Vb2.t13 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X84 VOUT+.t34 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 bgr_0.V_TOP.t20 VDDA.t437 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 GNDA.t50 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_21_0.V_source.t23 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X87 bgr_0.1st_Vout_2.t1 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t3 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X88 VDDA.t421 VDDA.t419 two_stage_opamp_dummy_magic_21_0.V_err_p.t20 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X89 VDDA.t35 two_stage_opamp_dummy_magic_21_0.Y.t28 VOUT+.t2 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X90 VDDA.t418 VDDA.t416 VOUT+.t18 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X91 two_stage_opamp_dummy_magic_21_0.V_err_p.t0 two_stage_opamp_dummy_magic_21_0.V_tot.t4 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t0 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X92 GNDA.t308 GNDA.t307 two_stage_opamp_dummy_magic_21_0.VD1.t9 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X93 VOUT-.t31 two_stage_opamp_dummy_magic_21_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 VOUT-.t32 two_stage_opamp_dummy_magic_21_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 VOUT+.t35 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT-.t33 two_stage_opamp_dummy_magic_21_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 two_stage_opamp_dummy_magic_21_0.X.t1 two_stage_opamp_dummy_magic_21_0.Vb1.t15 two_stage_opamp_dummy_magic_21_0.VD1.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X98 two_stage_opamp_dummy_magic_21_0.VD3.t25 two_stage_opamp_dummy_magic_21_0.VD3.t23 two_stage_opamp_dummy_magic_21_0.X.t17 two_stage_opamp_dummy_magic_21_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X99 VOUT+.t36 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 VOUT+.t9 a_5710_2046.t1 GNDA.t136 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X101 two_stage_opamp_dummy_magic_21_0.VD3.t34 two_stage_opamp_dummy_magic_21_0.Vb3.t9 VDDA.t312 VDDA.t311 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X102 VDDA.t467 two_stage_opamp_dummy_magic_21_0.X.t28 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t9 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X103 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t0 a_14240_2056.t0 GNDA.t48 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X104 bgr_0.PFET_GATE_10uA.t9 bgr_0.1st_Vout_2.t13 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X105 GNDA.t306 GNDA.t305 two_stage_opamp_dummy_magic_21_0.VD2.t14 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X106 VOUT-.t34 two_stage_opamp_dummy_magic_21_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 bgr_0.V_TOP.t21 VDDA.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t157 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X109 two_stage_opamp_dummy_magic_21_0.Y.t0 two_stage_opamp_dummy_magic_21_0.Vb1.t16 two_stage_opamp_dummy_magic_21_0.VD2.t3 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X110 a_5190_5068.t1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t0 GNDA.t128 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X111 GNDA.t133 two_stage_opamp_dummy_magic_21_0.X.t29 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t12 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X112 a_14560_4968.t1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t14 GNDA.t339 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X113 VOUT+.t37 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 bgr_0.V_TOP.t22 VDDA.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 GNDA.t218 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t12 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t11 bgr_0.NFET_GATE_10uA.t8 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X117 two_stage_opamp_dummy_magic_21_0.err_amp_out.t2 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_21_0.V_err_p.t10 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X118 VOUT-.t35 two_stage_opamp_dummy_magic_21_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT-.t36 two_stage_opamp_dummy_magic_21_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT-.t37 two_stage_opamp_dummy_magic_21_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 VOUT-.t38 two_stage_opamp_dummy_magic_21_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT-.t39 two_stage_opamp_dummy_magic_21_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 GNDA.t304 GNDA.t302 two_stage_opamp_dummy_magic_21_0.X.t19 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X125 VOUT+.t38 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT+.t39 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_21_0.Y.t29 VDDA.t36 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X128 VOUT+.t40 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 two_stage_opamp_dummy_magic_21_0.V_err_gate.t9 two_stage_opamp_dummy_magic_21_0.V_tot.t5 a_8570_6900.t4 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X130 VOUT+.t41 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 two_stage_opamp_dummy_magic_21_0.V_err_p.t19 VDDA.t413 VDDA.t415 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X132 VOUT+.t42 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 a_12530_23988.t1 bgr_0.Vin-.t7 GNDA.t335 sky130_fd_pr__res_xhigh_po_0p35 l=6
X134 two_stage_opamp_dummy_magic_21_0.V_source.t22 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t17 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X135 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t13 two_stage_opamp_dummy_magic_21_0.Y.t30 GNDA.t7 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X136 GNDA.t301 GNDA.t299 two_stage_opamp_dummy_magic_21_0.Y.t18 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X137 two_stage_opamp_dummy_magic_21_0.VD4.t37 VDDA.t410 VDDA.t412 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X138 bgr_0.1st_Vout_2.t9 bgr_0.V_mir2.t18 VDDA.t240 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X139 two_stage_opamp_dummy_magic_21_0.VD4.t21 two_stage_opamp_dummy_magic_21_0.Vb2.t14 two_stage_opamp_dummy_magic_21_0.Y.t24 two_stage_opamp_dummy_magic_21_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X140 VOUT-.t40 two_stage_opamp_dummy_magic_21_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 GNDA.t32 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_21_0.V_source.t21 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X142 VDDA.t16 two_stage_opamp_dummy_magic_21_0.V_err_gate.t14 two_stage_opamp_dummy_magic_21_0.V_err_p.t3 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X143 VOUT-.t41 two_stage_opamp_dummy_magic_21_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 two_stage_opamp_dummy_magic_21_0.VD3.t33 two_stage_opamp_dummy_magic_21_0.Vb3.t10 VDDA.t310 VDDA.t309 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X146 VDDA.t109 two_stage_opamp_dummy_magic_21_0.V_err_gate.t15 a_8570_6900.t19 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X147 VDDA.t409 VDDA.t406 VDDA.t408 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X148 VOUT-.t42 two_stage_opamp_dummy_magic_21_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t43 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VDDA.t10 two_stage_opamp_dummy_magic_21_0.Y.t31 VOUT+.t0 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X151 two_stage_opamp_dummy_magic_21_0.V_source.t40 VIN-.t1 two_stage_opamp_dummy_magic_21_0.VD1.t11 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X152 VOUT-.t43 two_stage_opamp_dummy_magic_21_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT+.t44 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VOUT+.t45 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 bgr_0.V_mir1.t3 bgr_0.Vin-.t8 bgr_0.V_p_1.t4 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X157 bgr_0.V_mir1.t15 bgr_0.V_mir1.t14 VDDA.t453 VDDA.t452 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X158 GNDA.t34 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_21_0.V_source.t20 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X159 a_14680_4968.t0 two_stage_opamp_dummy_magic_21_0.V_tot.t1 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X160 VDDA.t199 two_stage_opamp_dummy_magic_21_0.X.t30 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t8 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X161 GNDA.t332 a_7580_22380.t1 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X162 GNDA.t160 two_stage_opamp_dummy_magic_21_0.Y.t32 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t12 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X163 two_stage_opamp_dummy_magic_21_0.V_source.t37 VIN+.t1 two_stage_opamp_dummy_magic_21_0.VD2.t17 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X164 VOUT-.t44 two_stage_opamp_dummy_magic_21_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT-.t45 two_stage_opamp_dummy_magic_21_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+.t46 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT-.t46 two_stage_opamp_dummy_magic_21_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VOUT-.t47 two_stage_opamp_dummy_magic_21_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VDDA.t104 bgr_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_21_0.Vb1.t1 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X170 VOUT-.t48 two_stage_opamp_dummy_magic_21_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 two_stage_opamp_dummy_magic_21_0.VD4.t19 two_stage_opamp_dummy_magic_21_0.Vb2.t15 two_stage_opamp_dummy_magic_21_0.Y.t16 two_stage_opamp_dummy_magic_21_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X172 two_stage_opamp_dummy_magic_21_0.Vb1.t11 two_stage_opamp_dummy_magic_21_0.Vb1.t10 a_9370_2200.t4 GNDA.t327 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X173 GNDA.t330 two_stage_opamp_dummy_magic_21_0.X.t31 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t11 VDDA.t456 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X174 bgr_0.V_TOP.t23 VDDA.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VDDA.t405 VDDA.t403 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t15 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X176 GNDA.t336 two_stage_opamp_dummy_magic_21_0.X.t32 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t10 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X177 VOUT-.t49 two_stage_opamp_dummy_magic_21_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VOUT-.t50 two_stage_opamp_dummy_magic_21_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 two_stage_opamp_dummy_magic_21_0.V_source.t19 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t20 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X180 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t3 bgr_0.PFET_GATE_10uA.t15 VDDA.t98 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X181 VOUT+.t47 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT+.t48 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 bgr_0.V_mir1.t16 bgr_0.Vin-.t9 bgr_0.V_p_1.t3 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X184 VOUT+.t49 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 two_stage_opamp_dummy_magic_21_0.Vb2.t10 two_stage_opamp_dummy_magic_21_0.Vb2_2.t3 two_stage_opamp_dummy_magic_21_0.Vb2_2.t5 two_stage_opamp_dummy_magic_21_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X186 VOUT+.t50 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 two_stage_opamp_dummy_magic_21_0.VD1.t19 two_stage_opamp_dummy_magic_21_0.Vb1.t17 two_stage_opamp_dummy_magic_21_0.X.t2 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X188 VDDA.t308 two_stage_opamp_dummy_magic_21_0.Vb3.t11 two_stage_opamp_dummy_magic_21_0.VD3.t32 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X189 VOUT-.t3 two_stage_opamp_dummy_magic_21_0.X.t33 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X190 bgr_0.START_UP.t2 bgr_0.V_TOP.t24 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X191 bgr_0.PFET_GATE_10uA.t8 bgr_0.1st_Vout_2.t16 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X192 VDDA.t42 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t4 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X193 two_stage_opamp_dummy_magic_21_0.V_err_gate.t7 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t9 a_8570_6900.t9 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X194 VOUT+.t51 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT-.t51 two_stage_opamp_dummy_magic_21_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 a_8570_6900.t18 two_stage_opamp_dummy_magic_21_0.V_err_gate.t16 VDDA.t140 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X197 VOUT-.t52 two_stage_opamp_dummy_magic_21_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 two_stage_opamp_dummy_magic_21_0.V_source.t18 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t21 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X199 two_stage_opamp_dummy_magic_21_0.Vb2.t7 bgr_0.NFET_GATE_10uA.t9 GNDA.t214 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X200 two_stage_opamp_dummy_magic_21_0.VD2.t7 two_stage_opamp_dummy_magic_21_0.Vb1.t18 two_stage_opamp_dummy_magic_21_0.Y.t4 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X201 GNDA.t212 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_21_0.Vb2.t6 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X202 VDDA.t402 VDDA.t400 two_stage_opamp_dummy_magic_21_0.Vb2_2.t9 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X203 VOUT+.t52 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 bgr_0.V_TOP.t25 VDDA.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 GNDA.t210 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_21_0.Vb2.t5 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X206 VOUT+.t53 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT-.t53 two_stage_opamp_dummy_magic_21_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+.t54 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT+.t55 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VDDA.t244 two_stage_opamp_dummy_magic_21_0.V_err_gate.t17 a_8570_6900.t17 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X211 VOUT+.t56 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 GNDA.t97 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_21_0.V_source.t17 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X213 VDDA.t120 bgr_0.V_TOP.t26 bgr_0.Vin+.t2 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X214 VDDA.t221 two_stage_opamp_dummy_magic_21_0.Y.t33 VOUT+.t14 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X215 bgr_0.1st_Vout_2.t10 bgr_0.V_mir2.t19 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X216 VDDA.t306 two_stage_opamp_dummy_magic_21_0.Vb3.t12 two_stage_opamp_dummy_magic_21_0.VD3.t31 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X217 bgr_0.V_TOP.t6 bgr_0.1st_Vout_1.t16 VDDA.t256 VDDA.t255 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X218 bgr_0.V_CUR_REF_REG.t2 VDDA.t397 VDDA.t399 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X219 two_stage_opamp_dummy_magic_21_0.VD4.t5 two_stage_opamp_dummy_magic_21_0.VD4.t3 two_stage_opamp_dummy_magic_21_0.Y.t11 two_stage_opamp_dummy_magic_21_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X220 VOUT-.t54 two_stage_opamp_dummy_magic_21_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 VOUT-.t55 two_stage_opamp_dummy_magic_21_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT-.t56 two_stage_opamp_dummy_magic_21_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT+.t57 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t2 bgr_0.PFET_GATE_10uA.t16 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X225 VOUT-.t57 two_stage_opamp_dummy_magic_21_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VOUT+.t13 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t3 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X227 two_stage_opamp_dummy_magic_21_0.V_source.t28 VIN+.t2 two_stage_opamp_dummy_magic_21_0.VD2.t5 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X228 VOUT+.t58 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 GNDA.t111 two_stage_opamp_dummy_magic_21_0.Y.t34 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t11 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X230 VDDA.t455 two_stage_opamp_dummy_magic_21_0.X.t34 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t7 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X231 two_stage_opamp_dummy_magic_21_0.V_source.t29 VIN+.t3 two_stage_opamp_dummy_magic_21_0.VD2.t6 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X232 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t10 GNDA.t297 GNDA.t298 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X233 VOUT+.t59 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 a_14680_4968.t1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t16 GNDA.t338 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X235 VOUT+.t60 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 a_6810_23838.t1 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t6 GNDA.t113 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X238 bgr_0.Vin+.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t62 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X239 GNDA.t143 VDDA.t394 VDDA.t396 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X240 two_stage_opamp_dummy_magic_21_0.Vb1.t7 two_stage_opamp_dummy_magic_21_0.Vb1.t6 a_9370_2200.t3 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X241 VOUT+.t61 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 VOUT+.t62 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 VOUT-.t58 two_stage_opamp_dummy_magic_21_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT-.t59 two_stage_opamp_dummy_magic_21_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 bgr_0.Vin+.t1 bgr_0.V_TOP.t27 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X247 VDDA.t393 VDDA.t391 bgr_0.PFET_GATE_10uA.t3 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X248 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t3 two_stage_opamp_dummy_magic_21_0.V_tot.t6 two_stage_opamp_dummy_magic_21_0.V_err_p.t15 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X249 VOUT+.t63 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VDDA.t77 bgr_0.V_TOP.t28 bgr_0.Vin+.t0 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X251 VOUT+.t64 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 GNDA.t54 a_12410_22380.t0 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X254 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_21_0.Y.t35 VDDA.t138 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X255 GNDA.t208 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_21_0.Vb3.t7 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X256 VOUT-.t60 two_stage_opamp_dummy_magic_21_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 VOUT-.t61 two_stage_opamp_dummy_magic_21_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VOUT-.t18 two_stage_opamp_dummy_magic_21_0.X.t35 VDDA.t463 VDDA.t462 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X259 VOUT+.t65 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 two_stage_opamp_dummy_magic_21_0.V_err_gate.t4 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t10 a_8570_6900.t8 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X261 VOUT+.t66 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VOUT-.t62 two_stage_opamp_dummy_magic_21_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 bgr_0.cap_res1.t20 bgr_0.V_TOP.t1 GNDA.t150 sky130_fd_pr__res_high_po_0p35 l=2.05
X264 two_stage_opamp_dummy_magic_21_0.Vb3.t6 bgr_0.NFET_GATE_10uA.t13 GNDA.t206 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X265 bgr_0.V_mir2.t9 bgr_0.V_mir2.t8 VDDA.t268 VDDA.t267 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X266 VOUT-.t63 two_stage_opamp_dummy_magic_21_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VDDA.t304 two_stage_opamp_dummy_magic_21_0.Vb3.t13 two_stage_opamp_dummy_magic_21_0.VD4.t35 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X268 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t11 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t10 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X269 VDDA.t390 VDDA.t388 bgr_0.V_TOP.t12 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X270 VOUT+.t67 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 VOUT+.t68 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 two_stage_opamp_dummy_magic_21_0.V_err_p.t5 two_stage_opamp_dummy_magic_21_0.V_err_gate.t18 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X273 two_stage_opamp_dummy_magic_21_0.VD2.t9 two_stage_opamp_dummy_magic_21_0.Vb1.t19 two_stage_opamp_dummy_magic_21_0.Y.t6 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X274 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 two_stage_opamp_dummy_magic_21_0.Y.t17 two_stage_opamp_dummy_magic_21_0.Vb2.t16 two_stage_opamp_dummy_magic_21_0.VD4.t17 two_stage_opamp_dummy_magic_21_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X276 two_stage_opamp_dummy_magic_21_0.VD2.t19 two_stage_opamp_dummy_magic_21_0.Vb1.t20 two_stage_opamp_dummy_magic_21_0.Y.t20 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X277 VOUT-.t64 two_stage_opamp_dummy_magic_21_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VOUT+.t69 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t2 bgr_0.V_TOP.t29 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X280 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 VOUT-.t65 two_stage_opamp_dummy_magic_21_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 GNDA.t326 a_13060_22630.t0 GNDA.t325 sky130_fd_pr__res_xhigh_po_0p35 l=4
X283 VDDA.t387 VDDA.t385 two_stage_opamp_dummy_magic_21_0.VD3.t37 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X284 VOUT+.t70 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 GNDA.t296 GNDA.t294 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t14 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X286 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t19 VDDA.t461 VDDA.t460 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X287 VDDA.t246 two_stage_opamp_dummy_magic_21_0.V_err_gate.t19 two_stage_opamp_dummy_magic_21_0.V_err_p.t18 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X288 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t8 VIN-.t2 two_stage_opamp_dummy_magic_21_0.V_p_mir.t3 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X290 two_stage_opamp_dummy_magic_21_0.V_source.t5 VIN-.t3 two_stage_opamp_dummy_magic_21_0.VD1.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X291 VOUT-.t66 two_stage_opamp_dummy_magic_21_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VDDA.t217 two_stage_opamp_dummy_magic_21_0.Y.t36 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t7 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X293 VOUT+.t71 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VOUT-.t67 two_stage_opamp_dummy_magic_21_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 VOUT-.t68 two_stage_opamp_dummy_magic_21_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 a_14560_4968.t0 two_stage_opamp_dummy_magic_21_0.V_tot.t2 GNDA.t127 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X297 bgr_0.NFET_GATE_10uA.t4 bgr_0.PFET_GATE_10uA.t17 VDDA.t459 VDDA.t458 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X298 GNDA.t152 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t4 VOUT-.t8 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X299 VDDA.t465 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t11 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X300 VOUT+.t72 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT+.t73 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 bgr_0.V_p_2.t5 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t11 bgr_0.V_mir2.t16 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X304 VDDA.t302 two_stage_opamp_dummy_magic_21_0.Vb3.t14 two_stage_opamp_dummy_magic_21_0.VD4.t34 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X305 VDDA.t150 two_stage_opamp_dummy_magic_21_0.X.t36 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t6 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X306 VDDA.t206 two_stage_opamp_dummy_magic_21_0.V_err_gate.t20 two_stage_opamp_dummy_magic_21_0.V_err_p.t16 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X307 two_stage_opamp_dummy_magic_21_0.V_source.t38 VIN+.t4 two_stage_opamp_dummy_magic_21_0.VD2.t18 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X308 two_stage_opamp_dummy_magic_21_0.Y.t2 two_stage_opamp_dummy_magic_21_0.Vb2.t17 two_stage_opamp_dummy_magic_21_0.VD4.t15 two_stage_opamp_dummy_magic_21_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X309 GNDA.t159 two_stage_opamp_dummy_magic_21_0.Y.t37 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t10 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X310 VDDA.t157 two_stage_opamp_dummy_magic_21_0.X.t37 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t5 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X311 VDDA.t232 bgr_0.V_TOP.t30 bgr_0.START_UP.t1 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X312 GNDA.t22 two_stage_opamp_dummy_magic_21_0.Y.t38 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t9 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X313 VOUT+.t74 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VOUT-.t69 two_stage_opamp_dummy_magic_21_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT-.t70 two_stage_opamp_dummy_magic_21_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT+.t75 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VOUT+.t76 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 bgr_0.V_TOP.t31 VDDA.t233 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 bgr_0.V_TOP.t4 bgr_0.1st_Vout_1.t21 VDDA.t252 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X320 two_stage_opamp_dummy_magic_21_0.Vb1.t3 GNDA.t291 GNDA.t293 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X321 two_stage_opamp_dummy_magic_21_0.Vb2_2.t7 two_stage_opamp_dummy_magic_21_0.Vb2.t0 two_stage_opamp_dummy_magic_21_0.Vb2.t1 two_stage_opamp_dummy_magic_21_0.Vb2_2.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X322 a_8570_6900.t16 two_stage_opamp_dummy_magic_21_0.V_err_gate.t21 VDDA.t451 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X323 GNDA.t290 GNDA.t288 VOUT-.t14 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X324 two_stage_opamp_dummy_magic_21_0.err_amp_out.t10 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_21_0.V_err_p.t9 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X325 VOUT+.t77 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT-.t71 two_stage_opamp_dummy_magic_21_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VOUT-.t72 two_stage_opamp_dummy_magic_21_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT-.t73 two_stage_opamp_dummy_magic_21_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT-.t74 two_stage_opamp_dummy_magic_21_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 bgr_0.V_TOP.t5 bgr_0.1st_Vout_1.t22 VDDA.t254 VDDA.t253 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X331 two_stage_opamp_dummy_magic_21_0.VD1.t18 two_stage_opamp_dummy_magic_21_0.Vb1.t21 two_stage_opamp_dummy_magic_21_0.X.t0 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X332 VOUT+.t78 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VOUT+.t79 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT+.t80 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 bgr_0.NFET_GATE_10uA.t3 bgr_0.NFET_GATE_10uA.t2 GNDA.t204 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X336 GNDA.t26 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t5 VOUT+.t12 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X337 GNDA.t202 bgr_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_21_0.Vb3.t5 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X338 two_stage_opamp_dummy_magic_21_0.V_err_gate.t2 two_stage_opamp_dummy_magic_21_0.V_tot.t7 a_8570_6900.t3 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X339 VOUT-.t17 two_stage_opamp_dummy_magic_21_0.X.t38 VDDA.t445 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X340 VOUT+.t81 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 bgr_0.V_TOP.t32 VDDA.t234 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 two_stage_opamp_dummy_magic_21_0.err_amp_out.t8 GNDA.t285 GNDA.t287 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X343 two_stage_opamp_dummy_magic_21_0.VD3.t19 two_stage_opamp_dummy_magic_21_0.Vb2.t18 two_stage_opamp_dummy_magic_21_0.X.t14 two_stage_opamp_dummy_magic_21_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X344 a_8570_6900.t15 two_stage_opamp_dummy_magic_21_0.V_err_gate.t22 VDDA.t248 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X345 two_stage_opamp_dummy_magic_21_0.VD2.t11 two_stage_opamp_dummy_magic_21_0.Vb1.t22 two_stage_opamp_dummy_magic_21_0.Y.t12 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X346 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VOUT-.t75 two_stage_opamp_dummy_magic_21_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT-.t76 two_stage_opamp_dummy_magic_21_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT+.t82 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VDDA.t384 VDDA.t382 GNDA.t182 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X351 VDDA.t159 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t4 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X352 VOUT-.t77 two_stage_opamp_dummy_magic_21_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 bgr_0.V_mir1.t13 bgr_0.V_mir1.t12 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X355 GNDA.t93 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t18 two_stage_opamp_dummy_magic_21_0.err_amp_out.t6 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X356 GNDA.t101 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t6 VOUT+.t11 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X357 VDDA.t228 bgr_0.V_TOP.t33 bgr_0.START_UP.t0 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X358 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_21_0.Y.t21 GNDA.t324 sky130_fd_pr__res_high_po_1p41 l=1.41
X359 VOUT-.t78 two_stage_opamp_dummy_magic_21_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 VDDA.t300 two_stage_opamp_dummy_magic_21_0.Vb3.t15 two_stage_opamp_dummy_magic_21_0.VD4.t33 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X362 VDDA.t447 two_stage_opamp_dummy_magic_21_0.V_err_gate.t23 a_8570_6900.t14 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X363 VOUT-.t79 two_stage_opamp_dummy_magic_21_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VDDA.t33 two_stage_opamp_dummy_magic_21_0.Y.t39 VOUT+.t1 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X365 VOUT+.t83 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 VOUT+.t84 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 two_stage_opamp_dummy_magic_21_0.V_source.t39 VIN-.t4 two_stage_opamp_dummy_magic_21_0.VD1.t10 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X368 VOUT+.t85 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 a_7460_23988.t0 a_7580_22380.t0 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X370 bgr_0.V_p_2.t2 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t2 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X371 VDDA.t89 two_stage_opamp_dummy_magic_21_0.Y.t40 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t6 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X372 VOUT-.t80 two_stage_opamp_dummy_magic_21_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VDDA.t318 GNDA.t282 GNDA.t284 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X374 two_stage_opamp_dummy_magic_21_0.V_source.t36 VIN+.t5 two_stage_opamp_dummy_magic_21_0.VD2.t16 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X375 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 GNDA.t65 two_stage_opamp_dummy_magic_21_0.Y.t41 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t8 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X377 bgr_0.1st_Vout_1.t6 bgr_0.Vin+.t8 bgr_0.V_p_1.t8 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X378 VDDA.t7 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X379 VOUT-.t81 two_stage_opamp_dummy_magic_21_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VOUT-.t82 two_stage_opamp_dummy_magic_21_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 GNDA.t230 GNDA.t232 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X383 VOUT-.t83 two_stage_opamp_dummy_magic_21_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VOUT-.t84 two_stage_opamp_dummy_magic_21_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 GNDA.t200 bgr_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_21_0.Vb2.t4 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X387 two_stage_opamp_dummy_magic_21_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t16 GNDA.t198 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X388 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t13 GNDA.t279 GNDA.t281 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X389 VOUT+.t86 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 two_stage_opamp_dummy_magic_21_0.V_source.t8 two_stage_opamp_dummy_magic_21_0.err_amp_out.t12 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X391 GNDA.t227 GNDA.t266 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X392 GNDA.t265 GNDA.t263 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t14 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X393 GNDA.t269 GNDA.t267 two_stage_opamp_dummy_magic_21_0.Vb2.t9 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X394 VOUT+.t7 two_stage_opamp_dummy_magic_21_0.Y.t42 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X395 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t15 VDDA.t379 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X396 VOUT-.t85 two_stage_opamp_dummy_magic_21_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t16 two_stage_opamp_dummy_magic_21_0.V_tot.t8 two_stage_opamp_dummy_magic_21_0.V_err_p.t21 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X398 VOUT+.t87 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 bgr_0.PFET_GATE_10uA.t2 VDDA.t376 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X400 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t20 VDDA.t264 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X401 VOUT-.t13 GNDA.t276 GNDA.t278 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X402 two_stage_opamp_dummy_magic_21_0.VD1.t17 two_stage_opamp_dummy_magic_21_0.Vb1.t23 two_stage_opamp_dummy_magic_21_0.X.t24 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X403 VOUT-.t86 two_stage_opamp_dummy_magic_21_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 two_stage_opamp_dummy_magic_21_0.VD4.t32 two_stage_opamp_dummy_magic_21_0.Vb3.t16 VDDA.t298 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X405 VOUT-.t0 two_stage_opamp_dummy_magic_21_0.X.t39 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X406 bgr_0.V_p_2.t1 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t3 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X407 two_stage_opamp_dummy_magic_21_0.VD4.t13 two_stage_opamp_dummy_magic_21_0.Vb2.t19 two_stage_opamp_dummy_magic_21_0.Y.t15 two_stage_opamp_dummy_magic_21_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X408 two_stage_opamp_dummy_magic_21_0.V_err_gate.t13 VDDA.t373 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X409 VOUT-.t2 two_stage_opamp_dummy_magic_21_0.X.t40 VDDA.t81 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X410 VOUT-.t87 two_stage_opamp_dummy_magic_21_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VOUT+.t88 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 GNDA.t227 GNDA.t275 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X413 VOUT-.t88 two_stage_opamp_dummy_magic_21_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 two_stage_opamp_dummy_magic_21_0.VD2.t4 two_stage_opamp_dummy_magic_21_0.Vb1.t24 two_stage_opamp_dummy_magic_21_0.Y.t1 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X415 VOUT+.t89 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 GNDA.t227 GNDA.t274 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X417 VOUT-.t89 two_stage_opamp_dummy_magic_21_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_21_0.X.t41 GNDA.t138 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X419 VDDA.t242 bgr_0.V_mir2.t6 bgr_0.V_mir2.t7 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X420 VOUT+.t90 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+.t91 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 GNDA.t155 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t9 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X423 bgr_0.V_p_2.t0 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t4 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X424 VOUT+.t92 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VDDA.t136 two_stage_opamp_dummy_magic_21_0.Y.t43 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t5 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X426 two_stage_opamp_dummy_magic_21_0.V_source.t1 VIN-.t5 two_stage_opamp_dummy_magic_21_0.VD1.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X427 a_13180_23838.t0 bgr_0.V_CUR_REF_REG.t1 GNDA.t126 sky130_fd_pr__res_xhigh_po_0p35 l=4
X428 two_stage_opamp_dummy_magic_21_0.VD4.t31 two_stage_opamp_dummy_magic_21_0.Vb3.t17 VDDA.t296 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X429 VDDA.t86 two_stage_opamp_dummy_magic_21_0.Y.t44 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t4 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X430 VOUT-.t90 two_stage_opamp_dummy_magic_21_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 bgr_0.V_TOP.t34 VDDA.t229 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_21_0.X.t3 two_stage_opamp_dummy_magic_21_0.VD3.t20 two_stage_opamp_dummy_magic_21_0.VD3.t22 two_stage_opamp_dummy_magic_21_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X433 VOUT-.t91 two_stage_opamp_dummy_magic_21_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT-.t92 two_stage_opamp_dummy_magic_21_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 GNDA.t56 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t6 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t7 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X436 VOUT-.t93 two_stage_opamp_dummy_magic_21_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT-.t94 two_stage_opamp_dummy_magic_21_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 GNDA.t273 GNDA.t270 GNDA.t272 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X439 VOUT-.t95 two_stage_opamp_dummy_magic_21_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 GNDA.t99 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_21_0.V_source.t16 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X441 VOUT+.t93 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 bgr_0.V_TOP.t35 VDDA.t230 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 VDDA.t167 bgr_0.1st_Vout_2.t24 bgr_0.PFET_GATE_10uA.t7 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X444 VDDA.t372 VDDA.t370 two_stage_opamp_dummy_magic_21_0.Vb1.t5 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X445 VOUT+.t94 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 two_stage_opamp_dummy_magic_21_0.Vb1.t4 VDDA.t367 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X447 two_stage_opamp_dummy_magic_21_0.Vb2_2.t2 two_stage_opamp_dummy_magic_21_0.Vb2_2.t0 two_stage_opamp_dummy_magic_21_0.Vb2_2.t2 two_stage_opamp_dummy_magic_21_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X448 VOUT-.t96 two_stage_opamp_dummy_magic_21_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VOUT+.t95 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 two_stage_opamp_dummy_magic_21_0.VD4.t30 two_stage_opamp_dummy_magic_21_0.Vb3.t18 VDDA.t294 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X451 VOUT+.t96 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t2 bgr_0.PFET_GATE_10uA.t20 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X453 VOUT-.t97 two_stage_opamp_dummy_magic_21_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VOUT-.t98 two_stage_opamp_dummy_magic_21_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VDDA.t62 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t1 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X456 two_stage_opamp_dummy_magic_21_0.V_source.t15 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t24 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X457 VOUT+.t6 two_stage_opamp_dummy_magic_21_0.Y.t45 VDDA.t88 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X458 two_stage_opamp_dummy_magic_21_0.err_amp_out.t11 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_21_0.V_err_p.t8 VDDA.t439 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X459 VOUT-.t99 two_stage_opamp_dummy_magic_21_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 bgr_0.V_TOP.t36 VDDA.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VOUT-.t100 two_stage_opamp_dummy_magic_21_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 two_stage_opamp_dummy_magic_21_0.X.t11 two_stage_opamp_dummy_magic_21_0.Vb2.t20 two_stage_opamp_dummy_magic_21_0.VD3.t17 two_stage_opamp_dummy_magic_21_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X463 VOUT-.t16 VDDA.t364 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X464 two_stage_opamp_dummy_magic_21_0.VD1.t16 two_stage_opamp_dummy_magic_21_0.Vb1.t25 two_stage_opamp_dummy_magic_21_0.X.t22 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X465 bgr_0.Vin-.t2 bgr_0.V_TOP.t37 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X466 VOUT-.t101 two_stage_opamp_dummy_magic_21_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 two_stage_opamp_dummy_magic_21_0.V_err_gate.t1 two_stage_opamp_dummy_magic_21_0.V_tot.t9 a_8570_6900.t2 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X468 GNDA.t262 GNDA.t260 VDDA.t317 GNDA.t261 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X469 VOUT+.t97 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VOUT+.t98 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT+.t99 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 GNDA.t196 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t13 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X473 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t260 VDDA.t259 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X474 two_stage_opamp_dummy_magic_21_0.Vb2.t8 GNDA.t257 GNDA.t259 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X475 VOUT+.t100 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VOUT+.t101 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VOUT-.t102 two_stage_opamp_dummy_magic_21_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 two_stage_opamp_dummy_magic_21_0.VD4.t29 two_stage_opamp_dummy_magic_21_0.Vb3.t19 VDDA.t292 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X481 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_21_0.X.t42 GNDA.t132 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X482 VOUT+.t102 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VDDA.t363 VDDA.t361 two_stage_opamp_dummy_magic_21_0.err_amp_out.t9 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X484 GNDA.t95 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_21_0.err_amp_out.t5 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X485 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 VOUT-.t103 two_stage_opamp_dummy_magic_21_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT-.t104 two_stage_opamp_dummy_magic_21_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VOUT-.t105 two_stage_opamp_dummy_magic_21_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 two_stage_opamp_dummy_magic_21_0.V_source.t27 VIN-.t6 two_stage_opamp_dummy_magic_21_0.VD1.t4 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X490 VDDA.t45 two_stage_opamp_dummy_magic_21_0.Y.t46 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t3 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X491 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t4 bgr_0.PFET_GATE_10uA.t22 VDDA.t185 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X492 VOUT-.t106 two_stage_opamp_dummy_magic_21_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t1 bgr_0.V_TOP.t38 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X494 VOUT+.t103 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VDDA.t163 bgr_0.V_mir2.t4 bgr_0.V_mir2.t5 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X496 VDDA.t360 VDDA.t358 two_stage_opamp_dummy_magic_21_0.V_err_gate.t12 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X497 VOUT+.t104 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 VDDA.t60 bgr_0.V_mir1.t10 bgr_0.V_mir1.t11 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X499 VDDA.t201 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t5 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X500 bgr_0.V_p_1.t2 bgr_0.Vin-.t10 bgr_0.V_mir1.t1 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X501 GNDA.t61 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_21_0.V_source.t14 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X502 VOUT+.t105 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 VOUT+.t106 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 bgr_0.V_TOP.t11 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X507 two_stage_opamp_dummy_magic_21_0.X.t13 two_stage_opamp_dummy_magic_21_0.Vb2.t21 two_stage_opamp_dummy_magic_21_0.VD3.t15 two_stage_opamp_dummy_magic_21_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X508 VOUT+.t107 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT-.t107 two_stage_opamp_dummy_magic_21_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 two_stage_opamp_dummy_magic_21_0.V_source.t13 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t26 GNDA.t68 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X512 VDDA.t354 VDDA.t352 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t5 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X513 VDDA.t290 two_stage_opamp_dummy_magic_21_0.Vb3.t20 two_stage_opamp_dummy_magic_21_0.VD3.t30 VDDA.t289 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X514 VOUT+.t3 two_stage_opamp_dummy_magic_21_0.Y.t47 VDDA.t47 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X515 two_stage_opamp_dummy_magic_21_0.V_err_p.t1 two_stage_opamp_dummy_magic_21_0.V_err_gate.t24 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X516 VOUT-.t108 two_stage_opamp_dummy_magic_21_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VDDA.t288 two_stage_opamp_dummy_magic_21_0.Vb3.t21 two_stage_opamp_dummy_magic_21_0.VD4.t28 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X518 VOUT+.t4 two_stage_opamp_dummy_magic_21_0.Y.t48 VDDA.t83 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X519 VOUT-.t109 two_stage_opamp_dummy_magic_21_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 two_stage_opamp_dummy_magic_21_0.VD1.t7 VIN-.t7 two_stage_opamp_dummy_magic_21_0.V_source.t34 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X521 bgr_0.V_p_1.t1 bgr_0.Vin-.t11 bgr_0.V_mir1.t2 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X522 VOUT+.t108 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VOUT+.t109 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 VOUT-.t110 two_stage_opamp_dummy_magic_21_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VOUT+.t110 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 VOUT+.t111 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 VOUT+.t112 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 two_stage_opamp_dummy_magic_21_0.Vb3.t2 GNDA.t254 GNDA.t256 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X530 VOUT+.t113 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 two_stage_opamp_dummy_magic_21_0.VD1.t15 two_stage_opamp_dummy_magic_21_0.Vb1.t26 two_stage_opamp_dummy_magic_21_0.X.t23 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X532 bgr_0.Vin-.t4 bgr_0.START_UP.t6 bgr_0.V_TOP.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X533 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X534 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_21_0.X.t43 VDDA.t235 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X535 bgr_0.V_TOP.t2 bgr_0.START_UP.t7 bgr_0.Vin-.t5 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X536 two_stage_opamp_dummy_magic_21_0.VD2.t13 VIN+.t6 two_stage_opamp_dummy_magic_21_0.V_source.t31 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X537 VOUT-.t111 two_stage_opamp_dummy_magic_21_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VOUT+.t114 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VOUT+.t115 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VDDA.t154 bgr_0.1st_Vout_2.t27 bgr_0.PFET_GATE_10uA.t6 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X541 bgr_0.V_mir1.t9 bgr_0.V_mir1.t8 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X542 VOUT-.t112 two_stage_opamp_dummy_magic_21_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VOUT-.t113 two_stage_opamp_dummy_magic_21_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 GNDA.t227 GNDA.t228 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X545 bgr_0.START_UP.t5 bgr_0.START_UP.t4 bgr_0.START_UP_NFET1.t0 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X546 GNDA.t253 GNDA.t251 two_stage_opamp_dummy_magic_21_0.Vb1.t2 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X547 bgr_0.V_p_2.t7 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t14 bgr_0.V_mir2.t15 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X548 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_21_0.X.t44 GNDA.t146 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X549 two_stage_opamp_dummy_magic_21_0.cap_res_X.t138 two_stage_opamp_dummy_magic_21_0.X.t18 GNDA.t181 sky130_fd_pr__res_high_po_1p41 l=1.41
X550 VOUT+.t116 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VOUT-.t114 two_stage_opamp_dummy_magic_21_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 two_stage_opamp_dummy_magic_21_0.V_err_p.t13 two_stage_opamp_dummy_magic_21_0.V_tot.t10 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t2 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X553 VOUT+.t117 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 VOUT+.t118 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VOUT-.t115 two_stage_opamp_dummy_magic_21_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 two_stage_opamp_dummy_magic_21_0.VD3.t13 two_stage_opamp_dummy_magic_21_0.Vb2.t22 two_stage_opamp_dummy_magic_21_0.X.t12 two_stage_opamp_dummy_magic_21_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X558 two_stage_opamp_dummy_magic_21_0.X.t16 two_stage_opamp_dummy_magic_21_0.Vb1.t27 two_stage_opamp_dummy_magic_21_0.VD1.t14 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X559 VOUT+.t119 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VDDA.t216 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t7 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X561 VDDA.t351 VDDA.t349 VOUT-.t15 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X562 VDDA.t111 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t5 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X563 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t25 VDDA.t214 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X564 VOUT-.t116 two_stage_opamp_dummy_magic_21_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VOUT-.t117 two_stage_opamp_dummy_magic_21_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 bgr_0.V_p_1.t0 bgr_0.Vin-.t12 bgr_0.V_mir1.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X567 a_8570_6900.t7 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_21_0.V_err_gate.t8 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X568 GNDA.t227 GNDA.t239 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X569 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t10 VDDA.t346 VDDA.t348 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X570 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 VDDA.t449 two_stage_opamp_dummy_magic_21_0.V_err_gate.t25 a_8570_6900.t13 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X572 VOUT-.t118 two_stage_opamp_dummy_magic_21_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VOUT-.t119 two_stage_opamp_dummy_magic_21_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 GNDA.t70 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_21_0.V_source.t12 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X575 VOUT+.t120 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 GNDA.t72 VDDA.t343 VDDA.t345 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X577 two_stage_opamp_dummy_magic_21_0.Y.t22 two_stage_opamp_dummy_magic_21_0.Vb1.t28 two_stage_opamp_dummy_magic_21_0.VD2.t20 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X578 VDDA.t286 two_stage_opamp_dummy_magic_21_0.Vb3.t22 two_stage_opamp_dummy_magic_21_0.VD4.t27 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X579 VOUT-.t120 two_stage_opamp_dummy_magic_21_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 VOUT+.t121 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 GNDA.t230 GNDA.t229 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X583 VOUT+.t122 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 a_6810_23838.t0 a_6930_22564.t0 GNDA.t113 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X585 VOUT-.t121 two_stage_opamp_dummy_magic_21_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 VOUT+.t123 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 GNDA.t227 GNDA.t231 bgr_0.Vin-.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X588 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_21_0.Vb3.t0 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X589 two_stage_opamp_dummy_magic_21_0.V_err_p.t2 two_stage_opamp_dummy_magic_21_0.V_err_gate.t26 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X590 VOUT+.t124 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 two_stage_opamp_dummy_magic_21_0.V_source.t11 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t28 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X593 two_stage_opamp_dummy_magic_21_0.VD3.t11 two_stage_opamp_dummy_magic_21_0.Vb2.t23 two_stage_opamp_dummy_magic_21_0.X.t8 two_stage_opamp_dummy_magic_21_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X594 VOUT+.t5 two_stage_opamp_dummy_magic_21_0.Y.t49 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X595 two_stage_opamp_dummy_magic_21_0.VD3.t29 two_stage_opamp_dummy_magic_21_0.Vb3.t23 VDDA.t284 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X596 VOUT+.t125 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 GNDA.t186 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_21_0.V_err_gate.t10 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X598 bgr_0.Vin-.t1 bgr_0.V_TOP.t39 VDDA.t147 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X599 two_stage_opamp_dummy_magic_21_0.Y.t14 two_stage_opamp_dummy_magic_21_0.Vb2.t24 two_stage_opamp_dummy_magic_21_0.VD4.t11 two_stage_opamp_dummy_magic_21_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X600 a_12530_23988.t0 a_12410_22380.t1 GNDA.t82 sky130_fd_pr__res_xhigh_po_0p35 l=6
X601 two_stage_opamp_dummy_magic_21_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t19 GNDA.t194 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X602 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 two_stage_opamp_dummy_magic_21_0.V_source.t10 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t29 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X604 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_21_0.X.t45 VDDA.t20 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X605 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_21_0.Y.t50 GNDA.t108 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X606 two_stage_opamp_dummy_magic_21_0.VD2.t1 VIN+.t7 two_stage_opamp_dummy_magic_21_0.V_source.t2 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X607 VOUT-.t122 two_stage_opamp_dummy_magic_21_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 VDDA.t203 bgr_0.V_mir2.t2 bgr_0.V_mir2.t3 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X609 VDDA.t342 VDDA.t340 two_stage_opamp_dummy_magic_21_0.VD4.t36 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X610 VOUT+.t126 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 bgr_0.V_p_1.t5 VDDA.t470 GNDA.t168 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X614 VOUT-.t123 two_stage_opamp_dummy_magic_21_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 two_stage_opamp_dummy_magic_21_0.VD3.t9 two_stage_opamp_dummy_magic_21_0.Vb2.t25 two_stage_opamp_dummy_magic_21_0.X.t10 two_stage_opamp_dummy_magic_21_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X616 a_9370_2200.t2 two_stage_opamp_dummy_magic_21_0.Vb1.t12 two_stage_opamp_dummy_magic_21_0.Vb1.t13 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X617 VDDA.t339 VDDA.t337 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t15 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X618 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_21_0.X.t46 GNDA.t145 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X619 VOUT+.t127 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t1 bgr_0.PFET_GATE_10uA.t26 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X621 two_stage_opamp_dummy_magic_21_0.VD3.t36 VDDA.t334 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X622 VOUT-.t124 two_stage_opamp_dummy_magic_21_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 VOUT-.t125 two_stage_opamp_dummy_magic_21_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_21_0.X.t47 GNDA.t3 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X625 a_13180_23838.t1 a_13060_22630.t1 GNDA.t333 sky130_fd_pr__res_xhigh_po_0p35 l=4
X626 VOUT+.t128 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 bgr_0.V_p_1.t7 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t9 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X628 VDDA.t262 bgr_0.V_mir1.t22 bgr_0.1st_Vout_1.t0 VDDA.t261 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X629 bgr_0.V_TOP.t40 VDDA.t148 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 a_8570_6900.t6 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_21_0.V_err_gate.t5 VDDA.t441 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X631 VDDA.t196 two_stage_opamp_dummy_magic_21_0.X.t48 VOUT-.t5 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X632 VOUT-.t126 two_stage_opamp_dummy_magic_21_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 a_8570_6900.t1 two_stage_opamp_dummy_magic_21_0.V_tot.t11 two_stage_opamp_dummy_magic_21_0.V_err_gate.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X634 VOUT-.t127 two_stage_opamp_dummy_magic_21_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VOUT-.t128 two_stage_opamp_dummy_magic_21_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 VOUT+.t129 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 GNDA.t118 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_21_0.V_p_mir.t1 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X638 VDDA.t194 two_stage_opamp_dummy_magic_21_0.V_err_gate.t27 two_stage_opamp_dummy_magic_21_0.V_err_p.t14 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X639 VOUT-.t129 two_stage_opamp_dummy_magic_21_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 two_stage_opamp_dummy_magic_21_0.Y.t23 two_stage_opamp_dummy_magic_21_0.Vb1.t29 two_stage_opamp_dummy_magic_21_0.VD2.t21 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X641 two_stage_opamp_dummy_magic_21_0.VD3.t7 two_stage_opamp_dummy_magic_21_0.Vb2.t26 two_stage_opamp_dummy_magic_21_0.X.t5 two_stage_opamp_dummy_magic_21_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X642 GNDA.t250 GNDA.t248 VOUT+.t16 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X643 VOUT+.t130 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 VOUT+.t131 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 two_stage_opamp_dummy_magic_21_0.VD3.t28 two_stage_opamp_dummy_magic_21_0.Vb3.t24 VDDA.t282 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X646 bgr_0.V_TOP.t41 VDDA.t149 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 bgr_0.V_p_1.t6 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t10 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X648 VDDA.t333 VDDA.t331 bgr_0.V_TOP.t10 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X649 VOUT-.t130 two_stage_opamp_dummy_magic_21_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 two_stage_opamp_dummy_magic_21_0.Vb2.t2 bgr_0.NFET_GATE_10uA.t20 GNDA.t192 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X651 GNDA.t190 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t10 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X652 VOUT-.t131 two_stage_opamp_dummy_magic_21_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 a_8570_6900.t12 two_stage_opamp_dummy_magic_21_0.V_err_gate.t28 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X654 two_stage_opamp_dummy_magic_21_0.V_source.t9 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t31 GNDA.t119 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X655 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t12 bgr_0.NFET_GATE_10uA.t22 GNDA.t188 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X656 bgr_0.V_TOP.t42 VDDA.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 two_stage_opamp_dummy_magic_21_0.VD1.t3 VIN-.t8 two_stage_opamp_dummy_magic_21_0.V_source.t7 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X658 GNDA.t247 GNDA.t246 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t9 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X659 two_stage_opamp_dummy_magic_21_0.Vb3.t1 two_stage_opamp_dummy_magic_21_0.Vb2.t27 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X660 a_5310_5068.t1 two_stage_opamp_dummy_magic_21_0.V_tot.t3 GNDA.t164 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X661 bgr_0.V_TOP.t43 VDDA.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 VOUT-.t132 two_stage_opamp_dummy_magic_21_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 VOUT-.t133 two_stage_opamp_dummy_magic_21_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 VDDA.t171 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t7 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X665 VOUT-.t134 two_stage_opamp_dummy_magic_21_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 VDDA.t250 bgr_0.1st_Vout_1.t32 bgr_0.V_TOP.t3 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X667 VOUT+.t132 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 VOUT-.t135 two_stage_opamp_dummy_magic_21_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 VOUT-.t136 two_stage_opamp_dummy_magic_21_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 two_stage_opamp_dummy_magic_21_0.VD2.t2 VIN+.t8 two_stage_opamp_dummy_magic_21_0.V_source.t3 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X671 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_21_0.X.t49 VDDA.t443 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X672 VOUT+.t133 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_21_0.Y.t51 GNDA.t109 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X674 VDDA.t330 VDDA.t328 GNDA.t71 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X675 bgr_0.V_TOP.t44 VDDA.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 a_9370_2200.t1 two_stage_opamp_dummy_magic_21_0.Vb1.t8 two_stage_opamp_dummy_magic_21_0.Vb1.t9 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X677 two_stage_opamp_dummy_magic_21_0.X.t9 two_stage_opamp_dummy_magic_21_0.Vb2.t28 two_stage_opamp_dummy_magic_21_0.VD3.t5 two_stage_opamp_dummy_magic_21_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X678 VOUT-.t7 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t7 GNDA.t103 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X679 two_stage_opamp_dummy_magic_21_0.V_err_p.t7 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t17 two_stage_opamp_dummy_magic_21_0.err_amp_out.t0 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X680 bgr_0.V_TOP.t45 VDDA.t187 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 bgr_0.V_mir2.t1 bgr_0.V_mir2.t0 VDDA.t161 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X682 VDDA.t96 bgr_0.V_mir1.t6 bgr_0.V_mir1.t7 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X683 VOUT-.t137 two_stage_opamp_dummy_magic_21_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 two_stage_opamp_dummy_magic_21_0.VD4.t9 two_stage_opamp_dummy_magic_21_0.Vb2.t29 two_stage_opamp_dummy_magic_21_0.Y.t8 two_stage_opamp_dummy_magic_21_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X685 VOUT-.t138 two_stage_opamp_dummy_magic_21_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 two_stage_opamp_dummy_magic_21_0.X.t15 two_stage_opamp_dummy_magic_21_0.Vb1.t30 two_stage_opamp_dummy_magic_21_0.VD1.t13 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X687 VDDA.t280 two_stage_opamp_dummy_magic_21_0.Vb3.t25 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t9 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X688 VDDA.t316 GNDA.t243 GNDA.t245 GNDA.t244 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X689 VOUT-.t139 two_stage_opamp_dummy_magic_21_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 bgr_0.V_mir2.t14 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t18 bgr_0.V_p_2.t9 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X691 VOUT+.t134 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 VDDA.t73 two_stage_opamp_dummy_magic_21_0.X.t50 VOUT-.t1 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X693 a_8570_6900.t0 two_stage_opamp_dummy_magic_21_0.V_tot.t12 two_stage_opamp_dummy_magic_21_0.V_err_gate.t3 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X694 VOUT+.t135 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 bgr_0.PFET_GATE_10uA.t1 VDDA.t471 GNDA.t169 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X696 VOUT+.t136 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 two_stage_opamp_dummy_magic_21_0.VD4.t26 two_stage_opamp_dummy_magic_21_0.Vb3.t26 VDDA.t278 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X698 GNDA.t89 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_21_0.err_amp_out.t4 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X699 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X700 VDDA.t4 two_stage_opamp_dummy_magic_21_0.V_err_gate.t29 a_8570_6900.t11 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X701 two_stage_opamp_dummy_magic_21_0.Y.t5 two_stage_opamp_dummy_magic_21_0.Vb1.t31 two_stage_opamp_dummy_magic_21_0.VD2.t8 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X702 VOUT-.t140 two_stage_opamp_dummy_magic_21_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 VOUT-.t6 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t8 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X704 two_stage_opamp_dummy_magic_21_0.Vb1.t0 bgr_0.PFET_GATE_10uA.t27 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X705 VDDA.t189 bgr_0.V_TOP.t46 bgr_0.Vin-.t0 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X706 VOUT+.t137 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t33 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X708 VOUT+.t138 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VDDA.t165 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t0 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X710 VOUT+.t15 GNDA.t240 GNDA.t242 GNDA.t241 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X711 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t14 VDDA.t325 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X712 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t5 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t4 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X713 VOUT-.t141 two_stage_opamp_dummy_magic_21_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 two_stage_opamp_dummy_magic_21_0.V_err_p.t12 two_stage_opamp_dummy_magic_21_0.V_err_gate.t30 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X715 two_stage_opamp_dummy_magic_21_0.VD4.t7 two_stage_opamp_dummy_magic_21_0.Vb2.t30 two_stage_opamp_dummy_magic_21_0.Y.t9 two_stage_opamp_dummy_magic_21_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X716 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_21_0.Y.t52 VDDA.t43 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X717 two_stage_opamp_dummy_magic_21_0.V_p_mir.t0 VIN+.t9 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t0 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X718 two_stage_opamp_dummy_magic_21_0.VD1.t6 VIN-.t9 two_stage_opamp_dummy_magic_21_0.V_source.t33 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X719 VOUT-.t142 two_stage_opamp_dummy_magic_21_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT+.t139 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VDDA.t68 bgr_0.1st_Vout_2.t34 bgr_0.PFET_GATE_10uA.t4 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X722 VOUT+.t140 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 VOUT+.t141 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VOUT+.t142 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VOUT+.t143 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 a_5190_5068.t0 two_stage_opamp_dummy_magic_21_0.V_tot.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X728 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 two_stage_opamp_dummy_magic_21_0.V_err_p.t4 two_stage_opamp_dummy_magic_21_0.V_err_gate.t31 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X730 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_21_0.X.t51 VDDA.t191 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X731 VOUT-.t143 two_stage_opamp_dummy_magic_21_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 bgr_0.V_mir2.t13 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t19 bgr_0.V_p_2.t8 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X733 two_stage_opamp_dummy_magic_21_0.VD2.t12 VIN+.t10 two_stage_opamp_dummy_magic_21_0.V_source.t30 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X734 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_21_0.X.t52 VDDA.t468 GNDA.t340 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X735 two_stage_opamp_dummy_magic_21_0.X.t6 two_stage_opamp_dummy_magic_21_0.Vb2.t31 two_stage_opamp_dummy_magic_21_0.VD3.t3 two_stage_opamp_dummy_magic_21_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X736 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_21_0.Y.t53 GNDA.t42 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X737 VOUT+.t10 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t9 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X738 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t11 bgr_0.NFET_GATE_10uA.t23 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X739 VOUT-.t144 two_stage_opamp_dummy_magic_21_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 GNDA.t227 GNDA.t226 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X741 VDDA.t276 two_stage_opamp_dummy_magic_21_0.Vb3.t27 two_stage_opamp_dummy_magic_21_0.VD3.t27 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X742 VOUT-.t145 two_stage_opamp_dummy_magic_21_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 VOUT+.t144 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VOUT-.t146 two_stage_opamp_dummy_magic_21_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 VDDA.t266 bgr_0.1st_Vout_1.t36 bgr_0.V_TOP.t8 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X747 GNDA.t170 VDDA.t472 bgr_0.V_TOP.t9 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X748 bgr_0.V_TOP.t47 VDDA.t190 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 GNDA.t238 GNDA.t236 two_stage_opamp_dummy_magic_21_0.V_source.t35 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X750 two_stage_opamp_dummy_magic_21_0.V_err_p.t6 two_stage_opamp_dummy_magic_21_0.V_tot.t13 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t1 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X751 VOUT-.t147 two_stage_opamp_dummy_magic_21_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VDDA.t223 bgr_0.V_TOP.t48 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t0 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X753 VOUT+.t145 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VOUT+.t146 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VOUT+.t147 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 VOUT-.t148 two_stage_opamp_dummy_magic_21_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 VOUT-.t149 two_stage_opamp_dummy_magic_21_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 two_stage_opamp_dummy_magic_21_0.X.t21 two_stage_opamp_dummy_magic_21_0.Vb1.t32 two_stage_opamp_dummy_magic_21_0.VD1.t12 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X759 bgr_0.V_mir2.t12 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t20 bgr_0.V_p_2.t6 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X760 VOUT+.t148 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 two_stage_opamp_dummy_magic_21_0.V_source.t4 two_stage_opamp_dummy_magic_21_0.Vb1.t33 a_9370_2200.t0 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X762 VDDA.t152 bgr_0.PFET_GATE_10uA.t29 bgr_0.V_CUR_REF_REG.t0 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X763 two_stage_opamp_dummy_magic_21_0.Y.t13 two_stage_opamp_dummy_magic_21_0.VD4.t0 two_stage_opamp_dummy_magic_21_0.VD4.t2 two_stage_opamp_dummy_magic_21_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X764 VDDA.t226 two_stage_opamp_dummy_magic_21_0.X.t53 VOUT-.t12 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X765 VOUT+.t149 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 VOUT-.t150 two_stage_opamp_dummy_magic_21_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 a_8570_6900.t5 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_21_0.V_err_gate.t6 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X768 VOUT+.t150 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 two_stage_opamp_dummy_magic_21_0.X.t7 two_stage_opamp_dummy_magic_21_0.Vb2.t32 two_stage_opamp_dummy_magic_21_0.VD3.t1 two_stage_opamp_dummy_magic_21_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X770 VOUT-.t151 two_stage_opamp_dummy_magic_21_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 VDDA.t237 two_stage_opamp_dummy_magic_21_0.V_err_gate.t32 two_stage_opamp_dummy_magic_21_0.V_err_p.t17 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X772 two_stage_opamp_dummy_magic_21_0.Y.t10 two_stage_opamp_dummy_magic_21_0.Vb1.t34 two_stage_opamp_dummy_magic_21_0.VD2.t10 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X773 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t1 a_5710_2046.t0 GNDA.t87 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X774 VDDA.t274 two_stage_opamp_dummy_magic_21_0.Vb3.t28 two_stage_opamp_dummy_magic_21_0.VD3.t26 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X775 VOUT+.t151 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 VOUT-.t152 two_stage_opamp_dummy_magic_21_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 VOUT-.t10 a_14240_2056.t1 GNDA.t153 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X778 VOUT-.t153 two_stage_opamp_dummy_magic_21_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 GNDA.t328 two_stage_opamp_dummy_magic_21_0.X.t54 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t4 VDDA.t454 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X780 VOUT+.t152 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 bgr_0.V_TOP.t49 VDDA.t224 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t4 VDDA.t322 VDDA.t324 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X783 VOUT+.t153 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 two_stage_opamp_dummy_magic_21_0.err_amp_out.t3 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t21 GNDA.t91 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X785 VOUT+.t154 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 VOUT-.t154 two_stage_opamp_dummy_magic_21_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 VOUT-.t155 two_stage_opamp_dummy_magic_21_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X788 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X789 a_5310_5068.t0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t0 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X790 VDDA.t156 bgr_0.V_mir1.t4 bgr_0.V_mir1.t5 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X791 a_8570_6900.t10 two_stage_opamp_dummy_magic_21_0.V_err_gate.t33 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X792 VOUT+.t155 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 VOUT+.t17 VDDA.t319 VDDA.t321 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X794 two_stage_opamp_dummy_magic_21_0.VD1.t8 GNDA.t233 GNDA.t235 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X795 VOUT+.t156 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_21_0.Y.t54 VDDA.t2 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X797 GNDA.t225 GNDA.t223 VDDA.t315 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X798 two_stage_opamp_dummy_magic_21_0.VD1.t5 VIN-.t10 two_stage_opamp_dummy_magic_21_0.V_source.t32 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X799 VOUT-.t156 two_stage_opamp_dummy_magic_21_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t2 384.967
R1 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t10 369.534
R2 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t22 369.534
R3 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t7 369.534
R4 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t16 369.534
R5 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t12 369.534
R6 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.n18 369.534
R7 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 366.553
R8 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t9 192.8
R9 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t17 192.8
R10 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t23 192.8
R11 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t11 192.8
R12 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t20 192.8
R13 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t21 192.8
R14 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t8 192.8
R15 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t15 192.8
R16 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t19 192.8
R17 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t5 192.8
R18 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 192.8
R19 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t18 192.8
R20 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t6 192.8
R21 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t14 192.8
R22 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R23 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R24 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R25 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R26 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R27 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R28 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R29 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R30 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R31 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R32 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R33 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R34 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t0 39.4005
R41 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 39.4005
R42 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t1 24.0005
R44 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t3 24.0005
R45 two_stage_opamp_dummy_magic_21_0.Vb3.n25 two_stage_opamp_dummy_magic_21_0.Vb3.t25 768.551
R46 two_stage_opamp_dummy_magic_21_0.Vb3.n19 two_stage_opamp_dummy_magic_21_0.Vb3.t19 611.739
R47 two_stage_opamp_dummy_magic_21_0.Vb3.n15 two_stage_opamp_dummy_magic_21_0.Vb3.t13 611.739
R48 two_stage_opamp_dummy_magic_21_0.Vb3.n10 two_stage_opamp_dummy_magic_21_0.Vb3.t10 611.739
R49 two_stage_opamp_dummy_magic_21_0.Vb3.n6 two_stage_opamp_dummy_magic_21_0.Vb3.t27 611.739
R50 two_stage_opamp_dummy_magic_21_0.Vb3.n24 two_stage_opamp_dummy_magic_21_0.Vb3.n23 428.976
R51 two_stage_opamp_dummy_magic_21_0.Vb3.n24 two_stage_opamp_dummy_magic_21_0.Vb3.n14 428.445
R52 two_stage_opamp_dummy_magic_21_0.Vb3.n19 two_stage_opamp_dummy_magic_21_0.Vb3.t15 421.75
R53 two_stage_opamp_dummy_magic_21_0.Vb3.n20 two_stage_opamp_dummy_magic_21_0.Vb3.t17 421.75
R54 two_stage_opamp_dummy_magic_21_0.Vb3.n21 two_stage_opamp_dummy_magic_21_0.Vb3.t14 421.75
R55 two_stage_opamp_dummy_magic_21_0.Vb3.n22 two_stage_opamp_dummy_magic_21_0.Vb3.t26 421.75
R56 two_stage_opamp_dummy_magic_21_0.Vb3.n15 two_stage_opamp_dummy_magic_21_0.Vb3.t16 421.75
R57 two_stage_opamp_dummy_magic_21_0.Vb3.n16 two_stage_opamp_dummy_magic_21_0.Vb3.t21 421.75
R58 two_stage_opamp_dummy_magic_21_0.Vb3.n17 two_stage_opamp_dummy_magic_21_0.Vb3.t18 421.75
R59 two_stage_opamp_dummy_magic_21_0.Vb3.n18 two_stage_opamp_dummy_magic_21_0.Vb3.t22 421.75
R60 two_stage_opamp_dummy_magic_21_0.Vb3.n10 two_stage_opamp_dummy_magic_21_0.Vb3.t12 421.75
R61 two_stage_opamp_dummy_magic_21_0.Vb3.n11 two_stage_opamp_dummy_magic_21_0.Vb3.t9 421.75
R62 two_stage_opamp_dummy_magic_21_0.Vb3.n12 two_stage_opamp_dummy_magic_21_0.Vb3.t28 421.75
R63 two_stage_opamp_dummy_magic_21_0.Vb3.n13 two_stage_opamp_dummy_magic_21_0.Vb3.t24 421.75
R64 two_stage_opamp_dummy_magic_21_0.Vb3.n6 two_stage_opamp_dummy_magic_21_0.Vb3.t8 421.75
R65 two_stage_opamp_dummy_magic_21_0.Vb3.n7 two_stage_opamp_dummy_magic_21_0.Vb3.t11 421.75
R66 two_stage_opamp_dummy_magic_21_0.Vb3.n8 two_stage_opamp_dummy_magic_21_0.Vb3.t23 421.75
R67 two_stage_opamp_dummy_magic_21_0.Vb3.n9 two_stage_opamp_dummy_magic_21_0.Vb3.t20 421.75
R68 two_stage_opamp_dummy_magic_21_0.Vb3.n20 two_stage_opamp_dummy_magic_21_0.Vb3.n19 167.094
R69 two_stage_opamp_dummy_magic_21_0.Vb3.n21 two_stage_opamp_dummy_magic_21_0.Vb3.n20 167.094
R70 two_stage_opamp_dummy_magic_21_0.Vb3.n22 two_stage_opamp_dummy_magic_21_0.Vb3.n21 167.094
R71 two_stage_opamp_dummy_magic_21_0.Vb3.n16 two_stage_opamp_dummy_magic_21_0.Vb3.n15 167.094
R72 two_stage_opamp_dummy_magic_21_0.Vb3.n17 two_stage_opamp_dummy_magic_21_0.Vb3.n16 167.094
R73 two_stage_opamp_dummy_magic_21_0.Vb3.n18 two_stage_opamp_dummy_magic_21_0.Vb3.n17 167.094
R74 two_stage_opamp_dummy_magic_21_0.Vb3.n11 two_stage_opamp_dummy_magic_21_0.Vb3.n10 167.094
R75 two_stage_opamp_dummy_magic_21_0.Vb3.n12 two_stage_opamp_dummy_magic_21_0.Vb3.n11 167.094
R76 two_stage_opamp_dummy_magic_21_0.Vb3.n13 two_stage_opamp_dummy_magic_21_0.Vb3.n12 167.094
R77 two_stage_opamp_dummy_magic_21_0.Vb3.n7 two_stage_opamp_dummy_magic_21_0.Vb3.n6 167.094
R78 two_stage_opamp_dummy_magic_21_0.Vb3.n8 two_stage_opamp_dummy_magic_21_0.Vb3.n7 167.094
R79 two_stage_opamp_dummy_magic_21_0.Vb3.n9 two_stage_opamp_dummy_magic_21_0.Vb3.n8 167.094
R80 two_stage_opamp_dummy_magic_21_0.Vb3.n2 two_stage_opamp_dummy_magic_21_0.Vb3.n0 139.639
R81 two_stage_opamp_dummy_magic_21_0.Vb3.n2 two_stage_opamp_dummy_magic_21_0.Vb3.n1 139.638
R82 two_stage_opamp_dummy_magic_21_0.Vb3.n4 two_stage_opamp_dummy_magic_21_0.Vb3.n3 134.577
R83 two_stage_opamp_dummy_magic_21_0.Vb3.n26 two_stage_opamp_dummy_magic_21_0.Vb3.n5 73.3151
R84 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_21_0.Vb3.n26 47.563
R85 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_21_0.Vb3.n4 41.063
R86 two_stage_opamp_dummy_magic_21_0.Vb3.n23 two_stage_opamp_dummy_magic_21_0.Vb3.n22 35.3472
R87 two_stage_opamp_dummy_magic_21_0.Vb3.n23 two_stage_opamp_dummy_magic_21_0.Vb3.n18 35.3472
R88 two_stage_opamp_dummy_magic_21_0.Vb3.n14 two_stage_opamp_dummy_magic_21_0.Vb3.n13 35.3472
R89 two_stage_opamp_dummy_magic_21_0.Vb3.n14 two_stage_opamp_dummy_magic_21_0.Vb3.n9 35.3472
R90 two_stage_opamp_dummy_magic_21_0.Vb3.n3 two_stage_opamp_dummy_magic_21_0.Vb3.t4 24.0005
R91 two_stage_opamp_dummy_magic_21_0.Vb3.n3 two_stage_opamp_dummy_magic_21_0.Vb3.t6 24.0005
R92 two_stage_opamp_dummy_magic_21_0.Vb3.n1 two_stage_opamp_dummy_magic_21_0.Vb3.t7 24.0005
R93 two_stage_opamp_dummy_magic_21_0.Vb3.n1 two_stage_opamp_dummy_magic_21_0.Vb3.t2 24.0005
R94 two_stage_opamp_dummy_magic_21_0.Vb3.n0 two_stage_opamp_dummy_magic_21_0.Vb3.t5 24.0005
R95 two_stage_opamp_dummy_magic_21_0.Vb3.n0 two_stage_opamp_dummy_magic_21_0.Vb3.t3 24.0005
R96 two_stage_opamp_dummy_magic_21_0.Vb3.n25 two_stage_opamp_dummy_magic_21_0.Vb3.n24 14.3443
R97 two_stage_opamp_dummy_magic_21_0.Vb3.n5 two_stage_opamp_dummy_magic_21_0.Vb3.t0 11.2576
R98 two_stage_opamp_dummy_magic_21_0.Vb3.n5 two_stage_opamp_dummy_magic_21_0.Vb3.t1 11.2576
R99 two_stage_opamp_dummy_magic_21_0.Vb3.n4 two_stage_opamp_dummy_magic_21_0.Vb3.n2 4.5005
R100 two_stage_opamp_dummy_magic_21_0.Vb3.n26 two_stage_opamp_dummy_magic_21_0.Vb3.n25 1.21925
R101 GNDA.n2244 GNDA.n33 197450
R102 GNDA.n281 GNDA.n33 146899
R103 GNDA.n2244 GNDA.n34 127050
R104 GNDA.n266 GNDA.n148 14938
R105 GNDA.n2245 GNDA.n32 14922.8
R106 GNDA.n267 GNDA.n147 13700
R107 GNDA.n147 GNDA.n146 13700
R108 GNDA.n275 GNDA.n140 13200
R109 GNDA.n273 GNDA.n137 13132.3
R110 GNDA.n401 GNDA.n400 11953.3
R111 GNDA.n400 GNDA.n281 11890.5
R112 GNDA.n144 GNDA.n143 11440
R113 GNDA.n138 GNDA.n31 11404.3
R114 GNDA.n270 GNDA.n269 11377.2
R115 GNDA.n281 GNDA.n280 9950.42
R116 GNDA.n401 GNDA.n136 9950.42
R117 GNDA.n269 GNDA.n142 9371.43
R118 GNDA.n2245 GNDA.n31 9371.43
R119 GNDA.n139 GNDA.n138 9265.27
R120 GNDA.n138 GNDA.n34 8497.25
R121 GNDA.n271 GNDA.n270 8420
R122 GNDA.n268 GNDA.n144 7648.94
R123 GNDA.n145 GNDA.n144 7630.38
R124 GNDA.n143 GNDA.n140 7385.71
R125 GNDA.n279 GNDA.n278 6922.94
R126 GNDA.n272 GNDA.n141 6860
R127 GNDA.n273 GNDA.n136 6858.08
R128 GNDA.n280 GNDA.n137 6858.08
R129 GNDA.n270 GNDA.n140 6364.29
R130 GNDA.n276 GNDA.n139 5313.76
R131 GNDA.n402 GNDA.n401 4497.78
R132 GNDA.n277 GNDA.n137 4106.67
R133 GNDA.n274 GNDA.n273 4106.67
R134 GNDA.n400 GNDA.n399 3974.19
R135 GNDA.t2 GNDA.n2244 3883.81
R136 GNDA.n146 GNDA.n145 3498
R137 GNDA.n268 GNDA.n267 3463.37
R138 GNDA.n2244 GNDA.t37 3033.02
R139 GNDA.n143 GNDA.n139 2900.98
R140 GNDA.n278 GNDA.n34 2704.59
R141 GNDA.n272 GNDA.n271 2680
R142 GNDA.n271 GNDA.n142 2570.64
R143 GNDA.n146 GNDA.n32 2520.94
R144 GNDA.n267 GNDA.n266 2481.49
R145 GNDA.t127 GNDA.n148 2095.78
R146 GNDA.n271 GNDA.n135 1987.75
R147 GNDA.n276 GNDA.n275 1808.75
R148 GNDA.n196 GNDA.n147 1800
R149 GNDA.n141 GNDA.n135 1460.18
R150 GNDA.n141 GNDA.n136 1460.18
R151 GNDA.n266 GNDA.t303 1441.38
R152 GNDA.n280 GNDA.n279 1440.71
R153 GNDA.n279 GNDA.n33 1440.71
R154 GNDA.n32 GNDA.t313 1426.21
R155 GNDA.t150 GNDA.n402 1360.43
R156 GNDA.n1630 GNDA.n1629 1224.73
R157 GNDA.n965 GNDA.n958 1214.72
R158 GNDA.n996 GNDA.n965 1214.72
R159 GNDA.n996 GNDA.n995 1214.72
R160 GNDA.n995 GNDA.n994 1214.72
R161 GNDA.n994 GNDA.n434 1214.72
R162 GNDA.n987 GNDA.n433 1214.72
R163 GNDA.n987 GNDA.n986 1214.72
R164 GNDA.n986 GNDA.n985 1214.72
R165 GNDA.n985 GNDA.n976 1214.72
R166 GNDA.n976 GNDA.n432 1214.72
R167 GNDA.n1716 GNDA.n1715 1214.72
R168 GNDA.n1715 GNDA.n1714 1214.72
R169 GNDA.n1714 GNDA.n1684 1214.72
R170 GNDA.n1708 GNDA.n1684 1214.72
R171 GNDA.n1708 GNDA.n426 1214.72
R172 GNDA.n1696 GNDA.n425 1214.72
R173 GNDA.n1701 GNDA.n1696 1214.72
R174 GNDA.n1701 GNDA.n1700 1214.72
R175 GNDA.n1700 GNDA.n1699 1214.72
R176 GNDA.n1699 GNDA.n424 1214.72
R177 GNDA.n2153 GNDA.n2152 1185.07
R178 GNDA.n2152 GNDA.n2151 1185.07
R179 GNDA.n260 GNDA.n259 1182.8
R180 GNDA.n245 GNDA.n244 1182.8
R181 GNDA.n2062 GNDA.n36 1109.51
R182 GNDA.n274 GNDA.n272 1000.58
R183 GNDA.n278 GNDA.n277 1000.58
R184 GNDA.n402 GNDA.n135 872.588
R185 GNDA.t227 GNDA.n434 823.313
R186 GNDA.t227 GNDA.n426 823.313
R187 GNDA.n148 GNDA.t181 796.269
R188 GNDA.t181 GNDA.n142 779.851
R189 GNDA.n186 GNDA.t282 749.742
R190 GNDA.n158 GNDA.t260 749.742
R191 GNDA.n2250 GNDA.t223 749.742
R192 GNDA.n2248 GNDA.t243 749.742
R193 GNDA.n2232 GNDA.n2231 686.717
R194 GNDA.n2235 GNDA.n36 686.717
R195 GNDA.n2235 GNDA.n35 686.717
R196 GNDA.n2223 GNDA.n47 686.717
R197 GNDA.n416 GNDA.n405 686.717
R198 GNDA.n949 GNDA.n944 669.307
R199 GNDA.n238 GNDA.t270 659.367
R200 GNDA.n213 GNDA.t236 659.367
R201 GNDA.n277 GNDA.n276 641.399
R202 GNDA.n134 GNDA.n133 585.001
R203 GNDA.n2167 GNDA.n2166 585.001
R204 GNDA.n2179 GNDA.n2178 585.001
R205 GNDA.n2181 GNDA.n2180 585.001
R206 GNDA.n2191 GNDA.n2190 585.001
R207 GNDA.n2242 GNDA.n2241 585.001
R208 GNDA.n1989 GNDA.n1988 585
R209 GNDA.n2067 GNDA.n2066 585
R210 GNDA.n2068 GNDA.n2067 585
R211 GNDA.n1986 GNDA.n1985 585
R212 GNDA.n2069 GNDA.n1986 585
R213 GNDA.n2072 GNDA.n2071 585
R214 GNDA.n2071 GNDA.n2070 585
R215 GNDA.n2073 GNDA.n1984 585
R216 GNDA.n1987 GNDA.n1984 585
R217 GNDA.n2075 GNDA.n2074 585
R218 GNDA.n2075 GNDA.n50 585
R219 GNDA.n2076 GNDA.n1983 585
R220 GNDA.n2076 GNDA.n49 585
R221 GNDA.n2079 GNDA.n2078 585
R222 GNDA.n2078 GNDA.n2077 585
R223 GNDA.n2080 GNDA.n1981 585
R224 GNDA.n1981 GNDA.n1980 585
R225 GNDA.n2082 GNDA.n2081 585
R226 GNDA.n2083 GNDA.n2082 585
R227 GNDA.n1982 GNDA.n125 585
R228 GNDA.n2084 GNDA.n125 585
R229 GNDA.n2086 GNDA.n123 585
R230 GNDA.n2086 GNDA.n2085 585
R231 GNDA.n2063 GNDA.n2062 585
R232 GNDA.n1174 GNDA.n1173 585
R233 GNDA.n1584 GNDA.n1170 585
R234 GNDA.n1170 GNDA.n1169 585
R235 GNDA.n1586 GNDA.n1585 585
R236 GNDA.n1587 GNDA.n1586 585
R237 GNDA.n1171 GNDA.n1168 585
R238 GNDA.n1588 GNDA.n1168 585
R239 GNDA.n1590 GNDA.n1167 585
R240 GNDA.n1590 GNDA.n1589 585
R241 GNDA.n1592 GNDA.n1591 585
R242 GNDA.n1591 GNDA.n428 585
R243 GNDA.n1593 GNDA.n1166 585
R244 GNDA.n1166 GNDA.n429 585
R245 GNDA.n1595 GNDA.n1594 585
R246 GNDA.n1596 GNDA.n1595 585
R247 GNDA.n1165 GNDA.n1164 585
R248 GNDA.n1597 GNDA.n1165 585
R249 GNDA.n1600 GNDA.n1599 585
R250 GNDA.n1599 GNDA.n1598 585
R251 GNDA.n1601 GNDA.n1142 585
R252 GNDA.n1142 GNDA.n1140 585
R253 GNDA.n1603 GNDA.n1602 585
R254 GNDA.n1604 GNDA.n1603 585
R255 GNDA.n1581 GNDA.n427 585
R256 GNDA.n1139 GNDA.n1137 585
R257 GNDA.n1606 GNDA.n1605 585
R258 GNDA.n1609 GNDA.n1021 585
R259 GNDA.n1021 GNDA.n1020 585
R260 GNDA.n1611 GNDA.n1610 585
R261 GNDA.n1612 GNDA.n1611 585
R262 GNDA.n1022 GNDA.n1019 585
R263 GNDA.n1613 GNDA.n1019 585
R264 GNDA.n1615 GNDA.n1018 585
R265 GNDA.n1615 GNDA.n1614 585
R266 GNDA.n1617 GNDA.n1616 585
R267 GNDA.n1616 GNDA.n430 585
R268 GNDA.n1618 GNDA.n1017 585
R269 GNDA.n1017 GNDA.n431 585
R270 GNDA.n1620 GNDA.n1619 585
R271 GNDA.n1621 GNDA.n1620 585
R272 GNDA.n1016 GNDA.n1015 585
R273 GNDA.n1622 GNDA.n1016 585
R274 GNDA.n1625 GNDA.n1624 585
R275 GNDA.n1624 GNDA.n1623 585
R276 GNDA.n1626 GNDA.n1014 585
R277 GNDA.n1014 GNDA.n1013 585
R278 GNDA.n1628 GNDA.n1627 585
R279 GNDA.n1629 GNDA.n1628 585
R280 GNDA.n981 GNDA.n980 585
R281 GNDA.n980 GNDA.n432 585
R282 GNDA.n982 GNDA.n979 585
R283 GNDA.n979 GNDA.n976 585
R284 GNDA.n983 GNDA.n975 585
R285 GNDA.n985 GNDA.n975 585
R286 GNDA.n978 GNDA.n974 585
R287 GNDA.n986 GNDA.n974 585
R288 GNDA.n973 GNDA.n971 585
R289 GNDA.n987 GNDA.n973 585
R290 GNDA.n990 GNDA.n970 585
R291 GNDA.n970 GNDA.n433 585
R292 GNDA.n991 GNDA.n969 585
R293 GNDA.n969 GNDA.n434 585
R294 GNDA.n992 GNDA.n967 585
R295 GNDA.n994 GNDA.n967 585
R296 GNDA.n966 GNDA.n963 585
R297 GNDA.n995 GNDA.n966 585
R298 GNDA.n998 GNDA.n962 585
R299 GNDA.n996 GNDA.n962 585
R300 GNDA.n999 GNDA.n961 585
R301 GNDA.n965 GNDA.n961 585
R302 GNDA.n1000 GNDA.n957 585
R303 GNDA.n958 GNDA.n957 585
R304 GNDA.n1001 GNDA.n1000 585
R305 GNDA.n1001 GNDA.n958 585
R306 GNDA.n999 GNDA.n960 585
R307 GNDA.n965 GNDA.n960 585
R308 GNDA.n998 GNDA.n997 585
R309 GNDA.n997 GNDA.n996 585
R310 GNDA.n964 GNDA.n963 585
R311 GNDA.n995 GNDA.n964 585
R312 GNDA.n993 GNDA.n992 585
R313 GNDA.n994 GNDA.n993 585
R314 GNDA.n991 GNDA.n968 585
R315 GNDA.n968 GNDA.n434 585
R316 GNDA.n990 GNDA.n989 585
R317 GNDA.n989 GNDA.n433 585
R318 GNDA.n988 GNDA.n971 585
R319 GNDA.n988 GNDA.n987 585
R320 GNDA.n978 GNDA.n972 585
R321 GNDA.n986 GNDA.n972 585
R322 GNDA.n984 GNDA.n983 585
R323 GNDA.n985 GNDA.n984 585
R324 GNDA.n982 GNDA.n977 585
R325 GNDA.n977 GNDA.n976 585
R326 GNDA.n981 GNDA.n512 585
R327 GNDA.n512 GNDA.n432 585
R328 GNDA.n1945 GNDA.n1944 585
R329 GNDA.n1942 GNDA.n493 585
R330 GNDA.n1941 GNDA.n494 585
R331 GNDA.n1939 GNDA.n1938 585
R332 GNDA.n496 GNDA.n495 585
R333 GNDA.n504 GNDA.n500 585
R334 GNDA.n1931 GNDA.n1930 585
R335 GNDA.n1928 GNDA.n502 585
R336 GNDA.n1927 GNDA.n505 585
R337 GNDA.n1925 GNDA.n1924 585
R338 GNDA.n507 GNDA.n506 585
R339 GNDA.n1917 GNDA.n1916 585
R340 GNDA.n1918 GNDA.n1917 585
R341 GNDA.n1920 GNDA.n507 585
R342 GNDA.n1924 GNDA.n1923 585
R343 GNDA.n1923 GNDA.n435 585
R344 GNDA.n1922 GNDA.n505 585
R345 GNDA.n502 GNDA.n501 585
R346 GNDA.n1932 GNDA.n1931 585
R347 GNDA.n1934 GNDA.n500 585
R348 GNDA.n1935 GNDA.n496 585
R349 GNDA.n1938 GNDA.n1937 585
R350 GNDA.n499 GNDA.n494 585
R351 GNDA.n497 GNDA.n493 585
R352 GNDA.n1945 GNDA.n489 585
R353 GNDA.n489 GNDA.n435 585
R354 GNDA.n2138 GNDA.n102 585
R355 GNDA.n2141 GNDA.n2140 585
R356 GNDA.n2137 GNDA.n104 585
R357 GNDA.n2135 GNDA.n2134 585
R358 GNDA.n106 GNDA.n105 585
R359 GNDA.n2128 GNDA.n2127 585
R360 GNDA.n2125 GNDA.n108 585
R361 GNDA.n2123 GNDA.n2122 585
R362 GNDA.n110 GNDA.n109 585
R363 GNDA.n2116 GNDA.n2115 585
R364 GNDA.n2113 GNDA.n112 585
R365 GNDA.n2111 GNDA.n2110 585
R366 GNDA.n2110 GNDA.n2109 585
R367 GNDA.n112 GNDA.n111 585
R368 GNDA.n2117 GNDA.n2116 585
R369 GNDA.n2119 GNDA.n110 585
R370 GNDA.n2122 GNDA.n2121 585
R371 GNDA.n108 GNDA.n107 585
R372 GNDA.n2129 GNDA.n2128 585
R373 GNDA.n2131 GNDA.n106 585
R374 GNDA.n2134 GNDA.n2133 585
R375 GNDA.n104 GNDA.n103 585
R376 GNDA.n2142 GNDA.n2141 585
R377 GNDA.n2144 GNDA.n102 585
R378 GNDA.n2163 GNDA.n90 585
R379 GNDA.n2161 GNDA.n2160 585
R380 GNDA.n92 GNDA.n91 585
R381 GNDA.n728 GNDA.n727 585
R382 GNDA.n733 GNDA.n725 585
R383 GNDA.n734 GNDA.n723 585
R384 GNDA.n735 GNDA.n722 585
R385 GNDA.n720 GNDA.n718 585
R386 GNDA.n740 GNDA.n717 585
R387 GNDA.n741 GNDA.n715 585
R388 GNDA.n714 GNDA.n683 585
R389 GNDA.n746 GNDA.n681 585
R390 GNDA.n746 GNDA.n745 585
R391 GNDA.n743 GNDA.n683 585
R392 GNDA.n742 GNDA.n741 585
R393 GNDA.n740 GNDA.n739 585
R394 GNDA.n738 GNDA.n718 585
R395 GNDA.n736 GNDA.n735 585
R396 GNDA.n734 GNDA.n719 585
R397 GNDA.n733 GNDA.n732 585
R398 GNDA.n730 GNDA.n728 585
R399 GNDA.n93 GNDA.n92 585
R400 GNDA.n2160 GNDA.n2159 585
R401 GNDA.n2157 GNDA.n90 585
R402 GNDA.n1952 GNDA.n483 585
R403 GNDA.n1953 GNDA.n474 585
R404 GNDA.n1956 GNDA.n473 585
R405 GNDA.n1957 GNDA.n472 585
R406 GNDA.n1960 GNDA.n471 585
R407 GNDA.n1961 GNDA.n470 585
R408 GNDA.n1964 GNDA.n469 585
R409 GNDA.n1966 GNDA.n468 585
R410 GNDA.n1967 GNDA.n467 585
R411 GNDA.n1968 GNDA.n466 585
R412 GNDA.n475 GNDA.n458 585
R413 GNDA.n1974 GNDA.n454 585
R414 GNDA.n1974 GNDA.n1973 585
R415 GNDA.n460 GNDA.n458 585
R416 GNDA.n1969 GNDA.n1968 585
R417 GNDA.n1967 GNDA.n465 585
R418 GNDA.n1966 GNDA.n1965 585
R419 GNDA.n1964 GNDA.n1963 585
R420 GNDA.n1962 GNDA.n1961 585
R421 GNDA.n1960 GNDA.n1959 585
R422 GNDA.n1958 GNDA.n1957 585
R423 GNDA.n1956 GNDA.n1955 585
R424 GNDA.n1954 GNDA.n1953 585
R425 GNDA.n1952 GNDA.n1951 585
R426 GNDA.n1887 GNDA.n1886 585
R427 GNDA.n1887 GNDA.n424 585
R428 GNDA.n517 GNDA.n516 585
R429 GNDA.n1699 GNDA.n516 585
R430 GNDA.n1697 GNDA.n1694 585
R431 GNDA.n1700 GNDA.n1697 585
R432 GNDA.n1703 GNDA.n1693 585
R433 GNDA.n1701 GNDA.n1693 585
R434 GNDA.n1704 GNDA.n1692 585
R435 GNDA.n1696 GNDA.n1692 585
R436 GNDA.n1705 GNDA.n1691 585
R437 GNDA.n1691 GNDA.n425 585
R438 GNDA.n1690 GNDA.n1688 585
R439 GNDA.n1690 GNDA.n426 585
R440 GNDA.n1710 GNDA.n1687 585
R441 GNDA.n1708 GNDA.n1687 585
R442 GNDA.n1711 GNDA.n1686 585
R443 GNDA.n1686 GNDA.n1684 585
R444 GNDA.n1712 GNDA.n1683 585
R445 GNDA.n1714 GNDA.n1683 585
R446 GNDA.n1682 GNDA.n937 585
R447 GNDA.n1715 GNDA.n1682 585
R448 GNDA.n1718 GNDA.n935 585
R449 GNDA.n1716 GNDA.n935 585
R450 GNDA.n1718 GNDA.n1717 585
R451 GNDA.n1717 GNDA.n1716 585
R452 GNDA.n1681 GNDA.n937 585
R453 GNDA.n1715 GNDA.n1681 585
R454 GNDA.n1713 GNDA.n1712 585
R455 GNDA.n1714 GNDA.n1713 585
R456 GNDA.n1711 GNDA.n1685 585
R457 GNDA.n1685 GNDA.n1684 585
R458 GNDA.n1710 GNDA.n1709 585
R459 GNDA.n1709 GNDA.n1708 585
R460 GNDA.n1707 GNDA.n1688 585
R461 GNDA.n1707 GNDA.n426 585
R462 GNDA.n1706 GNDA.n1705 585
R463 GNDA.n1706 GNDA.n425 585
R464 GNDA.n1704 GNDA.n1689 585
R465 GNDA.n1696 GNDA.n1689 585
R466 GNDA.n1703 GNDA.n1702 585
R467 GNDA.n1702 GNDA.n1701 585
R468 GNDA.n1695 GNDA.n1694 585
R469 GNDA.n1700 GNDA.n1695 585
R470 GNDA.n1698 GNDA.n517 585
R471 GNDA.n1699 GNDA.n1698 585
R472 GNDA.n1886 GNDA.n518 585
R473 GNDA.n518 GNDA.n424 585
R474 GNDA.n1721 GNDA.n1720 585
R475 GNDA.n1722 GNDA.n1721 585
R476 GNDA.n933 GNDA.n932 585
R477 GNDA.n1723 GNDA.n933 585
R478 GNDA.n1726 GNDA.n1725 585
R479 GNDA.n1725 GNDA.n1724 585
R480 GNDA.n1727 GNDA.n931 585
R481 GNDA.n931 GNDA.n930 585
R482 GNDA.n1729 GNDA.n1728 585
R483 GNDA.n1730 GNDA.n1729 585
R484 GNDA.n929 GNDA.n928 585
R485 GNDA.n1731 GNDA.n929 585
R486 GNDA.n1734 GNDA.n1733 585
R487 GNDA.n1733 GNDA.n1732 585
R488 GNDA.n1735 GNDA.n927 585
R489 GNDA.n927 GNDA.n926 585
R490 GNDA.n1737 GNDA.n1736 585
R491 GNDA.n1738 GNDA.n1737 585
R492 GNDA.n925 GNDA.n924 585
R493 GNDA.n1739 GNDA.n925 585
R494 GNDA.n1742 GNDA.n1741 585
R495 GNDA.n1741 GNDA.n1740 585
R496 GNDA.n1743 GNDA.n923 585
R497 GNDA.n923 GNDA.n423 585
R498 GNDA.n1657 GNDA.n1656 585
R499 GNDA.n1656 GNDA.n1655 585
R500 GNDA.n1658 GNDA.n954 585
R501 GNDA.n954 GNDA.n953 585
R502 GNDA.n1660 GNDA.n1659 585
R503 GNDA.n1661 GNDA.n1660 585
R504 GNDA.n955 GNDA.n952 585
R505 GNDA.n1662 GNDA.n952 585
R506 GNDA.n1664 GNDA.n951 585
R507 GNDA.n1664 GNDA.n1663 585
R508 GNDA.n1666 GNDA.n1665 585
R509 GNDA.n1665 GNDA.n945 585
R510 GNDA.n943 GNDA.n942 585
R511 GNDA.n1670 GNDA.n943 585
R512 GNDA.n1673 GNDA.n1672 585
R513 GNDA.n1672 GNDA.n1671 585
R514 GNDA.n1674 GNDA.n940 585
R515 GNDA.n940 GNDA.n939 585
R516 GNDA.n1676 GNDA.n1675 585
R517 GNDA.n1677 GNDA.n1676 585
R518 GNDA.n941 GNDA.n938 585
R519 GNDA.n1678 GNDA.n938 585
R520 GNDA.n1680 GNDA.n936 585
R521 GNDA.n1680 GNDA.n1679 585
R522 GNDA.n1012 GNDA.n1011 585
R523 GNDA.n1630 GNDA.n1012 585
R524 GNDA.n1633 GNDA.n1632 585
R525 GNDA.n1632 GNDA.n1631 585
R526 GNDA.n1634 GNDA.n1010 585
R527 GNDA.n1010 GNDA.n1009 585
R528 GNDA.n1636 GNDA.n1635 585
R529 GNDA.n1637 GNDA.n1636 585
R530 GNDA.n1008 GNDA.n1007 585
R531 GNDA.n1638 GNDA.n1008 585
R532 GNDA.n1641 GNDA.n1640 585
R533 GNDA.n1640 GNDA.n1639 585
R534 GNDA.n1642 GNDA.n1006 585
R535 GNDA.n1006 GNDA.n1005 585
R536 GNDA.n1644 GNDA.n1643 585
R537 GNDA.n1645 GNDA.n1644 585
R538 GNDA.n1004 GNDA.n1003 585
R539 GNDA.n1646 GNDA.n1004 585
R540 GNDA.n1649 GNDA.n1648 585
R541 GNDA.n1648 GNDA.n1647 585
R542 GNDA.n1650 GNDA.n1002 585
R543 GNDA.n1002 GNDA.n959 585
R544 GNDA.n1652 GNDA.n1651 585
R545 GNDA.n1653 GNDA.n1652 585
R546 GNDA.n950 GNDA.n946 585
R547 GNDA.n1669 GNDA.n1668 585
R548 GNDA.t227 GNDA.n1669 585
R549 GNDA.n1977 GNDA.n1976 585
R550 GNDA.n455 GNDA.n453 585
R551 GNDA.n1302 GNDA.n1301 585
R552 GNDA.n1304 GNDA.n1303 585
R553 GNDA.n1306 GNDA.n1305 585
R554 GNDA.n1308 GNDA.n1307 585
R555 GNDA.n1310 GNDA.n1309 585
R556 GNDA.n1312 GNDA.n1311 585
R557 GNDA.n1314 GNDA.n1313 585
R558 GNDA.n1316 GNDA.n1315 585
R559 GNDA.n1318 GNDA.n1317 585
R560 GNDA.n1320 GNDA.n1319 585
R561 GNDA.n1914 GNDA.n1913 585
R562 GNDA.n1912 GNDA.n1911 585
R563 GNDA.n1910 GNDA.n1909 585
R564 GNDA.n1908 GNDA.n1907 585
R565 GNDA.n1906 GNDA.n1905 585
R566 GNDA.n1904 GNDA.n1903 585
R567 GNDA.n1902 GNDA.n1901 585
R568 GNDA.n1900 GNDA.n1899 585
R569 GNDA.n1898 GNDA.n1897 585
R570 GNDA.n1896 GNDA.n1895 585
R571 GNDA.n1894 GNDA.n1893 585
R572 GNDA.n459 GNDA.n456 585
R573 GNDA.n1163 GNDA.n1141 585
R574 GNDA.n1162 GNDA.n1161 585
R575 GNDA.n1160 GNDA.n1159 585
R576 GNDA.n1158 GNDA.n1157 585
R577 GNDA.n1156 GNDA.n1155 585
R578 GNDA.n1154 GNDA.n1153 585
R579 GNDA.n1152 GNDA.n1151 585
R580 GNDA.n1150 GNDA.n1149 585
R581 GNDA.n1148 GNDA.n1147 585
R582 GNDA.n1146 GNDA.n1145 585
R583 GNDA.n1144 GNDA.n1143 585
R584 GNDA.n509 GNDA.n508 585
R585 GNDA.n1888 GNDA.n457 585
R586 GNDA.n1889 GNDA.n1888 585
R587 GNDA.n1879 GNDA.n1878 585
R588 GNDA.n1876 GNDA.n650 585
R589 GNDA.n1769 GNDA.n1768 585
R590 GNDA.n1871 GNDA.n1870 585
R591 GNDA.n1869 GNDA.n1868 585
R592 GNDA.n1795 GNDA.n1773 585
R593 GNDA.n1797 GNDA.n1796 585
R594 GNDA.n1802 GNDA.n1801 585
R595 GNDA.n1800 GNDA.n1793 585
R596 GNDA.n1808 GNDA.n1807 585
R597 GNDA.n1810 GNDA.n1809 585
R598 GNDA.n519 GNDA.n515 585
R599 GNDA.n1891 GNDA.n511 585
R600 GNDA.n1889 GNDA.n511 585
R601 GNDA.n514 GNDA.n457 585
R602 GNDA.n1889 GNDA.n514 585
R603 GNDA.n1884 GNDA.n1883 585
R604 GNDA.n533 GNDA.n521 585
R605 GNDA.n643 GNDA.n642 585
R606 GNDA.n535 GNDA.n532 585
R607 GNDA.n561 GNDA.n560 585
R608 GNDA.n565 GNDA.n564 585
R609 GNDA.n567 GNDA.n566 585
R610 GNDA.n574 GNDA.n573 585
R611 GNDA.n572 GNDA.n558 585
R612 GNDA.n580 GNDA.n579 585
R613 GNDA.n582 GNDA.n581 585
R614 GNDA.n556 GNDA.n555 585
R615 GNDA.n1891 GNDA.n1890 585
R616 GNDA.n1890 GNDA.n1889 585
R617 GNDA.n1098 GNDA.n513 585
R618 GNDA.n1122 GNDA.n1100 585
R619 GNDA.n1124 GNDA.n1123 585
R620 GNDA.n1120 GNDA.n1119 585
R621 GNDA.n1118 GNDA.n1117 585
R622 GNDA.n1113 GNDA.n1112 585
R623 GNDA.n1111 GNDA.n1110 585
R624 GNDA.n1106 GNDA.n1105 585
R625 GNDA.n1104 GNDA.n1025 585
R626 GNDA.n1132 GNDA.n1131 585
R627 GNDA.n1134 GNDA.n1133 585
R628 GNDA.n1138 GNDA.n1136 585
R629 GNDA.n749 GNDA.n748 585
R630 GNDA.n751 GNDA.n679 585
R631 GNDA.n753 GNDA.n752 585
R632 GNDA.n754 GNDA.n678 585
R633 GNDA.n756 GNDA.n755 585
R634 GNDA.n758 GNDA.n676 585
R635 GNDA.n760 GNDA.n759 585
R636 GNDA.n761 GNDA.n675 585
R637 GNDA.n763 GNDA.n762 585
R638 GNDA.n765 GNDA.n673 585
R639 GNDA.n767 GNDA.n766 585
R640 GNDA.n768 GNDA.n672 585
R641 GNDA.n692 GNDA.n113 585
R642 GNDA.n693 GNDA.n691 585
R643 GNDA.n695 GNDA.n694 585
R644 GNDA.n697 GNDA.n688 585
R645 GNDA.n699 GNDA.n698 585
R646 GNDA.n700 GNDA.n687 585
R647 GNDA.n702 GNDA.n701 585
R648 GNDA.n704 GNDA.n685 585
R649 GNDA.n706 GNDA.n705 585
R650 GNDA.n707 GNDA.n684 585
R651 GNDA.n709 GNDA.n708 585
R652 GNDA.n711 GNDA.n682 585
R653 GNDA.n2088 GNDA.n2087 585
R654 GNDA.n2089 GNDA.n122 585
R655 GNDA.n2091 GNDA.n2090 585
R656 GNDA.n2093 GNDA.n120 585
R657 GNDA.n2095 GNDA.n2094 585
R658 GNDA.n2096 GNDA.n119 585
R659 GNDA.n2098 GNDA.n2097 585
R660 GNDA.n2100 GNDA.n117 585
R661 GNDA.n2102 GNDA.n2101 585
R662 GNDA.n2103 GNDA.n116 585
R663 GNDA.n2105 GNDA.n2104 585
R664 GNDA.n2107 GNDA.n115 585
R665 GNDA.n487 GNDA.n486 585
R666 GNDA.n1949 GNDA.n487 585
R667 GNDA.n1459 GNDA.n1458 585
R668 GNDA.n1456 GNDA.n1300 585
R669 GNDA.n1347 GNDA.n1346 585
R670 GNDA.n1451 GNDA.n1450 585
R671 GNDA.n1449 GNDA.n1448 585
R672 GNDA.n1375 GNDA.n1351 585
R673 GNDA.n1377 GNDA.n1376 585
R674 GNDA.n1382 GNDA.n1381 585
R675 GNDA.n1380 GNDA.n1373 585
R676 GNDA.n1388 GNDA.n1387 585
R677 GNDA.n1390 GNDA.n1389 585
R678 GNDA.n1371 GNDA.n1370 585
R679 GNDA.n1947 GNDA.n488 585
R680 GNDA.n1949 GNDA.n488 585
R681 GNDA.n1950 GNDA.n486 585
R682 GNDA.n1950 GNDA.n1949 585
R683 GNDA.n1182 GNDA.n485 585
R684 GNDA.n1293 GNDA.n1292 585
R685 GNDA.n1184 GNDA.n1181 585
R686 GNDA.n1287 GNDA.n1286 585
R687 GNDA.n1285 GNDA.n1284 585
R688 GNDA.n1210 GNDA.n1188 585
R689 GNDA.n1212 GNDA.n1211 585
R690 GNDA.n1217 GNDA.n1216 585
R691 GNDA.n1215 GNDA.n1208 585
R692 GNDA.n1223 GNDA.n1222 585
R693 GNDA.n1225 GNDA.n1224 585
R694 GNDA.n1175 GNDA.n491 585
R695 GNDA.n1948 GNDA.n1947 585
R696 GNDA.n1949 GNDA.n1948 585
R697 GNDA.n492 GNDA.n490 585
R698 GNDA.n1538 GNDA.n1475 585
R699 GNDA.n1548 GNDA.n1547 585
R700 GNDA.n1550 GNDA.n1473 585
R701 GNDA.n1553 GNDA.n1552 585
R702 GNDA.n1554 GNDA.n1469 585
R703 GNDA.n1563 GNDA.n1562 585
R704 GNDA.n1565 GNDA.n1468 585
R705 GNDA.n1568 GNDA.n1567 585
R706 GNDA.n1569 GNDA.n1462 585
R707 GNDA.n1578 GNDA.n1577 585
R708 GNDA.n1580 GNDA.n1172 585
R709 GNDA.n919 GNDA.n918 585
R710 GNDA.n917 GNDA.n671 585
R711 GNDA.n916 GNDA.n915 585
R712 GNDA.n914 GNDA.n913 585
R713 GNDA.n912 GNDA.n911 585
R714 GNDA.n910 GNDA.n909 585
R715 GNDA.n908 GNDA.n907 585
R716 GNDA.n906 GNDA.n905 585
R717 GNDA.n904 GNDA.n903 585
R718 GNDA.n902 GNDA.n901 585
R719 GNDA.n900 GNDA.n899 585
R720 GNDA.n1763 GNDA.n665 585
R721 GNDA.n1322 GNDA.n1321 585
R722 GNDA.n1324 GNDA.n1323 585
R723 GNDA.n1326 GNDA.n1325 585
R724 GNDA.n1328 GNDA.n1327 585
R725 GNDA.n1330 GNDA.n1329 585
R726 GNDA.n1332 GNDA.n1331 585
R727 GNDA.n1334 GNDA.n1333 585
R728 GNDA.n1336 GNDA.n1335 585
R729 GNDA.n1338 GNDA.n1337 585
R730 GNDA.n1340 GNDA.n1339 585
R731 GNDA.n1342 GNDA.n1341 585
R732 GNDA.n1763 GNDA.n664 585
R733 GNDA.n1761 GNDA.n1760 585
R734 GNDA.n1759 GNDA.n922 585
R735 GNDA.n1758 GNDA.n921 585
R736 GNDA.n1763 GNDA.n921 585
R737 GNDA.n1757 GNDA.n1756 585
R738 GNDA.n1755 GNDA.n1754 585
R739 GNDA.n1753 GNDA.n1752 585
R740 GNDA.n1751 GNDA.n1750 585
R741 GNDA.n1749 GNDA.n1748 585
R742 GNDA.n1747 GNDA.n1746 585
R743 GNDA.n1745 GNDA.n1744 585
R744 GNDA.n653 GNDA.n652 585
R745 GNDA.n1766 GNDA.n1765 585
R746 GNDA.n1766 GNDA.n651 585
R747 GNDA.n2226 GNDA.n46 585
R748 GNDA.n2229 GNDA.n2228 585
R749 GNDA.n2230 GNDA.n2229 585
R750 GNDA.n2221 GNDA.n2220 585
R751 GNDA.n2164 GNDA.n89 585
R752 GNDA.n2165 GNDA.n2164 585
R753 GNDA.n897 GNDA.n896 585
R754 GNDA.n896 GNDA.n895 585
R755 GNDA.n773 GNDA.n771 585
R756 GNDA.n894 GNDA.n771 585
R757 GNDA.n892 GNDA.n891 585
R758 GNDA.n893 GNDA.n892 585
R759 GNDA.n775 GNDA.n772 585
R760 GNDA.n807 GNDA.n772 585
R761 GNDA.n806 GNDA.n805 585
R762 GNDA.n808 GNDA.n806 585
R763 GNDA.n811 GNDA.n810 585
R764 GNDA.n810 GNDA.n809 585
R765 GNDA.n812 GNDA.n801 585
R766 GNDA.n801 GNDA.n800 585
R767 GNDA.n823 GNDA.n822 585
R768 GNDA.n824 GNDA.n823 585
R769 GNDA.n817 GNDA.n799 585
R770 GNDA.n825 GNDA.n799 585
R771 GNDA.n827 GNDA.n798 585
R772 GNDA.n827 GNDA.n826 585
R773 GNDA.n831 GNDA.n830 585
R774 GNDA.n830 GNDA.n829 585
R775 GNDA.n796 GNDA.n88 585
R776 GNDA.n828 GNDA.n88 585
R777 GNDA.n2146 GNDA.n99 585
R778 GNDA.n99 GNDA.n80 585
R779 GNDA.n2156 GNDA.n89 585
R780 GNDA.n2156 GNDA.n85 585
R781 GNDA.n2155 GNDA.n95 585
R782 GNDA.n2155 GNDA.n2154 585
R783 GNDA.n372 GNDA.n94 585
R784 GNDA.n96 GNDA.n94 585
R785 GNDA.n389 GNDA.n388 585
R786 GNDA.n388 GNDA.n387 585
R787 GNDA.n376 GNDA.n374 585
R788 GNDA.n386 GNDA.n374 585
R789 GNDA.n384 GNDA.n383 585
R790 GNDA.n385 GNDA.n384 585
R791 GNDA.n379 GNDA.n282 585
R792 GNDA.n375 GNDA.n282 585
R793 GNDA.n397 GNDA.n396 585
R794 GNDA.n398 GNDA.n397 585
R795 GNDA.n284 GNDA.n283 585
R796 GNDA.n310 GNDA.n283 585
R797 GNDA.n309 GNDA.n308 585
R798 GNDA.n311 GNDA.n309 585
R799 GNDA.n314 GNDA.n313 585
R800 GNDA.n313 GNDA.n312 585
R801 GNDA.n315 GNDA.n98 585
R802 GNDA.n98 GNDA.n97 585
R803 GNDA.n2149 GNDA.n2148 585
R804 GNDA.n2150 GNDA.n2149 585
R805 GNDA.n2146 GNDA.n2145 585
R806 GNDA.n2145 GNDA.n77 585
R807 GNDA.n101 GNDA.n76 585
R808 GNDA.n2192 GNDA.n76 585
R809 GNDA.n2194 GNDA.n74 585
R810 GNDA.n2194 GNDA.n2193 585
R811 GNDA.n2210 GNDA.n2209 585
R812 GNDA.n2209 GNDA.n2208 585
R813 GNDA.n2197 GNDA.n2195 585
R814 GNDA.n2207 GNDA.n2195 585
R815 GNDA.n2205 GNDA.n2204 585
R816 GNDA.n2206 GNDA.n2205 585
R817 GNDA.n2200 GNDA.n51 585
R818 GNDA.n2196 GNDA.n51 585
R819 GNDA.n2218 GNDA.n2217 585
R820 GNDA.n2219 GNDA.n2218 585
R821 GNDA.n53 GNDA.n52 585
R822 GNDA.n1993 GNDA.n52 585
R823 GNDA.n2056 GNDA.n2055 585
R824 GNDA.n2057 GNDA.n2056 585
R825 GNDA.n2052 GNDA.n1991 585
R826 GNDA.n2058 GNDA.n1991 585
R827 GNDA.n2060 GNDA.n1992 585
R828 GNDA.n2060 GNDA.n2059 585
R829 GNDA.n2061 GNDA.n1990 585
R830 GNDA.n2061 GNDA.n37 585
R831 GNDA.n419 GNDA.n418 585
R832 GNDA.n420 GNDA.n419 585
R833 GNDA.n408 GNDA.n406 585
R834 GNDA.n412 GNDA.n411 585
R835 GNDA.n414 GNDA.n413 585
R836 GNDA.n184 GNDA.n149 553.051
R837 GNDA.n2253 GNDA.n2252 544.918
R838 GNDA.n174 GNDA.t288 524.808
R839 GNDA.n181 GNDA.t276 524.808
R840 GNDA.n10 GNDA.t248 524.808
R841 GNDA.n28 GNDA.t240 524.808
R842 GNDA.t227 GNDA.n432 512.884
R843 GNDA.t227 GNDA.n424 512.884
R844 GNDA.n2262 GNDA.t251 508.743
R845 GNDA.n155 GNDA.t291 508.743
R846 GNDA.n198 GNDA.t315 508.743
R847 GNDA.n2257 GNDA.t299 508.743
R848 GNDA.n208 GNDA.t307 499.442
R849 GNDA.n188 GNDA.t317 499.442
R850 GNDA.n152 GNDA.t302 499.442
R851 GNDA.n2255 GNDA.t312 499.442
R852 GNDA.n204 GNDA.t246 475.976
R853 GNDA.n204 GNDA.t233 475.976
R854 GNDA.n192 GNDA.t305 475.976
R855 GNDA.n192 GNDA.t297 475.976
R856 GNDA.n132 GNDA.t267 409.067
R857 GNDA.n2168 GNDA.t279 409.067
R858 GNDA.n2177 GNDA.t309 409.067
R859 GNDA.n2182 GNDA.t254 409.067
R860 GNDA.n2189 GNDA.t263 409.067
R861 GNDA.n2240 GNDA.t257 409.067
R862 GNDA.t37 GNDA.n35 396.445
R863 GNDA.t227 GNDA.n433 391.411
R864 GNDA.t227 GNDA.n425 391.411
R865 GNDA.n258 GNDA.t294 338.034
R866 GNDA.n246 GNDA.t285 338.034
R867 GNDA.t90 GNDA.t92 333.793
R868 GNDA.t154 GNDA.t90 333.793
R869 GNDA.t179 GNDA.t154 333.793
R870 GNDA.t94 GNDA.t129 333.793
R871 GNDA.t129 GNDA.t55 333.793
R872 GNDA.t55 GNDA.t14 333.793
R873 GNDA.t8 GNDA.t114 333.793
R874 GNDA.t114 GNDA.t0 333.793
R875 GNDA.t227 GNDA.n81 172.876
R876 GNDA.t227 GNDA.n83 172.876
R877 GNDA.t227 GNDA.n84 172.615
R878 GNDA.t227 GNDA.n48 172.615
R879 GNDA.n2261 GNDA.n2260 296.158
R880 GNDA.n157 GNDA.n156 296.158
R881 GNDA.n200 GNDA.n199 296.158
R882 GNDA.n2259 GNDA.n2258 296.158
R883 GNDA.t227 GNDA.t131 294.625
R884 GNDA.n207 GNDA.n149 292.5
R885 GNDA.n201 GNDA.n200 292.5
R886 GNDA.n2259 GNDA.n3 292.5
R887 GNDA.n2253 GNDA.n5 292.5
R888 GNDA.n151 GNDA.n149 292.5
R889 GNDA.n2254 GNDA.n2253 292.5
R890 GNDA.n1764 GNDA.n1763 264.301
R891 GNDA.n2065 GNDA.n2064 264.301
R892 GNDA.n1583 GNDA.n1582 264.301
R893 GNDA.n1608 GNDA.n1607 264.301
R894 GNDA.n898 GNDA.n769 264.301
R895 GNDA.n1344 GNDA.n1343 264.301
R896 GNDA.n1721 GNDA.n935 259.416
R897 GNDA.n1977 GNDA.n454 259.416
R898 GNDA.n749 GNDA.n681 259.416
R899 GNDA.n2111 GNDA.n113 259.416
R900 GNDA.n1916 GNDA.n1914 259.416
R901 GNDA.n1656 GNDA.n957 259.416
R902 GNDA.n1603 GNDA.n1141 259.416
R903 GNDA.n2087 GNDA.n2086 259.416
R904 GNDA.n1628 GNDA.n1012 259.416
R905 GNDA.n1847 GNDA.n1790 258.334
R906 GNDA.n1427 GNDA.n1368 258.334
R907 GNDA.n870 GNDA.n869 258.334
R908 GNDA.n354 GNDA.n353 258.334
R909 GNDA.n1262 GNDA.n1205 258.334
R910 GNDA.n621 GNDA.n620 258.334
R911 GNDA.n1523 GNDA.n1481 258.334
R912 GNDA.n2013 GNDA.n2012 258.334
R913 GNDA.n1081 GNDA.n1080 258.334
R914 GNDA.n260 GNDA.t176 257.932
R915 GNDA.n244 GNDA.t124 257.932
R916 GNDA.n1943 GNDA.n127 254.34
R917 GNDA.n1940 GNDA.n127 254.34
R918 GNDA.n503 GNDA.n127 254.34
R919 GNDA.n1929 GNDA.n127 254.34
R920 GNDA.n1926 GNDA.n127 254.34
R921 GNDA.n1915 GNDA.n127 254.34
R922 GNDA.n1919 GNDA.n435 254.34
R923 GNDA.n1921 GNDA.n435 254.34
R924 GNDA.n1933 GNDA.n435 254.34
R925 GNDA.n1936 GNDA.n435 254.34
R926 GNDA.n498 GNDA.n435 254.34
R927 GNDA.n2139 GNDA.n83 254.34
R928 GNDA.n2136 GNDA.n83 254.34
R929 GNDA.n2126 GNDA.n83 254.34
R930 GNDA.n2124 GNDA.n83 254.34
R931 GNDA.n2114 GNDA.n83 254.34
R932 GNDA.n2112 GNDA.n83 254.34
R933 GNDA.n2108 GNDA.n48 254.34
R934 GNDA.n2118 GNDA.n48 254.34
R935 GNDA.n2120 GNDA.n48 254.34
R936 GNDA.n2130 GNDA.n48 254.34
R937 GNDA.n2132 GNDA.n48 254.34
R938 GNDA.n2143 GNDA.n48 254.34
R939 GNDA.n2162 GNDA.n81 254.34
R940 GNDA.n726 GNDA.n81 254.34
R941 GNDA.n724 GNDA.n81 254.34
R942 GNDA.n721 GNDA.n81 254.34
R943 GNDA.n716 GNDA.n81 254.34
R944 GNDA.n713 GNDA.n81 254.34
R945 GNDA.n744 GNDA.n84 254.34
R946 GNDA.n712 GNDA.n84 254.34
R947 GNDA.n737 GNDA.n84 254.34
R948 GNDA.n731 GNDA.n84 254.34
R949 GNDA.n729 GNDA.n84 254.34
R950 GNDA.n2158 GNDA.n84 254.34
R951 GNDA.n482 GNDA.n481 254.34
R952 GNDA.n481 GNDA.n480 254.34
R953 GNDA.n481 GNDA.n479 254.34
R954 GNDA.n481 GNDA.n478 254.34
R955 GNDA.n481 GNDA.n477 254.34
R956 GNDA.n481 GNDA.n476 254.34
R957 GNDA.n1972 GNDA.n1971 254.34
R958 GNDA.n1971 GNDA.n1970 254.34
R959 GNDA.n1971 GNDA.n464 254.34
R960 GNDA.n1971 GNDA.n463 254.34
R961 GNDA.n1971 GNDA.n462 254.34
R962 GNDA.n1971 GNDA.n461 254.34
R963 GNDA.n1979 GNDA.n1978 254.34
R964 GNDA.n1979 GNDA.n452 254.34
R965 GNDA.n1979 GNDA.n451 254.34
R966 GNDA.n1979 GNDA.n450 254.34
R967 GNDA.n1979 GNDA.n449 254.34
R968 GNDA.n1979 GNDA.n448 254.34
R969 GNDA.n1979 GNDA.n447 254.34
R970 GNDA.n1979 GNDA.n446 254.34
R971 GNDA.n1979 GNDA.n445 254.34
R972 GNDA.n1979 GNDA.n444 254.34
R973 GNDA.n1979 GNDA.n443 254.34
R974 GNDA.n1979 GNDA.n442 254.34
R975 GNDA.n1979 GNDA.n441 254.34
R976 GNDA.n1979 GNDA.n440 254.34
R977 GNDA.n1979 GNDA.n439 254.34
R978 GNDA.n1979 GNDA.n438 254.34
R979 GNDA.n1979 GNDA.n437 254.34
R980 GNDA.n1979 GNDA.n436 254.34
R981 GNDA.n1881 GNDA.n1880 254.34
R982 GNDA.n1881 GNDA.n649 254.34
R983 GNDA.n1881 GNDA.n648 254.34
R984 GNDA.n1881 GNDA.n647 254.34
R985 GNDA.n1881 GNDA.n646 254.34
R986 GNDA.n1881 GNDA.n645 254.34
R987 GNDA.n1882 GNDA.n1881 254.34
R988 GNDA.n1881 GNDA.n644 254.34
R989 GNDA.n1881 GNDA.n531 254.34
R990 GNDA.n1881 GNDA.n530 254.34
R991 GNDA.n1881 GNDA.n529 254.34
R992 GNDA.n1881 GNDA.n528 254.34
R993 GNDA.n1881 GNDA.n527 254.34
R994 GNDA.n1881 GNDA.n526 254.34
R995 GNDA.n1881 GNDA.n525 254.34
R996 GNDA.n1881 GNDA.n524 254.34
R997 GNDA.n1881 GNDA.n523 254.34
R998 GNDA.n1881 GNDA.n522 254.34
R999 GNDA.n750 GNDA.n82 254.34
R1000 GNDA.n680 GNDA.n82 254.34
R1001 GNDA.n757 GNDA.n82 254.34
R1002 GNDA.n677 GNDA.n82 254.34
R1003 GNDA.n764 GNDA.n82 254.34
R1004 GNDA.n674 GNDA.n82 254.34
R1005 GNDA.n690 GNDA.n82 254.34
R1006 GNDA.n696 GNDA.n82 254.34
R1007 GNDA.n689 GNDA.n82 254.34
R1008 GNDA.n703 GNDA.n82 254.34
R1009 GNDA.n686 GNDA.n82 254.34
R1010 GNDA.n710 GNDA.n82 254.34
R1011 GNDA.n124 GNDA.n82 254.34
R1012 GNDA.n2092 GNDA.n82 254.34
R1013 GNDA.n121 GNDA.n82 254.34
R1014 GNDA.n2099 GNDA.n82 254.34
R1015 GNDA.n118 GNDA.n82 254.34
R1016 GNDA.n2106 GNDA.n82 254.34
R1017 GNDA.n1461 GNDA.n1460 254.34
R1018 GNDA.n1461 GNDA.n1299 254.34
R1019 GNDA.n1461 GNDA.n1298 254.34
R1020 GNDA.n1461 GNDA.n1297 254.34
R1021 GNDA.n1461 GNDA.n1296 254.34
R1022 GNDA.n1461 GNDA.n1295 254.34
R1023 GNDA.n1461 GNDA.n1294 254.34
R1024 GNDA.n1461 GNDA.n1180 254.34
R1025 GNDA.n1461 GNDA.n1179 254.34
R1026 GNDA.n1461 GNDA.n1178 254.34
R1027 GNDA.n1461 GNDA.n1177 254.34
R1028 GNDA.n1461 GNDA.n1176 254.34
R1029 GNDA.n1474 GNDA.n1461 254.34
R1030 GNDA.n1549 GNDA.n1461 254.34
R1031 GNDA.n1551 GNDA.n1461 254.34
R1032 GNDA.n1564 GNDA.n1461 254.34
R1033 GNDA.n1566 GNDA.n1461 254.34
R1034 GNDA.n1579 GNDA.n1461 254.34
R1035 GNDA.n1763 GNDA.n920 254.34
R1036 GNDA.n1763 GNDA.n670 254.34
R1037 GNDA.n1763 GNDA.n669 254.34
R1038 GNDA.n1763 GNDA.n668 254.34
R1039 GNDA.n1763 GNDA.n667 254.34
R1040 GNDA.n1763 GNDA.n666 254.34
R1041 GNDA.n1763 GNDA.n658 254.34
R1042 GNDA.n1763 GNDA.n659 254.34
R1043 GNDA.n1763 GNDA.n660 254.34
R1044 GNDA.n1763 GNDA.n661 254.34
R1045 GNDA.n1763 GNDA.n662 254.34
R1046 GNDA.n1763 GNDA.n663 254.34
R1047 GNDA.n1763 GNDA.n1762 254.34
R1048 GNDA.n1763 GNDA.n654 254.34
R1049 GNDA.n1763 GNDA.n655 254.34
R1050 GNDA.n1763 GNDA.n656 254.34
R1051 GNDA.n1763 GNDA.n657 254.34
R1052 GNDA.t227 GNDA.n944 250.349
R1053 GNDA.n1761 GNDA.n923 249.663
R1054 GNDA.n1321 GNDA.n1320 249.663
R1055 GNDA.n919 GNDA.n672 249.663
R1056 GNDA.n745 GNDA.n711 249.663
R1057 GNDA.n1973 GNDA.n459 249.663
R1058 GNDA.n1717 GNDA.n1680 249.663
R1059 GNDA.n1918 GNDA.n508 249.663
R1060 GNDA.n2109 GNDA.n2107 249.663
R1061 GNDA.n1652 GNDA.n1001 249.663
R1062 GNDA.n2229 GNDA.n46 246.25
R1063 GNDA.n2229 GNDA.n2220 246.25
R1064 GNDA.n419 GNDA.n406 246.25
R1065 GNDA.n413 GNDA.n412 246.25
R1066 GNDA.n2236 GNDA.n2235 241.643
R1067 GNDA.n2231 GNDA.n2230 241.643
R1068 GNDA.n2230 GNDA.n47 241.643
R1069 GNDA.n420 GNDA.n404 241.643
R1070 GNDA.n420 GNDA.n405 241.643
R1071 GNDA.n259 GNDA.t296 233
R1072 GNDA.n245 GNDA.t287 233
R1073 GNDA.n265 GNDA.n150 200.456
R1074 GNDA.n240 GNDA.n239 200.456
R1075 GNDA.n171 GNDA.t153 199.262
R1076 GNDA.n256 GNDA.n255 199.03
R1077 GNDA.n254 GNDA.n253 199.03
R1078 GNDA.n252 GNDA.n251 199.03
R1079 GNDA.n250 GNDA.n249 199.03
R1080 GNDA.n248 GNDA.n247 199.03
R1081 GNDA.n1669 GNDA.n946 197
R1082 GNDA.n1888 GNDA.n515 197
R1083 GNDA.n1370 GNDA.n487 197
R1084 GNDA.n2164 GNDA.n88 197
R1085 GNDA.n2149 GNDA.n99 197
R1086 GNDA.n1175 GNDA.n488 197
R1087 GNDA.n555 GNDA.n511 197
R1088 GNDA.n1581 GNDA.n1580 197
R1089 GNDA.n2063 GNDA.n2061 197
R1090 GNDA.n1606 GNDA.n1138 197
R1091 GNDA.n1879 GNDA.n651 187.249
R1092 GNDA.n1459 GNDA.n664 187.249
R1093 GNDA.n896 GNDA.n665 187.249
R1094 GNDA.n2156 GNDA.n2155 187.249
R1095 GNDA.n1950 GNDA.n485 187.249
R1096 GNDA.n1883 GNDA.n514 187.249
R1097 GNDA.n1948 GNDA.n490 187.249
R1098 GNDA.n2145 GNDA.n76 187.249
R1099 GNDA.n1890 GNDA.n513 187.249
R1100 GNDA.n2232 GNDA.n45 185
R1101 GNDA.n2224 GNDA.n2223 185
R1102 GNDA.n1849 GNDA.n1790 185
R1103 GNDA.n1863 GNDA.n1862 185
R1104 GNDA.n1861 GNDA.n1791 185
R1105 GNDA.n1860 GNDA.n1859 185
R1106 GNDA.n1858 GNDA.n1857 185
R1107 GNDA.n1856 GNDA.n1855 185
R1108 GNDA.n1854 GNDA.n1853 185
R1109 GNDA.n1852 GNDA.n1851 185
R1110 GNDA.n1850 GNDA.n1767 185
R1111 GNDA.n1832 GNDA.n1831 185
R1112 GNDA.n1834 GNDA.n1833 185
R1113 GNDA.n1836 GNDA.n1835 185
R1114 GNDA.n1838 GNDA.n1837 185
R1115 GNDA.n1840 GNDA.n1839 185
R1116 GNDA.n1842 GNDA.n1841 185
R1117 GNDA.n1844 GNDA.n1843 185
R1118 GNDA.n1846 GNDA.n1845 185
R1119 GNDA.n1848 GNDA.n1847 185
R1120 GNDA.n1814 GNDA.n1813 185
R1121 GNDA.n1816 GNDA.n1815 185
R1122 GNDA.n1818 GNDA.n1817 185
R1123 GNDA.n1820 GNDA.n1819 185
R1124 GNDA.n1822 GNDA.n1821 185
R1125 GNDA.n1824 GNDA.n1823 185
R1126 GNDA.n1826 GNDA.n1825 185
R1127 GNDA.n1828 GNDA.n1827 185
R1128 GNDA.n1830 GNDA.n1829 185
R1129 GNDA.n1812 GNDA.n1811 185
R1130 GNDA.n1806 GNDA.n1805 185
R1131 GNDA.n1804 GNDA.n1803 185
R1132 GNDA.n1799 GNDA.n1798 185
R1133 GNDA.n1794 GNDA.n1775 185
R1134 GNDA.n1867 GNDA.n1866 185
R1135 GNDA.n1774 GNDA.n1772 185
R1136 GNDA.n1873 GNDA.n1872 185
R1137 GNDA.n1875 GNDA.n1874 185
R1138 GNDA.n1429 GNDA.n1368 185
R1139 GNDA.n1443 GNDA.n1442 185
R1140 GNDA.n1441 GNDA.n1369 185
R1141 GNDA.n1440 GNDA.n1439 185
R1142 GNDA.n1438 GNDA.n1437 185
R1143 GNDA.n1436 GNDA.n1435 185
R1144 GNDA.n1434 GNDA.n1433 185
R1145 GNDA.n1432 GNDA.n1431 185
R1146 GNDA.n1430 GNDA.n1345 185
R1147 GNDA.n1412 GNDA.n1411 185
R1148 GNDA.n1414 GNDA.n1413 185
R1149 GNDA.n1416 GNDA.n1415 185
R1150 GNDA.n1418 GNDA.n1417 185
R1151 GNDA.n1420 GNDA.n1419 185
R1152 GNDA.n1422 GNDA.n1421 185
R1153 GNDA.n1424 GNDA.n1423 185
R1154 GNDA.n1426 GNDA.n1425 185
R1155 GNDA.n1428 GNDA.n1427 185
R1156 GNDA.n1394 GNDA.n1393 185
R1157 GNDA.n1396 GNDA.n1395 185
R1158 GNDA.n1398 GNDA.n1397 185
R1159 GNDA.n1400 GNDA.n1399 185
R1160 GNDA.n1402 GNDA.n1401 185
R1161 GNDA.n1404 GNDA.n1403 185
R1162 GNDA.n1406 GNDA.n1405 185
R1163 GNDA.n1408 GNDA.n1407 185
R1164 GNDA.n1410 GNDA.n1409 185
R1165 GNDA.n1392 GNDA.n1391 185
R1166 GNDA.n1386 GNDA.n1385 185
R1167 GNDA.n1384 GNDA.n1383 185
R1168 GNDA.n1379 GNDA.n1378 185
R1169 GNDA.n1374 GNDA.n1353 185
R1170 GNDA.n1447 GNDA.n1446 185
R1171 GNDA.n1352 GNDA.n1350 185
R1172 GNDA.n1453 GNDA.n1452 185
R1173 GNDA.n1455 GNDA.n1454 185
R1174 GNDA.n871 GNDA.n870 185
R1175 GNDA.n873 GNDA.n872 185
R1176 GNDA.n875 GNDA.n874 185
R1177 GNDA.n877 GNDA.n876 185
R1178 GNDA.n879 GNDA.n878 185
R1179 GNDA.n881 GNDA.n880 185
R1180 GNDA.n883 GNDA.n882 185
R1181 GNDA.n884 GNDA.n794 185
R1182 GNDA.n886 GNDA.n885 185
R1183 GNDA.n853 GNDA.n852 185
R1184 GNDA.n855 GNDA.n854 185
R1185 GNDA.n857 GNDA.n856 185
R1186 GNDA.n859 GNDA.n858 185
R1187 GNDA.n861 GNDA.n860 185
R1188 GNDA.n863 GNDA.n862 185
R1189 GNDA.n865 GNDA.n864 185
R1190 GNDA.n867 GNDA.n866 185
R1191 GNDA.n869 GNDA.n868 185
R1192 GNDA.n835 GNDA.n834 185
R1193 GNDA.n837 GNDA.n836 185
R1194 GNDA.n839 GNDA.n838 185
R1195 GNDA.n841 GNDA.n840 185
R1196 GNDA.n843 GNDA.n842 185
R1197 GNDA.n845 GNDA.n844 185
R1198 GNDA.n847 GNDA.n846 185
R1199 GNDA.n849 GNDA.n848 185
R1200 GNDA.n851 GNDA.n850 185
R1201 GNDA.n833 GNDA.n832 185
R1202 GNDA.n819 GNDA.n818 185
R1203 GNDA.n821 GNDA.n820 185
R1204 GNDA.n816 GNDA.n815 185
R1205 GNDA.n814 GNDA.n813 185
R1206 GNDA.n803 GNDA.n802 185
R1207 GNDA.n804 GNDA.n777 185
R1208 GNDA.n890 GNDA.n889 185
R1209 GNDA.n776 GNDA.n774 185
R1210 GNDA.n355 GNDA.n354 185
R1211 GNDA.n357 GNDA.n356 185
R1212 GNDA.n359 GNDA.n358 185
R1213 GNDA.n361 GNDA.n360 185
R1214 GNDA.n363 GNDA.n362 185
R1215 GNDA.n365 GNDA.n364 185
R1216 GNDA.n367 GNDA.n366 185
R1217 GNDA.n369 GNDA.n368 185
R1218 GNDA.n370 GNDA.n303 185
R1219 GNDA.n337 GNDA.n336 185
R1220 GNDA.n339 GNDA.n338 185
R1221 GNDA.n341 GNDA.n340 185
R1222 GNDA.n343 GNDA.n342 185
R1223 GNDA.n345 GNDA.n344 185
R1224 GNDA.n347 GNDA.n346 185
R1225 GNDA.n349 GNDA.n348 185
R1226 GNDA.n351 GNDA.n350 185
R1227 GNDA.n353 GNDA.n352 185
R1228 GNDA.n319 GNDA.n318 185
R1229 GNDA.n321 GNDA.n320 185
R1230 GNDA.n323 GNDA.n322 185
R1231 GNDA.n325 GNDA.n324 185
R1232 GNDA.n327 GNDA.n326 185
R1233 GNDA.n329 GNDA.n328 185
R1234 GNDA.n331 GNDA.n330 185
R1235 GNDA.n333 GNDA.n332 185
R1236 GNDA.n335 GNDA.n334 185
R1237 GNDA.n317 GNDA.n316 185
R1238 GNDA.n306 GNDA.n305 185
R1239 GNDA.n307 GNDA.n286 185
R1240 GNDA.n395 GNDA.n394 185
R1241 GNDA.n378 GNDA.n285 185
R1242 GNDA.n382 GNDA.n381 185
R1243 GNDA.n380 GNDA.n377 185
R1244 GNDA.n373 GNDA.n304 185
R1245 GNDA.n391 GNDA.n390 185
R1246 GNDA.n1264 GNDA.n1205 185
R1247 GNDA.n1279 GNDA.n1278 185
R1248 GNDA.n1277 GNDA.n1206 185
R1249 GNDA.n1276 GNDA.n1275 185
R1250 GNDA.n1274 GNDA.n1273 185
R1251 GNDA.n1272 GNDA.n1271 185
R1252 GNDA.n1270 GNDA.n1269 185
R1253 GNDA.n1268 GNDA.n1267 185
R1254 GNDA.n1266 GNDA.n1265 185
R1255 GNDA.n1247 GNDA.n1246 185
R1256 GNDA.n1249 GNDA.n1248 185
R1257 GNDA.n1251 GNDA.n1250 185
R1258 GNDA.n1253 GNDA.n1252 185
R1259 GNDA.n1255 GNDA.n1254 185
R1260 GNDA.n1257 GNDA.n1256 185
R1261 GNDA.n1259 GNDA.n1258 185
R1262 GNDA.n1261 GNDA.n1260 185
R1263 GNDA.n1263 GNDA.n1262 185
R1264 GNDA.n1229 GNDA.n1228 185
R1265 GNDA.n1231 GNDA.n1230 185
R1266 GNDA.n1233 GNDA.n1232 185
R1267 GNDA.n1235 GNDA.n1234 185
R1268 GNDA.n1237 GNDA.n1236 185
R1269 GNDA.n1239 GNDA.n1238 185
R1270 GNDA.n1241 GNDA.n1240 185
R1271 GNDA.n1243 GNDA.n1242 185
R1272 GNDA.n1245 GNDA.n1244 185
R1273 GNDA.n1227 GNDA.n1226 185
R1274 GNDA.n1221 GNDA.n1220 185
R1275 GNDA.n1219 GNDA.n1218 185
R1276 GNDA.n1214 GNDA.n1213 185
R1277 GNDA.n1209 GNDA.n1190 185
R1278 GNDA.n1283 GNDA.n1282 185
R1279 GNDA.n1189 GNDA.n1187 185
R1280 GNDA.n1289 GNDA.n1288 185
R1281 GNDA.n1291 GNDA.n1290 185
R1282 GNDA.n622 GNDA.n621 185
R1283 GNDA.n624 GNDA.n623 185
R1284 GNDA.n626 GNDA.n625 185
R1285 GNDA.n628 GNDA.n627 185
R1286 GNDA.n630 GNDA.n629 185
R1287 GNDA.n632 GNDA.n631 185
R1288 GNDA.n634 GNDA.n633 185
R1289 GNDA.n635 GNDA.n554 185
R1290 GNDA.n637 GNDA.n636 185
R1291 GNDA.n604 GNDA.n603 185
R1292 GNDA.n606 GNDA.n605 185
R1293 GNDA.n608 GNDA.n607 185
R1294 GNDA.n610 GNDA.n609 185
R1295 GNDA.n612 GNDA.n611 185
R1296 GNDA.n614 GNDA.n613 185
R1297 GNDA.n616 GNDA.n615 185
R1298 GNDA.n618 GNDA.n617 185
R1299 GNDA.n620 GNDA.n619 185
R1300 GNDA.n586 GNDA.n585 185
R1301 GNDA.n588 GNDA.n587 185
R1302 GNDA.n590 GNDA.n589 185
R1303 GNDA.n592 GNDA.n591 185
R1304 GNDA.n594 GNDA.n593 185
R1305 GNDA.n596 GNDA.n595 185
R1306 GNDA.n598 GNDA.n597 185
R1307 GNDA.n600 GNDA.n599 185
R1308 GNDA.n602 GNDA.n601 185
R1309 GNDA.n584 GNDA.n583 185
R1310 GNDA.n578 GNDA.n577 185
R1311 GNDA.n576 GNDA.n575 185
R1312 GNDA.n571 GNDA.n570 185
R1313 GNDA.n569 GNDA.n568 185
R1314 GNDA.n563 GNDA.n562 185
R1315 GNDA.n559 GNDA.n537 185
R1316 GNDA.n641 GNDA.n640 185
R1317 GNDA.n536 GNDA.n534 185
R1318 GNDA.n1523 GNDA.n1522 185
R1319 GNDA.n1525 GNDA.n1480 185
R1320 GNDA.n1528 GNDA.n1527 185
R1321 GNDA.n1529 GNDA.n1479 185
R1322 GNDA.n1531 GNDA.n1530 185
R1323 GNDA.n1533 GNDA.n1478 185
R1324 GNDA.n1536 GNDA.n1535 185
R1325 GNDA.n1537 GNDA.n1477 185
R1326 GNDA.n1541 GNDA.n1540 185
R1327 GNDA.n1505 GNDA.n1485 185
R1328 GNDA.n1507 GNDA.n1506 185
R1329 GNDA.n1509 GNDA.n1484 185
R1330 GNDA.n1512 GNDA.n1511 185
R1331 GNDA.n1513 GNDA.n1483 185
R1332 GNDA.n1515 GNDA.n1514 185
R1333 GNDA.n1517 GNDA.n1482 185
R1334 GNDA.n1520 GNDA.n1519 185
R1335 GNDA.n1521 GNDA.n1481 185
R1336 GNDA.n1575 GNDA.n1574 185
R1337 GNDA.n1490 GNDA.n1464 185
R1338 GNDA.n1492 GNDA.n1491 185
R1339 GNDA.n1494 GNDA.n1488 185
R1340 GNDA.n1496 GNDA.n1495 185
R1341 GNDA.n1497 GNDA.n1487 185
R1342 GNDA.n1499 GNDA.n1498 185
R1343 GNDA.n1501 GNDA.n1486 185
R1344 GNDA.n1504 GNDA.n1503 185
R1345 GNDA.n1573 GNDA.n1463 185
R1346 GNDA.n1571 GNDA.n1570 185
R1347 GNDA.n1467 GNDA.n1466 185
R1348 GNDA.n1561 GNDA.n1560 185
R1349 GNDA.n1558 GNDA.n1470 185
R1350 GNDA.n1556 GNDA.n1555 185
R1351 GNDA.n1472 GNDA.n1471 185
R1352 GNDA.n1546 GNDA.n1545 185
R1353 GNDA.n1543 GNDA.n1476 185
R1354 GNDA.n2012 GNDA.n2011 185
R1355 GNDA.n2010 GNDA.n2009 185
R1356 GNDA.n2008 GNDA.n2007 185
R1357 GNDA.n2006 GNDA.n2005 185
R1358 GNDA.n2004 GNDA.n2003 185
R1359 GNDA.n2002 GNDA.n2001 185
R1360 GNDA.n2000 GNDA.n1999 185
R1361 GNDA.n1998 GNDA.n1997 185
R1362 GNDA.n1996 GNDA.n72 185
R1363 GNDA.n2030 GNDA.n2029 185
R1364 GNDA.n2028 GNDA.n2027 185
R1365 GNDA.n2026 GNDA.n2025 185
R1366 GNDA.n2024 GNDA.n2023 185
R1367 GNDA.n2022 GNDA.n2021 185
R1368 GNDA.n2020 GNDA.n2019 185
R1369 GNDA.n2018 GNDA.n2017 185
R1370 GNDA.n2016 GNDA.n2015 185
R1371 GNDA.n2014 GNDA.n2013 185
R1372 GNDA.n2049 GNDA.n2048 185
R1373 GNDA.n2046 GNDA.n2045 185
R1374 GNDA.n2044 GNDA.n2043 185
R1375 GNDA.n2042 GNDA.n2041 185
R1376 GNDA.n2040 GNDA.n2039 185
R1377 GNDA.n2038 GNDA.n2037 185
R1378 GNDA.n2036 GNDA.n2035 185
R1379 GNDA.n2034 GNDA.n2033 185
R1380 GNDA.n2032 GNDA.n2031 185
R1381 GNDA.n2051 GNDA.n2050 185
R1382 GNDA.n2054 GNDA.n2053 185
R1383 GNDA.n1994 GNDA.n55 185
R1384 GNDA.n2216 GNDA.n2215 185
R1385 GNDA.n2199 GNDA.n54 185
R1386 GNDA.n2203 GNDA.n2202 185
R1387 GNDA.n2201 GNDA.n2198 185
R1388 GNDA.n75 GNDA.n73 185
R1389 GNDA.n2212 GNDA.n2211 185
R1390 GNDA.n1082 GNDA.n1081 185
R1391 GNDA.n1084 GNDA.n1083 185
R1392 GNDA.n1086 GNDA.n1085 185
R1393 GNDA.n1088 GNDA.n1087 185
R1394 GNDA.n1090 GNDA.n1089 185
R1395 GNDA.n1092 GNDA.n1091 185
R1396 GNDA.n1094 GNDA.n1093 185
R1397 GNDA.n1096 GNDA.n1095 185
R1398 GNDA.n1097 GNDA.n1045 185
R1399 GNDA.n1064 GNDA.n1063 185
R1400 GNDA.n1066 GNDA.n1065 185
R1401 GNDA.n1068 GNDA.n1067 185
R1402 GNDA.n1070 GNDA.n1069 185
R1403 GNDA.n1072 GNDA.n1071 185
R1404 GNDA.n1074 GNDA.n1073 185
R1405 GNDA.n1076 GNDA.n1075 185
R1406 GNDA.n1078 GNDA.n1077 185
R1407 GNDA.n1080 GNDA.n1079 185
R1408 GNDA.n1037 GNDA.n1023 185
R1409 GNDA.n1048 GNDA.n1047 185
R1410 GNDA.n1050 GNDA.n1049 185
R1411 GNDA.n1052 GNDA.n1051 185
R1412 GNDA.n1054 GNDA.n1053 185
R1413 GNDA.n1056 GNDA.n1055 185
R1414 GNDA.n1058 GNDA.n1057 185
R1415 GNDA.n1060 GNDA.n1059 185
R1416 GNDA.n1062 GNDA.n1061 185
R1417 GNDA.n1027 GNDA.n1024 185
R1418 GNDA.n1130 GNDA.n1129 185
R1419 GNDA.n1103 GNDA.n1026 185
R1420 GNDA.n1109 GNDA.n1108 185
R1421 GNDA.n1107 GNDA.n1102 185
R1422 GNDA.n1116 GNDA.n1115 185
R1423 GNDA.n1114 GNDA.n1101 185
R1424 GNDA.n1121 GNDA.n1046 185
R1425 GNDA.n1126 GNDA.n1125 185
R1426 GNDA.n418 GNDA.n407 185
R1427 GNDA.n411 GNDA.n407 185
R1428 GNDA.n418 GNDA.n417 185
R1429 GNDA.n417 GNDA.n416 185
R1430 GNDA.n1722 GNDA.n934 183.948
R1431 GNDA.n1655 GNDA.n1654 183.948
R1432 GNDA.t322 GNDA.t295 182.07
R1433 GNDA.t234 GNDA.t104 182.07
R1434 GNDA.t300 GNDA.t88 182.07
R1435 GNDA.t175 GNDA.t286 182.07
R1436 GNDA.n1679 GNDA.n934 180.013
R1437 GNDA.n1654 GNDA.n1653 180.013
R1438 GNDA.n922 GNDA.n921 175.546
R1439 GNDA.n1756 GNDA.n921 175.546
R1440 GNDA.n1754 GNDA.n1753 175.546
R1441 GNDA.n1750 GNDA.n1749 175.546
R1442 GNDA.n1746 GNDA.n1745 175.546
R1443 GNDA.n1765 GNDA.n653 175.546
R1444 GNDA.n1741 GNDA.n923 175.546
R1445 GNDA.n1741 GNDA.n925 175.546
R1446 GNDA.n1737 GNDA.n925 175.546
R1447 GNDA.n1737 GNDA.n927 175.546
R1448 GNDA.n1733 GNDA.n927 175.546
R1449 GNDA.n1733 GNDA.n929 175.546
R1450 GNDA.n1729 GNDA.n929 175.546
R1451 GNDA.n1729 GNDA.n931 175.546
R1452 GNDA.n1725 GNDA.n931 175.546
R1453 GNDA.n1725 GNDA.n933 175.546
R1454 GNDA.n1721 GNDA.n933 175.546
R1455 GNDA.n1768 GNDA.n650 175.546
R1456 GNDA.n1870 GNDA.n1869 175.546
R1457 GNDA.n1796 GNDA.n1795 175.546
R1458 GNDA.n1801 GNDA.n1800 175.546
R1459 GNDA.n1809 GNDA.n1808 175.546
R1460 GNDA.n1682 GNDA.n935 175.546
R1461 GNDA.n1683 GNDA.n1682 175.546
R1462 GNDA.n1686 GNDA.n1683 175.546
R1463 GNDA.n1687 GNDA.n1686 175.546
R1464 GNDA.n1690 GNDA.n1687 175.546
R1465 GNDA.n1691 GNDA.n1690 175.546
R1466 GNDA.n1692 GNDA.n1691 175.546
R1467 GNDA.n1693 GNDA.n1692 175.546
R1468 GNDA.n1697 GNDA.n1693 175.546
R1469 GNDA.n1697 GNDA.n516 175.546
R1470 GNDA.n1887 GNDA.n516 175.546
R1471 GNDA.n1325 GNDA.n1324 175.546
R1472 GNDA.n1329 GNDA.n1328 175.546
R1473 GNDA.n1333 GNDA.n1332 175.546
R1474 GNDA.n1337 GNDA.n1336 175.546
R1475 GNDA.n1341 GNDA.n1340 175.546
R1476 GNDA.n1317 GNDA.n1316 175.546
R1477 GNDA.n1313 GNDA.n1312 175.546
R1478 GNDA.n1309 GNDA.n1308 175.546
R1479 GNDA.n1305 GNDA.n1304 175.546
R1480 GNDA.n1301 GNDA.n453 175.546
R1481 GNDA.n1346 GNDA.n1300 175.546
R1482 GNDA.n1450 GNDA.n1449 175.546
R1483 GNDA.n1376 GNDA.n1375 175.546
R1484 GNDA.n1381 GNDA.n1380 175.546
R1485 GNDA.n1389 GNDA.n1388 175.546
R1486 GNDA.n475 GNDA.n466 175.546
R1487 GNDA.n468 GNDA.n467 175.546
R1488 GNDA.n470 GNDA.n469 175.546
R1489 GNDA.n472 GNDA.n471 175.546
R1490 GNDA.n474 GNDA.n473 175.546
R1491 GNDA.n915 GNDA.n671 175.546
R1492 GNDA.n913 GNDA.n912 175.546
R1493 GNDA.n909 GNDA.n908 175.546
R1494 GNDA.n905 GNDA.n904 175.546
R1495 GNDA.n901 GNDA.n900 175.546
R1496 GNDA.n766 GNDA.n765 175.546
R1497 GNDA.n763 GNDA.n675 175.546
R1498 GNDA.n759 GNDA.n758 175.546
R1499 GNDA.n756 GNDA.n678 175.546
R1500 GNDA.n752 GNDA.n751 175.546
R1501 GNDA.n896 GNDA.n771 175.546
R1502 GNDA.n892 GNDA.n771 175.546
R1503 GNDA.n892 GNDA.n772 175.546
R1504 GNDA.n806 GNDA.n772 175.546
R1505 GNDA.n810 GNDA.n806 175.546
R1506 GNDA.n810 GNDA.n801 175.546
R1507 GNDA.n823 GNDA.n801 175.546
R1508 GNDA.n823 GNDA.n799 175.546
R1509 GNDA.n827 GNDA.n799 175.546
R1510 GNDA.n830 GNDA.n827 175.546
R1511 GNDA.n830 GNDA.n88 175.546
R1512 GNDA.n715 GNDA.n714 175.546
R1513 GNDA.n720 GNDA.n717 175.546
R1514 GNDA.n723 GNDA.n722 175.546
R1515 GNDA.n727 GNDA.n725 175.546
R1516 GNDA.n2161 GNDA.n91 175.546
R1517 GNDA.n743 GNDA.n742 175.546
R1518 GNDA.n739 GNDA.n738 175.546
R1519 GNDA.n736 GNDA.n719 175.546
R1520 GNDA.n732 GNDA.n730 175.546
R1521 GNDA.n2159 GNDA.n93 175.546
R1522 GNDA.n709 GNDA.n684 175.546
R1523 GNDA.n705 GNDA.n704 175.546
R1524 GNDA.n702 GNDA.n687 175.546
R1525 GNDA.n698 GNDA.n697 175.546
R1526 GNDA.n695 GNDA.n691 175.546
R1527 GNDA.n2155 GNDA.n94 175.546
R1528 GNDA.n388 GNDA.n94 175.546
R1529 GNDA.n388 GNDA.n374 175.546
R1530 GNDA.n384 GNDA.n374 175.546
R1531 GNDA.n384 GNDA.n282 175.546
R1532 GNDA.n397 GNDA.n282 175.546
R1533 GNDA.n397 GNDA.n283 175.546
R1534 GNDA.n309 GNDA.n283 175.546
R1535 GNDA.n313 GNDA.n309 175.546
R1536 GNDA.n313 GNDA.n98 175.546
R1537 GNDA.n2149 GNDA.n98 175.546
R1538 GNDA.n2115 GNDA.n2113 175.546
R1539 GNDA.n2123 GNDA.n109 175.546
R1540 GNDA.n2127 GNDA.n2125 175.546
R1541 GNDA.n2135 GNDA.n105 175.546
R1542 GNDA.n2140 GNDA.n2137 175.546
R1543 GNDA.n1969 GNDA.n460 175.546
R1544 GNDA.n1965 GNDA.n465 175.546
R1545 GNDA.n1963 GNDA.n1962 175.546
R1546 GNDA.n1959 GNDA.n1958 175.546
R1547 GNDA.n1955 GNDA.n1954 175.546
R1548 GNDA.n1895 GNDA.n1894 175.546
R1549 GNDA.n1899 GNDA.n1898 175.546
R1550 GNDA.n1903 GNDA.n1902 175.546
R1551 GNDA.n1907 GNDA.n1906 175.546
R1552 GNDA.n1911 GNDA.n1910 175.546
R1553 GNDA.n1293 GNDA.n1181 175.546
R1554 GNDA.n1286 GNDA.n1285 175.546
R1555 GNDA.n1211 GNDA.n1210 175.546
R1556 GNDA.n1216 GNDA.n1215 175.546
R1557 GNDA.n1224 GNDA.n1223 175.546
R1558 GNDA.n1925 GNDA.n506 175.546
R1559 GNDA.n1928 GNDA.n1927 175.546
R1560 GNDA.n1930 GNDA.n504 175.546
R1561 GNDA.n1939 GNDA.n495 175.546
R1562 GNDA.n1942 GNDA.n1941 175.546
R1563 GNDA.n1717 GNDA.n1681 175.546
R1564 GNDA.n1713 GNDA.n1681 175.546
R1565 GNDA.n1713 GNDA.n1685 175.546
R1566 GNDA.n1709 GNDA.n1685 175.546
R1567 GNDA.n1709 GNDA.n1707 175.546
R1568 GNDA.n1707 GNDA.n1706 175.546
R1569 GNDA.n1706 GNDA.n1689 175.546
R1570 GNDA.n1702 GNDA.n1689 175.546
R1571 GNDA.n1702 GNDA.n1695 175.546
R1572 GNDA.n1698 GNDA.n1695 175.546
R1573 GNDA.n1698 GNDA.n518 175.546
R1574 GNDA.n1680 GNDA.n938 175.546
R1575 GNDA.n1676 GNDA.n938 175.546
R1576 GNDA.n1676 GNDA.n940 175.546
R1577 GNDA.n1672 GNDA.n940 175.546
R1578 GNDA.n1672 GNDA.n943 175.546
R1579 GNDA.n1665 GNDA.n943 175.546
R1580 GNDA.n1665 GNDA.n1664 175.546
R1581 GNDA.n1664 GNDA.n952 175.546
R1582 GNDA.n1660 GNDA.n952 175.546
R1583 GNDA.n1660 GNDA.n954 175.546
R1584 GNDA.n1656 GNDA.n954 175.546
R1585 GNDA.n643 GNDA.n521 175.546
R1586 GNDA.n560 GNDA.n532 175.546
R1587 GNDA.n566 GNDA.n565 175.546
R1588 GNDA.n573 GNDA.n572 175.546
R1589 GNDA.n581 GNDA.n580 175.546
R1590 GNDA.n961 GNDA.n957 175.546
R1591 GNDA.n962 GNDA.n961 175.546
R1592 GNDA.n966 GNDA.n962 175.546
R1593 GNDA.n967 GNDA.n966 175.546
R1594 GNDA.n969 GNDA.n967 175.546
R1595 GNDA.n970 GNDA.n969 175.546
R1596 GNDA.n973 GNDA.n970 175.546
R1597 GNDA.n974 GNDA.n973 175.546
R1598 GNDA.n975 GNDA.n974 175.546
R1599 GNDA.n979 GNDA.n975 175.546
R1600 GNDA.n980 GNDA.n979 175.546
R1601 GNDA.n1923 GNDA.n1920 175.546
R1602 GNDA.n1923 GNDA.n1922 175.546
R1603 GNDA.n1932 GNDA.n501 175.546
R1604 GNDA.n1935 GNDA.n1934 175.546
R1605 GNDA.n1937 GNDA.n499 175.546
R1606 GNDA.n497 GNDA.n489 175.546
R1607 GNDA.n1145 GNDA.n1144 175.546
R1608 GNDA.n1149 GNDA.n1148 175.546
R1609 GNDA.n1153 GNDA.n1152 175.546
R1610 GNDA.n1157 GNDA.n1156 175.546
R1611 GNDA.n1161 GNDA.n1160 175.546
R1612 GNDA.n1548 GNDA.n1475 175.546
R1613 GNDA.n1552 GNDA.n1550 175.546
R1614 GNDA.n1563 GNDA.n1469 175.546
R1615 GNDA.n1567 GNDA.n1565 175.546
R1616 GNDA.n1578 GNDA.n1462 175.546
R1617 GNDA.n1603 GNDA.n1142 175.546
R1618 GNDA.n1599 GNDA.n1142 175.546
R1619 GNDA.n1599 GNDA.n1165 175.546
R1620 GNDA.n1595 GNDA.n1165 175.546
R1621 GNDA.n1595 GNDA.n1166 175.546
R1622 GNDA.n1591 GNDA.n1166 175.546
R1623 GNDA.n1591 GNDA.n1590 175.546
R1624 GNDA.n1590 GNDA.n1168 175.546
R1625 GNDA.n1586 GNDA.n1168 175.546
R1626 GNDA.n1586 GNDA.n1170 175.546
R1627 GNDA.n1174 GNDA.n1170 175.546
R1628 GNDA.n2117 GNDA.n111 175.546
R1629 GNDA.n2121 GNDA.n2119 175.546
R1630 GNDA.n2129 GNDA.n107 175.546
R1631 GNDA.n2133 GNDA.n2131 175.546
R1632 GNDA.n2142 GNDA.n103 175.546
R1633 GNDA.n2105 GNDA.n116 175.546
R1634 GNDA.n2101 GNDA.n2100 175.546
R1635 GNDA.n2098 GNDA.n119 175.546
R1636 GNDA.n2094 GNDA.n2093 175.546
R1637 GNDA.n2091 GNDA.n122 175.546
R1638 GNDA.n2194 GNDA.n76 175.546
R1639 GNDA.n2209 GNDA.n2194 175.546
R1640 GNDA.n2209 GNDA.n2195 175.546
R1641 GNDA.n2205 GNDA.n2195 175.546
R1642 GNDA.n2205 GNDA.n51 175.546
R1643 GNDA.n2218 GNDA.n51 175.546
R1644 GNDA.n2218 GNDA.n52 175.546
R1645 GNDA.n2056 GNDA.n52 175.546
R1646 GNDA.n2056 GNDA.n1991 175.546
R1647 GNDA.n2060 GNDA.n1991 175.546
R1648 GNDA.n2061 GNDA.n2060 175.546
R1649 GNDA.n2086 GNDA.n125 175.546
R1650 GNDA.n2082 GNDA.n125 175.546
R1651 GNDA.n2082 GNDA.n1981 175.546
R1652 GNDA.n2078 GNDA.n1981 175.546
R1653 GNDA.n2078 GNDA.n2076 175.546
R1654 GNDA.n2076 GNDA.n2075 175.546
R1655 GNDA.n2075 GNDA.n1984 175.546
R1656 GNDA.n2071 GNDA.n1984 175.546
R1657 GNDA.n2071 GNDA.n1986 175.546
R1658 GNDA.n2067 GNDA.n1986 175.546
R1659 GNDA.n2067 GNDA.n1989 175.546
R1660 GNDA.n1001 GNDA.n960 175.546
R1661 GNDA.n997 GNDA.n960 175.546
R1662 GNDA.n997 GNDA.n964 175.546
R1663 GNDA.n993 GNDA.n964 175.546
R1664 GNDA.n993 GNDA.n968 175.546
R1665 GNDA.n989 GNDA.n968 175.546
R1666 GNDA.n989 GNDA.n988 175.546
R1667 GNDA.n988 GNDA.n972 175.546
R1668 GNDA.n984 GNDA.n972 175.546
R1669 GNDA.n984 GNDA.n977 175.546
R1670 GNDA.n977 GNDA.n512 175.546
R1671 GNDA.n1652 GNDA.n1002 175.546
R1672 GNDA.n1648 GNDA.n1002 175.546
R1673 GNDA.n1648 GNDA.n1004 175.546
R1674 GNDA.n1644 GNDA.n1004 175.546
R1675 GNDA.n1644 GNDA.n1006 175.546
R1676 GNDA.n1640 GNDA.n1006 175.546
R1677 GNDA.n1640 GNDA.n1008 175.546
R1678 GNDA.n1636 GNDA.n1008 175.546
R1679 GNDA.n1636 GNDA.n1010 175.546
R1680 GNDA.n1632 GNDA.n1010 175.546
R1681 GNDA.n1632 GNDA.n1012 175.546
R1682 GNDA.n1123 GNDA.n1122 175.546
R1683 GNDA.n1119 GNDA.n1118 175.546
R1684 GNDA.n1112 GNDA.n1111 175.546
R1685 GNDA.n1105 GNDA.n1104 175.546
R1686 GNDA.n1133 GNDA.n1132 175.546
R1687 GNDA.n1628 GNDA.n1014 175.546
R1688 GNDA.n1624 GNDA.n1014 175.546
R1689 GNDA.n1624 GNDA.n1016 175.546
R1690 GNDA.n1620 GNDA.n1016 175.546
R1691 GNDA.n1620 GNDA.n1017 175.546
R1692 GNDA.n1616 GNDA.n1017 175.546
R1693 GNDA.n1616 GNDA.n1615 175.546
R1694 GNDA.n1615 GNDA.n1019 175.546
R1695 GNDA.n1611 GNDA.n1019 175.546
R1696 GNDA.n1611 GNDA.n1021 175.546
R1697 GNDA.n1137 GNDA.n1021 175.546
R1698 GNDA.n481 GNDA.n126 173.881
R1699 GNDA.t227 GNDA.n127 172.876
R1700 GNDA.t227 GNDA.n435 172.615
R1701 GNDA.n1971 GNDA.n126 171.624
R1702 GNDA.n196 GNDA.t94 166.898
R1703 GNDA.n1813 GNDA.n1812 163.333
R1704 GNDA.n1393 GNDA.n1392 163.333
R1705 GNDA.n834 GNDA.n833 163.333
R1706 GNDA.n318 GNDA.n317 163.333
R1707 GNDA.n1228 GNDA.n1227 163.333
R1708 GNDA.n585 GNDA.n584 163.333
R1709 GNDA.n1574 GNDA.n1573 163.333
R1710 GNDA.n2050 GNDA.n2049 163.333
R1711 GNDA.n1037 GNDA.n1027 163.333
R1712 GNDA.t48 GNDA.t339 162.662
R1713 GNDA.n205 GNDA.n204 161.3
R1714 GNDA.n193 GNDA.n192 161.3
R1715 GNDA.t295 GNDA.t176 151.725
R1716 GNDA.t104 GNDA.t322 151.725
R1717 GNDA.t92 GNDA.t234 151.725
R1718 GNDA.n197 GNDA.t179 151.725
R1719 GNDA.t14 GNDA.t300 151.725
R1720 GNDA.t88 GNDA.t175 151.725
R1721 GNDA.t286 GNDA.t124 151.725
R1722 GNDA.n1845 GNDA.n1844 150
R1723 GNDA.n1841 GNDA.n1840 150
R1724 GNDA.n1837 GNDA.n1836 150
R1725 GNDA.n1833 GNDA.n1832 150
R1726 GNDA.n1829 GNDA.n1828 150
R1727 GNDA.n1825 GNDA.n1824 150
R1728 GNDA.n1821 GNDA.n1820 150
R1729 GNDA.n1817 GNDA.n1816 150
R1730 GNDA.n1874 GNDA.n1873 150
R1731 GNDA.n1866 GNDA.n1774 150
R1732 GNDA.n1798 GNDA.n1775 150
R1733 GNDA.n1805 GNDA.n1804 150
R1734 GNDA.n1863 GNDA.n1791 150
R1735 GNDA.n1859 GNDA.n1858 150
R1736 GNDA.n1855 GNDA.n1854 150
R1737 GNDA.n1851 GNDA.n1850 150
R1738 GNDA.n1425 GNDA.n1424 150
R1739 GNDA.n1421 GNDA.n1420 150
R1740 GNDA.n1417 GNDA.n1416 150
R1741 GNDA.n1413 GNDA.n1412 150
R1742 GNDA.n1409 GNDA.n1408 150
R1743 GNDA.n1405 GNDA.n1404 150
R1744 GNDA.n1401 GNDA.n1400 150
R1745 GNDA.n1397 GNDA.n1396 150
R1746 GNDA.n1454 GNDA.n1453 150
R1747 GNDA.n1446 GNDA.n1352 150
R1748 GNDA.n1378 GNDA.n1353 150
R1749 GNDA.n1385 GNDA.n1384 150
R1750 GNDA.n1443 GNDA.n1369 150
R1751 GNDA.n1439 GNDA.n1438 150
R1752 GNDA.n1435 GNDA.n1434 150
R1753 GNDA.n1431 GNDA.n1430 150
R1754 GNDA.n866 GNDA.n865 150
R1755 GNDA.n862 GNDA.n861 150
R1756 GNDA.n858 GNDA.n857 150
R1757 GNDA.n854 GNDA.n853 150
R1758 GNDA.n850 GNDA.n849 150
R1759 GNDA.n846 GNDA.n845 150
R1760 GNDA.n842 GNDA.n841 150
R1761 GNDA.n838 GNDA.n837 150
R1762 GNDA.n889 GNDA.n776 150
R1763 GNDA.n802 GNDA.n777 150
R1764 GNDA.n815 GNDA.n814 150
R1765 GNDA.n820 GNDA.n819 150
R1766 GNDA.n874 GNDA.n873 150
R1767 GNDA.n878 GNDA.n877 150
R1768 GNDA.n882 GNDA.n881 150
R1769 GNDA.n886 GNDA.n794 150
R1770 GNDA.n350 GNDA.n349 150
R1771 GNDA.n346 GNDA.n345 150
R1772 GNDA.n342 GNDA.n341 150
R1773 GNDA.n338 GNDA.n337 150
R1774 GNDA.n334 GNDA.n333 150
R1775 GNDA.n330 GNDA.n329 150
R1776 GNDA.n326 GNDA.n325 150
R1777 GNDA.n322 GNDA.n321 150
R1778 GNDA.n391 GNDA.n304 150
R1779 GNDA.n381 GNDA.n380 150
R1780 GNDA.n394 GNDA.n285 150
R1781 GNDA.n305 GNDA.n286 150
R1782 GNDA.n358 GNDA.n357 150
R1783 GNDA.n362 GNDA.n361 150
R1784 GNDA.n366 GNDA.n365 150
R1785 GNDA.n368 GNDA.n303 150
R1786 GNDA.n1260 GNDA.n1259 150
R1787 GNDA.n1256 GNDA.n1255 150
R1788 GNDA.n1252 GNDA.n1251 150
R1789 GNDA.n1248 GNDA.n1247 150
R1790 GNDA.n1244 GNDA.n1243 150
R1791 GNDA.n1240 GNDA.n1239 150
R1792 GNDA.n1236 GNDA.n1235 150
R1793 GNDA.n1232 GNDA.n1231 150
R1794 GNDA.n1290 GNDA.n1289 150
R1795 GNDA.n1282 GNDA.n1189 150
R1796 GNDA.n1213 GNDA.n1190 150
R1797 GNDA.n1220 GNDA.n1219 150
R1798 GNDA.n1279 GNDA.n1206 150
R1799 GNDA.n1275 GNDA.n1274 150
R1800 GNDA.n1271 GNDA.n1270 150
R1801 GNDA.n1267 GNDA.n1266 150
R1802 GNDA.n617 GNDA.n616 150
R1803 GNDA.n613 GNDA.n612 150
R1804 GNDA.n609 GNDA.n608 150
R1805 GNDA.n605 GNDA.n604 150
R1806 GNDA.n601 GNDA.n600 150
R1807 GNDA.n597 GNDA.n596 150
R1808 GNDA.n593 GNDA.n592 150
R1809 GNDA.n589 GNDA.n588 150
R1810 GNDA.n640 GNDA.n536 150
R1811 GNDA.n562 GNDA.n537 150
R1812 GNDA.n570 GNDA.n569 150
R1813 GNDA.n577 GNDA.n576 150
R1814 GNDA.n625 GNDA.n624 150
R1815 GNDA.n629 GNDA.n628 150
R1816 GNDA.n633 GNDA.n632 150
R1817 GNDA.n637 GNDA.n554 150
R1818 GNDA.n1519 GNDA.n1517 150
R1819 GNDA.n1515 GNDA.n1483 150
R1820 GNDA.n1511 GNDA.n1509 150
R1821 GNDA.n1507 GNDA.n1485 150
R1822 GNDA.n1503 GNDA.n1501 150
R1823 GNDA.n1499 GNDA.n1487 150
R1824 GNDA.n1495 GNDA.n1494 150
R1825 GNDA.n1492 GNDA.n1490 150
R1826 GNDA.n1545 GNDA.n1543 150
R1827 GNDA.n1556 GNDA.n1471 150
R1828 GNDA.n1560 GNDA.n1558 150
R1829 GNDA.n1571 GNDA.n1466 150
R1830 GNDA.n1527 GNDA.n1525 150
R1831 GNDA.n1531 GNDA.n1479 150
R1832 GNDA.n1535 GNDA.n1533 150
R1833 GNDA.n1541 GNDA.n1477 150
R1834 GNDA.n2017 GNDA.n2016 150
R1835 GNDA.n2021 GNDA.n2020 150
R1836 GNDA.n2025 GNDA.n2024 150
R1837 GNDA.n2029 GNDA.n2028 150
R1838 GNDA.n2033 GNDA.n2032 150
R1839 GNDA.n2037 GNDA.n2036 150
R1840 GNDA.n2041 GNDA.n2040 150
R1841 GNDA.n2045 GNDA.n2044 150
R1842 GNDA.n2212 GNDA.n73 150
R1843 GNDA.n2202 GNDA.n2201 150
R1844 GNDA.n2215 GNDA.n54 150
R1845 GNDA.n2053 GNDA.n55 150
R1846 GNDA.n2009 GNDA.n2008 150
R1847 GNDA.n2005 GNDA.n2004 150
R1848 GNDA.n2001 GNDA.n2000 150
R1849 GNDA.n1997 GNDA.n72 150
R1850 GNDA.n1077 GNDA.n1076 150
R1851 GNDA.n1073 GNDA.n1072 150
R1852 GNDA.n1069 GNDA.n1068 150
R1853 GNDA.n1065 GNDA.n1064 150
R1854 GNDA.n1061 GNDA.n1060 150
R1855 GNDA.n1057 GNDA.n1056 150
R1856 GNDA.n1053 GNDA.n1052 150
R1857 GNDA.n1049 GNDA.n1048 150
R1858 GNDA.n1126 GNDA.n1046 150
R1859 GNDA.n1115 GNDA.n1114 150
R1860 GNDA.n1108 GNDA.n1107 150
R1861 GNDA.n1129 GNDA.n1026 150
R1862 GNDA.n1085 GNDA.n1084 150
R1863 GNDA.n1089 GNDA.n1088 150
R1864 GNDA.n1093 GNDA.n1092 150
R1865 GNDA.n1095 GNDA.n1045 150
R1866 GNDA.n185 GNDA.n184 148.017
R1867 GNDA.n171 GNDA.n170 148.017
R1868 GNDA.n2252 GNDA.n2251 148.017
R1869 GNDA.n2247 GNDA.n2246 148.017
R1870 GNDA.t126 GNDA.t150 147.84
R1871 GNDA.t335 GNDA.t325 144.321
R1872 GNDA.n131 GNDA.n130 139.077
R1873 GNDA.n129 GNDA.n128 139.077
R1874 GNDA.n87 GNDA.n86 139.077
R1875 GNDA.n2175 GNDA.n2174 139.077
R1876 GNDA.n2173 GNDA.n2172 139.077
R1877 GNDA.n2171 GNDA.n2170 139.077
R1878 GNDA.n79 GNDA.n78 139.077
R1879 GNDA.n2187 GNDA.n2186 139.077
R1880 GNDA.n2185 GNDA.n2184 139.077
R1881 GNDA.n39 GNDA.n38 139.077
R1882 GNDA.t167 GNDA.t53 139.041
R1883 GNDA.n2236 GNDA.t157 135.69
R1884 GNDA.n409 GNDA.n407 134.268
R1885 GNDA.n417 GNDA.n409 134.268
R1886 GNDA.n1343 GNDA.n663 132.721
R1887 GNDA.n769 GNDA.n666 132.721
R1888 GNDA.n2241 GNDA.t259 130.001
R1889 GNDA.n2190 GNDA.t265 130.001
R1890 GNDA.n2181 GNDA.t256 130.001
R1891 GNDA.n2178 GNDA.t311 130.001
R1892 GNDA.n2167 GNDA.t281 130.001
R1893 GNDA.n133 GNDA.t269 130.001
R1894 GNDA.n1888 GNDA.n1887 124.832
R1895 GNDA.n487 GNDA.n483 124.832
R1896 GNDA.n2164 GNDA.n2163 124.832
R1897 GNDA.n2157 GNDA.n2156 124.832
R1898 GNDA.n2138 GNDA.n99 124.832
R1899 GNDA.n1951 GNDA.n1950 124.832
R1900 GNDA.n1944 GNDA.n488 124.832
R1901 GNDA.n518 GNDA.n514 124.832
R1902 GNDA.n980 GNDA.n511 124.832
R1903 GNDA.n1948 GNDA.n489 124.832
R1904 GNDA.n2145 GNDA.n2144 124.832
R1905 GNDA.n1890 GNDA.n512 124.832
R1906 GNDA.n18 GNDA.n16 124.59
R1907 GNDA.n161 GNDA.n159 124.59
R1908 GNDA.n26 GNDA.n25 124.028
R1909 GNDA.n24 GNDA.n23 124.028
R1910 GNDA.n22 GNDA.n21 124.028
R1911 GNDA.n20 GNDA.n19 124.028
R1912 GNDA.n18 GNDA.n17 124.028
R1913 GNDA.n169 GNDA.n168 124.028
R1914 GNDA.n167 GNDA.n166 124.028
R1915 GNDA.n165 GNDA.n164 124.028
R1916 GNDA.n163 GNDA.n162 124.028
R1917 GNDA.n161 GNDA.n160 124.028
R1918 GNDA.n41 GNDA.t54 115.948
R1919 GNDA.n947 GNDA.t148 115.105
R1920 GNDA.n41 GNDA.t326 114.635
R1921 GNDA.n948 GNDA.t332 114.635
R1922 GNDA.n2245 GNDA.t136 111.954
R1923 GNDA.t303 GNDA.n149 109.797
R1924 GNDA.n2253 GNDA.t313 109.797
R1925 GNDA.t255 GNDA.n80 101.942
R1926 GNDA.n2220 GNDA.n47 101.718
R1927 GNDA.n2231 GNDA.n46 101.718
R1928 GNDA.n406 GNDA.n404 101.718
R1929 GNDA.n413 GNDA.n405 101.718
R1930 GNDA.n412 GNDA.n404 101.718
R1931 GNDA.t227 GNDA.n82 47.6748
R1932 GNDA.n2154 GNDA.n85 98.8538
R1933 GNDA.t20 GNDA.t127 97.5975
R1934 GNDA.t338 GNDA.t20 97.5975
R1935 GNDA.t339 GNDA.t338 97.5975
R1936 GNDA.t153 GNDA.t48 97.5975
R1937 GNDA.n2193 GNDA.n2192 92.6754
R1938 GNDA.n2227 GNDA.n45 91.069
R1939 GNDA.n2222 GNDA.n45 91.069
R1940 GNDA.n2224 GNDA.n44 91.069
R1941 GNDA.n2225 GNDA.n2224 91.069
R1942 GNDA.n415 GNDA.n407 91.069
R1943 GNDA.n417 GNDA.n410 91.069
R1944 GNDA.t280 GNDA.n828 90.616
R1945 GNDA.n2085 GNDA.t227 90.5399
R1946 GNDA.t337 GNDA.t165 89.4645
R1947 GNDA.t147 GNDA.t13 89.4645
R1948 GNDA.t329 GNDA.t323 89.4645
R1949 GNDA.t125 GNDA.t340 89.4645
R1950 GNDA.t116 GNDA.t137 89.4645
R1951 GNDA.t31 GNDA.t171 89.4645
R1952 GNDA.t171 GNDA.t96 89.4645
R1953 GNDA.t33 GNDA.t173 89.4645
R1954 GNDA.t115 GNDA.t63 89.4645
R1955 GNDA.t28 GNDA.t43 89.4645
R1956 GNDA.t41 GNDA.t158 89.4645
R1957 GNDA.t4 GNDA.t64 89.4645
R1958 GNDA.t112 GNDA.t110 89.4645
R1959 GNDA.n1740 GNDA.n423 88.5317
R1960 GNDA.n1740 GNDA.n1739 88.5317
R1961 GNDA.n1739 GNDA.n1738 88.5317
R1962 GNDA.n1738 GNDA.n926 88.5317
R1963 GNDA.n1732 GNDA.n926 88.5317
R1964 GNDA.n1731 GNDA.n1730 88.5317
R1965 GNDA.n1730 GNDA.n930 88.5317
R1966 GNDA.n1724 GNDA.n930 88.5317
R1967 GNDA.n1724 GNDA.n1723 88.5317
R1968 GNDA.n1723 GNDA.n1722 88.5317
R1969 GNDA.n1679 GNDA.n1678 88.5317
R1970 GNDA.n1678 GNDA.n1677 88.5317
R1971 GNDA.n1677 GNDA.n939 88.5317
R1972 GNDA.n1671 GNDA.n939 88.5317
R1973 GNDA.n1671 GNDA.n1670 88.5317
R1974 GNDA.n1663 GNDA.n945 88.5317
R1975 GNDA.n1663 GNDA.n1662 88.5317
R1976 GNDA.n1662 GNDA.n1661 88.5317
R1977 GNDA.n1661 GNDA.n953 88.5317
R1978 GNDA.n1655 GNDA.n953 88.5317
R1979 GNDA.n1653 GNDA.n959 88.5317
R1980 GNDA.n1647 GNDA.n959 88.5317
R1981 GNDA.n1647 GNDA.n1646 88.5317
R1982 GNDA.n1646 GNDA.n1645 88.5317
R1983 GNDA.n1645 GNDA.n1005 88.5317
R1984 GNDA.n1639 GNDA.n1638 88.5317
R1985 GNDA.n1638 GNDA.n1637 88.5317
R1986 GNDA.n1637 GNDA.n1009 88.5317
R1987 GNDA.n1631 GNDA.n1009 88.5317
R1988 GNDA.n1631 GNDA.n1630 88.5317
R1989 GNDA.t37 GNDA.n2243 85.4674
R1990 GNDA.t261 GNDA.t289 85.3979
R1991 GNDA.t277 GNDA.t283 85.3979
R1992 GNDA.n2260 GNDA.t35 85.3979
R1993 GNDA.t249 GNDA.t224 85.3979
R1994 GNDA.t244 GNDA.t241 85.3979
R1995 GNDA.n385 GNDA.t201 84.4377
R1996 GNDA.n946 GNDA.n944 84.306
R1997 GNDA.t87 GNDA.t128 83.3141
R1998 GNDA.t23 GNDA.t131 82.3782
R1999 GNDA.t144 GNDA.t156 82.3782
R2000 GNDA.t16 GNDA.n1604 81.9681
R2001 GNDA.n1654 GNDA.n958 80.9821
R2002 GNDA.n1716 GNDA.n934 80.9821
R2003 GNDA.n310 GNDA.t193 80.3188
R2004 GNDA.t227 GNDA.n126 76.3879
R2005 GNDA.n1762 GNDA.n1761 76.3222
R2006 GNDA.n1756 GNDA.n654 76.3222
R2007 GNDA.n1753 GNDA.n655 76.3222
R2008 GNDA.n1749 GNDA.n656 76.3222
R2009 GNDA.n1745 GNDA.n657 76.3222
R2010 GNDA.n1880 GNDA.n1879 76.3222
R2011 GNDA.n1768 GNDA.n649 76.3222
R2012 GNDA.n1869 GNDA.n648 76.3222
R2013 GNDA.n1796 GNDA.n647 76.3222
R2014 GNDA.n1800 GNDA.n646 76.3222
R2015 GNDA.n1809 GNDA.n645 76.3222
R2016 GNDA.n1321 GNDA.n658 76.3222
R2017 GNDA.n1325 GNDA.n659 76.3222
R2018 GNDA.n1329 GNDA.n660 76.3222
R2019 GNDA.n1333 GNDA.n661 76.3222
R2020 GNDA.n1337 GNDA.n662 76.3222
R2021 GNDA.n1341 GNDA.n663 76.3222
R2022 GNDA.n1317 GNDA.n448 76.3222
R2023 GNDA.n1313 GNDA.n449 76.3222
R2024 GNDA.n1309 GNDA.n450 76.3222
R2025 GNDA.n1305 GNDA.n451 76.3222
R2026 GNDA.n1301 GNDA.n452 76.3222
R2027 GNDA.n1978 GNDA.n1977 76.3222
R2028 GNDA.n1460 GNDA.n1459 76.3222
R2029 GNDA.n1346 GNDA.n1299 76.3222
R2030 GNDA.n1449 GNDA.n1298 76.3222
R2031 GNDA.n1376 GNDA.n1297 76.3222
R2032 GNDA.n1380 GNDA.n1296 76.3222
R2033 GNDA.n1389 GNDA.n1295 76.3222
R2034 GNDA.n476 GNDA.n454 76.3222
R2035 GNDA.n477 GNDA.n466 76.3222
R2036 GNDA.n478 GNDA.n468 76.3222
R2037 GNDA.n479 GNDA.n470 76.3222
R2038 GNDA.n480 GNDA.n472 76.3222
R2039 GNDA.n482 GNDA.n474 76.3222
R2040 GNDA.n920 GNDA.n919 76.3222
R2041 GNDA.n915 GNDA.n670 76.3222
R2042 GNDA.n912 GNDA.n669 76.3222
R2043 GNDA.n908 GNDA.n668 76.3222
R2044 GNDA.n904 GNDA.n667 76.3222
R2045 GNDA.n900 GNDA.n666 76.3222
R2046 GNDA.n766 GNDA.n674 76.3222
R2047 GNDA.n764 GNDA.n763 76.3222
R2048 GNDA.n759 GNDA.n677 76.3222
R2049 GNDA.n757 GNDA.n756 76.3222
R2050 GNDA.n752 GNDA.n680 76.3222
R2051 GNDA.n750 GNDA.n749 76.3222
R2052 GNDA.n713 GNDA.n681 76.3222
R2053 GNDA.n716 GNDA.n715 76.3222
R2054 GNDA.n721 GNDA.n720 76.3222
R2055 GNDA.n724 GNDA.n723 76.3222
R2056 GNDA.n727 GNDA.n726 76.3222
R2057 GNDA.n2162 GNDA.n2161 76.3222
R2058 GNDA.n745 GNDA.n744 76.3222
R2059 GNDA.n742 GNDA.n712 76.3222
R2060 GNDA.n738 GNDA.n737 76.3222
R2061 GNDA.n731 GNDA.n719 76.3222
R2062 GNDA.n730 GNDA.n729 76.3222
R2063 GNDA.n2159 GNDA.n2158 76.3222
R2064 GNDA.n710 GNDA.n709 76.3222
R2065 GNDA.n705 GNDA.n686 76.3222
R2066 GNDA.n703 GNDA.n702 76.3222
R2067 GNDA.n698 GNDA.n689 76.3222
R2068 GNDA.n696 GNDA.n695 76.3222
R2069 GNDA.n690 GNDA.n113 76.3222
R2070 GNDA.n2112 GNDA.n2111 76.3222
R2071 GNDA.n2115 GNDA.n2114 76.3222
R2072 GNDA.n2124 GNDA.n2123 76.3222
R2073 GNDA.n2127 GNDA.n2126 76.3222
R2074 GNDA.n2136 GNDA.n2135 76.3222
R2075 GNDA.n2140 GNDA.n2139 76.3222
R2076 GNDA.n1973 GNDA.n1972 76.3222
R2077 GNDA.n1970 GNDA.n1969 76.3222
R2078 GNDA.n1965 GNDA.n464 76.3222
R2079 GNDA.n1962 GNDA.n463 76.3222
R2080 GNDA.n1958 GNDA.n462 76.3222
R2081 GNDA.n1954 GNDA.n461 76.3222
R2082 GNDA.n1894 GNDA.n442 76.3222
R2083 GNDA.n1898 GNDA.n443 76.3222
R2084 GNDA.n1902 GNDA.n444 76.3222
R2085 GNDA.n1906 GNDA.n445 76.3222
R2086 GNDA.n1910 GNDA.n446 76.3222
R2087 GNDA.n1914 GNDA.n447 76.3222
R2088 GNDA.n1294 GNDA.n485 76.3222
R2089 GNDA.n1181 GNDA.n1180 76.3222
R2090 GNDA.n1285 GNDA.n1179 76.3222
R2091 GNDA.n1211 GNDA.n1178 76.3222
R2092 GNDA.n1215 GNDA.n1177 76.3222
R2093 GNDA.n1224 GNDA.n1176 76.3222
R2094 GNDA.n1916 GNDA.n1915 76.3222
R2095 GNDA.n1926 GNDA.n1925 76.3222
R2096 GNDA.n1929 GNDA.n1928 76.3222
R2097 GNDA.n504 GNDA.n503 76.3222
R2098 GNDA.n1940 GNDA.n1939 76.3222
R2099 GNDA.n1943 GNDA.n1942 76.3222
R2100 GNDA.n1883 GNDA.n1882 76.3222
R2101 GNDA.n644 GNDA.n643 76.3222
R2102 GNDA.n560 GNDA.n531 76.3222
R2103 GNDA.n566 GNDA.n530 76.3222
R2104 GNDA.n572 GNDA.n529 76.3222
R2105 GNDA.n581 GNDA.n528 76.3222
R2106 GNDA.n1919 GNDA.n1918 76.3222
R2107 GNDA.n1922 GNDA.n1921 76.3222
R2108 GNDA.n1933 GNDA.n1932 76.3222
R2109 GNDA.n1936 GNDA.n1935 76.3222
R2110 GNDA.n499 GNDA.n498 76.3222
R2111 GNDA.n1144 GNDA.n436 76.3222
R2112 GNDA.n1148 GNDA.n437 76.3222
R2113 GNDA.n1152 GNDA.n438 76.3222
R2114 GNDA.n1156 GNDA.n439 76.3222
R2115 GNDA.n1160 GNDA.n440 76.3222
R2116 GNDA.n1141 GNDA.n441 76.3222
R2117 GNDA.n1474 GNDA.n490 76.3222
R2118 GNDA.n1549 GNDA.n1548 76.3222
R2119 GNDA.n1552 GNDA.n1551 76.3222
R2120 GNDA.n1564 GNDA.n1563 76.3222
R2121 GNDA.n1567 GNDA.n1566 76.3222
R2122 GNDA.n1579 GNDA.n1578 76.3222
R2123 GNDA.n2109 GNDA.n2108 76.3222
R2124 GNDA.n2118 GNDA.n2117 76.3222
R2125 GNDA.n2121 GNDA.n2120 76.3222
R2126 GNDA.n2130 GNDA.n2129 76.3222
R2127 GNDA.n2133 GNDA.n2132 76.3222
R2128 GNDA.n2143 GNDA.n2142 76.3222
R2129 GNDA.n2106 GNDA.n2105 76.3222
R2130 GNDA.n2101 GNDA.n118 76.3222
R2131 GNDA.n2099 GNDA.n2098 76.3222
R2132 GNDA.n2094 GNDA.n121 76.3222
R2133 GNDA.n2092 GNDA.n2091 76.3222
R2134 GNDA.n2087 GNDA.n124 76.3222
R2135 GNDA.n527 GNDA.n513 76.3222
R2136 GNDA.n1123 GNDA.n526 76.3222
R2137 GNDA.n1118 GNDA.n525 76.3222
R2138 GNDA.n1111 GNDA.n524 76.3222
R2139 GNDA.n1104 GNDA.n523 76.3222
R2140 GNDA.n1133 GNDA.n522 76.3222
R2141 GNDA.n1944 GNDA.n1943 76.3222
R2142 GNDA.n1941 GNDA.n1940 76.3222
R2143 GNDA.n503 GNDA.n495 76.3222
R2144 GNDA.n1930 GNDA.n1929 76.3222
R2145 GNDA.n1927 GNDA.n1926 76.3222
R2146 GNDA.n1915 GNDA.n506 76.3222
R2147 GNDA.n1920 GNDA.n1919 76.3222
R2148 GNDA.n1921 GNDA.n501 76.3222
R2149 GNDA.n1934 GNDA.n1933 76.3222
R2150 GNDA.n1937 GNDA.n1936 76.3222
R2151 GNDA.n498 GNDA.n497 76.3222
R2152 GNDA.n2139 GNDA.n2138 76.3222
R2153 GNDA.n2137 GNDA.n2136 76.3222
R2154 GNDA.n2126 GNDA.n105 76.3222
R2155 GNDA.n2125 GNDA.n2124 76.3222
R2156 GNDA.n2114 GNDA.n109 76.3222
R2157 GNDA.n2113 GNDA.n2112 76.3222
R2158 GNDA.n2108 GNDA.n111 76.3222
R2159 GNDA.n2119 GNDA.n2118 76.3222
R2160 GNDA.n2120 GNDA.n107 76.3222
R2161 GNDA.n2131 GNDA.n2130 76.3222
R2162 GNDA.n2132 GNDA.n103 76.3222
R2163 GNDA.n2144 GNDA.n2143 76.3222
R2164 GNDA.n2163 GNDA.n2162 76.3222
R2165 GNDA.n726 GNDA.n91 76.3222
R2166 GNDA.n725 GNDA.n724 76.3222
R2167 GNDA.n722 GNDA.n721 76.3222
R2168 GNDA.n717 GNDA.n716 76.3222
R2169 GNDA.n714 GNDA.n713 76.3222
R2170 GNDA.n744 GNDA.n743 76.3222
R2171 GNDA.n739 GNDA.n712 76.3222
R2172 GNDA.n737 GNDA.n736 76.3222
R2173 GNDA.n732 GNDA.n731 76.3222
R2174 GNDA.n729 GNDA.n93 76.3222
R2175 GNDA.n2158 GNDA.n2157 76.3222
R2176 GNDA.n483 GNDA.n482 76.3222
R2177 GNDA.n480 GNDA.n473 76.3222
R2178 GNDA.n479 GNDA.n471 76.3222
R2179 GNDA.n478 GNDA.n469 76.3222
R2180 GNDA.n477 GNDA.n467 76.3222
R2181 GNDA.n476 GNDA.n475 76.3222
R2182 GNDA.n1972 GNDA.n460 76.3222
R2183 GNDA.n1970 GNDA.n465 76.3222
R2184 GNDA.n1963 GNDA.n464 76.3222
R2185 GNDA.n1959 GNDA.n463 76.3222
R2186 GNDA.n1955 GNDA.n462 76.3222
R2187 GNDA.n1951 GNDA.n461 76.3222
R2188 GNDA.n1978 GNDA.n453 76.3222
R2189 GNDA.n1304 GNDA.n452 76.3222
R2190 GNDA.n1308 GNDA.n451 76.3222
R2191 GNDA.n1312 GNDA.n450 76.3222
R2192 GNDA.n1316 GNDA.n449 76.3222
R2193 GNDA.n1320 GNDA.n448 76.3222
R2194 GNDA.n1911 GNDA.n447 76.3222
R2195 GNDA.n1907 GNDA.n446 76.3222
R2196 GNDA.n1903 GNDA.n445 76.3222
R2197 GNDA.n1899 GNDA.n444 76.3222
R2198 GNDA.n1895 GNDA.n443 76.3222
R2199 GNDA.n459 GNDA.n442 76.3222
R2200 GNDA.n1161 GNDA.n441 76.3222
R2201 GNDA.n1157 GNDA.n440 76.3222
R2202 GNDA.n1153 GNDA.n439 76.3222
R2203 GNDA.n1149 GNDA.n438 76.3222
R2204 GNDA.n1145 GNDA.n437 76.3222
R2205 GNDA.n508 GNDA.n436 76.3222
R2206 GNDA.n1880 GNDA.n650 76.3222
R2207 GNDA.n1870 GNDA.n649 76.3222
R2208 GNDA.n1795 GNDA.n648 76.3222
R2209 GNDA.n1801 GNDA.n647 76.3222
R2210 GNDA.n1808 GNDA.n646 76.3222
R2211 GNDA.n645 GNDA.n515 76.3222
R2212 GNDA.n1882 GNDA.n521 76.3222
R2213 GNDA.n644 GNDA.n532 76.3222
R2214 GNDA.n565 GNDA.n531 76.3222
R2215 GNDA.n573 GNDA.n530 76.3222
R2216 GNDA.n580 GNDA.n529 76.3222
R2217 GNDA.n555 GNDA.n528 76.3222
R2218 GNDA.n1122 GNDA.n527 76.3222
R2219 GNDA.n1119 GNDA.n526 76.3222
R2220 GNDA.n1112 GNDA.n525 76.3222
R2221 GNDA.n1105 GNDA.n524 76.3222
R2222 GNDA.n1132 GNDA.n523 76.3222
R2223 GNDA.n1138 GNDA.n522 76.3222
R2224 GNDA.n751 GNDA.n750 76.3222
R2225 GNDA.n680 GNDA.n678 76.3222
R2226 GNDA.n758 GNDA.n757 76.3222
R2227 GNDA.n677 GNDA.n675 76.3222
R2228 GNDA.n765 GNDA.n764 76.3222
R2229 GNDA.n674 GNDA.n672 76.3222
R2230 GNDA.n691 GNDA.n690 76.3222
R2231 GNDA.n697 GNDA.n696 76.3222
R2232 GNDA.n689 GNDA.n687 76.3222
R2233 GNDA.n704 GNDA.n703 76.3222
R2234 GNDA.n686 GNDA.n684 76.3222
R2235 GNDA.n711 GNDA.n710 76.3222
R2236 GNDA.n124 GNDA.n122 76.3222
R2237 GNDA.n2093 GNDA.n2092 76.3222
R2238 GNDA.n121 GNDA.n119 76.3222
R2239 GNDA.n2100 GNDA.n2099 76.3222
R2240 GNDA.n118 GNDA.n116 76.3222
R2241 GNDA.n2107 GNDA.n2106 76.3222
R2242 GNDA.n1460 GNDA.n1300 76.3222
R2243 GNDA.n1450 GNDA.n1299 76.3222
R2244 GNDA.n1375 GNDA.n1298 76.3222
R2245 GNDA.n1381 GNDA.n1297 76.3222
R2246 GNDA.n1388 GNDA.n1296 76.3222
R2247 GNDA.n1370 GNDA.n1295 76.3222
R2248 GNDA.n1294 GNDA.n1293 76.3222
R2249 GNDA.n1286 GNDA.n1180 76.3222
R2250 GNDA.n1210 GNDA.n1179 76.3222
R2251 GNDA.n1216 GNDA.n1178 76.3222
R2252 GNDA.n1223 GNDA.n1177 76.3222
R2253 GNDA.n1176 GNDA.n1175 76.3222
R2254 GNDA.n1475 GNDA.n1474 76.3222
R2255 GNDA.n1550 GNDA.n1549 76.3222
R2256 GNDA.n1551 GNDA.n1469 76.3222
R2257 GNDA.n1565 GNDA.n1564 76.3222
R2258 GNDA.n1566 GNDA.n1462 76.3222
R2259 GNDA.n1580 GNDA.n1579 76.3222
R2260 GNDA.n920 GNDA.n671 76.3222
R2261 GNDA.n913 GNDA.n670 76.3222
R2262 GNDA.n909 GNDA.n669 76.3222
R2263 GNDA.n905 GNDA.n668 76.3222
R2264 GNDA.n901 GNDA.n667 76.3222
R2265 GNDA.n1324 GNDA.n658 76.3222
R2266 GNDA.n1328 GNDA.n659 76.3222
R2267 GNDA.n1332 GNDA.n660 76.3222
R2268 GNDA.n1336 GNDA.n661 76.3222
R2269 GNDA.n1340 GNDA.n662 76.3222
R2270 GNDA.n1762 GNDA.n922 76.3222
R2271 GNDA.n1754 GNDA.n654 76.3222
R2272 GNDA.n1750 GNDA.n655 76.3222
R2273 GNDA.n1746 GNDA.n656 76.3222
R2274 GNDA.n657 GNDA.n653 76.3222
R2275 GNDA.t18 GNDA.n260 75.8626
R2276 GNDA.n244 GNDA.t8 75.8626
R2277 GNDA.n1832 GNDA.n1780 74.5978
R2278 GNDA.n1829 GNDA.n1780 74.5978
R2279 GNDA.n1412 GNDA.n1358 74.5978
R2280 GNDA.n1409 GNDA.n1358 74.5978
R2281 GNDA.n853 GNDA.n783 74.5978
R2282 GNDA.n850 GNDA.n783 74.5978
R2283 GNDA.n337 GNDA.n292 74.5978
R2284 GNDA.n334 GNDA.n292 74.5978
R2285 GNDA.n1247 GNDA.n1195 74.5978
R2286 GNDA.n1244 GNDA.n1195 74.5978
R2287 GNDA.n604 GNDA.n543 74.5978
R2288 GNDA.n601 GNDA.n543 74.5978
R2289 GNDA.n1502 GNDA.n1485 74.5978
R2290 GNDA.n1503 GNDA.n1502 74.5978
R2291 GNDA.n2029 GNDA.n61 74.5978
R2292 GNDA.n2032 GNDA.n61 74.5978
R2293 GNDA.n1064 GNDA.n1033 74.5978
R2294 GNDA.n1061 GNDA.n1033 74.5978
R2295 GNDA.n312 GNDA.t207 74.1404
R2296 GNDA.t303 GNDA.t135 70.5544
R2297 GNDA.t135 GNDA.t36 70.5544
R2298 GNDA.t36 GNDA.t75 70.5544
R2299 GNDA.t134 GNDA.t27 70.5544
R2300 GNDA.t27 GNDA.t313 70.5544
R2301 GNDA.n387 GNDA.t203 70.0216
R2302 GNDA.n1874 GNDA.n1770 69.3109
R2303 GNDA.n1850 GNDA.n1770 69.3109
R2304 GNDA.n1454 GNDA.n1348 69.3109
R2305 GNDA.n1430 GNDA.n1348 69.3109
R2306 GNDA.n887 GNDA.n776 69.3109
R2307 GNDA.n887 GNDA.n886 69.3109
R2308 GNDA.n392 GNDA.n391 69.3109
R2309 GNDA.n392 GNDA.n303 69.3109
R2310 GNDA.n1290 GNDA.n1185 69.3109
R2311 GNDA.n1266 GNDA.n1185 69.3109
R2312 GNDA.n638 GNDA.n536 69.3109
R2313 GNDA.n638 GNDA.n637 69.3109
R2314 GNDA.n1543 GNDA.n1542 69.3109
R2315 GNDA.n1542 GNDA.n1541 69.3109
R2316 GNDA.n2213 GNDA.n2212 69.3109
R2317 GNDA.n2213 GNDA.n72 69.3109
R2318 GNDA.n1127 GNDA.n1126 69.3109
R2319 GNDA.n1127 GNDA.n1045 69.3109
R2320 GNDA.t165 GNDA.t45 69.1317
R2321 GNDA.t9 GNDA.t116 69.1317
R2322 GNDA.n2259 GNDA.t98 69.1317
R2323 GNDA.t29 GNDA.t115 69.1317
R2324 GNDA.t110 GNDA.t25 69.1317
R2325 GNDA.t239 GNDA.n1864 65.8183
R2326 GNDA.t239 GNDA.n1789 65.8183
R2327 GNDA.t239 GNDA.n1788 65.8183
R2328 GNDA.t239 GNDA.n1787 65.8183
R2329 GNDA.t239 GNDA.n1778 65.8183
R2330 GNDA.t239 GNDA.n1785 65.8183
R2331 GNDA.t239 GNDA.n1776 65.8183
R2332 GNDA.t239 GNDA.n1786 65.8183
R2333 GNDA.t239 GNDA.n1784 65.8183
R2334 GNDA.t239 GNDA.n1783 65.8183
R2335 GNDA.t239 GNDA.n1782 65.8183
R2336 GNDA.t239 GNDA.n1781 65.8183
R2337 GNDA.t239 GNDA.n1779 65.8183
R2338 GNDA.t239 GNDA.n1777 65.8183
R2339 GNDA.n1865 GNDA.t239 65.8183
R2340 GNDA.t239 GNDA.n1771 65.8183
R2341 GNDA.t274 GNDA.n1444 65.8183
R2342 GNDA.t274 GNDA.n1367 65.8183
R2343 GNDA.t274 GNDA.n1366 65.8183
R2344 GNDA.t274 GNDA.n1365 65.8183
R2345 GNDA.t274 GNDA.n1356 65.8183
R2346 GNDA.t274 GNDA.n1363 65.8183
R2347 GNDA.t274 GNDA.n1354 65.8183
R2348 GNDA.t274 GNDA.n1364 65.8183
R2349 GNDA.t274 GNDA.n1362 65.8183
R2350 GNDA.t274 GNDA.n1361 65.8183
R2351 GNDA.t274 GNDA.n1360 65.8183
R2352 GNDA.t274 GNDA.n1359 65.8183
R2353 GNDA.t274 GNDA.n1357 65.8183
R2354 GNDA.t274 GNDA.n1355 65.8183
R2355 GNDA.n1445 GNDA.t274 65.8183
R2356 GNDA.t274 GNDA.n1349 65.8183
R2357 GNDA.t275 GNDA.n793 65.8183
R2358 GNDA.t275 GNDA.n792 65.8183
R2359 GNDA.t275 GNDA.n791 65.8183
R2360 GNDA.t275 GNDA.n790 65.8183
R2361 GNDA.t275 GNDA.n781 65.8183
R2362 GNDA.t275 GNDA.n788 65.8183
R2363 GNDA.t275 GNDA.n778 65.8183
R2364 GNDA.t275 GNDA.n789 65.8183
R2365 GNDA.t275 GNDA.n787 65.8183
R2366 GNDA.t275 GNDA.n786 65.8183
R2367 GNDA.t275 GNDA.n785 65.8183
R2368 GNDA.t275 GNDA.n784 65.8183
R2369 GNDA.t275 GNDA.n782 65.8183
R2370 GNDA.t275 GNDA.n780 65.8183
R2371 GNDA.t275 GNDA.n779 65.8183
R2372 GNDA.n888 GNDA.t275 65.8183
R2373 GNDA.t229 GNDA.n302 65.8183
R2374 GNDA.t229 GNDA.n301 65.8183
R2375 GNDA.t229 GNDA.n300 65.8183
R2376 GNDA.t229 GNDA.n299 65.8183
R2377 GNDA.t229 GNDA.n290 65.8183
R2378 GNDA.t229 GNDA.n297 65.8183
R2379 GNDA.t229 GNDA.n288 65.8183
R2380 GNDA.t229 GNDA.n298 65.8183
R2381 GNDA.t229 GNDA.n296 65.8183
R2382 GNDA.t229 GNDA.n295 65.8183
R2383 GNDA.t229 GNDA.n294 65.8183
R2384 GNDA.t229 GNDA.n293 65.8183
R2385 GNDA.t229 GNDA.n291 65.8183
R2386 GNDA.n393 GNDA.t229 65.8183
R2387 GNDA.t229 GNDA.n289 65.8183
R2388 GNDA.t229 GNDA.n287 65.8183
R2389 GNDA.t231 GNDA.n1280 65.8183
R2390 GNDA.t231 GNDA.n1204 65.8183
R2391 GNDA.t231 GNDA.n1203 65.8183
R2392 GNDA.t231 GNDA.n1202 65.8183
R2393 GNDA.t231 GNDA.n1193 65.8183
R2394 GNDA.t231 GNDA.n1200 65.8183
R2395 GNDA.t231 GNDA.n1191 65.8183
R2396 GNDA.t231 GNDA.n1201 65.8183
R2397 GNDA.t231 GNDA.n1199 65.8183
R2398 GNDA.t231 GNDA.n1198 65.8183
R2399 GNDA.t231 GNDA.n1197 65.8183
R2400 GNDA.t231 GNDA.n1196 65.8183
R2401 GNDA.t231 GNDA.n1194 65.8183
R2402 GNDA.t231 GNDA.n1192 65.8183
R2403 GNDA.n1281 GNDA.t231 65.8183
R2404 GNDA.t231 GNDA.n1186 65.8183
R2405 GNDA.t226 GNDA.n553 65.8183
R2406 GNDA.t226 GNDA.n552 65.8183
R2407 GNDA.t226 GNDA.n551 65.8183
R2408 GNDA.t226 GNDA.n550 65.8183
R2409 GNDA.t226 GNDA.n541 65.8183
R2410 GNDA.t226 GNDA.n548 65.8183
R2411 GNDA.t226 GNDA.n538 65.8183
R2412 GNDA.t226 GNDA.n549 65.8183
R2413 GNDA.t226 GNDA.n547 65.8183
R2414 GNDA.t226 GNDA.n546 65.8183
R2415 GNDA.t226 GNDA.n545 65.8183
R2416 GNDA.t226 GNDA.n544 65.8183
R2417 GNDA.t226 GNDA.n542 65.8183
R2418 GNDA.t226 GNDA.n540 65.8183
R2419 GNDA.t226 GNDA.n539 65.8183
R2420 GNDA.n639 GNDA.t226 65.8183
R2421 GNDA.n1524 GNDA.t266 65.8183
R2422 GNDA.n1526 GNDA.t266 65.8183
R2423 GNDA.n1532 GNDA.t266 65.8183
R2424 GNDA.n1534 GNDA.t266 65.8183
R2425 GNDA.n1508 GNDA.t266 65.8183
R2426 GNDA.n1510 GNDA.t266 65.8183
R2427 GNDA.n1516 GNDA.t266 65.8183
R2428 GNDA.n1518 GNDA.t266 65.8183
R2429 GNDA.t266 GNDA.n1465 65.8183
R2430 GNDA.n1493 GNDA.t266 65.8183
R2431 GNDA.n1489 GNDA.t266 65.8183
R2432 GNDA.n1500 GNDA.t266 65.8183
R2433 GNDA.n1572 GNDA.t266 65.8183
R2434 GNDA.n1559 GNDA.t266 65.8183
R2435 GNDA.n1557 GNDA.t266 65.8183
R2436 GNDA.n1544 GNDA.t266 65.8183
R2437 GNDA.t232 GNDA.n71 65.8183
R2438 GNDA.t232 GNDA.n70 65.8183
R2439 GNDA.t232 GNDA.n69 65.8183
R2440 GNDA.t232 GNDA.n68 65.8183
R2441 GNDA.t232 GNDA.n59 65.8183
R2442 GNDA.t232 GNDA.n66 65.8183
R2443 GNDA.t232 GNDA.n57 65.8183
R2444 GNDA.t232 GNDA.n67 65.8183
R2445 GNDA.t232 GNDA.n65 65.8183
R2446 GNDA.t232 GNDA.n64 65.8183
R2447 GNDA.t232 GNDA.n63 65.8183
R2448 GNDA.t232 GNDA.n62 65.8183
R2449 GNDA.t232 GNDA.n60 65.8183
R2450 GNDA.n2214 GNDA.t232 65.8183
R2451 GNDA.t232 GNDA.n58 65.8183
R2452 GNDA.t232 GNDA.n56 65.8183
R2453 GNDA.t228 GNDA.n1044 65.8183
R2454 GNDA.t228 GNDA.n1043 65.8183
R2455 GNDA.t228 GNDA.n1042 65.8183
R2456 GNDA.t228 GNDA.n1041 65.8183
R2457 GNDA.t228 GNDA.n1032 65.8183
R2458 GNDA.t228 GNDA.n1039 65.8183
R2459 GNDA.t228 GNDA.n1029 65.8183
R2460 GNDA.t228 GNDA.n1040 65.8183
R2461 GNDA.t228 GNDA.n1038 65.8183
R2462 GNDA.t228 GNDA.n1036 65.8183
R2463 GNDA.t228 GNDA.n1035 65.8183
R2464 GNDA.t228 GNDA.n1034 65.8183
R2465 GNDA.n1128 GNDA.t228 65.8183
R2466 GNDA.t228 GNDA.n1031 65.8183
R2467 GNDA.t228 GNDA.n1030 65.8183
R2468 GNDA.t228 GNDA.n1028 65.8183
R2469 GNDA.n2246 GNDA.n2245 65.0652
R2470 GNDA.n893 GNDA.t197 63.8432
R2471 GNDA.n386 GNDA.t219 63.8432
R2472 GNDA.n2206 GNDA.t213 63.8432
R2473 GNDA.t136 GNDA.t87 62.4857
R2474 GNDA.t1 GNDA.t164 62.4857
R2475 GNDA.t164 GNDA.t2 62.4857
R2476 GNDA.n2261 GNDA.t253 62.2505
R2477 GNDA.n156 GNDA.t293 62.2505
R2478 GNDA.n207 GNDA.t308 62.2505
R2479 GNDA.n202 GNDA.t247 62.2505
R2480 GNDA.n195 GNDA.t235 62.2505
R2481 GNDA.n190 GNDA.t306 62.2505
R2482 GNDA.n189 GNDA.t298 62.2505
R2483 GNDA.n5 GNDA.t318 62.2505
R2484 GNDA.n151 GNDA.t304 62.2505
R2485 GNDA.n199 GNDA.t316 62.2505
R2486 GNDA.n2258 GNDA.t301 62.2505
R2487 GNDA.n2254 GNDA.t314 62.2505
R2488 GNDA.n172 GNDA.t261 60.9987
R2489 GNDA.n183 GNDA.t283 60.9987
R2490 GNDA.t224 GNDA.n6 60.9987
R2491 GNDA.n30 GNDA.t244 60.9987
R2492 GNDA.n824 GNDA.t199 59.7243
R2493 GNDA.n311 GNDA.t221 59.7243
R2494 GNDA.n2058 GNDA.t211 59.7243
R2495 GNDA.t227 GNDA.n427 59.4672
R2496 GNDA.n183 GNDA.n182 59.2425
R2497 GNDA.n9 GNDA.n6 59.2425
R2498 GNDA.n30 GNDA.n29 59.2425
R2499 GNDA.n173 GNDA.n172 59.2425
R2500 GNDA.n895 GNDA.t162 58.6946
R2501 GNDA.t24 GNDA.n808 58.6946
R2502 GNDA.t44 GNDA.n825 58.6946
R2503 GNDA.t239 GNDA.n1770 57.8461
R2504 GNDA.t274 GNDA.n1348 57.8461
R2505 GNDA.t275 GNDA.n887 57.8461
R2506 GNDA.t229 GNDA.n392 57.8461
R2507 GNDA.t231 GNDA.n1185 57.8461
R2508 GNDA.t226 GNDA.n638 57.8461
R2509 GNDA.n1542 GNDA.t266 57.8461
R2510 GNDA.t232 GNDA.n2213 57.8461
R2511 GNDA.t228 GNDA.n1127 57.8461
R2512 GNDA.t189 GNDA.t319 56.6352
R2513 GNDA.t310 GNDA.n2153 56.6352
R2514 GNDA.t321 GNDA.t183 56.6352
R2515 GNDA.n1765 GNDA.n1764 56.3995
R2516 GNDA.n1764 GNDA.n651 56.3995
R2517 GNDA.n1582 GNDA.n1174 56.3995
R2518 GNDA.n2064 GNDA.n1989 56.3995
R2519 GNDA.n2064 GNDA.n2063 56.3995
R2520 GNDA.n1582 GNDA.n1581 56.3995
R2521 GNDA.n1607 GNDA.n1137 56.3995
R2522 GNDA.n1607 GNDA.n1606 56.3995
R2523 GNDA.n769 GNDA.n665 56.3995
R2524 GNDA.n1343 GNDA.n664 56.3995
R2525 GNDA.n2166 GNDA.n2165 55.6055
R2526 GNDA.t239 GNDA.n1780 55.2026
R2527 GNDA.t274 GNDA.n1358 55.2026
R2528 GNDA.t275 GNDA.n783 55.2026
R2529 GNDA.t229 GNDA.n292 55.2026
R2530 GNDA.t231 GNDA.n1195 55.2026
R2531 GNDA.t226 GNDA.n543 55.2026
R2532 GNDA.n1502 GNDA.t266 55.2026
R2533 GNDA.t232 GNDA.n61 55.2026
R2534 GNDA.t228 GNDA.n1033 55.2026
R2535 GNDA.n2151 GNDA.n2150 54.5757
R2536 GNDA.n2191 GNDA.n77 54.5757
R2537 GNDA.t320 GNDA.n2207 54.5757
R2538 GNDA.n1993 GNDA.t39 54.5757
R2539 GNDA.t77 GNDA.n37 54.5757
R2540 GNDA.n265 GNDA.t6 54.5199
R2541 GNDA.t149 GNDA.n240 54.5199
R2542 GNDA.t205 GNDA.n311 53.546
R2543 GNDA.n1847 GNDA.n1786 53.3664
R2544 GNDA.n1844 GNDA.n1776 53.3664
R2545 GNDA.n1840 GNDA.n1785 53.3664
R2546 GNDA.n1836 GNDA.n1778 53.3664
R2547 GNDA.n1825 GNDA.n1781 53.3664
R2548 GNDA.n1821 GNDA.n1782 53.3664
R2549 GNDA.n1817 GNDA.n1783 53.3664
R2550 GNDA.n1813 GNDA.n1784 53.3664
R2551 GNDA.n1873 GNDA.n1771 53.3664
R2552 GNDA.n1866 GNDA.n1865 53.3664
R2553 GNDA.n1798 GNDA.n1777 53.3664
R2554 GNDA.n1805 GNDA.n1779 53.3664
R2555 GNDA.n1864 GNDA.n1863 53.3664
R2556 GNDA.n1791 GNDA.n1789 53.3664
R2557 GNDA.n1858 GNDA.n1788 53.3664
R2558 GNDA.n1854 GNDA.n1787 53.3664
R2559 GNDA.n1864 GNDA.n1790 53.3664
R2560 GNDA.n1859 GNDA.n1789 53.3664
R2561 GNDA.n1855 GNDA.n1788 53.3664
R2562 GNDA.n1851 GNDA.n1787 53.3664
R2563 GNDA.n1833 GNDA.n1778 53.3664
R2564 GNDA.n1837 GNDA.n1785 53.3664
R2565 GNDA.n1841 GNDA.n1776 53.3664
R2566 GNDA.n1845 GNDA.n1786 53.3664
R2567 GNDA.n1816 GNDA.n1784 53.3664
R2568 GNDA.n1820 GNDA.n1783 53.3664
R2569 GNDA.n1824 GNDA.n1782 53.3664
R2570 GNDA.n1828 GNDA.n1781 53.3664
R2571 GNDA.n1812 GNDA.n1779 53.3664
R2572 GNDA.n1804 GNDA.n1777 53.3664
R2573 GNDA.n1865 GNDA.n1775 53.3664
R2574 GNDA.n1774 GNDA.n1771 53.3664
R2575 GNDA.n1427 GNDA.n1364 53.3664
R2576 GNDA.n1424 GNDA.n1354 53.3664
R2577 GNDA.n1420 GNDA.n1363 53.3664
R2578 GNDA.n1416 GNDA.n1356 53.3664
R2579 GNDA.n1405 GNDA.n1359 53.3664
R2580 GNDA.n1401 GNDA.n1360 53.3664
R2581 GNDA.n1397 GNDA.n1361 53.3664
R2582 GNDA.n1393 GNDA.n1362 53.3664
R2583 GNDA.n1453 GNDA.n1349 53.3664
R2584 GNDA.n1446 GNDA.n1445 53.3664
R2585 GNDA.n1378 GNDA.n1355 53.3664
R2586 GNDA.n1385 GNDA.n1357 53.3664
R2587 GNDA.n1444 GNDA.n1443 53.3664
R2588 GNDA.n1369 GNDA.n1367 53.3664
R2589 GNDA.n1438 GNDA.n1366 53.3664
R2590 GNDA.n1434 GNDA.n1365 53.3664
R2591 GNDA.n1444 GNDA.n1368 53.3664
R2592 GNDA.n1439 GNDA.n1367 53.3664
R2593 GNDA.n1435 GNDA.n1366 53.3664
R2594 GNDA.n1431 GNDA.n1365 53.3664
R2595 GNDA.n1413 GNDA.n1356 53.3664
R2596 GNDA.n1417 GNDA.n1363 53.3664
R2597 GNDA.n1421 GNDA.n1354 53.3664
R2598 GNDA.n1425 GNDA.n1364 53.3664
R2599 GNDA.n1396 GNDA.n1362 53.3664
R2600 GNDA.n1400 GNDA.n1361 53.3664
R2601 GNDA.n1404 GNDA.n1360 53.3664
R2602 GNDA.n1408 GNDA.n1359 53.3664
R2603 GNDA.n1392 GNDA.n1357 53.3664
R2604 GNDA.n1384 GNDA.n1355 53.3664
R2605 GNDA.n1445 GNDA.n1353 53.3664
R2606 GNDA.n1352 GNDA.n1349 53.3664
R2607 GNDA.n869 GNDA.n789 53.3664
R2608 GNDA.n865 GNDA.n778 53.3664
R2609 GNDA.n861 GNDA.n788 53.3664
R2610 GNDA.n857 GNDA.n781 53.3664
R2611 GNDA.n846 GNDA.n784 53.3664
R2612 GNDA.n842 GNDA.n785 53.3664
R2613 GNDA.n838 GNDA.n786 53.3664
R2614 GNDA.n834 GNDA.n787 53.3664
R2615 GNDA.n889 GNDA.n888 53.3664
R2616 GNDA.n802 GNDA.n779 53.3664
R2617 GNDA.n815 GNDA.n780 53.3664
R2618 GNDA.n819 GNDA.n782 53.3664
R2619 GNDA.n873 GNDA.n793 53.3664
R2620 GNDA.n874 GNDA.n792 53.3664
R2621 GNDA.n878 GNDA.n791 53.3664
R2622 GNDA.n882 GNDA.n790 53.3664
R2623 GNDA.n870 GNDA.n793 53.3664
R2624 GNDA.n877 GNDA.n792 53.3664
R2625 GNDA.n881 GNDA.n791 53.3664
R2626 GNDA.n794 GNDA.n790 53.3664
R2627 GNDA.n854 GNDA.n781 53.3664
R2628 GNDA.n858 GNDA.n788 53.3664
R2629 GNDA.n862 GNDA.n778 53.3664
R2630 GNDA.n866 GNDA.n789 53.3664
R2631 GNDA.n837 GNDA.n787 53.3664
R2632 GNDA.n841 GNDA.n786 53.3664
R2633 GNDA.n845 GNDA.n785 53.3664
R2634 GNDA.n849 GNDA.n784 53.3664
R2635 GNDA.n833 GNDA.n782 53.3664
R2636 GNDA.n820 GNDA.n780 53.3664
R2637 GNDA.n814 GNDA.n779 53.3664
R2638 GNDA.n888 GNDA.n777 53.3664
R2639 GNDA.n353 GNDA.n298 53.3664
R2640 GNDA.n349 GNDA.n288 53.3664
R2641 GNDA.n345 GNDA.n297 53.3664
R2642 GNDA.n341 GNDA.n290 53.3664
R2643 GNDA.n330 GNDA.n293 53.3664
R2644 GNDA.n326 GNDA.n294 53.3664
R2645 GNDA.n322 GNDA.n295 53.3664
R2646 GNDA.n318 GNDA.n296 53.3664
R2647 GNDA.n304 GNDA.n287 53.3664
R2648 GNDA.n381 GNDA.n289 53.3664
R2649 GNDA.n394 GNDA.n393 53.3664
R2650 GNDA.n305 GNDA.n291 53.3664
R2651 GNDA.n357 GNDA.n302 53.3664
R2652 GNDA.n358 GNDA.n301 53.3664
R2653 GNDA.n362 GNDA.n300 53.3664
R2654 GNDA.n366 GNDA.n299 53.3664
R2655 GNDA.n354 GNDA.n302 53.3664
R2656 GNDA.n361 GNDA.n301 53.3664
R2657 GNDA.n365 GNDA.n300 53.3664
R2658 GNDA.n368 GNDA.n299 53.3664
R2659 GNDA.n338 GNDA.n290 53.3664
R2660 GNDA.n342 GNDA.n297 53.3664
R2661 GNDA.n346 GNDA.n288 53.3664
R2662 GNDA.n350 GNDA.n298 53.3664
R2663 GNDA.n321 GNDA.n296 53.3664
R2664 GNDA.n325 GNDA.n295 53.3664
R2665 GNDA.n329 GNDA.n294 53.3664
R2666 GNDA.n333 GNDA.n293 53.3664
R2667 GNDA.n317 GNDA.n291 53.3664
R2668 GNDA.n393 GNDA.n286 53.3664
R2669 GNDA.n289 GNDA.n285 53.3664
R2670 GNDA.n380 GNDA.n287 53.3664
R2671 GNDA.n1262 GNDA.n1201 53.3664
R2672 GNDA.n1259 GNDA.n1191 53.3664
R2673 GNDA.n1255 GNDA.n1200 53.3664
R2674 GNDA.n1251 GNDA.n1193 53.3664
R2675 GNDA.n1240 GNDA.n1196 53.3664
R2676 GNDA.n1236 GNDA.n1197 53.3664
R2677 GNDA.n1232 GNDA.n1198 53.3664
R2678 GNDA.n1228 GNDA.n1199 53.3664
R2679 GNDA.n1289 GNDA.n1186 53.3664
R2680 GNDA.n1282 GNDA.n1281 53.3664
R2681 GNDA.n1213 GNDA.n1192 53.3664
R2682 GNDA.n1220 GNDA.n1194 53.3664
R2683 GNDA.n1280 GNDA.n1279 53.3664
R2684 GNDA.n1206 GNDA.n1204 53.3664
R2685 GNDA.n1274 GNDA.n1203 53.3664
R2686 GNDA.n1270 GNDA.n1202 53.3664
R2687 GNDA.n1280 GNDA.n1205 53.3664
R2688 GNDA.n1275 GNDA.n1204 53.3664
R2689 GNDA.n1271 GNDA.n1203 53.3664
R2690 GNDA.n1267 GNDA.n1202 53.3664
R2691 GNDA.n1248 GNDA.n1193 53.3664
R2692 GNDA.n1252 GNDA.n1200 53.3664
R2693 GNDA.n1256 GNDA.n1191 53.3664
R2694 GNDA.n1260 GNDA.n1201 53.3664
R2695 GNDA.n1231 GNDA.n1199 53.3664
R2696 GNDA.n1235 GNDA.n1198 53.3664
R2697 GNDA.n1239 GNDA.n1197 53.3664
R2698 GNDA.n1243 GNDA.n1196 53.3664
R2699 GNDA.n1227 GNDA.n1194 53.3664
R2700 GNDA.n1219 GNDA.n1192 53.3664
R2701 GNDA.n1281 GNDA.n1190 53.3664
R2702 GNDA.n1189 GNDA.n1186 53.3664
R2703 GNDA.n620 GNDA.n549 53.3664
R2704 GNDA.n616 GNDA.n538 53.3664
R2705 GNDA.n612 GNDA.n548 53.3664
R2706 GNDA.n608 GNDA.n541 53.3664
R2707 GNDA.n597 GNDA.n544 53.3664
R2708 GNDA.n593 GNDA.n545 53.3664
R2709 GNDA.n589 GNDA.n546 53.3664
R2710 GNDA.n585 GNDA.n547 53.3664
R2711 GNDA.n640 GNDA.n639 53.3664
R2712 GNDA.n562 GNDA.n539 53.3664
R2713 GNDA.n570 GNDA.n540 53.3664
R2714 GNDA.n577 GNDA.n542 53.3664
R2715 GNDA.n624 GNDA.n553 53.3664
R2716 GNDA.n625 GNDA.n552 53.3664
R2717 GNDA.n629 GNDA.n551 53.3664
R2718 GNDA.n633 GNDA.n550 53.3664
R2719 GNDA.n621 GNDA.n553 53.3664
R2720 GNDA.n628 GNDA.n552 53.3664
R2721 GNDA.n632 GNDA.n551 53.3664
R2722 GNDA.n554 GNDA.n550 53.3664
R2723 GNDA.n605 GNDA.n541 53.3664
R2724 GNDA.n609 GNDA.n548 53.3664
R2725 GNDA.n613 GNDA.n538 53.3664
R2726 GNDA.n617 GNDA.n549 53.3664
R2727 GNDA.n588 GNDA.n547 53.3664
R2728 GNDA.n592 GNDA.n546 53.3664
R2729 GNDA.n596 GNDA.n545 53.3664
R2730 GNDA.n600 GNDA.n544 53.3664
R2731 GNDA.n584 GNDA.n542 53.3664
R2732 GNDA.n576 GNDA.n540 53.3664
R2733 GNDA.n569 GNDA.n539 53.3664
R2734 GNDA.n639 GNDA.n537 53.3664
R2735 GNDA.n1518 GNDA.n1481 53.3664
R2736 GNDA.n1517 GNDA.n1516 53.3664
R2737 GNDA.n1510 GNDA.n1483 53.3664
R2738 GNDA.n1509 GNDA.n1508 53.3664
R2739 GNDA.n1500 GNDA.n1499 53.3664
R2740 GNDA.n1495 GNDA.n1489 53.3664
R2741 GNDA.n1493 GNDA.n1492 53.3664
R2742 GNDA.n1574 GNDA.n1465 53.3664
R2743 GNDA.n1545 GNDA.n1544 53.3664
R2744 GNDA.n1557 GNDA.n1556 53.3664
R2745 GNDA.n1560 GNDA.n1559 53.3664
R2746 GNDA.n1572 GNDA.n1571 53.3664
R2747 GNDA.n1525 GNDA.n1524 53.3664
R2748 GNDA.n1527 GNDA.n1526 53.3664
R2749 GNDA.n1532 GNDA.n1531 53.3664
R2750 GNDA.n1535 GNDA.n1534 53.3664
R2751 GNDA.n1524 GNDA.n1523 53.3664
R2752 GNDA.n1526 GNDA.n1479 53.3664
R2753 GNDA.n1533 GNDA.n1532 53.3664
R2754 GNDA.n1534 GNDA.n1477 53.3664
R2755 GNDA.n1508 GNDA.n1507 53.3664
R2756 GNDA.n1511 GNDA.n1510 53.3664
R2757 GNDA.n1516 GNDA.n1515 53.3664
R2758 GNDA.n1519 GNDA.n1518 53.3664
R2759 GNDA.n1490 GNDA.n1465 53.3664
R2760 GNDA.n1494 GNDA.n1493 53.3664
R2761 GNDA.n1489 GNDA.n1487 53.3664
R2762 GNDA.n1501 GNDA.n1500 53.3664
R2763 GNDA.n1573 GNDA.n1572 53.3664
R2764 GNDA.n1559 GNDA.n1466 53.3664
R2765 GNDA.n1558 GNDA.n1557 53.3664
R2766 GNDA.n1544 GNDA.n1471 53.3664
R2767 GNDA.n2013 GNDA.n67 53.3664
R2768 GNDA.n2017 GNDA.n57 53.3664
R2769 GNDA.n2021 GNDA.n66 53.3664
R2770 GNDA.n2025 GNDA.n59 53.3664
R2771 GNDA.n2036 GNDA.n62 53.3664
R2772 GNDA.n2040 GNDA.n63 53.3664
R2773 GNDA.n2044 GNDA.n64 53.3664
R2774 GNDA.n2049 GNDA.n65 53.3664
R2775 GNDA.n73 GNDA.n56 53.3664
R2776 GNDA.n2202 GNDA.n58 53.3664
R2777 GNDA.n2215 GNDA.n2214 53.3664
R2778 GNDA.n2053 GNDA.n60 53.3664
R2779 GNDA.n2009 GNDA.n71 53.3664
R2780 GNDA.n2008 GNDA.n70 53.3664
R2781 GNDA.n2004 GNDA.n69 53.3664
R2782 GNDA.n2000 GNDA.n68 53.3664
R2783 GNDA.n2012 GNDA.n71 53.3664
R2784 GNDA.n2005 GNDA.n70 53.3664
R2785 GNDA.n2001 GNDA.n69 53.3664
R2786 GNDA.n1997 GNDA.n68 53.3664
R2787 GNDA.n2028 GNDA.n59 53.3664
R2788 GNDA.n2024 GNDA.n66 53.3664
R2789 GNDA.n2020 GNDA.n57 53.3664
R2790 GNDA.n2016 GNDA.n67 53.3664
R2791 GNDA.n2045 GNDA.n65 53.3664
R2792 GNDA.n2041 GNDA.n64 53.3664
R2793 GNDA.n2037 GNDA.n63 53.3664
R2794 GNDA.n2033 GNDA.n62 53.3664
R2795 GNDA.n2050 GNDA.n60 53.3664
R2796 GNDA.n2214 GNDA.n55 53.3664
R2797 GNDA.n58 GNDA.n54 53.3664
R2798 GNDA.n2201 GNDA.n56 53.3664
R2799 GNDA.n1080 GNDA.n1040 53.3664
R2800 GNDA.n1076 GNDA.n1029 53.3664
R2801 GNDA.n1072 GNDA.n1039 53.3664
R2802 GNDA.n1068 GNDA.n1032 53.3664
R2803 GNDA.n1057 GNDA.n1034 53.3664
R2804 GNDA.n1053 GNDA.n1035 53.3664
R2805 GNDA.n1049 GNDA.n1036 53.3664
R2806 GNDA.n1038 GNDA.n1037 53.3664
R2807 GNDA.n1046 GNDA.n1028 53.3664
R2808 GNDA.n1115 GNDA.n1030 53.3664
R2809 GNDA.n1108 GNDA.n1031 53.3664
R2810 GNDA.n1129 GNDA.n1128 53.3664
R2811 GNDA.n1084 GNDA.n1044 53.3664
R2812 GNDA.n1085 GNDA.n1043 53.3664
R2813 GNDA.n1089 GNDA.n1042 53.3664
R2814 GNDA.n1093 GNDA.n1041 53.3664
R2815 GNDA.n1081 GNDA.n1044 53.3664
R2816 GNDA.n1088 GNDA.n1043 53.3664
R2817 GNDA.n1092 GNDA.n1042 53.3664
R2818 GNDA.n1095 GNDA.n1041 53.3664
R2819 GNDA.n1065 GNDA.n1032 53.3664
R2820 GNDA.n1069 GNDA.n1039 53.3664
R2821 GNDA.n1073 GNDA.n1029 53.3664
R2822 GNDA.n1077 GNDA.n1040 53.3664
R2823 GNDA.n1048 GNDA.n1038 53.3664
R2824 GNDA.n1052 GNDA.n1036 53.3664
R2825 GNDA.n1056 GNDA.n1035 53.3664
R2826 GNDA.n1060 GNDA.n1034 53.3664
R2827 GNDA.n1128 GNDA.n1027 53.3664
R2828 GNDA.n1031 GNDA.n1026 53.3664
R2829 GNDA.n1107 GNDA.n1030 53.3664
R2830 GNDA.n1114 GNDA.n1028 53.3664
R2831 GNDA.t13 GNDA.t151 52.8656
R2832 GNDA.t102 GNDA.t125 52.8656
R2833 GNDA.t67 GNDA.t17 52.8656
R2834 GNDA.t100 GNDA.t28 52.8656
R2835 GNDA.t64 GNDA.t177 52.8656
R2836 GNDA.t227 GNDA.n2179 51.4866
R2837 GNDA.n2180 GNDA.t227 51.4866
R2838 GNDA.t185 GNDA.n386 49.4271
R2839 GNDA.n172 GNDA.n171 48.799
R2840 GNDA.n184 GNDA.n183 48.799
R2841 GNDA.t176 GNDA.t122 48.799
R2842 GNDA.t322 GNDA.t58 48.799
R2843 GNDA.t234 GNDA.t49 48.799
R2844 GNDA.n197 GNDA.t35 48.799
R2845 GNDA.t300 GNDA.t141 48.799
R2846 GNDA.t175 GNDA.t60 48.799
R2847 GNDA.t51 GNDA.t124 48.799
R2848 GNDA.t8 GNDA.t69 48.799
R2849 GNDA.t114 GNDA.t85 48.799
R2850 GNDA.n2252 GNDA.n6 48.799
R2851 GNDA.n2246 GNDA.n30 48.799
R2852 GNDA.t81 GNDA.n77 48.3974
R2853 GNDA.n1629 GNDA.n1013 48.2167
R2854 GNDA.n1623 GNDA.n1013 48.2167
R2855 GNDA.n1623 GNDA.n1622 48.2167
R2856 GNDA.n1622 GNDA.n1621 48.2167
R2857 GNDA.n1621 GNDA.n431 48.2167
R2858 GNDA.n1614 GNDA.n430 48.2167
R2859 GNDA.n1614 GNDA.n1613 48.2167
R2860 GNDA.n1613 GNDA.n1612 48.2167
R2861 GNDA.n1612 GNDA.n1020 48.2167
R2862 GNDA.n1139 GNDA.n1020 48.2167
R2863 GNDA.n1605 GNDA.n1139 48.2167
R2864 GNDA.n1605 GNDA.t57 48.2167
R2865 GNDA.n1604 GNDA.n1140 48.2167
R2866 GNDA.n1598 GNDA.n1140 48.2167
R2867 GNDA.n1598 GNDA.n1597 48.2167
R2868 GNDA.n1597 GNDA.n1596 48.2167
R2869 GNDA.n1596 GNDA.n429 48.2167
R2870 GNDA.n1589 GNDA.n428 48.2167
R2871 GNDA.n1589 GNDA.n1588 48.2167
R2872 GNDA.n1588 GNDA.n1587 48.2167
R2873 GNDA.n1587 GNDA.n1169 48.2167
R2874 GNDA.n1173 GNDA.n1169 48.2167
R2875 GNDA.n1173 GNDA.n427 48.2167
R2876 GNDA.n2085 GNDA.n2084 48.2167
R2877 GNDA.n2084 GNDA.n2083 48.2167
R2878 GNDA.n2083 GNDA.n1980 48.2167
R2879 GNDA.n2077 GNDA.n1980 48.2167
R2880 GNDA.n2077 GNDA.n49 48.2167
R2881 GNDA.n1987 GNDA.n50 48.2167
R2882 GNDA.n2070 GNDA.n1987 48.2167
R2883 GNDA.n2070 GNDA.n2069 48.2167
R2884 GNDA.n2069 GNDA.n2068 48.2167
R2885 GNDA.n2068 GNDA.n1988 48.2167
R2886 GNDA.n2062 GNDA.n1988 48.2167
R2887 GNDA.n255 GNDA.t105 48.0005
R2888 GNDA.n255 GNDA.t93 48.0005
R2889 GNDA.n253 GNDA.t91 48.0005
R2890 GNDA.n253 GNDA.t155 48.0005
R2891 GNDA.n251 GNDA.t180 48.0005
R2892 GNDA.n251 GNDA.t95 48.0005
R2893 GNDA.n249 GNDA.t130 48.0005
R2894 GNDA.n249 GNDA.t56 48.0005
R2895 GNDA.n247 GNDA.t15 48.0005
R2896 GNDA.n247 GNDA.t89 48.0005
R2897 GNDA.t227 GNDA.n1979 47.6748
R2898 GNDA.n2165 GNDA.t5 47.3677
R2899 GNDA.t268 GNDA.t21 46.338
R2900 GNDA.t258 GNDA.t79 46.338
R2901 GNDA.n1732 GNDA.t227 46.2335
R2902 GNDA.n1670 GNDA.t227 46.2335
R2903 GNDA.t227 GNDA.n1005 46.2335
R2904 GNDA.n145 GNDA.n31 44.0005
R2905 GNDA.n269 GNDA.n268 43.5649
R2906 GNDA.n894 GNDA.t268 43.2488
R2907 GNDA.n387 GNDA.t185 43.2488
R2908 GNDA.n2207 GNDA.t209 43.2488
R2909 GNDA.t227 GNDA.n1731 42.2987
R2910 GNDA.t227 GNDA.n945 42.2987
R2911 GNDA.n1639 GNDA.t227 42.2987
R2912 GNDA.t333 GNDA.t126 42.2405
R2913 GNDA.t325 GNDA.t333 42.2405
R2914 GNDA.t82 GNDA.t335 42.2405
R2915 GNDA.t53 GNDA.t82 42.2405
R2916 GNDA.n375 GNDA.t62 42.2191
R2917 GNDA.t227 GNDA.t5 41.1894
R2918 GNDA.t227 GNDA.t81 41.1894
R2919 GNDA.t18 GNDA.t122 40.6659
R2920 GNDA.t58 GNDA.t176 40.6659
R2921 GNDA.t322 GNDA.t49 40.6659
R2922 GNDA.t234 GNDA.t67 40.6659
R2923 GNDA.t96 GNDA.n197 40.6659
R2924 GNDA.n239 GNDA.t273 40.4338
R2925 GNDA.n150 GNDA.t238 40.4338
R2926 GNDA.n418 GNDA.n43 39.3903
R2927 GNDA.n825 GNDA.t191 39.1299
R2928 GNDA.n399 GNDA.n398 39.1299
R2929 GNDA.n312 GNDA.t205 39.1299
R2930 GNDA.n2059 GNDA.t258 39.1299
R2931 GNDA.t324 GNDA.t1 38.533
R2932 GNDA.n264 GNDA.t19 38.485
R2933 GNDA.t107 GNDA.n242 38.485
R2934 GNDA.t11 GNDA.n241 38.485
R2935 GNDA.n263 GNDA.t106 38.485
R2936 GNDA.n262 GNDA.t47 38.485
R2937 GNDA.n261 GNDA.t18 38.485
R2938 GNDA.t0 GNDA.n243 38.485
R2939 GNDA.n275 GNDA.n274 38.4845
R2940 GNDA.n2179 GNDA.n85 38.1002
R2941 GNDA.n2151 GNDA.n97 38.1002
R2942 GNDA.n2219 GNDA.t39 38.1002
R2943 GNDA.n2059 GNDA.t77 38.1002
R2944 GNDA.n236 GNDA.n235 37.5297
R2945 GNDA.n234 GNDA.n233 37.5297
R2946 GNDA.n232 GNDA.n231 37.5297
R2947 GNDA.n230 GNDA.n229 37.5297
R2948 GNDA.n228 GNDA.n227 37.5297
R2949 GNDA.n226 GNDA.n225 37.5297
R2950 GNDA.n224 GNDA.n223 37.5297
R2951 GNDA.n222 GNDA.n221 37.5297
R2952 GNDA.n220 GNDA.n219 37.5297
R2953 GNDA.n218 GNDA.n217 37.5297
R2954 GNDA.n216 GNDA.n215 37.5297
R2955 GNDA.n2180 GNDA.n80 37.0705
R2956 GNDA.t151 GNDA.t329 36.5994
R2957 GNDA.t323 GNDA.t102 36.5994
R2958 GNDA.n157 GNDA.t85 36.5994
R2959 GNDA.t158 GNDA.t100 36.5994
R2960 GNDA.t177 GNDA.t41 36.5994
R2961 GNDA.t227 GNDA.t215 36.0408
R2962 GNDA.t227 GNDA.t195 36.0408
R2963 GNDA.n2233 GNDA.n2232 35.3278
R2964 GNDA.t162 GNDA.n894 33.9813
R2965 GNDA.n809 GNDA.t24 33.9813
R2966 GNDA.n2153 GNDA.n96 33.9813
R2967 GNDA.n800 GNDA.t199 32.9516
R2968 GNDA.t221 GNDA.n310 32.9516
R2969 GNDA.t211 GNDA.n2057 32.9516
R2970 GNDA.t227 GNDA.n422 32.9056
R2971 GNDA.t227 GNDA.n421 32.9056
R2972 GNDA.t227 GNDA.n431 32.6804
R2973 GNDA.t227 GNDA.n429 32.6804
R2974 GNDA.t227 GNDA.n49 32.6804
R2975 GNDA.n2237 GNDA.n2236 32.3063
R2976 GNDA.t19 GNDA.n263 32.071
R2977 GNDA.t106 GNDA.n262 32.071
R2978 GNDA.t47 GNDA.n261 32.071
R2979 GNDA.n243 GNDA.t107 32.071
R2980 GNDA.t6 GNDA.n264 32.071
R2981 GNDA.n242 GNDA.t11 32.071
R2982 GNDA.n241 GNDA.t149 32.071
R2983 GNDA.n188 GNDA.n5 31.5738
R2984 GNDA.n185 GNDA.t284 31.1255
R2985 GNDA.n170 GNDA.t262 31.1255
R2986 GNDA.n2251 GNDA.t225 31.1255
R2987 GNDA.n2247 GNDA.t245 31.1255
R2988 GNDA.n27 GNDA.n26 30.8755
R2989 GNDA.n175 GNDA.n169 30.813
R2990 GNDA.n2265 GNDA.n0 30.4627
R2991 GNDA.n208 GNDA.n207 29.8672
R2992 GNDA.n152 GNDA.n151 29.8672
R2993 GNDA.n2255 GNDA.n2254 29.8672
R2994 GNDA.n807 GNDA.t197 28.8327
R2995 GNDA.t219 GNDA.n385 28.8327
R2996 GNDA.t213 GNDA.n2196 28.8327
R2997 GNDA.t319 GNDA.n807 27.803
R2998 GNDA.t12 GNDA.n824 27.803
R2999 GNDA.n828 GNDA.t163 27.803
R3000 GNDA.n1849 GNDA.n1848 27.5561
R3001 GNDA.n1429 GNDA.n1428 27.5561
R3002 GNDA.n871 GNDA.n868 27.5561
R3003 GNDA.n355 GNDA.n352 27.5561
R3004 GNDA.n1264 GNDA.n1263 27.5561
R3005 GNDA.n622 GNDA.n619 27.5561
R3006 GNDA.n1522 GNDA.n1521 27.5561
R3007 GNDA.n2014 GNDA.n2011 27.5561
R3008 GNDA.n1082 GNDA.n1079 27.5561
R3009 GNDA.t156 GNDA.n35 26.7873
R3010 GNDA.n1831 GNDA.n1830 26.6672
R3011 GNDA.n1411 GNDA.n1410 26.6672
R3012 GNDA.n852 GNDA.n851 26.6672
R3013 GNDA.n336 GNDA.n335 26.6672
R3014 GNDA.n1246 GNDA.n1245 26.6672
R3015 GNDA.n603 GNDA.n602 26.6672
R3016 GNDA.n1505 GNDA.n1504 26.6672
R3017 GNDA.n2031 GNDA.n2030 26.6672
R3018 GNDA.n1063 GNDA.n1062 26.6672
R3019 GNDA.t191 GNDA.t12 25.7435
R3020 GNDA.t209 GNDA.t80 25.7435
R3021 GNDA.n409 GNDA.n408 25.3679
R3022 GNDA.t300 GNDA.t327 24.3998
R3023 GNDA.t175 GNDA.t76 24.3998
R3024 GNDA.t166 GNDA.t124 24.3998
R3025 GNDA.t8 GNDA.t334 24.3998
R3026 GNDA.t114 GNDA.t292 24.3998
R3027 GNDA.n130 GNDA.t198 24.0005
R3028 GNDA.n130 GNDA.t190 24.0005
R3029 GNDA.n128 GNDA.t216 24.0005
R3030 GNDA.n128 GNDA.t200 24.0005
R3031 GNDA.n86 GNDA.t192 24.0005
R3032 GNDA.n86 GNDA.t218 24.0005
R3033 GNDA.n2174 GNDA.t204 24.0005
R3034 GNDA.n2174 GNDA.t186 24.0005
R3035 GNDA.n2172 GNDA.t220 24.0005
R3036 GNDA.n2172 GNDA.t202 24.0005
R3037 GNDA.n2170 GNDA.t194 24.0005
R3038 GNDA.n2170 GNDA.t222 24.0005
R3039 GNDA.n78 GNDA.t206 24.0005
R3040 GNDA.n78 GNDA.t208 24.0005
R3041 GNDA.n2186 GNDA.t188 24.0005
R3042 GNDA.n2186 GNDA.t210 24.0005
R3043 GNDA.n2184 GNDA.t214 24.0005
R3044 GNDA.n2184 GNDA.t196 24.0005
R3045 GNDA.n38 GNDA.t184 24.0005
R3046 GNDA.n38 GNDA.t212 24.0005
R3047 GNDA.t128 GNDA.t324 23.9532
R3048 GNDA.n2192 GNDA.t40 23.6841
R3049 GNDA.t80 GNDA.n2206 23.6841
R3050 GNDA.n2057 GNDA.t321 23.6841
R3051 GNDA.t203 GNDA.n96 22.6544
R3052 GNDA.n2208 GNDA.t187 22.6544
R3053 GNDA.n2265 GNDA.n2264 21.383
R3054 GNDA.n949 GNDA.n948 21.0192
R3055 GNDA.n133 GNDA.n132 20.8233
R3056 GNDA.n2168 GNDA.n2167 20.8233
R3057 GNDA.n2178 GNDA.n2177 20.8233
R3058 GNDA.n2182 GNDA.n2181 20.8233
R3059 GNDA.n2190 GNDA.n2189 20.8233
R3060 GNDA.n2241 GNDA.n2240 20.8233
R3061 GNDA.t227 GNDA.n420 20.5949
R3062 GNDA.t161 GNDA.n420 20.5949
R3063 GNDA.n2166 GNDA.t163 20.5949
R3064 GNDA.t40 GNDA.n2191 20.5949
R3065 GNDA.n2230 GNDA.t78 20.5949
R3066 GNDA.n2230 GNDA.t227 20.5949
R3067 GNDA.t45 GNDA.t147 20.3332
R3068 GNDA.t340 GNDA.t9 20.3332
R3069 GNDA.n200 GNDA.t31 20.3332
R3070 GNDA.t43 GNDA.t29 20.3332
R3071 GNDA.t25 GNDA.t4 20.3332
R3072 GNDA.t227 GNDA.n403 19.9378
R3073 GNDA.n25 GNDA.t7 19.7005
R3074 GNDA.n25 GNDA.t72 19.7005
R3075 GNDA.n23 GNDA.t109 19.7005
R3076 GNDA.n23 GNDA.t159 19.7005
R3077 GNDA.n21 GNDA.t108 19.7005
R3078 GNDA.n21 GNDA.t111 19.7005
R3079 GNDA.n19 GNDA.t66 19.7005
R3080 GNDA.n19 GNDA.t160 19.7005
R3081 GNDA.n17 GNDA.t42 19.7005
R3082 GNDA.n17 GNDA.t65 19.7005
R3083 GNDA.n16 GNDA.t71 19.7005
R3084 GNDA.n16 GNDA.t22 19.7005
R3085 GNDA.n168 GNDA.t182 19.7005
R3086 GNDA.n168 GNDA.t328 19.7005
R3087 GNDA.n166 GNDA.t138 19.7005
R3088 GNDA.n166 GNDA.t331 19.7005
R3089 GNDA.n164 GNDA.t132 19.7005
R3090 GNDA.n164 GNDA.t133 19.7005
R3091 GNDA.n162 GNDA.t146 19.7005
R3092 GNDA.n162 GNDA.t336 19.7005
R3093 GNDA.n160 GNDA.t3 19.7005
R3094 GNDA.n160 GNDA.t330 19.7005
R3095 GNDA.n159 GNDA.t145 19.7005
R3096 GNDA.n159 GNDA.t143 19.7005
R3097 GNDA.t227 GNDA.n423 19.6741
R3098 GNDA.n2243 GNDA.t156 19.287
R3099 GNDA.n1668 GNDA.n1667 18.5605
R3100 GNDA.n826 GNDA.t217 18.5355
R3101 GNDA.t207 GNDA.n97 18.5355
R3102 GNDA.n194 GNDA.n188 18.4151
R3103 GNDA GNDA.n42 18.1546
R3104 GNDA.n2256 GNDA.n2255 18.0922
R3105 GNDA.n1602 GNDA.n1163 17.5843
R3106 GNDA.n2088 GNDA.n123 17.5843
R3107 GNDA.n1627 GNDA.n1011 17.5843
R3108 GNDA.t227 GNDA.n134 17.5058
R3109 GNDA.n2243 GNDA.n2242 17.5058
R3110 GNDA.n1760 GNDA.n1743 16.9379
R3111 GNDA.n1322 GNDA.n1319 16.9379
R3112 GNDA.n918 GNDA.n768 16.9379
R3113 GNDA.n1892 GNDA.n1891 16.7709
R3114 GNDA.n1947 GNDA.n114 16.7709
R3115 GNDA.n747 GNDA.n486 16.7709
R3116 GNDA.n1975 GNDA.n457 16.7709
R3117 GNDA.n200 GNDA.t17 16.2667
R3118 GNDA.t173 GNDA.t252 16.2667
R3119 GNDA.t327 GNDA.t98 16.2667
R3120 GNDA.t76 GNDA.t141 16.2667
R3121 GNDA.t60 GNDA.t166 16.2667
R3122 GNDA.t334 GNDA.t51 16.2667
R3123 GNDA.t292 GNDA.t69 16.2667
R3124 GNDA.n177 GNDA.n176 16.2608
R3125 GNDA.n179 GNDA.n178 16.2608
R3126 GNDA.n13 GNDA.n12 16.2608
R3127 GNDA.n15 GNDA.n14 16.2608
R3128 GNDA.t75 GNDA.n265 16.036
R3129 GNDA.n240 GNDA.t134 16.036
R3130 GNDA.n1862 GNDA.n1849 16.0005
R3131 GNDA.n1862 GNDA.n1861 16.0005
R3132 GNDA.n1861 GNDA.n1860 16.0005
R3133 GNDA.n1860 GNDA.n1857 16.0005
R3134 GNDA.n1857 GNDA.n1856 16.0005
R3135 GNDA.n1856 GNDA.n1853 16.0005
R3136 GNDA.n1853 GNDA.n1852 16.0005
R3137 GNDA.n1852 GNDA.n1767 16.0005
R3138 GNDA.n1848 GNDA.n1846 16.0005
R3139 GNDA.n1846 GNDA.n1843 16.0005
R3140 GNDA.n1843 GNDA.n1842 16.0005
R3141 GNDA.n1842 GNDA.n1839 16.0005
R3142 GNDA.n1839 GNDA.n1838 16.0005
R3143 GNDA.n1838 GNDA.n1835 16.0005
R3144 GNDA.n1835 GNDA.n1834 16.0005
R3145 GNDA.n1834 GNDA.n1831 16.0005
R3146 GNDA.n1830 GNDA.n1827 16.0005
R3147 GNDA.n1827 GNDA.n1826 16.0005
R3148 GNDA.n1826 GNDA.n1823 16.0005
R3149 GNDA.n1823 GNDA.n1822 16.0005
R3150 GNDA.n1822 GNDA.n1819 16.0005
R3151 GNDA.n1819 GNDA.n1818 16.0005
R3152 GNDA.n1818 GNDA.n1815 16.0005
R3153 GNDA.n1815 GNDA.n1814 16.0005
R3154 GNDA.n1442 GNDA.n1429 16.0005
R3155 GNDA.n1442 GNDA.n1441 16.0005
R3156 GNDA.n1441 GNDA.n1440 16.0005
R3157 GNDA.n1440 GNDA.n1437 16.0005
R3158 GNDA.n1437 GNDA.n1436 16.0005
R3159 GNDA.n1436 GNDA.n1433 16.0005
R3160 GNDA.n1433 GNDA.n1432 16.0005
R3161 GNDA.n1432 GNDA.n1345 16.0005
R3162 GNDA.n1428 GNDA.n1426 16.0005
R3163 GNDA.n1426 GNDA.n1423 16.0005
R3164 GNDA.n1423 GNDA.n1422 16.0005
R3165 GNDA.n1422 GNDA.n1419 16.0005
R3166 GNDA.n1419 GNDA.n1418 16.0005
R3167 GNDA.n1418 GNDA.n1415 16.0005
R3168 GNDA.n1415 GNDA.n1414 16.0005
R3169 GNDA.n1414 GNDA.n1411 16.0005
R3170 GNDA.n1410 GNDA.n1407 16.0005
R3171 GNDA.n1407 GNDA.n1406 16.0005
R3172 GNDA.n1406 GNDA.n1403 16.0005
R3173 GNDA.n1403 GNDA.n1402 16.0005
R3174 GNDA.n1402 GNDA.n1399 16.0005
R3175 GNDA.n1399 GNDA.n1398 16.0005
R3176 GNDA.n1398 GNDA.n1395 16.0005
R3177 GNDA.n1395 GNDA.n1394 16.0005
R3178 GNDA.n872 GNDA.n871 16.0005
R3179 GNDA.n875 GNDA.n872 16.0005
R3180 GNDA.n876 GNDA.n875 16.0005
R3181 GNDA.n879 GNDA.n876 16.0005
R3182 GNDA.n880 GNDA.n879 16.0005
R3183 GNDA.n883 GNDA.n880 16.0005
R3184 GNDA.n884 GNDA.n883 16.0005
R3185 GNDA.n885 GNDA.n884 16.0005
R3186 GNDA.n868 GNDA.n867 16.0005
R3187 GNDA.n867 GNDA.n864 16.0005
R3188 GNDA.n864 GNDA.n863 16.0005
R3189 GNDA.n863 GNDA.n860 16.0005
R3190 GNDA.n860 GNDA.n859 16.0005
R3191 GNDA.n859 GNDA.n856 16.0005
R3192 GNDA.n856 GNDA.n855 16.0005
R3193 GNDA.n855 GNDA.n852 16.0005
R3194 GNDA.n851 GNDA.n848 16.0005
R3195 GNDA.n848 GNDA.n847 16.0005
R3196 GNDA.n847 GNDA.n844 16.0005
R3197 GNDA.n844 GNDA.n843 16.0005
R3198 GNDA.n843 GNDA.n840 16.0005
R3199 GNDA.n840 GNDA.n839 16.0005
R3200 GNDA.n839 GNDA.n836 16.0005
R3201 GNDA.n836 GNDA.n835 16.0005
R3202 GNDA.n356 GNDA.n355 16.0005
R3203 GNDA.n359 GNDA.n356 16.0005
R3204 GNDA.n360 GNDA.n359 16.0005
R3205 GNDA.n363 GNDA.n360 16.0005
R3206 GNDA.n364 GNDA.n363 16.0005
R3207 GNDA.n367 GNDA.n364 16.0005
R3208 GNDA.n369 GNDA.n367 16.0005
R3209 GNDA.n370 GNDA.n369 16.0005
R3210 GNDA.n352 GNDA.n351 16.0005
R3211 GNDA.n351 GNDA.n348 16.0005
R3212 GNDA.n348 GNDA.n347 16.0005
R3213 GNDA.n347 GNDA.n344 16.0005
R3214 GNDA.n344 GNDA.n343 16.0005
R3215 GNDA.n343 GNDA.n340 16.0005
R3216 GNDA.n340 GNDA.n339 16.0005
R3217 GNDA.n339 GNDA.n336 16.0005
R3218 GNDA.n335 GNDA.n332 16.0005
R3219 GNDA.n332 GNDA.n331 16.0005
R3220 GNDA.n331 GNDA.n328 16.0005
R3221 GNDA.n328 GNDA.n327 16.0005
R3222 GNDA.n327 GNDA.n324 16.0005
R3223 GNDA.n324 GNDA.n323 16.0005
R3224 GNDA.n323 GNDA.n320 16.0005
R3225 GNDA.n320 GNDA.n319 16.0005
R3226 GNDA.n1278 GNDA.n1264 16.0005
R3227 GNDA.n1278 GNDA.n1277 16.0005
R3228 GNDA.n1277 GNDA.n1276 16.0005
R3229 GNDA.n1276 GNDA.n1273 16.0005
R3230 GNDA.n1273 GNDA.n1272 16.0005
R3231 GNDA.n1272 GNDA.n1269 16.0005
R3232 GNDA.n1269 GNDA.n1268 16.0005
R3233 GNDA.n1268 GNDA.n1265 16.0005
R3234 GNDA.n1263 GNDA.n1261 16.0005
R3235 GNDA.n1261 GNDA.n1258 16.0005
R3236 GNDA.n1258 GNDA.n1257 16.0005
R3237 GNDA.n1257 GNDA.n1254 16.0005
R3238 GNDA.n1254 GNDA.n1253 16.0005
R3239 GNDA.n1253 GNDA.n1250 16.0005
R3240 GNDA.n1250 GNDA.n1249 16.0005
R3241 GNDA.n1249 GNDA.n1246 16.0005
R3242 GNDA.n1245 GNDA.n1242 16.0005
R3243 GNDA.n1242 GNDA.n1241 16.0005
R3244 GNDA.n1241 GNDA.n1238 16.0005
R3245 GNDA.n1238 GNDA.n1237 16.0005
R3246 GNDA.n1237 GNDA.n1234 16.0005
R3247 GNDA.n1234 GNDA.n1233 16.0005
R3248 GNDA.n1233 GNDA.n1230 16.0005
R3249 GNDA.n1230 GNDA.n1229 16.0005
R3250 GNDA.n623 GNDA.n622 16.0005
R3251 GNDA.n626 GNDA.n623 16.0005
R3252 GNDA.n627 GNDA.n626 16.0005
R3253 GNDA.n630 GNDA.n627 16.0005
R3254 GNDA.n631 GNDA.n630 16.0005
R3255 GNDA.n634 GNDA.n631 16.0005
R3256 GNDA.n635 GNDA.n634 16.0005
R3257 GNDA.n636 GNDA.n635 16.0005
R3258 GNDA.n619 GNDA.n618 16.0005
R3259 GNDA.n618 GNDA.n615 16.0005
R3260 GNDA.n615 GNDA.n614 16.0005
R3261 GNDA.n614 GNDA.n611 16.0005
R3262 GNDA.n611 GNDA.n610 16.0005
R3263 GNDA.n610 GNDA.n607 16.0005
R3264 GNDA.n607 GNDA.n606 16.0005
R3265 GNDA.n606 GNDA.n603 16.0005
R3266 GNDA.n602 GNDA.n599 16.0005
R3267 GNDA.n599 GNDA.n598 16.0005
R3268 GNDA.n598 GNDA.n595 16.0005
R3269 GNDA.n595 GNDA.n594 16.0005
R3270 GNDA.n594 GNDA.n591 16.0005
R3271 GNDA.n591 GNDA.n590 16.0005
R3272 GNDA.n590 GNDA.n587 16.0005
R3273 GNDA.n587 GNDA.n586 16.0005
R3274 GNDA.n950 GNDA.n949 16.0005
R3275 GNDA.n1668 GNDA.n950 16.0005
R3276 GNDA.n1522 GNDA.n1480 16.0005
R3277 GNDA.n1528 GNDA.n1480 16.0005
R3278 GNDA.n1529 GNDA.n1528 16.0005
R3279 GNDA.n1530 GNDA.n1529 16.0005
R3280 GNDA.n1530 GNDA.n1478 16.0005
R3281 GNDA.n1536 GNDA.n1478 16.0005
R3282 GNDA.n1537 GNDA.n1536 16.0005
R3283 GNDA.n1540 GNDA.n1537 16.0005
R3284 GNDA.n1521 GNDA.n1520 16.0005
R3285 GNDA.n1520 GNDA.n1482 16.0005
R3286 GNDA.n1514 GNDA.n1482 16.0005
R3287 GNDA.n1514 GNDA.n1513 16.0005
R3288 GNDA.n1513 GNDA.n1512 16.0005
R3289 GNDA.n1512 GNDA.n1484 16.0005
R3290 GNDA.n1506 GNDA.n1484 16.0005
R3291 GNDA.n1506 GNDA.n1505 16.0005
R3292 GNDA.n1504 GNDA.n1486 16.0005
R3293 GNDA.n1498 GNDA.n1486 16.0005
R3294 GNDA.n1498 GNDA.n1497 16.0005
R3295 GNDA.n1497 GNDA.n1496 16.0005
R3296 GNDA.n1496 GNDA.n1488 16.0005
R3297 GNDA.n1491 GNDA.n1488 16.0005
R3298 GNDA.n1491 GNDA.n1464 16.0005
R3299 GNDA.n1575 GNDA.n1464 16.0005
R3300 GNDA.n2011 GNDA.n2010 16.0005
R3301 GNDA.n2010 GNDA.n2007 16.0005
R3302 GNDA.n2007 GNDA.n2006 16.0005
R3303 GNDA.n2006 GNDA.n2003 16.0005
R3304 GNDA.n2003 GNDA.n2002 16.0005
R3305 GNDA.n2002 GNDA.n1999 16.0005
R3306 GNDA.n1999 GNDA.n1998 16.0005
R3307 GNDA.n1998 GNDA.n1996 16.0005
R3308 GNDA.n2015 GNDA.n2014 16.0005
R3309 GNDA.n2018 GNDA.n2015 16.0005
R3310 GNDA.n2019 GNDA.n2018 16.0005
R3311 GNDA.n2022 GNDA.n2019 16.0005
R3312 GNDA.n2023 GNDA.n2022 16.0005
R3313 GNDA.n2026 GNDA.n2023 16.0005
R3314 GNDA.n2027 GNDA.n2026 16.0005
R3315 GNDA.n2030 GNDA.n2027 16.0005
R3316 GNDA.n2034 GNDA.n2031 16.0005
R3317 GNDA.n2035 GNDA.n2034 16.0005
R3318 GNDA.n2038 GNDA.n2035 16.0005
R3319 GNDA.n2039 GNDA.n2038 16.0005
R3320 GNDA.n2042 GNDA.n2039 16.0005
R3321 GNDA.n2043 GNDA.n2042 16.0005
R3322 GNDA.n2046 GNDA.n2043 16.0005
R3323 GNDA.n2048 GNDA.n2046 16.0005
R3324 GNDA.n1083 GNDA.n1082 16.0005
R3325 GNDA.n1086 GNDA.n1083 16.0005
R3326 GNDA.n1087 GNDA.n1086 16.0005
R3327 GNDA.n1090 GNDA.n1087 16.0005
R3328 GNDA.n1091 GNDA.n1090 16.0005
R3329 GNDA.n1094 GNDA.n1091 16.0005
R3330 GNDA.n1096 GNDA.n1094 16.0005
R3331 GNDA.n1097 GNDA.n1096 16.0005
R3332 GNDA.n1079 GNDA.n1078 16.0005
R3333 GNDA.n1078 GNDA.n1075 16.0005
R3334 GNDA.n1075 GNDA.n1074 16.0005
R3335 GNDA.n1074 GNDA.n1071 16.0005
R3336 GNDA.n1071 GNDA.n1070 16.0005
R3337 GNDA.n1070 GNDA.n1067 16.0005
R3338 GNDA.n1067 GNDA.n1066 16.0005
R3339 GNDA.n1066 GNDA.n1063 16.0005
R3340 GNDA.n1062 GNDA.n1059 16.0005
R3341 GNDA.n1059 GNDA.n1058 16.0005
R3342 GNDA.n1058 GNDA.n1055 16.0005
R3343 GNDA.n1055 GNDA.n1054 16.0005
R3344 GNDA.n1054 GNDA.n1051 16.0005
R3345 GNDA.n1051 GNDA.n1050 16.0005
R3346 GNDA.n1050 GNDA.n1047 16.0005
R3347 GNDA.n1047 GNDA.n1023 16.0005
R3348 GNDA.t227 GNDA.n430 15.5368
R3349 GNDA.t227 GNDA.n428 15.5368
R3350 GNDA.t227 GNDA.n50 15.5368
R3351 GNDA.t217 GNDA.t44 15.4463
R3352 GNDA.t187 GNDA.t320 15.4463
R3353 GNDA.n197 GNDA.n196 15.1729
R3354 GNDA.n1881 GNDA.n422 14.555
R3355 GNDA.n1461 GNDA.n421 14.555
R3356 GNDA.n132 GNDA.n131 14.363
R3357 GNDA.n209 GNDA.n208 14.1651
R3358 GNDA.n153 GNDA.n152 14.0922
R3359 GNDA.n2169 GNDA.n2168 13.8005
R3360 GNDA.n2177 GNDA.n2176 13.8005
R3361 GNDA.n2183 GNDA.n2182 13.8005
R3362 GNDA.n2189 GNDA.n2188 13.8005
R3363 GNDA.n2240 GNDA.n2239 13.8005
R3364 GNDA.n2234 GNDA.n2233 12.7542
R3365 GNDA.n173 GNDA.t290 12.6791
R3366 GNDA.n182 GNDA.t278 12.6791
R3367 GNDA.n9 GNDA.t250 12.6791
R3368 GNDA.n29 GNDA.t242 12.6791
R3369 GNDA.n809 GNDA.t215 12.3572
R3370 GNDA.n398 GNDA.t193 12.3572
R3371 GNDA.t183 GNDA.n1993 12.3572
R3372 GNDA.n257 GNDA.n154 12.2505
R3373 GNDA.n2152 GNDA.n43 12.2193
R3374 GNDA.n1760 GNDA.n1759 11.6369
R3375 GNDA.n1759 GNDA.n1758 11.6369
R3376 GNDA.n1758 GNDA.n1757 11.6369
R3377 GNDA.n1757 GNDA.n1755 11.6369
R3378 GNDA.n1755 GNDA.n1752 11.6369
R3379 GNDA.n1752 GNDA.n1751 11.6369
R3380 GNDA.n1751 GNDA.n1748 11.6369
R3381 GNDA.n1748 GNDA.n1747 11.6369
R3382 GNDA.n1747 GNDA.n1744 11.6369
R3383 GNDA.n1744 GNDA.n652 11.6369
R3384 GNDA.n1743 GNDA.n1742 11.6369
R3385 GNDA.n1742 GNDA.n924 11.6369
R3386 GNDA.n1736 GNDA.n924 11.6369
R3387 GNDA.n1736 GNDA.n1735 11.6369
R3388 GNDA.n1735 GNDA.n1734 11.6369
R3389 GNDA.n1734 GNDA.n928 11.6369
R3390 GNDA.n1728 GNDA.n928 11.6369
R3391 GNDA.n1728 GNDA.n1727 11.6369
R3392 GNDA.n1727 GNDA.n1726 11.6369
R3393 GNDA.n1726 GNDA.n932 11.6369
R3394 GNDA.n1720 GNDA.n932 11.6369
R3395 GNDA.n1323 GNDA.n1322 11.6369
R3396 GNDA.n1326 GNDA.n1323 11.6369
R3397 GNDA.n1327 GNDA.n1326 11.6369
R3398 GNDA.n1330 GNDA.n1327 11.6369
R3399 GNDA.n1331 GNDA.n1330 11.6369
R3400 GNDA.n1334 GNDA.n1331 11.6369
R3401 GNDA.n1335 GNDA.n1334 11.6369
R3402 GNDA.n1338 GNDA.n1335 11.6369
R3403 GNDA.n1339 GNDA.n1338 11.6369
R3404 GNDA.n1342 GNDA.n1339 11.6369
R3405 GNDA.n1319 GNDA.n1318 11.6369
R3406 GNDA.n1318 GNDA.n1315 11.6369
R3407 GNDA.n1315 GNDA.n1314 11.6369
R3408 GNDA.n1314 GNDA.n1311 11.6369
R3409 GNDA.n1311 GNDA.n1310 11.6369
R3410 GNDA.n1310 GNDA.n1307 11.6369
R3411 GNDA.n1307 GNDA.n1306 11.6369
R3412 GNDA.n1306 GNDA.n1303 11.6369
R3413 GNDA.n1303 GNDA.n1302 11.6369
R3414 GNDA.n1302 GNDA.n455 11.6369
R3415 GNDA.n1976 GNDA.n455 11.6369
R3416 GNDA.n918 GNDA.n917 11.6369
R3417 GNDA.n917 GNDA.n916 11.6369
R3418 GNDA.n916 GNDA.n914 11.6369
R3419 GNDA.n914 GNDA.n911 11.6369
R3420 GNDA.n911 GNDA.n910 11.6369
R3421 GNDA.n910 GNDA.n907 11.6369
R3422 GNDA.n907 GNDA.n906 11.6369
R3423 GNDA.n906 GNDA.n903 11.6369
R3424 GNDA.n903 GNDA.n902 11.6369
R3425 GNDA.n902 GNDA.n899 11.6369
R3426 GNDA.n1893 GNDA.n456 11.6369
R3427 GNDA.n1896 GNDA.n1893 11.6369
R3428 GNDA.n1897 GNDA.n1896 11.6369
R3429 GNDA.n1900 GNDA.n1897 11.6369
R3430 GNDA.n1901 GNDA.n1900 11.6369
R3431 GNDA.n1904 GNDA.n1901 11.6369
R3432 GNDA.n1905 GNDA.n1904 11.6369
R3433 GNDA.n1908 GNDA.n1905 11.6369
R3434 GNDA.n1909 GNDA.n1908 11.6369
R3435 GNDA.n1912 GNDA.n1909 11.6369
R3436 GNDA.n1913 GNDA.n1912 11.6369
R3437 GNDA.n1143 GNDA.n509 11.6369
R3438 GNDA.n1146 GNDA.n1143 11.6369
R3439 GNDA.n1147 GNDA.n1146 11.6369
R3440 GNDA.n1150 GNDA.n1147 11.6369
R3441 GNDA.n1151 GNDA.n1150 11.6369
R3442 GNDA.n1154 GNDA.n1151 11.6369
R3443 GNDA.n1155 GNDA.n1154 11.6369
R3444 GNDA.n1158 GNDA.n1155 11.6369
R3445 GNDA.n1159 GNDA.n1158 11.6369
R3446 GNDA.n1162 GNDA.n1159 11.6369
R3447 GNDA.n1163 GNDA.n1162 11.6369
R3448 GNDA.n1602 GNDA.n1601 11.6369
R3449 GNDA.n1601 GNDA.n1600 11.6369
R3450 GNDA.n1600 GNDA.n1164 11.6369
R3451 GNDA.n1594 GNDA.n1164 11.6369
R3452 GNDA.n1594 GNDA.n1593 11.6369
R3453 GNDA.n1593 GNDA.n1592 11.6369
R3454 GNDA.n1592 GNDA.n1167 11.6369
R3455 GNDA.n1171 GNDA.n1167 11.6369
R3456 GNDA.n1585 GNDA.n1171 11.6369
R3457 GNDA.n1585 GNDA.n1584 11.6369
R3458 GNDA.n2104 GNDA.n115 11.6369
R3459 GNDA.n2104 GNDA.n2103 11.6369
R3460 GNDA.n2103 GNDA.n2102 11.6369
R3461 GNDA.n2102 GNDA.n117 11.6369
R3462 GNDA.n2097 GNDA.n117 11.6369
R3463 GNDA.n2097 GNDA.n2096 11.6369
R3464 GNDA.n2096 GNDA.n2095 11.6369
R3465 GNDA.n2095 GNDA.n120 11.6369
R3466 GNDA.n2090 GNDA.n120 11.6369
R3467 GNDA.n2090 GNDA.n2089 11.6369
R3468 GNDA.n2089 GNDA.n2088 11.6369
R3469 GNDA.n1982 GNDA.n123 11.6369
R3470 GNDA.n2081 GNDA.n1982 11.6369
R3471 GNDA.n2081 GNDA.n2080 11.6369
R3472 GNDA.n2080 GNDA.n2079 11.6369
R3473 GNDA.n2079 GNDA.n1983 11.6369
R3474 GNDA.n2074 GNDA.n1983 11.6369
R3475 GNDA.n2074 GNDA.n2073 11.6369
R3476 GNDA.n2073 GNDA.n2072 11.6369
R3477 GNDA.n2072 GNDA.n1985 11.6369
R3478 GNDA.n2066 GNDA.n1985 11.6369
R3479 GNDA.n1627 GNDA.n1626 11.6369
R3480 GNDA.n1626 GNDA.n1625 11.6369
R3481 GNDA.n1625 GNDA.n1015 11.6369
R3482 GNDA.n1619 GNDA.n1015 11.6369
R3483 GNDA.n1619 GNDA.n1618 11.6369
R3484 GNDA.n1618 GNDA.n1617 11.6369
R3485 GNDA.n1617 GNDA.n1018 11.6369
R3486 GNDA.n1022 GNDA.n1018 11.6369
R3487 GNDA.n1610 GNDA.n1022 11.6369
R3488 GNDA.n1610 GNDA.n1609 11.6369
R3489 GNDA.n1651 GNDA.n1650 11.6369
R3490 GNDA.n1650 GNDA.n1649 11.6369
R3491 GNDA.n1649 GNDA.n1003 11.6369
R3492 GNDA.n1643 GNDA.n1003 11.6369
R3493 GNDA.n1643 GNDA.n1642 11.6369
R3494 GNDA.n1642 GNDA.n1641 11.6369
R3495 GNDA.n1641 GNDA.n1007 11.6369
R3496 GNDA.n1635 GNDA.n1007 11.6369
R3497 GNDA.n1635 GNDA.n1634 11.6369
R3498 GNDA.n1634 GNDA.n1633 11.6369
R3499 GNDA.n1633 GNDA.n1011 11.6369
R3500 GNDA.n941 GNDA.n936 11.6369
R3501 GNDA.n1675 GNDA.n941 11.6369
R3502 GNDA.n1675 GNDA.n1674 11.6369
R3503 GNDA.n1674 GNDA.n1673 11.6369
R3504 GNDA.n1673 GNDA.n942 11.6369
R3505 GNDA.n1666 GNDA.n951 11.6369
R3506 GNDA.n955 GNDA.n951 11.6369
R3507 GNDA.n1659 GNDA.n955 11.6369
R3508 GNDA.n1659 GNDA.n1658 11.6369
R3509 GNDA.n1658 GNDA.n1657 11.6369
R3510 GNDA.n708 GNDA.n682 11.6369
R3511 GNDA.n708 GNDA.n707 11.6369
R3512 GNDA.n707 GNDA.n706 11.6369
R3513 GNDA.n706 GNDA.n685 11.6369
R3514 GNDA.n701 GNDA.n685 11.6369
R3515 GNDA.n701 GNDA.n700 11.6369
R3516 GNDA.n700 GNDA.n699 11.6369
R3517 GNDA.n699 GNDA.n688 11.6369
R3518 GNDA.n694 GNDA.n688 11.6369
R3519 GNDA.n694 GNDA.n693 11.6369
R3520 GNDA.n693 GNDA.n692 11.6369
R3521 GNDA.n768 GNDA.n767 11.6369
R3522 GNDA.n767 GNDA.n673 11.6369
R3523 GNDA.n762 GNDA.n673 11.6369
R3524 GNDA.n762 GNDA.n761 11.6369
R3525 GNDA.n761 GNDA.n760 11.6369
R3526 GNDA.n760 GNDA.n676 11.6369
R3527 GNDA.n755 GNDA.n676 11.6369
R3528 GNDA.n755 GNDA.n754 11.6369
R3529 GNDA.n754 GNDA.n753 11.6369
R3530 GNDA.n753 GNDA.n679 11.6369
R3531 GNDA.n748 GNDA.n679 11.6369
R3532 GNDA.n2239 GNDA.n2238 11.3792
R3533 GNDA.t57 GNDA.t113 10.7152
R3534 GNDA.n40 GNDA.n0 9.75668
R3535 GNDA.n417 GNDA.t168 9.6005
R3536 GNDA.n407 GNDA.t170 9.6005
R3537 GNDA.n2224 GNDA.t38 9.6005
R3538 GNDA.n45 GNDA.t169 9.6005
R3539 GNDA.n235 GNDA.t121 9.6005
R3540 GNDA.n235 GNDA.t272 9.6005
R3541 GNDA.n233 GNDA.t86 9.6005
R3542 GNDA.n233 GNDA.t118 9.6005
R3543 GNDA.n231 GNDA.t52 9.6005
R3544 GNDA.n231 GNDA.t70 9.6005
R3545 GNDA.n229 GNDA.t142 9.6005
R3546 GNDA.n229 GNDA.t61 9.6005
R3547 GNDA.n227 GNDA.t174 9.6005
R3548 GNDA.n227 GNDA.t99 9.6005
R3549 GNDA.n225 GNDA.t119 9.6005
R3550 GNDA.n225 GNDA.t34 9.6005
R3551 GNDA.n223 GNDA.t172 9.6005
R3552 GNDA.n223 GNDA.t97 9.6005
R3553 GNDA.n221 GNDA.t68 9.6005
R3554 GNDA.n221 GNDA.t32 9.6005
R3555 GNDA.n219 GNDA.t59 9.6005
R3556 GNDA.n219 GNDA.t50 9.6005
R3557 GNDA.n217 GNDA.t84 9.6005
R3558 GNDA.n217 GNDA.t123 9.6005
R3559 GNDA.n215 GNDA.t74 9.6005
R3560 GNDA.n215 GNDA.t140 9.6005
R3561 GNDA.n259 GNDA.n258 9.52967
R3562 GNDA.n246 GNDA.n245 9.52967
R3563 GNDA.t113 GNDA.t16 9.10801
R3564 GNDA.n187 GNDA.n158 9.0005
R3565 GNDA.n2249 GNDA.n2248 9.0005
R3566 GNDA.n2249 GNDA.n7 8.90675
R3567 GNDA.n1889 GNDA.n422 8.60107
R3568 GNDA.n1949 GNDA.n421 8.60107
R3569 GNDA.n808 GNDA.t189 8.23827
R3570 GNDA.t201 GNDA.n375 8.23827
R3571 GNDA.t195 GNDA.n2219 8.23827
R3572 GNDA.n42 GNDA.n41 7.56675
R3573 GNDA.n947 GNDA.n40 7.56675
R3574 GNDA.n2243 GNDA.n36 7.5008
R3575 GNDA.n8 GNDA.n7 7.46925
R3576 GNDA.n212 GNDA.n1 7.40675
R3577 GNDA.n826 GNDA.t131 7.20855
R3578 GNDA.n2196 GNDA.t78 7.20855
R3579 GNDA.t79 GNDA.n2058 7.20855
R3580 GNDA.n2242 GNDA.n37 7.20855
R3581 GNDA.n237 GNDA.n7 7.09425
R3582 GNDA.n214 GNDA.n212 7.03175
R3583 GNDA.n1720 GNDA.n1719 6.72373
R3584 GNDA.n1976 GNDA.n1975 6.72373
R3585 GNDA.n1913 GNDA.n1892 6.72373
R3586 GNDA.n1657 GNDA.n956 6.72373
R3587 GNDA.n692 GNDA.n114 6.72373
R3588 GNDA.n748 GNDA.n747 6.72373
R3589 GNDA.n2264 GNDA.n1 6.313
R3590 GNDA.n1975 GNDA.n456 6.20656
R3591 GNDA.n1892 GNDA.n509 6.20656
R3592 GNDA.n115 GNDA.n114 6.20656
R3593 GNDA.n1651 GNDA.n956 6.20656
R3594 GNDA.n1719 GNDA.n936 6.20656
R3595 GNDA.n747 GNDA.n682 6.20656
R3596 GNDA.t62 GNDA.t227 6.17883
R3597 GNDA.n1667 GNDA.n942 6.07727
R3598 GNDA.n418 GNDA.n408 5.81868
R3599 GNDA.n411 GNDA.n408 5.81868
R3600 GNDA.n42 GNDA.n0 5.737
R3601 GNDA.n1667 GNDA.n1666 5.5601
R3602 GNDA.n1814 GNDA.n1792 5.51161
R3603 GNDA.n1394 GNDA.n1372 5.51161
R3604 GNDA.n835 GNDA.n797 5.51161
R3605 GNDA.n319 GNDA.n100 5.51161
R3606 GNDA.n1229 GNDA.n1207 5.51161
R3607 GNDA.n586 GNDA.n557 5.51161
R3608 GNDA.n1576 GNDA.n1575 5.51161
R3609 GNDA.n2048 GNDA.n2047 5.51161
R3610 GNDA.n1135 GNDA.n1023 5.51161
R3611 GNDA.n154 GNDA.n153 5.5005
R3612 GNDA.n1583 GNDA.n1172 5.1717
R3613 GNDA.n2065 GNDA.n1990 5.1717
R3614 GNDA.n1608 GNDA.n1136 5.1717
R3615 GNDA.n399 GNDA.t227 5.14911
R3616 GNDA.t264 GNDA.t144 5.14911
R3617 GNDA.n248 GNDA.n246 5.063
R3618 GNDA.n2263 GNDA.n2262 5.02133
R3619 GNDA.n155 GNDA.n2 5.02133
R3620 GNDA.n187 GNDA.n186 5.0005
R3621 GNDA.n2250 GNDA.n2249 5.0005
R3622 GNDA.n181 GNDA.n180 4.91717
R3623 GNDA.n11 GNDA.n10 4.91717
R3624 GNDA.n28 GNDA.n27 4.91717
R3625 GNDA.n175 GNDA.n174 4.91717
R3626 GNDA.n1878 GNDA.n1766 4.9157
R3627 GNDA.n1458 GNDA.n1344 4.9157
R3628 GNDA.n898 GNDA.n897 4.9157
R3629 GNDA.n206 GNDA.n205 4.86508
R3630 GNDA.n194 GNDA.n193 4.86508
R3631 GNDA.n198 GNDA.n4 4.79217
R3632 GNDA.n2257 GNDA.n2256 4.79217
R3633 GNDA.n264 GNDA.t237 4.68943
R3634 GNDA.n263 GNDA.t73 4.68943
R3635 GNDA.n262 GNDA.t139 4.68943
R3636 GNDA.n261 GNDA.t83 4.68943
R3637 GNDA.n243 GNDA.t117 4.68943
R3638 GNDA.n242 GNDA.t120 4.68943
R3639 GNDA.n241 GNDA.t271 4.68943
R3640 GNDA.n258 GNDA.n257 4.5005
R3641 GNDA.n211 GNDA.n210 4.5005
R3642 GNDA.n214 GNDA.n213 4.5005
R3643 GNDA.n238 GNDA.n237 4.5005
R3644 GNDA.n1000 GNDA.n999 4.26717
R3645 GNDA.n999 GNDA.n998 4.26717
R3646 GNDA.n998 GNDA.n963 4.26717
R3647 GNDA.n992 GNDA.n963 4.26717
R3648 GNDA.n992 GNDA.n991 4.26717
R3649 GNDA.n991 GNDA.n990 4.26717
R3650 GNDA.n990 GNDA.n971 4.26717
R3651 GNDA.n978 GNDA.n971 4.26717
R3652 GNDA.n983 GNDA.n978 4.26717
R3653 GNDA.n983 GNDA.n982 4.26717
R3654 GNDA.n982 GNDA.n981 4.26717
R3655 GNDA.n1917 GNDA.n507 4.26717
R3656 GNDA.n1924 GNDA.n507 4.26717
R3657 GNDA.n1924 GNDA.n505 4.26717
R3658 GNDA.n505 GNDA.n502 4.26717
R3659 GNDA.n1931 GNDA.n502 4.26717
R3660 GNDA.n1931 GNDA.n500 4.26717
R3661 GNDA.n500 GNDA.n496 4.26717
R3662 GNDA.n1938 GNDA.n496 4.26717
R3663 GNDA.n1938 GNDA.n494 4.26717
R3664 GNDA.n494 GNDA.n493 4.26717
R3665 GNDA.n1945 GNDA.n493 4.26717
R3666 GNDA.n2110 GNDA.n112 4.26717
R3667 GNDA.n2116 GNDA.n112 4.26717
R3668 GNDA.n2116 GNDA.n110 4.26717
R3669 GNDA.n2122 GNDA.n110 4.26717
R3670 GNDA.n2122 GNDA.n108 4.26717
R3671 GNDA.n2128 GNDA.n108 4.26717
R3672 GNDA.n2128 GNDA.n106 4.26717
R3673 GNDA.n2134 GNDA.n106 4.26717
R3674 GNDA.n2134 GNDA.n104 4.26717
R3675 GNDA.n2141 GNDA.n104 4.26717
R3676 GNDA.n2141 GNDA.n102 4.26717
R3677 GNDA.n746 GNDA.n683 4.26717
R3678 GNDA.n741 GNDA.n683 4.26717
R3679 GNDA.n741 GNDA.n740 4.26717
R3680 GNDA.n740 GNDA.n718 4.26717
R3681 GNDA.n735 GNDA.n718 4.26717
R3682 GNDA.n735 GNDA.n734 4.26717
R3683 GNDA.n734 GNDA.n733 4.26717
R3684 GNDA.n733 GNDA.n728 4.26717
R3685 GNDA.n728 GNDA.n92 4.26717
R3686 GNDA.n2160 GNDA.n92 4.26717
R3687 GNDA.n2160 GNDA.n90 4.26717
R3688 GNDA.n1974 GNDA.n458 4.26717
R3689 GNDA.n1968 GNDA.n458 4.26717
R3690 GNDA.n1968 GNDA.n1967 4.26717
R3691 GNDA.n1967 GNDA.n1966 4.26717
R3692 GNDA.n1966 GNDA.n1964 4.26717
R3693 GNDA.n1964 GNDA.n1961 4.26717
R3694 GNDA.n1961 GNDA.n1960 4.26717
R3695 GNDA.n1960 GNDA.n1957 4.26717
R3696 GNDA.n1957 GNDA.n1956 4.26717
R3697 GNDA.n1956 GNDA.n1953 4.26717
R3698 GNDA.n1953 GNDA.n1952 4.26717
R3699 GNDA.n1718 GNDA.n937 4.26717
R3700 GNDA.n1712 GNDA.n937 4.26717
R3701 GNDA.n1712 GNDA.n1711 4.26717
R3702 GNDA.n1711 GNDA.n1710 4.26717
R3703 GNDA.n1710 GNDA.n1688 4.26717
R3704 GNDA.n1705 GNDA.n1688 4.26717
R3705 GNDA.n1705 GNDA.n1704 4.26717
R3706 GNDA.n1704 GNDA.n1703 4.26717
R3707 GNDA.n1703 GNDA.n1694 4.26717
R3708 GNDA.n1694 GNDA.n517 4.26717
R3709 GNDA.n1886 GNDA.n517 4.26717
R3710 GNDA.n209 GNDA.n206 4.2505
R3711 GNDA GNDA.n2265 4.2117
R3712 GNDA.t289 GNDA.t337 4.06704
R3713 GNDA.t137 GNDA.t277 4.06704
R3714 GNDA.n2260 GNDA.t33 4.06704
R3715 GNDA.t252 GNDA.n2259 4.06704
R3716 GNDA.t0 GNDA.n157 4.06704
R3717 GNDA.t63 GNDA.t249 4.06704
R3718 GNDA.t241 GNDA.t112 4.06704
R3719 GNDA.n2233 GNDA.n43 4.063
R3720 GNDA.n153 GNDA.n4 4.0005
R3721 GNDA.n1000 GNDA.n956 3.93531
R3722 GNDA.n1917 GNDA.n1892 3.93531
R3723 GNDA.n2110 GNDA.n114 3.93531
R3724 GNDA.n747 GNDA.n746 3.93531
R3725 GNDA.n1975 GNDA.n1974 3.93531
R3726 GNDA.n1719 GNDA.n1718 3.93531
R3727 GNDA.n8 GNDA.n2 3.90675
R3728 GNDA.n1876 GNDA.n1875 3.7893
R3729 GNDA.n1872 GNDA.n1769 3.7893
R3730 GNDA.n1871 GNDA.n1772 3.7893
R3731 GNDA.n1868 GNDA.n1867 3.7893
R3732 GNDA.n1794 GNDA.n1773 3.7893
R3733 GNDA.n1803 GNDA.n1802 3.7893
R3734 GNDA.n1806 GNDA.n1793 3.7893
R3735 GNDA.n1811 GNDA.n1807 3.7893
R3736 GNDA.n1456 GNDA.n1455 3.7893
R3737 GNDA.n1452 GNDA.n1347 3.7893
R3738 GNDA.n1451 GNDA.n1350 3.7893
R3739 GNDA.n1448 GNDA.n1447 3.7893
R3740 GNDA.n1374 GNDA.n1351 3.7893
R3741 GNDA.n1383 GNDA.n1382 3.7893
R3742 GNDA.n1386 GNDA.n1373 3.7893
R3743 GNDA.n1391 GNDA.n1387 3.7893
R3744 GNDA.n774 GNDA.n773 3.7893
R3745 GNDA.n891 GNDA.n890 3.7893
R3746 GNDA.n804 GNDA.n775 3.7893
R3747 GNDA.n805 GNDA.n803 3.7893
R3748 GNDA.n813 GNDA.n811 3.7893
R3749 GNDA.n822 GNDA.n821 3.7893
R3750 GNDA.n818 GNDA.n817 3.7893
R3751 GNDA.n832 GNDA.n798 3.7893
R3752 GNDA.n390 GNDA.n372 3.7893
R3753 GNDA.n389 GNDA.n373 3.7893
R3754 GNDA.n377 GNDA.n376 3.7893
R3755 GNDA.n383 GNDA.n382 3.7893
R3756 GNDA.n379 GNDA.n378 3.7893
R3757 GNDA.n307 GNDA.n284 3.7893
R3758 GNDA.n308 GNDA.n306 3.7893
R3759 GNDA.n316 GNDA.n314 3.7893
R3760 GNDA.n1292 GNDA.n1291 3.7893
R3761 GNDA.n1288 GNDA.n1184 3.7893
R3762 GNDA.n1287 GNDA.n1187 3.7893
R3763 GNDA.n1284 GNDA.n1283 3.7893
R3764 GNDA.n1209 GNDA.n1188 3.7893
R3765 GNDA.n1218 GNDA.n1217 3.7893
R3766 GNDA.n1221 GNDA.n1208 3.7893
R3767 GNDA.n1226 GNDA.n1222 3.7893
R3768 GNDA.n534 GNDA.n533 3.7893
R3769 GNDA.n642 GNDA.n641 3.7893
R3770 GNDA.n559 GNDA.n535 3.7893
R3771 GNDA.n563 GNDA.n561 3.7893
R3772 GNDA.n568 GNDA.n564 3.7893
R3773 GNDA.n575 GNDA.n574 3.7893
R3774 GNDA.n578 GNDA.n558 3.7893
R3775 GNDA.n583 GNDA.n579 3.7893
R3776 GNDA.n1538 GNDA.n1476 3.7893
R3777 GNDA.n1547 GNDA.n1546 3.7893
R3778 GNDA.n1473 GNDA.n1472 3.7893
R3779 GNDA.n1555 GNDA.n1553 3.7893
R3780 GNDA.n1554 GNDA.n1470 3.7893
R3781 GNDA.n1468 GNDA.n1467 3.7893
R3782 GNDA.n1570 GNDA.n1568 3.7893
R3783 GNDA.n1569 GNDA.n1463 3.7893
R3784 GNDA.n2211 GNDA.n74 3.7893
R3785 GNDA.n2210 GNDA.n75 3.7893
R3786 GNDA.n2198 GNDA.n2197 3.7893
R3787 GNDA.n2204 GNDA.n2203 3.7893
R3788 GNDA.n2200 GNDA.n2199 3.7893
R3789 GNDA.n1994 GNDA.n53 3.7893
R3790 GNDA.n2055 GNDA.n2054 3.7893
R3791 GNDA.n2052 GNDA.n2051 3.7893
R3792 GNDA.n1125 GNDA.n1100 3.7893
R3793 GNDA.n1124 GNDA.n1121 3.7893
R3794 GNDA.n1120 GNDA.n1101 3.7893
R3795 GNDA.n1117 GNDA.n1116 3.7893
R3796 GNDA.n1113 GNDA.n1102 3.7893
R3797 GNDA.n1106 GNDA.n1103 3.7893
R3798 GNDA.n1130 GNDA.n1025 3.7893
R3799 GNDA.n1131 GNDA.n1024 3.7893
R3800 GNDA.n1799 GNDA 3.7381
R3801 GNDA.n1379 GNDA 3.7381
R3802 GNDA.n816 GNDA 3.7381
R3803 GNDA GNDA.n395 3.7381
R3804 GNDA.n1214 GNDA 3.7381
R3805 GNDA.n571 GNDA 3.7381
R3806 GNDA GNDA.n1561 3.7381
R3807 GNDA GNDA.n2216 3.7381
R3808 GNDA GNDA.n1109 3.7381
R3809 GNDA.n201 GNDA.n195 3.65764
R3810 GNDA.n202 GNDA.n201 3.65764
R3811 GNDA.n189 GNDA.n3 3.65764
R3812 GNDA.n190 GNDA.n3 3.65764
R3813 GNDA.n212 GNDA.n211 3.53175
R3814 GNDA.n2238 GNDA.n40 3.51962
R3815 GNDA.n176 GNDA.t46 3.42907
R3816 GNDA.n176 GNDA.t152 3.42907
R3817 GNDA.n178 GNDA.t103 3.42907
R3818 GNDA.n178 GNDA.t10 3.42907
R3819 GNDA.n12 GNDA.t30 3.42907
R3820 GNDA.n12 GNDA.t101 3.42907
R3821 GNDA.n14 GNDA.t178 3.42907
R3822 GNDA.n14 GNDA.t26 3.42907
R3823 GNDA.n2262 GNDA.n2261 3.39217
R3824 GNDA.n156 GNDA.n155 3.39217
R3825 GNDA.n199 GNDA.n198 3.39217
R3826 GNDA.n2258 GNDA.n2257 3.39217
R3827 GNDA.n203 GNDA.n195 3.13621
R3828 GNDA.n203 GNDA.n202 3.13621
R3829 GNDA.n191 GNDA.n189 3.13621
R3830 GNDA.n191 GNDA.n190 3.13621
R3831 GNDA.n895 GNDA.n134 3.08966
R3832 GNDA.t21 GNDA.n893 3.08966
R3833 GNDA.n800 GNDA.t161 3.08966
R3834 GNDA.n829 GNDA.t23 3.08966
R3835 GNDA.n2208 GNDA.t156 3.08966
R3836 GNDA.n2226 GNDA.n44 2.86505
R3837 GNDA.n2227 GNDA.n2226 2.86505
R3838 GNDA.n2225 GNDA.n2221 2.86505
R3839 GNDA.n2222 GNDA.n2221 2.86505
R3840 GNDA.n2228 GNDA.n2227 2.86505
R3841 GNDA.n2223 GNDA.n2222 2.86505
R3842 GNDA.n2232 GNDA.n44 2.86505
R3843 GNDA.n2228 GNDA.n2225 2.86505
R3844 GNDA.n414 GNDA.n410 2.86505
R3845 GNDA.n415 GNDA.n414 2.86505
R3846 GNDA.n416 GNDA.n415 2.86505
R3847 GNDA.n411 GNDA.n410 2.86505
R3848 GNDA.n211 GNDA.n154 2.813
R3849 GNDA.n1878 GNDA.n1877 2.6629
R3850 GNDA.n1885 GNDA.n519 2.6629
R3851 GNDA.n1458 GNDA.n1457 2.6629
R3852 GNDA.n1371 GNDA.n484 2.6629
R3853 GNDA.n897 GNDA.n770 2.6629
R3854 GNDA.n796 GNDA.n795 2.6629
R3855 GNDA.n371 GNDA.n95 2.6629
R3856 GNDA.n2148 GNDA.n2147 2.6629
R3857 GNDA.n1183 GNDA.n1182 2.6629
R3858 GNDA.n1946 GNDA.n491 2.6629
R3859 GNDA.n1884 GNDA.n520 2.6629
R3860 GNDA.n556 GNDA.n510 2.6629
R3861 GNDA.n1539 GNDA.n492 2.6629
R3862 GNDA.n1995 GNDA.n101 2.6629
R3863 GNDA.n1099 GNDA.n1098 2.6629
R3864 GNDA.n1792 GNDA.n519 2.4581
R3865 GNDA.n1372 GNDA.n1371 2.4581
R3866 GNDA.n797 GNDA.n796 2.4581
R3867 GNDA.n795 GNDA.n95 2.4581
R3868 GNDA.n2148 GNDA.n100 2.4581
R3869 GNDA.n1182 GNDA.n484 2.4581
R3870 GNDA.n1207 GNDA.n491 2.4581
R3871 GNDA.n1885 GNDA.n1884 2.4581
R3872 GNDA.n557 GNDA.n556 2.4581
R3873 GNDA.n1946 GNDA.n492 2.4581
R3874 GNDA.n1576 GNDA.n1172 2.4581
R3875 GNDA.n2147 GNDA.n101 2.4581
R3876 GNDA.n2047 GNDA.n1990 2.4581
R3877 GNDA.n1098 GNDA.n510 2.4581
R3878 GNDA.n1136 GNDA.n1135 2.4581
R3879 GNDA.n2256 GNDA.n4 2.2505
R3880 GNDA.n213 GNDA.n150 2.19633
R3881 GNDA.n981 GNDA.n510 2.18124
R3882 GNDA.n1946 GNDA.n1945 2.18124
R3883 GNDA.n2147 GNDA.n102 2.18124
R3884 GNDA.n795 GNDA.n90 2.18124
R3885 GNDA.n1952 GNDA.n484 2.18124
R3886 GNDA.n1886 GNDA.n1885 2.18124
R3887 GNDA.n1810 GNDA.n1792 2.1509
R3888 GNDA.n1390 GNDA.n1372 2.1509
R3889 GNDA.n831 GNDA.n797 2.1509
R3890 GNDA.n315 GNDA.n100 2.1509
R3891 GNDA.n1225 GNDA.n1207 2.1509
R3892 GNDA.n582 GNDA.n557 2.1509
R3893 GNDA.n1577 GNDA.n1576 2.1509
R3894 GNDA.n2047 GNDA.n1992 2.1509
R3895 GNDA.n1135 GNDA.n1134 2.1509
R3896 GNDA.n1877 GNDA.n1767 2.13383
R3897 GNDA.n1457 GNDA.n1345 2.13383
R3898 GNDA.n885 GNDA.n770 2.13383
R3899 GNDA.n371 GNDA.n370 2.13383
R3900 GNDA.n1265 GNDA.n1183 2.13383
R3901 GNDA.n636 GNDA.n520 2.13383
R3902 GNDA.n1540 GNDA.n1539 2.13383
R3903 GNDA.n1996 GNDA.n1995 2.13383
R3904 GNDA.n1099 GNDA.n1097 2.13383
R3905 GNDA.n2234 GNDA 2.09787
R3906 GNDA.n182 GNDA.n181 2.09414
R3907 GNDA.n10 GNDA.n9 2.09414
R3908 GNDA.n29 GNDA.n28 2.09414
R3909 GNDA.n174 GNDA.n173 2.09414
R3910 GNDA.n1891 GNDA.n510 2.08643
R3911 GNDA.n1947 GNDA.n1946 2.08643
R3912 GNDA.n2147 GNDA.n2146 2.08643
R3913 GNDA.n795 GNDA.n89 2.08643
R3914 GNDA.n486 GNDA.n484 2.08643
R3915 GNDA.n1885 GNDA.n457 2.08643
R3916 GNDA.n829 GNDA.t280 2.05994
R3917 GNDA.n2154 GNDA.t310 2.05994
R3918 GNDA.n2150 GNDA.t255 2.05994
R3919 GNDA.n2193 GNDA.t264 2.05994
R3920 GNDA.n1877 GNDA.n1876 1.9461
R3921 GNDA.n1457 GNDA.n1456 1.9461
R3922 GNDA.n773 GNDA.n770 1.9461
R3923 GNDA.n372 GNDA.n371 1.9461
R3924 GNDA.n1292 GNDA.n1183 1.9461
R3925 GNDA.n533 GNDA.n520 1.9461
R3926 GNDA.n1539 GNDA.n1538 1.9461
R3927 GNDA.n1995 GNDA.n74 1.9461
R3928 GNDA.n1100 GNDA.n1099 1.9461
R3929 GNDA.n2263 GNDA.n2 1.938
R3930 GNDA.n186 GNDA.n185 1.93383
R3931 GNDA.n170 GNDA.n158 1.93383
R3932 GNDA.n2251 GNDA.n2250 1.93383
R3933 GNDA.n2248 GNDA.n2247 1.93383
R3934 GNDA.n239 GNDA.n238 1.91062
R3935 GNDA.n948 GNDA.n947 1.90675
R3936 GNDA.n403 GNDA.t167 1.83728
R3937 GNDA.n206 GNDA.n194 1.7505
R3938 GNDA.n180 GNDA.n1 1.563
R3939 GNDA.n1766 GNDA.n652 1.47392
R3940 GNDA.n1344 GNDA.n1342 1.47392
R3941 GNDA.n899 GNDA.n898 1.47392
R3942 GNDA.n1584 GNDA.n1583 1.47392
R3943 GNDA.n2066 GNDA.n2065 1.47392
R3944 GNDA.n1609 GNDA.n1608 1.47392
R3945 GNDA.n210 GNDA.n187 1.3755
R3946 GNDA.n27 GNDA.n15 1.1255
R3947 GNDA.n15 GNDA.n13 1.1255
R3948 GNDA.n13 GNDA.n11 1.1255
R3949 GNDA.n11 GNDA.n8 1.1255
R3950 GNDA.n180 GNDA.n179 1.1255
R3951 GNDA.n179 GNDA.n177 1.1255
R3952 GNDA.n177 GNDA.n175 1.1255
R3953 GNDA.n210 GNDA.n209 1.0005
R3954 GNDA.n2188 GNDA.n2183 0.96925
R3955 GNDA.n2176 GNDA.n2169 0.96925
R3956 GNDA.n1875 GNDA.n1769 0.8197
R3957 GNDA.n1872 GNDA.n1871 0.8197
R3958 GNDA.n1868 GNDA.n1772 0.8197
R3959 GNDA.n1867 GNDA.n1773 0.8197
R3960 GNDA.n1802 GNDA.n1799 0.8197
R3961 GNDA.n1803 GNDA.n1793 0.8197
R3962 GNDA.n1807 GNDA.n1806 0.8197
R3963 GNDA.n1811 GNDA.n1810 0.8197
R3964 GNDA.n1455 GNDA.n1347 0.8197
R3965 GNDA.n1452 GNDA.n1451 0.8197
R3966 GNDA.n1448 GNDA.n1350 0.8197
R3967 GNDA.n1447 GNDA.n1351 0.8197
R3968 GNDA.n1382 GNDA.n1379 0.8197
R3969 GNDA.n1383 GNDA.n1373 0.8197
R3970 GNDA.n1387 GNDA.n1386 0.8197
R3971 GNDA.n1391 GNDA.n1390 0.8197
R3972 GNDA.n891 GNDA.n774 0.8197
R3973 GNDA.n890 GNDA.n775 0.8197
R3974 GNDA.n805 GNDA.n804 0.8197
R3975 GNDA.n811 GNDA.n803 0.8197
R3976 GNDA.n822 GNDA.n816 0.8197
R3977 GNDA.n821 GNDA.n817 0.8197
R3978 GNDA.n818 GNDA.n798 0.8197
R3979 GNDA.n832 GNDA.n831 0.8197
R3980 GNDA.n390 GNDA.n389 0.8197
R3981 GNDA.n376 GNDA.n373 0.8197
R3982 GNDA.n383 GNDA.n377 0.8197
R3983 GNDA.n382 GNDA.n379 0.8197
R3984 GNDA.n395 GNDA.n284 0.8197
R3985 GNDA.n308 GNDA.n307 0.8197
R3986 GNDA.n314 GNDA.n306 0.8197
R3987 GNDA.n316 GNDA.n315 0.8197
R3988 GNDA.n1291 GNDA.n1184 0.8197
R3989 GNDA.n1288 GNDA.n1287 0.8197
R3990 GNDA.n1284 GNDA.n1187 0.8197
R3991 GNDA.n1283 GNDA.n1188 0.8197
R3992 GNDA.n1217 GNDA.n1214 0.8197
R3993 GNDA.n1218 GNDA.n1208 0.8197
R3994 GNDA.n1222 GNDA.n1221 0.8197
R3995 GNDA.n1226 GNDA.n1225 0.8197
R3996 GNDA.n642 GNDA.n534 0.8197
R3997 GNDA.n641 GNDA.n535 0.8197
R3998 GNDA.n561 GNDA.n559 0.8197
R3999 GNDA.n564 GNDA.n563 0.8197
R4000 GNDA.n574 GNDA.n571 0.8197
R4001 GNDA.n575 GNDA.n558 0.8197
R4002 GNDA.n579 GNDA.n578 0.8197
R4003 GNDA.n583 GNDA.n582 0.8197
R4004 GNDA.n1547 GNDA.n1476 0.8197
R4005 GNDA.n1546 GNDA.n1473 0.8197
R4006 GNDA.n1553 GNDA.n1472 0.8197
R4007 GNDA.n1555 GNDA.n1554 0.8197
R4008 GNDA.n1561 GNDA.n1468 0.8197
R4009 GNDA.n1568 GNDA.n1467 0.8197
R4010 GNDA.n1570 GNDA.n1569 0.8197
R4011 GNDA.n1577 GNDA.n1463 0.8197
R4012 GNDA.n2211 GNDA.n2210 0.8197
R4013 GNDA.n2197 GNDA.n75 0.8197
R4014 GNDA.n2204 GNDA.n2198 0.8197
R4015 GNDA.n2203 GNDA.n2200 0.8197
R4016 GNDA.n2216 GNDA.n53 0.8197
R4017 GNDA.n2055 GNDA.n1994 0.8197
R4018 GNDA.n2054 GNDA.n2052 0.8197
R4019 GNDA.n2051 GNDA.n1992 0.8197
R4020 GNDA.n1125 GNDA.n1124 0.8197
R4021 GNDA.n1121 GNDA.n1120 0.8197
R4022 GNDA.n1117 GNDA.n1101 0.8197
R4023 GNDA.n1116 GNDA.n1113 0.8197
R4024 GNDA.n1109 GNDA.n1106 0.8197
R4025 GNDA.n1103 GNDA.n1025 0.8197
R4026 GNDA.n1131 GNDA.n1130 0.8197
R4027 GNDA.n1134 GNDA.n1024 0.8197
R4028 GNDA.n2264 GNDA.n2263 0.6255
R4029 GNDA.n1763 GNDA.n403 0.575776
R4030 GNDA GNDA.n1794 0.5637
R4031 GNDA GNDA.n1374 0.5637
R4032 GNDA.n813 GNDA 0.5637
R4033 GNDA.n378 GNDA 0.5637
R4034 GNDA GNDA.n1209 0.5637
R4035 GNDA.n568 GNDA 0.5637
R4036 GNDA.n1470 GNDA 0.5637
R4037 GNDA.n2199 GNDA 0.5637
R4038 GNDA GNDA.n1102 0.5637
R4039 GNDA.n2239 GNDA.n39 0.563
R4040 GNDA.n2185 GNDA.n39 0.563
R4041 GNDA.n2187 GNDA.n2185 0.563
R4042 GNDA.n2188 GNDA.n2187 0.563
R4043 GNDA.n2183 GNDA.n79 0.563
R4044 GNDA.n2171 GNDA.n79 0.563
R4045 GNDA.n2173 GNDA.n2171 0.563
R4046 GNDA.n2175 GNDA.n2173 0.563
R4047 GNDA.n2176 GNDA.n2175 0.563
R4048 GNDA.n2169 GNDA.n87 0.563
R4049 GNDA.n129 GNDA.n87 0.563
R4050 GNDA.n131 GNDA.n129 0.563
R4051 GNDA.n250 GNDA.n248 0.563
R4052 GNDA.n252 GNDA.n250 0.563
R4053 GNDA.n254 GNDA.n252 0.563
R4054 GNDA.n256 GNDA.n254 0.563
R4055 GNDA.n257 GNDA.n256 0.563
R4056 GNDA.n216 GNDA.n214 0.563
R4057 GNDA.n218 GNDA.n216 0.563
R4058 GNDA.n220 GNDA.n218 0.563
R4059 GNDA.n222 GNDA.n220 0.563
R4060 GNDA.n224 GNDA.n222 0.563
R4061 GNDA.n226 GNDA.n224 0.563
R4062 GNDA.n228 GNDA.n226 0.563
R4063 GNDA.n230 GNDA.n228 0.563
R4064 GNDA.n232 GNDA.n230 0.563
R4065 GNDA.n234 GNDA.n232 0.563
R4066 GNDA.n236 GNDA.n234 0.563
R4067 GNDA.n20 GNDA.n18 0.563
R4068 GNDA.n22 GNDA.n20 0.563
R4069 GNDA.n24 GNDA.n22 0.563
R4070 GNDA.n26 GNDA.n24 0.563
R4071 GNDA.n163 GNDA.n161 0.563
R4072 GNDA.n165 GNDA.n163 0.563
R4073 GNDA.n167 GNDA.n165 0.563
R4074 GNDA.n169 GNDA.n167 0.563
R4075 GNDA.n2237 GNDA.n2234 0.276625
R4076 GNDA.n1797 GNDA 0.2565
R4077 GNDA.n1377 GNDA 0.2565
R4078 GNDA GNDA.n812 0.2565
R4079 GNDA.n396 GNDA 0.2565
R4080 GNDA.n1212 GNDA 0.2565
R4081 GNDA GNDA.n567 0.2565
R4082 GNDA.n1562 GNDA 0.2565
R4083 GNDA.n2217 GNDA 0.2565
R4084 GNDA.n1110 GNDA 0.2565
R4085 GNDA.n2238 GNDA.n2237 0.22375
R4086 GNDA.n237 GNDA.n236 0.21925
R4087 GNDA.n205 GNDA.n203 0.208833
R4088 GNDA.n193 GNDA.n191 0.208833
R4089 GNDA GNDA.n1797 0.0517
R4090 GNDA GNDA.n1377 0.0517
R4091 GNDA.n812 GNDA 0.0517
R4092 GNDA.n396 GNDA 0.0517
R4093 GNDA GNDA.n1212 0.0517
R4094 GNDA.n567 GNDA 0.0517
R4095 GNDA.n1562 GNDA 0.0517
R4096 GNDA.n2217 GNDA 0.0517
R4097 GNDA.n1110 GNDA 0.0517
R4098 VDDA.n129 VDDA.t319 1231.74
R4099 VDDA.n132 VDDA.t416 1231.74
R4100 VDDA.n48 VDDA.t349 1231.74
R4101 VDDA.n51 VDDA.t364 1231.74
R4102 VDDA.t359 VDDA.n114 1095.3
R4103 VDDA.n115 VDDA.t374 1095.3
R4104 VDDA.n75 VDDA.t420 1095.3
R4105 VDDA.t414 VDDA.n74 1095.3
R4106 VDDA.n34 VDDA.t362 1095.3
R4107 VDDA.t380 VDDA.n33 1095.3
R4108 VDDA.n212 VDDA.t393 708.125
R4109 VDDA.t393 VDDA.n168 708.125
R4110 VDDA.n189 VDDA.t333 708.125
R4111 VDDA.t333 VDDA.n171 708.125
R4112 VDDA.n234 VDDA.t432 676.966
R4113 VDDA.n86 VDDA.t340 672.293
R4114 VDDA.n89 VDDA.t410 672.293
R4115 VDDA.n5 VDDA.t385 672.293
R4116 VDDA.n8 VDDA.t334 672.293
R4117 VDDA.n114 VDDA.t360 663.801
R4118 VDDA.n115 VDDA.t375 663.801
R4119 VDDA.n75 VDDA.t421 663.801
R4120 VDDA.n74 VDDA.t415 663.801
R4121 VDDA.n34 VDDA.t363 663.801
R4122 VDDA.n33 VDDA.t381 663.801
R4123 VDDA.n147 VDDA.t428 661.375
R4124 VDDA.n150 VDDA.t346 661.375
R4125 VDDA.n191 VDDA.t356 660.001
R4126 VDDA.t392 VDDA.n213 657.76
R4127 VDDA.t332 VDDA.n190 657.76
R4128 VDDA.t426 VDDA.n311 645.231
R4129 VDDA.n312 VDDA.t398 645.231
R4130 VDDA.t371 VDDA.n280 643.038
R4131 VDDA.t389 VDDA.n233 643.038
R4132 VDDA.n281 VDDA.t368 643.038
R4133 VDDA.t338 VDDA.n319 643.037
R4134 VDDA.n320 VDDA.t423 643.037
R4135 VDDA.t404 VDDA.n297 643.037
R4136 VDDA.n298 VDDA.t326 643.037
R4137 VDDA.n54 VDDA.n53 599.342
R4138 VDDA.n56 VDDA.n55 599.342
R4139 VDDA.n58 VDDA.n57 599.342
R4140 VDDA.n60 VDDA.n59 599.342
R4141 VDDA.n62 VDDA.n61 599.342
R4142 VDDA.n64 VDDA.n63 599.342
R4143 VDDA.n66 VDDA.n65 599.342
R4144 VDDA.n68 VDDA.n67 599.342
R4145 VDDA.n70 VDDA.n69 599.342
R4146 VDDA.n72 VDDA.n71 599.342
R4147 VDDA.n107 VDDA.t343 589.076
R4148 VDDA.n110 VDDA.t328 589.076
R4149 VDDA.n26 VDDA.t382 589.076
R4150 VDDA.n29 VDDA.t394 589.076
R4151 VDDA.n259 VDDA.n227 587.407
R4152 VDDA.n255 VDDA.n254 587.407
R4153 VDDA.n272 VDDA.n271 587.407
R4154 VDDA.n266 VDDA.n221 587.407
R4155 VDDA.n271 VDDA.n270 585
R4156 VDDA.n269 VDDA.n266 585
R4157 VDDA.n257 VDDA.n227 585
R4158 VDDA.n256 VDDA.n255 585
R4159 VDDA.t107 VDDA.t359 580.557
R4160 VDDA.t440 VDDA.t107 580.557
R4161 VDDA.t209 VDDA.t440 580.557
R4162 VDDA.t17 VDDA.t209 580.557
R4163 VDDA.t92 VDDA.t17 580.557
R4164 VDDA.t441 VDDA.t92 580.557
R4165 VDDA.t210 VDDA.t441 580.557
R4166 VDDA.t100 VDDA.t210 580.557
R4167 VDDA.t99 VDDA.t100 580.557
R4168 VDDA.t127 VDDA.t99 580.557
R4169 VDDA.t374 VDDA.t127 580.557
R4170 VDDA.t420 VDDA.t11 580.557
R4171 VDDA.t11 VDDA.t108 580.557
R4172 VDDA.t108 VDDA.t450 580.557
R4173 VDDA.t450 VDDA.t15 580.557
R4174 VDDA.t15 VDDA.t13 580.557
R4175 VDDA.t13 VDDA.t243 580.557
R4176 VDDA.t243 VDDA.t123 580.557
R4177 VDDA.t123 VDDA.t245 580.557
R4178 VDDA.t245 VDDA.t105 580.557
R4179 VDDA.t105 VDDA.t446 580.557
R4180 VDDA.t446 VDDA.t172 580.557
R4181 VDDA.t172 VDDA.t205 580.557
R4182 VDDA.t205 VDDA.t27 580.557
R4183 VDDA.t27 VDDA.t448 580.557
R4184 VDDA.t448 VDDA.t139 580.557
R4185 VDDA.t139 VDDA.t193 580.557
R4186 VDDA.t193 VDDA.t29 580.557
R4187 VDDA.t29 VDDA.t3 580.557
R4188 VDDA.t3 VDDA.t247 580.557
R4189 VDDA.t247 VDDA.t236 580.557
R4190 VDDA.t236 VDDA.t414 580.557
R4191 VDDA.t362 VDDA.t208 580.557
R4192 VDDA.t208 VDDA.t186 580.557
R4193 VDDA.t186 VDDA.t442 580.557
R4194 VDDA.t442 VDDA.t207 580.557
R4195 VDDA.t207 VDDA.t439 580.557
R4196 VDDA.t439 VDDA.t1 580.557
R4197 VDDA.t1 VDDA.t204 580.557
R4198 VDDA.t204 VDDA.t112 580.557
R4199 VDDA.t112 VDDA.t438 580.557
R4200 VDDA.t438 VDDA.t48 580.557
R4201 VDDA.t48 VDDA.t380 580.557
R4202 VDDA.n214 VDDA.t377 540.818
R4203 VDDA.n139 VDDA.t406 456.526
R4204 VDDA.n142 VDDA.t400 456.526
R4205 VDDA.n279 VDDA.t370 419.108
R4206 VDDA.n282 VDDA.t367 419.108
R4207 VDDA.n232 VDDA.t388 413.084
R4208 VDDA.n235 VDDA.t431 413.084
R4209 VDDA.n318 VDDA.t337 409.067
R4210 VDDA.n321 VDDA.t422 409.067
R4211 VDDA.n310 VDDA.t425 409.067
R4212 VDDA.n313 VDDA.t397 409.067
R4213 VDDA.n296 VDDA.t403 409.067
R4214 VDDA.t65 VDDA.t392 407.144
R4215 VDDA.t6 VDDA.t65 407.144
R4216 VDDA.t141 VDDA.t6 407.144
R4217 VDDA.t162 VDDA.t141 407.144
R4218 VDDA.t160 VDDA.t162 407.144
R4219 VDDA.t166 VDDA.t160 407.144
R4220 VDDA.t93 VDDA.t166 407.144
R4221 VDDA.t110 VDDA.t93 407.144
R4222 VDDA.t269 VDDA.t110 407.144
R4223 VDDA.t241 VDDA.t269 407.144
R4224 VDDA.t271 VDDA.t241 407.144
R4225 VDDA.t153 VDDA.t271 407.144
R4226 VDDA.t168 VDDA.t153 407.144
R4227 VDDA.t170 VDDA.t168 407.144
R4228 VDDA.t239 VDDA.t170 407.144
R4229 VDDA.t202 VDDA.t239 407.144
R4230 VDDA.t267 VDDA.t202 407.144
R4231 VDDA.t67 VDDA.t267 407.144
R4232 VDDA.t377 VDDA.t67 407.144
R4233 VDDA.t251 VDDA.t332 407.144
R4234 VDDA.t59 VDDA.t251 407.144
R4235 VDDA.t452 VDDA.t59 407.144
R4236 VDDA.t261 VDDA.t452 407.144
R4237 VDDA.t460 VDDA.t261 407.144
R4238 VDDA.t265 VDDA.t460 407.144
R4239 VDDA.t255 VDDA.t265 407.144
R4240 VDDA.t95 VDDA.t255 407.144
R4241 VDDA.t176 VDDA.t95 407.144
R4242 VDDA.t18 VDDA.t176 407.144
R4243 VDDA.t259 VDDA.t18 407.144
R4244 VDDA.t249 VDDA.t259 407.144
R4245 VDDA.t253 VDDA.t249 407.144
R4246 VDDA.t155 VDDA.t253 407.144
R4247 VDDA.t101 VDDA.t155 407.144
R4248 VDDA.t41 VDDA.t101 407.144
R4249 VDDA.t263 VDDA.t41 407.144
R4250 VDDA.t257 VDDA.t263 407.144
R4251 VDDA.t356 VDDA.t257 407.144
R4252 VDDA.n141 VDDA.t401 397.784
R4253 VDDA.t407 VDDA.n140 397.784
R4254 VDDA.n299 VDDA.t325 390.322
R4255 VDDA.n212 VDDA.t391 379.582
R4256 VDDA.n189 VDDA.t331 379.582
R4257 VDDA.t376 VDDA.n215 379.277
R4258 VDDA.t37 VDDA.t371 373.214
R4259 VDDA.t103 VDDA.t37 373.214
R4260 VDDA.t368 VDDA.t103 373.214
R4261 VDDA.t238 VDDA.t389 373.214
R4262 VDDA.t5 VDDA.t238 373.214
R4263 VDDA.t432 VDDA.t5 373.214
R4264 VDDA.t39 VDDA.t338 373.214
R4265 VDDA.t158 VDDA.t39 373.214
R4266 VDDA.t23 VDDA.t158 373.214
R4267 VDDA.t125 VDDA.t23 373.214
R4268 VDDA.t423 VDDA.t125 373.214
R4269 VDDA.t458 VDDA.t426 373.214
R4270 VDDA.t215 VDDA.t458 373.214
R4271 VDDA.t130 VDDA.t215 373.214
R4272 VDDA.t464 VDDA.t130 373.214
R4273 VDDA.t213 VDDA.t464 373.214
R4274 VDDA.t63 VDDA.t213 373.214
R4275 VDDA.t128 VDDA.t63 373.214
R4276 VDDA.t200 VDDA.t128 373.214
R4277 VDDA.t184 VDDA.t200 373.214
R4278 VDDA.t151 VDDA.t184 373.214
R4279 VDDA.t398 VDDA.t151 373.214
R4280 VDDA.t25 VDDA.t404 373.214
R4281 VDDA.t164 VDDA.t25 373.214
R4282 VDDA.t97 VDDA.t164 373.214
R4283 VDDA.t61 VDDA.t97 373.214
R4284 VDDA.t326 VDDA.t61 373.214
R4285 VDDA.n252 VDDA.t352 360.868
R4286 VDDA.n277 VDDA.t322 360.868
R4287 VDDA.n216 VDDA.t376 358.858
R4288 VDDA.t391 VDDA.n211 358.858
R4289 VDDA.n192 VDDA.t355 358.858
R4290 VDDA.t331 VDDA.n188 358.858
R4291 VDDA.n311 VDDA.t427 354.154
R4292 VDDA.n312 VDDA.t399 354.154
R4293 VDDA.n191 VDDA.t357 354.065
R4294 VDDA.n281 VDDA.t369 354.065
R4295 VDDA.n280 VDDA.t372 354.063
R4296 VDDA.n233 VDDA.t390 354.063
R4297 VDDA.n167 VDDA.t378 351.793
R4298 VDDA.n73 VDDA.t413 348.325
R4299 VDDA.n76 VDDA.t419 348.325
R4300 VDDA.n113 VDDA.t358 348.075
R4301 VDDA.n116 VDDA.t373 348.075
R4302 VDDA.n32 VDDA.t379 348.075
R4303 VDDA.n35 VDDA.t361 348.075
R4304 VDDA.n234 VDDA.t433 347.224
R4305 VDDA.n293 VDDA.n292 345.127
R4306 VDDA.n295 VDDA.n294 345.127
R4307 VDDA.n289 VDDA.n288 344.7
R4308 VDDA.n316 VDDA.n315 344.7
R4309 VDDA.n109 VDDA.t329 343.882
R4310 VDDA.t344 VDDA.n108 343.882
R4311 VDDA.t383 VDDA.n27 343.882
R4312 VDDA.n28 VDDA.t395 343.882
R4313 VDDA.n165 VDDA.n164 341.675
R4314 VDDA.n195 VDDA.n194 341.675
R4315 VDDA.n197 VDDA.n196 341.675
R4316 VDDA.n199 VDDA.n198 341.675
R4317 VDDA.n201 VDDA.n200 341.675
R4318 VDDA.n203 VDDA.n202 341.675
R4319 VDDA.n205 VDDA.n204 341.675
R4320 VDDA.n207 VDDA.n206 341.675
R4321 VDDA.n209 VDDA.n208 341.675
R4322 VDDA.n170 VDDA.n169 341.675
R4323 VDDA.n173 VDDA.n172 341.675
R4324 VDDA.n175 VDDA.n174 341.675
R4325 VDDA.n177 VDDA.n176 341.675
R4326 VDDA.n179 VDDA.n178 341.675
R4327 VDDA.n181 VDDA.n180 341.675
R4328 VDDA.n183 VDDA.n182 341.675
R4329 VDDA.n185 VDDA.n184 341.675
R4330 VDDA.n187 VDDA.n186 341.675
R4331 VDDA.n291 VDDA.n290 339.272
R4332 VDDA.n302 VDDA.n301 339.272
R4333 VDDA.n304 VDDA.n303 339.272
R4334 VDDA.n306 VDDA.n305 339.272
R4335 VDDA.n308 VDDA.n307 339.272
R4336 VDDA.n285 VDDA.n284 334.772
R4337 VDDA.n297 VDDA.t405 332.267
R4338 VDDA.n298 VDDA.t327 332.267
R4339 VDDA.n319 VDDA.t339 332.084
R4340 VDDA.n320 VDDA.t424 332.084
R4341 VDDA.t401 VDDA.t174 259.091
R4342 VDDA.t174 VDDA.t407 259.091
R4343 VDDA.t78 VDDA.t353 251.471
R4344 VDDA.t231 VDDA.t78 251.471
R4345 VDDA.t434 VDDA.t231 251.471
R4346 VDDA.t188 VDDA.t434 251.471
R4347 VDDA.t50 VDDA.t188 251.471
R4348 VDDA.t119 VDDA.t50 251.471
R4349 VDDA.t74 VDDA.t119 251.471
R4350 VDDA.t121 VDDA.t74 251.471
R4351 VDDA.t52 VDDA.t121 251.471
R4352 VDDA.t76 VDDA.t52 251.471
R4353 VDDA.t54 VDDA.t76 251.471
R4354 VDDA.t56 VDDA.t54 251.471
R4355 VDDA.t146 VDDA.t56 251.471
R4356 VDDA.t227 VDDA.t146 251.471
R4357 VDDA.t116 VDDA.t227 251.471
R4358 VDDA.t222 VDDA.t116 251.471
R4359 VDDA.t323 VDDA.t222 251.471
R4360 VDDA.n273 VDDA.n272 243.698
R4361 VDDA.n215 VDDA.n214 238.367
R4362 VDDA.n214 VDDA.n166 238.367
R4363 VDDA.t353 VDDA.n261 237.5
R4364 VDDA.n274 VDDA.t323 237.5
R4365 VDDA.t329 VDDA.t31 217.708
R4366 VDDA.t31 VDDA.t44 217.708
R4367 VDDA.t44 VDDA.t90 217.708
R4368 VDDA.t90 VDDA.t91 217.708
R4369 VDDA.t91 VDDA.t219 217.708
R4370 VDDA.t219 VDDA.t132 217.708
R4371 VDDA.t132 VDDA.t137 217.708
R4372 VDDA.t137 VDDA.t133 217.708
R4373 VDDA.t133 VDDA.t218 217.708
R4374 VDDA.t218 VDDA.t8 217.708
R4375 VDDA.t8 VDDA.t344 217.708
R4376 VDDA.t454 VDDA.t383 217.708
R4377 VDDA.t192 VDDA.t454 217.708
R4378 VDDA.t457 VDDA.t192 217.708
R4379 VDDA.t178 VDDA.t457 217.708
R4380 VDDA.t181 VDDA.t178 217.708
R4381 VDDA.t198 VDDA.t181 217.708
R4382 VDDA.t466 VDDA.t198 217.708
R4383 VDDA.t0 VDDA.t466 217.708
R4384 VDDA.t456 VDDA.t0 217.708
R4385 VDDA.t197 VDDA.t456 217.708
R4386 VDDA.t395 VDDA.t197 217.708
R4387 VDDA.t429 VDDA.n148 213.131
R4388 VDDA.n149 VDDA.t347 213.131
R4389 VDDA.t341 VDDA.n87 213.131
R4390 VDDA.n88 VDDA.t411 213.131
R4391 VDDA.t386 VDDA.n6 213.131
R4392 VDDA.n7 VDDA.t335 213.131
R4393 VDDA.n260 VDDA.n259 190.333
R4394 VDDA.n265 VDDA.n264 185
R4395 VDDA.n270 VDDA.n263 185
R4396 VDDA.n274 VDDA.n263 185
R4397 VDDA.n269 VDDA.n268 185
R4398 VDDA.n267 VDDA.n222 185
R4399 VDDA.n276 VDDA.n275 185
R4400 VDDA.n275 VDDA.n274 185
R4401 VDDA.n261 VDDA.n260 185
R4402 VDDA.n258 VDDA.n226 185
R4403 VDDA.n257 VDDA.n228 185
R4404 VDDA.n256 VDDA.n229 185
R4405 VDDA.n231 VDDA.n230 185
R4406 VDDA.n253 VDDA.n225 185
R4407 VDDA.n261 VDDA.n225 185
R4408 VDDA.n220 VDDA.n219 168.435
R4409 VDDA.n238 VDDA.n237 168.435
R4410 VDDA.n240 VDDA.n239 168.435
R4411 VDDA.n242 VDDA.n241 168.435
R4412 VDDA.n244 VDDA.n243 168.435
R4413 VDDA.n246 VDDA.n245 168.435
R4414 VDDA.n248 VDDA.n247 168.435
R4415 VDDA.n250 VDDA.n249 168.435
R4416 VDDA.n141 VDDA.t402 168.139
R4417 VDDA.n140 VDDA.t409 168.139
R4418 VDDA.n138 VDDA.n137 153.576
R4419 VDDA.n264 VDDA.n263 150
R4420 VDDA.n268 VDDA.n263 150
R4421 VDDA.n275 VDDA.n222 150
R4422 VDDA.n260 VDDA.n226 150
R4423 VDDA.n229 VDDA.n228 150
R4424 VDDA.n230 VDDA.n225 150
R4425 VDDA.t279 VDDA.t429 146.155
R4426 VDDA.t347 VDDA.t279 146.155
R4427 VDDA.t291 VDDA.t341 146.155
R4428 VDDA.t299 VDDA.t291 146.155
R4429 VDDA.t295 VDDA.t299 146.155
R4430 VDDA.t301 VDDA.t295 146.155
R4431 VDDA.t277 VDDA.t301 146.155
R4432 VDDA.t285 VDDA.t277 146.155
R4433 VDDA.t293 VDDA.t285 146.155
R4434 VDDA.t287 VDDA.t293 146.155
R4435 VDDA.t297 VDDA.t287 146.155
R4436 VDDA.t303 VDDA.t297 146.155
R4437 VDDA.t411 VDDA.t303 146.155
R4438 VDDA.t309 VDDA.t386 146.155
R4439 VDDA.t305 VDDA.t309 146.155
R4440 VDDA.t311 VDDA.t305 146.155
R4441 VDDA.t273 VDDA.t311 146.155
R4442 VDDA.t281 VDDA.t273 146.155
R4443 VDDA.t289 VDDA.t281 146.155
R4444 VDDA.t283 VDDA.t289 146.155
R4445 VDDA.t307 VDDA.t283 146.155
R4446 VDDA.t313 VDDA.t307 146.155
R4447 VDDA.t275 VDDA.t313 146.155
R4448 VDDA.t335 VDDA.t275 146.155
R4449 VDDA.n109 VDDA.t330 136.701
R4450 VDDA.n108 VDDA.t345 136.701
R4451 VDDA.n27 VDDA.t384 136.701
R4452 VDDA.n28 VDDA.t396 136.701
R4453 VDDA.t354 VDDA.n227 123.126
R4454 VDDA.n255 VDDA.t354 123.126
R4455 VDDA.n271 VDDA.t324 123.126
R4456 VDDA.n266 VDDA.t324 123.126
R4457 VDDA.n131 VDDA.t417 122.829
R4458 VDDA.t320 VDDA.n130 122.829
R4459 VDDA.t350 VDDA.n49 122.829
R4460 VDDA.n50 VDDA.t365 122.829
R4461 VDDA.t417 VDDA.t82 81.6411
R4462 VDDA.t82 VDDA.t9 81.6411
R4463 VDDA.t9 VDDA.t84 81.6411
R4464 VDDA.t84 VDDA.t220 81.6411
R4465 VDDA.t220 VDDA.t134 81.6411
R4466 VDDA.t134 VDDA.t143 81.6411
R4467 VDDA.t143 VDDA.t87 81.6411
R4468 VDDA.t87 VDDA.t34 81.6411
R4469 VDDA.t34 VDDA.t46 81.6411
R4470 VDDA.t46 VDDA.t32 81.6411
R4471 VDDA.t32 VDDA.t320 81.6411
R4472 VDDA.t179 VDDA.t350 81.6411
R4473 VDDA.t195 VDDA.t179 81.6411
R4474 VDDA.t462 VDDA.t195 81.6411
R4475 VDDA.t72 VDDA.t462 81.6411
R4476 VDDA.t444 VDDA.t72 81.6411
R4477 VDDA.t225 VDDA.t444 81.6411
R4478 VDDA.t80 VDDA.t225 81.6411
R4479 VDDA.t211 VDDA.t80 81.6411
R4480 VDDA.t21 VDDA.t211 81.6411
R4481 VDDA.t182 VDDA.t21 81.6411
R4482 VDDA.t365 VDDA.t182 81.6411
R4483 VDDA.n53 VDDA.t12 78.8005
R4484 VDDA.n53 VDDA.t109 78.8005
R4485 VDDA.n55 VDDA.t451 78.8005
R4486 VDDA.n55 VDDA.t16 78.8005
R4487 VDDA.n57 VDDA.t14 78.8005
R4488 VDDA.n57 VDDA.t244 78.8005
R4489 VDDA.n59 VDDA.t124 78.8005
R4490 VDDA.n59 VDDA.t246 78.8005
R4491 VDDA.n61 VDDA.t106 78.8005
R4492 VDDA.n61 VDDA.t447 78.8005
R4493 VDDA.n63 VDDA.t173 78.8005
R4494 VDDA.n63 VDDA.t206 78.8005
R4495 VDDA.n65 VDDA.t28 78.8005
R4496 VDDA.n65 VDDA.t449 78.8005
R4497 VDDA.n67 VDDA.t140 78.8005
R4498 VDDA.n67 VDDA.t194 78.8005
R4499 VDDA.n69 VDDA.t30 78.8005
R4500 VDDA.n69 VDDA.t4 78.8005
R4501 VDDA.n71 VDDA.t248 78.8005
R4502 VDDA.n71 VDDA.t237 78.8005
R4503 VDDA.n148 VDDA.t430 76.2576
R4504 VDDA.n149 VDDA.t348 76.2576
R4505 VDDA.n87 VDDA.t342 76.2576
R4506 VDDA.n88 VDDA.t412 76.2576
R4507 VDDA.n6 VDDA.t387 76.2576
R4508 VDDA.n7 VDDA.t336 76.2576
R4509 VDDA.n83 VDDA.n82 71.513
R4510 VDDA.n85 VDDA.n84 71.513
R4511 VDDA.n91 VDDA.n90 71.513
R4512 VDDA.n93 VDDA.n92 71.513
R4513 VDDA.n2 VDDA.n1 71.513
R4514 VDDA.n4 VDDA.n3 71.513
R4515 VDDA.n10 VDDA.n9 71.513
R4516 VDDA.n12 VDDA.n11 71.513
R4517 VDDA.n146 VDDA.n145 71.388
R4518 VDDA.n95 VDDA.n81 67.013
R4519 VDDA.n14 VDDA.n0 67.013
R4520 VDDA.n274 VDDA.n273 65.8183
R4521 VDDA.n274 VDDA.n262 65.8183
R4522 VDDA.n261 VDDA.n223 65.8183
R4523 VDDA.n261 VDDA.n224 65.8183
R4524 VDDA.n161 VDDA.t471 59.5681
R4525 VDDA.n160 VDDA.t472 59.5681
R4526 VDDA.n268 VDDA.n262 53.3664
R4527 VDDA.n273 VDDA.n264 53.3664
R4528 VDDA.n262 VDDA.n222 53.3664
R4529 VDDA.n226 VDDA.n223 53.3664
R4530 VDDA.n229 VDDA.n224 53.3664
R4531 VDDA.n228 VDDA.n223 53.3664
R4532 VDDA.n230 VDDA.n224 53.3664
R4533 VDDA.n160 VDDA.t470 52.3888
R4534 VDDA.n162 VDDA.t469 48.9557
R4535 VDDA.n120 VDDA.n119 41.1393
R4536 VDDA.n122 VDDA.n121 41.1393
R4537 VDDA.n124 VDDA.n123 41.1393
R4538 VDDA.n126 VDDA.n125 41.1393
R4539 VDDA.n128 VDDA.n127 41.1393
R4540 VDDA.n39 VDDA.n38 41.1393
R4541 VDDA.n41 VDDA.n40 41.1393
R4542 VDDA.n43 VDDA.n42 41.1393
R4543 VDDA.n45 VDDA.n44 41.1393
R4544 VDDA.n47 VDDA.n46 41.1393
R4545 VDDA.n131 VDDA.t418 40.9789
R4546 VDDA.n130 VDDA.t321 40.9789
R4547 VDDA.n49 VDDA.t351 40.9789
R4548 VDDA.n50 VDDA.t366 40.9789
R4549 VDDA.n164 VDDA.t268 39.4005
R4550 VDDA.n164 VDDA.t68 39.4005
R4551 VDDA.n194 VDDA.t240 39.4005
R4552 VDDA.n194 VDDA.t203 39.4005
R4553 VDDA.n196 VDDA.t169 39.4005
R4554 VDDA.n196 VDDA.t171 39.4005
R4555 VDDA.n198 VDDA.t272 39.4005
R4556 VDDA.n198 VDDA.t154 39.4005
R4557 VDDA.n200 VDDA.t270 39.4005
R4558 VDDA.n200 VDDA.t242 39.4005
R4559 VDDA.n202 VDDA.t94 39.4005
R4560 VDDA.n202 VDDA.t111 39.4005
R4561 VDDA.n204 VDDA.t161 39.4005
R4562 VDDA.n204 VDDA.t167 39.4005
R4563 VDDA.n206 VDDA.t142 39.4005
R4564 VDDA.n206 VDDA.t163 39.4005
R4565 VDDA.n208 VDDA.t66 39.4005
R4566 VDDA.n208 VDDA.t7 39.4005
R4567 VDDA.n169 VDDA.t264 39.4005
R4568 VDDA.n169 VDDA.t258 39.4005
R4569 VDDA.n172 VDDA.t102 39.4005
R4570 VDDA.n172 VDDA.t42 39.4005
R4571 VDDA.n174 VDDA.t254 39.4005
R4572 VDDA.n174 VDDA.t156 39.4005
R4573 VDDA.n176 VDDA.t260 39.4005
R4574 VDDA.n176 VDDA.t250 39.4005
R4575 VDDA.n178 VDDA.t177 39.4005
R4576 VDDA.n178 VDDA.t19 39.4005
R4577 VDDA.n180 VDDA.t256 39.4005
R4578 VDDA.n180 VDDA.t96 39.4005
R4579 VDDA.n182 VDDA.t461 39.4005
R4580 VDDA.n182 VDDA.t266 39.4005
R4581 VDDA.n184 VDDA.t453 39.4005
R4582 VDDA.n184 VDDA.t262 39.4005
R4583 VDDA.n186 VDDA.t252 39.4005
R4584 VDDA.n186 VDDA.t60 39.4005
R4585 VDDA.n284 VDDA.t38 39.4005
R4586 VDDA.n284 VDDA.t104 39.4005
R4587 VDDA.n288 VDDA.t24 39.4005
R4588 VDDA.n288 VDDA.t126 39.4005
R4589 VDDA.n315 VDDA.t40 39.4005
R4590 VDDA.n315 VDDA.t159 39.4005
R4591 VDDA.n290 VDDA.t185 39.4005
R4592 VDDA.n290 VDDA.t152 39.4005
R4593 VDDA.n301 VDDA.t129 39.4005
R4594 VDDA.n301 VDDA.t201 39.4005
R4595 VDDA.n303 VDDA.t214 39.4005
R4596 VDDA.n303 VDDA.t64 39.4005
R4597 VDDA.n305 VDDA.t131 39.4005
R4598 VDDA.n305 VDDA.t465 39.4005
R4599 VDDA.n307 VDDA.t459 39.4005
R4600 VDDA.n307 VDDA.t216 39.4005
R4601 VDDA.n292 VDDA.t98 39.4005
R4602 VDDA.n292 VDDA.t62 39.4005
R4603 VDDA.n294 VDDA.t26 39.4005
R4604 VDDA.n294 VDDA.t165 39.4005
R4605 VDDA.n98 VDDA.n96 30.2255
R4606 VDDA.n17 VDDA.n15 30.2255
R4607 VDDA.n106 VDDA.n105 29.663
R4608 VDDA.n104 VDDA.n103 29.663
R4609 VDDA.n102 VDDA.n101 29.663
R4610 VDDA.n100 VDDA.n99 29.663
R4611 VDDA.n98 VDDA.n97 29.663
R4612 VDDA.n25 VDDA.n24 29.663
R4613 VDDA.n23 VDDA.n22 29.663
R4614 VDDA.n21 VDDA.n20 29.663
R4615 VDDA.n19 VDDA.n18 29.663
R4616 VDDA.n17 VDDA.n16 29.663
R4617 VDDA.n159 VDDA.n153 27.9413
R4618 VDDA.n321 VDDA.n320 27.2462
R4619 VDDA.n319 VDDA.n318 27.2462
R4620 VDDA.n299 VDDA.n298 27.2462
R4621 VDDA.n297 VDDA.n296 27.2462
R4622 VDDA.n280 VDDA.n279 25.087
R4623 VDDA.n282 VDDA.n281 25.087
R4624 VDDA.n313 VDDA.n312 25.0384
R4625 VDDA.n311 VDDA.n310 25.0384
R4626 VDDA.n233 VDDA.n232 22.9536
R4627 VDDA.n192 VDDA.n191 22.9536
R4628 VDDA.n277 VDDA.n276 22.8576
R4629 VDDA.n253 VDDA.n252 22.8576
R4630 VDDA.n137 VDDA.t175 21.8894
R4631 VDDA.n137 VDDA.t408 21.8894
R4632 VDDA.n216 VDDA.n166 20.7243
R4633 VDDA.n211 VDDA.n168 20.7243
R4634 VDDA.n188 VDDA.n171 20.7243
R4635 VDDA.n235 VDDA.n234 20.4312
R4636 VDDA.n153 VDDA.n152 20.1017
R4637 VDDA.n159 VDDA.t149 19.9244
R4638 VDDA.n236 VDDA.n232 15.488
R4639 VDDA.n188 VDDA.n187 14.6963
R4640 VDDA.n283 VDDA.n282 14.363
R4641 VDDA.n283 VDDA.n279 14.363
R4642 VDDA.n296 VDDA.n295 14.363
R4643 VDDA.n236 VDDA.n235 14.238
R4644 VDDA.n211 VDDA.n210 14.0713
R4645 VDDA.n217 VDDA.n216 14.0713
R4646 VDDA.n193 VDDA.n192 14.0713
R4647 VDDA.n252 VDDA.n251 13.8005
R4648 VDDA.n278 VDDA.n277 13.8005
R4649 VDDA.n318 VDDA.n317 13.8005
R4650 VDDA.n310 VDDA.n309 13.8005
R4651 VDDA.n300 VDDA.n299 13.8005
R4652 VDDA.n314 VDDA.n313 13.8005
R4653 VDDA.n322 VDDA.n321 13.8005
R4654 VDDA.n219 VDDA.t117 13.1338
R4655 VDDA.n219 VDDA.t223 13.1338
R4656 VDDA.n237 VDDA.t147 13.1338
R4657 VDDA.n237 VDDA.t228 13.1338
R4658 VDDA.n239 VDDA.t55 13.1338
R4659 VDDA.n239 VDDA.t57 13.1338
R4660 VDDA.n241 VDDA.t53 13.1338
R4661 VDDA.n241 VDDA.t77 13.1338
R4662 VDDA.n243 VDDA.t75 13.1338
R4663 VDDA.n243 VDDA.t122 13.1338
R4664 VDDA.n245 VDDA.t51 13.1338
R4665 VDDA.n245 VDDA.t120 13.1338
R4666 VDDA.n247 VDDA.t435 13.1338
R4667 VDDA.n247 VDDA.t189 13.1338
R4668 VDDA.n249 VDDA.t79 13.1338
R4669 VDDA.n249 VDDA.t232 13.1338
R4670 VDDA.n323 VDDA.n322 11.4105
R4671 VDDA.n112 VDDA.n106 11.3443
R4672 VDDA.n31 VDDA.n25 11.3443
R4673 VDDA.t430 VDDA.n146 11.2576
R4674 VDDA.n146 VDDA.t280 11.2576
R4675 VDDA.n82 VDDA.t296 11.2576
R4676 VDDA.n82 VDDA.t302 11.2576
R4677 VDDA.n84 VDDA.t292 11.2576
R4678 VDDA.n84 VDDA.t300 11.2576
R4679 VDDA.n90 VDDA.t298 11.2576
R4680 VDDA.n90 VDDA.t304 11.2576
R4681 VDDA.n92 VDDA.t294 11.2576
R4682 VDDA.n92 VDDA.t288 11.2576
R4683 VDDA.n81 VDDA.t278 11.2576
R4684 VDDA.n81 VDDA.t286 11.2576
R4685 VDDA.n1 VDDA.t312 11.2576
R4686 VDDA.n1 VDDA.t274 11.2576
R4687 VDDA.n3 VDDA.t310 11.2576
R4688 VDDA.n3 VDDA.t306 11.2576
R4689 VDDA.n9 VDDA.t314 11.2576
R4690 VDDA.n9 VDDA.t276 11.2576
R4691 VDDA.n11 VDDA.t284 11.2576
R4692 VDDA.n11 VDDA.t308 11.2576
R4693 VDDA.n0 VDDA.t282 11.2576
R4694 VDDA.n0 VDDA.t290 11.2576
R4695 VDDA.n163 VDDA.n162 11.1572
R4696 VDDA.n287 VDDA.n286 9.7855
R4697 VDDA.n116 VDDA.n115 9.5505
R4698 VDDA.n114 VDDA.n113 9.5505
R4699 VDDA.n35 VDDA.n34 9.5505
R4700 VDDA.n33 VDDA.n32 9.5505
R4701 VDDA.n135 VDDA.n134 9.5005
R4702 VDDA.n80 VDDA.n79 9.5005
R4703 VDDA.n76 VDDA.n75 9.3005
R4704 VDDA.n74 VDDA.n73 9.3005
R4705 VDDA.n270 VDDA.n265 9.14336
R4706 VDDA.n270 VDDA.n269 9.14336
R4707 VDDA.n269 VDDA.n267 9.14336
R4708 VDDA.n258 VDDA.n257 9.14336
R4709 VDDA.n257 VDDA.n256 9.14336
R4710 VDDA.n256 VDDA.n231 9.14336
R4711 VDDA.n117 VDDA.n113 9.02133
R4712 VDDA.n36 VDDA.n32 9.02133
R4713 VDDA.n218 VDDA.n217 8.973
R4714 VDDA.n111 VDDA.n107 8.79217
R4715 VDDA.n30 VDDA.n26 8.79217
R4716 VDDA.n105 VDDA.t315 8.0005
R4717 VDDA.n105 VDDA.t86 8.0005
R4718 VDDA.n103 VDDA.t145 8.0005
R4719 VDDA.n103 VDDA.t45 8.0005
R4720 VDDA.n101 VDDA.t36 8.0005
R4721 VDDA.n101 VDDA.t217 8.0005
R4722 VDDA.n99 VDDA.t43 8.0005
R4723 VDDA.n99 VDDA.t89 8.0005
R4724 VDDA.n97 VDDA.t2 8.0005
R4725 VDDA.n97 VDDA.t136 8.0005
R4726 VDDA.n96 VDDA.t138 8.0005
R4727 VDDA.n96 VDDA.t316 8.0005
R4728 VDDA.n24 VDDA.t191 8.0005
R4729 VDDA.n24 VDDA.t318 8.0005
R4730 VDDA.n22 VDDA.t468 8.0005
R4731 VDDA.n22 VDDA.t150 8.0005
R4732 VDDA.n20 VDDA.t443 8.0005
R4733 VDDA.n20 VDDA.t157 8.0005
R4734 VDDA.n18 VDDA.t20 8.0005
R4735 VDDA.n18 VDDA.t455 8.0005
R4736 VDDA.n16 VDDA.t235 8.0005
R4737 VDDA.n16 VDDA.t199 8.0005
R4738 VDDA.n15 VDDA.t317 8.0005
R4739 VDDA.n15 VDDA.t467 8.0005
R4740 VDDA.n135 VDDA.n95 7.71925
R4741 VDDA.n80 VDDA.n14 7.71925
R4742 VDDA.n136 VDDA.n80 6.90675
R4743 VDDA.n136 VDDA.n135 6.8755
R4744 VDDA.n144 VDDA.n136 6.813
R4745 VDDA.n119 VDDA.t83 6.56717
R4746 VDDA.n119 VDDA.t10 6.56717
R4747 VDDA.n121 VDDA.t85 6.56717
R4748 VDDA.n121 VDDA.t221 6.56717
R4749 VDDA.n123 VDDA.t135 6.56717
R4750 VDDA.n123 VDDA.t144 6.56717
R4751 VDDA.n125 VDDA.t88 6.56717
R4752 VDDA.n125 VDDA.t35 6.56717
R4753 VDDA.n127 VDDA.t47 6.56717
R4754 VDDA.n127 VDDA.t33 6.56717
R4755 VDDA.n38 VDDA.t22 6.56717
R4756 VDDA.n38 VDDA.t183 6.56717
R4757 VDDA.n40 VDDA.t81 6.56717
R4758 VDDA.n40 VDDA.t212 6.56717
R4759 VDDA.n42 VDDA.t445 6.56717
R4760 VDDA.n42 VDDA.t226 6.56717
R4761 VDDA.n44 VDDA.t463 6.56717
R4762 VDDA.n44 VDDA.t73 6.56717
R4763 VDDA.n46 VDDA.t180 6.56717
R4764 VDDA.n46 VDDA.t196 6.56717
R4765 VDDA.n91 VDDA.n89 6.10467
R4766 VDDA.n86 VDDA.n85 6.10467
R4767 VDDA.n10 VDDA.n8 6.10467
R4768 VDDA.n5 VDDA.n4 6.10467
R4769 VDDA.n37 VDDA.n36 6.09425
R4770 VDDA.n118 VDDA.n117 6.063
R4771 VDDA.n73 VDDA.n72 5.60467
R4772 VDDA.n276 VDDA.n221 5.33286
R4773 VDDA.n254 VDDA.n253 5.33286
R4774 VDDA.n129 VDDA.n128 5.313
R4775 VDDA.n48 VDDA.n47 5.313
R4776 VDDA.n152 VDDA.n151 5.28175
R4777 VDDA.n144 VDDA.n143 5.28175
R4778 VDDA.n134 VDDA.n133 5.28175
R4779 VDDA.n112 VDDA.n111 5.28175
R4780 VDDA.n31 VDDA.n30 5.28175
R4781 VDDA.n77 VDDA.n76 5.04217
R4782 VDDA.n117 VDDA.n116 5.02133
R4783 VDDA.n36 VDDA.n35 5.02133
R4784 VDDA.n286 VDDA.n285 5.0005
R4785 VDDA.n111 VDDA.n110 4.79217
R4786 VDDA.n30 VDDA.n29 4.79217
R4787 VDDA.n147 VDDA.n145 4.7505
R4788 VDDA.n139 VDDA.n138 4.7505
R4789 VDDA.n133 VDDA.n132 4.7505
R4790 VDDA.n52 VDDA.n51 4.7505
R4791 VDDA.n163 VDDA.n159 4.5595
R4792 VDDA.n167 VDDA.n166 4.54311
R4793 VDDA.n215 VDDA.n167 4.54311
R4794 VDDA.n151 VDDA.n150 4.5005
R4795 VDDA.n143 VDDA.n142 4.5005
R4796 VDDA.n95 VDDA.n94 4.5005
R4797 VDDA.n79 VDDA.n78 4.5005
R4798 VDDA.n14 VDDA.n13 4.5005
R4799 VDDA.n285 VDDA.n283 4.5005
R4800 VDDA.n213 VDDA.n168 4.48641
R4801 VDDA.n213 VDDA.n212 4.48641
R4802 VDDA.n190 VDDA.n171 4.48641
R4803 VDDA.n190 VDDA.n189 4.48641
R4804 VDDA.n161 VDDA.n160 4.12334
R4805 VDDA.n134 VDDA.n118 3.84425
R4806 VDDA.n79 VDDA.n37 3.84425
R4807 VDDA.n272 VDDA.n265 3.75335
R4808 VDDA.n267 VDDA.n221 3.75335
R4809 VDDA.n259 VDDA.n258 3.75335
R4810 VDDA.n254 VDDA.n231 3.75335
R4811 VDDA.n324 VDDA.n323 3.71013
R4812 VDDA.n162 VDDA.n161 3.43377
R4813 VDDA.n78 VDDA.n77 3.1255
R4814 VDDA.n142 VDDA.n141 2.8255
R4815 VDDA.n140 VDDA.n139 2.8255
R4816 VDDA.n286 VDDA.n278 2.5005
R4817 VDDA.n110 VDDA.n109 2.423
R4818 VDDA.n108 VDDA.n107 2.423
R4819 VDDA.n29 VDDA.n28 2.423
R4820 VDDA.n27 VDDA.n26 2.423
R4821 VDDA.n324 VDDA.n153 2.1343
R4822 VDDA VDDA.n324 2.0779
R4823 VDDA.n132 VDDA.n131 1.97758
R4824 VDDA.n130 VDDA.n129 1.97758
R4825 VDDA.n51 VDDA.n50 1.97758
R4826 VDDA.n49 VDDA.n48 1.97758
R4827 VDDA.n150 VDDA.n149 1.888
R4828 VDDA.n148 VDDA.n147 1.888
R4829 VDDA.n210 VDDA.n193 1.8755
R4830 VDDA.n251 VDDA.n236 1.84425
R4831 VDDA.n309 VDDA.n300 1.813
R4832 VDDA.n317 VDDA.n314 1.813
R4833 VDDA.n118 VDDA.n112 1.438
R4834 VDDA.n37 VDDA.n31 1.438
R4835 VDDA.n89 VDDA.n88 1.03383
R4836 VDDA.n87 VDDA.n86 1.03383
R4837 VDDA.n8 VDDA.n7 1.03383
R4838 VDDA.n6 VDDA.n5 1.03383
R4839 VDDA.n251 VDDA.n250 1.0005
R4840 VDDA.n250 VDDA.n248 1.0005
R4841 VDDA.n248 VDDA.n246 1.0005
R4842 VDDA.n246 VDDA.n244 1.0005
R4843 VDDA.n244 VDDA.n242 1.0005
R4844 VDDA.n242 VDDA.n240 1.0005
R4845 VDDA.n240 VDDA.n238 1.0005
R4846 VDDA.n238 VDDA.n220 1.0005
R4847 VDDA.n278 VDDA.n220 1.0005
R4848 VDDA.n152 VDDA.n144 0.938
R4849 VDDA.n218 VDDA.n163 0.840625
R4850 VDDA.n78 VDDA.n52 0.78175
R4851 VDDA.n287 VDDA.n218 0.74075
R4852 VDDA.n151 VDDA.n145 0.6255
R4853 VDDA.n143 VDDA.n138 0.6255
R4854 VDDA.n94 VDDA.n93 0.6255
R4855 VDDA.n93 VDDA.n91 0.6255
R4856 VDDA.n85 VDDA.n83 0.6255
R4857 VDDA.n94 VDDA.n83 0.6255
R4858 VDDA.n13 VDDA.n12 0.6255
R4859 VDDA.n12 VDDA.n10 0.6255
R4860 VDDA.n4 VDDA.n2 0.6255
R4861 VDDA.n13 VDDA.n2 0.6255
R4862 VDDA.n187 VDDA.n185 0.6255
R4863 VDDA.n185 VDDA.n183 0.6255
R4864 VDDA.n183 VDDA.n181 0.6255
R4865 VDDA.n181 VDDA.n179 0.6255
R4866 VDDA.n179 VDDA.n177 0.6255
R4867 VDDA.n177 VDDA.n175 0.6255
R4868 VDDA.n175 VDDA.n173 0.6255
R4869 VDDA.n173 VDDA.n170 0.6255
R4870 VDDA.n193 VDDA.n170 0.6255
R4871 VDDA.n210 VDDA.n209 0.6255
R4872 VDDA.n209 VDDA.n207 0.6255
R4873 VDDA.n207 VDDA.n205 0.6255
R4874 VDDA.n205 VDDA.n203 0.6255
R4875 VDDA.n203 VDDA.n201 0.6255
R4876 VDDA.n201 VDDA.n199 0.6255
R4877 VDDA.n199 VDDA.n197 0.6255
R4878 VDDA.n197 VDDA.n195 0.6255
R4879 VDDA.n195 VDDA.n165 0.6255
R4880 VDDA.n217 VDDA.n165 0.6255
R4881 VDDA.n128 VDDA.n126 0.563
R4882 VDDA.n126 VDDA.n124 0.563
R4883 VDDA.n124 VDDA.n122 0.563
R4884 VDDA.n122 VDDA.n120 0.563
R4885 VDDA.n133 VDDA.n120 0.563
R4886 VDDA.n100 VDDA.n98 0.563
R4887 VDDA.n102 VDDA.n100 0.563
R4888 VDDA.n104 VDDA.n102 0.563
R4889 VDDA.n106 VDDA.n104 0.563
R4890 VDDA.n72 VDDA.n70 0.563
R4891 VDDA.n70 VDDA.n68 0.563
R4892 VDDA.n68 VDDA.n66 0.563
R4893 VDDA.n66 VDDA.n64 0.563
R4894 VDDA.n64 VDDA.n62 0.563
R4895 VDDA.n62 VDDA.n60 0.563
R4896 VDDA.n60 VDDA.n58 0.563
R4897 VDDA.n58 VDDA.n56 0.563
R4898 VDDA.n56 VDDA.n54 0.563
R4899 VDDA.n77 VDDA.n54 0.563
R4900 VDDA.n47 VDDA.n45 0.563
R4901 VDDA.n45 VDDA.n43 0.563
R4902 VDDA.n43 VDDA.n41 0.563
R4903 VDDA.n41 VDDA.n39 0.563
R4904 VDDA.n52 VDDA.n39 0.563
R4905 VDDA.n19 VDDA.n17 0.563
R4906 VDDA.n21 VDDA.n19 0.563
R4907 VDDA.n23 VDDA.n21 0.563
R4908 VDDA.n25 VDDA.n23 0.563
R4909 VDDA.n295 VDDA.n293 0.563
R4910 VDDA.n300 VDDA.n293 0.563
R4911 VDDA.n309 VDDA.n308 0.563
R4912 VDDA.n308 VDDA.n306 0.563
R4913 VDDA.n306 VDDA.n304 0.563
R4914 VDDA.n304 VDDA.n302 0.563
R4915 VDDA.n302 VDDA.n291 0.563
R4916 VDDA.n314 VDDA.n291 0.563
R4917 VDDA.n317 VDDA.n316 0.563
R4918 VDDA.n316 VDDA.n289 0.563
R4919 VDDA.n322 VDDA.n289 0.563
R4920 VDDA VDDA.n287 0.41175
R4921 VDDA.t190 VDDA.t148 0.1603
R4922 VDDA.t115 VDDA.t58 0.1603
R4923 VDDA.t224 VDDA.t69 0.1603
R4924 VDDA.t118 VDDA.t437 0.1603
R4925 VDDA.t230 VDDA.t233 0.1603
R4926 VDDA.n155 VDDA.t234 0.159278
R4927 VDDA.n156 VDDA.t113 0.159278
R4928 VDDA.n157 VDDA.t71 0.159278
R4929 VDDA.n158 VDDA.t436 0.159278
R4930 VDDA.n158 VDDA.t229 0.1368
R4931 VDDA.n158 VDDA.t190 0.1368
R4932 VDDA.n157 VDDA.t70 0.1368
R4933 VDDA.n157 VDDA.t115 0.1368
R4934 VDDA.n156 VDDA.t49 0.1368
R4935 VDDA.n156 VDDA.t224 0.1368
R4936 VDDA.n155 VDDA.t187 0.1368
R4937 VDDA.n155 VDDA.t118 0.1368
R4938 VDDA.n154 VDDA.t114 0.1368
R4939 VDDA.n154 VDDA.t230 0.1368
R4940 VDDA.n323 VDDA 0.135625
R4941 VDDA.t234 VDDA.n154 0.00152174
R4942 VDDA.t113 VDDA.n155 0.00152174
R4943 VDDA.t71 VDDA.n156 0.00152174
R4944 VDDA.t436 VDDA.n157 0.00152174
R4945 VDDA.t149 VDDA.n158 0.00152174
R4946 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 369.534
R4947 bgr_0.V_TOP.n23 bgr_0.V_TOP.n21 339.961
R4948 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 339.272
R4949 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 339.272
R4950 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 339.272
R4951 bgr_0.V_TOP.n29 bgr_0.V_TOP.n28 339.272
R4952 bgr_0.V_TOP.n24 bgr_0.V_TOP.n20 334.772
R4953 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 224.934
R4954 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 224.934
R4955 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 224.934
R4956 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 224.934
R4957 bgr_0.V_TOP.n35 bgr_0.V_TOP.n34 224.934
R4958 bgr_0.V_TOP.n34 bgr_0.V_TOP.n33 224.934
R4959 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 224.934
R4960 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R4961 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R4962 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R4963 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R4964 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R4965 bgr_0.V_TOP bgr_0.V_TOP.t48 214.222
R4966 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 163.175
R4967 bgr_0.V_TOP.n39 bgr_0.V_TOP.t24 144.601
R4968 bgr_0.V_TOP.n38 bgr_0.V_TOP.t33 144.601
R4969 bgr_0.V_TOP.n37 bgr_0.V_TOP.t39 144.601
R4970 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 144.601
R4971 bgr_0.V_TOP.n35 bgr_0.V_TOP.t15 144.601
R4972 bgr_0.V_TOP.n34 bgr_0.V_TOP.t28 144.601
R4973 bgr_0.V_TOP.n33 bgr_0.V_TOP.t38 144.601
R4974 bgr_0.V_TOP.n32 bgr_0.V_TOP.t14 144.601
R4975 bgr_0.V_TOP.n0 bgr_0.V_TOP.t30 144.601
R4976 bgr_0.V_TOP.n1 bgr_0.V_TOP.t18 144.601
R4977 bgr_0.V_TOP.n2 bgr_0.V_TOP.t46 144.601
R4978 bgr_0.V_TOP.n3 bgr_0.V_TOP.t37 144.601
R4979 bgr_0.V_TOP.n4 bgr_0.V_TOP.t26 144.601
R4980 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R4981 bgr_0.V_TOP.n17 bgr_0.V_TOP.t1 108.424
R4982 bgr_0.V_TOP.n30 bgr_0.V_TOP.t9 95.4467
R4983 bgr_0.V_TOP bgr_0.V_TOP.n39 69.6227
R4984 bgr_0.V_TOP.n32 bgr_0.V_TOP.n31 69.6227
R4985 bgr_0.V_TOP.n31 bgr_0.V_TOP.n5 69.6227
R4986 bgr_0.V_TOP.n18 bgr_0.V_TOP.t10 39.4005
R4987 bgr_0.V_TOP.n18 bgr_0.V_TOP.t4 39.4005
R4988 bgr_0.V_TOP.n20 bgr_0.V_TOP.t8 39.4005
R4989 bgr_0.V_TOP.n20 bgr_0.V_TOP.t6 39.4005
R4990 bgr_0.V_TOP.n22 bgr_0.V_TOP.t0 39.4005
R4991 bgr_0.V_TOP.n22 bgr_0.V_TOP.t13 39.4005
R4992 bgr_0.V_TOP.n21 bgr_0.V_TOP.t12 39.4005
R4993 bgr_0.V_TOP.n21 bgr_0.V_TOP.t2 39.4005
R4994 bgr_0.V_TOP.n26 bgr_0.V_TOP.t3 39.4005
R4995 bgr_0.V_TOP.n26 bgr_0.V_TOP.t5 39.4005
R4996 bgr_0.V_TOP.n28 bgr_0.V_TOP.t7 39.4005
R4997 bgr_0.V_TOP.n28 bgr_0.V_TOP.t11 39.4005
R4998 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 37.1479
R4999 bgr_0.V_TOP.n19 bgr_0.V_TOP.n17 27.8371
R5000 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 8.313
R5001 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 5.188
R5002 bgr_0.V_TOP.n6 bgr_0.V_TOP.t31 4.8295
R5003 bgr_0.V_TOP.n7 bgr_0.V_TOP.t22 4.8295
R5004 bgr_0.V_TOP.n8 bgr_0.V_TOP.t20 4.8295
R5005 bgr_0.V_TOP.n9 bgr_0.V_TOP.t45 4.8295
R5006 bgr_0.V_TOP.n10 bgr_0.V_TOP.t42 4.8295
R5007 bgr_0.V_TOP.n11 bgr_0.V_TOP.t36 4.8295
R5008 bgr_0.V_TOP.n12 bgr_0.V_TOP.t17 4.8295
R5009 bgr_0.V_TOP.n13 bgr_0.V_TOP.t43 4.8295
R5010 bgr_0.V_TOP.n14 bgr_0.V_TOP.t34 4.8295
R5011 bgr_0.V_TOP.n6 bgr_0.V_TOP.t35 4.5005
R5012 bgr_0.V_TOP.n7 bgr_0.V_TOP.t32 4.5005
R5013 bgr_0.V_TOP.n8 bgr_0.V_TOP.t25 4.5005
R5014 bgr_0.V_TOP.n9 bgr_0.V_TOP.t21 4.5005
R5015 bgr_0.V_TOP.n10 bgr_0.V_TOP.t49 4.5005
R5016 bgr_0.V_TOP.n11 bgr_0.V_TOP.t44 4.5005
R5017 bgr_0.V_TOP.n12 bgr_0.V_TOP.t23 4.5005
R5018 bgr_0.V_TOP.n13 bgr_0.V_TOP.t19 4.5005
R5019 bgr_0.V_TOP.n16 bgr_0.V_TOP.t40 4.5005
R5020 bgr_0.V_TOP.n15 bgr_0.V_TOP.t47 4.5005
R5021 bgr_0.V_TOP.n14 bgr_0.V_TOP.t41 4.5005
R5022 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 4.5005
R5023 bgr_0.V_TOP.n29 bgr_0.V_TOP.n27 2.1255
R5024 bgr_0.V_TOP.n27 bgr_0.V_TOP.n25 2.1255
R5025 bgr_0.V_TOP.n25 bgr_0.V_TOP.n19 2.1255
R5026 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 0.3295
R5027 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R5028 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 0.3295
R5029 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 0.3295
R5030 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 0.3295
R5031 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 0.3295
R5032 bgr_0.V_TOP.n9 bgr_0.V_TOP.n7 0.2825
R5033 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 0.2825
R5034 bgr_0.V_TOP.n13 bgr_0.V_TOP.n11 0.2825
R5035 bgr_0.V_TOP.n14 bgr_0.V_TOP.n13 0.2825
R5036 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n15 594.301
R5037 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n16 594.301
R5038 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n19 594.301
R5039 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t20 289.2
R5040 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t4 289.2
R5041 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n3 194.3
R5042 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n24 194.3
R5043 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n1 194.3
R5044 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n5 176.733
R5045 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n6 176.733
R5046 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n9 176.733
R5047 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n10 176.733
R5048 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n11 176.733
R5049 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n1 161.3
R5050 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n14 161.3
R5051 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t10 112.468
R5052 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t8 112.468
R5053 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t21 112.468
R5054 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t18 112.468
R5055 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t6 112.468
R5056 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t17 112.468
R5057 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t19 112.468
R5058 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t12 112.468
R5059 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t0 78.8005
R5060 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t3 78.8005
R5061 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t2 78.8005
R5062 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t16 78.8005
R5063 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t1 78.8005
R5064 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t15 78.8005
R5065 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t14 48.0005
R5066 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t5 48.0005
R5067 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t7 48.0005
R5068 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t11 48.0005
R5069 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t9 48.0005
R5070 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n26 48.0005
R5071 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n13 45.5227
R5072 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n7 45.5227
R5073 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n8 45.5227
R5074 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n12 45.5227
R5075 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n2 6.39633
R5076 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n0 6.39633
R5077 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n4 6.39633
R5078 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n20 6.10467
R5079 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n17 6.10467
R5080 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n23 5.97967
R5081 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n18 5.91717
R5082 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n17 5.91717
R5083 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n25 5.14633
R5084 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n21 4.85467
R5085 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n4 4.72967
R5086 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n1 4.72967
R5087 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n0 4.66717
R5088 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n22 1.2505
R5089 two_stage_opamp_dummy_magic_21_0.err_amp_out.n10 two_stage_opamp_dummy_magic_21_0.err_amp_out.t12 840.595
R5090 two_stage_opamp_dummy_magic_21_0.err_amp_out.n2 two_stage_opamp_dummy_magic_21_0.err_amp_out.n0 601.051
R5091 two_stage_opamp_dummy_magic_21_0.err_amp_out two_stage_opamp_dummy_magic_21_0.err_amp_out.n3 599.801
R5092 two_stage_opamp_dummy_magic_21_0.err_amp_out.n2 two_stage_opamp_dummy_magic_21_0.err_amp_out.n1 599.801
R5093 two_stage_opamp_dummy_magic_21_0.err_amp_out.n12 two_stage_opamp_dummy_magic_21_0.err_amp_out.n11 194.3
R5094 two_stage_opamp_dummy_magic_21_0.err_amp_out.n6 two_stage_opamp_dummy_magic_21_0.err_amp_out.n5 194.3
R5095 two_stage_opamp_dummy_magic_21_0.err_amp_out.n8 two_stage_opamp_dummy_magic_21_0.err_amp_out.n7 194.3
R5096 two_stage_opamp_dummy_magic_21_0.err_amp_out.n3 two_stage_opamp_dummy_magic_21_0.err_amp_out.t0 78.8005
R5097 two_stage_opamp_dummy_magic_21_0.err_amp_out.n3 two_stage_opamp_dummy_magic_21_0.err_amp_out.t10 78.8005
R5098 two_stage_opamp_dummy_magic_21_0.err_amp_out.n1 two_stage_opamp_dummy_magic_21_0.err_amp_out.t1 78.8005
R5099 two_stage_opamp_dummy_magic_21_0.err_amp_out.n1 two_stage_opamp_dummy_magic_21_0.err_amp_out.t11 78.8005
R5100 two_stage_opamp_dummy_magic_21_0.err_amp_out.n0 two_stage_opamp_dummy_magic_21_0.err_amp_out.t9 78.8005
R5101 two_stage_opamp_dummy_magic_21_0.err_amp_out.n0 two_stage_opamp_dummy_magic_21_0.err_amp_out.t2 78.8005
R5102 two_stage_opamp_dummy_magic_21_0.err_amp_out.n11 two_stage_opamp_dummy_magic_21_0.err_amp_out.t6 48.0005
R5103 two_stage_opamp_dummy_magic_21_0.err_amp_out.n11 two_stage_opamp_dummy_magic_21_0.err_amp_out.t3 48.0005
R5104 two_stage_opamp_dummy_magic_21_0.err_amp_out.n5 two_stage_opamp_dummy_magic_21_0.err_amp_out.t4 48.0005
R5105 two_stage_opamp_dummy_magic_21_0.err_amp_out.n5 two_stage_opamp_dummy_magic_21_0.err_amp_out.t8 48.0005
R5106 two_stage_opamp_dummy_magic_21_0.err_amp_out.n7 two_stage_opamp_dummy_magic_21_0.err_amp_out.t5 48.0005
R5107 two_stage_opamp_dummy_magic_21_0.err_amp_out.n7 two_stage_opamp_dummy_magic_21_0.err_amp_out.t7 48.0005
R5108 two_stage_opamp_dummy_magic_21_0.err_amp_out.n9 two_stage_opamp_dummy_magic_21_0.err_amp_out.n6 6.20883
R5109 two_stage_opamp_dummy_magic_21_0.err_amp_out.n6 two_stage_opamp_dummy_magic_21_0.err_amp_out.n4 6.20883
R5110 two_stage_opamp_dummy_magic_21_0.err_amp_out.n8 two_stage_opamp_dummy_magic_21_0.err_amp_out.n4 4.95883
R5111 two_stage_opamp_dummy_magic_21_0.err_amp_out.n13 two_stage_opamp_dummy_magic_21_0.err_amp_out.n12 4.95883
R5112 two_stage_opamp_dummy_magic_21_0.err_amp_out.n12 two_stage_opamp_dummy_magic_21_0.err_amp_out.n10 4.95883
R5113 two_stage_opamp_dummy_magic_21_0.err_amp_out.n9 two_stage_opamp_dummy_magic_21_0.err_amp_out.n8 4.95883
R5114 two_stage_opamp_dummy_magic_21_0.err_amp_out.n13 two_stage_opamp_dummy_magic_21_0.err_amp_out.n4 1.2505
R5115 two_stage_opamp_dummy_magic_21_0.err_amp_out two_stage_opamp_dummy_magic_21_0.err_amp_out.n2 1.2505
R5116 two_stage_opamp_dummy_magic_21_0.err_amp_out.n10 two_stage_opamp_dummy_magic_21_0.err_amp_out.n9 1.2505
R5117 two_stage_opamp_dummy_magic_21_0.err_amp_out two_stage_opamp_dummy_magic_21_0.err_amp_out.n13 1.063
R5118 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t12 610.534
R5119 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t14 610.534
R5120 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t30 433.8
R5121 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t21 433.8
R5122 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t27 433.8
R5123 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t17 433.8
R5124 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t25 433.8
R5125 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t15 433.8
R5126 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t23 433.8
R5127 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t29 433.8
R5128 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t19 433.8
R5129 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t31 433.8
R5130 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t22 433.8
R5131 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t28 433.8
R5132 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t18 433.8
R5133 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t26 433.8
R5134 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t16 433.8
R5135 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t24 433.8
R5136 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t13 433.8
R5137 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t20 433.8
R5138 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n0 339.836
R5139 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n1 339.834
R5140 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n2 339.272
R5141 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n5 287.264
R5142 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n24 176.733
R5143 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n23 176.733
R5144 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n22 176.733
R5145 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n21 176.733
R5146 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n20 176.733
R5147 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n19 176.733
R5148 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n18 176.733
R5149 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n17 176.733
R5150 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n8 176.733
R5151 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n9 176.733
R5152 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n10 176.733
R5153 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n11 176.733
R5154 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n12 176.733
R5155 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n13 176.733
R5156 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n14 176.733
R5157 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n15 176.733
R5158 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n26 162.508
R5159 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n25 56.2338
R5160 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n16 56.2338
R5161 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n4 52.01
R5162 two_stage_opamp_dummy_magic_21_0.V_tail_gate two_stage_opamp_dummy_magic_21_0.V_tail_gate.n6 51.6642
R5163 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n7 50.5797
R5164 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n28 49.3505
R5165 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t11 39.4005
R5166 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t6 39.4005
R5167 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t1 39.4005
R5168 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t2 39.4005
R5169 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t5 39.4005
R5170 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t4 39.4005
R5171 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t7 39.4005
R5172 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t3 39.4005
R5173 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t9 16.0005
R5174 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t8 16.0005
R5175 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t0 16.0005
R5176 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t10 16.0005
R5177 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n27 10.7922
R5178 two_stage_opamp_dummy_magic_21_0.V_tail_gate two_stage_opamp_dummy_magic_21_0.V_tail_gate.n29 1.04217
R5179 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n3 0.563
R5180 two_stage_opamp_dummy_magic_21_0.V_p_mir.n1 two_stage_opamp_dummy_magic_21_0.V_p_mir.n0 97.1193
R5181 two_stage_opamp_dummy_magic_21_0.V_p_mir.n0 two_stage_opamp_dummy_magic_21_0.V_p_mir.t3 16.0005
R5182 two_stage_opamp_dummy_magic_21_0.V_p_mir.n0 two_stage_opamp_dummy_magic_21_0.V_p_mir.t0 16.0005
R5183 two_stage_opamp_dummy_magic_21_0.V_p_mir.n1 two_stage_opamp_dummy_magic_21_0.V_p_mir.t1 9.6005
R5184 two_stage_opamp_dummy_magic_21_0.V_p_mir.t2 two_stage_opamp_dummy_magic_21_0.V_p_mir.n1 9.6005
R5185 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t8 525.38
R5186 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t5 525.38
R5187 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t2 483.608
R5188 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t3 360.43
R5189 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t7 291.209
R5190 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t4 281.168
R5191 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t9 281.168
R5192 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t6 281.168
R5193 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n0 244.214
R5194 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n4 202.44
R5195 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n5 202.159
R5196 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n2 165.972
R5197 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t1 117.754
R5198 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n6 117.254
R5199 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n1 79.2627
R5200 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n3 18.9067
R5201 VOUT-.n110 VOUT-.t10 113.16
R5202 VOUT-.n1 VOUT-.n0 34.9935
R5203 VOUT-.n5 VOUT-.n4 34.9935
R5204 VOUT-.n7 VOUT-.n6 34.9935
R5205 VOUT-.n11 VOUT-.n10 34.9935
R5206 VOUT-.n14 VOUT-.n13 34.9935
R5207 VOUT-.n18 VOUT-.n17 34.9935
R5208 VOUT-.n100 VOUT-.n20 20.4693
R5209 VOUT-.n100 VOUT-.n99 11.6871
R5210 VOUT- VOUT-.n100 9.8755
R5211 VOUT-.n103 VOUT-.n102 9.73997
R5212 VOUT-.n105 VOUT-.n104 9.73997
R5213 VOUT-.n108 VOUT-.n107 9.73997
R5214 VOUT-.n108 VOUT-.n106 7.14633
R5215 VOUT-.n106 VOUT-.n103 7.14633
R5216 VOUT-.n103 VOUT-.n101 7.14633
R5217 VOUT-.n0 VOUT-.t11 6.56717
R5218 VOUT-.n0 VOUT-.t0 6.56717
R5219 VOUT-.n4 VOUT-.t15 6.56717
R5220 VOUT-.n4 VOUT-.t3 6.56717
R5221 VOUT-.n6 VOUT-.t5 6.56717
R5222 VOUT-.n6 VOUT-.t18 6.56717
R5223 VOUT-.n10 VOUT-.t1 6.56717
R5224 VOUT-.n10 VOUT-.t17 6.56717
R5225 VOUT-.n13 VOUT-.t12 6.56717
R5226 VOUT-.n13 VOUT-.t2 6.56717
R5227 VOUT-.n17 VOUT-.t4 6.56717
R5228 VOUT-.n17 VOUT-.t16 6.56717
R5229 VOUT-.n18 VOUT-.n16 6.3755
R5230 VOUT-.n19 VOUT-.n18 6.3755
R5231 VOUT-.n8 VOUT-.n5 6.3755
R5232 VOUT-.n5 VOUT-.n3 6.3755
R5233 VOUT-.n105 VOUT-.n101 6.02133
R5234 VOUT-.n106 VOUT-.n105 6.02133
R5235 VOUT-.n109 VOUT-.n108 6.02133
R5236 VOUT-.n7 VOUT-.n3 5.813
R5237 VOUT-.n8 VOUT-.n7 5.813
R5238 VOUT-.n12 VOUT-.n11 5.813
R5239 VOUT-.n11 VOUT-.n9 5.813
R5240 VOUT-.n15 VOUT-.n14 5.813
R5241 VOUT-.n14 VOUT-.n2 5.813
R5242 VOUT-.n16 VOUT-.n1 5.813
R5243 VOUT-.n47 VOUT-.t108 4.8295
R5244 VOUT-.n56 VOUT-.t65 4.8295
R5245 VOUT-.n54 VOUT-.t118 4.8295
R5246 VOUT-.n52 VOUT-.t151 4.8295
R5247 VOUT-.n50 VOUT-.t44 4.8295
R5248 VOUT-.n49 VOUT-.t67 4.8295
R5249 VOUT-.n69 VOUT-.t27 4.8295
R5250 VOUT-.n70 VOUT-.t76 4.8295
R5251 VOUT-.n72 VOUT-.t62 4.8295
R5252 VOUT-.n73 VOUT-.t112 4.8295
R5253 VOUT-.n75 VOUT-.t114 4.8295
R5254 VOUT-.n76 VOUT-.t99 4.8295
R5255 VOUT-.n78 VOUT-.t74 4.8295
R5256 VOUT-.n79 VOUT-.t55 4.8295
R5257 VOUT-.n81 VOUT-.t109 4.8295
R5258 VOUT-.n82 VOUT-.t91 4.8295
R5259 VOUT-.n84 VOUT-.t68 4.8295
R5260 VOUT-.n85 VOUT-.t52 4.8295
R5261 VOUT-.n87 VOUT-.t29 4.8295
R5262 VOUT-.n88 VOUT-.t153 4.8295
R5263 VOUT-.n90 VOUT-.t63 4.8295
R5264 VOUT-.n91 VOUT-.t46 4.8295
R5265 VOUT-.n93 VOUT-.t22 4.8295
R5266 VOUT-.n94 VOUT-.t146 4.8295
R5267 VOUT-.n21 VOUT-.t117 4.8295
R5268 VOUT-.n23 VOUT-.t72 4.8295
R5269 VOUT-.n35 VOUT-.t37 4.8295
R5270 VOUT-.n36 VOUT-.t20 4.8295
R5271 VOUT-.n38 VOUT-.t79 4.8295
R5272 VOUT-.n39 VOUT-.t60 4.8295
R5273 VOUT-.n41 VOUT-.t121 4.8295
R5274 VOUT-.n42 VOUT-.t104 4.8295
R5275 VOUT-.n44 VOUT-.t84 4.8295
R5276 VOUT-.n45 VOUT-.t66 4.8295
R5277 VOUT-.n96 VOUT-.t123 4.8295
R5278 VOUT-.n58 VOUT-.t95 4.8154
R5279 VOUT-.n59 VOUT-.t70 4.8154
R5280 VOUT-.n60 VOUT-.t110 4.8154
R5281 VOUT-.n61 VOUT-.t145 4.8154
R5282 VOUT-.n58 VOUT-.t32 4.806
R5283 VOUT-.n59 VOUT-.t150 4.806
R5284 VOUT-.n60 VOUT-.t50 4.806
R5285 VOUT-.n61 VOUT-.t87 4.806
R5286 VOUT-.n62 VOUT-.t125 4.806
R5287 VOUT-.n63 VOUT-.t105 4.806
R5288 VOUT-.n64 VOUT-.t140 4.806
R5289 VOUT-.n65 VOUT-.t36 4.806
R5290 VOUT-.n66 VOUT-.t156 4.806
R5291 VOUT-.n67 VOUT-.t53 4.806
R5292 VOUT-.n24 VOUT-.t73 4.806
R5293 VOUT-.n25 VOUT-.t116 4.806
R5294 VOUT-.n26 VOUT-.t64 4.806
R5295 VOUT-.n27 VOUT-.t154 4.806
R5296 VOUT-.n28 VOUT-.t106 4.806
R5297 VOUT-.n29 VOUT-.t143 4.806
R5298 VOUT-.n30 VOUT-.t96 4.806
R5299 VOUT-.n31 VOUT-.t42 4.806
R5300 VOUT-.n32 VOUT-.t86 4.806
R5301 VOUT-.n33 VOUT-.t34 4.806
R5302 VOUT-.n47 VOUT-.t69 4.5005
R5303 VOUT-.n48 VOUT-.t90 4.5005
R5304 VOUT-.n56 VOUT-.t80 4.5005
R5305 VOUT-.n57 VOUT-.t43 4.5005
R5306 VOUT-.n54 VOUT-.t56 4.5005
R5307 VOUT-.n55 VOUT-.t21 4.5005
R5308 VOUT-.n52 VOUT-.t98 4.5005
R5309 VOUT-.n53 VOUT-.t59 4.5005
R5310 VOUT-.n50 VOUT-.t136 4.5005
R5311 VOUT-.n51 VOUT-.t101 4.5005
R5312 VOUT-.n49 VOUT-.t30 4.5005
R5313 VOUT-.n68 VOUT-.t51 4.5005
R5314 VOUT-.n67 VOUT-.t155 4.5005
R5315 VOUT-.n66 VOUT-.t119 4.5005
R5316 VOUT-.n65 VOUT-.t139 4.5005
R5317 VOUT-.n64 VOUT-.t102 4.5005
R5318 VOUT-.n63 VOUT-.t61 4.5005
R5319 VOUT-.n62 VOUT-.t85 4.5005
R5320 VOUT-.n61 VOUT-.t45 4.5005
R5321 VOUT-.n60 VOUT-.t147 4.5005
R5322 VOUT-.n59 VOUT-.t111 4.5005
R5323 VOUT-.n58 VOUT-.t134 4.5005
R5324 VOUT-.n69 VOUT-.t130 4.5005
R5325 VOUT-.n71 VOUT-.t152 4.5005
R5326 VOUT-.n70 VOUT-.t115 4.5005
R5327 VOUT-.n72 VOUT-.t23 4.5005
R5328 VOUT-.n74 VOUT-.t47 4.5005
R5329 VOUT-.n73 VOUT-.t148 4.5005
R5330 VOUT-.n75 VOUT-.t78 4.5005
R5331 VOUT-.n77 VOUT-.t26 4.5005
R5332 VOUT-.n76 VOUT-.t132 4.5005
R5333 VOUT-.n78 VOUT-.t39 4.5005
R5334 VOUT-.n80 VOUT-.t128 4.5005
R5335 VOUT-.n79 VOUT-.t92 4.5005
R5336 VOUT-.n81 VOUT-.t71 4.5005
R5337 VOUT-.n83 VOUT-.t19 4.5005
R5338 VOUT-.n82 VOUT-.t126 4.5005
R5339 VOUT-.n84 VOUT-.t33 4.5005
R5340 VOUT-.n86 VOUT-.t122 4.5005
R5341 VOUT-.n85 VOUT-.t88 4.5005
R5342 VOUT-.n87 VOUT-.t135 4.5005
R5343 VOUT-.n89 VOUT-.t82 4.5005
R5344 VOUT-.n88 VOUT-.t48 4.5005
R5345 VOUT-.n90 VOUT-.t28 4.5005
R5346 VOUT-.n92 VOUT-.t120 4.5005
R5347 VOUT-.n91 VOUT-.t81 4.5005
R5348 VOUT-.n93 VOUT-.t129 4.5005
R5349 VOUT-.n95 VOUT-.t77 4.5005
R5350 VOUT-.n94 VOUT-.t40 4.5005
R5351 VOUT-.n21 VOUT-.t25 4.5005
R5352 VOUT-.n22 VOUT-.t124 4.5005
R5353 VOUT-.n23 VOUT-.t38 4.5005
R5354 VOUT-.n34 VOUT-.t127 4.5005
R5355 VOUT-.n33 VOUT-.t94 4.5005
R5356 VOUT-.n32 VOUT-.t54 4.5005
R5357 VOUT-.n31 VOUT-.t144 4.5005
R5358 VOUT-.n30 VOUT-.t113 4.5005
R5359 VOUT-.n29 VOUT-.t75 4.5005
R5360 VOUT-.n28 VOUT-.t24 4.5005
R5361 VOUT-.n27 VOUT-.t131 4.5005
R5362 VOUT-.n26 VOUT-.t97 4.5005
R5363 VOUT-.n25 VOUT-.t58 4.5005
R5364 VOUT-.n24 VOUT-.t149 4.5005
R5365 VOUT-.n35 VOUT-.t142 4.5005
R5366 VOUT-.n37 VOUT-.t93 4.5005
R5367 VOUT-.n36 VOUT-.t57 4.5005
R5368 VOUT-.n38 VOUT-.t41 4.5005
R5369 VOUT-.n40 VOUT-.t133 4.5005
R5370 VOUT-.n39 VOUT-.t100 4.5005
R5371 VOUT-.n41 VOUT-.t83 4.5005
R5372 VOUT-.n43 VOUT-.t31 4.5005
R5373 VOUT-.n42 VOUT-.t137 4.5005
R5374 VOUT-.n44 VOUT-.t49 4.5005
R5375 VOUT-.n46 VOUT-.t138 4.5005
R5376 VOUT-.n45 VOUT-.t103 4.5005
R5377 VOUT-.n96 VOUT-.t89 4.5005
R5378 VOUT-.n97 VOUT-.t35 4.5005
R5379 VOUT-.n98 VOUT-.t141 4.5005
R5380 VOUT-.n99 VOUT-.t107 4.5005
R5381 VOUT-.n20 VOUT-.n19 4.5005
R5382 VOUT-.n102 VOUT-.t9 3.42907
R5383 VOUT-.n102 VOUT-.t13 3.42907
R5384 VOUT-.n104 VOUT-.t8 3.42907
R5385 VOUT-.n104 VOUT-.t7 3.42907
R5386 VOUT-.n107 VOUT-.t14 3.42907
R5387 VOUT-.n107 VOUT-.t6 3.42907
R5388 VOUT-.n110 VOUT-.n109 1.69693
R5389 VOUT- VOUT-.n110 1.53175
R5390 VOUT-.n20 VOUT-.n1 1.313
R5391 VOUT-.n109 VOUT-.n101 1.13443
R5392 VOUT-.n19 VOUT-.n2 0.563
R5393 VOUT-.n9 VOUT-.n2 0.563
R5394 VOUT-.n9 VOUT-.n8 0.563
R5395 VOUT-.n12 VOUT-.n3 0.563
R5396 VOUT-.n15 VOUT-.n12 0.563
R5397 VOUT-.n16 VOUT-.n15 0.563
R5398 VOUT-.n48 VOUT-.n47 0.3295
R5399 VOUT-.n57 VOUT-.n56 0.3295
R5400 VOUT-.n55 VOUT-.n54 0.3295
R5401 VOUT-.n53 VOUT-.n52 0.3295
R5402 VOUT-.n51 VOUT-.n50 0.3295
R5403 VOUT-.n68 VOUT-.n49 0.3295
R5404 VOUT-.n68 VOUT-.n67 0.3295
R5405 VOUT-.n67 VOUT-.n66 0.3295
R5406 VOUT-.n66 VOUT-.n65 0.3295
R5407 VOUT-.n65 VOUT-.n64 0.3295
R5408 VOUT-.n64 VOUT-.n63 0.3295
R5409 VOUT-.n63 VOUT-.n62 0.3295
R5410 VOUT-.n62 VOUT-.n61 0.3295
R5411 VOUT-.n61 VOUT-.n60 0.3295
R5412 VOUT-.n60 VOUT-.n59 0.3295
R5413 VOUT-.n59 VOUT-.n58 0.3295
R5414 VOUT-.n71 VOUT-.n69 0.3295
R5415 VOUT-.n71 VOUT-.n70 0.3295
R5416 VOUT-.n74 VOUT-.n72 0.3295
R5417 VOUT-.n74 VOUT-.n73 0.3295
R5418 VOUT-.n77 VOUT-.n75 0.3295
R5419 VOUT-.n77 VOUT-.n76 0.3295
R5420 VOUT-.n80 VOUT-.n78 0.3295
R5421 VOUT-.n80 VOUT-.n79 0.3295
R5422 VOUT-.n83 VOUT-.n81 0.3295
R5423 VOUT-.n83 VOUT-.n82 0.3295
R5424 VOUT-.n86 VOUT-.n84 0.3295
R5425 VOUT-.n86 VOUT-.n85 0.3295
R5426 VOUT-.n89 VOUT-.n87 0.3295
R5427 VOUT-.n89 VOUT-.n88 0.3295
R5428 VOUT-.n92 VOUT-.n90 0.3295
R5429 VOUT-.n92 VOUT-.n91 0.3295
R5430 VOUT-.n95 VOUT-.n93 0.3295
R5431 VOUT-.n95 VOUT-.n94 0.3295
R5432 VOUT-.n22 VOUT-.n21 0.3295
R5433 VOUT-.n34 VOUT-.n23 0.3295
R5434 VOUT-.n34 VOUT-.n33 0.3295
R5435 VOUT-.n33 VOUT-.n32 0.3295
R5436 VOUT-.n32 VOUT-.n31 0.3295
R5437 VOUT-.n31 VOUT-.n30 0.3295
R5438 VOUT-.n30 VOUT-.n29 0.3295
R5439 VOUT-.n29 VOUT-.n28 0.3295
R5440 VOUT-.n28 VOUT-.n27 0.3295
R5441 VOUT-.n27 VOUT-.n26 0.3295
R5442 VOUT-.n26 VOUT-.n25 0.3295
R5443 VOUT-.n25 VOUT-.n24 0.3295
R5444 VOUT-.n37 VOUT-.n35 0.3295
R5445 VOUT-.n37 VOUT-.n36 0.3295
R5446 VOUT-.n40 VOUT-.n38 0.3295
R5447 VOUT-.n40 VOUT-.n39 0.3295
R5448 VOUT-.n43 VOUT-.n41 0.3295
R5449 VOUT-.n43 VOUT-.n42 0.3295
R5450 VOUT-.n46 VOUT-.n44 0.3295
R5451 VOUT-.n46 VOUT-.n45 0.3295
R5452 VOUT-.n97 VOUT-.n96 0.3295
R5453 VOUT-.n98 VOUT-.n97 0.3295
R5454 VOUT-.n99 VOUT-.n98 0.3295
R5455 VOUT-.n62 VOUT-.n57 0.306
R5456 VOUT-.n63 VOUT-.n55 0.306
R5457 VOUT-.n64 VOUT-.n53 0.306
R5458 VOUT-.n65 VOUT-.n51 0.306
R5459 VOUT-.n68 VOUT-.n48 0.2825
R5460 VOUT-.n71 VOUT-.n68 0.2825
R5461 VOUT-.n74 VOUT-.n71 0.2825
R5462 VOUT-.n77 VOUT-.n74 0.2825
R5463 VOUT-.n80 VOUT-.n77 0.2825
R5464 VOUT-.n83 VOUT-.n80 0.2825
R5465 VOUT-.n86 VOUT-.n83 0.2825
R5466 VOUT-.n89 VOUT-.n86 0.2825
R5467 VOUT-.n92 VOUT-.n89 0.2825
R5468 VOUT-.n95 VOUT-.n92 0.2825
R5469 VOUT-.n34 VOUT-.n22 0.2825
R5470 VOUT-.n37 VOUT-.n34 0.2825
R5471 VOUT-.n40 VOUT-.n37 0.2825
R5472 VOUT-.n43 VOUT-.n40 0.2825
R5473 VOUT-.n46 VOUT-.n43 0.2825
R5474 VOUT-.n97 VOUT-.n46 0.2825
R5475 VOUT-.n97 VOUT-.n95 0.2825
R5476 two_stage_opamp_dummy_magic_21_0.VD2.n20 two_stage_opamp_dummy_magic_21_0.VD2.n19 49.3505
R5477 two_stage_opamp_dummy_magic_21_0.VD2.n23 two_stage_opamp_dummy_magic_21_0.VD2.n22 49.3505
R5478 two_stage_opamp_dummy_magic_21_0.VD2.n26 two_stage_opamp_dummy_magic_21_0.VD2.n25 49.3505
R5479 two_stage_opamp_dummy_magic_21_0.VD2.n0 two_stage_opamp_dummy_magic_21_0.VD2.n3 49.3505
R5480 two_stage_opamp_dummy_magic_21_0.VD2.n8 two_stage_opamp_dummy_magic_21_0.VD2.n7 49.3505
R5481 two_stage_opamp_dummy_magic_21_0.VD2.n10 two_stage_opamp_dummy_magic_21_0.VD2.n9 49.3505
R5482 two_stage_opamp_dummy_magic_21_0.VD2.n6 two_stage_opamp_dummy_magic_21_0.VD2.n5 49.3505
R5483 two_stage_opamp_dummy_magic_21_0.VD2.n15 two_stage_opamp_dummy_magic_21_0.VD2.n14 49.3505
R5484 two_stage_opamp_dummy_magic_21_0.VD2.n35 two_stage_opamp_dummy_magic_21_0.VD2.n34 49.3505
R5485 two_stage_opamp_dummy_magic_21_0.VD2.n31 two_stage_opamp_dummy_magic_21_0.VD2.n30 49.3505
R5486 two_stage_opamp_dummy_magic_21_0.VD2.n29 two_stage_opamp_dummy_magic_21_0.VD2.n28 49.3505
R5487 two_stage_opamp_dummy_magic_21_0.VD2.n19 two_stage_opamp_dummy_magic_21_0.VD2.t14 16.0005
R5488 two_stage_opamp_dummy_magic_21_0.VD2.n19 two_stage_opamp_dummy_magic_21_0.VD2.t13 16.0005
R5489 two_stage_opamp_dummy_magic_21_0.VD2.n22 two_stage_opamp_dummy_magic_21_0.VD2.t17 16.0005
R5490 two_stage_opamp_dummy_magic_21_0.VD2.n22 two_stage_opamp_dummy_magic_21_0.VD2.t1 16.0005
R5491 two_stage_opamp_dummy_magic_21_0.VD2.n25 two_stage_opamp_dummy_magic_21_0.VD2.t6 16.0005
R5492 two_stage_opamp_dummy_magic_21_0.VD2.n25 two_stage_opamp_dummy_magic_21_0.VD2.t0 16.0005
R5493 two_stage_opamp_dummy_magic_21_0.VD2.n3 two_stage_opamp_dummy_magic_21_0.VD2.t3 16.0005
R5494 two_stage_opamp_dummy_magic_21_0.VD2.n3 two_stage_opamp_dummy_magic_21_0.VD2.t9 16.0005
R5495 two_stage_opamp_dummy_magic_21_0.VD2.n7 two_stage_opamp_dummy_magic_21_0.VD2.t20 16.0005
R5496 two_stage_opamp_dummy_magic_21_0.VD2.n7 two_stage_opamp_dummy_magic_21_0.VD2.t7 16.0005
R5497 two_stage_opamp_dummy_magic_21_0.VD2.n9 two_stage_opamp_dummy_magic_21_0.VD2.t21 16.0005
R5498 two_stage_opamp_dummy_magic_21_0.VD2.n9 two_stage_opamp_dummy_magic_21_0.VD2.t19 16.0005
R5499 two_stage_opamp_dummy_magic_21_0.VD2.n5 two_stage_opamp_dummy_magic_21_0.VD2.t10 16.0005
R5500 two_stage_opamp_dummy_magic_21_0.VD2.n5 two_stage_opamp_dummy_magic_21_0.VD2.t4 16.0005
R5501 two_stage_opamp_dummy_magic_21_0.VD2.n14 two_stage_opamp_dummy_magic_21_0.VD2.t8 16.0005
R5502 two_stage_opamp_dummy_magic_21_0.VD2.n14 two_stage_opamp_dummy_magic_21_0.VD2.t11 16.0005
R5503 two_stage_opamp_dummy_magic_21_0.VD2.n34 two_stage_opamp_dummy_magic_21_0.VD2.t5 16.0005
R5504 two_stage_opamp_dummy_magic_21_0.VD2.n34 two_stage_opamp_dummy_magic_21_0.VD2.t2 16.0005
R5505 two_stage_opamp_dummy_magic_21_0.VD2.n30 two_stage_opamp_dummy_magic_21_0.VD2.t18 16.0005
R5506 two_stage_opamp_dummy_magic_21_0.VD2.n30 two_stage_opamp_dummy_magic_21_0.VD2.t12 16.0005
R5507 two_stage_opamp_dummy_magic_21_0.VD2.n28 two_stage_opamp_dummy_magic_21_0.VD2.t16 16.0005
R5508 two_stage_opamp_dummy_magic_21_0.VD2.n28 two_stage_opamp_dummy_magic_21_0.VD2.t15 16.0005
R5509 two_stage_opamp_dummy_magic_21_0.VD2.n29 two_stage_opamp_dummy_magic_21_0.VD2.n18 5.64633
R5510 two_stage_opamp_dummy_magic_21_0.VD2.n21 two_stage_opamp_dummy_magic_21_0.VD2.n20 5.64633
R5511 two_stage_opamp_dummy_magic_21_0.VD2.n13 two_stage_opamp_dummy_magic_21_0.VD2.n6 5.6255
R5512 two_stage_opamp_dummy_magic_21_0.VD2.n11 two_stage_opamp_dummy_magic_21_0.VD2.n8 5.6255
R5513 two_stage_opamp_dummy_magic_21_0.VD2.n16 two_stage_opamp_dummy_magic_21_0.VD2.n6 5.438
R5514 two_stage_opamp_dummy_magic_21_0.VD2.n8 two_stage_opamp_dummy_magic_21_0.VD2.n4 5.438
R5515 two_stage_opamp_dummy_magic_21_0.VD2.n24 two_stage_opamp_dummy_magic_21_0.VD2.n20 5.438
R5516 two_stage_opamp_dummy_magic_21_0.VD2.n32 two_stage_opamp_dummy_magic_21_0.VD2.n29 5.438
R5517 two_stage_opamp_dummy_magic_21_0.VD2.n23 two_stage_opamp_dummy_magic_21_0.VD2.n21 5.08383
R5518 two_stage_opamp_dummy_magic_21_0.VD2.n26 two_stage_opamp_dummy_magic_21_0.VD2.n2 5.08383
R5519 two_stage_opamp_dummy_magic_21_0.VD2.n1 two_stage_opamp_dummy_magic_21_0.VD2.n35 5.08383
R5520 two_stage_opamp_dummy_magic_21_0.VD2.n31 two_stage_opamp_dummy_magic_21_0.VD2.n18 5.08383
R5521 two_stage_opamp_dummy_magic_21_0.VD2.n11 two_stage_opamp_dummy_magic_21_0.VD2.n10 5.063
R5522 two_stage_opamp_dummy_magic_21_0.VD2.n15 two_stage_opamp_dummy_magic_21_0.VD2.n13 5.063
R5523 two_stage_opamp_dummy_magic_21_0.VD2.n12 two_stage_opamp_dummy_magic_21_0.VD2.n0 5.063
R5524 two_stage_opamp_dummy_magic_21_0.VD2 two_stage_opamp_dummy_magic_21_0.VD2.n2 5.02133
R5525 two_stage_opamp_dummy_magic_21_0.VD2.n24 two_stage_opamp_dummy_magic_21_0.VD2.n23 4.8755
R5526 two_stage_opamp_dummy_magic_21_0.VD2.n27 two_stage_opamp_dummy_magic_21_0.VD2.n26 4.8755
R5527 two_stage_opamp_dummy_magic_21_0.VD2.n10 two_stage_opamp_dummy_magic_21_0.VD2.n4 4.8755
R5528 two_stage_opamp_dummy_magic_21_0.VD2.n16 two_stage_opamp_dummy_magic_21_0.VD2.n15 4.8755
R5529 two_stage_opamp_dummy_magic_21_0.VD2.n35 two_stage_opamp_dummy_magic_21_0.VD2.n33 4.8755
R5530 two_stage_opamp_dummy_magic_21_0.VD2.n32 two_stage_opamp_dummy_magic_21_0.VD2.n31 4.8755
R5531 two_stage_opamp_dummy_magic_21_0.VD2.n0 two_stage_opamp_dummy_magic_21_0.VD2.n17 4.5005
R5532 two_stage_opamp_dummy_magic_21_0.VD2 two_stage_opamp_dummy_magic_21_0.VD2.n0 1.1255
R5533 two_stage_opamp_dummy_magic_21_0.VD2.n13 two_stage_opamp_dummy_magic_21_0.VD2.n12 0.563
R5534 two_stage_opamp_dummy_magic_21_0.VD2.n17 two_stage_opamp_dummy_magic_21_0.VD2.n16 0.563
R5535 two_stage_opamp_dummy_magic_21_0.VD2.n17 two_stage_opamp_dummy_magic_21_0.VD2.n4 0.563
R5536 two_stage_opamp_dummy_magic_21_0.VD2.n12 two_stage_opamp_dummy_magic_21_0.VD2.n11 0.563
R5537 two_stage_opamp_dummy_magic_21_0.VD2.n1 two_stage_opamp_dummy_magic_21_0.VD2.n18 0.563
R5538 two_stage_opamp_dummy_magic_21_0.VD2.n21 two_stage_opamp_dummy_magic_21_0.VD2.n2 0.563
R5539 two_stage_opamp_dummy_magic_21_0.VD2.n27 two_stage_opamp_dummy_magic_21_0.VD2.n24 0.563
R5540 two_stage_opamp_dummy_magic_21_0.VD2.n33 two_stage_opamp_dummy_magic_21_0.VD2.n27 0.563
R5541 two_stage_opamp_dummy_magic_21_0.VD2.n33 two_stage_opamp_dummy_magic_21_0.VD2.n32 0.563
R5542 two_stage_opamp_dummy_magic_21_0.VD2.n2 two_stage_opamp_dummy_magic_21_0.VD2.n1 0.46925
R5543 VOUT+.n9 VOUT+.t9 113.192
R5544 VOUT+.n11 VOUT+.n10 34.9935
R5545 VOUT+.n13 VOUT+.n12 34.9935
R5546 VOUT+.n17 VOUT+.n16 34.9935
R5547 VOUT+.n20 VOUT+.n19 34.9935
R5548 VOUT+.n23 VOUT+.n22 34.9935
R5549 VOUT+.n27 VOUT+.n26 34.9935
R5550 VOUT+.n110 VOUT+.n30 20.5005
R5551 VOUT+.n110 VOUT+.n109 11.6871
R5552 VOUT+.n2 VOUT+.n1 9.73997
R5553 VOUT+.n4 VOUT+.n3 9.73997
R5554 VOUT+.n7 VOUT+.n6 9.73997
R5555 VOUT+ VOUT+.n110 9.53033
R5556 VOUT+.n7 VOUT+.n5 7.14633
R5557 VOUT+.n5 VOUT+.n2 7.14633
R5558 VOUT+.n2 VOUT+.n0 7.14633
R5559 VOUT+.n10 VOUT+.t0 6.56717
R5560 VOUT+.n10 VOUT+.t5 6.56717
R5561 VOUT+.n12 VOUT+.t18 6.56717
R5562 VOUT+.n12 VOUT+.t4 6.56717
R5563 VOUT+.n16 VOUT+.t1 6.56717
R5564 VOUT+.n16 VOUT+.t17 6.56717
R5565 VOUT+.n19 VOUT+.t2 6.56717
R5566 VOUT+.n19 VOUT+.t3 6.56717
R5567 VOUT+.n22 VOUT+.t8 6.56717
R5568 VOUT+.n22 VOUT+.t6 6.56717
R5569 VOUT+.n26 VOUT+.t14 6.56717
R5570 VOUT+.n26 VOUT+.t7 6.56717
R5571 VOUT+.n21 VOUT+.n17 6.3755
R5572 VOUT+.n18 VOUT+.n17 6.3755
R5573 VOUT+.n29 VOUT+.n13 6.3755
R5574 VOUT+.n15 VOUT+.n13 6.3755
R5575 VOUT+.n4 VOUT+.n0 6.02133
R5576 VOUT+.n5 VOUT+.n4 6.02133
R5577 VOUT+.n8 VOUT+.n7 6.02133
R5578 VOUT+.n20 VOUT+.n18 5.813
R5579 VOUT+.n21 VOUT+.n20 5.813
R5580 VOUT+.n23 VOUT+.n14 5.813
R5581 VOUT+.n24 VOUT+.n23 5.813
R5582 VOUT+.n28 VOUT+.n27 5.813
R5583 VOUT+.n27 VOUT+.n25 5.813
R5584 VOUT+.n15 VOUT+.n11 5.813
R5585 VOUT+.n57 VOUT+.t85 4.8295
R5586 VOUT+.n59 VOUT+.t131 4.8295
R5587 VOUT+.n61 VOUT+.t31 4.8295
R5588 VOUT+.n63 VOUT+.t62 4.8295
R5589 VOUT+.n65 VOUT+.t114 4.8295
R5590 VOUT+.n77 VOUT+.t40 4.8295
R5591 VOUT+.n79 VOUT+.t34 4.8295
R5592 VOUT+.n80 VOUT+.t136 4.8295
R5593 VOUT+.n82 VOUT+.t70 4.8295
R5594 VOUT+.n83 VOUT+.t36 4.8295
R5595 VOUT+.n85 VOUT+.t95 4.8295
R5596 VOUT+.n86 VOUT+.t66 4.8295
R5597 VOUT+.n88 VOUT+.t55 4.8295
R5598 VOUT+.n89 VOUT+.t29 4.8295
R5599 VOUT+.n91 VOUT+.t91 4.8295
R5600 VOUT+.n92 VOUT+.t58 4.8295
R5601 VOUT+.n94 VOUT+.t49 4.8295
R5602 VOUT+.n95 VOUT+.t20 4.8295
R5603 VOUT+.n97 VOUT+.t148 4.8295
R5604 VOUT+.n98 VOUT+.t122 4.8295
R5605 VOUT+.n100 VOUT+.t44 4.8295
R5606 VOUT+.n101 VOUT+.t152 4.8295
R5607 VOUT+.n103 VOUT+.t142 4.8295
R5608 VOUT+.n104 VOUT+.t116 4.8295
R5609 VOUT+.n31 VOUT+.t108 4.8295
R5610 VOUT+.n43 VOUT+.t28 4.8295
R5611 VOUT+.n45 VOUT+.t24 4.8295
R5612 VOUT+.n46 VOUT+.t129 4.8295
R5613 VOUT+.n48 VOUT+.t61 4.8295
R5614 VOUT+.n49 VOUT+.t32 4.8295
R5615 VOUT+.n51 VOUT+.t100 4.8295
R5616 VOUT+.n52 VOUT+.t71 4.8295
R5617 VOUT+.n54 VOUT+.t69 4.8295
R5618 VOUT+.n55 VOUT+.t35 4.8295
R5619 VOUT+.n106 VOUT+.t77 4.8295
R5620 VOUT+.n70 VOUT+.t26 4.8154
R5621 VOUT+.n69 VOUT+.t59 4.8154
R5622 VOUT+.n68 VOUT+.t37 4.8154
R5623 VOUT+.n67 VOUT+.t81 4.8154
R5624 VOUT+.n76 VOUT+.t132 4.806
R5625 VOUT+.n75 VOUT+.t115 4.806
R5626 VOUT+.n74 VOUT+.t146 4.806
R5627 VOUT+.n73 VOUT+.t46 4.806
R5628 VOUT+.n72 VOUT+.t87 4.806
R5629 VOUT+.n71 VOUT+.t65 4.806
R5630 VOUT+.n70 VOUT+.t102 4.806
R5631 VOUT+.n69 VOUT+.t134 4.806
R5632 VOUT+.n68 VOUT+.t120 4.806
R5633 VOUT+.n67 VOUT+.t155 4.806
R5634 VOUT+.n42 VOUT+.t48 4.806
R5635 VOUT+.n41 VOUT+.t92 4.806
R5636 VOUT+.n40 VOUT+.t42 4.806
R5637 VOUT+.n39 VOUT+.t130 4.806
R5638 VOUT+.n38 VOUT+.t84 4.806
R5639 VOUT+.n37 VOUT+.t125 4.806
R5640 VOUT+.n36 VOUT+.t74 4.806
R5641 VOUT+.n35 VOUT+.t23 4.806
R5642 VOUT+.n34 VOUT+.t64 4.806
R5643 VOUT+.n33 VOUT+.t150 4.806
R5644 VOUT+.n58 VOUT+.t96 4.5005
R5645 VOUT+.n57 VOUT+.t57 4.5005
R5646 VOUT+.n59 VOUT+.t104 4.5005
R5647 VOUT+.n60 VOUT+.t73 4.5005
R5648 VOUT+.n61 VOUT+.t138 4.5005
R5649 VOUT+.n62 VOUT+.t107 4.5005
R5650 VOUT+.n63 VOUT+.t41 4.5005
R5651 VOUT+.n64 VOUT+.t143 4.5005
R5652 VOUT+.n65 VOUT+.t21 4.5005
R5653 VOUT+.n66 VOUT+.t126 4.5005
R5654 VOUT+.n67 VOUT+.t119 4.5005
R5655 VOUT+.n68 VOUT+.t82 4.5005
R5656 VOUT+.n69 VOUT+.t97 4.5005
R5657 VOUT+.n70 VOUT+.t63 4.5005
R5658 VOUT+.n71 VOUT+.t27 4.5005
R5659 VOUT+.n72 VOUT+.t45 4.5005
R5660 VOUT+.n73 VOUT+.t144 4.5005
R5661 VOUT+.n74 VOUT+.t112 4.5005
R5662 VOUT+.n75 VOUT+.t76 4.5005
R5663 VOUT+.n76 VOUT+.t93 4.5005
R5664 VOUT+.n78 VOUT+.t56 4.5005
R5665 VOUT+.n77 VOUT+.t19 4.5005
R5666 VOUT+.n79 VOUT+.t52 4.5005
R5667 VOUT+.n81 VOUT+.t156 4.5005
R5668 VOUT+.n80 VOUT+.t121 4.5005
R5669 VOUT+.n82 VOUT+.t89 4.5005
R5670 VOUT+.n84 VOUT+.t50 4.5005
R5671 VOUT+.n83 VOUT+.t151 4.5005
R5672 VOUT+.n85 VOUT+.t43 4.5005
R5673 VOUT+.n87 VOUT+.t145 4.5005
R5674 VOUT+.n86 VOUT+.t118 4.5005
R5675 VOUT+.n88 VOUT+.t141 4.5005
R5676 VOUT+.n90 VOUT+.t111 4.5005
R5677 VOUT+.n89 VOUT+.t80 4.5005
R5678 VOUT+.n91 VOUT+.t39 4.5005
R5679 VOUT+.n93 VOUT+.t139 4.5005
R5680 VOUT+.n92 VOUT+.t109 4.5005
R5681 VOUT+.n94 VOUT+.t135 4.5005
R5682 VOUT+.n96 VOUT+.t103 4.5005
R5683 VOUT+.n95 VOUT+.t72 4.5005
R5684 VOUT+.n97 VOUT+.t99 4.5005
R5685 VOUT+.n99 VOUT+.t68 4.5005
R5686 VOUT+.n98 VOUT+.t33 4.5005
R5687 VOUT+.n100 VOUT+.t133 4.5005
R5688 VOUT+.n102 VOUT+.t98 4.5005
R5689 VOUT+.n101 VOUT+.t67 4.5005
R5690 VOUT+.n103 VOUT+.t94 4.5005
R5691 VOUT+.n105 VOUT+.t60 4.5005
R5692 VOUT+.n104 VOUT+.t30 4.5005
R5693 VOUT+.n32 VOUT+.t101 4.5005
R5694 VOUT+.n31 VOUT+.t149 4.5005
R5695 VOUT+.n33 VOUT+.t88 4.5005
R5696 VOUT+.n34 VOUT+.t51 4.5005
R5697 VOUT+.n35 VOUT+.t137 4.5005
R5698 VOUT+.n36 VOUT+.t106 4.5005
R5699 VOUT+.n37 VOUT+.t75 4.5005
R5700 VOUT+.n38 VOUT+.t25 4.5005
R5701 VOUT+.n39 VOUT+.t128 4.5005
R5702 VOUT+.n40 VOUT+.t90 4.5005
R5703 VOUT+.n41 VOUT+.t54 4.5005
R5704 VOUT+.n42 VOUT+.t140 4.5005
R5705 VOUT+.n44 VOUT+.t110 4.5005
R5706 VOUT+.n43 VOUT+.t79 4.5005
R5707 VOUT+.n45 VOUT+.t113 4.5005
R5708 VOUT+.n47 VOUT+.t78 4.5005
R5709 VOUT+.n46 VOUT+.t38 4.5005
R5710 VOUT+.n48 VOUT+.t147 4.5005
R5711 VOUT+.n50 VOUT+.t117 4.5005
R5712 VOUT+.n49 VOUT+.t83 4.5005
R5713 VOUT+.n51 VOUT+.t47 4.5005
R5714 VOUT+.n53 VOUT+.t153 4.5005
R5715 VOUT+.n52 VOUT+.t123 4.5005
R5716 VOUT+.n54 VOUT+.t154 4.5005
R5717 VOUT+.n56 VOUT+.t124 4.5005
R5718 VOUT+.n55 VOUT+.t86 4.5005
R5719 VOUT+.n109 VOUT+.t105 4.5005
R5720 VOUT+.n108 VOUT+.t53 4.5005
R5721 VOUT+.n107 VOUT+.t22 4.5005
R5722 VOUT+.n106 VOUT+.t127 4.5005
R5723 VOUT+.n30 VOUT+.n29 4.5005
R5724 VOUT+.n1 VOUT+.t16 3.42907
R5725 VOUT+.n1 VOUT+.t13 3.42907
R5726 VOUT+.n3 VOUT+.t11 3.42907
R5727 VOUT+.n3 VOUT+.t10 3.42907
R5728 VOUT+.n6 VOUT+.t12 3.42907
R5729 VOUT+.n6 VOUT+.t15 3.42907
R5730 VOUT+.n9 VOUT+.n8 1.84425
R5731 VOUT+ VOUT+.n9 1.688
R5732 VOUT+.n30 VOUT+.n11 1.313
R5733 VOUT+.n8 VOUT+.n0 1.1255
R5734 VOUT+.n25 VOUT+.n15 0.563
R5735 VOUT+.n25 VOUT+.n24 0.563
R5736 VOUT+.n24 VOUT+.n21 0.563
R5737 VOUT+.n18 VOUT+.n14 0.563
R5738 VOUT+.n28 VOUT+.n14 0.563
R5739 VOUT+.n29 VOUT+.n28 0.563
R5740 VOUT+.n58 VOUT+.n57 0.3295
R5741 VOUT+.n60 VOUT+.n59 0.3295
R5742 VOUT+.n62 VOUT+.n61 0.3295
R5743 VOUT+.n64 VOUT+.n63 0.3295
R5744 VOUT+.n66 VOUT+.n65 0.3295
R5745 VOUT+.n68 VOUT+.n67 0.3295
R5746 VOUT+.n69 VOUT+.n68 0.3295
R5747 VOUT+.n70 VOUT+.n69 0.3295
R5748 VOUT+.n71 VOUT+.n70 0.3295
R5749 VOUT+.n72 VOUT+.n71 0.3295
R5750 VOUT+.n73 VOUT+.n72 0.3295
R5751 VOUT+.n74 VOUT+.n73 0.3295
R5752 VOUT+.n75 VOUT+.n74 0.3295
R5753 VOUT+.n76 VOUT+.n75 0.3295
R5754 VOUT+.n78 VOUT+.n76 0.3295
R5755 VOUT+.n78 VOUT+.n77 0.3295
R5756 VOUT+.n81 VOUT+.n79 0.3295
R5757 VOUT+.n81 VOUT+.n80 0.3295
R5758 VOUT+.n84 VOUT+.n82 0.3295
R5759 VOUT+.n84 VOUT+.n83 0.3295
R5760 VOUT+.n87 VOUT+.n85 0.3295
R5761 VOUT+.n87 VOUT+.n86 0.3295
R5762 VOUT+.n90 VOUT+.n88 0.3295
R5763 VOUT+.n90 VOUT+.n89 0.3295
R5764 VOUT+.n93 VOUT+.n91 0.3295
R5765 VOUT+.n93 VOUT+.n92 0.3295
R5766 VOUT+.n96 VOUT+.n94 0.3295
R5767 VOUT+.n96 VOUT+.n95 0.3295
R5768 VOUT+.n99 VOUT+.n97 0.3295
R5769 VOUT+.n99 VOUT+.n98 0.3295
R5770 VOUT+.n102 VOUT+.n100 0.3295
R5771 VOUT+.n102 VOUT+.n101 0.3295
R5772 VOUT+.n105 VOUT+.n103 0.3295
R5773 VOUT+.n105 VOUT+.n104 0.3295
R5774 VOUT+.n32 VOUT+.n31 0.3295
R5775 VOUT+.n34 VOUT+.n33 0.3295
R5776 VOUT+.n35 VOUT+.n34 0.3295
R5777 VOUT+.n36 VOUT+.n35 0.3295
R5778 VOUT+.n37 VOUT+.n36 0.3295
R5779 VOUT+.n38 VOUT+.n37 0.3295
R5780 VOUT+.n39 VOUT+.n38 0.3295
R5781 VOUT+.n40 VOUT+.n39 0.3295
R5782 VOUT+.n41 VOUT+.n40 0.3295
R5783 VOUT+.n42 VOUT+.n41 0.3295
R5784 VOUT+.n44 VOUT+.n42 0.3295
R5785 VOUT+.n44 VOUT+.n43 0.3295
R5786 VOUT+.n47 VOUT+.n45 0.3295
R5787 VOUT+.n47 VOUT+.n46 0.3295
R5788 VOUT+.n50 VOUT+.n48 0.3295
R5789 VOUT+.n50 VOUT+.n49 0.3295
R5790 VOUT+.n53 VOUT+.n51 0.3295
R5791 VOUT+.n53 VOUT+.n52 0.3295
R5792 VOUT+.n56 VOUT+.n54 0.3295
R5793 VOUT+.n56 VOUT+.n55 0.3295
R5794 VOUT+.n109 VOUT+.n108 0.3295
R5795 VOUT+.n108 VOUT+.n107 0.3295
R5796 VOUT+.n107 VOUT+.n106 0.3295
R5797 VOUT+.n74 VOUT+.n60 0.306
R5798 VOUT+.n73 VOUT+.n62 0.306
R5799 VOUT+.n72 VOUT+.n64 0.306
R5800 VOUT+.n71 VOUT+.n66 0.306
R5801 VOUT+.n78 VOUT+.n58 0.2825
R5802 VOUT+.n81 VOUT+.n78 0.2825
R5803 VOUT+.n84 VOUT+.n81 0.2825
R5804 VOUT+.n87 VOUT+.n84 0.2825
R5805 VOUT+.n90 VOUT+.n87 0.2825
R5806 VOUT+.n93 VOUT+.n90 0.2825
R5807 VOUT+.n96 VOUT+.n93 0.2825
R5808 VOUT+.n99 VOUT+.n96 0.2825
R5809 VOUT+.n102 VOUT+.n99 0.2825
R5810 VOUT+.n105 VOUT+.n102 0.2825
R5811 VOUT+.n44 VOUT+.n32 0.2825
R5812 VOUT+.n47 VOUT+.n44 0.2825
R5813 VOUT+.n50 VOUT+.n47 0.2825
R5814 VOUT+.n53 VOUT+.n50 0.2825
R5815 VOUT+.n56 VOUT+.n53 0.2825
R5816 VOUT+.n107 VOUT+.n56 0.2825
R5817 VOUT+.n107 VOUT+.n105 0.2825
R5818 two_stage_opamp_dummy_magic_21_0.cap_res_Y two_stage_opamp_dummy_magic_21_0.cap_res_Y.t138 49.2388
R5819 two_stage_opamp_dummy_magic_21_0.cap_res_Y two_stage_opamp_dummy_magic_21_0.cap_res_Y.t125 0.922875
R5820 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t116 0.1603
R5821 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t71 0.1603
R5822 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t20 0.1603
R5823 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t122 0.1603
R5824 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t120 0.1603
R5825 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t86 0.1603
R5826 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t90 0.1603
R5827 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t61 0.1603
R5828 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t127 0.1603
R5829 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t101 0.1603
R5830 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t98 0.1603
R5831 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t65 0.1603
R5832 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t136 0.1603
R5833 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t107 0.1603
R5834 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t34 0.1603
R5835 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t8 0.1603
R5836 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t4 0.1603
R5837 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t112 0.1603
R5838 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t40 0.1603
R5839 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t14 0.1603
R5840 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t79 0.1603
R5841 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t51 0.1603
R5842 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t121 0.1603
R5843 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t87 0.1603
R5844 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t85 0.1603
R5845 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t56 0.1603
R5846 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t124 0.1603
R5847 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t95 0.1603
R5848 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t27 0.1603
R5849 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t132 0.1603
R5850 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t128 0.1603
R5851 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t6 0.1603
R5852 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t92 0.1603
R5853 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t133 0.1603
R5854 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t82 0.1603
R5855 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t31 0.1603
R5856 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t72 0.1603
R5857 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t26 0.1603
R5858 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t114 0.1603
R5859 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t64 0.1603
R5860 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t108 0.1603
R5861 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t48 0.1603
R5862 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t25 0.1603
R5863 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t52 0.1603
R5864 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t83 0.1603
R5865 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t75 0.1603
R5866 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t119 0.1603
R5867 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t97 0.1603
R5868 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t130 0.1603
R5869 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t42 0.1603
R5870 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t135 0.1603
R5871 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t30 0.1603
R5872 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t94 0.1603
R5873 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t115 0.1603
R5874 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t13 0.1603
R5875 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t12 0.1603
R5876 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t49 0.1603
R5877 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t18 0.1603
R5878 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t60 0.159278
R5879 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n15 0.159278
R5880 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n16 0.159278
R5881 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n17 0.159278
R5882 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n18 0.159278
R5883 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n19 0.159278
R5884 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n20 0.159278
R5885 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n21 0.159278
R5886 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n22 0.159278
R5887 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n23 0.159278
R5888 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n24 0.159278
R5889 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n25 0.159278
R5890 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n26 0.159278
R5891 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n27 0.159278
R5892 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n28 0.159278
R5893 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n29 0.159278
R5894 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n30 0.159278
R5895 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t24 0.159278
R5896 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t41 0.159278
R5897 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t10 0.159278
R5898 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t1 0.159278
R5899 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t36 0.159278
R5900 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t22 0.159278
R5901 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t54 0.159278
R5902 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t91 0.159278
R5903 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t69 0.159278
R5904 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t110 0.159278
R5905 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t99 0.137822
R5906 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t137 0.1368
R5907 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t35 0.1368
R5908 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t104 0.1368
R5909 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t5 0.1368
R5910 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t67 0.1368
R5911 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t38 0.1368
R5912 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t113 0.1368
R5913 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t76 0.1368
R5914 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t15 0.1368
R5915 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t47 0.1368
R5916 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t117 0.1368
R5917 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t84 0.1368
R5918 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t21 0.1368
R5919 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t123 0.1368
R5920 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t57 0.1368
R5921 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t89 0.1368
R5922 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t23 0.1368
R5923 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t126 0.1368
R5924 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t62 0.1368
R5925 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t29 0.1368
R5926 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t103 0.1368
R5927 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t70 0.1368
R5928 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t2 0.1368
R5929 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t33 0.1368
R5930 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t109 0.1368
R5931 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t73 0.1368
R5932 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t9 0.1368
R5933 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t118 0.1368
R5934 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t43 0.1368
R5935 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t77 0.1368
R5936 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t7 0.1368
R5937 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t68 0.114322
R5938 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n6 0.1133
R5939 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n7 0.1133
R5940 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n8 0.1133
R5941 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n9 0.1133
R5942 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n10 0.1133
R5943 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n11 0.1133
R5944 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n12 0.1133
R5945 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n13 0.1133
R5946 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n14 0.1133
R5947 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n31 0.1133
R5948 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n32 0.1133
R5949 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n33 0.1133
R5950 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n0 0.1133
R5951 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n1 0.1133
R5952 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n2 0.1133
R5953 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n3 0.1133
R5954 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n4 0.1133
R5955 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n5 0.1133
R5956 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n34 0.1133
R5957 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t105 0.00152174
R5958 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t19 0.00152174
R5959 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t50 0.00152174
R5960 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t81 0.00152174
R5961 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t131 0.00152174
R5962 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t28 0.00152174
R5963 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t66 0.00152174
R5964 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t102 0.00152174
R5965 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t16 0.00152174
R5966 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t55 0.00152174
R5967 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t46 0.00152174
R5968 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t78 0.00152174
R5969 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t39 0.00152174
R5970 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t3 0.00152174
R5971 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t32 0.00152174
R5972 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t134 0.00152174
R5973 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t96 0.00152174
R5974 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t58 0.00152174
R5975 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t88 0.00152174
R5976 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t53 0.00152174
R5977 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t17 0.00152174
R5978 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t45 0.00152174
R5979 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t11 0.00152174
R5980 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t106 0.00152174
R5981 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t0 0.00152174
R5982 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t100 0.00152174
R5983 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t63 0.00152174
R5984 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t80 0.00152174
R5985 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t44 0.00152174
R5986 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t37 0.00152174
R5987 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t74 0.00152174
R5988 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t59 0.00152174
R5989 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t93 0.00152174
R5990 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t129 0.00152174
R5991 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t111 0.00152174
R5992 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n35 0.00152174
R5993 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t8 739.067
R5994 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n3 724.936
R5995 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t18 688.859
R5996 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n1 530.201
R5997 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n5 530.201
R5998 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n7 530.201
R5999 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n10 514.134
R6000 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n8 361.5
R6001 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n12 214.056
R6002 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t21 208.868
R6003 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t12 208.868
R6004 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t7 208.868
R6005 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t13 208.868
R6006 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t17 208.868
R6007 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t15 208.868
R6008 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t9 208.868
R6009 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t16 208.868
R6010 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t10 208.868
R6011 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n0 176.733
R6012 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n2 176.733
R6013 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n4 176.733
R6014 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n6 176.733
R6015 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t11 174.726
R6016 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t20 174.726
R6017 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t14 174.726
R6018 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t19 174.726
R6019 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n14 173.591
R6020 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n17 169.216
R6021 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n15 169.216
R6022 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n9 128.534
R6023 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n11 128.534
R6024 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t6 125.736
R6025 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n19 46.2505
R6026 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t0 13.1338
R6027 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t4 13.1338
R6028 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t3 13.1338
R6029 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t1 13.1338
R6030 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t5 13.1338
R6031 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t2 13.1338
R6032 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n18 10.0317
R6033 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n16 4.3755
R6034 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n13 3.03175
R6035 two_stage_opamp_dummy_magic_21_0.Y.n65 two_stage_opamp_dummy_magic_21_0.Y.t48 1172.87
R6036 two_stage_opamp_dummy_magic_21_0.Y.n63 two_stage_opamp_dummy_magic_21_0.Y.t39 1172.87
R6037 two_stage_opamp_dummy_magic_21_0.Y.n65 two_stage_opamp_dummy_magic_21_0.Y.t31 996.134
R6038 two_stage_opamp_dummy_magic_21_0.Y.n66 two_stage_opamp_dummy_magic_21_0.Y.t49 996.134
R6039 two_stage_opamp_dummy_magic_21_0.Y.n67 two_stage_opamp_dummy_magic_21_0.Y.t33 996.134
R6040 two_stage_opamp_dummy_magic_21_0.Y.n68 two_stage_opamp_dummy_magic_21_0.Y.t42 996.134
R6041 two_stage_opamp_dummy_magic_21_0.Y.n69 two_stage_opamp_dummy_magic_21_0.Y.t26 996.134
R6042 two_stage_opamp_dummy_magic_21_0.Y.n70 two_stage_opamp_dummy_magic_21_0.Y.t45 996.134
R6043 two_stage_opamp_dummy_magic_21_0.Y.n64 two_stage_opamp_dummy_magic_21_0.Y.t28 996.134
R6044 two_stage_opamp_dummy_magic_21_0.Y.n63 two_stage_opamp_dummy_magic_21_0.Y.t47 996.134
R6045 two_stage_opamp_dummy_magic_21_0.Y.n58 two_stage_opamp_dummy_magic_21_0.Y.t44 690.867
R6046 two_stage_opamp_dummy_magic_21_0.Y.n51 two_stage_opamp_dummy_magic_21_0.Y.t35 690.867
R6047 two_stage_opamp_dummy_magic_21_0.Y.n49 two_stage_opamp_dummy_magic_21_0.Y.t38 530.201
R6048 two_stage_opamp_dummy_magic_21_0.Y.n42 two_stage_opamp_dummy_magic_21_0.Y.t30 530.201
R6049 two_stage_opamp_dummy_magic_21_0.Y.n58 two_stage_opamp_dummy_magic_21_0.Y.t27 514.134
R6050 two_stage_opamp_dummy_magic_21_0.Y.n51 two_stage_opamp_dummy_magic_21_0.Y.t43 514.134
R6051 two_stage_opamp_dummy_magic_21_0.Y.n52 two_stage_opamp_dummy_magic_21_0.Y.t54 514.134
R6052 two_stage_opamp_dummy_magic_21_0.Y.n53 two_stage_opamp_dummy_magic_21_0.Y.t40 514.134
R6053 two_stage_opamp_dummy_magic_21_0.Y.n54 two_stage_opamp_dummy_magic_21_0.Y.t52 514.134
R6054 two_stage_opamp_dummy_magic_21_0.Y.n55 two_stage_opamp_dummy_magic_21_0.Y.t36 514.134
R6055 two_stage_opamp_dummy_magic_21_0.Y.n56 two_stage_opamp_dummy_magic_21_0.Y.t29 514.134
R6056 two_stage_opamp_dummy_magic_21_0.Y.n57 two_stage_opamp_dummy_magic_21_0.Y.t46 514.134
R6057 two_stage_opamp_dummy_magic_21_0.Y.n49 two_stage_opamp_dummy_magic_21_0.Y.t53 353.467
R6058 two_stage_opamp_dummy_magic_21_0.Y.n48 two_stage_opamp_dummy_magic_21_0.Y.t41 353.467
R6059 two_stage_opamp_dummy_magic_21_0.Y.n47 two_stage_opamp_dummy_magic_21_0.Y.t25 353.467
R6060 two_stage_opamp_dummy_magic_21_0.Y.n46 two_stage_opamp_dummy_magic_21_0.Y.t32 353.467
R6061 two_stage_opamp_dummy_magic_21_0.Y.n45 two_stage_opamp_dummy_magic_21_0.Y.t50 353.467
R6062 two_stage_opamp_dummy_magic_21_0.Y.n44 two_stage_opamp_dummy_magic_21_0.Y.t34 353.467
R6063 two_stage_opamp_dummy_magic_21_0.Y.n43 two_stage_opamp_dummy_magic_21_0.Y.t51 353.467
R6064 two_stage_opamp_dummy_magic_21_0.Y.n42 two_stage_opamp_dummy_magic_21_0.Y.t37 353.467
R6065 two_stage_opamp_dummy_magic_21_0.Y.n72 two_stage_opamp_dummy_magic_21_0.Y.n71 304.375
R6066 two_stage_opamp_dummy_magic_21_0.Y.n60 two_stage_opamp_dummy_magic_21_0.Y.n50 216.9
R6067 two_stage_opamp_dummy_magic_21_0.Y.n60 two_stage_opamp_dummy_magic_21_0.Y.n59 216.9
R6068 two_stage_opamp_dummy_magic_21_0.Y.n64 two_stage_opamp_dummy_magic_21_0.Y.n63 176.733
R6069 two_stage_opamp_dummy_magic_21_0.Y.n66 two_stage_opamp_dummy_magic_21_0.Y.n65 176.733
R6070 two_stage_opamp_dummy_magic_21_0.Y.n67 two_stage_opamp_dummy_magic_21_0.Y.n66 176.733
R6071 two_stage_opamp_dummy_magic_21_0.Y.n68 two_stage_opamp_dummy_magic_21_0.Y.n67 176.733
R6072 two_stage_opamp_dummy_magic_21_0.Y.n69 two_stage_opamp_dummy_magic_21_0.Y.n68 176.733
R6073 two_stage_opamp_dummy_magic_21_0.Y.n70 two_stage_opamp_dummy_magic_21_0.Y.n69 176.733
R6074 two_stage_opamp_dummy_magic_21_0.Y.n48 two_stage_opamp_dummy_magic_21_0.Y.n47 176.733
R6075 two_stage_opamp_dummy_magic_21_0.Y.n47 two_stage_opamp_dummy_magic_21_0.Y.n46 176.733
R6076 two_stage_opamp_dummy_magic_21_0.Y.n46 two_stage_opamp_dummy_magic_21_0.Y.n45 176.733
R6077 two_stage_opamp_dummy_magic_21_0.Y.n45 two_stage_opamp_dummy_magic_21_0.Y.n44 176.733
R6078 two_stage_opamp_dummy_magic_21_0.Y.n44 two_stage_opamp_dummy_magic_21_0.Y.n43 176.733
R6079 two_stage_opamp_dummy_magic_21_0.Y.n43 two_stage_opamp_dummy_magic_21_0.Y.n42 176.733
R6080 two_stage_opamp_dummy_magic_21_0.Y.n57 two_stage_opamp_dummy_magic_21_0.Y.n56 176.733
R6081 two_stage_opamp_dummy_magic_21_0.Y.n56 two_stage_opamp_dummy_magic_21_0.Y.n55 176.733
R6082 two_stage_opamp_dummy_magic_21_0.Y.n55 two_stage_opamp_dummy_magic_21_0.Y.n54 176.733
R6083 two_stage_opamp_dummy_magic_21_0.Y.n54 two_stage_opamp_dummy_magic_21_0.Y.n53 176.733
R6084 two_stage_opamp_dummy_magic_21_0.Y.n53 two_stage_opamp_dummy_magic_21_0.Y.n52 176.733
R6085 two_stage_opamp_dummy_magic_21_0.Y.n52 two_stage_opamp_dummy_magic_21_0.Y.n51 176.733
R6086 two_stage_opamp_dummy_magic_21_0.Y.n61 two_stage_opamp_dummy_magic_21_0.Y.n60 175.05
R6087 two_stage_opamp_dummy_magic_21_0.Y.n22 two_stage_opamp_dummy_magic_21_0.Y.n21 66.0338
R6088 two_stage_opamp_dummy_magic_21_0.Y.n26 two_stage_opamp_dummy_magic_21_0.Y.n25 66.0338
R6089 two_stage_opamp_dummy_magic_21_0.Y.n28 two_stage_opamp_dummy_magic_21_0.Y.n27 66.0338
R6090 two_stage_opamp_dummy_magic_21_0.Y.n32 two_stage_opamp_dummy_magic_21_0.Y.n31 66.0338
R6091 two_stage_opamp_dummy_magic_21_0.Y.n35 two_stage_opamp_dummy_magic_21_0.Y.n34 66.0338
R6092 two_stage_opamp_dummy_magic_21_0.Y.n39 two_stage_opamp_dummy_magic_21_0.Y.n38 66.0338
R6093 two_stage_opamp_dummy_magic_21_0.Y.t21 two_stage_opamp_dummy_magic_21_0.Y.n72 49.4802
R6094 two_stage_opamp_dummy_magic_21_0.Y.n1 two_stage_opamp_dummy_magic_21_0.Y.n0 49.3505
R6095 two_stage_opamp_dummy_magic_21_0.Y.n6 two_stage_opamp_dummy_magic_21_0.Y.n5 49.3505
R6096 two_stage_opamp_dummy_magic_21_0.Y.n9 two_stage_opamp_dummy_magic_21_0.Y.n8 49.3505
R6097 two_stage_opamp_dummy_magic_21_0.Y.n12 two_stage_opamp_dummy_magic_21_0.Y.n11 49.3505
R6098 two_stage_opamp_dummy_magic_21_0.Y.n4 two_stage_opamp_dummy_magic_21_0.Y.n3 49.3505
R6099 two_stage_opamp_dummy_magic_21_0.Y.n17 two_stage_opamp_dummy_magic_21_0.Y.n16 49.3505
R6100 two_stage_opamp_dummy_magic_21_0.Y.n71 two_stage_opamp_dummy_magic_21_0.Y.n64 40.1672
R6101 two_stage_opamp_dummy_magic_21_0.Y.n71 two_stage_opamp_dummy_magic_21_0.Y.n70 40.1672
R6102 two_stage_opamp_dummy_magic_21_0.Y.n50 two_stage_opamp_dummy_magic_21_0.Y.n48 40.1672
R6103 two_stage_opamp_dummy_magic_21_0.Y.n50 two_stage_opamp_dummy_magic_21_0.Y.n49 40.1672
R6104 two_stage_opamp_dummy_magic_21_0.Y.n59 two_stage_opamp_dummy_magic_21_0.Y.n57 40.1672
R6105 two_stage_opamp_dummy_magic_21_0.Y.n59 two_stage_opamp_dummy_magic_21_0.Y.n58 40.1672
R6106 two_stage_opamp_dummy_magic_21_0.Y.n61 two_stage_opamp_dummy_magic_21_0.Y.n41 17.6567
R6107 two_stage_opamp_dummy_magic_21_0.Y.n0 two_stage_opamp_dummy_magic_21_0.Y.t6 16.0005
R6108 two_stage_opamp_dummy_magic_21_0.Y.n0 two_stage_opamp_dummy_magic_21_0.Y.t5 16.0005
R6109 two_stage_opamp_dummy_magic_21_0.Y.n5 two_stage_opamp_dummy_magic_21_0.Y.t18 16.0005
R6110 two_stage_opamp_dummy_magic_21_0.Y.n5 two_stage_opamp_dummy_magic_21_0.Y.t22 16.0005
R6111 two_stage_opamp_dummy_magic_21_0.Y.n8 two_stage_opamp_dummy_magic_21_0.Y.t4 16.0005
R6112 two_stage_opamp_dummy_magic_21_0.Y.n8 two_stage_opamp_dummy_magic_21_0.Y.t23 16.0005
R6113 two_stage_opamp_dummy_magic_21_0.Y.n11 two_stage_opamp_dummy_magic_21_0.Y.t20 16.0005
R6114 two_stage_opamp_dummy_magic_21_0.Y.n11 two_stage_opamp_dummy_magic_21_0.Y.t0 16.0005
R6115 two_stage_opamp_dummy_magic_21_0.Y.n3 two_stage_opamp_dummy_magic_21_0.Y.t1 16.0005
R6116 two_stage_opamp_dummy_magic_21_0.Y.n3 two_stage_opamp_dummy_magic_21_0.Y.t19 16.0005
R6117 two_stage_opamp_dummy_magic_21_0.Y.n16 two_stage_opamp_dummy_magic_21_0.Y.t12 16.0005
R6118 two_stage_opamp_dummy_magic_21_0.Y.n16 two_stage_opamp_dummy_magic_21_0.Y.t10 16.0005
R6119 two_stage_opamp_dummy_magic_21_0.Y.n21 two_stage_opamp_dummy_magic_21_0.Y.t8 11.2576
R6120 two_stage_opamp_dummy_magic_21_0.Y.n21 two_stage_opamp_dummy_magic_21_0.Y.t13 11.2576
R6121 two_stage_opamp_dummy_magic_21_0.Y.n25 two_stage_opamp_dummy_magic_21_0.Y.t11 11.2576
R6122 two_stage_opamp_dummy_magic_21_0.Y.n25 two_stage_opamp_dummy_magic_21_0.Y.t2 11.2576
R6123 two_stage_opamp_dummy_magic_21_0.Y.n27 two_stage_opamp_dummy_magic_21_0.Y.t16 11.2576
R6124 two_stage_opamp_dummy_magic_21_0.Y.n27 two_stage_opamp_dummy_magic_21_0.Y.t7 11.2576
R6125 two_stage_opamp_dummy_magic_21_0.Y.n31 two_stage_opamp_dummy_magic_21_0.Y.t9 11.2576
R6126 two_stage_opamp_dummy_magic_21_0.Y.n31 two_stage_opamp_dummy_magic_21_0.Y.t14 11.2576
R6127 two_stage_opamp_dummy_magic_21_0.Y.n34 two_stage_opamp_dummy_magic_21_0.Y.t15 11.2576
R6128 two_stage_opamp_dummy_magic_21_0.Y.n34 two_stage_opamp_dummy_magic_21_0.Y.t17 11.2576
R6129 two_stage_opamp_dummy_magic_21_0.Y.n38 two_stage_opamp_dummy_magic_21_0.Y.t24 11.2576
R6130 two_stage_opamp_dummy_magic_21_0.Y.n38 two_stage_opamp_dummy_magic_21_0.Y.t3 11.2576
R6131 two_stage_opamp_dummy_magic_21_0.Y.n62 two_stage_opamp_dummy_magic_21_0.Y.n20 10.2817
R6132 two_stage_opamp_dummy_magic_21_0.Y.n29 two_stage_opamp_dummy_magic_21_0.Y.n26 5.91717
R6133 two_stage_opamp_dummy_magic_21_0.Y.n26 two_stage_opamp_dummy_magic_21_0.Y.n24 5.91717
R6134 two_stage_opamp_dummy_magic_21_0.Y.n37 two_stage_opamp_dummy_magic_21_0.Y.n22 5.91717
R6135 two_stage_opamp_dummy_magic_21_0.Y.n15 two_stage_opamp_dummy_magic_21_0.Y.n4 5.6255
R6136 two_stage_opamp_dummy_magic_21_0.Y.n10 two_stage_opamp_dummy_magic_21_0.Y.n6 5.6255
R6137 two_stage_opamp_dummy_magic_21_0.Y.n18 two_stage_opamp_dummy_magic_21_0.Y.n4 5.438
R6138 two_stage_opamp_dummy_magic_21_0.Y.n7 two_stage_opamp_dummy_magic_21_0.Y.n6 5.438
R6139 two_stage_opamp_dummy_magic_21_0.Y.n28 two_stage_opamp_dummy_magic_21_0.Y.n24 5.29217
R6140 two_stage_opamp_dummy_magic_21_0.Y.n29 two_stage_opamp_dummy_magic_21_0.Y.n28 5.29217
R6141 two_stage_opamp_dummy_magic_21_0.Y.n33 two_stage_opamp_dummy_magic_21_0.Y.n32 5.29217
R6142 two_stage_opamp_dummy_magic_21_0.Y.n32 two_stage_opamp_dummy_magic_21_0.Y.n30 5.29217
R6143 two_stage_opamp_dummy_magic_21_0.Y.n36 two_stage_opamp_dummy_magic_21_0.Y.n35 5.29217
R6144 two_stage_opamp_dummy_magic_21_0.Y.n35 two_stage_opamp_dummy_magic_21_0.Y.n23 5.29217
R6145 two_stage_opamp_dummy_magic_21_0.Y.n39 two_stage_opamp_dummy_magic_21_0.Y.n37 5.29217
R6146 two_stage_opamp_dummy_magic_21_0.Y.n40 two_stage_opamp_dummy_magic_21_0.Y.n39 5.29217
R6147 two_stage_opamp_dummy_magic_21_0.Y.n41 two_stage_opamp_dummy_magic_21_0.Y.n40 5.1255
R6148 two_stage_opamp_dummy_magic_21_0.Y.n10 two_stage_opamp_dummy_magic_21_0.Y.n9 5.063
R6149 two_stage_opamp_dummy_magic_21_0.Y.n13 two_stage_opamp_dummy_magic_21_0.Y.n12 5.063
R6150 two_stage_opamp_dummy_magic_21_0.Y.n17 two_stage_opamp_dummy_magic_21_0.Y.n15 5.063
R6151 two_stage_opamp_dummy_magic_21_0.Y.n14 two_stage_opamp_dummy_magic_21_0.Y.n1 5.063
R6152 two_stage_opamp_dummy_magic_21_0.Y.n9 two_stage_opamp_dummy_magic_21_0.Y.n7 4.8755
R6153 two_stage_opamp_dummy_magic_21_0.Y.n12 two_stage_opamp_dummy_magic_21_0.Y.n2 4.8755
R6154 two_stage_opamp_dummy_magic_21_0.Y.n18 two_stage_opamp_dummy_magic_21_0.Y.n17 4.8755
R6155 two_stage_opamp_dummy_magic_21_0.Y.n20 two_stage_opamp_dummy_magic_21_0.Y.n19 4.5005
R6156 two_stage_opamp_dummy_magic_21_0.Y.n62 two_stage_opamp_dummy_magic_21_0.Y.n61 4.5005
R6157 two_stage_opamp_dummy_magic_21_0.Y.n72 two_stage_opamp_dummy_magic_21_0.Y.n62 3.27133
R6158 two_stage_opamp_dummy_magic_21_0.Y.n41 two_stage_opamp_dummy_magic_21_0.Y.n22 0.792167
R6159 two_stage_opamp_dummy_magic_21_0.Y.n40 two_stage_opamp_dummy_magic_21_0.Y.n23 0.6255
R6160 two_stage_opamp_dummy_magic_21_0.Y.n30 two_stage_opamp_dummy_magic_21_0.Y.n23 0.6255
R6161 two_stage_opamp_dummy_magic_21_0.Y.n30 two_stage_opamp_dummy_magic_21_0.Y.n29 0.6255
R6162 two_stage_opamp_dummy_magic_21_0.Y.n33 two_stage_opamp_dummy_magic_21_0.Y.n24 0.6255
R6163 two_stage_opamp_dummy_magic_21_0.Y.n36 two_stage_opamp_dummy_magic_21_0.Y.n33 0.6255
R6164 two_stage_opamp_dummy_magic_21_0.Y.n37 two_stage_opamp_dummy_magic_21_0.Y.n36 0.6255
R6165 two_stage_opamp_dummy_magic_21_0.Y.n15 two_stage_opamp_dummy_magic_21_0.Y.n14 0.563
R6166 two_stage_opamp_dummy_magic_21_0.Y.n19 two_stage_opamp_dummy_magic_21_0.Y.n18 0.563
R6167 two_stage_opamp_dummy_magic_21_0.Y.n19 two_stage_opamp_dummy_magic_21_0.Y.n2 0.563
R6168 two_stage_opamp_dummy_magic_21_0.Y.n7 two_stage_opamp_dummy_magic_21_0.Y.n2 0.563
R6169 two_stage_opamp_dummy_magic_21_0.Y.n13 two_stage_opamp_dummy_magic_21_0.Y.n10 0.563
R6170 two_stage_opamp_dummy_magic_21_0.Y.n14 two_stage_opamp_dummy_magic_21_0.Y.n13 0.563
R6171 two_stage_opamp_dummy_magic_21_0.Y.n20 two_stage_opamp_dummy_magic_21_0.Y.n1 0.3755
R6172 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n0 345.264
R6173 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n1 344.7
R6174 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n3 292.5
R6175 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t0 122.442
R6176 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n7 118.861
R6177 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n9 118.861
R6178 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n13 118.861
R6179 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n16 118.861
R6180 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n19 118.861
R6181 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n2 52.763
R6182 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n4 51.7297
R6183 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n22 42.3755
R6184 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t15 39.4005
R6185 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t2 39.4005
R6186 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t4 39.4005
R6187 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t1 39.4005
R6188 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t3 39.4005
R6189 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t16 39.4005
R6190 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t9 19.7005
R6191 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t5 19.7005
R6192 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t8 19.7005
R6193 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t14 19.7005
R6194 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t12 19.7005
R6195 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t7 19.7005
R6196 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t11 19.7005
R6197 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t6 19.7005
R6198 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t10 19.7005
R6199 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t13 19.7005
R6200 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n21 6.28175
R6201 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n8 5.60467
R6202 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n18 5.54217
R6203 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n6 5.54217
R6204 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n10 5.04217
R6205 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n12 5.04217
R6206 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n5 5.04217
R6207 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n20 5.04217
R6208 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n6 4.97967
R6209 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n14 4.97967
R6210 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n17 4.97967
R6211 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n15 0.563
R6212 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n6 0.563
R6213 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n11 0.563
R6214 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n5 0.563
R6215 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n5 0.563
R6216 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R6217 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R6218 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R6219 bgr_0.Vin+.n5 bgr_0.Vin+.n3 227.169
R6220 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R6221 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R6222 bgr_0.Vin+.n2 bgr_0.Vin+.t10 174.726
R6223 bgr_0.Vin+.n7 bgr_0.Vin+.n6 168.435
R6224 bgr_0.Vin+.n5 bgr_0.Vin+.n4 168.435
R6225 bgr_0.Vin+.t4 bgr_0.Vin+.n8 158.989
R6226 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R6227 bgr_0.Vin+.n8 bgr_0.Vin+.t5 119.067
R6228 bgr_0.Vin+.n3 bgr_0.Vin+.t7 96.4005
R6229 bgr_0.Vin+.n8 bgr_0.Vin+.n7 35.0317
R6230 bgr_0.Vin+.n6 bgr_0.Vin+.t0 13.1338
R6231 bgr_0.Vin+.n6 bgr_0.Vin+.t3 13.1338
R6232 bgr_0.Vin+.n4 bgr_0.Vin+.t2 13.1338
R6233 bgr_0.Vin+.n4 bgr_0.Vin+.t1 13.1338
R6234 bgr_0.Vin+.n7 bgr_0.Vin+.n5 2.1255
R6235 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R6236 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R6237 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R6238 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R6239 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R6240 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R6241 bgr_0.V_mir1.n7 bgr_0.V_mir1.t0 278.312
R6242 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R6243 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R6244 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R6245 bgr_0.V_mir1.n11 bgr_0.V_mir1.t6 184.097
R6246 bgr_0.V_mir1.n2 bgr_0.V_mir1.t4 184.097
R6247 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R6248 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R6249 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R6250 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R6251 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R6252 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R6253 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 120.501
R6254 bgr_0.V_mir1.n17 bgr_0.V_mir1.t14 120.501
R6255 bgr_0.V_mir1.n9 bgr_0.V_mir1.t17 120.501
R6256 bgr_0.V_mir1.n10 bgr_0.V_mir1.t12 120.501
R6257 bgr_0.V_mir1.n0 bgr_0.V_mir1.t18 120.501
R6258 bgr_0.V_mir1.n1 bgr_0.V_mir1.t8 120.501
R6259 bgr_0.V_mir1.n6 bgr_0.V_mir1.t1 48.0005
R6260 bgr_0.V_mir1.n6 bgr_0.V_mir1.t3 48.0005
R6261 bgr_0.V_mir1.n5 bgr_0.V_mir1.t2 48.0005
R6262 bgr_0.V_mir1.n5 bgr_0.V_mir1.t16 48.0005
R6263 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R6264 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R6265 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R6266 bgr_0.V_mir1.n12 bgr_0.V_mir1.t7 39.4005
R6267 bgr_0.V_mir1.n12 bgr_0.V_mir1.t13 39.4005
R6268 bgr_0.V_mir1.n3 bgr_0.V_mir1.t5 39.4005
R6269 bgr_0.V_mir1.n3 bgr_0.V_mir1.t9 39.4005
R6270 bgr_0.V_mir1.n20 bgr_0.V_mir1.t11 39.4005
R6271 bgr_0.V_mir1.t15 bgr_0.V_mir1.n20 39.4005
R6272 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R6273 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R6274 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R6275 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R6276 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R6277 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R6278 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t13 354.854
R6279 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t21 346.8
R6280 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 339.522
R6281 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 339.522
R6282 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 335.022
R6283 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t7 275.909
R6284 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.n10 227.909
R6285 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n12 222.034
R6286 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t22 184.097
R6287 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t32 184.097
R6288 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t16 184.097
R6289 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t36 184.097
R6290 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n17 166.05
R6291 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n8 166.05
R6292 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n4 54.2759
R6293 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t10 48.0005
R6294 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t8 48.0005
R6295 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t9 48.0005
R6296 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t6 48.0005
R6297 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t4 39.4005
R6298 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t2 39.4005
R6299 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t0 39.4005
R6300 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 39.4005
R6301 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t5 39.4005
R6302 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t1 39.4005
R6303 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t11 4.8295
R6304 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t29 4.8295
R6305 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t31 4.8295
R6306 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R6307 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.8295
R6308 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.8295
R6309 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t30 4.8295
R6310 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t18 4.8295
R6311 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t23 4.8295
R6312 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t15 4.5005
R6313 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t35 4.5005
R6314 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t34 4.5005
R6315 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t28 4.5005
R6316 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t27 4.5005
R6317 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t19 4.5005
R6318 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t33 4.5005
R6319 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t26 4.5005
R6320 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t25 4.5005
R6321 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t17 4.5005
R6322 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t12 4.5005
R6323 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n11 4.5005
R6324 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n15 4.5005
R6325 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n18 1.3755
R6326 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n9 1.3755
R6327 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n5 1.188
R6328 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.8935
R6329 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n0 0.8935
R6330 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n13 0.78175
R6331 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.6585
R6332 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 0.6585
R6333 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n16 0.6255
R6334 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n7 0.6255
R6335 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n20 0.438
R6336 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t33 355.293
R6337 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t34 346.8
R6338 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 339.522
R6339 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n5 339.522
R6340 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n10 335.022
R6341 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t3 275.909
R6342 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.n7 227.909
R6343 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n9 222.034
R6344 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t13 184.097
R6345 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t24 184.097
R6346 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t16 184.097
R6347 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t27 184.097
R6348 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n11 166.05
R6349 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n6 166.05
R6350 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n4 52.9634
R6351 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t4 48.0005
R6352 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t1 48.0005
R6353 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t2 48.0005
R6354 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t8 48.0005
R6355 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t5 39.4005
R6356 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t10 39.4005
R6357 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t7 39.4005
R6358 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t9 39.4005
R6359 bgr_0.1st_Vout_2.t0 bgr_0.1st_Vout_2.n13 39.4005
R6360 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t6 39.4005
R6361 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n3 5.28175
R6362 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t17 4.8295
R6363 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t35 4.8295
R6364 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.8295
R6365 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t26 4.8295
R6366 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.8295
R6367 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.8295
R6368 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t36 4.8295
R6369 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.8295
R6370 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t18 4.8295
R6371 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n8 4.5005
R6372 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t12 4.5005
R6373 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t32 4.5005
R6374 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R6375 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t23 4.5005
R6376 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.5005
R6377 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t15 4.5005
R6378 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t29 4.5005
R6379 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t21 4.5005
R6380 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t28 4.5005
R6381 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R6382 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t14 4.5005
R6383 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 3.188
R6384 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 3.1025
R6385 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n1 2.0005
R6386 bgr_0.cap_res2.t0 bgr_0.cap_res2.t18 121.245
R6387 bgr_0.cap_res2.t13 bgr_0.cap_res2.t7 0.1603
R6388 bgr_0.cap_res2.t6 bgr_0.cap_res2.t1 0.1603
R6389 bgr_0.cap_res2.t11 bgr_0.cap_res2.t5 0.1603
R6390 bgr_0.cap_res2.t4 bgr_0.cap_res2.t20 0.1603
R6391 bgr_0.cap_res2.t19 bgr_0.cap_res2.t16 0.1603
R6392 bgr_0.cap_res2.n1 bgr_0.cap_res2.t3 0.159278
R6393 bgr_0.cap_res2.n2 bgr_0.cap_res2.t10 0.159278
R6394 bgr_0.cap_res2.n3 bgr_0.cap_res2.t17 0.159278
R6395 bgr_0.cap_res2.n4 bgr_0.cap_res2.t12 0.159278
R6396 bgr_0.cap_res2.n4 bgr_0.cap_res2.t15 0.1368
R6397 bgr_0.cap_res2.n4 bgr_0.cap_res2.t13 0.1368
R6398 bgr_0.cap_res2.n3 bgr_0.cap_res2.t9 0.1368
R6399 bgr_0.cap_res2.n3 bgr_0.cap_res2.t6 0.1368
R6400 bgr_0.cap_res2.n2 bgr_0.cap_res2.t14 0.1368
R6401 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.1368
R6402 bgr_0.cap_res2.n1 bgr_0.cap_res2.t8 0.1368
R6403 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R6404 bgr_0.cap_res2.n0 bgr_0.cap_res2.t2 0.1368
R6405 bgr_0.cap_res2.n0 bgr_0.cap_res2.t19 0.1368
R6406 bgr_0.cap_res2.t3 bgr_0.cap_res2.n0 0.00152174
R6407 bgr_0.cap_res2.t10 bgr_0.cap_res2.n1 0.00152174
R6408 bgr_0.cap_res2.t17 bgr_0.cap_res2.n2 0.00152174
R6409 bgr_0.cap_res2.t12 bgr_0.cap_res2.n3 0.00152174
R6410 bgr_0.cap_res2.t18 bgr_0.cap_res2.n4 0.00152174
R6411 two_stage_opamp_dummy_magic_21_0.V_source.n70 two_stage_opamp_dummy_magic_21_0.V_source.t4 66.2047
R6412 two_stage_opamp_dummy_magic_21_0.V_source.n1 two_stage_opamp_dummy_magic_21_0.V_source.n0 49.3505
R6413 two_stage_opamp_dummy_magic_21_0.V_source.n4 two_stage_opamp_dummy_magic_21_0.V_source.n3 49.3505
R6414 two_stage_opamp_dummy_magic_21_0.V_source.n7 two_stage_opamp_dummy_magic_21_0.V_source.n6 49.3505
R6415 two_stage_opamp_dummy_magic_21_0.V_source.n10 two_stage_opamp_dummy_magic_21_0.V_source.n9 49.3505
R6416 two_stage_opamp_dummy_magic_21_0.V_source.n14 two_stage_opamp_dummy_magic_21_0.V_source.n13 49.3505
R6417 two_stage_opamp_dummy_magic_21_0.V_source.n19 two_stage_opamp_dummy_magic_21_0.V_source.n18 49.3505
R6418 two_stage_opamp_dummy_magic_21_0.V_source.n21 two_stage_opamp_dummy_magic_21_0.V_source.n20 49.3505
R6419 two_stage_opamp_dummy_magic_21_0.V_source.n25 two_stage_opamp_dummy_magic_21_0.V_source.n24 49.3505
R6420 two_stage_opamp_dummy_magic_21_0.V_source.n28 two_stage_opamp_dummy_magic_21_0.V_source.n27 49.3505
R6421 two_stage_opamp_dummy_magic_21_0.V_source.n31 two_stage_opamp_dummy_magic_21_0.V_source.n30 49.3505
R6422 two_stage_opamp_dummy_magic_21_0.V_source.n39 two_stage_opamp_dummy_magic_21_0.V_source.n38 32.3838
R6423 two_stage_opamp_dummy_magic_21_0.V_source.n41 two_stage_opamp_dummy_magic_21_0.V_source.n40 32.3838
R6424 two_stage_opamp_dummy_magic_21_0.V_source.n47 two_stage_opamp_dummy_magic_21_0.V_source.n46 32.3838
R6425 two_stage_opamp_dummy_magic_21_0.V_source.n49 two_stage_opamp_dummy_magic_21_0.V_source.n48 32.3838
R6426 two_stage_opamp_dummy_magic_21_0.V_source.n53 two_stage_opamp_dummy_magic_21_0.V_source.n52 32.3838
R6427 two_stage_opamp_dummy_magic_21_0.V_source.n56 two_stage_opamp_dummy_magic_21_0.V_source.n55 32.3838
R6428 two_stage_opamp_dummy_magic_21_0.V_source.n60 two_stage_opamp_dummy_magic_21_0.V_source.n59 32.3838
R6429 two_stage_opamp_dummy_magic_21_0.V_source.n63 two_stage_opamp_dummy_magic_21_0.V_source.n62 32.3838
R6430 two_stage_opamp_dummy_magic_21_0.V_source.n67 two_stage_opamp_dummy_magic_21_0.V_source.n66 32.3838
R6431 two_stage_opamp_dummy_magic_21_0.V_source.n72 two_stage_opamp_dummy_magic_21_0.V_source.n71 32.3838
R6432 two_stage_opamp_dummy_magic_21_0.V_source.n0 two_stage_opamp_dummy_magic_21_0.V_source.t33 16.0005
R6433 two_stage_opamp_dummy_magic_21_0.V_source.n0 two_stage_opamp_dummy_magic_21_0.V_source.t39 16.0005
R6434 two_stage_opamp_dummy_magic_21_0.V_source.n3 two_stage_opamp_dummy_magic_21_0.V_source.t34 16.0005
R6435 two_stage_opamp_dummy_magic_21_0.V_source.n3 two_stage_opamp_dummy_magic_21_0.V_source.t40 16.0005
R6436 two_stage_opamp_dummy_magic_21_0.V_source.n6 two_stage_opamp_dummy_magic_21_0.V_source.t32 16.0005
R6437 two_stage_opamp_dummy_magic_21_0.V_source.n6 two_stage_opamp_dummy_magic_21_0.V_source.t1 16.0005
R6438 two_stage_opamp_dummy_magic_21_0.V_source.n9 two_stage_opamp_dummy_magic_21_0.V_source.t6 16.0005
R6439 two_stage_opamp_dummy_magic_21_0.V_source.n9 two_stage_opamp_dummy_magic_21_0.V_source.t27 16.0005
R6440 two_stage_opamp_dummy_magic_21_0.V_source.n13 two_stage_opamp_dummy_magic_21_0.V_source.t7 16.0005
R6441 two_stage_opamp_dummy_magic_21_0.V_source.n13 two_stage_opamp_dummy_magic_21_0.V_source.t5 16.0005
R6442 two_stage_opamp_dummy_magic_21_0.V_source.n18 two_stage_opamp_dummy_magic_21_0.V_source.t30 16.0005
R6443 two_stage_opamp_dummy_magic_21_0.V_source.n18 two_stage_opamp_dummy_magic_21_0.V_source.t36 16.0005
R6444 two_stage_opamp_dummy_magic_21_0.V_source.n20 two_stage_opamp_dummy_magic_21_0.V_source.t3 16.0005
R6445 two_stage_opamp_dummy_magic_21_0.V_source.n20 two_stage_opamp_dummy_magic_21_0.V_source.t38 16.0005
R6446 two_stage_opamp_dummy_magic_21_0.V_source.n24 two_stage_opamp_dummy_magic_21_0.V_source.t0 16.0005
R6447 two_stage_opamp_dummy_magic_21_0.V_source.n24 two_stage_opamp_dummy_magic_21_0.V_source.t28 16.0005
R6448 two_stage_opamp_dummy_magic_21_0.V_source.n27 two_stage_opamp_dummy_magic_21_0.V_source.t2 16.0005
R6449 two_stage_opamp_dummy_magic_21_0.V_source.n27 two_stage_opamp_dummy_magic_21_0.V_source.t29 16.0005
R6450 two_stage_opamp_dummy_magic_21_0.V_source.n30 two_stage_opamp_dummy_magic_21_0.V_source.t31 16.0005
R6451 two_stage_opamp_dummy_magic_21_0.V_source.n30 two_stage_opamp_dummy_magic_21_0.V_source.t37 16.0005
R6452 two_stage_opamp_dummy_magic_21_0.V_source.n38 two_stage_opamp_dummy_magic_21_0.V_source.t35 9.6005
R6453 two_stage_opamp_dummy_magic_21_0.V_source.n38 two_stage_opamp_dummy_magic_21_0.V_source.t8 9.6005
R6454 two_stage_opamp_dummy_magic_21_0.V_source.n40 two_stage_opamp_dummy_magic_21_0.V_source.t25 9.6005
R6455 two_stage_opamp_dummy_magic_21_0.V_source.n40 two_stage_opamp_dummy_magic_21_0.V_source.t19 9.6005
R6456 two_stage_opamp_dummy_magic_21_0.V_source.n46 two_stage_opamp_dummy_magic_21_0.V_source.t12 9.6005
R6457 two_stage_opamp_dummy_magic_21_0.V_source.n46 two_stage_opamp_dummy_magic_21_0.V_source.t18 9.6005
R6458 two_stage_opamp_dummy_magic_21_0.V_source.n48 two_stage_opamp_dummy_magic_21_0.V_source.t14 9.6005
R6459 two_stage_opamp_dummy_magic_21_0.V_source.n48 two_stage_opamp_dummy_magic_21_0.V_source.t22 9.6005
R6460 two_stage_opamp_dummy_magic_21_0.V_source.n52 two_stage_opamp_dummy_magic_21_0.V_source.t16 9.6005
R6461 two_stage_opamp_dummy_magic_21_0.V_source.n52 two_stage_opamp_dummy_magic_21_0.V_source.t24 9.6005
R6462 two_stage_opamp_dummy_magic_21_0.V_source.n55 two_stage_opamp_dummy_magic_21_0.V_source.t20 9.6005
R6463 two_stage_opamp_dummy_magic_21_0.V_source.n55 two_stage_opamp_dummy_magic_21_0.V_source.t10 9.6005
R6464 two_stage_opamp_dummy_magic_21_0.V_source.n59 two_stage_opamp_dummy_magic_21_0.V_source.t17 9.6005
R6465 two_stage_opamp_dummy_magic_21_0.V_source.n59 two_stage_opamp_dummy_magic_21_0.V_source.t9 9.6005
R6466 two_stage_opamp_dummy_magic_21_0.V_source.n62 two_stage_opamp_dummy_magic_21_0.V_source.t21 9.6005
R6467 two_stage_opamp_dummy_magic_21_0.V_source.n62 two_stage_opamp_dummy_magic_21_0.V_source.t11 9.6005
R6468 two_stage_opamp_dummy_magic_21_0.V_source.n66 two_stage_opamp_dummy_magic_21_0.V_source.t23 9.6005
R6469 two_stage_opamp_dummy_magic_21_0.V_source.n66 two_stage_opamp_dummy_magic_21_0.V_source.t13 9.6005
R6470 two_stage_opamp_dummy_magic_21_0.V_source.t26 two_stage_opamp_dummy_magic_21_0.V_source.n72 9.6005
R6471 two_stage_opamp_dummy_magic_21_0.V_source.n72 two_stage_opamp_dummy_magic_21_0.V_source.t15 9.6005
R6472 two_stage_opamp_dummy_magic_21_0.V_source.n47 two_stage_opamp_dummy_magic_21_0.V_source.n45 5.89633
R6473 two_stage_opamp_dummy_magic_21_0.V_source.n39 two_stage_opamp_dummy_magic_21_0.V_source.n36 5.89633
R6474 two_stage_opamp_dummy_magic_21_0.V_source.n50 two_stage_opamp_dummy_magic_21_0.V_source.n47 5.70883
R6475 two_stage_opamp_dummy_magic_21_0.V_source.n42 two_stage_opamp_dummy_magic_21_0.V_source.n39 5.70883
R6476 two_stage_opamp_dummy_magic_21_0.V_source.n22 two_stage_opamp_dummy_magic_21_0.V_source.n19 5.6255
R6477 two_stage_opamp_dummy_magic_21_0.V_source.n5 two_stage_opamp_dummy_magic_21_0.V_source.n4 5.6255
R6478 two_stage_opamp_dummy_magic_21_0.V_source.n31 two_stage_opamp_dummy_magic_21_0.V_source.n29 5.45883
R6479 two_stage_opamp_dummy_magic_21_0.V_source.n19 two_stage_opamp_dummy_magic_21_0.V_source.n17 5.45883
R6480 two_stage_opamp_dummy_magic_21_0.V_source.n8 two_stage_opamp_dummy_magic_21_0.V_source.n4 5.45883
R6481 two_stage_opamp_dummy_magic_21_0.V_source.n12 two_stage_opamp_dummy_magic_21_0.V_source.n1 5.45883
R6482 two_stage_opamp_dummy_magic_21_0.V_source.n41 two_stage_opamp_dummy_magic_21_0.V_source.n36 5.33383
R6483 two_stage_opamp_dummy_magic_21_0.V_source.n49 two_stage_opamp_dummy_magic_21_0.V_source.n45 5.33383
R6484 two_stage_opamp_dummy_magic_21_0.V_source.n54 two_stage_opamp_dummy_magic_21_0.V_source.n53 5.33383
R6485 two_stage_opamp_dummy_magic_21_0.V_source.n57 two_stage_opamp_dummy_magic_21_0.V_source.n56 5.33383
R6486 two_stage_opamp_dummy_magic_21_0.V_source.n60 two_stage_opamp_dummy_magic_21_0.V_source.n58 5.33383
R6487 two_stage_opamp_dummy_magic_21_0.V_source.n63 two_stage_opamp_dummy_magic_21_0.V_source.n37 5.33383
R6488 two_stage_opamp_dummy_magic_21_0.V_source.n68 two_stage_opamp_dummy_magic_21_0.V_source.n67 5.33383
R6489 two_stage_opamp_dummy_magic_21_0.V_source.n42 two_stage_opamp_dummy_magic_21_0.V_source.n41 5.14633
R6490 two_stage_opamp_dummy_magic_21_0.V_source.n50 two_stage_opamp_dummy_magic_21_0.V_source.n49 5.14633
R6491 two_stage_opamp_dummy_magic_21_0.V_source.n53 two_stage_opamp_dummy_magic_21_0.V_source.n51 5.14633
R6492 two_stage_opamp_dummy_magic_21_0.V_source.n56 two_stage_opamp_dummy_magic_21_0.V_source.n44 5.14633
R6493 two_stage_opamp_dummy_magic_21_0.V_source.n61 two_stage_opamp_dummy_magic_21_0.V_source.n60 5.14633
R6494 two_stage_opamp_dummy_magic_21_0.V_source.n64 two_stage_opamp_dummy_magic_21_0.V_source.n63 5.14633
R6495 two_stage_opamp_dummy_magic_21_0.V_source.n67 two_stage_opamp_dummy_magic_21_0.V_source.n65 5.14633
R6496 two_stage_opamp_dummy_magic_21_0.V_source.n7 two_stage_opamp_dummy_magic_21_0.V_source.n5 5.063
R6497 two_stage_opamp_dummy_magic_21_0.V_source.n10 two_stage_opamp_dummy_magic_21_0.V_source.n2 5.063
R6498 two_stage_opamp_dummy_magic_21_0.V_source.n15 two_stage_opamp_dummy_magic_21_0.V_source.n14 5.063
R6499 two_stage_opamp_dummy_magic_21_0.V_source.n22 two_stage_opamp_dummy_magic_21_0.V_source.n21 5.063
R6500 two_stage_opamp_dummy_magic_21_0.V_source.n25 two_stage_opamp_dummy_magic_21_0.V_source.n23 5.063
R6501 two_stage_opamp_dummy_magic_21_0.V_source.n28 two_stage_opamp_dummy_magic_21_0.V_source.n16 5.063
R6502 two_stage_opamp_dummy_magic_21_0.V_source.n32 two_stage_opamp_dummy_magic_21_0.V_source.n31 5.063
R6503 two_stage_opamp_dummy_magic_21_0.V_source.n8 two_stage_opamp_dummy_magic_21_0.V_source.n7 4.89633
R6504 two_stage_opamp_dummy_magic_21_0.V_source.n11 two_stage_opamp_dummy_magic_21_0.V_source.n10 4.89633
R6505 two_stage_opamp_dummy_magic_21_0.V_source.n14 two_stage_opamp_dummy_magic_21_0.V_source.n12 4.89633
R6506 two_stage_opamp_dummy_magic_21_0.V_source.n21 two_stage_opamp_dummy_magic_21_0.V_source.n17 4.89633
R6507 two_stage_opamp_dummy_magic_21_0.V_source.n26 two_stage_opamp_dummy_magic_21_0.V_source.n25 4.89633
R6508 two_stage_opamp_dummy_magic_21_0.V_source.n29 two_stage_opamp_dummy_magic_21_0.V_source.n28 4.89633
R6509 two_stage_opamp_dummy_magic_21_0.V_source.n34 two_stage_opamp_dummy_magic_21_0.V_source.n33 4.5005
R6510 two_stage_opamp_dummy_magic_21_0.V_source.n43 two_stage_opamp_dummy_magic_21_0.V_source.n35 4.5005
R6511 two_stage_opamp_dummy_magic_21_0.V_source.n70 two_stage_opamp_dummy_magic_21_0.V_source.n69 4.5005
R6512 two_stage_opamp_dummy_magic_21_0.V_source.n33 two_stage_opamp_dummy_magic_21_0.V_source.n32 3.6255
R6513 two_stage_opamp_dummy_magic_21_0.V_source.n35 two_stage_opamp_dummy_magic_21_0.V_source.n34 1.738
R6514 two_stage_opamp_dummy_magic_21_0.V_source.n71 two_stage_opamp_dummy_magic_21_0.V_source.n70 0.833833
R6515 two_stage_opamp_dummy_magic_21_0.V_source.n71 two_stage_opamp_dummy_magic_21_0.V_source.n35 0.633833
R6516 two_stage_opamp_dummy_magic_21_0.V_source.n29 two_stage_opamp_dummy_magic_21_0.V_source.n26 0.563
R6517 two_stage_opamp_dummy_magic_21_0.V_source.n26 two_stage_opamp_dummy_magic_21_0.V_source.n17 0.563
R6518 two_stage_opamp_dummy_magic_21_0.V_source.n23 two_stage_opamp_dummy_magic_21_0.V_source.n22 0.563
R6519 two_stage_opamp_dummy_magic_21_0.V_source.n23 two_stage_opamp_dummy_magic_21_0.V_source.n16 0.563
R6520 two_stage_opamp_dummy_magic_21_0.V_source.n32 two_stage_opamp_dummy_magic_21_0.V_source.n16 0.563
R6521 two_stage_opamp_dummy_magic_21_0.V_source.n33 two_stage_opamp_dummy_magic_21_0.V_source.n15 0.563
R6522 two_stage_opamp_dummy_magic_21_0.V_source.n15 two_stage_opamp_dummy_magic_21_0.V_source.n2 0.563
R6523 two_stage_opamp_dummy_magic_21_0.V_source.n5 two_stage_opamp_dummy_magic_21_0.V_source.n2 0.563
R6524 two_stage_opamp_dummy_magic_21_0.V_source.n11 two_stage_opamp_dummy_magic_21_0.V_source.n8 0.563
R6525 two_stage_opamp_dummy_magic_21_0.V_source.n12 two_stage_opamp_dummy_magic_21_0.V_source.n11 0.563
R6526 two_stage_opamp_dummy_magic_21_0.V_source.n34 two_stage_opamp_dummy_magic_21_0.V_source.n1 0.563
R6527 two_stage_opamp_dummy_magic_21_0.V_source.n69 two_stage_opamp_dummy_magic_21_0.V_source.n68 0.563
R6528 two_stage_opamp_dummy_magic_21_0.V_source.n68 two_stage_opamp_dummy_magic_21_0.V_source.n37 0.563
R6529 two_stage_opamp_dummy_magic_21_0.V_source.n58 two_stage_opamp_dummy_magic_21_0.V_source.n37 0.563
R6530 two_stage_opamp_dummy_magic_21_0.V_source.n58 two_stage_opamp_dummy_magic_21_0.V_source.n57 0.563
R6531 two_stage_opamp_dummy_magic_21_0.V_source.n57 two_stage_opamp_dummy_magic_21_0.V_source.n54 0.563
R6532 two_stage_opamp_dummy_magic_21_0.V_source.n54 two_stage_opamp_dummy_magic_21_0.V_source.n45 0.563
R6533 two_stage_opamp_dummy_magic_21_0.V_source.n51 two_stage_opamp_dummy_magic_21_0.V_source.n50 0.563
R6534 two_stage_opamp_dummy_magic_21_0.V_source.n51 two_stage_opamp_dummy_magic_21_0.V_source.n44 0.563
R6535 two_stage_opamp_dummy_magic_21_0.V_source.n61 two_stage_opamp_dummy_magic_21_0.V_source.n44 0.563
R6536 two_stage_opamp_dummy_magic_21_0.V_source.n64 two_stage_opamp_dummy_magic_21_0.V_source.n61 0.563
R6537 two_stage_opamp_dummy_magic_21_0.V_source.n65 two_stage_opamp_dummy_magic_21_0.V_source.n64 0.563
R6538 two_stage_opamp_dummy_magic_21_0.V_source.n65 two_stage_opamp_dummy_magic_21_0.V_source.n43 0.563
R6539 two_stage_opamp_dummy_magic_21_0.V_source.n43 two_stage_opamp_dummy_magic_21_0.V_source.n42 0.563
R6540 two_stage_opamp_dummy_magic_21_0.V_source.n69 two_stage_opamp_dummy_magic_21_0.V_source.n36 0.563
R6541 two_stage_opamp_dummy_magic_21_0.Vb2.n23 two_stage_opamp_dummy_magic_21_0.Vb2.t27 746.673
R6542 two_stage_opamp_dummy_magic_21_0.Vb2.n1 two_stage_opamp_dummy_magic_21_0.Vb2.t0 721.625
R6543 two_stage_opamp_dummy_magic_21_0.Vb2.n16 two_stage_opamp_dummy_magic_21_0.Vb2.t17 611.739
R6544 two_stage_opamp_dummy_magic_21_0.Vb2.n12 two_stage_opamp_dummy_magic_21_0.Vb2.t29 611.739
R6545 two_stage_opamp_dummy_magic_21_0.Vb2.n7 two_stage_opamp_dummy_magic_21_0.Vb2.t32 611.739
R6546 two_stage_opamp_dummy_magic_21_0.Vb2.n3 two_stage_opamp_dummy_magic_21_0.Vb2.t22 611.739
R6547 two_stage_opamp_dummy_magic_21_0.Vb2.n2 two_stage_opamp_dummy_magic_21_0.Vb2.t13 563.451
R6548 two_stage_opamp_dummy_magic_21_0.Vb2.n16 two_stage_opamp_dummy_magic_21_0.Vb2.t15 421.75
R6549 two_stage_opamp_dummy_magic_21_0.Vb2.n17 two_stage_opamp_dummy_magic_21_0.Vb2.t12 421.75
R6550 two_stage_opamp_dummy_magic_21_0.Vb2.n18 two_stage_opamp_dummy_magic_21_0.Vb2.t30 421.75
R6551 two_stage_opamp_dummy_magic_21_0.Vb2.n19 two_stage_opamp_dummy_magic_21_0.Vb2.t24 421.75
R6552 two_stage_opamp_dummy_magic_21_0.Vb2.n12 two_stage_opamp_dummy_magic_21_0.Vb2.t11 421.75
R6553 two_stage_opamp_dummy_magic_21_0.Vb2.n13 two_stage_opamp_dummy_magic_21_0.Vb2.t14 421.75
R6554 two_stage_opamp_dummy_magic_21_0.Vb2.n14 two_stage_opamp_dummy_magic_21_0.Vb2.t16 421.75
R6555 two_stage_opamp_dummy_magic_21_0.Vb2.n15 two_stage_opamp_dummy_magic_21_0.Vb2.t19 421.75
R6556 two_stage_opamp_dummy_magic_21_0.Vb2.n7 two_stage_opamp_dummy_magic_21_0.Vb2.t26 421.75
R6557 two_stage_opamp_dummy_magic_21_0.Vb2.n8 two_stage_opamp_dummy_magic_21_0.Vb2.t21 421.75
R6558 two_stage_opamp_dummy_magic_21_0.Vb2.n9 two_stage_opamp_dummy_magic_21_0.Vb2.t23 421.75
R6559 two_stage_opamp_dummy_magic_21_0.Vb2.n10 two_stage_opamp_dummy_magic_21_0.Vb2.t20 421.75
R6560 two_stage_opamp_dummy_magic_21_0.Vb2.n3 two_stage_opamp_dummy_magic_21_0.Vb2.t28 421.75
R6561 two_stage_opamp_dummy_magic_21_0.Vb2.n4 two_stage_opamp_dummy_magic_21_0.Vb2.t25 421.75
R6562 two_stage_opamp_dummy_magic_21_0.Vb2.n5 two_stage_opamp_dummy_magic_21_0.Vb2.t31 421.75
R6563 two_stage_opamp_dummy_magic_21_0.Vb2.n6 two_stage_opamp_dummy_magic_21_0.Vb2.t18 421.75
R6564 two_stage_opamp_dummy_magic_21_0.Vb2.n21 two_stage_opamp_dummy_magic_21_0.Vb2.n11 313.776
R6565 two_stage_opamp_dummy_magic_21_0.Vb2.n21 two_stage_opamp_dummy_magic_21_0.Vb2.n20 313.212
R6566 two_stage_opamp_dummy_magic_21_0.Vb2.n17 two_stage_opamp_dummy_magic_21_0.Vb2.n16 167.094
R6567 two_stage_opamp_dummy_magic_21_0.Vb2.n18 two_stage_opamp_dummy_magic_21_0.Vb2.n17 167.094
R6568 two_stage_opamp_dummy_magic_21_0.Vb2.n19 two_stage_opamp_dummy_magic_21_0.Vb2.n18 167.094
R6569 two_stage_opamp_dummy_magic_21_0.Vb2.n13 two_stage_opamp_dummy_magic_21_0.Vb2.n12 167.094
R6570 two_stage_opamp_dummy_magic_21_0.Vb2.n14 two_stage_opamp_dummy_magic_21_0.Vb2.n13 167.094
R6571 two_stage_opamp_dummy_magic_21_0.Vb2.n15 two_stage_opamp_dummy_magic_21_0.Vb2.n14 167.094
R6572 two_stage_opamp_dummy_magic_21_0.Vb2.n8 two_stage_opamp_dummy_magic_21_0.Vb2.n7 167.094
R6573 two_stage_opamp_dummy_magic_21_0.Vb2.n9 two_stage_opamp_dummy_magic_21_0.Vb2.n8 167.094
R6574 two_stage_opamp_dummy_magic_21_0.Vb2.n10 two_stage_opamp_dummy_magic_21_0.Vb2.n9 167.094
R6575 two_stage_opamp_dummy_magic_21_0.Vb2.n4 two_stage_opamp_dummy_magic_21_0.Vb2.n3 167.094
R6576 two_stage_opamp_dummy_magic_21_0.Vb2.n5 two_stage_opamp_dummy_magic_21_0.Vb2.n4 167.094
R6577 two_stage_opamp_dummy_magic_21_0.Vb2.n6 two_stage_opamp_dummy_magic_21_0.Vb2.n5 167.094
R6578 two_stage_opamp_dummy_magic_21_0.Vb2.n29 two_stage_opamp_dummy_magic_21_0.Vb2.n28 140.857
R6579 two_stage_opamp_dummy_magic_21_0.Vb2.n27 two_stage_opamp_dummy_magic_21_0.Vb2.n26 139.608
R6580 two_stage_opamp_dummy_magic_21_0.Vb2.n25 two_stage_opamp_dummy_magic_21_0.Vb2.n24 139.608
R6581 two_stage_opamp_dummy_magic_21_0.Vb2.n30 two_stage_opamp_dummy_magic_21_0.Vb2.n29 139.608
R6582 two_stage_opamp_dummy_magic_21_0.Vb2.n1 two_stage_opamp_dummy_magic_21_0.Vb2.n0 67.013
R6583 two_stage_opamp_dummy_magic_21_0.Vb2.n25 two_stage_opamp_dummy_magic_21_0.Vb2.n23 60.7286
R6584 two_stage_opamp_dummy_magic_21_0.Vb2.n20 two_stage_opamp_dummy_magic_21_0.Vb2.n19 35.3472
R6585 two_stage_opamp_dummy_magic_21_0.Vb2.n20 two_stage_opamp_dummy_magic_21_0.Vb2.n15 35.3472
R6586 two_stage_opamp_dummy_magic_21_0.Vb2.n11 two_stage_opamp_dummy_magic_21_0.Vb2.n10 35.3472
R6587 two_stage_opamp_dummy_magic_21_0.Vb2.n11 two_stage_opamp_dummy_magic_21_0.Vb2.n6 35.3472
R6588 two_stage_opamp_dummy_magic_21_0.Vb2.n28 two_stage_opamp_dummy_magic_21_0.Vb2.t6 24.0005
R6589 two_stage_opamp_dummy_magic_21_0.Vb2.n28 two_stage_opamp_dummy_magic_21_0.Vb2.t8 24.0005
R6590 two_stage_opamp_dummy_magic_21_0.Vb2.n26 two_stage_opamp_dummy_magic_21_0.Vb2.t4 24.0005
R6591 two_stage_opamp_dummy_magic_21_0.Vb2.n26 two_stage_opamp_dummy_magic_21_0.Vb2.t2 24.0005
R6592 two_stage_opamp_dummy_magic_21_0.Vb2.n24 two_stage_opamp_dummy_magic_21_0.Vb2.t9 24.0005
R6593 two_stage_opamp_dummy_magic_21_0.Vb2.n24 two_stage_opamp_dummy_magic_21_0.Vb2.t3 24.0005
R6594 two_stage_opamp_dummy_magic_21_0.Vb2.n30 two_stage_opamp_dummy_magic_21_0.Vb2.t5 24.0005
R6595 two_stage_opamp_dummy_magic_21_0.Vb2.t7 two_stage_opamp_dummy_magic_21_0.Vb2.n30 24.0005
R6596 two_stage_opamp_dummy_magic_21_0.Vb2.n22 two_stage_opamp_dummy_magic_21_0.Vb2.n21 13.2817
R6597 two_stage_opamp_dummy_magic_21_0.Vb2.n0 two_stage_opamp_dummy_magic_21_0.Vb2.t1 11.2576
R6598 two_stage_opamp_dummy_magic_21_0.Vb2.n0 two_stage_opamp_dummy_magic_21_0.Vb2.t10 11.2576
R6599 two_stage_opamp_dummy_magic_21_0.Vb2.n29 two_stage_opamp_dummy_magic_21_0.Vb2.n27 7.563
R6600 two_stage_opamp_dummy_magic_21_0.Vb2.n2 two_stage_opamp_dummy_magic_21_0.Vb2.n1 7.35988
R6601 two_stage_opamp_dummy_magic_21_0.Vb2.n23 two_stage_opamp_dummy_magic_21_0.Vb2.n22 4.55362
R6602 two_stage_opamp_dummy_magic_21_0.Vb2.n27 two_stage_opamp_dummy_magic_21_0.Vb2.n25 1.2505
R6603 two_stage_opamp_dummy_magic_21_0.Vb2.n22 two_stage_opamp_dummy_magic_21_0.Vb2.n2 1.14112
R6604 two_stage_opamp_dummy_magic_21_0.VD4.n10 two_stage_opamp_dummy_magic_21_0.VD4.t3 672.293
R6605 two_stage_opamp_dummy_magic_21_0.VD4.n13 two_stage_opamp_dummy_magic_21_0.VD4.t0 672.293
R6606 two_stage_opamp_dummy_magic_21_0.VD4.t4 two_stage_opamp_dummy_magic_21_0.VD4.n11 213.131
R6607 two_stage_opamp_dummy_magic_21_0.VD4.n12 two_stage_opamp_dummy_magic_21_0.VD4.t1 213.131
R6608 two_stage_opamp_dummy_magic_21_0.VD4.t14 two_stage_opamp_dummy_magic_21_0.VD4.t4 146.155
R6609 two_stage_opamp_dummy_magic_21_0.VD4.t18 two_stage_opamp_dummy_magic_21_0.VD4.t14 146.155
R6610 two_stage_opamp_dummy_magic_21_0.VD4.t22 two_stage_opamp_dummy_magic_21_0.VD4.t18 146.155
R6611 two_stage_opamp_dummy_magic_21_0.VD4.t6 two_stage_opamp_dummy_magic_21_0.VD4.t22 146.155
R6612 two_stage_opamp_dummy_magic_21_0.VD4.t10 two_stage_opamp_dummy_magic_21_0.VD4.t6 146.155
R6613 two_stage_opamp_dummy_magic_21_0.VD4.t12 two_stage_opamp_dummy_magic_21_0.VD4.t10 146.155
R6614 two_stage_opamp_dummy_magic_21_0.VD4.t16 two_stage_opamp_dummy_magic_21_0.VD4.t12 146.155
R6615 two_stage_opamp_dummy_magic_21_0.VD4.t20 two_stage_opamp_dummy_magic_21_0.VD4.t16 146.155
R6616 two_stage_opamp_dummy_magic_21_0.VD4.t24 two_stage_opamp_dummy_magic_21_0.VD4.t20 146.155
R6617 two_stage_opamp_dummy_magic_21_0.VD4.t8 two_stage_opamp_dummy_magic_21_0.VD4.t24 146.155
R6618 two_stage_opamp_dummy_magic_21_0.VD4.t1 two_stage_opamp_dummy_magic_21_0.VD4.t8 146.155
R6619 two_stage_opamp_dummy_magic_21_0.VD4.n11 two_stage_opamp_dummy_magic_21_0.VD4.t5 76.2576
R6620 two_stage_opamp_dummy_magic_21_0.VD4.n12 two_stage_opamp_dummy_magic_21_0.VD4.t2 76.2576
R6621 two_stage_opamp_dummy_magic_21_0.VD4.n3 two_stage_opamp_dummy_magic_21_0.VD4.n2 71.513
R6622 two_stage_opamp_dummy_magic_21_0.VD4.n5 two_stage_opamp_dummy_magic_21_0.VD4.n4 71.513
R6623 two_stage_opamp_dummy_magic_21_0.VD4.n7 two_stage_opamp_dummy_magic_21_0.VD4.n6 71.513
R6624 two_stage_opamp_dummy_magic_21_0.VD4.n9 two_stage_opamp_dummy_magic_21_0.VD4.n8 71.513
R6625 two_stage_opamp_dummy_magic_21_0.VD4.n1 two_stage_opamp_dummy_magic_21_0.VD4.n0 71.513
R6626 two_stage_opamp_dummy_magic_21_0.VD4.n18 two_stage_opamp_dummy_magic_21_0.VD4.n17 66.0338
R6627 two_stage_opamp_dummy_magic_21_0.VD4.n21 two_stage_opamp_dummy_magic_21_0.VD4.n20 66.0338
R6628 two_stage_opamp_dummy_magic_21_0.VD4.n24 two_stage_opamp_dummy_magic_21_0.VD4.n23 66.0338
R6629 two_stage_opamp_dummy_magic_21_0.VD4.n28 two_stage_opamp_dummy_magic_21_0.VD4.n27 66.0338
R6630 two_stage_opamp_dummy_magic_21_0.VD4.n31 two_stage_opamp_dummy_magic_21_0.VD4.n30 66.0338
R6631 two_stage_opamp_dummy_magic_21_0.VD4.n34 two_stage_opamp_dummy_magic_21_0.VD4.n33 66.0338
R6632 two_stage_opamp_dummy_magic_21_0.VD4.n2 two_stage_opamp_dummy_magic_21_0.VD4.t17 11.2576
R6633 two_stage_opamp_dummy_magic_21_0.VD4.n2 two_stage_opamp_dummy_magic_21_0.VD4.t21 11.2576
R6634 two_stage_opamp_dummy_magic_21_0.VD4.n4 two_stage_opamp_dummy_magic_21_0.VD4.t11 11.2576
R6635 two_stage_opamp_dummy_magic_21_0.VD4.n4 two_stage_opamp_dummy_magic_21_0.VD4.t13 11.2576
R6636 two_stage_opamp_dummy_magic_21_0.VD4.n6 two_stage_opamp_dummy_magic_21_0.VD4.t23 11.2576
R6637 two_stage_opamp_dummy_magic_21_0.VD4.n6 two_stage_opamp_dummy_magic_21_0.VD4.t7 11.2576
R6638 two_stage_opamp_dummy_magic_21_0.VD4.n8 two_stage_opamp_dummy_magic_21_0.VD4.t15 11.2576
R6639 two_stage_opamp_dummy_magic_21_0.VD4.n8 two_stage_opamp_dummy_magic_21_0.VD4.t19 11.2576
R6640 two_stage_opamp_dummy_magic_21_0.VD4.n17 two_stage_opamp_dummy_magic_21_0.VD4.t35 11.2576
R6641 two_stage_opamp_dummy_magic_21_0.VD4.n17 two_stage_opamp_dummy_magic_21_0.VD4.t37 11.2576
R6642 two_stage_opamp_dummy_magic_21_0.VD4.n20 two_stage_opamp_dummy_magic_21_0.VD4.t28 11.2576
R6643 two_stage_opamp_dummy_magic_21_0.VD4.n20 two_stage_opamp_dummy_magic_21_0.VD4.t32 11.2576
R6644 two_stage_opamp_dummy_magic_21_0.VD4.n23 two_stage_opamp_dummy_magic_21_0.VD4.t27 11.2576
R6645 two_stage_opamp_dummy_magic_21_0.VD4.n23 two_stage_opamp_dummy_magic_21_0.VD4.t30 11.2576
R6646 two_stage_opamp_dummy_magic_21_0.VD4.n27 two_stage_opamp_dummy_magic_21_0.VD4.t34 11.2576
R6647 two_stage_opamp_dummy_magic_21_0.VD4.n27 two_stage_opamp_dummy_magic_21_0.VD4.t26 11.2576
R6648 two_stage_opamp_dummy_magic_21_0.VD4.n30 two_stage_opamp_dummy_magic_21_0.VD4.t33 11.2576
R6649 two_stage_opamp_dummy_magic_21_0.VD4.n30 two_stage_opamp_dummy_magic_21_0.VD4.t31 11.2576
R6650 two_stage_opamp_dummy_magic_21_0.VD4.n33 two_stage_opamp_dummy_magic_21_0.VD4.t36 11.2576
R6651 two_stage_opamp_dummy_magic_21_0.VD4.n33 two_stage_opamp_dummy_magic_21_0.VD4.t29 11.2576
R6652 two_stage_opamp_dummy_magic_21_0.VD4.n0 two_stage_opamp_dummy_magic_21_0.VD4.t25 11.2576
R6653 two_stage_opamp_dummy_magic_21_0.VD4.n0 two_stage_opamp_dummy_magic_21_0.VD4.t9 11.2576
R6654 two_stage_opamp_dummy_magic_21_0.VD4 two_stage_opamp_dummy_magic_21_0.VD4.n35 8.59425
R6655 two_stage_opamp_dummy_magic_21_0.VD4.n10 two_stage_opamp_dummy_magic_21_0.VD4.n9 6.10467
R6656 two_stage_opamp_dummy_magic_21_0.VD4.n34 two_stage_opamp_dummy_magic_21_0.VD4.n32 5.91717
R6657 two_stage_opamp_dummy_magic_21_0.VD4.n19 two_stage_opamp_dummy_magic_21_0.VD4.n18 5.91717
R6658 two_stage_opamp_dummy_magic_21_0.VD4.n22 two_stage_opamp_dummy_magic_21_0.VD4.n18 5.91717
R6659 two_stage_opamp_dummy_magic_21_0.VD4.n14 two_stage_opamp_dummy_magic_21_0.VD4.n13 5.47967
R6660 two_stage_opamp_dummy_magic_21_0.VD4 two_stage_opamp_dummy_magic_21_0.VD4.n14 5.3755
R6661 two_stage_opamp_dummy_magic_21_0.VD4.n22 two_stage_opamp_dummy_magic_21_0.VD4.n21 5.29217
R6662 two_stage_opamp_dummy_magic_21_0.VD4.n21 two_stage_opamp_dummy_magic_21_0.VD4.n19 5.29217
R6663 two_stage_opamp_dummy_magic_21_0.VD4.n25 two_stage_opamp_dummy_magic_21_0.VD4.n24 5.29217
R6664 two_stage_opamp_dummy_magic_21_0.VD4.n24 two_stage_opamp_dummy_magic_21_0.VD4.n16 5.29217
R6665 two_stage_opamp_dummy_magic_21_0.VD4.n28 two_stage_opamp_dummy_magic_21_0.VD4.n26 5.29217
R6666 two_stage_opamp_dummy_magic_21_0.VD4.n29 two_stage_opamp_dummy_magic_21_0.VD4.n28 5.29217
R6667 two_stage_opamp_dummy_magic_21_0.VD4.n31 two_stage_opamp_dummy_magic_21_0.VD4.n15 5.29217
R6668 two_stage_opamp_dummy_magic_21_0.VD4.n32 two_stage_opamp_dummy_magic_21_0.VD4.n31 5.29217
R6669 two_stage_opamp_dummy_magic_21_0.VD4.n35 two_stage_opamp_dummy_magic_21_0.VD4.n34 5.29217
R6670 two_stage_opamp_dummy_magic_21_0.VD4.n13 two_stage_opamp_dummy_magic_21_0.VD4.n12 1.03383
R6671 two_stage_opamp_dummy_magic_21_0.VD4.n11 two_stage_opamp_dummy_magic_21_0.VD4.n10 1.03383
R6672 two_stage_opamp_dummy_magic_21_0.VD4.n32 two_stage_opamp_dummy_magic_21_0.VD4.n29 0.6255
R6673 two_stage_opamp_dummy_magic_21_0.VD4.n29 two_stage_opamp_dummy_magic_21_0.VD4.n16 0.6255
R6674 two_stage_opamp_dummy_magic_21_0.VD4.n19 two_stage_opamp_dummy_magic_21_0.VD4.n16 0.6255
R6675 two_stage_opamp_dummy_magic_21_0.VD4.n25 two_stage_opamp_dummy_magic_21_0.VD4.n22 0.6255
R6676 two_stage_opamp_dummy_magic_21_0.VD4.n26 two_stage_opamp_dummy_magic_21_0.VD4.n25 0.6255
R6677 two_stage_opamp_dummy_magic_21_0.VD4.n26 two_stage_opamp_dummy_magic_21_0.VD4.n15 0.6255
R6678 two_stage_opamp_dummy_magic_21_0.VD4.n35 two_stage_opamp_dummy_magic_21_0.VD4.n15 0.6255
R6679 two_stage_opamp_dummy_magic_21_0.VD4.n14 two_stage_opamp_dummy_magic_21_0.VD4.n1 0.6255
R6680 two_stage_opamp_dummy_magic_21_0.VD4.n9 two_stage_opamp_dummy_magic_21_0.VD4.n7 0.6255
R6681 two_stage_opamp_dummy_magic_21_0.VD4.n7 two_stage_opamp_dummy_magic_21_0.VD4.n5 0.6255
R6682 two_stage_opamp_dummy_magic_21_0.VD4.n5 two_stage_opamp_dummy_magic_21_0.VD4.n3 0.6255
R6683 two_stage_opamp_dummy_magic_21_0.VD4.n3 two_stage_opamp_dummy_magic_21_0.VD4.n1 0.6255
R6684 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.n3 526.183
R6685 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 514.134
R6686 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n0 360.586
R6687 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 303.259
R6688 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 210.169
R6689 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t3 174.726
R6690 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t7 174.726
R6691 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 174.726
R6692 bgr_0.V_CUR_REF_REG.t1 bgr_0.V_CUR_REF_REG.n5 153.474
R6693 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 128.534
R6694 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t6 96.4005
R6695 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t0 39.4005
R6696 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t2 39.4005
R6697 bgr_0.V_p_2.n1 bgr_0.V_p_2.n2 229.562
R6698 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R6699 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R6700 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R6701 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R6702 bgr_0.V_p_2.n0 bgr_0.V_p_2.t10 98.7279
R6703 bgr_0.V_p_2.n5 bgr_0.V_p_2.t6 48.0005
R6704 bgr_0.V_p_2.n5 bgr_0.V_p_2.t0 48.0005
R6705 bgr_0.V_p_2.n4 bgr_0.V_p_2.t3 48.0005
R6706 bgr_0.V_p_2.n4 bgr_0.V_p_2.t7 48.0005
R6707 bgr_0.V_p_2.n3 bgr_0.V_p_2.t8 48.0005
R6708 bgr_0.V_p_2.n3 bgr_0.V_p_2.t1 48.0005
R6709 bgr_0.V_p_2.n2 bgr_0.V_p_2.t9 48.0005
R6710 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R6711 bgr_0.V_p_2.t4 bgr_0.V_p_2.n6 48.0005
R6712 bgr_0.V_p_2.n6 bgr_0.V_p_2.t5 48.0005
R6713 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R6714 a_7460_23988.t0 a_7460_23988.t1 178.133
R6715 two_stage_opamp_dummy_magic_21_0.V_err_p.n6 two_stage_opamp_dummy_magic_21_0.V_err_p.n5 594.301
R6716 two_stage_opamp_dummy_magic_21_0.V_err_p.n4 two_stage_opamp_dummy_magic_21_0.V_err_p.n7 594.301
R6717 two_stage_opamp_dummy_magic_21_0.V_err_p.n9 two_stage_opamp_dummy_magic_21_0.V_err_p.n8 594.301
R6718 two_stage_opamp_dummy_magic_21_0.V_err_p.n13 two_stage_opamp_dummy_magic_21_0.V_err_p.n12 594.301
R6719 two_stage_opamp_dummy_magic_21_0.V_err_p.n16 two_stage_opamp_dummy_magic_21_0.V_err_p.n15 594.301
R6720 two_stage_opamp_dummy_magic_21_0.V_err_p.n19 two_stage_opamp_dummy_magic_21_0.V_err_p.n18 594.301
R6721 two_stage_opamp_dummy_magic_21_0.V_err_p.n23 two_stage_opamp_dummy_magic_21_0.V_err_p.n22 594.301
R6722 two_stage_opamp_dummy_magic_21_0.V_err_p.n3 two_stage_opamp_dummy_magic_21_0.V_err_p.n26 594.301
R6723 two_stage_opamp_dummy_magic_21_0.V_err_p.n28 two_stage_opamp_dummy_magic_21_0.V_err_p.n27 594.301
R6724 two_stage_opamp_dummy_magic_21_0.V_err_p.n30 two_stage_opamp_dummy_magic_21_0.V_err_p.n29 594.301
R6725 two_stage_opamp_dummy_magic_21_0.V_err_p.n33 two_stage_opamp_dummy_magic_21_0.V_err_p.n32 594.301
R6726 two_stage_opamp_dummy_magic_21_0.V_err_p.n5 two_stage_opamp_dummy_magic_21_0.V_err_p.t10 78.8005
R6727 two_stage_opamp_dummy_magic_21_0.V_err_p.n5 two_stage_opamp_dummy_magic_21_0.V_err_p.t13 78.8005
R6728 two_stage_opamp_dummy_magic_21_0.V_err_p.n7 two_stage_opamp_dummy_magic_21_0.V_err_p.t3 78.8005
R6729 two_stage_opamp_dummy_magic_21_0.V_err_p.n7 two_stage_opamp_dummy_magic_21_0.V_err_p.t2 78.8005
R6730 two_stage_opamp_dummy_magic_21_0.V_err_p.n8 two_stage_opamp_dummy_magic_21_0.V_err_p.t20 78.8005
R6731 two_stage_opamp_dummy_magic_21_0.V_err_p.n8 two_stage_opamp_dummy_magic_21_0.V_err_p.t1 78.8005
R6732 two_stage_opamp_dummy_magic_21_0.V_err_p.n12 two_stage_opamp_dummy_magic_21_0.V_err_p.t17 78.8005
R6733 two_stage_opamp_dummy_magic_21_0.V_err_p.n12 two_stage_opamp_dummy_magic_21_0.V_err_p.t19 78.8005
R6734 two_stage_opamp_dummy_magic_21_0.V_err_p.n15 two_stage_opamp_dummy_magic_21_0.V_err_p.t14 78.8005
R6735 two_stage_opamp_dummy_magic_21_0.V_err_p.n15 two_stage_opamp_dummy_magic_21_0.V_err_p.t5 78.8005
R6736 two_stage_opamp_dummy_magic_21_0.V_err_p.n18 two_stage_opamp_dummy_magic_21_0.V_err_p.t16 78.8005
R6737 two_stage_opamp_dummy_magic_21_0.V_err_p.n18 two_stage_opamp_dummy_magic_21_0.V_err_p.t4 78.8005
R6738 two_stage_opamp_dummy_magic_21_0.V_err_p.n22 two_stage_opamp_dummy_magic_21_0.V_err_p.t18 78.8005
R6739 two_stage_opamp_dummy_magic_21_0.V_err_p.n22 two_stage_opamp_dummy_magic_21_0.V_err_p.t12 78.8005
R6740 two_stage_opamp_dummy_magic_21_0.V_err_p.n26 two_stage_opamp_dummy_magic_21_0.V_err_p.t9 78.8005
R6741 two_stage_opamp_dummy_magic_21_0.V_err_p.n26 two_stage_opamp_dummy_magic_21_0.V_err_p.t6 78.8005
R6742 two_stage_opamp_dummy_magic_21_0.V_err_p.n27 two_stage_opamp_dummy_magic_21_0.V_err_p.t15 78.8005
R6743 two_stage_opamp_dummy_magic_21_0.V_err_p.n27 two_stage_opamp_dummy_magic_21_0.V_err_p.t7 78.8005
R6744 two_stage_opamp_dummy_magic_21_0.V_err_p.n29 two_stage_opamp_dummy_magic_21_0.V_err_p.t8 78.8005
R6745 two_stage_opamp_dummy_magic_21_0.V_err_p.n29 two_stage_opamp_dummy_magic_21_0.V_err_p.t0 78.8005
R6746 two_stage_opamp_dummy_magic_21_0.V_err_p.n33 two_stage_opamp_dummy_magic_21_0.V_err_p.t21 78.8005
R6747 two_stage_opamp_dummy_magic_21_0.V_err_p.t11 two_stage_opamp_dummy_magic_21_0.V_err_p.n33 78.8005
R6748 two_stage_opamp_dummy_magic_21_0.V_err_p.n17 two_stage_opamp_dummy_magic_21_0.V_err_p.n13 6.10467
R6749 two_stage_opamp_dummy_magic_21_0.V_err_p.n11 two_stage_opamp_dummy_magic_21_0.V_err_p.n9 6.10467
R6750 two_stage_opamp_dummy_magic_21_0.V_err_p.n14 two_stage_opamp_dummy_magic_21_0.V_err_p.n13 5.91717
R6751 two_stage_opamp_dummy_magic_21_0.V_err_p.n25 two_stage_opamp_dummy_magic_21_0.V_err_p.n9 5.91717
R6752 two_stage_opamp_dummy_magic_21_0.V_err_p.n6 two_stage_opamp_dummy_magic_21_0.V_err_p.n2 5.41717
R6753 two_stage_opamp_dummy_magic_21_0.V_err_p.n3 two_stage_opamp_dummy_magic_21_0.V_err_p.n0 5.22967
R6754 two_stage_opamp_dummy_magic_21_0.V_err_p.n31 two_stage_opamp_dummy_magic_21_0.V_err_p.n6 5.22967
R6755 two_stage_opamp_dummy_magic_21_0.V_err_p.n1 two_stage_opamp_dummy_magic_21_0.V_err_p.n3 5.063
R6756 two_stage_opamp_dummy_magic_21_0.V_err_p.n32 two_stage_opamp_dummy_magic_21_0.V_err_p.n2 4.85467
R6757 two_stage_opamp_dummy_magic_21_0.V_err_p.n17 two_stage_opamp_dummy_magic_21_0.V_err_p.n16 4.85467
R6758 two_stage_opamp_dummy_magic_21_0.V_err_p.n20 two_stage_opamp_dummy_magic_21_0.V_err_p.n19 4.85467
R6759 two_stage_opamp_dummy_magic_21_0.V_err_p.n23 two_stage_opamp_dummy_magic_21_0.V_err_p.n21 4.85467
R6760 two_stage_opamp_dummy_magic_21_0.V_err_p.n11 two_stage_opamp_dummy_magic_21_0.V_err_p.n4 4.85467
R6761 two_stage_opamp_dummy_magic_21_0.V_err_p.n1 two_stage_opamp_dummy_magic_21_0.V_err_p.n28 4.85467
R6762 two_stage_opamp_dummy_magic_21_0.V_err_p.n30 two_stage_opamp_dummy_magic_21_0.V_err_p.n2 4.85467
R6763 two_stage_opamp_dummy_magic_21_0.V_err_p.n16 two_stage_opamp_dummy_magic_21_0.V_err_p.n14 4.66717
R6764 two_stage_opamp_dummy_magic_21_0.V_err_p.n19 two_stage_opamp_dummy_magic_21_0.V_err_p.n10 4.66717
R6765 two_stage_opamp_dummy_magic_21_0.V_err_p.n24 two_stage_opamp_dummy_magic_21_0.V_err_p.n23 4.66717
R6766 two_stage_opamp_dummy_magic_21_0.V_err_p.n28 two_stage_opamp_dummy_magic_21_0.V_err_p.n0 4.66717
R6767 two_stage_opamp_dummy_magic_21_0.V_err_p.n0 two_stage_opamp_dummy_magic_21_0.V_err_p.n30 4.66717
R6768 two_stage_opamp_dummy_magic_21_0.V_err_p.n32 two_stage_opamp_dummy_magic_21_0.V_err_p.n31 4.66717
R6769 two_stage_opamp_dummy_magic_21_0.V_err_p.n4 two_stage_opamp_dummy_magic_21_0.V_err_p.n25 4.5005
R6770 two_stage_opamp_dummy_magic_21_0.V_err_p.n3 two_stage_opamp_dummy_magic_21_0.V_err_p.n4 1.44842
R6771 two_stage_opamp_dummy_magic_21_0.V_err_p.n21 two_stage_opamp_dummy_magic_21_0.V_err_p.n11 1.2505
R6772 two_stage_opamp_dummy_magic_21_0.V_err_p.n21 two_stage_opamp_dummy_magic_21_0.V_err_p.n20 1.2505
R6773 two_stage_opamp_dummy_magic_21_0.V_err_p.n20 two_stage_opamp_dummy_magic_21_0.V_err_p.n17 1.2505
R6774 two_stage_opamp_dummy_magic_21_0.V_err_p.n14 two_stage_opamp_dummy_magic_21_0.V_err_p.n10 1.2505
R6775 two_stage_opamp_dummy_magic_21_0.V_err_p.n24 two_stage_opamp_dummy_magic_21_0.V_err_p.n10 1.2505
R6776 two_stage_opamp_dummy_magic_21_0.V_err_p.n25 two_stage_opamp_dummy_magic_21_0.V_err_p.n24 1.2505
R6777 two_stage_opamp_dummy_magic_21_0.V_err_p.n2 two_stage_opamp_dummy_magic_21_0.V_err_p.n1 1.1255
R6778 two_stage_opamp_dummy_magic_21_0.V_err_p.n31 two_stage_opamp_dummy_magic_21_0.V_err_p.n0 1.1255
R6779 two_stage_opamp_dummy_magic_21_0.X.n27 two_stage_opamp_dummy_magic_21_0.X.t33 1172.87
R6780 two_stage_opamp_dummy_magic_21_0.X.n21 two_stage_opamp_dummy_magic_21_0.X.t25 1172.87
R6781 two_stage_opamp_dummy_magic_21_0.X.n27 two_stage_opamp_dummy_magic_21_0.X.t48 996.134
R6782 two_stage_opamp_dummy_magic_21_0.X.n28 two_stage_opamp_dummy_magic_21_0.X.t35 996.134
R6783 two_stage_opamp_dummy_magic_21_0.X.n26 two_stage_opamp_dummy_magic_21_0.X.t50 996.134
R6784 two_stage_opamp_dummy_magic_21_0.X.n25 two_stage_opamp_dummy_magic_21_0.X.t38 996.134
R6785 two_stage_opamp_dummy_magic_21_0.X.n24 two_stage_opamp_dummy_magic_21_0.X.t53 996.134
R6786 two_stage_opamp_dummy_magic_21_0.X.n23 two_stage_opamp_dummy_magic_21_0.X.t40 996.134
R6787 two_stage_opamp_dummy_magic_21_0.X.n22 two_stage_opamp_dummy_magic_21_0.X.t26 996.134
R6788 two_stage_opamp_dummy_magic_21_0.X.n21 two_stage_opamp_dummy_magic_21_0.X.t39 996.134
R6789 two_stage_opamp_dummy_magic_21_0.X.n62 two_stage_opamp_dummy_magic_21_0.X.t28 690.867
R6790 two_stage_opamp_dummy_magic_21_0.X.n61 two_stage_opamp_dummy_magic_21_0.X.t51 690.867
R6791 two_stage_opamp_dummy_magic_21_0.X.n53 two_stage_opamp_dummy_magic_21_0.X.t54 530.201
R6792 two_stage_opamp_dummy_magic_21_0.X.n52 two_stage_opamp_dummy_magic_21_0.X.t46 530.201
R6793 two_stage_opamp_dummy_magic_21_0.X.n68 two_stage_opamp_dummy_magic_21_0.X.t52 514.134
R6794 two_stage_opamp_dummy_magic_21_0.X.n67 two_stage_opamp_dummy_magic_21_0.X.t37 514.134
R6795 two_stage_opamp_dummy_magic_21_0.X.n66 two_stage_opamp_dummy_magic_21_0.X.t49 514.134
R6796 two_stage_opamp_dummy_magic_21_0.X.n65 two_stage_opamp_dummy_magic_21_0.X.t34 514.134
R6797 two_stage_opamp_dummy_magic_21_0.X.n64 two_stage_opamp_dummy_magic_21_0.X.t45 514.134
R6798 two_stage_opamp_dummy_magic_21_0.X.n63 two_stage_opamp_dummy_magic_21_0.X.t30 514.134
R6799 two_stage_opamp_dummy_magic_21_0.X.n62 two_stage_opamp_dummy_magic_21_0.X.t43 514.134
R6800 two_stage_opamp_dummy_magic_21_0.X.n61 two_stage_opamp_dummy_magic_21_0.X.t36 514.134
R6801 two_stage_opamp_dummy_magic_21_0.X.n53 two_stage_opamp_dummy_magic_21_0.X.t41 353.467
R6802 two_stage_opamp_dummy_magic_21_0.X.n54 two_stage_opamp_dummy_magic_21_0.X.t27 353.467
R6803 two_stage_opamp_dummy_magic_21_0.X.n55 two_stage_opamp_dummy_magic_21_0.X.t42 353.467
R6804 two_stage_opamp_dummy_magic_21_0.X.n56 two_stage_opamp_dummy_magic_21_0.X.t29 353.467
R6805 two_stage_opamp_dummy_magic_21_0.X.n57 two_stage_opamp_dummy_magic_21_0.X.t44 353.467
R6806 two_stage_opamp_dummy_magic_21_0.X.n58 two_stage_opamp_dummy_magic_21_0.X.t32 353.467
R6807 two_stage_opamp_dummy_magic_21_0.X.n59 two_stage_opamp_dummy_magic_21_0.X.t47 353.467
R6808 two_stage_opamp_dummy_magic_21_0.X.n52 two_stage_opamp_dummy_magic_21_0.X.t31 353.467
R6809 two_stage_opamp_dummy_magic_21_0.X.n30 two_stage_opamp_dummy_magic_21_0.X.n29 304.375
R6810 two_stage_opamp_dummy_magic_21_0.X.n70 two_stage_opamp_dummy_magic_21_0.X.n60 216.9
R6811 two_stage_opamp_dummy_magic_21_0.X.n70 two_stage_opamp_dummy_magic_21_0.X.n69 216.9
R6812 two_stage_opamp_dummy_magic_21_0.X.n26 two_stage_opamp_dummy_magic_21_0.X.n25 176.733
R6813 two_stage_opamp_dummy_magic_21_0.X.n25 two_stage_opamp_dummy_magic_21_0.X.n24 176.733
R6814 two_stage_opamp_dummy_magic_21_0.X.n24 two_stage_opamp_dummy_magic_21_0.X.n23 176.733
R6815 two_stage_opamp_dummy_magic_21_0.X.n23 two_stage_opamp_dummy_magic_21_0.X.n22 176.733
R6816 two_stage_opamp_dummy_magic_21_0.X.n22 two_stage_opamp_dummy_magic_21_0.X.n21 176.733
R6817 two_stage_opamp_dummy_magic_21_0.X.n28 two_stage_opamp_dummy_magic_21_0.X.n27 176.733
R6818 two_stage_opamp_dummy_magic_21_0.X.n54 two_stage_opamp_dummy_magic_21_0.X.n53 176.733
R6819 two_stage_opamp_dummy_magic_21_0.X.n55 two_stage_opamp_dummy_magic_21_0.X.n54 176.733
R6820 two_stage_opamp_dummy_magic_21_0.X.n56 two_stage_opamp_dummy_magic_21_0.X.n55 176.733
R6821 two_stage_opamp_dummy_magic_21_0.X.n57 two_stage_opamp_dummy_magic_21_0.X.n56 176.733
R6822 two_stage_opamp_dummy_magic_21_0.X.n58 two_stage_opamp_dummy_magic_21_0.X.n57 176.733
R6823 two_stage_opamp_dummy_magic_21_0.X.n59 two_stage_opamp_dummy_magic_21_0.X.n58 176.733
R6824 two_stage_opamp_dummy_magic_21_0.X.n63 two_stage_opamp_dummy_magic_21_0.X.n62 176.733
R6825 two_stage_opamp_dummy_magic_21_0.X.n64 two_stage_opamp_dummy_magic_21_0.X.n63 176.733
R6826 two_stage_opamp_dummy_magic_21_0.X.n65 two_stage_opamp_dummy_magic_21_0.X.n64 176.733
R6827 two_stage_opamp_dummy_magic_21_0.X.n66 two_stage_opamp_dummy_magic_21_0.X.n65 176.733
R6828 two_stage_opamp_dummy_magic_21_0.X.n67 two_stage_opamp_dummy_magic_21_0.X.n66 176.733
R6829 two_stage_opamp_dummy_magic_21_0.X.n68 two_stage_opamp_dummy_magic_21_0.X.n67 176.733
R6830 two_stage_opamp_dummy_magic_21_0.X.n71 two_stage_opamp_dummy_magic_21_0.X.n70 175.05
R6831 two_stage_opamp_dummy_magic_21_0.X.n32 two_stage_opamp_dummy_magic_21_0.X.n31 66.0338
R6832 two_stage_opamp_dummy_magic_21_0.X.n36 two_stage_opamp_dummy_magic_21_0.X.n35 66.0338
R6833 two_stage_opamp_dummy_magic_21_0.X.n38 two_stage_opamp_dummy_magic_21_0.X.n37 66.0338
R6834 two_stage_opamp_dummy_magic_21_0.X.n42 two_stage_opamp_dummy_magic_21_0.X.n41 66.0338
R6835 two_stage_opamp_dummy_magic_21_0.X.n45 two_stage_opamp_dummy_magic_21_0.X.n44 66.0338
R6836 two_stage_opamp_dummy_magic_21_0.X.n49 two_stage_opamp_dummy_magic_21_0.X.n48 66.0338
R6837 two_stage_opamp_dummy_magic_21_0.X.n30 two_stage_opamp_dummy_magic_21_0.X.t18 49.4481
R6838 two_stage_opamp_dummy_magic_21_0.X.n1 two_stage_opamp_dummy_magic_21_0.X.n0 49.3505
R6839 two_stage_opamp_dummy_magic_21_0.X.n5 two_stage_opamp_dummy_magic_21_0.X.n4 49.3505
R6840 two_stage_opamp_dummy_magic_21_0.X.n7 two_stage_opamp_dummy_magic_21_0.X.n6 49.3505
R6841 two_stage_opamp_dummy_magic_21_0.X.n11 two_stage_opamp_dummy_magic_21_0.X.n10 49.3505
R6842 two_stage_opamp_dummy_magic_21_0.X.n13 two_stage_opamp_dummy_magic_21_0.X.n12 49.3505
R6843 two_stage_opamp_dummy_magic_21_0.X.n17 two_stage_opamp_dummy_magic_21_0.X.n16 49.3505
R6844 two_stage_opamp_dummy_magic_21_0.X.n29 two_stage_opamp_dummy_magic_21_0.X.n26 40.1672
R6845 two_stage_opamp_dummy_magic_21_0.X.n29 two_stage_opamp_dummy_magic_21_0.X.n28 40.1672
R6846 two_stage_opamp_dummy_magic_21_0.X.n60 two_stage_opamp_dummy_magic_21_0.X.n52 40.1672
R6847 two_stage_opamp_dummy_magic_21_0.X.n60 two_stage_opamp_dummy_magic_21_0.X.n59 40.1672
R6848 two_stage_opamp_dummy_magic_21_0.X.n69 two_stage_opamp_dummy_magic_21_0.X.n61 40.1672
R6849 two_stage_opamp_dummy_magic_21_0.X.n69 two_stage_opamp_dummy_magic_21_0.X.n68 40.1672
R6850 two_stage_opamp_dummy_magic_21_0.X.n71 two_stage_opamp_dummy_magic_21_0.X.n51 17.688
R6851 two_stage_opamp_dummy_magic_21_0.X.n0 two_stage_opamp_dummy_magic_21_0.X.t22 16.0005
R6852 two_stage_opamp_dummy_magic_21_0.X.n0 two_stage_opamp_dummy_magic_21_0.X.t1 16.0005
R6853 two_stage_opamp_dummy_magic_21_0.X.n4 two_stage_opamp_dummy_magic_21_0.X.t19 16.0005
R6854 two_stage_opamp_dummy_magic_21_0.X.n4 two_stage_opamp_dummy_magic_21_0.X.t16 16.0005
R6855 two_stage_opamp_dummy_magic_21_0.X.n6 two_stage_opamp_dummy_magic_21_0.X.t2 16.0005
R6856 two_stage_opamp_dummy_magic_21_0.X.n6 two_stage_opamp_dummy_magic_21_0.X.t4 16.0005
R6857 two_stage_opamp_dummy_magic_21_0.X.n10 two_stage_opamp_dummy_magic_21_0.X.t24 16.0005
R6858 two_stage_opamp_dummy_magic_21_0.X.n10 two_stage_opamp_dummy_magic_21_0.X.t20 16.0005
R6859 two_stage_opamp_dummy_magic_21_0.X.n12 two_stage_opamp_dummy_magic_21_0.X.t0 16.0005
R6860 two_stage_opamp_dummy_magic_21_0.X.n12 two_stage_opamp_dummy_magic_21_0.X.t21 16.0005
R6861 two_stage_opamp_dummy_magic_21_0.X.n16 two_stage_opamp_dummy_magic_21_0.X.t23 16.0005
R6862 two_stage_opamp_dummy_magic_21_0.X.n16 two_stage_opamp_dummy_magic_21_0.X.t15 16.0005
R6863 two_stage_opamp_dummy_magic_21_0.X.n31 two_stage_opamp_dummy_magic_21_0.X.t17 11.2576
R6864 two_stage_opamp_dummy_magic_21_0.X.n31 two_stage_opamp_dummy_magic_21_0.X.t7 11.2576
R6865 two_stage_opamp_dummy_magic_21_0.X.n35 two_stage_opamp_dummy_magic_21_0.X.t12 11.2576
R6866 two_stage_opamp_dummy_magic_21_0.X.n35 two_stage_opamp_dummy_magic_21_0.X.t3 11.2576
R6867 two_stage_opamp_dummy_magic_21_0.X.n37 two_stage_opamp_dummy_magic_21_0.X.t10 11.2576
R6868 two_stage_opamp_dummy_magic_21_0.X.n37 two_stage_opamp_dummy_magic_21_0.X.t9 11.2576
R6869 two_stage_opamp_dummy_magic_21_0.X.n41 two_stage_opamp_dummy_magic_21_0.X.t14 11.2576
R6870 two_stage_opamp_dummy_magic_21_0.X.n41 two_stage_opamp_dummy_magic_21_0.X.t6 11.2576
R6871 two_stage_opamp_dummy_magic_21_0.X.n44 two_stage_opamp_dummy_magic_21_0.X.t8 11.2576
R6872 two_stage_opamp_dummy_magic_21_0.X.n44 two_stage_opamp_dummy_magic_21_0.X.t11 11.2576
R6873 two_stage_opamp_dummy_magic_21_0.X.n48 two_stage_opamp_dummy_magic_21_0.X.t5 11.2576
R6874 two_stage_opamp_dummy_magic_21_0.X.n48 two_stage_opamp_dummy_magic_21_0.X.t13 11.2576
R6875 two_stage_opamp_dummy_magic_21_0.X.n73 two_stage_opamp_dummy_magic_21_0.X.n72 8.09425
R6876 two_stage_opamp_dummy_magic_21_0.X.n39 two_stage_opamp_dummy_magic_21_0.X.n36 5.91717
R6877 two_stage_opamp_dummy_magic_21_0.X.n36 two_stage_opamp_dummy_magic_21_0.X.n34 5.91717
R6878 two_stage_opamp_dummy_magic_21_0.X.n47 two_stage_opamp_dummy_magic_21_0.X.n32 5.91717
R6879 two_stage_opamp_dummy_magic_21_0.X.n14 two_stage_opamp_dummy_magic_21_0.X.n11 5.6255
R6880 two_stage_opamp_dummy_magic_21_0.X.n8 two_stage_opamp_dummy_magic_21_0.X.n5 5.6255
R6881 two_stage_opamp_dummy_magic_21_0.X.n11 two_stage_opamp_dummy_magic_21_0.X.n3 5.438
R6882 two_stage_opamp_dummy_magic_21_0.X.n5 two_stage_opamp_dummy_magic_21_0.X.n2 5.438
R6883 two_stage_opamp_dummy_magic_21_0.X.n38 two_stage_opamp_dummy_magic_21_0.X.n34 5.29217
R6884 two_stage_opamp_dummy_magic_21_0.X.n39 two_stage_opamp_dummy_magic_21_0.X.n38 5.29217
R6885 two_stage_opamp_dummy_magic_21_0.X.n43 two_stage_opamp_dummy_magic_21_0.X.n42 5.29217
R6886 two_stage_opamp_dummy_magic_21_0.X.n42 two_stage_opamp_dummy_magic_21_0.X.n40 5.29217
R6887 two_stage_opamp_dummy_magic_21_0.X.n46 two_stage_opamp_dummy_magic_21_0.X.n45 5.29217
R6888 two_stage_opamp_dummy_magic_21_0.X.n45 two_stage_opamp_dummy_magic_21_0.X.n33 5.29217
R6889 two_stage_opamp_dummy_magic_21_0.X.n49 two_stage_opamp_dummy_magic_21_0.X.n47 5.29217
R6890 two_stage_opamp_dummy_magic_21_0.X.n50 two_stage_opamp_dummy_magic_21_0.X.n49 5.29217
R6891 two_stage_opamp_dummy_magic_21_0.X.n51 two_stage_opamp_dummy_magic_21_0.X.n50 5.1255
R6892 two_stage_opamp_dummy_magic_21_0.X.n8 two_stage_opamp_dummy_magic_21_0.X.n7 5.063
R6893 two_stage_opamp_dummy_magic_21_0.X.n14 two_stage_opamp_dummy_magic_21_0.X.n13 5.063
R6894 two_stage_opamp_dummy_magic_21_0.X.n17 two_stage_opamp_dummy_magic_21_0.X.n15 5.063
R6895 two_stage_opamp_dummy_magic_21_0.X.n9 two_stage_opamp_dummy_magic_21_0.X.n1 5.063
R6896 two_stage_opamp_dummy_magic_21_0.X.n7 two_stage_opamp_dummy_magic_21_0.X.n2 4.8755
R6897 two_stage_opamp_dummy_magic_21_0.X.n13 two_stage_opamp_dummy_magic_21_0.X.n3 4.8755
R6898 two_stage_opamp_dummy_magic_21_0.X.n18 two_stage_opamp_dummy_magic_21_0.X.n17 4.8755
R6899 two_stage_opamp_dummy_magic_21_0.X.n20 two_stage_opamp_dummy_magic_21_0.X.n19 4.5005
R6900 two_stage_opamp_dummy_magic_21_0.X.n72 two_stage_opamp_dummy_magic_21_0.X.n71 4.5005
R6901 two_stage_opamp_dummy_magic_21_0.X.n72 two_stage_opamp_dummy_magic_21_0.X.n30 3.27133
R6902 two_stage_opamp_dummy_magic_21_0.X.n73 two_stage_opamp_dummy_magic_21_0.X.n20 2.15675
R6903 two_stage_opamp_dummy_magic_21_0.X.n51 two_stage_opamp_dummy_magic_21_0.X.n32 0.792167
R6904 two_stage_opamp_dummy_magic_21_0.X.n50 two_stage_opamp_dummy_magic_21_0.X.n33 0.6255
R6905 two_stage_opamp_dummy_magic_21_0.X.n40 two_stage_opamp_dummy_magic_21_0.X.n33 0.6255
R6906 two_stage_opamp_dummy_magic_21_0.X.n40 two_stage_opamp_dummy_magic_21_0.X.n39 0.6255
R6907 two_stage_opamp_dummy_magic_21_0.X.n43 two_stage_opamp_dummy_magic_21_0.X.n34 0.6255
R6908 two_stage_opamp_dummy_magic_21_0.X.n46 two_stage_opamp_dummy_magic_21_0.X.n43 0.6255
R6909 two_stage_opamp_dummy_magic_21_0.X.n47 two_stage_opamp_dummy_magic_21_0.X.n46 0.6255
R6910 two_stage_opamp_dummy_magic_21_0.X.n15 two_stage_opamp_dummy_magic_21_0.X.n9 0.563
R6911 two_stage_opamp_dummy_magic_21_0.X.n15 two_stage_opamp_dummy_magic_21_0.X.n14 0.563
R6912 two_stage_opamp_dummy_magic_21_0.X.n18 two_stage_opamp_dummy_magic_21_0.X.n3 0.563
R6913 two_stage_opamp_dummy_magic_21_0.X.n19 two_stage_opamp_dummy_magic_21_0.X.n18 0.563
R6914 two_stage_opamp_dummy_magic_21_0.X.n19 two_stage_opamp_dummy_magic_21_0.X.n2 0.563
R6915 two_stage_opamp_dummy_magic_21_0.X.n9 two_stage_opamp_dummy_magic_21_0.X.n8 0.563
R6916 two_stage_opamp_dummy_magic_21_0.X.n20 two_stage_opamp_dummy_magic_21_0.X.n1 0.3755
R6917 two_stage_opamp_dummy_magic_21_0.X two_stage_opamp_dummy_magic_21_0.X.n73 0.063
R6918 two_stage_opamp_dummy_magic_21_0.Vb1.n25 two_stage_opamp_dummy_magic_21_0.Vb1.n24 611.782
R6919 two_stage_opamp_dummy_magic_21_0.Vb1.n9 two_stage_opamp_dummy_magic_21_0.Vb1.t8 449.868
R6920 two_stage_opamp_dummy_magic_21_0.Vb1.n8 two_stage_opamp_dummy_magic_21_0.Vb1.t10 449.868
R6921 two_stage_opamp_dummy_magic_21_0.Vb1.n16 two_stage_opamp_dummy_magic_21_0.Vb1.t27 449.868
R6922 two_stage_opamp_dummy_magic_21_0.Vb1.n4 two_stage_opamp_dummy_magic_21_0.Vb1.n2 339.961
R6923 two_stage_opamp_dummy_magic_21_0.Vb1.n4 two_stage_opamp_dummy_magic_21_0.Vb1.n3 339.272
R6924 two_stage_opamp_dummy_magic_21_0.Vb1.n35 two_stage_opamp_dummy_magic_21_0.Vb1.n34 310.392
R6925 two_stage_opamp_dummy_magic_21_0.Vb1.n9 two_stage_opamp_dummy_magic_21_0.Vb1.t6 273.134
R6926 two_stage_opamp_dummy_magic_21_0.Vb1.n8 two_stage_opamp_dummy_magic_21_0.Vb1.t12 273.134
R6927 two_stage_opamp_dummy_magic_21_0.Vb1.n34 two_stage_opamp_dummy_magic_21_0.Vb1.t24 273.134
R6928 two_stage_opamp_dummy_magic_21_0.Vb1.n25 two_stage_opamp_dummy_magic_21_0.Vb1.t28 273.134
R6929 two_stage_opamp_dummy_magic_21_0.Vb1.n24 two_stage_opamp_dummy_magic_21_0.Vb1.t23 273.134
R6930 two_stage_opamp_dummy_magic_21_0.Vb1.n23 two_stage_opamp_dummy_magic_21_0.Vb1.t32 273.134
R6931 two_stage_opamp_dummy_magic_21_0.Vb1.n22 two_stage_opamp_dummy_magic_21_0.Vb1.t21 273.134
R6932 two_stage_opamp_dummy_magic_21_0.Vb1.n21 two_stage_opamp_dummy_magic_21_0.Vb1.t30 273.134
R6933 two_stage_opamp_dummy_magic_21_0.Vb1.n20 two_stage_opamp_dummy_magic_21_0.Vb1.t26 273.134
R6934 two_stage_opamp_dummy_magic_21_0.Vb1.n19 two_stage_opamp_dummy_magic_21_0.Vb1.t15 273.134
R6935 two_stage_opamp_dummy_magic_21_0.Vb1.n18 two_stage_opamp_dummy_magic_21_0.Vb1.t25 273.134
R6936 two_stage_opamp_dummy_magic_21_0.Vb1.n17 two_stage_opamp_dummy_magic_21_0.Vb1.t14 273.134
R6937 two_stage_opamp_dummy_magic_21_0.Vb1.n16 two_stage_opamp_dummy_magic_21_0.Vb1.t17 273.134
R6938 two_stage_opamp_dummy_magic_21_0.Vb1.n33 two_stage_opamp_dummy_magic_21_0.Vb1.t34 273.134
R6939 two_stage_opamp_dummy_magic_21_0.Vb1.n32 two_stage_opamp_dummy_magic_21_0.Vb1.t22 273.134
R6940 two_stage_opamp_dummy_magic_21_0.Vb1.n31 two_stage_opamp_dummy_magic_21_0.Vb1.t31 273.134
R6941 two_stage_opamp_dummy_magic_21_0.Vb1.n30 two_stage_opamp_dummy_magic_21_0.Vb1.t19 273.134
R6942 two_stage_opamp_dummy_magic_21_0.Vb1.n29 two_stage_opamp_dummy_magic_21_0.Vb1.t16 273.134
R6943 two_stage_opamp_dummy_magic_21_0.Vb1.n28 two_stage_opamp_dummy_magic_21_0.Vb1.t20 273.134
R6944 two_stage_opamp_dummy_magic_21_0.Vb1.n27 two_stage_opamp_dummy_magic_21_0.Vb1.t29 273.134
R6945 two_stage_opamp_dummy_magic_21_0.Vb1.n26 two_stage_opamp_dummy_magic_21_0.Vb1.t18 273.134
R6946 two_stage_opamp_dummy_magic_21_0.Vb1.n17 two_stage_opamp_dummy_magic_21_0.Vb1.n16 176.733
R6947 two_stage_opamp_dummy_magic_21_0.Vb1.n18 two_stage_opamp_dummy_magic_21_0.Vb1.n17 176.733
R6948 two_stage_opamp_dummy_magic_21_0.Vb1.n19 two_stage_opamp_dummy_magic_21_0.Vb1.n18 176.733
R6949 two_stage_opamp_dummy_magic_21_0.Vb1.n20 two_stage_opamp_dummy_magic_21_0.Vb1.n19 176.733
R6950 two_stage_opamp_dummy_magic_21_0.Vb1.n21 two_stage_opamp_dummy_magic_21_0.Vb1.n20 176.733
R6951 two_stage_opamp_dummy_magic_21_0.Vb1.n22 two_stage_opamp_dummy_magic_21_0.Vb1.n21 176.733
R6952 two_stage_opamp_dummy_magic_21_0.Vb1.n23 two_stage_opamp_dummy_magic_21_0.Vb1.n22 176.733
R6953 two_stage_opamp_dummy_magic_21_0.Vb1.n24 two_stage_opamp_dummy_magic_21_0.Vb1.n23 176.733
R6954 two_stage_opamp_dummy_magic_21_0.Vb1.n26 two_stage_opamp_dummy_magic_21_0.Vb1.n25 176.733
R6955 two_stage_opamp_dummy_magic_21_0.Vb1.n27 two_stage_opamp_dummy_magic_21_0.Vb1.n26 176.733
R6956 two_stage_opamp_dummy_magic_21_0.Vb1.n28 two_stage_opamp_dummy_magic_21_0.Vb1.n27 176.733
R6957 two_stage_opamp_dummy_magic_21_0.Vb1.n29 two_stage_opamp_dummy_magic_21_0.Vb1.n28 176.733
R6958 two_stage_opamp_dummy_magic_21_0.Vb1.n30 two_stage_opamp_dummy_magic_21_0.Vb1.n29 176.733
R6959 two_stage_opamp_dummy_magic_21_0.Vb1.n31 two_stage_opamp_dummy_magic_21_0.Vb1.n30 176.733
R6960 two_stage_opamp_dummy_magic_21_0.Vb1.n32 two_stage_opamp_dummy_magic_21_0.Vb1.n31 176.733
R6961 two_stage_opamp_dummy_magic_21_0.Vb1.n33 two_stage_opamp_dummy_magic_21_0.Vb1.n32 176.733
R6962 two_stage_opamp_dummy_magic_21_0.Vb1.n34 two_stage_opamp_dummy_magic_21_0.Vb1.n33 176.733
R6963 two_stage_opamp_dummy_magic_21_0.Vb1.n5 two_stage_opamp_dummy_magic_21_0.Vb1.t33 167.769
R6964 two_stage_opamp_dummy_magic_21_0.Vb1.n1 two_stage_opamp_dummy_magic_21_0.Vb1.n10 161.3
R6965 two_stage_opamp_dummy_magic_21_0.Vb1.n7 two_stage_opamp_dummy_magic_21_0.Vb1.n6 49.3505
R6966 two_stage_opamp_dummy_magic_21_0.Vb1.n1 two_stage_opamp_dummy_magic_21_0.Vb1.n11 49.3505
R6967 two_stage_opamp_dummy_magic_21_0.Vb1.n14 two_stage_opamp_dummy_magic_21_0.Vb1.n13 49.3505
R6968 two_stage_opamp_dummy_magic_21_0.Vb1.n10 two_stage_opamp_dummy_magic_21_0.Vb1.n9 45.5227
R6969 two_stage_opamp_dummy_magic_21_0.Vb1.n10 two_stage_opamp_dummy_magic_21_0.Vb1.n8 45.5227
R6970 two_stage_opamp_dummy_magic_21_0.Vb1.n3 two_stage_opamp_dummy_magic_21_0.Vb1.t1 39.4005
R6971 two_stage_opamp_dummy_magic_21_0.Vb1.n3 two_stage_opamp_dummy_magic_21_0.Vb1.t4 39.4005
R6972 two_stage_opamp_dummy_magic_21_0.Vb1.n2 two_stage_opamp_dummy_magic_21_0.Vb1.t5 39.4005
R6973 two_stage_opamp_dummy_magic_21_0.Vb1.n2 two_stage_opamp_dummy_magic_21_0.Vb1.t0 39.4005
R6974 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_21_0.Vb1.n35 35.5734
R6975 two_stage_opamp_dummy_magic_21_0.Vb1.n35 two_stage_opamp_dummy_magic_21_0.Vb1.n15 17.8547
R6976 two_stage_opamp_dummy_magic_21_0.Vb1.n6 two_stage_opamp_dummy_magic_21_0.Vb1.t2 16.0005
R6977 two_stage_opamp_dummy_magic_21_0.Vb1.n6 two_stage_opamp_dummy_magic_21_0.Vb1.t11 16.0005
R6978 two_stage_opamp_dummy_magic_21_0.Vb1.n11 two_stage_opamp_dummy_magic_21_0.Vb1.t13 16.0005
R6979 two_stage_opamp_dummy_magic_21_0.Vb1.n11 two_stage_opamp_dummy_magic_21_0.Vb1.t7 16.0005
R6980 two_stage_opamp_dummy_magic_21_0.Vb1.n13 two_stage_opamp_dummy_magic_21_0.Vb1.t9 16.0005
R6981 two_stage_opamp_dummy_magic_21_0.Vb1.n13 two_stage_opamp_dummy_magic_21_0.Vb1.t3 16.0005
R6982 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_21_0.Vb1.n4 12.1255
R6983 two_stage_opamp_dummy_magic_21_0.Vb1.n12 two_stage_opamp_dummy_magic_21_0.Vb1.n7 5.6255
R6984 two_stage_opamp_dummy_magic_21_0.Vb1.n14 two_stage_opamp_dummy_magic_21_0.Vb1.n12 5.6255
R6985 two_stage_opamp_dummy_magic_21_0.Vb1.n12 two_stage_opamp_dummy_magic_21_0.Vb1.n1 5.063
R6986 two_stage_opamp_dummy_magic_21_0.Vb1.n15 two_stage_opamp_dummy_magic_21_0.Vb1.n14 4.938
R6987 two_stage_opamp_dummy_magic_21_0.Vb1.n7 two_stage_opamp_dummy_magic_21_0.Vb1.n5 4.938
R6988 two_stage_opamp_dummy_magic_21_0.Vb1.n1 two_stage_opamp_dummy_magic_21_0.Vb1.n0 4.938
R6989 two_stage_opamp_dummy_magic_21_0.Vb1.n15 two_stage_opamp_dummy_magic_21_0.Vb1.n0 0.563
R6990 two_stage_opamp_dummy_magic_21_0.Vb1.n5 two_stage_opamp_dummy_magic_21_0.Vb1.n0 0.563
R6991 two_stage_opamp_dummy_magic_21_0.VD1.n23 two_stage_opamp_dummy_magic_21_0.VD1.n22 49.3505
R6992 two_stage_opamp_dummy_magic_21_0.VD1.n26 two_stage_opamp_dummy_magic_21_0.VD1.n25 49.3505
R6993 two_stage_opamp_dummy_magic_21_0.VD1.n29 two_stage_opamp_dummy_magic_21_0.VD1.n28 49.3505
R6994 two_stage_opamp_dummy_magic_21_0.VD1.n32 two_stage_opamp_dummy_magic_21_0.VD1.n31 49.3505
R6995 two_stage_opamp_dummy_magic_21_0.VD1.n4 two_stage_opamp_dummy_magic_21_0.VD1.n3 49.3505
R6996 two_stage_opamp_dummy_magic_21_0.VD1.n7 two_stage_opamp_dummy_magic_21_0.VD1.n6 49.3505
R6997 two_stage_opamp_dummy_magic_21_0.VD1.n10 two_stage_opamp_dummy_magic_21_0.VD1.n9 49.3505
R6998 two_stage_opamp_dummy_magic_21_0.VD1.n13 two_stage_opamp_dummy_magic_21_0.VD1.n12 49.3505
R6999 two_stage_opamp_dummy_magic_21_0.VD1.n15 two_stage_opamp_dummy_magic_21_0.VD1.n14 49.3505
R7000 two_stage_opamp_dummy_magic_21_0.VD1.n19 two_stage_opamp_dummy_magic_21_0.VD1.n18 49.3505
R7001 two_stage_opamp_dummy_magic_21_0.VD1.n37 two_stage_opamp_dummy_magic_21_0.VD1.n36 49.3505
R7002 two_stage_opamp_dummy_magic_21_0.VD1.n22 two_stage_opamp_dummy_magic_21_0.VD1.t14 16.0005
R7003 two_stage_opamp_dummy_magic_21_0.VD1.n22 two_stage_opamp_dummy_magic_21_0.VD1.t19 16.0005
R7004 two_stage_opamp_dummy_magic_21_0.VD1.n25 two_stage_opamp_dummy_magic_21_0.VD1.t21 16.0005
R7005 two_stage_opamp_dummy_magic_21_0.VD1.n25 two_stage_opamp_dummy_magic_21_0.VD1.t16 16.0005
R7006 two_stage_opamp_dummy_magic_21_0.VD1.n28 two_stage_opamp_dummy_magic_21_0.VD1.t12 16.0005
R7007 two_stage_opamp_dummy_magic_21_0.VD1.n28 two_stage_opamp_dummy_magic_21_0.VD1.t17 16.0005
R7008 two_stage_opamp_dummy_magic_21_0.VD1.n31 two_stage_opamp_dummy_magic_21_0.VD1.t13 16.0005
R7009 two_stage_opamp_dummy_magic_21_0.VD1.n31 two_stage_opamp_dummy_magic_21_0.VD1.t18 16.0005
R7010 two_stage_opamp_dummy_magic_21_0.VD1.n3 two_stage_opamp_dummy_magic_21_0.VD1.t9 16.0005
R7011 two_stage_opamp_dummy_magic_21_0.VD1.n3 two_stage_opamp_dummy_magic_21_0.VD1.t7 16.0005
R7012 two_stage_opamp_dummy_magic_21_0.VD1.n6 two_stage_opamp_dummy_magic_21_0.VD1.t11 16.0005
R7013 two_stage_opamp_dummy_magic_21_0.VD1.n6 two_stage_opamp_dummy_magic_21_0.VD1.t5 16.0005
R7014 two_stage_opamp_dummy_magic_21_0.VD1.n9 two_stage_opamp_dummy_magic_21_0.VD1.t0 16.0005
R7015 two_stage_opamp_dummy_magic_21_0.VD1.n9 two_stage_opamp_dummy_magic_21_0.VD1.t2 16.0005
R7016 two_stage_opamp_dummy_magic_21_0.VD1.n12 two_stage_opamp_dummy_magic_21_0.VD1.t10 16.0005
R7017 two_stage_opamp_dummy_magic_21_0.VD1.n12 two_stage_opamp_dummy_magic_21_0.VD1.t8 16.0005
R7018 two_stage_opamp_dummy_magic_21_0.VD1.n14 two_stage_opamp_dummy_magic_21_0.VD1.t1 16.0005
R7019 two_stage_opamp_dummy_magic_21_0.VD1.n14 two_stage_opamp_dummy_magic_21_0.VD1.t6 16.0005
R7020 two_stage_opamp_dummy_magic_21_0.VD1.n18 two_stage_opamp_dummy_magic_21_0.VD1.t4 16.0005
R7021 two_stage_opamp_dummy_magic_21_0.VD1.n18 two_stage_opamp_dummy_magic_21_0.VD1.t3 16.0005
R7022 two_stage_opamp_dummy_magic_21_0.VD1.t20 two_stage_opamp_dummy_magic_21_0.VD1.n37 16.0005
R7023 two_stage_opamp_dummy_magic_21_0.VD1.n37 two_stage_opamp_dummy_magic_21_0.VD1.t15 16.0005
R7024 two_stage_opamp_dummy_magic_21_0.VD1.n35 two_stage_opamp_dummy_magic_21_0.VD1.n21 5.77133
R7025 two_stage_opamp_dummy_magic_21_0.VD1.n13 two_stage_opamp_dummy_magic_21_0.VD1.n2 5.64633
R7026 two_stage_opamp_dummy_magic_21_0.VD1.n5 two_stage_opamp_dummy_magic_21_0.VD1.n4 5.64633
R7027 two_stage_opamp_dummy_magic_21_0.VD1.n30 two_stage_opamp_dummy_magic_21_0.VD1.n29 5.6255
R7028 two_stage_opamp_dummy_magic_21_0.VD1.n24 two_stage_opamp_dummy_magic_21_0.VD1.n23 5.6255
R7029 two_stage_opamp_dummy_magic_21_0.VD1.n33 two_stage_opamp_dummy_magic_21_0.VD1.n29 5.438
R7030 two_stage_opamp_dummy_magic_21_0.VD1.n27 two_stage_opamp_dummy_magic_21_0.VD1.n23 5.438
R7031 two_stage_opamp_dummy_magic_21_0.VD1.n16 two_stage_opamp_dummy_magic_21_0.VD1.n13 5.438
R7032 two_stage_opamp_dummy_magic_21_0.VD1.n8 two_stage_opamp_dummy_magic_21_0.VD1.n4 5.438
R7033 two_stage_opamp_dummy_magic_21_0.VD1.n7 two_stage_opamp_dummy_magic_21_0.VD1.n5 5.08383
R7034 two_stage_opamp_dummy_magic_21_0.VD1.n10 two_stage_opamp_dummy_magic_21_0.VD1.n1 5.08383
R7035 two_stage_opamp_dummy_magic_21_0.VD1.n15 two_stage_opamp_dummy_magic_21_0.VD1.n2 5.08383
R7036 two_stage_opamp_dummy_magic_21_0.VD1.n20 two_stage_opamp_dummy_magic_21_0.VD1.n19 5.08383
R7037 two_stage_opamp_dummy_magic_21_0.VD1.n26 two_stage_opamp_dummy_magic_21_0.VD1.n24 5.063
R7038 two_stage_opamp_dummy_magic_21_0.VD1.n36 two_stage_opamp_dummy_magic_21_0.VD1.n0 5.063
R7039 two_stage_opamp_dummy_magic_21_0.VD1.n32 two_stage_opamp_dummy_magic_21_0.VD1.n30 5.063
R7040 two_stage_opamp_dummy_magic_21_0.VD1.n27 two_stage_opamp_dummy_magic_21_0.VD1.n26 4.8755
R7041 two_stage_opamp_dummy_magic_21_0.VD1.n33 two_stage_opamp_dummy_magic_21_0.VD1.n32 4.8755
R7042 two_stage_opamp_dummy_magic_21_0.VD1.n8 two_stage_opamp_dummy_magic_21_0.VD1.n7 4.8755
R7043 two_stage_opamp_dummy_magic_21_0.VD1.n11 two_stage_opamp_dummy_magic_21_0.VD1.n10 4.8755
R7044 two_stage_opamp_dummy_magic_21_0.VD1.n16 two_stage_opamp_dummy_magic_21_0.VD1.n15 4.8755
R7045 two_stage_opamp_dummy_magic_21_0.VD1.n19 two_stage_opamp_dummy_magic_21_0.VD1.n17 4.8755
R7046 two_stage_opamp_dummy_magic_21_0.VD1.n35 two_stage_opamp_dummy_magic_21_0.VD1.n34 4.5005
R7047 two_stage_opamp_dummy_magic_21_0.VD1.n34 two_stage_opamp_dummy_magic_21_0.VD1.n33 0.563
R7048 two_stage_opamp_dummy_magic_21_0.VD1.n30 two_stage_opamp_dummy_magic_21_0.VD1.n0 0.563
R7049 two_stage_opamp_dummy_magic_21_0.VD1.n24 two_stage_opamp_dummy_magic_21_0.VD1.n0 0.563
R7050 two_stage_opamp_dummy_magic_21_0.VD1.n34 two_stage_opamp_dummy_magic_21_0.VD1.n27 0.563
R7051 two_stage_opamp_dummy_magic_21_0.VD1.n20 two_stage_opamp_dummy_magic_21_0.VD1.n2 0.563
R7052 two_stage_opamp_dummy_magic_21_0.VD1.n17 two_stage_opamp_dummy_magic_21_0.VD1.n16 0.563
R7053 two_stage_opamp_dummy_magic_21_0.VD1.n17 two_stage_opamp_dummy_magic_21_0.VD1.n11 0.563
R7054 two_stage_opamp_dummy_magic_21_0.VD1.n11 two_stage_opamp_dummy_magic_21_0.VD1.n8 0.563
R7055 two_stage_opamp_dummy_magic_21_0.VD1.n5 two_stage_opamp_dummy_magic_21_0.VD1.n1 0.563
R7056 two_stage_opamp_dummy_magic_21_0.VD1.n36 two_stage_opamp_dummy_magic_21_0.VD1.n35 0.3755
R7057 two_stage_opamp_dummy_magic_21_0.VD1.n21 two_stage_opamp_dummy_magic_21_0.VD1.n20 0.234875
R7058 two_stage_opamp_dummy_magic_21_0.VD1.n21 two_stage_opamp_dummy_magic_21_0.VD1.n1 0.234875
R7059 a_6930_22564.t0 a_6930_22564.t1 178.133
R7060 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t13 369.534
R7061 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t12 369.534
R7062 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t29 369.534
R7063 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t17 369.534
R7064 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R7065 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t20 369.534
R7066 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7067 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7068 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7069 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7070 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t14 238.322
R7071 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t27 238.322
R7072 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t26 192.8
R7073 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t19 192.8
R7074 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t16 192.8
R7075 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t23 192.8
R7076 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t22 192.8
R7077 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t24 192.8
R7078 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t10 192.8
R7079 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t18 192.8
R7080 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t25 192.8
R7081 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t11 192.8
R7082 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t15 192.8
R7083 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t28 192.8
R7084 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7085 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7086 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7087 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7088 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7089 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7090 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7091 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7092 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n14 167.519
R7093 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7094 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t0 137.48
R7095 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t1 100.635
R7096 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7097 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7098 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7099 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7100 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7101 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7102 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t3 39.4005
R7103 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t5 39.4005
R7104 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t7 39.4005
R7105 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t9 39.4005
R7106 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t6 39.4005
R7107 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t8 39.4005
R7108 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t4 39.4005
R7109 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t2 39.4005
R7110 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 27.5005
R7111 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n13 9.53175
R7112 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7113 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 2.34425
R7114 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7115 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7116 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 1.688
R7117 two_stage_opamp_dummy_magic_21_0.cap_res_X.t138 two_stage_opamp_dummy_magic_21_0.cap_res_X.t5 50.1603
R7118 two_stage_opamp_dummy_magic_21_0.cap_res_X.t22 two_stage_opamp_dummy_magic_21_0.cap_res_X.t61 0.1603
R7119 two_stage_opamp_dummy_magic_21_0.cap_res_X.t45 two_stage_opamp_dummy_magic_21_0.cap_res_X.t86 0.1603
R7120 two_stage_opamp_dummy_magic_21_0.cap_res_X.t9 two_stage_opamp_dummy_magic_21_0.cap_res_X.t46 0.1603
R7121 two_stage_opamp_dummy_magic_21_0.cap_res_X.t111 two_stage_opamp_dummy_magic_21_0.cap_res_X.t11 0.1603
R7122 two_stage_opamp_dummy_magic_21_0.cap_res_X.t76 two_stage_opamp_dummy_magic_21_0.cap_res_X.t91 0.1603
R7123 two_stage_opamp_dummy_magic_21_0.cap_res_X.t113 two_stage_opamp_dummy_magic_21_0.cap_res_X.t76 0.1603
R7124 two_stage_opamp_dummy_magic_21_0.cap_res_X.t71 two_stage_opamp_dummy_magic_21_0.cap_res_X.t113 0.1603
R7125 two_stage_opamp_dummy_magic_21_0.cap_res_X.t100 two_stage_opamp_dummy_magic_21_0.cap_res_X.t38 0.1603
R7126 two_stage_opamp_dummy_magic_21_0.cap_res_X.t135 two_stage_opamp_dummy_magic_21_0.cap_res_X.t100 0.1603
R7127 two_stage_opamp_dummy_magic_21_0.cap_res_X.t95 two_stage_opamp_dummy_magic_21_0.cap_res_X.t135 0.1603
R7128 two_stage_opamp_dummy_magic_21_0.cap_res_X.t126 two_stage_opamp_dummy_magic_21_0.cap_res_X.t89 0.1603
R7129 two_stage_opamp_dummy_magic_21_0.cap_res_X.t87 two_stage_opamp_dummy_magic_21_0.cap_res_X.t48 0.1603
R7130 two_stage_opamp_dummy_magic_21_0.cap_res_X.t41 two_stage_opamp_dummy_magic_21_0.cap_res_X.t80 0.1603
R7131 two_stage_opamp_dummy_magic_21_0.cap_res_X.t26 two_stage_opamp_dummy_magic_21_0.cap_res_X.t129 0.1603
R7132 two_stage_opamp_dummy_magic_21_0.cap_res_X.t8 two_stage_opamp_dummy_magic_21_0.cap_res_X.t44 0.1603
R7133 two_stage_opamp_dummy_magic_21_0.cap_res_X.t133 two_stage_opamp_dummy_magic_21_0.cap_res_X.t94 0.1603
R7134 two_stage_opamp_dummy_magic_21_0.cap_res_X.t24 two_stage_opamp_dummy_magic_21_0.cap_res_X.t57 0.1603
R7135 two_stage_opamp_dummy_magic_21_0.cap_res_X.t78 two_stage_opamp_dummy_magic_21_0.cap_res_X.t42 0.1603
R7136 two_stage_opamp_dummy_magic_21_0.cap_res_X.t64 two_stage_opamp_dummy_magic_21_0.cap_res_X.t101 0.1603
R7137 two_stage_opamp_dummy_magic_21_0.cap_res_X.t117 two_stage_opamp_dummy_magic_21_0.cap_res_X.t82 0.1603
R7138 two_stage_opamp_dummy_magic_21_0.cap_res_X.t30 two_stage_opamp_dummy_magic_21_0.cap_res_X.t65 0.1603
R7139 two_stage_opamp_dummy_magic_21_0.cap_res_X.t85 two_stage_opamp_dummy_magic_21_0.cap_res_X.t47 0.1603
R7140 two_stage_opamp_dummy_magic_21_0.cap_res_X.t68 two_stage_opamp_dummy_magic_21_0.cap_res_X.t104 0.1603
R7141 two_stage_opamp_dummy_magic_21_0.cap_res_X.t123 two_stage_opamp_dummy_magic_21_0.cap_res_X.t88 0.1603
R7142 two_stage_opamp_dummy_magic_21_0.cap_res_X.t108 two_stage_opamp_dummy_magic_21_0.cap_res_X.t3 0.1603
R7143 two_stage_opamp_dummy_magic_21_0.cap_res_X.t21 two_stage_opamp_dummy_magic_21_0.cap_res_X.t127 0.1603
R7144 two_stage_opamp_dummy_magic_21_0.cap_res_X.t75 two_stage_opamp_dummy_magic_21_0.cap_res_X.t110 0.1603
R7145 two_stage_opamp_dummy_magic_21_0.cap_res_X.t128 two_stage_opamp_dummy_magic_21_0.cap_res_X.t93 0.1603
R7146 two_stage_opamp_dummy_magic_21_0.cap_res_X.t116 two_stage_opamp_dummy_magic_21_0.cap_res_X.t10 0.1603
R7147 two_stage_opamp_dummy_magic_21_0.cap_res_X.t27 two_stage_opamp_dummy_magic_21_0.cap_res_X.t134 0.1603
R7148 two_stage_opamp_dummy_magic_21_0.cap_res_X.t15 two_stage_opamp_dummy_magic_21_0.cap_res_X.t49 0.1603
R7149 two_stage_opamp_dummy_magic_21_0.cap_res_X.t67 two_stage_opamp_dummy_magic_21_0.cap_res_X.t33 0.1603
R7150 two_stage_opamp_dummy_magic_21_0.cap_res_X.t53 two_stage_opamp_dummy_magic_21_0.cap_res_X.t90 0.1603
R7151 two_stage_opamp_dummy_magic_21_0.cap_res_X.t107 two_stage_opamp_dummy_magic_21_0.cap_res_X.t72 0.1603
R7152 two_stage_opamp_dummy_magic_21_0.cap_res_X.t19 two_stage_opamp_dummy_magic_21_0.cap_res_X.t52 0.1603
R7153 two_stage_opamp_dummy_magic_21_0.cap_res_X.t73 two_stage_opamp_dummy_magic_21_0.cap_res_X.t35 0.1603
R7154 two_stage_opamp_dummy_magic_21_0.cap_res_X.t56 two_stage_opamp_dummy_magic_21_0.cap_res_X.t96 0.1603
R7155 two_stage_opamp_dummy_magic_21_0.cap_res_X.t115 two_stage_opamp_dummy_magic_21_0.cap_res_X.t77 0.1603
R7156 two_stage_opamp_dummy_magic_21_0.cap_res_X.t99 two_stage_opamp_dummy_magic_21_0.cap_res_X.t136 0.1603
R7157 two_stage_opamp_dummy_magic_21_0.cap_res_X.t14 two_stage_opamp_dummy_magic_21_0.cap_res_X.t119 0.1603
R7158 two_stage_opamp_dummy_magic_21_0.cap_res_X.t7 two_stage_opamp_dummy_magic_21_0.cap_res_X.t83 0.1603
R7159 two_stage_opamp_dummy_magic_21_0.cap_res_X.t98 two_stage_opamp_dummy_magic_21_0.cap_res_X.t40 0.1603
R7160 two_stage_opamp_dummy_magic_21_0.cap_res_X.t59 two_stage_opamp_dummy_magic_21_0.cap_res_X.t92 0.1603
R7161 two_stage_opamp_dummy_magic_21_0.cap_res_X.t25 two_stage_opamp_dummy_magic_21_0.cap_res_X.t2 0.1603
R7162 two_stage_opamp_dummy_magic_21_0.cap_res_X.t132 two_stage_opamp_dummy_magic_21_0.cap_res_X.t50 0.1603
R7163 two_stage_opamp_dummy_magic_21_0.cap_res_X.t81 two_stage_opamp_dummy_magic_21_0.cap_res_X.t13 0.1603
R7164 two_stage_opamp_dummy_magic_21_0.cap_res_X.t43 two_stage_opamp_dummy_magic_21_0.cap_res_X.t60 0.1603
R7165 two_stage_opamp_dummy_magic_21_0.cap_res_X.t12 two_stage_opamp_dummy_magic_21_0.cap_res_X.t114 0.1603
R7166 two_stage_opamp_dummy_magic_21_0.cap_res_X.t102 two_stage_opamp_dummy_magic_21_0.cap_res_X.t70 0.1603
R7167 two_stage_opamp_dummy_magic_21_0.cap_res_X.t62 two_stage_opamp_dummy_magic_21_0.cap_res_X.t122 0.1603
R7168 two_stage_opamp_dummy_magic_21_0.cap_res_X.t118 two_stage_opamp_dummy_magic_21_0.cap_res_X.t84 0.1603
R7169 two_stage_opamp_dummy_magic_21_0.cap_res_X.t131 two_stage_opamp_dummy_magic_21_0.cap_res_X.t39 0.1603
R7170 two_stage_opamp_dummy_magic_21_0.cap_res_X.t20 two_stage_opamp_dummy_magic_21_0.cap_res_X.t112 0.1603
R7171 two_stage_opamp_dummy_magic_21_0.cap_res_X.t55 two_stage_opamp_dummy_magic_21_0.cap_res_X.t20 0.1603
R7172 two_stage_opamp_dummy_magic_21_0.cap_res_X.t17 two_stage_opamp_dummy_magic_21_0.cap_res_X.t55 0.1603
R7173 two_stage_opamp_dummy_magic_21_0.cap_res_X.t97 two_stage_opamp_dummy_magic_21_0.cap_res_X.t54 0.1603
R7174 two_stage_opamp_dummy_magic_21_0.cap_res_X.t58 two_stage_opamp_dummy_magic_21_0.cap_res_X.t97 0.1603
R7175 two_stage_opamp_dummy_magic_21_0.cap_res_X.t5 two_stage_opamp_dummy_magic_21_0.cap_res_X.t58 0.1603
R7176 two_stage_opamp_dummy_magic_21_0.cap_res_X.n29 two_stage_opamp_dummy_magic_21_0.cap_res_X.t124 0.159278
R7177 two_stage_opamp_dummy_magic_21_0.cap_res_X.n30 two_stage_opamp_dummy_magic_21_0.cap_res_X.t6 0.159278
R7178 two_stage_opamp_dummy_magic_21_0.cap_res_X.n31 two_stage_opamp_dummy_magic_21_0.cap_res_X.t106 0.159278
R7179 two_stage_opamp_dummy_magic_21_0.cap_res_X.n32 two_stage_opamp_dummy_magic_21_0.cap_res_X.t69 0.159278
R7180 two_stage_opamp_dummy_magic_21_0.cap_res_X.n33 two_stage_opamp_dummy_magic_21_0.cap_res_X.t31 0.159278
R7181 two_stage_opamp_dummy_magic_21_0.cap_res_X.n34 two_stage_opamp_dummy_magic_21_0.cap_res_X.t51 0.159278
R7182 two_stage_opamp_dummy_magic_21_0.cap_res_X.n25 two_stage_opamp_dummy_magic_21_0.cap_res_X.t66 0.159278
R7183 two_stage_opamp_dummy_magic_21_0.cap_res_X.t29 two_stage_opamp_dummy_magic_21_0.cap_res_X.n9 0.159278
R7184 two_stage_opamp_dummy_magic_21_0.cap_res_X.t63 two_stage_opamp_dummy_magic_21_0.cap_res_X.n10 0.159278
R7185 two_stage_opamp_dummy_magic_21_0.cap_res_X.t23 two_stage_opamp_dummy_magic_21_0.cap_res_X.n11 0.159278
R7186 two_stage_opamp_dummy_magic_21_0.cap_res_X.t125 two_stage_opamp_dummy_magic_21_0.cap_res_X.n12 0.159278
R7187 two_stage_opamp_dummy_magic_21_0.cap_res_X.t18 two_stage_opamp_dummy_magic_21_0.cap_res_X.n13 0.159278
R7188 two_stage_opamp_dummy_magic_21_0.cap_res_X.t121 two_stage_opamp_dummy_magic_21_0.cap_res_X.n14 0.159278
R7189 two_stage_opamp_dummy_magic_21_0.cap_res_X.t79 two_stage_opamp_dummy_magic_21_0.cap_res_X.n15 0.159278
R7190 two_stage_opamp_dummy_magic_21_0.cap_res_X.t36 two_stage_opamp_dummy_magic_21_0.cap_res_X.n16 0.159278
R7191 two_stage_opamp_dummy_magic_21_0.cap_res_X.t74 two_stage_opamp_dummy_magic_21_0.cap_res_X.n17 0.159278
R7192 two_stage_opamp_dummy_magic_21_0.cap_res_X.t34 two_stage_opamp_dummy_magic_21_0.cap_res_X.n18 0.159278
R7193 two_stage_opamp_dummy_magic_21_0.cap_res_X.t137 two_stage_opamp_dummy_magic_21_0.cap_res_X.n19 0.159278
R7194 two_stage_opamp_dummy_magic_21_0.cap_res_X.t28 two_stage_opamp_dummy_magic_21_0.cap_res_X.n20 0.159278
R7195 two_stage_opamp_dummy_magic_21_0.cap_res_X.t130 two_stage_opamp_dummy_magic_21_0.cap_res_X.n21 0.159278
R7196 two_stage_opamp_dummy_magic_21_0.cap_res_X.t109 two_stage_opamp_dummy_magic_21_0.cap_res_X.n22 0.159278
R7197 two_stage_opamp_dummy_magic_21_0.cap_res_X.t4 two_stage_opamp_dummy_magic_21_0.cap_res_X.n23 0.159278
R7198 two_stage_opamp_dummy_magic_21_0.cap_res_X.t105 two_stage_opamp_dummy_magic_21_0.cap_res_X.n24 0.159278
R7199 two_stage_opamp_dummy_magic_21_0.cap_res_X.n26 two_stage_opamp_dummy_magic_21_0.cap_res_X.t103 0.159278
R7200 two_stage_opamp_dummy_magic_21_0.cap_res_X.n27 two_stage_opamp_dummy_magic_21_0.cap_res_X.t0 0.159278
R7201 two_stage_opamp_dummy_magic_21_0.cap_res_X.n28 two_stage_opamp_dummy_magic_21_0.cap_res_X.t120 0.159278
R7202 two_stage_opamp_dummy_magic_21_0.cap_res_X.n35 two_stage_opamp_dummy_magic_21_0.cap_res_X.t16 0.159278
R7203 two_stage_opamp_dummy_magic_21_0.cap_res_X.t66 two_stage_opamp_dummy_magic_21_0.cap_res_X.t87 0.137822
R7204 two_stage_opamp_dummy_magic_21_0.cap_res_X.n25 two_stage_opamp_dummy_magic_21_0.cap_res_X.t126 0.1368
R7205 two_stage_opamp_dummy_magic_21_0.cap_res_X.n24 two_stage_opamp_dummy_magic_21_0.cap_res_X.t41 0.1368
R7206 two_stage_opamp_dummy_magic_21_0.cap_res_X.n24 two_stage_opamp_dummy_magic_21_0.cap_res_X.t26 0.1368
R7207 two_stage_opamp_dummy_magic_21_0.cap_res_X.n23 two_stage_opamp_dummy_magic_21_0.cap_res_X.t8 0.1368
R7208 two_stage_opamp_dummy_magic_21_0.cap_res_X.n23 two_stage_opamp_dummy_magic_21_0.cap_res_X.t133 0.1368
R7209 two_stage_opamp_dummy_magic_21_0.cap_res_X.n22 two_stage_opamp_dummy_magic_21_0.cap_res_X.t24 0.1368
R7210 two_stage_opamp_dummy_magic_21_0.cap_res_X.n22 two_stage_opamp_dummy_magic_21_0.cap_res_X.t78 0.1368
R7211 two_stage_opamp_dummy_magic_21_0.cap_res_X.n21 two_stage_opamp_dummy_magic_21_0.cap_res_X.t64 0.1368
R7212 two_stage_opamp_dummy_magic_21_0.cap_res_X.n21 two_stage_opamp_dummy_magic_21_0.cap_res_X.t117 0.1368
R7213 two_stage_opamp_dummy_magic_21_0.cap_res_X.n20 two_stage_opamp_dummy_magic_21_0.cap_res_X.t30 0.1368
R7214 two_stage_opamp_dummy_magic_21_0.cap_res_X.n20 two_stage_opamp_dummy_magic_21_0.cap_res_X.t85 0.1368
R7215 two_stage_opamp_dummy_magic_21_0.cap_res_X.n19 two_stage_opamp_dummy_magic_21_0.cap_res_X.t68 0.1368
R7216 two_stage_opamp_dummy_magic_21_0.cap_res_X.n19 two_stage_opamp_dummy_magic_21_0.cap_res_X.t123 0.1368
R7217 two_stage_opamp_dummy_magic_21_0.cap_res_X.n18 two_stage_opamp_dummy_magic_21_0.cap_res_X.t108 0.1368
R7218 two_stage_opamp_dummy_magic_21_0.cap_res_X.n18 two_stage_opamp_dummy_magic_21_0.cap_res_X.t21 0.1368
R7219 two_stage_opamp_dummy_magic_21_0.cap_res_X.n17 two_stage_opamp_dummy_magic_21_0.cap_res_X.t75 0.1368
R7220 two_stage_opamp_dummy_magic_21_0.cap_res_X.n17 two_stage_opamp_dummy_magic_21_0.cap_res_X.t128 0.1368
R7221 two_stage_opamp_dummy_magic_21_0.cap_res_X.n16 two_stage_opamp_dummy_magic_21_0.cap_res_X.t116 0.1368
R7222 two_stage_opamp_dummy_magic_21_0.cap_res_X.n16 two_stage_opamp_dummy_magic_21_0.cap_res_X.t27 0.1368
R7223 two_stage_opamp_dummy_magic_21_0.cap_res_X.n15 two_stage_opamp_dummy_magic_21_0.cap_res_X.t15 0.1368
R7224 two_stage_opamp_dummy_magic_21_0.cap_res_X.n15 two_stage_opamp_dummy_magic_21_0.cap_res_X.t67 0.1368
R7225 two_stage_opamp_dummy_magic_21_0.cap_res_X.n14 two_stage_opamp_dummy_magic_21_0.cap_res_X.t53 0.1368
R7226 two_stage_opamp_dummy_magic_21_0.cap_res_X.n14 two_stage_opamp_dummy_magic_21_0.cap_res_X.t107 0.1368
R7227 two_stage_opamp_dummy_magic_21_0.cap_res_X.n13 two_stage_opamp_dummy_magic_21_0.cap_res_X.t19 0.1368
R7228 two_stage_opamp_dummy_magic_21_0.cap_res_X.n13 two_stage_opamp_dummy_magic_21_0.cap_res_X.t73 0.1368
R7229 two_stage_opamp_dummy_magic_21_0.cap_res_X.n12 two_stage_opamp_dummy_magic_21_0.cap_res_X.t56 0.1368
R7230 two_stage_opamp_dummy_magic_21_0.cap_res_X.n12 two_stage_opamp_dummy_magic_21_0.cap_res_X.t115 0.1368
R7231 two_stage_opamp_dummy_magic_21_0.cap_res_X.n11 two_stage_opamp_dummy_magic_21_0.cap_res_X.t99 0.1368
R7232 two_stage_opamp_dummy_magic_21_0.cap_res_X.n11 two_stage_opamp_dummy_magic_21_0.cap_res_X.t14 0.1368
R7233 two_stage_opamp_dummy_magic_21_0.cap_res_X.n10 two_stage_opamp_dummy_magic_21_0.cap_res_X.t118 0.1368
R7234 two_stage_opamp_dummy_magic_21_0.cap_res_X.n9 two_stage_opamp_dummy_magic_21_0.cap_res_X.t131 0.1368
R7235 two_stage_opamp_dummy_magic_21_0.cap_res_X.n0 two_stage_opamp_dummy_magic_21_0.cap_res_X.t7 0.114322
R7236 two_stage_opamp_dummy_magic_21_0.cap_res_X.n30 two_stage_opamp_dummy_magic_21_0.cap_res_X.n29 0.1133
R7237 two_stage_opamp_dummy_magic_21_0.cap_res_X.n31 two_stage_opamp_dummy_magic_21_0.cap_res_X.n30 0.1133
R7238 two_stage_opamp_dummy_magic_21_0.cap_res_X.n32 two_stage_opamp_dummy_magic_21_0.cap_res_X.n31 0.1133
R7239 two_stage_opamp_dummy_magic_21_0.cap_res_X.n33 two_stage_opamp_dummy_magic_21_0.cap_res_X.n32 0.1133
R7240 two_stage_opamp_dummy_magic_21_0.cap_res_X.n34 two_stage_opamp_dummy_magic_21_0.cap_res_X.n33 0.1133
R7241 two_stage_opamp_dummy_magic_21_0.cap_res_X.n1 two_stage_opamp_dummy_magic_21_0.cap_res_X.n0 0.1133
R7242 two_stage_opamp_dummy_magic_21_0.cap_res_X.n2 two_stage_opamp_dummy_magic_21_0.cap_res_X.n1 0.1133
R7243 two_stage_opamp_dummy_magic_21_0.cap_res_X.n3 two_stage_opamp_dummy_magic_21_0.cap_res_X.n2 0.1133
R7244 two_stage_opamp_dummy_magic_21_0.cap_res_X.n4 two_stage_opamp_dummy_magic_21_0.cap_res_X.n3 0.1133
R7245 two_stage_opamp_dummy_magic_21_0.cap_res_X.n5 two_stage_opamp_dummy_magic_21_0.cap_res_X.n4 0.1133
R7246 two_stage_opamp_dummy_magic_21_0.cap_res_X.n6 two_stage_opamp_dummy_magic_21_0.cap_res_X.n5 0.1133
R7247 two_stage_opamp_dummy_magic_21_0.cap_res_X.n7 two_stage_opamp_dummy_magic_21_0.cap_res_X.n6 0.1133
R7248 two_stage_opamp_dummy_magic_21_0.cap_res_X.n8 two_stage_opamp_dummy_magic_21_0.cap_res_X.n7 0.1133
R7249 two_stage_opamp_dummy_magic_21_0.cap_res_X.n10 two_stage_opamp_dummy_magic_21_0.cap_res_X.n8 0.1133
R7250 two_stage_opamp_dummy_magic_21_0.cap_res_X.n26 two_stage_opamp_dummy_magic_21_0.cap_res_X.n25 0.1133
R7251 two_stage_opamp_dummy_magic_21_0.cap_res_X.n27 two_stage_opamp_dummy_magic_21_0.cap_res_X.n26 0.1133
R7252 two_stage_opamp_dummy_magic_21_0.cap_res_X.n28 two_stage_opamp_dummy_magic_21_0.cap_res_X.n27 0.1133
R7253 two_stage_opamp_dummy_magic_21_0.cap_res_X.n35 two_stage_opamp_dummy_magic_21_0.cap_res_X.n28 0.1133
R7254 two_stage_opamp_dummy_magic_21_0.cap_res_X.n35 two_stage_opamp_dummy_magic_21_0.cap_res_X.n34 0.1133
R7255 two_stage_opamp_dummy_magic_21_0.cap_res_X.n29 two_stage_opamp_dummy_magic_21_0.cap_res_X.t22 0.00152174
R7256 two_stage_opamp_dummy_magic_21_0.cap_res_X.n30 two_stage_opamp_dummy_magic_21_0.cap_res_X.t45 0.00152174
R7257 two_stage_opamp_dummy_magic_21_0.cap_res_X.n31 two_stage_opamp_dummy_magic_21_0.cap_res_X.t9 0.00152174
R7258 two_stage_opamp_dummy_magic_21_0.cap_res_X.n32 two_stage_opamp_dummy_magic_21_0.cap_res_X.t111 0.00152174
R7259 two_stage_opamp_dummy_magic_21_0.cap_res_X.n33 two_stage_opamp_dummy_magic_21_0.cap_res_X.t71 0.00152174
R7260 two_stage_opamp_dummy_magic_21_0.cap_res_X.n34 two_stage_opamp_dummy_magic_21_0.cap_res_X.t95 0.00152174
R7261 two_stage_opamp_dummy_magic_21_0.cap_res_X.n0 two_stage_opamp_dummy_magic_21_0.cap_res_X.t98 0.00152174
R7262 two_stage_opamp_dummy_magic_21_0.cap_res_X.n1 two_stage_opamp_dummy_magic_21_0.cap_res_X.t59 0.00152174
R7263 two_stage_opamp_dummy_magic_21_0.cap_res_X.n2 two_stage_opamp_dummy_magic_21_0.cap_res_X.t25 0.00152174
R7264 two_stage_opamp_dummy_magic_21_0.cap_res_X.n3 two_stage_opamp_dummy_magic_21_0.cap_res_X.t132 0.00152174
R7265 two_stage_opamp_dummy_magic_21_0.cap_res_X.n4 two_stage_opamp_dummy_magic_21_0.cap_res_X.t81 0.00152174
R7266 two_stage_opamp_dummy_magic_21_0.cap_res_X.n5 two_stage_opamp_dummy_magic_21_0.cap_res_X.t43 0.00152174
R7267 two_stage_opamp_dummy_magic_21_0.cap_res_X.n6 two_stage_opamp_dummy_magic_21_0.cap_res_X.t12 0.00152174
R7268 two_stage_opamp_dummy_magic_21_0.cap_res_X.n7 two_stage_opamp_dummy_magic_21_0.cap_res_X.t102 0.00152174
R7269 two_stage_opamp_dummy_magic_21_0.cap_res_X.n8 two_stage_opamp_dummy_magic_21_0.cap_res_X.t62 0.00152174
R7270 two_stage_opamp_dummy_magic_21_0.cap_res_X.n9 two_stage_opamp_dummy_magic_21_0.cap_res_X.t32 0.00152174
R7271 two_stage_opamp_dummy_magic_21_0.cap_res_X.n10 two_stage_opamp_dummy_magic_21_0.cap_res_X.t29 0.00152174
R7272 two_stage_opamp_dummy_magic_21_0.cap_res_X.n11 two_stage_opamp_dummy_magic_21_0.cap_res_X.t63 0.00152174
R7273 two_stage_opamp_dummy_magic_21_0.cap_res_X.n12 two_stage_opamp_dummy_magic_21_0.cap_res_X.t23 0.00152174
R7274 two_stage_opamp_dummy_magic_21_0.cap_res_X.n13 two_stage_opamp_dummy_magic_21_0.cap_res_X.t125 0.00152174
R7275 two_stage_opamp_dummy_magic_21_0.cap_res_X.n14 two_stage_opamp_dummy_magic_21_0.cap_res_X.t18 0.00152174
R7276 two_stage_opamp_dummy_magic_21_0.cap_res_X.n15 two_stage_opamp_dummy_magic_21_0.cap_res_X.t121 0.00152174
R7277 two_stage_opamp_dummy_magic_21_0.cap_res_X.n16 two_stage_opamp_dummy_magic_21_0.cap_res_X.t79 0.00152174
R7278 two_stage_opamp_dummy_magic_21_0.cap_res_X.n17 two_stage_opamp_dummy_magic_21_0.cap_res_X.t36 0.00152174
R7279 two_stage_opamp_dummy_magic_21_0.cap_res_X.n18 two_stage_opamp_dummy_magic_21_0.cap_res_X.t74 0.00152174
R7280 two_stage_opamp_dummy_magic_21_0.cap_res_X.n19 two_stage_opamp_dummy_magic_21_0.cap_res_X.t34 0.00152174
R7281 two_stage_opamp_dummy_magic_21_0.cap_res_X.n20 two_stage_opamp_dummy_magic_21_0.cap_res_X.t137 0.00152174
R7282 two_stage_opamp_dummy_magic_21_0.cap_res_X.n21 two_stage_opamp_dummy_magic_21_0.cap_res_X.t28 0.00152174
R7283 two_stage_opamp_dummy_magic_21_0.cap_res_X.n22 two_stage_opamp_dummy_magic_21_0.cap_res_X.t130 0.00152174
R7284 two_stage_opamp_dummy_magic_21_0.cap_res_X.n23 two_stage_opamp_dummy_magic_21_0.cap_res_X.t109 0.00152174
R7285 two_stage_opamp_dummy_magic_21_0.cap_res_X.n24 two_stage_opamp_dummy_magic_21_0.cap_res_X.t4 0.00152174
R7286 two_stage_opamp_dummy_magic_21_0.cap_res_X.n25 two_stage_opamp_dummy_magic_21_0.cap_res_X.t105 0.00152174
R7287 two_stage_opamp_dummy_magic_21_0.cap_res_X.n26 two_stage_opamp_dummy_magic_21_0.cap_res_X.t1 0.00152174
R7288 two_stage_opamp_dummy_magic_21_0.cap_res_X.n27 two_stage_opamp_dummy_magic_21_0.cap_res_X.t37 0.00152174
R7289 two_stage_opamp_dummy_magic_21_0.cap_res_X.n28 two_stage_opamp_dummy_magic_21_0.cap_res_X.t17 0.00152174
R7290 two_stage_opamp_dummy_magic_21_0.cap_res_X.t54 two_stage_opamp_dummy_magic_21_0.cap_res_X.n35 0.00152174
R7291 bgr_0.cap_res1.t20 bgr_0.cap_res1.t9 121.245
R7292 bgr_0.cap_res1.t15 bgr_0.cap_res1.t18 0.1603
R7293 bgr_0.cap_res1.t8 bgr_0.cap_res1.t14 0.1603
R7294 bgr_0.cap_res1.t13 bgr_0.cap_res1.t17 0.1603
R7295 bgr_0.cap_res1.t6 bgr_0.cap_res1.t12 0.1603
R7296 bgr_0.cap_res1.t0 bgr_0.cap_res1.t5 0.1603
R7297 bgr_0.cap_res1.n1 bgr_0.cap_res1.t16 0.159278
R7298 bgr_0.cap_res1.n2 bgr_0.cap_res1.t1 0.159278
R7299 bgr_0.cap_res1.n3 bgr_0.cap_res1.t7 0.159278
R7300 bgr_0.cap_res1.n4 bgr_0.cap_res1.t2 0.159278
R7301 bgr_0.cap_res1.n4 bgr_0.cap_res1.t15 0.1368
R7302 bgr_0.cap_res1.n4 bgr_0.cap_res1.t11 0.1368
R7303 bgr_0.cap_res1.n3 bgr_0.cap_res1.t8 0.1368
R7304 bgr_0.cap_res1.n3 bgr_0.cap_res1.t4 0.1368
R7305 bgr_0.cap_res1.n2 bgr_0.cap_res1.t13 0.1368
R7306 bgr_0.cap_res1.n2 bgr_0.cap_res1.t10 0.1368
R7307 bgr_0.cap_res1.n1 bgr_0.cap_res1.t6 0.1368
R7308 bgr_0.cap_res1.n1 bgr_0.cap_res1.t3 0.1368
R7309 bgr_0.cap_res1.n0 bgr_0.cap_res1.t0 0.1368
R7310 bgr_0.cap_res1.n0 bgr_0.cap_res1.t19 0.1368
R7311 bgr_0.cap_res1.t16 bgr_0.cap_res1.n0 0.00152174
R7312 bgr_0.cap_res1.t1 bgr_0.cap_res1.n1 0.00152174
R7313 bgr_0.cap_res1.t7 bgr_0.cap_res1.n2 0.00152174
R7314 bgr_0.cap_res1.t2 bgr_0.cap_res1.n3 0.00152174
R7315 bgr_0.cap_res1.t9 bgr_0.cap_res1.n4 0.00152174
R7316 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R7317 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R7318 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R7319 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 310.488
R7320 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R7321 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R7322 bgr_0.V_mir2.n2 bgr_0.V_mir2.t14 278.312
R7323 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R7324 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R7325 bgr_0.V_mir2.n18 bgr_0.V_mir2.t10 184.097
R7326 bgr_0.V_mir2.n11 bgr_0.V_mir2.t8 184.097
R7327 bgr_0.V_mir2.n6 bgr_0.V_mir2.t0 184.097
R7328 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R7329 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R7330 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R7331 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R7332 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R7333 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R7334 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R7335 bgr_0.V_mir2.n17 bgr_0.V_mir2.t6 120.501
R7336 bgr_0.V_mir2.n9 bgr_0.V_mir2.t18 120.501
R7337 bgr_0.V_mir2.n10 bgr_0.V_mir2.t2 120.501
R7338 bgr_0.V_mir2.n4 bgr_0.V_mir2.t17 120.501
R7339 bgr_0.V_mir2.n5 bgr_0.V_mir2.t4 120.501
R7340 bgr_0.V_mir2.n1 bgr_0.V_mir2.t16 48.0005
R7341 bgr_0.V_mir2.n1 bgr_0.V_mir2.t12 48.0005
R7342 bgr_0.V_mir2.n0 bgr_0.V_mir2.t15 48.0005
R7343 bgr_0.V_mir2.n0 bgr_0.V_mir2.t13 48.0005
R7344 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R7345 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R7346 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R7347 bgr_0.V_mir2.n12 bgr_0.V_mir2.t3 39.4005
R7348 bgr_0.V_mir2.n12 bgr_0.V_mir2.t9 39.4005
R7349 bgr_0.V_mir2.n7 bgr_0.V_mir2.t5 39.4005
R7350 bgr_0.V_mir2.n7 bgr_0.V_mir2.t1 39.4005
R7351 bgr_0.V_mir2.n20 bgr_0.V_mir2.t7 39.4005
R7352 bgr_0.V_mir2.t11 bgr_0.V_mir2.n20 39.4005
R7353 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R7354 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R7355 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R7356 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R7357 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R7358 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R7359 bgr_0.Vin-.n8 bgr_0.Vin-.t12 688.859
R7360 bgr_0.Vin-.n10 bgr_0.Vin-.n9 514.134
R7361 bgr_0.Vin-.n7 bgr_0.Vin-.n6 351.522
R7362 bgr_0.Vin-.n12 bgr_0.Vin-.n11 213.4
R7363 bgr_0.Vin-.n8 bgr_0.Vin-.t8 174.726
R7364 bgr_0.Vin-.n9 bgr_0.Vin-.t10 174.726
R7365 bgr_0.Vin-.n10 bgr_0.Vin-.t9 174.726
R7366 bgr_0.Vin-.n11 bgr_0.Vin-.t11 174.726
R7367 bgr_0.Vin-.n5 bgr_0.Vin-.n3 173.029
R7368 bgr_0.Vin-.n5 bgr_0.Vin-.n4 168.654
R7369 bgr_0.Vin-.n22 bgr_0.Vin-.n21 141.667
R7370 bgr_0.Vin-.n9 bgr_0.Vin-.n8 128.534
R7371 bgr_0.Vin-.n11 bgr_0.Vin-.n10 128.534
R7372 bgr_0.Vin-.n13 bgr_0.Vin-.t7 119.099
R7373 bgr_0.Vin-.n23 bgr_0.Vin-.n22 84.0884
R7374 bgr_0.Vin-.n18 bgr_0.Vin-.n17 83.5719
R7375 bgr_0.Vin-.n19 bgr_0.Vin-.n0 83.5719
R7376 bgr_0.Vin-.n20 bgr_0.Vin-.n1 83.5719
R7377 bgr_0.Vin-.n15 bgr_0.Vin-.t6 65.0299
R7378 bgr_0.Vin-.n6 bgr_0.Vin-.t5 39.4005
R7379 bgr_0.Vin-.n6 bgr_0.Vin-.t4 39.4005
R7380 bgr_0.Vin-.n14 bgr_0.Vin-.n13 28.813
R7381 bgr_0.Vin-.n19 bgr_0.Vin-.n18 26.074
R7382 bgr_0.Vin-.n20 bgr_0.Vin-.n19 26.074
R7383 bgr_0.Vin-.n22 bgr_0.Vin-.n20 26.074
R7384 bgr_0.Vin-.n13 bgr_0.Vin-.n12 16.188
R7385 bgr_0.Vin-.n4 bgr_0.Vin-.t0 13.1338
R7386 bgr_0.Vin-.n4 bgr_0.Vin-.t2 13.1338
R7387 bgr_0.Vin-.n3 bgr_0.Vin-.t3 13.1338
R7388 bgr_0.Vin-.n3 bgr_0.Vin-.t1 13.1338
R7389 bgr_0.Vin-.n12 bgr_0.Vin-.n7 11.2193
R7390 bgr_0.Vin-.n7 bgr_0.Vin-.n5 3.8755
R7391 bgr_0.Vin-.n24 bgr_0.Vin-.n23 1.56836
R7392 bgr_0.Vin-.n17 bgr_0.Vin-.n15 1.56363
R7393 bgr_0.Vin-.n25 bgr_0.Vin-.n24 1.5505
R7394 bgr_0.Vin-.n16 bgr_0.Vin-.n2 1.5505
R7395 bgr_0.Vin-.n23 bgr_0.Vin-.n1 1.14402
R7396 bgr_0.Vin-.n16 bgr_0.Vin-.n0 0.885803
R7397 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.77514
R7398 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n0 0.756696
R7399 bgr_0.Vin-.n25 bgr_0.Vin-.n1 0.701365
R7400 bgr_0.Vin-.n15 bgr_0.Vin-.n14 0.530034
R7401 bgr_0.Vin-.n18 bgr_0.Vin-.t6 0.290206
R7402 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n25 0.203382
R7403 bgr_0.Vin-.n24 bgr_0.Vin-.n2 0.0183571
R7404 bgr_0.Vin-.n14 bgr_0.Vin-.n2 0.00817857
R7405 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 229.562
R7406 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R7407 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R7408 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R7409 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 228.938
R7410 bgr_0.V_p_1.n0 bgr_0.V_p_1.t5 98.7279
R7411 bgr_0.V_p_1.n5 bgr_0.V_p_1.t8 48.0005
R7412 bgr_0.V_p_1.n5 bgr_0.V_p_1.t0 48.0005
R7413 bgr_0.V_p_1.n4 bgr_0.V_p_1.t10 48.0005
R7414 bgr_0.V_p_1.n4 bgr_0.V_p_1.t2 48.0005
R7415 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R7416 bgr_0.V_p_1.n3 bgr_0.V_p_1.t6 48.0005
R7417 bgr_0.V_p_1.n2 bgr_0.V_p_1.t9 48.0005
R7418 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R7419 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R7420 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R7421 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R7422 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n0 344.837
R7423 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n1 344.274
R7424 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n3 292.5
R7425 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t16 122.754
R7426 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n7 118.861
R7427 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n9 118.861
R7428 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n13 118.861
R7429 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n16 118.861
R7430 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n19 118.861
R7431 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n2 52.3363
R7432 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n4 52.1563
R7433 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n22 42.3755
R7434 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t1 39.4005
R7435 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t14 39.4005
R7436 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t0 39.4005
R7437 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t3 39.4005
R7438 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t15 39.4005
R7439 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t2 39.4005
R7440 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t11 19.7005
R7441 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t6 19.7005
R7442 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t10 19.7005
R7443 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t5 19.7005
R7444 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t12 19.7005
R7445 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t7 19.7005
R7446 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t13 19.7005
R7447 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t8 19.7005
R7448 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t4 19.7005
R7449 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t9 19.7005
R7450 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n21 6.2505
R7451 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n8 5.60467
R7452 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n18 5.54217
R7453 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n6 5.54217
R7454 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n10 5.04217
R7455 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n12 5.04217
R7456 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n5 5.04217
R7457 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n20 5.04217
R7458 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n6 4.97967
R7459 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n14 4.97967
R7460 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n17 4.97967
R7461 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n15 0.563
R7462 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n6 0.563
R7463 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n11 0.563
R7464 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n5 0.563
R7465 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n5 0.563
R7466 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n0 144.827
R7467 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n1 134.577
R7468 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t0 120.504
R7469 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n2 37.4067
R7470 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n20 35.4067
R7471 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n5 24.288
R7472 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n7 24.288
R7473 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n11 24.288
R7474 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n14 24.288
R7475 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n17 24.288
R7476 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t13 24.0005
R7477 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t11 24.0005
R7478 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t14 24.0005
R7479 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t12 24.0005
R7480 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t4 8.0005
R7481 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t10 8.0005
R7482 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t3 8.0005
R7483 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t9 8.0005
R7484 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t7 8.0005
R7485 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t2 8.0005
R7486 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t6 8.0005
R7487 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t1 8.0005
R7488 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t5 8.0005
R7489 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t8 8.0005
R7490 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n19 6.0005
R7491 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n16 5.7505
R7492 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n4 5.7505
R7493 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n6 5.7505
R7494 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n8 5.188
R7495 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n4 5.188
R7496 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n10 5.188
R7497 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n12 5.188
R7498 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n3 5.188
R7499 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n15 5.188
R7500 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n18 5.188
R7501 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n13 0.563
R7502 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n4 0.563
R7503 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n9 0.563
R7504 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n3 0.563
R7505 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n3 0.563
R7506 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n21 0.047375
R7507 VIN-.n0 VIN-.t2 1000.38
R7508 VIN- VIN-.n9 433.019
R7509 VIN-.n9 VIN-.t7 273.134
R7510 VIN-.n0 VIN-.t4 273.134
R7511 VIN-.n1 VIN-.t9 273.134
R7512 VIN-.n2 VIN-.t3 273.134
R7513 VIN-.n3 VIN-.t8 273.134
R7514 VIN-.n4 VIN-.t6 273.134
R7515 VIN-.n5 VIN-.t0 273.134
R7516 VIN-.n6 VIN-.t5 273.134
R7517 VIN-.n7 VIN-.t10 273.134
R7518 VIN-.n8 VIN-.t1 273.134
R7519 VIN-.n9 VIN-.n8 176.733
R7520 VIN-.n8 VIN-.n7 176.733
R7521 VIN-.n7 VIN-.n6 176.733
R7522 VIN-.n6 VIN-.n5 176.733
R7523 VIN-.n5 VIN-.n4 176.733
R7524 VIN-.n4 VIN-.n3 176.733
R7525 VIN-.n3 VIN-.n2 176.733
R7526 VIN-.n2 VIN-.n1 176.733
R7527 VIN-.n1 VIN-.n0 176.733
R7528 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R7529 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R7530 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R7531 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R7532 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R7533 bgr_0.START_UP.n0 bgr_0.START_UP.t5 130.001
R7534 bgr_0.START_UP.n0 bgr_0.START_UP.t4 81.7074
R7535 bgr_0.START_UP bgr_0.START_UP.n0 36.9489
R7536 bgr_0.START_UP bgr_0.START_UP.n5 13.4693
R7537 bgr_0.START_UP.n1 bgr_0.START_UP.t0 13.1338
R7538 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R7539 bgr_0.START_UP.n2 bgr_0.START_UP.t1 13.1338
R7540 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R7541 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R7542 two_stage_opamp_dummy_magic_21_0.V_err_gate.n2 two_stage_opamp_dummy_magic_21_0.V_err_gate.n26 594.301
R7543 two_stage_opamp_dummy_magic_21_0.V_err_gate.n28 two_stage_opamp_dummy_magic_21_0.V_err_gate.n27 594.301
R7544 two_stage_opamp_dummy_magic_21_0.V_err_gate.n30 two_stage_opamp_dummy_magic_21_0.V_err_gate.n29 594.301
R7545 two_stage_opamp_dummy_magic_21_0.V_err_gate.n32 two_stage_opamp_dummy_magic_21_0.V_err_gate.n31 594.301
R7546 two_stage_opamp_dummy_magic_21_0.V_err_gate.n34 two_stage_opamp_dummy_magic_21_0.V_err_gate.n33 594.301
R7547 two_stage_opamp_dummy_magic_21_0.V_err_gate.n36 two_stage_opamp_dummy_magic_21_0.V_err_gate.n35 594.301
R7548 two_stage_opamp_dummy_magic_21_0.V_err_gate.n7 two_stage_opamp_dummy_magic_21_0.V_err_gate.t24 289.2
R7549 two_stage_opamp_dummy_magic_21_0.V_err_gate.n17 two_stage_opamp_dummy_magic_21_0.V_err_gate.t32 224.934
R7550 two_stage_opamp_dummy_magic_21_0.V_err_gate.n24 two_stage_opamp_dummy_magic_21_0.V_err_gate.n23 176.733
R7551 two_stage_opamp_dummy_magic_21_0.V_err_gate.n23 two_stage_opamp_dummy_magic_21_0.V_err_gate.n22 176.733
R7552 two_stage_opamp_dummy_magic_21_0.V_err_gate.n22 two_stage_opamp_dummy_magic_21_0.V_err_gate.n21 176.733
R7553 two_stage_opamp_dummy_magic_21_0.V_err_gate.n21 two_stage_opamp_dummy_magic_21_0.V_err_gate.n20 176.733
R7554 two_stage_opamp_dummy_magic_21_0.V_err_gate.n20 two_stage_opamp_dummy_magic_21_0.V_err_gate.n19 176.733
R7555 two_stage_opamp_dummy_magic_21_0.V_err_gate.n19 two_stage_opamp_dummy_magic_21_0.V_err_gate.n18 176.733
R7556 two_stage_opamp_dummy_magic_21_0.V_err_gate.n18 two_stage_opamp_dummy_magic_21_0.V_err_gate.n17 176.733
R7557 two_stage_opamp_dummy_magic_21_0.V_err_gate.n8 two_stage_opamp_dummy_magic_21_0.V_err_gate.n7 176.733
R7558 two_stage_opamp_dummy_magic_21_0.V_err_gate.n9 two_stage_opamp_dummy_magic_21_0.V_err_gate.n8 176.733
R7559 two_stage_opamp_dummy_magic_21_0.V_err_gate.n10 two_stage_opamp_dummy_magic_21_0.V_err_gate.n9 176.733
R7560 two_stage_opamp_dummy_magic_21_0.V_err_gate.n11 two_stage_opamp_dummy_magic_21_0.V_err_gate.n10 176.733
R7561 two_stage_opamp_dummy_magic_21_0.V_err_gate.n12 two_stage_opamp_dummy_magic_21_0.V_err_gate.n11 176.733
R7562 two_stage_opamp_dummy_magic_21_0.V_err_gate.n13 two_stage_opamp_dummy_magic_21_0.V_err_gate.n12 176.733
R7563 two_stage_opamp_dummy_magic_21_0.V_err_gate.n14 two_stage_opamp_dummy_magic_21_0.V_err_gate.n13 176.733
R7564 two_stage_opamp_dummy_magic_21_0.V_err_gate.n15 two_stage_opamp_dummy_magic_21_0.V_err_gate.n14 176.733
R7565 two_stage_opamp_dummy_magic_21_0.V_err_gate.n16 two_stage_opamp_dummy_magic_21_0.V_err_gate.n15 176.733
R7566 two_stage_opamp_dummy_magic_21_0.V_err_gate two_stage_opamp_dummy_magic_21_0.V_err_gate.n6 175.013
R7567 two_stage_opamp_dummy_magic_21_0.V_err_gate two_stage_opamp_dummy_magic_21_0.V_err_gate.n25 161.869
R7568 two_stage_opamp_dummy_magic_21_0.V_err_gate.n24 two_stage_opamp_dummy_magic_21_0.V_err_gate.t20 112.468
R7569 two_stage_opamp_dummy_magic_21_0.V_err_gate.n23 two_stage_opamp_dummy_magic_21_0.V_err_gate.t31 112.468
R7570 two_stage_opamp_dummy_magic_21_0.V_err_gate.n22 two_stage_opamp_dummy_magic_21_0.V_err_gate.t25 112.468
R7571 two_stage_opamp_dummy_magic_21_0.V_err_gate.n21 two_stage_opamp_dummy_magic_21_0.V_err_gate.t16 112.468
R7572 two_stage_opamp_dummy_magic_21_0.V_err_gate.n20 two_stage_opamp_dummy_magic_21_0.V_err_gate.t27 112.468
R7573 two_stage_opamp_dummy_magic_21_0.V_err_gate.n19 two_stage_opamp_dummy_magic_21_0.V_err_gate.t18 112.468
R7574 two_stage_opamp_dummy_magic_21_0.V_err_gate.n18 two_stage_opamp_dummy_magic_21_0.V_err_gate.t29 112.468
R7575 two_stage_opamp_dummy_magic_21_0.V_err_gate.n17 two_stage_opamp_dummy_magic_21_0.V_err_gate.t22 112.468
R7576 two_stage_opamp_dummy_magic_21_0.V_err_gate.n7 two_stage_opamp_dummy_magic_21_0.V_err_gate.t15 112.468
R7577 two_stage_opamp_dummy_magic_21_0.V_err_gate.n8 two_stage_opamp_dummy_magic_21_0.V_err_gate.t21 112.468
R7578 two_stage_opamp_dummy_magic_21_0.V_err_gate.n9 two_stage_opamp_dummy_magic_21_0.V_err_gate.t14 112.468
R7579 two_stage_opamp_dummy_magic_21_0.V_err_gate.n10 two_stage_opamp_dummy_magic_21_0.V_err_gate.t26 112.468
R7580 two_stage_opamp_dummy_magic_21_0.V_err_gate.n11 two_stage_opamp_dummy_magic_21_0.V_err_gate.t17 112.468
R7581 two_stage_opamp_dummy_magic_21_0.V_err_gate.n12 two_stage_opamp_dummy_magic_21_0.V_err_gate.t28 112.468
R7582 two_stage_opamp_dummy_magic_21_0.V_err_gate.n13 two_stage_opamp_dummy_magic_21_0.V_err_gate.t19 112.468
R7583 two_stage_opamp_dummy_magic_21_0.V_err_gate.n14 two_stage_opamp_dummy_magic_21_0.V_err_gate.t30 112.468
R7584 two_stage_opamp_dummy_magic_21_0.V_err_gate.n15 two_stage_opamp_dummy_magic_21_0.V_err_gate.t23 112.468
R7585 two_stage_opamp_dummy_magic_21_0.V_err_gate.n16 two_stage_opamp_dummy_magic_21_0.V_err_gate.t33 112.468
R7586 two_stage_opamp_dummy_magic_21_0.V_err_gate.n26 two_stage_opamp_dummy_magic_21_0.V_err_gate.t6 78.8005
R7587 two_stage_opamp_dummy_magic_21_0.V_err_gate.n26 two_stage_opamp_dummy_magic_21_0.V_err_gate.t13 78.8005
R7588 two_stage_opamp_dummy_magic_21_0.V_err_gate.n27 two_stage_opamp_dummy_magic_21_0.V_err_gate.t3 78.8005
R7589 two_stage_opamp_dummy_magic_21_0.V_err_gate.n27 two_stage_opamp_dummy_magic_21_0.V_err_gate.t2 78.8005
R7590 two_stage_opamp_dummy_magic_21_0.V_err_gate.n29 two_stage_opamp_dummy_magic_21_0.V_err_gate.t5 78.8005
R7591 two_stage_opamp_dummy_magic_21_0.V_err_gate.n29 two_stage_opamp_dummy_magic_21_0.V_err_gate.t4 78.8005
R7592 two_stage_opamp_dummy_magic_21_0.V_err_gate.n31 two_stage_opamp_dummy_magic_21_0.V_err_gate.t0 78.8005
R7593 two_stage_opamp_dummy_magic_21_0.V_err_gate.n31 two_stage_opamp_dummy_magic_21_0.V_err_gate.t1 78.8005
R7594 two_stage_opamp_dummy_magic_21_0.V_err_gate.n33 two_stage_opamp_dummy_magic_21_0.V_err_gate.t8 78.8005
R7595 two_stage_opamp_dummy_magic_21_0.V_err_gate.n33 two_stage_opamp_dummy_magic_21_0.V_err_gate.t7 78.8005
R7596 two_stage_opamp_dummy_magic_21_0.V_err_gate.n35 two_stage_opamp_dummy_magic_21_0.V_err_gate.t12 78.8005
R7597 two_stage_opamp_dummy_magic_21_0.V_err_gate.n35 two_stage_opamp_dummy_magic_21_0.V_err_gate.t9 78.8005
R7598 two_stage_opamp_dummy_magic_21_0.V_err_gate.n25 two_stage_opamp_dummy_magic_21_0.V_err_gate.n24 56.2338
R7599 two_stage_opamp_dummy_magic_21_0.V_err_gate.n25 two_stage_opamp_dummy_magic_21_0.V_err_gate.n16 56.2338
R7600 two_stage_opamp_dummy_magic_21_0.V_err_gate.n6 two_stage_opamp_dummy_magic_21_0.V_err_gate.t10 24.0005
R7601 two_stage_opamp_dummy_magic_21_0.V_err_gate.n6 two_stage_opamp_dummy_magic_21_0.V_err_gate.t11 24.0005
R7602 two_stage_opamp_dummy_magic_21_0.V_err_gate two_stage_opamp_dummy_magic_21_0.V_err_gate.n3 6.89112
R7603 two_stage_opamp_dummy_magic_21_0.V_err_gate.n4 two_stage_opamp_dummy_magic_21_0.V_err_gate.n2 5.41717
R7604 two_stage_opamp_dummy_magic_21_0.V_err_gate.n36 two_stage_opamp_dummy_magic_21_0.V_err_gate.n1 5.22967
R7605 two_stage_opamp_dummy_magic_21_0.V_err_gate.n0 two_stage_opamp_dummy_magic_21_0.V_err_gate.n2 5.22967
R7606 two_stage_opamp_dummy_magic_21_0.V_err_gate.n4 two_stage_opamp_dummy_magic_21_0.V_err_gate.n28 4.85467
R7607 two_stage_opamp_dummy_magic_21_0.V_err_gate.n5 two_stage_opamp_dummy_magic_21_0.V_err_gate.n30 4.85467
R7608 two_stage_opamp_dummy_magic_21_0.V_err_gate.n32 two_stage_opamp_dummy_magic_21_0.V_err_gate.n5 4.85467
R7609 two_stage_opamp_dummy_magic_21_0.V_err_gate.n34 two_stage_opamp_dummy_magic_21_0.V_err_gate.n3 4.85467
R7610 two_stage_opamp_dummy_magic_21_0.V_err_gate.n3 two_stage_opamp_dummy_magic_21_0.V_err_gate.n36 4.85467
R7611 two_stage_opamp_dummy_magic_21_0.V_err_gate.n28 two_stage_opamp_dummy_magic_21_0.V_err_gate.n0 4.66717
R7612 two_stage_opamp_dummy_magic_21_0.V_err_gate.n30 two_stage_opamp_dummy_magic_21_0.V_err_gate.n0 4.66717
R7613 two_stage_opamp_dummy_magic_21_0.V_err_gate.n1 two_stage_opamp_dummy_magic_21_0.V_err_gate.n32 4.66717
R7614 two_stage_opamp_dummy_magic_21_0.V_err_gate.n1 two_stage_opamp_dummy_magic_21_0.V_err_gate.n34 4.66717
R7615 two_stage_opamp_dummy_magic_21_0.V_err_gate.n1 two_stage_opamp_dummy_magic_21_0.V_err_gate.n0 1.688
R7616 two_stage_opamp_dummy_magic_21_0.V_err_gate.n5 two_stage_opamp_dummy_magic_21_0.V_err_gate.n3 1.1255
R7617 two_stage_opamp_dummy_magic_21_0.V_err_gate.n5 two_stage_opamp_dummy_magic_21_0.V_err_gate.n4 1.1255
R7618 two_stage_opamp_dummy_magic_21_0.VD3.n26 two_stage_opamp_dummy_magic_21_0.VD3.t23 672.293
R7619 two_stage_opamp_dummy_magic_21_0.VD3.n29 two_stage_opamp_dummy_magic_21_0.VD3.t20 672.293
R7620 two_stage_opamp_dummy_magic_21_0.VD3.t24 two_stage_opamp_dummy_magic_21_0.VD3.n27 213.131
R7621 two_stage_opamp_dummy_magic_21_0.VD3.n28 two_stage_opamp_dummy_magic_21_0.VD3.t21 213.131
R7622 two_stage_opamp_dummy_magic_21_0.VD3.t0 two_stage_opamp_dummy_magic_21_0.VD3.t24 146.155
R7623 two_stage_opamp_dummy_magic_21_0.VD3.t6 two_stage_opamp_dummy_magic_21_0.VD3.t0 146.155
R7624 two_stage_opamp_dummy_magic_21_0.VD3.t14 two_stage_opamp_dummy_magic_21_0.VD3.t6 146.155
R7625 two_stage_opamp_dummy_magic_21_0.VD3.t10 two_stage_opamp_dummy_magic_21_0.VD3.t14 146.155
R7626 two_stage_opamp_dummy_magic_21_0.VD3.t16 two_stage_opamp_dummy_magic_21_0.VD3.t10 146.155
R7627 two_stage_opamp_dummy_magic_21_0.VD3.t18 two_stage_opamp_dummy_magic_21_0.VD3.t16 146.155
R7628 two_stage_opamp_dummy_magic_21_0.VD3.t2 two_stage_opamp_dummy_magic_21_0.VD3.t18 146.155
R7629 two_stage_opamp_dummy_magic_21_0.VD3.t8 two_stage_opamp_dummy_magic_21_0.VD3.t2 146.155
R7630 two_stage_opamp_dummy_magic_21_0.VD3.t4 two_stage_opamp_dummy_magic_21_0.VD3.t8 146.155
R7631 two_stage_opamp_dummy_magic_21_0.VD3.t12 two_stage_opamp_dummy_magic_21_0.VD3.t4 146.155
R7632 two_stage_opamp_dummy_magic_21_0.VD3.t21 two_stage_opamp_dummy_magic_21_0.VD3.t12 146.155
R7633 two_stage_opamp_dummy_magic_21_0.VD3.n27 two_stage_opamp_dummy_magic_21_0.VD3.t25 76.2576
R7634 two_stage_opamp_dummy_magic_21_0.VD3.n28 two_stage_opamp_dummy_magic_21_0.VD3.t22 76.2576
R7635 two_stage_opamp_dummy_magic_21_0.VD3.n1 two_stage_opamp_dummy_magic_21_0.VD3.n0 71.513
R7636 two_stage_opamp_dummy_magic_21_0.VD3.n24 two_stage_opamp_dummy_magic_21_0.VD3.n23 71.513
R7637 two_stage_opamp_dummy_magic_21_0.VD3.n31 two_stage_opamp_dummy_magic_21_0.VD3.n30 71.513
R7638 two_stage_opamp_dummy_magic_21_0.VD3.n33 two_stage_opamp_dummy_magic_21_0.VD3.n32 71.513
R7639 two_stage_opamp_dummy_magic_21_0.VD3.n35 two_stage_opamp_dummy_magic_21_0.VD3.n34 71.513
R7640 two_stage_opamp_dummy_magic_21_0.VD3.n5 two_stage_opamp_dummy_magic_21_0.VD3.n4 66.0338
R7641 two_stage_opamp_dummy_magic_21_0.VD3.n8 two_stage_opamp_dummy_magic_21_0.VD3.n7 66.0338
R7642 two_stage_opamp_dummy_magic_21_0.VD3.n11 two_stage_opamp_dummy_magic_21_0.VD3.n10 66.0338
R7643 two_stage_opamp_dummy_magic_21_0.VD3.n15 two_stage_opamp_dummy_magic_21_0.VD3.n14 66.0338
R7644 two_stage_opamp_dummy_magic_21_0.VD3.n18 two_stage_opamp_dummy_magic_21_0.VD3.n17 66.0338
R7645 two_stage_opamp_dummy_magic_21_0.VD3.n21 two_stage_opamp_dummy_magic_21_0.VD3.n20 66.0338
R7646 two_stage_opamp_dummy_magic_21_0.VD3.n25 two_stage_opamp_dummy_magic_21_0.VD3.n22 14.0005
R7647 two_stage_opamp_dummy_magic_21_0.VD3.n0 two_stage_opamp_dummy_magic_21_0.VD3.t15 11.2576
R7648 two_stage_opamp_dummy_magic_21_0.VD3.n0 two_stage_opamp_dummy_magic_21_0.VD3.t11 11.2576
R7649 two_stage_opamp_dummy_magic_21_0.VD3.n23 two_stage_opamp_dummy_magic_21_0.VD3.t1 11.2576
R7650 two_stage_opamp_dummy_magic_21_0.VD3.n23 two_stage_opamp_dummy_magic_21_0.VD3.t7 11.2576
R7651 two_stage_opamp_dummy_magic_21_0.VD3.n30 two_stage_opamp_dummy_magic_21_0.VD3.t5 11.2576
R7652 two_stage_opamp_dummy_magic_21_0.VD3.n30 two_stage_opamp_dummy_magic_21_0.VD3.t13 11.2576
R7653 two_stage_opamp_dummy_magic_21_0.VD3.n32 two_stage_opamp_dummy_magic_21_0.VD3.t3 11.2576
R7654 two_stage_opamp_dummy_magic_21_0.VD3.n32 two_stage_opamp_dummy_magic_21_0.VD3.t9 11.2576
R7655 two_stage_opamp_dummy_magic_21_0.VD3.n4 two_stage_opamp_dummy_magic_21_0.VD3.t37 11.2576
R7656 two_stage_opamp_dummy_magic_21_0.VD3.n4 two_stage_opamp_dummy_magic_21_0.VD3.t33 11.2576
R7657 two_stage_opamp_dummy_magic_21_0.VD3.n7 two_stage_opamp_dummy_magic_21_0.VD3.t31 11.2576
R7658 two_stage_opamp_dummy_magic_21_0.VD3.n7 two_stage_opamp_dummy_magic_21_0.VD3.t34 11.2576
R7659 two_stage_opamp_dummy_magic_21_0.VD3.n10 two_stage_opamp_dummy_magic_21_0.VD3.t26 11.2576
R7660 two_stage_opamp_dummy_magic_21_0.VD3.n10 two_stage_opamp_dummy_magic_21_0.VD3.t28 11.2576
R7661 two_stage_opamp_dummy_magic_21_0.VD3.n14 two_stage_opamp_dummy_magic_21_0.VD3.t30 11.2576
R7662 two_stage_opamp_dummy_magic_21_0.VD3.n14 two_stage_opamp_dummy_magic_21_0.VD3.t29 11.2576
R7663 two_stage_opamp_dummy_magic_21_0.VD3.n17 two_stage_opamp_dummy_magic_21_0.VD3.t32 11.2576
R7664 two_stage_opamp_dummy_magic_21_0.VD3.n17 two_stage_opamp_dummy_magic_21_0.VD3.t35 11.2576
R7665 two_stage_opamp_dummy_magic_21_0.VD3.n20 two_stage_opamp_dummy_magic_21_0.VD3.t27 11.2576
R7666 two_stage_opamp_dummy_magic_21_0.VD3.n20 two_stage_opamp_dummy_magic_21_0.VD3.t36 11.2576
R7667 two_stage_opamp_dummy_magic_21_0.VD3.n35 two_stage_opamp_dummy_magic_21_0.VD3.t17 11.2576
R7668 two_stage_opamp_dummy_magic_21_0.VD3.t19 two_stage_opamp_dummy_magic_21_0.VD3.n35 11.2576
R7669 two_stage_opamp_dummy_magic_21_0.VD3.n31 two_stage_opamp_dummy_magic_21_0.VD3.n29 6.10467
R7670 two_stage_opamp_dummy_magic_21_0.VD3.n21 two_stage_opamp_dummy_magic_21_0.VD3.n19 5.91717
R7671 two_stage_opamp_dummy_magic_21_0.VD3.n6 two_stage_opamp_dummy_magic_21_0.VD3.n5 5.91717
R7672 two_stage_opamp_dummy_magic_21_0.VD3.n9 two_stage_opamp_dummy_magic_21_0.VD3.n5 5.91717
R7673 two_stage_opamp_dummy_magic_21_0.VD3.n26 two_stage_opamp_dummy_magic_21_0.VD3.n25 5.47967
R7674 two_stage_opamp_dummy_magic_21_0.VD3.n9 two_stage_opamp_dummy_magic_21_0.VD3.n8 5.29217
R7675 two_stage_opamp_dummy_magic_21_0.VD3.n8 two_stage_opamp_dummy_magic_21_0.VD3.n6 5.29217
R7676 two_stage_opamp_dummy_magic_21_0.VD3.n12 two_stage_opamp_dummy_magic_21_0.VD3.n11 5.29217
R7677 two_stage_opamp_dummy_magic_21_0.VD3.n11 two_stage_opamp_dummy_magic_21_0.VD3.n3 5.29217
R7678 two_stage_opamp_dummy_magic_21_0.VD3.n15 two_stage_opamp_dummy_magic_21_0.VD3.n13 5.29217
R7679 two_stage_opamp_dummy_magic_21_0.VD3.n16 two_stage_opamp_dummy_magic_21_0.VD3.n15 5.29217
R7680 two_stage_opamp_dummy_magic_21_0.VD3.n18 two_stage_opamp_dummy_magic_21_0.VD3.n2 5.29217
R7681 two_stage_opamp_dummy_magic_21_0.VD3.n19 two_stage_opamp_dummy_magic_21_0.VD3.n18 5.29217
R7682 two_stage_opamp_dummy_magic_21_0.VD3.n22 two_stage_opamp_dummy_magic_21_0.VD3.n21 5.29217
R7683 two_stage_opamp_dummy_magic_21_0.VD3.n29 two_stage_opamp_dummy_magic_21_0.VD3.n28 1.03383
R7684 two_stage_opamp_dummy_magic_21_0.VD3.n27 two_stage_opamp_dummy_magic_21_0.VD3.n26 1.03383
R7685 two_stage_opamp_dummy_magic_21_0.VD3.n34 two_stage_opamp_dummy_magic_21_0.VD3.n33 0.6255
R7686 two_stage_opamp_dummy_magic_21_0.VD3.n33 two_stage_opamp_dummy_magic_21_0.VD3.n31 0.6255
R7687 two_stage_opamp_dummy_magic_21_0.VD3.n19 two_stage_opamp_dummy_magic_21_0.VD3.n16 0.6255
R7688 two_stage_opamp_dummy_magic_21_0.VD3.n16 two_stage_opamp_dummy_magic_21_0.VD3.n3 0.6255
R7689 two_stage_opamp_dummy_magic_21_0.VD3.n6 two_stage_opamp_dummy_magic_21_0.VD3.n3 0.6255
R7690 two_stage_opamp_dummy_magic_21_0.VD3.n12 two_stage_opamp_dummy_magic_21_0.VD3.n9 0.6255
R7691 two_stage_opamp_dummy_magic_21_0.VD3.n13 two_stage_opamp_dummy_magic_21_0.VD3.n12 0.6255
R7692 two_stage_opamp_dummy_magic_21_0.VD3.n13 two_stage_opamp_dummy_magic_21_0.VD3.n2 0.6255
R7693 two_stage_opamp_dummy_magic_21_0.VD3.n22 two_stage_opamp_dummy_magic_21_0.VD3.n2 0.6255
R7694 two_stage_opamp_dummy_magic_21_0.VD3.n25 two_stage_opamp_dummy_magic_21_0.VD3.n24 0.6255
R7695 two_stage_opamp_dummy_magic_21_0.VD3.n24 two_stage_opamp_dummy_magic_21_0.VD3.n1 0.6255
R7696 two_stage_opamp_dummy_magic_21_0.VD3.n34 two_stage_opamp_dummy_magic_21_0.VD3.n1 0.6255
R7697 VIN+.n0 VIN+.t9 1001.28
R7698 VIN+ VIN+.n9 433.019
R7699 VIN+.n9 VIN+.t5 273.134
R7700 VIN+.n0 VIN+.t6 273.134
R7701 VIN+.n8 VIN+.t10 273.134
R7702 VIN+.n7 VIN+.t4 273.134
R7703 VIN+.n6 VIN+.t8 273.134
R7704 VIN+.n5 VIN+.t2 273.134
R7705 VIN+.n4 VIN+.t0 273.134
R7706 VIN+.n3 VIN+.t3 273.134
R7707 VIN+.n2 VIN+.t7 273.134
R7708 VIN+.n1 VIN+.t1 273.134
R7709 VIN+.n1 VIN+.n0 176.733
R7710 VIN+.n2 VIN+.n1 176.733
R7711 VIN+.n3 VIN+.n2 176.733
R7712 VIN+.n4 VIN+.n3 176.733
R7713 VIN+.n5 VIN+.n4 176.733
R7714 VIN+.n6 VIN+.n5 176.733
R7715 VIN+.n7 VIN+.n6 176.733
R7716 VIN+.n8 VIN+.n7 176.733
R7717 VIN+.n9 VIN+.n8 176.733
R7718 two_stage_opamp_dummy_magic_21_0.Vb2_2.n2 two_stage_opamp_dummy_magic_21_0.Vb2_2.t0 661.375
R7719 two_stage_opamp_dummy_magic_21_0.Vb2_2.n4 two_stage_opamp_dummy_magic_21_0.Vb2_2.t3 661.375
R7720 two_stage_opamp_dummy_magic_21_0.Vb2_2.t1 two_stage_opamp_dummy_magic_21_0.Vb2_2.n0 213.131
R7721 two_stage_opamp_dummy_magic_21_0.Vb2_2.n3 two_stage_opamp_dummy_magic_21_0.Vb2_2.t4 213.131
R7722 two_stage_opamp_dummy_magic_21_0.Vb2_2.n6 two_stage_opamp_dummy_magic_21_0.Vb2_2.n1 154.983
R7723 two_stage_opamp_dummy_magic_21_0.Vb2_2.t6 two_stage_opamp_dummy_magic_21_0.Vb2_2.t1 146.155
R7724 two_stage_opamp_dummy_magic_21_0.Vb2_2.t4 two_stage_opamp_dummy_magic_21_0.Vb2_2.t6 146.155
R7725 two_stage_opamp_dummy_magic_21_0.Vb2_2.t2 two_stage_opamp_dummy_magic_21_0.Vb2_2.n0 76.2576
R7726 two_stage_opamp_dummy_magic_21_0.Vb2_2.n3 two_stage_opamp_dummy_magic_21_0.Vb2_2.t5 76.2576
R7727 two_stage_opamp_dummy_magic_21_0.Vb2_2.n7 two_stage_opamp_dummy_magic_21_0.Vb2_2.n6 66.4421
R7728 two_stage_opamp_dummy_magic_21_0.Vb2_2.n1 two_stage_opamp_dummy_magic_21_0.Vb2_2.t9 21.8894
R7729 two_stage_opamp_dummy_magic_21_0.Vb2_2.n1 two_stage_opamp_dummy_magic_21_0.Vb2_2.t8 21.8894
R7730 two_stage_opamp_dummy_magic_21_0.Vb2_2.t2 two_stage_opamp_dummy_magic_21_0.Vb2_2.n7 11.2576
R7731 two_stage_opamp_dummy_magic_21_0.Vb2_2.n7 two_stage_opamp_dummy_magic_21_0.Vb2_2.t7 11.2576
R7732 two_stage_opamp_dummy_magic_21_0.Vb2_2.n5 two_stage_opamp_dummy_magic_21_0.Vb2_2.n4 5.1255
R7733 two_stage_opamp_dummy_magic_21_0.Vb2_2.n6 two_stage_opamp_dummy_magic_21_0.Vb2_2.n5 4.92067
R7734 two_stage_opamp_dummy_magic_21_0.Vb2_2.n5 two_stage_opamp_dummy_magic_21_0.Vb2_2.n2 4.7505
R7735 two_stage_opamp_dummy_magic_21_0.Vb2_2.n4 two_stage_opamp_dummy_magic_21_0.Vb2_2.n3 1.888
R7736 two_stage_opamp_dummy_magic_21_0.Vb2_2.n2 two_stage_opamp_dummy_magic_21_0.Vb2_2.n0 1.888
R7737 two_stage_opamp_dummy_magic_21_0.V_tot.n6 two_stage_opamp_dummy_magic_21_0.V_tot.n5 771.76
R7738 two_stage_opamp_dummy_magic_21_0.V_tot.n11 two_stage_opamp_dummy_magic_21_0.V_tot.n10 595.444
R7739 two_stage_opamp_dummy_magic_21_0.V_tot.n1 two_stage_opamp_dummy_magic_21_0.V_tot.n0 595.131
R7740 two_stage_opamp_dummy_magic_21_0.V_tot.n3 two_stage_opamp_dummy_magic_21_0.V_tot.n2 530.201
R7741 two_stage_opamp_dummy_magic_21_0.V_tot.n5 two_stage_opamp_dummy_magic_21_0.V_tot.n4 530.201
R7742 two_stage_opamp_dummy_magic_21_0.V_tot.n7 two_stage_opamp_dummy_magic_21_0.V_tot.n6 530.201
R7743 two_stage_opamp_dummy_magic_21_0.V_tot.n9 two_stage_opamp_dummy_magic_21_0.V_tot.n8 530.201
R7744 two_stage_opamp_dummy_magic_21_0.V_tot.n5 two_stage_opamp_dummy_magic_21_0.V_tot.t13 208.868
R7745 two_stage_opamp_dummy_magic_21_0.V_tot.n4 two_stage_opamp_dummy_magic_21_0.V_tot.t6 208.868
R7746 two_stage_opamp_dummy_magic_21_0.V_tot.n3 two_stage_opamp_dummy_magic_21_0.V_tot.t4 208.868
R7747 two_stage_opamp_dummy_magic_21_0.V_tot.n2 two_stage_opamp_dummy_magic_21_0.V_tot.t8 208.868
R7748 two_stage_opamp_dummy_magic_21_0.V_tot.n1 two_stage_opamp_dummy_magic_21_0.V_tot.t10 208.868
R7749 two_stage_opamp_dummy_magic_21_0.V_tot.n10 two_stage_opamp_dummy_magic_21_0.V_tot.t7 208.868
R7750 two_stage_opamp_dummy_magic_21_0.V_tot.n9 two_stage_opamp_dummy_magic_21_0.V_tot.t12 208.868
R7751 two_stage_opamp_dummy_magic_21_0.V_tot.n8 two_stage_opamp_dummy_magic_21_0.V_tot.t9 208.868
R7752 two_stage_opamp_dummy_magic_21_0.V_tot.n7 two_stage_opamp_dummy_magic_21_0.V_tot.t11 208.868
R7753 two_stage_opamp_dummy_magic_21_0.V_tot.n6 two_stage_opamp_dummy_magic_21_0.V_tot.t5 208.868
R7754 two_stage_opamp_dummy_magic_21_0.V_tot.n2 two_stage_opamp_dummy_magic_21_0.V_tot.n1 176.733
R7755 two_stage_opamp_dummy_magic_21_0.V_tot.n4 two_stage_opamp_dummy_magic_21_0.V_tot.n3 176.733
R7756 two_stage_opamp_dummy_magic_21_0.V_tot.n8 two_stage_opamp_dummy_magic_21_0.V_tot.n7 176.733
R7757 two_stage_opamp_dummy_magic_21_0.V_tot.n10 two_stage_opamp_dummy_magic_21_0.V_tot.n9 176.733
R7758 two_stage_opamp_dummy_magic_21_0.V_tot.n11 two_stage_opamp_dummy_magic_21_0.V_tot.t3 117.591
R7759 two_stage_opamp_dummy_magic_21_0.V_tot.n0 two_stage_opamp_dummy_magic_21_0.V_tot.t1 117.591
R7760 two_stage_opamp_dummy_magic_21_0.V_tot.n0 two_stage_opamp_dummy_magic_21_0.V_tot.t2 108.424
R7761 two_stage_opamp_dummy_magic_21_0.V_tot.t0 two_stage_opamp_dummy_magic_21_0.V_tot.n11 108.424
R7762 a_5710_2046.t0 a_5710_2046.t1 169.905
R7763 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n0 144.827
R7764 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n1 134.577
R7765 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t14 120.817
R7766 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n2 37.4067
R7767 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n21 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n20 35.4067
R7768 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n5 24.288
R7769 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n7 24.288
R7770 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n11 24.288
R7771 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n14 24.288
R7772 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n17 24.288
R7773 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t10 24.0005
R7774 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t11 24.0005
R7775 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t12 24.0005
R7776 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t13 24.0005
R7777 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t6 8.0005
R7778 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t1 8.0005
R7779 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t5 8.0005
R7780 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t0 8.0005
R7781 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t7 8.0005
R7782 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t2 8.0005
R7783 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t8 8.0005
R7784 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t3 8.0005
R7785 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t9 8.0005
R7786 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t4 8.0005
R7787 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n19 5.96925
R7788 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n16 5.7505
R7789 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n4 5.7505
R7790 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n6 5.7505
R7791 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n8 5.188
R7792 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n4 5.188
R7793 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n10 5.188
R7794 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n12 5.188
R7795 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n3 5.188
R7796 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n15 5.188
R7797 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n18 5.188
R7798 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n13 0.563
R7799 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n4 0.563
R7800 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n9 0.563
R7801 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n3 0.563
R7802 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n3 0.563
R7803 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n21 0.047375
R7804 a_14240_2056.t0 a_14240_2056.t1 169.905
R7805 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R7806 a_5190_5068.t0 a_5190_5068.t1 294.339
R7807 a_14560_4968.t0 a_14560_4968.t1 294.339
R7808 a_8570_6900.n3 a_8570_6900.n2 594.301
R7809 a_8570_6900.n5 a_8570_6900.n4 594.301
R7810 a_8570_6900.n9 a_8570_6900.n8 594.301
R7811 a_8570_6900.n12 a_8570_6900.n11 594.301
R7812 a_8570_6900.n14 a_8570_6900.n13 594.301
R7813 a_8570_6900.n16 a_8570_6900.n15 594.301
R7814 a_8570_6900.n20 a_8570_6900.n19 594.301
R7815 a_8570_6900.n22 a_8570_6900.n21 594.301
R7816 a_8570_6900.n26 a_8570_6900.n25 594.301
R7817 a_8570_6900.n33 a_8570_6900.n32 594.301
R7818 a_8570_6900.n2 a_8570_6900.t19 78.8005
R7819 a_8570_6900.n2 a_8570_6900.t16 78.8005
R7820 a_8570_6900.n4 a_8570_6900.t17 78.8005
R7821 a_8570_6900.n4 a_8570_6900.t12 78.8005
R7822 a_8570_6900.n8 a_8570_6900.t14 78.8005
R7823 a_8570_6900.n8 a_8570_6900.t10 78.8005
R7824 a_8570_6900.n11 a_8570_6900.t11 78.8005
R7825 a_8570_6900.n11 a_8570_6900.t15 78.8005
R7826 a_8570_6900.n13 a_8570_6900.t9 78.8005
R7827 a_8570_6900.n13 a_8570_6900.t1 78.8005
R7828 a_8570_6900.n15 a_8570_6900.t4 78.8005
R7829 a_8570_6900.n15 a_8570_6900.t7 78.8005
R7830 a_8570_6900.n19 a_8570_6900.t3 78.8005
R7831 a_8570_6900.n19 a_8570_6900.t5 78.8005
R7832 a_8570_6900.n21 a_8570_6900.t8 78.8005
R7833 a_8570_6900.n21 a_8570_6900.t0 78.8005
R7834 a_8570_6900.n25 a_8570_6900.t2 78.8005
R7835 a_8570_6900.n25 a_8570_6900.t6 78.8005
R7836 a_8570_6900.n33 a_8570_6900.t13 78.8005
R7837 a_8570_6900.t18 a_8570_6900.n33 78.8005
R7838 a_8570_6900.n3 a_8570_6900.n1 6.20883
R7839 a_8570_6900.n12 a_8570_6900.n0 5.91717
R7840 a_8570_6900.n6 a_8570_6900.n3 5.91717
R7841 a_8570_6900.n31 a_8570_6900.n30 5.7505
R7842 a_8570_6900.n20 a_8570_6900.n17 5.41717
R7843 a_8570_6900.n28 a_8570_6900.n16 5.41717
R7844 a_8570_6900.n23 a_8570_6900.n20 5.22967
R7845 a_8570_6900.n18 a_8570_6900.n16 5.22967
R7846 a_8570_6900.n5 a_8570_6900.n1 4.95883
R7847 a_8570_6900.n10 a_8570_6900.n9 4.95883
R7848 a_8570_6900.n32 a_8570_6900.n31 4.95883
R7849 a_8570_6900.n22 a_8570_6900.n17 4.85467
R7850 a_8570_6900.n27 a_8570_6900.n26 4.85467
R7851 a_8570_6900.n6 a_8570_6900.n5 4.66717
R7852 a_8570_6900.n9 a_8570_6900.n7 4.66717
R7853 a_8570_6900.n32 a_8570_6900.n0 4.66717
R7854 a_8570_6900.n23 a_8570_6900.n22 4.66717
R7855 a_8570_6900.n26 a_8570_6900.n24 4.66717
R7856 a_8570_6900.n18 a_8570_6900.n14 4.66717
R7857 a_8570_6900.n29 a_8570_6900.n28 4.5005
R7858 a_8570_6900.n7 a_8570_6900.n0 1.2505
R7859 a_8570_6900.n7 a_8570_6900.n6 1.2505
R7860 a_8570_6900.n10 a_8570_6900.n1 1.2505
R7861 a_8570_6900.n31 a_8570_6900.n10 1.2505
R7862 a_8570_6900.n24 a_8570_6900.n18 0.563
R7863 a_8570_6900.n24 a_8570_6900.n23 0.563
R7864 a_8570_6900.n27 a_8570_6900.n17 0.563
R7865 a_8570_6900.n28 a_8570_6900.n27 0.563
R7866 a_8570_6900.n30 a_8570_6900.n29 0.51925
R7867 a_8570_6900.n30 a_8570_6900.n12 0.446333
R7868 a_8570_6900.n29 a_8570_6900.n14 0.354667
R7869 a_12530_23988.t0 a_12530_23988.t1 178.133
R7870 a_14680_4968.t0 a_14680_4968.t1 169.905
R7871 a_7580_22380.t0 a_7580_22380.t1 178.133
R7872 a_9370_2200.n1 a_9370_2200.t0 65.3505
R7873 a_9370_2200.n3 a_9370_2200.n2 49.3505
R7874 a_9370_2200.n6 a_9370_2200.n5 49.3505
R7875 a_9370_2200.n2 a_9370_2200.t4 16.0005
R7876 a_9370_2200.n2 a_9370_2200.t2 16.0005
R7877 a_9370_2200.t3 a_9370_2200.n6 16.0005
R7878 a_9370_2200.n6 a_9370_2200.t1 16.0005
R7879 a_9370_2200.n1 a_9370_2200.n0 6.3755
R7880 a_9370_2200.n4 a_9370_2200.n1 6.1255
R7881 a_9370_2200.n5 a_9370_2200.n0 5.688
R7882 a_9370_2200.n5 a_9370_2200.n4 5.438
R7883 a_9370_2200.n3 a_9370_2200.n0 5.1255
R7884 a_9370_2200.n4 a_9370_2200.n3 4.8755
R7885 a_6810_23838.t0 a_6810_23838.t1 178.133
R7886 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R7887 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R7888 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R7889 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R7890 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R7891 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R7892 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R7893 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R7894 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R7895 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R7896 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R7897 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R7898 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R7899 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R7900 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R7901 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R7902 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R7903 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R7904 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R7905 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R7906 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R7907 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R7908 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R7909 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R7910 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R7911 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R7912 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R7913 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R7914 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R7915 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R7916 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R7917 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R7918 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R7919 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R7920 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R7921 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R7922 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R7923 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R7924 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R7925 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R7926 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R7927 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R7928 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R7929 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R7930 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R7931 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R7932 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R7933 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R7934 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R7935 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R7936 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R7937 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R7938 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R7939 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R7940 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7941 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7942 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R7943 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7944 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7945 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7946 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R7947 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7948 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7949 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7950 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7951 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R7952 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R7953 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7954 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7955 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7956 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R7957 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7958 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7959 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7960 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R7961 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7962 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7963 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7964 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R7965 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R7966 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R7967 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7968 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7969 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7970 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R7971 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7972 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7973 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7974 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R7975 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7976 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7977 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7978 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7979 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7980 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7981 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7982 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7983 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7984 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7985 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7986 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7987 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R7988 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R7989 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7990 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7991 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7992 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7993 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R7994 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R7995 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R7996 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R7997 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R7998 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R7999 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R8000 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R8001 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R8002 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R8003 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R8004 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R8005 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R8006 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R8007 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R8008 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R8009 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R8010 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R8011 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R8012 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R8013 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R8014 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R8015 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R8016 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R8017 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R8018 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R8019 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R8020 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R8021 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R8022 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R8023 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R8024 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R8025 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R8026 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R8027 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R8028 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R8029 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R8030 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R8031 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R8032 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R8033 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R8034 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R8035 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R8036 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R8037 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R8038 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R8039 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R8040 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R8041 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R8042 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R8043 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R8044 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R8045 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R8046 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R8047 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R8048 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R8049 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R8050 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R8051 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R8052 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R8053 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R8054 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R8055 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R8056 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R8057 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R8058 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R8059 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R8060 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R8061 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R8062 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R8063 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R8064 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R8065 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R8066 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R8067 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R8068 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R8069 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R8070 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R8071 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R8072 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R8073 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8074 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R8075 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R8076 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8077 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R8078 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8079 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R8080 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R8081 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R8082 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R8083 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R8084 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R8085 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R8086 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R8087 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R8088 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R8089 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R8090 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R8091 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R8092 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R8093 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R8094 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R8095 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R8096 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R8097 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R8098 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R8099 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R8100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R8101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R8102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R8106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R8108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R8109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R8110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R8111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R8112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R8113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R8114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R8115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R8116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R8117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R8118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R8121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R8124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R8125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R8130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R8133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R8134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R8135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R8136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R8137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R8138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R8139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R8141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8143 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8144 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R8145 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R8146 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R8147 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8148 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R8149 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8150 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8151 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8152 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8153 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R8154 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8155 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R8156 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R8157 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R8158 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R8159 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R8160 a_12410_22380.t0 a_12410_22380.t1 178.133
R8161 a_13060_22630.t0 a_13060_22630.t1 178.133
R8162 a_13180_23838.t0 a_13180_23838.t1 178.133
R8163 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t3 661.375
R8164 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t0 661.375
R8165 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n6 213.131
R8166 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t4 213.131
R8167 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t1 146.155
R8168 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t7 146.155
R8169 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t2 76.2576
R8170 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n7 76.2576
R8171 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n1 72.4424
R8172 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n2 66.4532
R8173 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t8 11.2576
R8174 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t5 11.2576
R8175 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t9 11.2576
R8176 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.t10 11.2576
R8177 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n4 5.1255
R8178 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n3 4.9096
R8179 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n0 4.7505
R8180 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n5 1.888
R8181 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_21_0.Vb2_Vb3.n0 1.888
R8182 a_5310_5068.t0 a_5310_5068.t1 169.905
C0 VIN- VIN+ 0.151796f
C1 VIN- two_stage_opamp_dummy_magic_21_0.V_tail_gate 0.135107f
C2 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref two_stage_opamp_dummy_magic_21_0.V_err_gate 0.492517f
C3 two_stage_opamp_dummy_magic_21_0.err_amp_out two_stage_opamp_dummy_magic_21_0.V_err_gate 0.026461f
C4 VDDA VOUT+ 13.868401f
C5 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref bgr_0.START_UP 1.36583f
C6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter m1_10050_19490# 0.013969f
C7 m2_10730_16580# bgr_0.V_TOP 0.012f
C8 two_stage_opamp_dummy_magic_21_0.VD4 VOUT+ 0.028865f
C9 m2_10730_16580# bgr_0.1st_Vout_1 0.075543f
C10 VDDA two_stage_opamp_dummy_magic_21_0.cap_res_Y 0.582903f
C11 VDDA VOUT- 13.8732f
C12 VDDA two_stage_opamp_dummy_magic_21_0.X 5.01789f
C13 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.052756f
C14 bgr_0.NFET_GATE_10uA bgr_0.1st_Vout_1 0.03875f
C15 bgr_0.V_TOP two_stage_opamp_dummy_magic_21_0.V_err_gate 0.08195f
C16 two_stage_opamp_dummy_magic_21_0.V_err_gate bgr_0.1st_Vout_1 0.041119f
C17 two_stage_opamp_dummy_magic_21_0.VD4 two_stage_opamp_dummy_magic_21_0.cap_res_Y 0.054393f
C18 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_21_0.cap_res_Y 0.010678f
C19 bgr_0.V_TOP bgr_0.START_UP 0.792764f
C20 VDDA two_stage_opamp_dummy_magic_21_0.V_tail_gate 3.83722f
C21 bgr_0.START_UP bgr_0.1st_Vout_1 0.04354f
C22 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref two_stage_opamp_dummy_magic_21_0.err_amp_out 0.289292f
C23 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_21_0.V_tail_gate 0.269369f
C24 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.351171f
C25 VOUT+ two_stage_opamp_dummy_magic_21_0.cap_res_Y 50.8468f
C26 VDDA bgr_0.NFET_GATE_10uA 0.818988f
C27 VOUT+ VOUT- 0.305434f
C28 VDDA two_stage_opamp_dummy_magic_21_0.V_err_gate 2.12648f
C29 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C30 VDDA bgr_0.START_UP 1.09181f
C31 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref bgr_0.V_TOP 0.583702f
C32 VOUT- two_stage_opamp_dummy_magic_21_0.cap_res_Y 0.028842f
C33 bgr_0.PFET_GATE_10uA bgr_0.NFET_GATE_10uA 0.012365f
C34 VOUT+ two_stage_opamp_dummy_magic_21_0.V_tail_gate 0.010408f
C35 VOUT- two_stage_opamp_dummy_magic_21_0.X 2.33193f
C36 two_stage_opamp_dummy_magic_21_0.V_tail_gate two_stage_opamp_dummy_magic_21_0.cap_res_Y 0.032733f
C37 VOUT- two_stage_opamp_dummy_magic_21_0.V_tail_gate 0.02527f
C38 two_stage_opamp_dummy_magic_21_0.V_tail_gate two_stage_opamp_dummy_magic_21_0.X 0.183919f
C39 bgr_0.V_TOP bgr_0.1st_Vout_1 2.47405f
C40 VDDA two_stage_opamp_dummy_magic_21_0.VD2 0.027746f
C41 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref VDDA 4.2164f
C42 VDDA two_stage_opamp_dummy_magic_21_0.err_amp_out 1.0994f
C43 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.V_TOP 0.055802f
C44 VIN+ two_stage_opamp_dummy_magic_21_0.V_tail_gate 0.056847f
C45 two_stage_opamp_dummy_magic_21_0.VD4 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref 0.04352f
C46 VOUT- two_stage_opamp_dummy_magic_21_0.V_err_gate 0.038208f
C47 two_stage_opamp_dummy_magic_21_0.X two_stage_opamp_dummy_magic_21_0.V_err_gate 0.161254f
C48 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_21_0.V_err_amp_ref 1.67032f
C49 two_stage_opamp_dummy_magic_21_0.V_tail_gate bgr_0.NFET_GATE_10uA 0.038519f
C50 m1_10050_19490# two_stage_opamp_dummy_magic_21_0.V_err_gate 0.091711f
C51 VDDA bgr_0.V_TOP 13.2374f
C52 two_stage_opamp_dummy_magic_21_0.V_tail_gate two_stage_opamp_dummy_magic_21_0.V_err_gate 1.43091f
C53 VDDA bgr_0.1st_Vout_1 0.896465f
C54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C55 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref VOUT+ 0.039353f
C56 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 0.221314f
C57 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_21_0.V_err_gate 3.51257f
C58 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref two_stage_opamp_dummy_magic_21_0.cap_res_Y 0.243204f
C59 bgr_0.PFET_GATE_10uA m2_9370_16580# 0.012f
C60 bgr_0.NFET_GATE_10uA bgr_0.START_UP 1.64177f
C61 two_stage_opamp_dummy_magic_21_0.X two_stage_opamp_dummy_magic_21_0.err_amp_out 0.205842f
C62 VDDA bgr_0.START_UP_NFET1 0.167059f
C63 VIN+ two_stage_opamp_dummy_magic_21_0.VD2 0.510937f
C64 two_stage_opamp_dummy_magic_21_0.VD2 two_stage_opamp_dummy_magic_21_0.V_tail_gate 0.02379f
C65 two_stage_opamp_dummy_magic_21_0.V_tail_gate two_stage_opamp_dummy_magic_21_0.err_amp_out 0.2961f
C66 two_stage_opamp_dummy_magic_21_0.VD4 VDDA 8.479321f
C67 bgr_0.PFET_GATE_10uA bgr_0.START_UP_NFET1 0.0108f
C68 bgr_0.PFET_GATE_10uA VDDA 7.97055f
C69 VIN- GNDA 1.92317f
C70 VIN+ GNDA 1.90963f
C71 VOUT- GNDA 19.93293f
C72 VOUT+ GNDA 19.982286f
C73 VDDA GNDA 0.125855p
C74 m2_10730_16580# GNDA 0.0105f $ **FLOATING
C75 m2_9370_16580# GNDA 0.010002f $ **FLOATING
C76 m1_10050_19490# GNDA 0.259273f $ **FLOATING
C77 two_stage_opamp_dummy_magic_21_0.VD2 GNDA 2.003606f
C78 two_stage_opamp_dummy_magic_21_0.err_amp_out GNDA 5.206694f
C79 two_stage_opamp_dummy_magic_21_0.cap_res_Y GNDA 33.62958f
C80 two_stage_opamp_dummy_magic_21_0.X GNDA 7.153171f
C81 two_stage_opamp_dummy_magic_21_0.V_tail_gate GNDA 8.9159f
C82 bgr_0.1st_Vout_1 GNDA 7.823503f
C83 bgr_0.START_UP GNDA 5.877827f
C84 bgr_0.START_UP_NFET1 GNDA 4.29564f
C85 two_stage_opamp_dummy_magic_21_0.V_err_gate GNDA 12.2626f
C86 bgr_0.NFET_GATE_10uA GNDA 7.923511f
C87 bgr_0.V_TOP GNDA 9.96016f
C88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.8955f
C89 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref GNDA 8.65596f
C90 bgr_0.PFET_GATE_10uA GNDA 6.602193f
C91 two_stage_opamp_dummy_magic_21_0.VD4 GNDA 5.12103f
C92 a_9370_2200.t1 GNDA 0.047649f
C93 a_9370_2200.n0 GNDA 0.318351f
C94 a_9370_2200.t0 GNDA 0.161927f
C95 a_9370_2200.n1 GNDA 0.491746f
C96 a_9370_2200.t4 GNDA 0.047649f
C97 a_9370_2200.t2 GNDA 0.047649f
C98 a_9370_2200.n2 GNDA 0.103679f
C99 a_9370_2200.n3 GNDA 0.407675f
C100 a_9370_2200.n4 GNDA 0.297965f
C101 a_9370_2200.n5 GNDA 0.42438f
C102 a_9370_2200.n6 GNDA 0.103679f
C103 a_9370_2200.t3 GNDA 0.047649f
C104 a_8570_6900.t13 GNDA 0.020006f
C105 a_8570_6900.n0 GNDA 0.319666f
C106 a_8570_6900.n1 GNDA 0.335179f
C107 a_8570_6900.t19 GNDA 0.020006f
C108 a_8570_6900.t16 GNDA 0.020006f
C109 a_8570_6900.n2 GNDA 0.040763f
C110 a_8570_6900.n3 GNDA 0.365375f
C111 a_8570_6900.t17 GNDA 0.020006f
C112 a_8570_6900.t12 GNDA 0.020006f
C113 a_8570_6900.n4 GNDA 0.040763f
C114 a_8570_6900.n5 GNDA 0.306668f
C115 a_8570_6900.n6 GNDA 0.319666f
C116 a_8570_6900.n7 GNDA 0.210468f
C117 a_8570_6900.t14 GNDA 0.020006f
C118 a_8570_6900.t10 GNDA 0.020006f
C119 a_8570_6900.n8 GNDA 0.040763f
C120 a_8570_6900.n9 GNDA 0.306668f
C121 a_8570_6900.n10 GNDA 0.218329f
C122 a_8570_6900.t11 GNDA 0.020006f
C123 a_8570_6900.t15 GNDA 0.020006f
C124 a_8570_6900.n11 GNDA 0.040763f
C125 a_8570_6900.n12 GNDA 0.233788f
C126 a_8570_6900.t9 GNDA 0.020006f
C127 a_8570_6900.t1 GNDA 0.020006f
C128 a_8570_6900.n13 GNDA 0.040763f
C129 a_8570_6900.n14 GNDA 0.191134f
C130 a_8570_6900.t4 GNDA 0.020006f
C131 a_8570_6900.t7 GNDA 0.020006f
C132 a_8570_6900.n15 GNDA 0.040763f
C133 a_8570_6900.n16 GNDA 0.300378f
C134 a_8570_6900.n17 GNDA 0.215758f
C135 a_8570_6900.n18 GNDA 0.206718f
C136 a_8570_6900.t3 GNDA 0.020006f
C137 a_8570_6900.t5 GNDA 0.020006f
C138 a_8570_6900.n19 GNDA 0.040763f
C139 a_8570_6900.n20 GNDA 0.300378f
C140 a_8570_6900.t8 GNDA 0.020006f
C141 a_8570_6900.t0 GNDA 0.020006f
C142 a_8570_6900.n21 GNDA 0.040763f
C143 a_8570_6900.n22 GNDA 0.279938f
C144 a_8570_6900.n23 GNDA 0.206718f
C145 a_8570_6900.n24 GNDA 0.122442f
C146 a_8570_6900.t2 GNDA 0.020006f
C147 a_8570_6900.t6 GNDA 0.020006f
C148 a_8570_6900.n25 GNDA 0.040763f
C149 a_8570_6900.n26 GNDA 0.279938f
C150 a_8570_6900.n27 GNDA 0.127024f
C151 a_8570_6900.n28 GNDA 0.208769f
C152 a_8570_6900.n29 GNDA 0.121174f
C153 a_8570_6900.n30 GNDA 0.18461f
C154 a_8570_6900.n31 GNDA 0.324795f
C155 a_8570_6900.n32 GNDA 0.306668f
C156 a_8570_6900.n33 GNDA 0.040763f
C157 a_8570_6900.t18 GNDA 0.020006f
C158 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t12 GNDA 0.026007f
C159 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t13 GNDA 0.026007f
C160 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n0 GNDA 0.09453f
C161 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t10 GNDA 0.026007f
C162 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t11 GNDA 0.026007f
C163 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n1 GNDA 0.078554f
C164 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n2 GNDA 1.53217f
C165 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t14 GNDA 0.324356f
C166 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n3 GNDA 0.090462f
C167 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n4 GNDA 0.155651f
C168 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t6 GNDA 0.078023f
C169 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t1 GNDA 0.078023f
C170 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n5 GNDA 0.166875f
C171 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n6 GNDA 0.521985f
C172 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t5 GNDA 0.078023f
C173 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t0 GNDA 0.078023f
C174 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n7 GNDA 0.166875f
C175 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n8 GNDA 0.507848f
C176 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n9 GNDA 0.155651f
C177 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n10 GNDA 0.090462f
C178 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t7 GNDA 0.078023f
C179 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t2 GNDA 0.078023f
C180 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n11 GNDA 0.166875f
C181 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n12 GNDA 0.507848f
C182 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n13 GNDA 0.090462f
C183 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t8 GNDA 0.078023f
C184 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t3 GNDA 0.078023f
C185 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n14 GNDA 0.166875f
C186 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n15 GNDA 0.507848f
C187 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n16 GNDA 0.155651f
C188 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t9 GNDA 0.078023f
C189 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.t4 GNDA 0.078023f
C190 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n17 GNDA 0.166875f
C191 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n18 GNDA 0.514916f
C192 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n19 GNDA 0.201702f
C193 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n20 GNDA 1.99814f
C194 two_stage_opamp_dummy_magic_21_0.V_CMFB_S2.n21 GNDA 2.34014f
C195 bgr_0.V_CMFB_S2 GNDA 0.013004f
C196 two_stage_opamp_dummy_magic_21_0.VD3.t17 GNDA 0.060837f
C197 two_stage_opamp_dummy_magic_21_0.VD3.t15 GNDA 0.060837f
C198 two_stage_opamp_dummy_magic_21_0.VD3.t11 GNDA 0.060837f
C199 two_stage_opamp_dummy_magic_21_0.VD3.n0 GNDA 0.154422f
C200 two_stage_opamp_dummy_magic_21_0.VD3.n1 GNDA 0.43135f
C201 two_stage_opamp_dummy_magic_21_0.VD3.t20 GNDA 0.106675f
C202 two_stage_opamp_dummy_magic_21_0.VD3.t25 GNDA 0.216405f
C203 two_stage_opamp_dummy_magic_21_0.VD3.n2 GNDA 0.065988f
C204 two_stage_opamp_dummy_magic_21_0.VD3.n3 GNDA 0.065988f
C205 two_stage_opamp_dummy_magic_21_0.VD3.t37 GNDA 0.060837f
C206 two_stage_opamp_dummy_magic_21_0.VD3.t33 GNDA 0.060837f
C207 two_stage_opamp_dummy_magic_21_0.VD3.n4 GNDA 0.124448f
C208 two_stage_opamp_dummy_magic_21_0.VD3.n5 GNDA 0.402926f
C209 two_stage_opamp_dummy_magic_21_0.VD3.n6 GNDA 0.112569f
C210 two_stage_opamp_dummy_magic_21_0.VD3.t31 GNDA 0.060837f
C211 two_stage_opamp_dummy_magic_21_0.VD3.t34 GNDA 0.060837f
C212 two_stage_opamp_dummy_magic_21_0.VD3.n7 GNDA 0.124448f
C213 two_stage_opamp_dummy_magic_21_0.VD3.n8 GNDA 0.391923f
C214 two_stage_opamp_dummy_magic_21_0.VD3.n9 GNDA 0.112569f
C215 two_stage_opamp_dummy_magic_21_0.VD3.t26 GNDA 0.060837f
C216 two_stage_opamp_dummy_magic_21_0.VD3.t28 GNDA 0.060837f
C217 two_stage_opamp_dummy_magic_21_0.VD3.n10 GNDA 0.124448f
C218 two_stage_opamp_dummy_magic_21_0.VD3.n11 GNDA 0.391923f
C219 two_stage_opamp_dummy_magic_21_0.VD3.n12 GNDA 0.065988f
C220 two_stage_opamp_dummy_magic_21_0.VD3.n13 GNDA 0.065988f
C221 two_stage_opamp_dummy_magic_21_0.VD3.t30 GNDA 0.060837f
C222 two_stage_opamp_dummy_magic_21_0.VD3.t29 GNDA 0.060837f
C223 two_stage_opamp_dummy_magic_21_0.VD3.n14 GNDA 0.124448f
C224 two_stage_opamp_dummy_magic_21_0.VD3.n15 GNDA 0.391923f
C225 two_stage_opamp_dummy_magic_21_0.VD3.n16 GNDA 0.065988f
C226 two_stage_opamp_dummy_magic_21_0.VD3.t32 GNDA 0.060837f
C227 two_stage_opamp_dummy_magic_21_0.VD3.t35 GNDA 0.060837f
C228 two_stage_opamp_dummy_magic_21_0.VD3.n17 GNDA 0.124448f
C229 two_stage_opamp_dummy_magic_21_0.VD3.n18 GNDA 0.391923f
C230 two_stage_opamp_dummy_magic_21_0.VD3.n19 GNDA 0.112569f
C231 two_stage_opamp_dummy_magic_21_0.VD3.t27 GNDA 0.060837f
C232 two_stage_opamp_dummy_magic_21_0.VD3.t36 GNDA 0.060837f
C233 two_stage_opamp_dummy_magic_21_0.VD3.n20 GNDA 0.124448f
C234 two_stage_opamp_dummy_magic_21_0.VD3.n21 GNDA 0.397425f
C235 two_stage_opamp_dummy_magic_21_0.VD3.n22 GNDA 0.257485f
C236 two_stage_opamp_dummy_magic_21_0.VD3.t1 GNDA 0.060837f
C237 two_stage_opamp_dummy_magic_21_0.VD3.t7 GNDA 0.060837f
C238 two_stage_opamp_dummy_magic_21_0.VD3.n23 GNDA 0.154422f
C239 two_stage_opamp_dummy_magic_21_0.VD3.n24 GNDA 0.43135f
C240 two_stage_opamp_dummy_magic_21_0.VD3.n25 GNDA 0.2193f
C241 two_stage_opamp_dummy_magic_21_0.VD3.t23 GNDA 0.106675f
C242 two_stage_opamp_dummy_magic_21_0.VD3.n26 GNDA 0.311214f
C243 two_stage_opamp_dummy_magic_21_0.VD3.n27 GNDA 0.627773f
C244 two_stage_opamp_dummy_magic_21_0.VD3.t24 GNDA 0.518568f
C245 two_stage_opamp_dummy_magic_21_0.VD3.t0 GNDA 0.406738f
C246 two_stage_opamp_dummy_magic_21_0.VD3.t6 GNDA 0.406738f
C247 two_stage_opamp_dummy_magic_21_0.VD3.t14 GNDA 0.406738f
C248 two_stage_opamp_dummy_magic_21_0.VD3.t10 GNDA 0.402972f
C249 two_stage_opamp_dummy_magic_21_0.VD3.t16 GNDA 0.399206f
C250 two_stage_opamp_dummy_magic_21_0.VD3.t18 GNDA 0.406738f
C251 two_stage_opamp_dummy_magic_21_0.VD3.t2 GNDA 0.406738f
C252 two_stage_opamp_dummy_magic_21_0.VD3.t8 GNDA 0.406738f
C253 two_stage_opamp_dummy_magic_21_0.VD3.t4 GNDA 0.406738f
C254 two_stage_opamp_dummy_magic_21_0.VD3.t12 GNDA 0.406738f
C255 two_stage_opamp_dummy_magic_21_0.VD3.t21 GNDA 0.518568f
C256 two_stage_opamp_dummy_magic_21_0.VD3.t22 GNDA 0.216405f
C257 two_stage_opamp_dummy_magic_21_0.VD3.n28 GNDA 0.627773f
C258 two_stage_opamp_dummy_magic_21_0.VD3.n29 GNDA 0.316969f
C259 two_stage_opamp_dummy_magic_21_0.VD3.t5 GNDA 0.060837f
C260 two_stage_opamp_dummy_magic_21_0.VD3.t13 GNDA 0.060837f
C261 two_stage_opamp_dummy_magic_21_0.VD3.n30 GNDA 0.154422f
C262 two_stage_opamp_dummy_magic_21_0.VD3.n31 GNDA 0.481799f
C263 two_stage_opamp_dummy_magic_21_0.VD3.t3 GNDA 0.060837f
C264 two_stage_opamp_dummy_magic_21_0.VD3.t9 GNDA 0.060837f
C265 two_stage_opamp_dummy_magic_21_0.VD3.n32 GNDA 0.154422f
C266 two_stage_opamp_dummy_magic_21_0.VD3.n33 GNDA 0.43135f
C267 two_stage_opamp_dummy_magic_21_0.VD3.n34 GNDA 0.43135f
C268 two_stage_opamp_dummy_magic_21_0.VD3.n35 GNDA 0.154422f
C269 two_stage_opamp_dummy_magic_21_0.VD3.t19 GNDA 0.060837f
C270 two_stage_opamp_dummy_magic_21_0.V_err_gate.n0 GNDA 0.27052f
C271 two_stage_opamp_dummy_magic_21_0.V_err_gate.n1 GNDA 0.27052f
C272 two_stage_opamp_dummy_magic_21_0.V_err_gate.n2 GNDA 0.246866f
C273 two_stage_opamp_dummy_magic_21_0.V_err_gate.n3 GNDA 0.343254f
C274 two_stage_opamp_dummy_magic_21_0.V_err_gate.n4 GNDA 0.177321f
C275 two_stage_opamp_dummy_magic_21_0.V_err_gate.n5 GNDA 0.20879f
C276 two_stage_opamp_dummy_magic_21_0.V_err_gate.t10 GNDA 0.032884f
C277 two_stage_opamp_dummy_magic_21_0.V_err_gate.t11 GNDA 0.032884f
C278 two_stage_opamp_dummy_magic_21_0.V_err_gate.n6 GNDA 0.500021f
C279 two_stage_opamp_dummy_magic_21_0.V_err_gate.t33 GNDA 0.013565f
C280 two_stage_opamp_dummy_magic_21_0.V_err_gate.t23 GNDA 0.013565f
C281 two_stage_opamp_dummy_magic_21_0.V_err_gate.t30 GNDA 0.013565f
C282 two_stage_opamp_dummy_magic_21_0.V_err_gate.t19 GNDA 0.013565f
C283 two_stage_opamp_dummy_magic_21_0.V_err_gate.t28 GNDA 0.013565f
C284 two_stage_opamp_dummy_magic_21_0.V_err_gate.t17 GNDA 0.013565f
C285 two_stage_opamp_dummy_magic_21_0.V_err_gate.t26 GNDA 0.013565f
C286 two_stage_opamp_dummy_magic_21_0.V_err_gate.t14 GNDA 0.013565f
C287 two_stage_opamp_dummy_magic_21_0.V_err_gate.t21 GNDA 0.013565f
C288 two_stage_opamp_dummy_magic_21_0.V_err_gate.t15 GNDA 0.013565f
C289 two_stage_opamp_dummy_magic_21_0.V_err_gate.t24 GNDA 0.02939f
C290 two_stage_opamp_dummy_magic_21_0.V_err_gate.n7 GNDA 0.045832f
C291 two_stage_opamp_dummy_magic_21_0.V_err_gate.n8 GNDA 0.035761f
C292 two_stage_opamp_dummy_magic_21_0.V_err_gate.n9 GNDA 0.035761f
C293 two_stage_opamp_dummy_magic_21_0.V_err_gate.n10 GNDA 0.035761f
C294 two_stage_opamp_dummy_magic_21_0.V_err_gate.n11 GNDA 0.035761f
C295 two_stage_opamp_dummy_magic_21_0.V_err_gate.n12 GNDA 0.035761f
C296 two_stage_opamp_dummy_magic_21_0.V_err_gate.n13 GNDA 0.035761f
C297 two_stage_opamp_dummy_magic_21_0.V_err_gate.n14 GNDA 0.035761f
C298 two_stage_opamp_dummy_magic_21_0.V_err_gate.n15 GNDA 0.035761f
C299 two_stage_opamp_dummy_magic_21_0.V_err_gate.n16 GNDA 0.029331f
C300 two_stage_opamp_dummy_magic_21_0.V_err_gate.t20 GNDA 0.013565f
C301 two_stage_opamp_dummy_magic_21_0.V_err_gate.t31 GNDA 0.013565f
C302 two_stage_opamp_dummy_magic_21_0.V_err_gate.t25 GNDA 0.013565f
C303 two_stage_opamp_dummy_magic_21_0.V_err_gate.t16 GNDA 0.013565f
C304 two_stage_opamp_dummy_magic_21_0.V_err_gate.t27 GNDA 0.013565f
C305 two_stage_opamp_dummy_magic_21_0.V_err_gate.t18 GNDA 0.013565f
C306 two_stage_opamp_dummy_magic_21_0.V_err_gate.t29 GNDA 0.013565f
C307 two_stage_opamp_dummy_magic_21_0.V_err_gate.t22 GNDA 0.013565f
C308 two_stage_opamp_dummy_magic_21_0.V_err_gate.t32 GNDA 0.033911f
C309 two_stage_opamp_dummy_magic_21_0.V_err_gate.n17 GNDA 0.070905f
C310 two_stage_opamp_dummy_magic_21_0.V_err_gate.n18 GNDA 0.035761f
C311 two_stage_opamp_dummy_magic_21_0.V_err_gate.n19 GNDA 0.035761f
C312 two_stage_opamp_dummy_magic_21_0.V_err_gate.n20 GNDA 0.035761f
C313 two_stage_opamp_dummy_magic_21_0.V_err_gate.n21 GNDA 0.035761f
C314 two_stage_opamp_dummy_magic_21_0.V_err_gate.n22 GNDA 0.035761f
C315 two_stage_opamp_dummy_magic_21_0.V_err_gate.n23 GNDA 0.035761f
C316 two_stage_opamp_dummy_magic_21_0.V_err_gate.n24 GNDA 0.029331f
C317 two_stage_opamp_dummy_magic_21_0.V_err_gate.n25 GNDA 0.045072f
C318 two_stage_opamp_dummy_magic_21_0.V_err_gate.t6 GNDA 0.016442f
C319 two_stage_opamp_dummy_magic_21_0.V_err_gate.t13 GNDA 0.016442f
C320 two_stage_opamp_dummy_magic_21_0.V_err_gate.n26 GNDA 0.033501f
C321 two_stage_opamp_dummy_magic_21_0.V_err_gate.t3 GNDA 0.016442f
C322 two_stage_opamp_dummy_magic_21_0.V_err_gate.t2 GNDA 0.016442f
C323 two_stage_opamp_dummy_magic_21_0.V_err_gate.n27 GNDA 0.033501f
C324 two_stage_opamp_dummy_magic_21_0.V_err_gate.n28 GNDA 0.230067f
C325 two_stage_opamp_dummy_magic_21_0.V_err_gate.t5 GNDA 0.016442f
C326 two_stage_opamp_dummy_magic_21_0.V_err_gate.t4 GNDA 0.016442f
C327 two_stage_opamp_dummy_magic_21_0.V_err_gate.n29 GNDA 0.033501f
C328 two_stage_opamp_dummy_magic_21_0.V_err_gate.n30 GNDA 0.230067f
C329 two_stage_opamp_dummy_magic_21_0.V_err_gate.t0 GNDA 0.016442f
C330 two_stage_opamp_dummy_magic_21_0.V_err_gate.t1 GNDA 0.016442f
C331 two_stage_opamp_dummy_magic_21_0.V_err_gate.n31 GNDA 0.033501f
C332 two_stage_opamp_dummy_magic_21_0.V_err_gate.n32 GNDA 0.230067f
C333 two_stage_opamp_dummy_magic_21_0.V_err_gate.t8 GNDA 0.016442f
C334 two_stage_opamp_dummy_magic_21_0.V_err_gate.t7 GNDA 0.016442f
C335 two_stage_opamp_dummy_magic_21_0.V_err_gate.n33 GNDA 0.033501f
C336 two_stage_opamp_dummy_magic_21_0.V_err_gate.n34 GNDA 0.230067f
C337 two_stage_opamp_dummy_magic_21_0.V_err_gate.t12 GNDA 0.016442f
C338 two_stage_opamp_dummy_magic_21_0.V_err_gate.t9 GNDA 0.016442f
C339 two_stage_opamp_dummy_magic_21_0.V_err_gate.n35 GNDA 0.033501f
C340 two_stage_opamp_dummy_magic_21_0.V_err_gate.n36 GNDA 0.238415f
C341 bgr_0.START_UP.t4 GNDA 1.06745f
C342 bgr_0.START_UP.t5 GNDA 0.02806f
C343 bgr_0.START_UP.n0 GNDA 0.714928f
C344 bgr_0.START_UP.t0 GNDA 0.026778f
C345 bgr_0.START_UP.t2 GNDA 0.026778f
C346 bgr_0.START_UP.n1 GNDA 0.097147f
C347 bgr_0.START_UP.t1 GNDA 0.026778f
C348 bgr_0.START_UP.t3 GNDA 0.026778f
C349 bgr_0.START_UP.n2 GNDA 0.08937f
C350 bgr_0.START_UP.n3 GNDA 0.462855f
C351 bgr_0.START_UP.t7 GNDA 0.010062f
C352 bgr_0.START_UP.t6 GNDA 0.010062f
C353 bgr_0.START_UP.n4 GNDA 0.028407f
C354 bgr_0.START_UP.n5 GNDA 0.260836f
C355 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t14 GNDA 0.026498f
C356 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t12 GNDA 0.026498f
C357 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n0 GNDA 0.096311f
C358 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t13 GNDA 0.026498f
C359 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t11 GNDA 0.026498f
C360 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n1 GNDA 0.080034f
C361 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n2 GNDA 1.56103f
C362 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t0 GNDA 0.329048f
C363 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n3 GNDA 0.092167f
C364 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n4 GNDA 0.158583f
C365 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t4 GNDA 0.079493f
C366 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t10 GNDA 0.079493f
C367 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n5 GNDA 0.170019f
C368 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n6 GNDA 0.531819f
C369 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t3 GNDA 0.079493f
C370 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t9 GNDA 0.079493f
C371 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n7 GNDA 0.170019f
C372 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n8 GNDA 0.517415f
C373 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n9 GNDA 0.158583f
C374 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n10 GNDA 0.092167f
C375 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t7 GNDA 0.079493f
C376 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t2 GNDA 0.079493f
C377 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n11 GNDA 0.170019f
C378 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n12 GNDA 0.517415f
C379 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n13 GNDA 0.092167f
C380 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t6 GNDA 0.079493f
C381 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t1 GNDA 0.079493f
C382 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n14 GNDA 0.170019f
C383 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n15 GNDA 0.517415f
C384 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n16 GNDA 0.158583f
C385 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t5 GNDA 0.079493f
C386 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.t8 GNDA 0.079493f
C387 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n17 GNDA 0.170019f
C388 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n18 GNDA 0.524617f
C389 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n19 GNDA 0.207431f
C390 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n20 GNDA 2.0121f
C391 two_stage_opamp_dummy_magic_21_0.V_CMFB_S4.n21 GNDA 2.38885f
C392 bgr_0.V_CMFB_S4 GNDA 0.013249f
C393 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t15 GNDA 0.014602f
C394 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t2 GNDA 0.014602f
C395 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n0 GNDA 0.036602f
C396 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t0 GNDA 0.014602f
C397 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t3 GNDA 0.014602f
C398 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n1 GNDA 0.036408f
C399 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n2 GNDA 0.323597f
C400 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t1 GNDA 0.014602f
C401 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t14 GNDA 0.014602f
C402 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n3 GNDA 0.029204f
C403 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n4 GNDA 0.054309f
C404 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t16 GNDA 0.187697f
C405 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n5 GNDA 0.046127f
C406 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n6 GNDA 0.081589f
C407 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t11 GNDA 0.029204f
C408 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t6 GNDA 0.029204f
C409 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n7 GNDA 0.059709f
C410 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n8 GNDA 0.200562f
C411 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t10 GNDA 0.029204f
C412 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t5 GNDA 0.029204f
C413 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n9 GNDA 0.059709f
C414 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n10 GNDA 0.193142f
C415 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n11 GNDA 0.078428f
C416 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n12 GNDA 0.046127f
C417 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t12 GNDA 0.029204f
C418 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t7 GNDA 0.029204f
C419 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n13 GNDA 0.059709f
C420 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n14 GNDA 0.193142f
C421 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n15 GNDA 0.047813f
C422 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t13 GNDA 0.029204f
C423 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t8 GNDA 0.029204f
C424 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n16 GNDA 0.059709f
C425 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n17 GNDA 0.193142f
C426 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n18 GNDA 0.081589f
C427 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t4 GNDA 0.029204f
C428 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.t9 GNDA 0.029204f
C429 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n19 GNDA 0.059709f
C430 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n20 GNDA 0.196958f
C431 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n21 GNDA 0.118026f
C432 two_stage_opamp_dummy_magic_21_0.V_CMFB_S1.n22 GNDA 1.33686f
C433 bgr_0.V_CMFB_S1 GNDA 0.840486f
C434 bgr_0.Vin-.n0 GNDA 0.069747f
C435 bgr_0.Vin-.n1 GNDA 0.078367f
C436 bgr_0.Vin-.n2 GNDA 0.113033f
C437 bgr_0.Vin-.t6 GNDA 0.261601f
C438 bgr_0.Vin-.t3 GNDA 0.027101f
C439 bgr_0.Vin-.t1 GNDA 0.027101f
C440 bgr_0.Vin-.n3 GNDA 0.094346f
C441 bgr_0.Vin-.t0 GNDA 0.027101f
C442 bgr_0.Vin-.t2 GNDA 0.027101f
C443 bgr_0.Vin-.n4 GNDA 0.090091f
C444 bgr_0.Vin-.n5 GNDA 0.386489f
C445 bgr_0.Vin-.n6 GNDA 0.027681f
C446 bgr_0.Vin-.n7 GNDA 0.366254f
C447 bgr_0.Vin-.t12 GNDA 0.022346f
C448 bgr_0.Vin-.n8 GNDA 0.026209f
C449 bgr_0.Vin-.n9 GNDA 0.021455f
C450 bgr_0.Vin-.n10 GNDA 0.021455f
C451 bgr_0.Vin-.n11 GNDA 0.036491f
C452 bgr_0.Vin-.n12 GNDA 0.497932f
C453 bgr_0.Vin-.t7 GNDA 0.117924f
C454 bgr_0.Vin-.n13 GNDA 0.65583f
C455 bgr_0.Vin-.n14 GNDA 1.073f
C456 bgr_0.Vin-.n15 GNDA 0.471409f
C457 bgr_0.Vin-.n16 GNDA 0.07053f
C458 bgr_0.Vin-.n17 GNDA 0.119504f
C459 bgr_0.Vin-.n18 GNDA 0.069875f
C460 bgr_0.Vin-.n19 GNDA 0.138215f
C461 bgr_0.Vin-.n20 GNDA 0.138215f
C462 bgr_0.Vin-.n21 GNDA -0.269519f
C463 bgr_0.Vin-.n22 GNDA 0.445457f
C464 bgr_0.Vin-.n23 GNDA 0.213551f
C465 bgr_0.Vin-.n24 GNDA 0.403461f
C466 bgr_0.Vin-.n25 GNDA 0.0384f
C467 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.040751f
C468 bgr_0.V_mir2.t7 GNDA 0.019293f
C469 bgr_0.V_mir2.n0 GNDA 0.025223f
C470 bgr_0.V_mir2.t14 GNDA 0.041163f
C471 bgr_0.V_mir2.n1 GNDA 0.027381f
C472 bgr_0.V_mir2.n2 GNDA 0.451535f
C473 bgr_0.V_mir2.n3 GNDA 0.146338f
C474 bgr_0.V_mir2.t4 GNDA 0.023151f
C475 bgr_0.V_mir2.t17 GNDA 0.023151f
C476 bgr_0.V_mir2.t20 GNDA 0.037369f
C477 bgr_0.V_mir2.n4 GNDA 0.041731f
C478 bgr_0.V_mir2.n5 GNDA 0.028507f
C479 bgr_0.V_mir2.t0 GNDA 0.02939f
C480 bgr_0.V_mir2.n6 GNDA 0.044354f
C481 bgr_0.V_mir2.t5 GNDA 0.019293f
C482 bgr_0.V_mir2.t1 GNDA 0.019293f
C483 bgr_0.V_mir2.n7 GNDA 0.044166f
C484 bgr_0.V_mir2.n8 GNDA 0.109943f
C485 bgr_0.V_mir2.t2 GNDA 0.023151f
C486 bgr_0.V_mir2.t18 GNDA 0.023151f
C487 bgr_0.V_mir2.t22 GNDA 0.037369f
C488 bgr_0.V_mir2.n9 GNDA 0.041731f
C489 bgr_0.V_mir2.n10 GNDA 0.028507f
C490 bgr_0.V_mir2.t8 GNDA 0.02939f
C491 bgr_0.V_mir2.n11 GNDA 0.044354f
C492 bgr_0.V_mir2.t3 GNDA 0.019293f
C493 bgr_0.V_mir2.t9 GNDA 0.019293f
C494 bgr_0.V_mir2.n12 GNDA 0.044166f
C495 bgr_0.V_mir2.n13 GNDA 0.111042f
C496 bgr_0.V_mir2.n14 GNDA 0.381359f
C497 bgr_0.V_mir2.n15 GNDA 0.051125f
C498 bgr_0.V_mir2.t6 GNDA 0.023151f
C499 bgr_0.V_mir2.t19 GNDA 0.023151f
C500 bgr_0.V_mir2.t21 GNDA 0.037369f
C501 bgr_0.V_mir2.n16 GNDA 0.041731f
C502 bgr_0.V_mir2.n17 GNDA 0.028507f
C503 bgr_0.V_mir2.t10 GNDA 0.02939f
C504 bgr_0.V_mir2.n18 GNDA 0.044354f
C505 bgr_0.V_mir2.n19 GNDA 0.085095f
C506 bgr_0.V_mir2.n20 GNDA 0.044166f
C507 bgr_0.V_mir2.t11 GNDA 0.019293f
C508 bgr_0.cap_res1.t11 GNDA 0.331712f
C509 bgr_0.cap_res1.t18 GNDA 0.349187f
C510 bgr_0.cap_res1.t15 GNDA 0.350452f
C511 bgr_0.cap_res1.t4 GNDA 0.331712f
C512 bgr_0.cap_res1.t14 GNDA 0.349187f
C513 bgr_0.cap_res1.t8 GNDA 0.350452f
C514 bgr_0.cap_res1.t10 GNDA 0.331712f
C515 bgr_0.cap_res1.t17 GNDA 0.349187f
C516 bgr_0.cap_res1.t13 GNDA 0.350452f
C517 bgr_0.cap_res1.t3 GNDA 0.331712f
C518 bgr_0.cap_res1.t12 GNDA 0.349187f
C519 bgr_0.cap_res1.t6 GNDA 0.350452f
C520 bgr_0.cap_res1.t19 GNDA 0.331712f
C521 bgr_0.cap_res1.t5 GNDA 0.349187f
C522 bgr_0.cap_res1.t0 GNDA 0.350452f
C523 bgr_0.cap_res1.n0 GNDA 0.23406f
C524 bgr_0.cap_res1.t16 GNDA 0.186395f
C525 bgr_0.cap_res1.n1 GNDA 0.253961f
C526 bgr_0.cap_res1.t1 GNDA 0.186395f
C527 bgr_0.cap_res1.n2 GNDA 0.253961f
C528 bgr_0.cap_res1.t7 GNDA 0.186395f
C529 bgr_0.cap_res1.n3 GNDA 0.253961f
C530 bgr_0.cap_res1.t2 GNDA 0.186395f
C531 bgr_0.cap_res1.n4 GNDA 0.253961f
C532 bgr_0.cap_res1.t9 GNDA 0.363549f
C533 bgr_0.cap_res1.t20 GNDA 0.08421f
C534 two_stage_opamp_dummy_magic_21_0.cap_res_X.t89 GNDA 0.344881f
C535 two_stage_opamp_dummy_magic_21_0.cap_res_X.t126 GNDA 0.346131f
C536 two_stage_opamp_dummy_magic_21_0.cap_res_X.t48 GNDA 0.344881f
C537 two_stage_opamp_dummy_magic_21_0.cap_res_X.t87 GNDA 0.347585f
C538 two_stage_opamp_dummy_magic_21_0.cap_res_X.t66 GNDA 0.378048f
C539 two_stage_opamp_dummy_magic_21_0.cap_res_X.t129 GNDA 0.344881f
C540 two_stage_opamp_dummy_magic_21_0.cap_res_X.t26 GNDA 0.346131f
C541 two_stage_opamp_dummy_magic_21_0.cap_res_X.t80 GNDA 0.344881f
C542 two_stage_opamp_dummy_magic_21_0.cap_res_X.t41 GNDA 0.346131f
C543 two_stage_opamp_dummy_magic_21_0.cap_res_X.t94 GNDA 0.344881f
C544 two_stage_opamp_dummy_magic_21_0.cap_res_X.t133 GNDA 0.346131f
C545 two_stage_opamp_dummy_magic_21_0.cap_res_X.t44 GNDA 0.344881f
C546 two_stage_opamp_dummy_magic_21_0.cap_res_X.t8 GNDA 0.346131f
C547 two_stage_opamp_dummy_magic_21_0.cap_res_X.t42 GNDA 0.344881f
C548 two_stage_opamp_dummy_magic_21_0.cap_res_X.t78 GNDA 0.346131f
C549 two_stage_opamp_dummy_magic_21_0.cap_res_X.t57 GNDA 0.344881f
C550 two_stage_opamp_dummy_magic_21_0.cap_res_X.t24 GNDA 0.346131f
C551 two_stage_opamp_dummy_magic_21_0.cap_res_X.t82 GNDA 0.344881f
C552 two_stage_opamp_dummy_magic_21_0.cap_res_X.t117 GNDA 0.346131f
C553 two_stage_opamp_dummy_magic_21_0.cap_res_X.t101 GNDA 0.344881f
C554 two_stage_opamp_dummy_magic_21_0.cap_res_X.t64 GNDA 0.346131f
C555 two_stage_opamp_dummy_magic_21_0.cap_res_X.t47 GNDA 0.344881f
C556 two_stage_opamp_dummy_magic_21_0.cap_res_X.t85 GNDA 0.346131f
C557 two_stage_opamp_dummy_magic_21_0.cap_res_X.t65 GNDA 0.344881f
C558 two_stage_opamp_dummy_magic_21_0.cap_res_X.t30 GNDA 0.346131f
C559 two_stage_opamp_dummy_magic_21_0.cap_res_X.t88 GNDA 0.344881f
C560 two_stage_opamp_dummy_magic_21_0.cap_res_X.t123 GNDA 0.346131f
C561 two_stage_opamp_dummy_magic_21_0.cap_res_X.t104 GNDA 0.344881f
C562 two_stage_opamp_dummy_magic_21_0.cap_res_X.t68 GNDA 0.346131f
C563 two_stage_opamp_dummy_magic_21_0.cap_res_X.t127 GNDA 0.344881f
C564 two_stage_opamp_dummy_magic_21_0.cap_res_X.t21 GNDA 0.346131f
C565 two_stage_opamp_dummy_magic_21_0.cap_res_X.t3 GNDA 0.344881f
C566 two_stage_opamp_dummy_magic_21_0.cap_res_X.t108 GNDA 0.346131f
C567 two_stage_opamp_dummy_magic_21_0.cap_res_X.t93 GNDA 0.344881f
C568 two_stage_opamp_dummy_magic_21_0.cap_res_X.t128 GNDA 0.346131f
C569 two_stage_opamp_dummy_magic_21_0.cap_res_X.t110 GNDA 0.344881f
C570 two_stage_opamp_dummy_magic_21_0.cap_res_X.t75 GNDA 0.346131f
C571 two_stage_opamp_dummy_magic_21_0.cap_res_X.t134 GNDA 0.344881f
C572 two_stage_opamp_dummy_magic_21_0.cap_res_X.t27 GNDA 0.346131f
C573 two_stage_opamp_dummy_magic_21_0.cap_res_X.t10 GNDA 0.344881f
C574 two_stage_opamp_dummy_magic_21_0.cap_res_X.t116 GNDA 0.346131f
C575 two_stage_opamp_dummy_magic_21_0.cap_res_X.t33 GNDA 0.344881f
C576 two_stage_opamp_dummy_magic_21_0.cap_res_X.t67 GNDA 0.346131f
C577 two_stage_opamp_dummy_magic_21_0.cap_res_X.t49 GNDA 0.344881f
C578 two_stage_opamp_dummy_magic_21_0.cap_res_X.t15 GNDA 0.346131f
C579 two_stage_opamp_dummy_magic_21_0.cap_res_X.t72 GNDA 0.344881f
C580 two_stage_opamp_dummy_magic_21_0.cap_res_X.t107 GNDA 0.346131f
C581 two_stage_opamp_dummy_magic_21_0.cap_res_X.t90 GNDA 0.344881f
C582 two_stage_opamp_dummy_magic_21_0.cap_res_X.t53 GNDA 0.346131f
C583 two_stage_opamp_dummy_magic_21_0.cap_res_X.t35 GNDA 0.344881f
C584 two_stage_opamp_dummy_magic_21_0.cap_res_X.t73 GNDA 0.346131f
C585 two_stage_opamp_dummy_magic_21_0.cap_res_X.t52 GNDA 0.344881f
C586 two_stage_opamp_dummy_magic_21_0.cap_res_X.t19 GNDA 0.346131f
C587 two_stage_opamp_dummy_magic_21_0.cap_res_X.t77 GNDA 0.344881f
C588 two_stage_opamp_dummy_magic_21_0.cap_res_X.t115 GNDA 0.346131f
C589 two_stage_opamp_dummy_magic_21_0.cap_res_X.t96 GNDA 0.344881f
C590 two_stage_opamp_dummy_magic_21_0.cap_res_X.t56 GNDA 0.346131f
C591 two_stage_opamp_dummy_magic_21_0.cap_res_X.t119 GNDA 0.344881f
C592 two_stage_opamp_dummy_magic_21_0.cap_res_X.t14 GNDA 0.346131f
C593 two_stage_opamp_dummy_magic_21_0.cap_res_X.t136 GNDA 0.344881f
C594 two_stage_opamp_dummy_magic_21_0.cap_res_X.t99 GNDA 0.346131f
C595 two_stage_opamp_dummy_magic_21_0.cap_res_X.t84 GNDA 0.344881f
C596 two_stage_opamp_dummy_magic_21_0.cap_res_X.t118 GNDA 0.346131f
C597 two_stage_opamp_dummy_magic_21_0.cap_res_X.t83 GNDA 0.344881f
C598 two_stage_opamp_dummy_magic_21_0.cap_res_X.t7 GNDA 0.361791f
C599 two_stage_opamp_dummy_magic_21_0.cap_res_X.t40 GNDA 0.344881f
C600 two_stage_opamp_dummy_magic_21_0.cap_res_X.t98 GNDA 0.185242f
C601 two_stage_opamp_dummy_magic_21_0.cap_res_X.n0 GNDA 0.198255f
C602 two_stage_opamp_dummy_magic_21_0.cap_res_X.t92 GNDA 0.344881f
C603 two_stage_opamp_dummy_magic_21_0.cap_res_X.t59 GNDA 0.185242f
C604 two_stage_opamp_dummy_magic_21_0.cap_res_X.n1 GNDA 0.196656f
C605 two_stage_opamp_dummy_magic_21_0.cap_res_X.t2 GNDA 0.344881f
C606 two_stage_opamp_dummy_magic_21_0.cap_res_X.t25 GNDA 0.185242f
C607 two_stage_opamp_dummy_magic_21_0.cap_res_X.n2 GNDA 0.196656f
C608 two_stage_opamp_dummy_magic_21_0.cap_res_X.t50 GNDA 0.344881f
C609 two_stage_opamp_dummy_magic_21_0.cap_res_X.t132 GNDA 0.185242f
C610 two_stage_opamp_dummy_magic_21_0.cap_res_X.n3 GNDA 0.196656f
C611 two_stage_opamp_dummy_magic_21_0.cap_res_X.t13 GNDA 0.344881f
C612 two_stage_opamp_dummy_magic_21_0.cap_res_X.t81 GNDA 0.185242f
C613 two_stage_opamp_dummy_magic_21_0.cap_res_X.n4 GNDA 0.196656f
C614 two_stage_opamp_dummy_magic_21_0.cap_res_X.t60 GNDA 0.344881f
C615 two_stage_opamp_dummy_magic_21_0.cap_res_X.t43 GNDA 0.185242f
C616 two_stage_opamp_dummy_magic_21_0.cap_res_X.n5 GNDA 0.196656f
C617 two_stage_opamp_dummy_magic_21_0.cap_res_X.t114 GNDA 0.344881f
C618 two_stage_opamp_dummy_magic_21_0.cap_res_X.t12 GNDA 0.185242f
C619 two_stage_opamp_dummy_magic_21_0.cap_res_X.n6 GNDA 0.196656f
C620 two_stage_opamp_dummy_magic_21_0.cap_res_X.t70 GNDA 0.344881f
C621 two_stage_opamp_dummy_magic_21_0.cap_res_X.t102 GNDA 0.185242f
C622 two_stage_opamp_dummy_magic_21_0.cap_res_X.n7 GNDA 0.196656f
C623 two_stage_opamp_dummy_magic_21_0.cap_res_X.t122 GNDA 0.344881f
C624 two_stage_opamp_dummy_magic_21_0.cap_res_X.t62 GNDA 0.185242f
C625 two_stage_opamp_dummy_magic_21_0.cap_res_X.n8 GNDA 0.196656f
C626 two_stage_opamp_dummy_magic_21_0.cap_res_X.t39 GNDA 0.344881f
C627 two_stage_opamp_dummy_magic_21_0.cap_res_X.t131 GNDA 0.346131f
C628 two_stage_opamp_dummy_magic_21_0.cap_res_X.t32 GNDA 0.166734f
C629 two_stage_opamp_dummy_magic_21_0.cap_res_X.n9 GNDA 0.215061f
C630 two_stage_opamp_dummy_magic_21_0.cap_res_X.t29 GNDA 0.184096f
C631 two_stage_opamp_dummy_magic_21_0.cap_res_X.n10 GNDA 0.23357f
C632 two_stage_opamp_dummy_magic_21_0.cap_res_X.t63 GNDA 0.184096f
C633 two_stage_opamp_dummy_magic_21_0.cap_res_X.n11 GNDA 0.250829f
C634 two_stage_opamp_dummy_magic_21_0.cap_res_X.t23 GNDA 0.184096f
C635 two_stage_opamp_dummy_magic_21_0.cap_res_X.n12 GNDA 0.250829f
C636 two_stage_opamp_dummy_magic_21_0.cap_res_X.t125 GNDA 0.184096f
C637 two_stage_opamp_dummy_magic_21_0.cap_res_X.n13 GNDA 0.250829f
C638 two_stage_opamp_dummy_magic_21_0.cap_res_X.t18 GNDA 0.184096f
C639 two_stage_opamp_dummy_magic_21_0.cap_res_X.n14 GNDA 0.250829f
C640 two_stage_opamp_dummy_magic_21_0.cap_res_X.t121 GNDA 0.184096f
C641 two_stage_opamp_dummy_magic_21_0.cap_res_X.n15 GNDA 0.250829f
C642 two_stage_opamp_dummy_magic_21_0.cap_res_X.t79 GNDA 0.184096f
C643 two_stage_opamp_dummy_magic_21_0.cap_res_X.n16 GNDA 0.250829f
C644 two_stage_opamp_dummy_magic_21_0.cap_res_X.t36 GNDA 0.184096f
C645 two_stage_opamp_dummy_magic_21_0.cap_res_X.n17 GNDA 0.250829f
C646 two_stage_opamp_dummy_magic_21_0.cap_res_X.t74 GNDA 0.184096f
C647 two_stage_opamp_dummy_magic_21_0.cap_res_X.n18 GNDA 0.250829f
C648 two_stage_opamp_dummy_magic_21_0.cap_res_X.t34 GNDA 0.184096f
C649 two_stage_opamp_dummy_magic_21_0.cap_res_X.n19 GNDA 0.250829f
C650 two_stage_opamp_dummy_magic_21_0.cap_res_X.t137 GNDA 0.184096f
C651 two_stage_opamp_dummy_magic_21_0.cap_res_X.n20 GNDA 0.250829f
C652 two_stage_opamp_dummy_magic_21_0.cap_res_X.t28 GNDA 0.184096f
C653 two_stage_opamp_dummy_magic_21_0.cap_res_X.n21 GNDA 0.250829f
C654 two_stage_opamp_dummy_magic_21_0.cap_res_X.t130 GNDA 0.184096f
C655 two_stage_opamp_dummy_magic_21_0.cap_res_X.n22 GNDA 0.250829f
C656 two_stage_opamp_dummy_magic_21_0.cap_res_X.t109 GNDA 0.184096f
C657 two_stage_opamp_dummy_magic_21_0.cap_res_X.n23 GNDA 0.250829f
C658 two_stage_opamp_dummy_magic_21_0.cap_res_X.t4 GNDA 0.184096f
C659 two_stage_opamp_dummy_magic_21_0.cap_res_X.n24 GNDA 0.250829f
C660 two_stage_opamp_dummy_magic_21_0.cap_res_X.t105 GNDA 0.184096f
C661 two_stage_opamp_dummy_magic_21_0.cap_res_X.n25 GNDA 0.23357f
C662 two_stage_opamp_dummy_magic_21_0.cap_res_X.t103 GNDA 0.343735f
C663 two_stage_opamp_dummy_magic_21_0.cap_res_X.t1 GNDA 0.166734f
C664 two_stage_opamp_dummy_magic_21_0.cap_res_X.n26 GNDA 0.216311f
C665 two_stage_opamp_dummy_magic_21_0.cap_res_X.t0 GNDA 0.343735f
C666 two_stage_opamp_dummy_magic_21_0.cap_res_X.t37 GNDA 0.166734f
C667 two_stage_opamp_dummy_magic_21_0.cap_res_X.n27 GNDA 0.216311f
C668 two_stage_opamp_dummy_magic_21_0.cap_res_X.t120 GNDA 0.343735f
C669 two_stage_opamp_dummy_magic_21_0.cap_res_X.t112 GNDA 0.344881f
C670 two_stage_opamp_dummy_magic_21_0.cap_res_X.t20 GNDA 0.36339f
C671 two_stage_opamp_dummy_magic_21_0.cap_res_X.t55 GNDA 0.36339f
C672 two_stage_opamp_dummy_magic_21_0.cap_res_X.t17 GNDA 0.185242f
C673 two_stage_opamp_dummy_magic_21_0.cap_res_X.n28 GNDA 0.216311f
C674 two_stage_opamp_dummy_magic_21_0.cap_res_X.t124 GNDA 0.343735f
C675 two_stage_opamp_dummy_magic_21_0.cap_res_X.t61 GNDA 0.344881f
C676 two_stage_opamp_dummy_magic_21_0.cap_res_X.t22 GNDA 0.185242f
C677 two_stage_opamp_dummy_magic_21_0.cap_res_X.n29 GNDA 0.197803f
C678 two_stage_opamp_dummy_magic_21_0.cap_res_X.t6 GNDA 0.343735f
C679 two_stage_opamp_dummy_magic_21_0.cap_res_X.t86 GNDA 0.344881f
C680 two_stage_opamp_dummy_magic_21_0.cap_res_X.t45 GNDA 0.185242f
C681 two_stage_opamp_dummy_magic_21_0.cap_res_X.n30 GNDA 0.216311f
C682 two_stage_opamp_dummy_magic_21_0.cap_res_X.t106 GNDA 0.343735f
C683 two_stage_opamp_dummy_magic_21_0.cap_res_X.t46 GNDA 0.344881f
C684 two_stage_opamp_dummy_magic_21_0.cap_res_X.t9 GNDA 0.185242f
C685 two_stage_opamp_dummy_magic_21_0.cap_res_X.n31 GNDA 0.216311f
C686 two_stage_opamp_dummy_magic_21_0.cap_res_X.t69 GNDA 0.343735f
C687 two_stage_opamp_dummy_magic_21_0.cap_res_X.t11 GNDA 0.344881f
C688 two_stage_opamp_dummy_magic_21_0.cap_res_X.t111 GNDA 0.185242f
C689 two_stage_opamp_dummy_magic_21_0.cap_res_X.n32 GNDA 0.216311f
C690 two_stage_opamp_dummy_magic_21_0.cap_res_X.t31 GNDA 0.343735f
C691 two_stage_opamp_dummy_magic_21_0.cap_res_X.t91 GNDA 0.344881f
C692 two_stage_opamp_dummy_magic_21_0.cap_res_X.t76 GNDA 0.36339f
C693 two_stage_opamp_dummy_magic_21_0.cap_res_X.t113 GNDA 0.36339f
C694 two_stage_opamp_dummy_magic_21_0.cap_res_X.t71 GNDA 0.185242f
C695 two_stage_opamp_dummy_magic_21_0.cap_res_X.n33 GNDA 0.216311f
C696 two_stage_opamp_dummy_magic_21_0.cap_res_X.t51 GNDA 0.343735f
C697 two_stage_opamp_dummy_magic_21_0.cap_res_X.t38 GNDA 0.344881f
C698 two_stage_opamp_dummy_magic_21_0.cap_res_X.t100 GNDA 0.36339f
C699 two_stage_opamp_dummy_magic_21_0.cap_res_X.t135 GNDA 0.36339f
C700 two_stage_opamp_dummy_magic_21_0.cap_res_X.t95 GNDA 0.185242f
C701 two_stage_opamp_dummy_magic_21_0.cap_res_X.n34 GNDA 0.216311f
C702 two_stage_opamp_dummy_magic_21_0.cap_res_X.t16 GNDA 0.343735f
C703 two_stage_opamp_dummy_magic_21_0.cap_res_X.n35 GNDA 0.216311f
C704 two_stage_opamp_dummy_magic_21_0.cap_res_X.t54 GNDA 0.185242f
C705 two_stage_opamp_dummy_magic_21_0.cap_res_X.t97 GNDA 0.36339f
C706 two_stage_opamp_dummy_magic_21_0.cap_res_X.t58 GNDA 0.36339f
C707 two_stage_opamp_dummy_magic_21_0.cap_res_X.t5 GNDA 0.736617f
C708 two_stage_opamp_dummy_magic_21_0.cap_res_X.t138 GNDA 0.297532f
C709 bgr_0.PFET_GATE_10uA.t28 GNDA 0.020856f
C710 bgr_0.PFET_GATE_10uA.t20 GNDA 0.030831f
C711 bgr_0.PFET_GATE_10uA.n0 GNDA 0.033972f
C712 bgr_0.PFET_GATE_10uA.t15 GNDA 0.020856f
C713 bgr_0.PFET_GATE_10uA.t21 GNDA 0.030831f
C714 bgr_0.PFET_GATE_10uA.n1 GNDA 0.033972f
C715 bgr_0.PFET_GATE_10uA.n2 GNDA 0.040878f
C716 bgr_0.PFET_GATE_10uA.t19 GNDA 0.020856f
C717 bgr_0.PFET_GATE_10uA.t12 GNDA 0.030831f
C718 bgr_0.PFET_GATE_10uA.n3 GNDA 0.033972f
C719 bgr_0.PFET_GATE_10uA.t26 GNDA 0.020856f
C720 bgr_0.PFET_GATE_10uA.t13 GNDA 0.030831f
C721 bgr_0.PFET_GATE_10uA.n4 GNDA 0.033972f
C722 bgr_0.PFET_GATE_10uA.n5 GNDA 0.034081f
C723 bgr_0.PFET_GATE_10uA.t1 GNDA 0.312465f
C724 bgr_0.PFET_GATE_10uA.t4 GNDA 0.021391f
C725 bgr_0.PFET_GATE_10uA.t2 GNDA 0.021391f
C726 bgr_0.PFET_GATE_10uA.n6 GNDA 0.054673f
C727 bgr_0.PFET_GATE_10uA.t6 GNDA 0.021391f
C728 bgr_0.PFET_GATE_10uA.t8 GNDA 0.021391f
C729 bgr_0.PFET_GATE_10uA.n7 GNDA 0.05326f
C730 bgr_0.PFET_GATE_10uA.n8 GNDA 0.520952f
C731 bgr_0.PFET_GATE_10uA.t7 GNDA 0.021391f
C732 bgr_0.PFET_GATE_10uA.t9 GNDA 0.021391f
C733 bgr_0.PFET_GATE_10uA.n9 GNDA 0.05326f
C734 bgr_0.PFET_GATE_10uA.n10 GNDA 0.295408f
C735 bgr_0.PFET_GATE_10uA.n11 GNDA 0.603055f
C736 bgr_0.PFET_GATE_10uA.t3 GNDA 0.021391f
C737 bgr_0.PFET_GATE_10uA.t5 GNDA 0.021391f
C738 bgr_0.PFET_GATE_10uA.n12 GNDA 0.05159f
C739 bgr_0.PFET_GATE_10uA.n13 GNDA 0.275411f
C740 bgr_0.PFET_GATE_10uA.t0 GNDA 0.464967f
C741 bgr_0.PFET_GATE_10uA.t27 GNDA 0.024114f
C742 bgr_0.PFET_GATE_10uA.t14 GNDA 0.024114f
C743 bgr_0.PFET_GATE_10uA.n14 GNDA 0.069715f
C744 bgr_0.PFET_GATE_10uA.n15 GNDA 1.91969f
C745 bgr_0.PFET_GATE_10uA.n16 GNDA 0.771508f
C746 bgr_0.PFET_GATE_10uA.n17 GNDA 0.759224f
C747 bgr_0.PFET_GATE_10uA.t11 GNDA 0.020856f
C748 bgr_0.PFET_GATE_10uA.t25 GNDA 0.020856f
C749 bgr_0.PFET_GATE_10uA.t18 GNDA 0.020856f
C750 bgr_0.PFET_GATE_10uA.t10 GNDA 0.020856f
C751 bgr_0.PFET_GATE_10uA.t24 GNDA 0.020856f
C752 bgr_0.PFET_GATE_10uA.t17 GNDA 0.030831f
C753 bgr_0.PFET_GATE_10uA.n18 GNDA 0.038154f
C754 bgr_0.PFET_GATE_10uA.n19 GNDA 0.027273f
C755 bgr_0.PFET_GATE_10uA.n20 GNDA 0.027273f
C756 bgr_0.PFET_GATE_10uA.n21 GNDA 0.027273f
C757 bgr_0.PFET_GATE_10uA.n22 GNDA 0.023091f
C758 bgr_0.PFET_GATE_10uA.t16 GNDA 0.020856f
C759 bgr_0.PFET_GATE_10uA.t23 GNDA 0.020856f
C760 bgr_0.PFET_GATE_10uA.t22 GNDA 0.020856f
C761 bgr_0.PFET_GATE_10uA.t29 GNDA 0.030831f
C762 bgr_0.PFET_GATE_10uA.n23 GNDA 0.038154f
C763 bgr_0.PFET_GATE_10uA.n24 GNDA 0.027273f
C764 bgr_0.PFET_GATE_10uA.n25 GNDA 0.023091f
C765 bgr_0.PFET_GATE_10uA.n26 GNDA 0.031695f
C766 two_stage_opamp_dummy_magic_21_0.VD1.t15 GNDA 0.053331f
C767 two_stage_opamp_dummy_magic_21_0.VD1.n0 GNDA 0.119128f
C768 two_stage_opamp_dummy_magic_21_0.VD1.n1 GNDA 0.099935f
C769 two_stage_opamp_dummy_magic_21_0.VD1.n2 GNDA 0.205342f
C770 two_stage_opamp_dummy_magic_21_0.VD1.t9 GNDA 0.053331f
C771 two_stage_opamp_dummy_magic_21_0.VD1.t7 GNDA 0.053331f
C772 two_stage_opamp_dummy_magic_21_0.VD1.n3 GNDA 0.116042f
C773 two_stage_opamp_dummy_magic_21_0.VD1.n4 GNDA 0.465721f
C774 two_stage_opamp_dummy_magic_21_0.VD1.n5 GNDA 0.205342f
C775 two_stage_opamp_dummy_magic_21_0.VD1.t11 GNDA 0.053331f
C776 two_stage_opamp_dummy_magic_21_0.VD1.t5 GNDA 0.053331f
C777 two_stage_opamp_dummy_magic_21_0.VD1.n6 GNDA 0.116042f
C778 two_stage_opamp_dummy_magic_21_0.VD1.n7 GNDA 0.447102f
C779 two_stage_opamp_dummy_magic_21_0.VD1.n8 GNDA 0.192793f
C780 two_stage_opamp_dummy_magic_21_0.VD1.t0 GNDA 0.053331f
C781 two_stage_opamp_dummy_magic_21_0.VD1.t2 GNDA 0.053331f
C782 two_stage_opamp_dummy_magic_21_0.VD1.n9 GNDA 0.116042f
C783 two_stage_opamp_dummy_magic_21_0.VD1.n10 GNDA 0.447102f
C784 two_stage_opamp_dummy_magic_21_0.VD1.n11 GNDA 0.113419f
C785 two_stage_opamp_dummy_magic_21_0.VD1.t10 GNDA 0.053331f
C786 two_stage_opamp_dummy_magic_21_0.VD1.t8 GNDA 0.053331f
C787 two_stage_opamp_dummy_magic_21_0.VD1.n12 GNDA 0.116042f
C788 two_stage_opamp_dummy_magic_21_0.VD1.n13 GNDA 0.465721f
C789 two_stage_opamp_dummy_magic_21_0.VD1.t1 GNDA 0.053331f
C790 two_stage_opamp_dummy_magic_21_0.VD1.t6 GNDA 0.053331f
C791 two_stage_opamp_dummy_magic_21_0.VD1.n14 GNDA 0.116042f
C792 two_stage_opamp_dummy_magic_21_0.VD1.n15 GNDA 0.447102f
C793 two_stage_opamp_dummy_magic_21_0.VD1.n16 GNDA 0.192793f
C794 two_stage_opamp_dummy_magic_21_0.VD1.n17 GNDA 0.113419f
C795 two_stage_opamp_dummy_magic_21_0.VD1.t4 GNDA 0.053331f
C796 two_stage_opamp_dummy_magic_21_0.VD1.t3 GNDA 0.053331f
C797 two_stage_opamp_dummy_magic_21_0.VD1.n18 GNDA 0.116042f
C798 two_stage_opamp_dummy_magic_21_0.VD1.n19 GNDA 0.447102f
C799 two_stage_opamp_dummy_magic_21_0.VD1.n20 GNDA 0.099935f
C800 two_stage_opamp_dummy_magic_21_0.VD1.n21 GNDA 0.08441f
C801 two_stage_opamp_dummy_magic_21_0.VD1.t14 GNDA 0.053331f
C802 two_stage_opamp_dummy_magic_21_0.VD1.t19 GNDA 0.053331f
C803 two_stage_opamp_dummy_magic_21_0.VD1.n22 GNDA 0.116042f
C804 two_stage_opamp_dummy_magic_21_0.VD1.n23 GNDA 0.461069f
C805 two_stage_opamp_dummy_magic_21_0.VD1.n24 GNDA 0.203944f
C806 two_stage_opamp_dummy_magic_21_0.VD1.t21 GNDA 0.053331f
C807 two_stage_opamp_dummy_magic_21_0.VD1.t16 GNDA 0.053331f
C808 two_stage_opamp_dummy_magic_21_0.VD1.n25 GNDA 0.116042f
C809 two_stage_opamp_dummy_magic_21_0.VD1.n26 GNDA 0.442486f
C810 two_stage_opamp_dummy_magic_21_0.VD1.n27 GNDA 0.192793f
C811 two_stage_opamp_dummy_magic_21_0.VD1.t12 GNDA 0.053331f
C812 two_stage_opamp_dummy_magic_21_0.VD1.t17 GNDA 0.053331f
C813 two_stage_opamp_dummy_magic_21_0.VD1.n28 GNDA 0.116042f
C814 two_stage_opamp_dummy_magic_21_0.VD1.n29 GNDA 0.461069f
C815 two_stage_opamp_dummy_magic_21_0.VD1.n30 GNDA 0.203944f
C816 two_stage_opamp_dummy_magic_21_0.VD1.t13 GNDA 0.053331f
C817 two_stage_opamp_dummy_magic_21_0.VD1.t18 GNDA 0.053331f
C818 two_stage_opamp_dummy_magic_21_0.VD1.n31 GNDA 0.116042f
C819 two_stage_opamp_dummy_magic_21_0.VD1.n32 GNDA 0.442486f
C820 two_stage_opamp_dummy_magic_21_0.VD1.n33 GNDA 0.192793f
C821 two_stage_opamp_dummy_magic_21_0.VD1.n34 GNDA 0.106662f
C822 two_stage_opamp_dummy_magic_21_0.VD1.n35 GNDA 0.235249f
C823 two_stage_opamp_dummy_magic_21_0.VD1.n36 GNDA 0.361396f
C824 two_stage_opamp_dummy_magic_21_0.VD1.n37 GNDA 0.116042f
C825 two_stage_opamp_dummy_magic_21_0.VD1.t20 GNDA 0.053331f
C826 two_stage_opamp_dummy_magic_21_0.Vb1.n0 GNDA 0.037919f
C827 two_stage_opamp_dummy_magic_21_0.Vb1.n1 GNDA 0.184455f
C828 two_stage_opamp_dummy_magic_21_0.Vb1.t5 GNDA 0.01264f
C829 two_stage_opamp_dummy_magic_21_0.Vb1.t0 GNDA 0.01264f
C830 two_stage_opamp_dummy_magic_21_0.Vb1.n2 GNDA 0.031684f
C831 two_stage_opamp_dummy_magic_21_0.Vb1.t1 GNDA 0.01264f
C832 two_stage_opamp_dummy_magic_21_0.Vb1.t4 GNDA 0.01264f
C833 two_stage_opamp_dummy_magic_21_0.Vb1.n3 GNDA 0.031471f
C834 two_stage_opamp_dummy_magic_21_0.Vb1.n4 GNDA 0.345583f
C835 two_stage_opamp_dummy_magic_21_0.Vb1.t33 GNDA 0.592366f
C836 two_stage_opamp_dummy_magic_21_0.Vb1.n5 GNDA 0.163985f
C837 two_stage_opamp_dummy_magic_21_0.Vb1.t2 GNDA 0.01896f
C838 two_stage_opamp_dummy_magic_21_0.Vb1.t11 GNDA 0.01896f
C839 two_stage_opamp_dummy_magic_21_0.Vb1.n6 GNDA 0.041254f
C840 two_stage_opamp_dummy_magic_21_0.Vb1.n7 GNDA 0.165724f
C841 two_stage_opamp_dummy_magic_21_0.Vb1.t12 GNDA 0.019434f
C842 two_stage_opamp_dummy_magic_21_0.Vb1.t10 GNDA 0.025206f
C843 two_stage_opamp_dummy_magic_21_0.Vb1.n8 GNDA 0.025915f
C844 two_stage_opamp_dummy_magic_21_0.Vb1.t6 GNDA 0.019434f
C845 two_stage_opamp_dummy_magic_21_0.Vb1.t8 GNDA 0.025206f
C846 two_stage_opamp_dummy_magic_21_0.Vb1.n9 GNDA 0.025915f
C847 two_stage_opamp_dummy_magic_21_0.Vb1.n10 GNDA 0.019317f
C848 two_stage_opamp_dummy_magic_21_0.Vb1.t13 GNDA 0.01896f
C849 two_stage_opamp_dummy_magic_21_0.Vb1.t7 GNDA 0.01896f
C850 two_stage_opamp_dummy_magic_21_0.Vb1.n11 GNDA 0.041254f
C851 two_stage_opamp_dummy_magic_21_0.Vb1.n12 GNDA 0.102656f
C852 two_stage_opamp_dummy_magic_21_0.Vb1.t9 GNDA 0.01896f
C853 two_stage_opamp_dummy_magic_21_0.Vb1.t3 GNDA 0.01896f
C854 two_stage_opamp_dummy_magic_21_0.Vb1.n13 GNDA 0.041254f
C855 two_stage_opamp_dummy_magic_21_0.Vb1.n14 GNDA 0.165724f
C856 two_stage_opamp_dummy_magic_21_0.Vb1.n15 GNDA 0.295093f
C857 two_stage_opamp_dummy_magic_21_0.Vb1.t24 GNDA 0.019434f
C858 two_stage_opamp_dummy_magic_21_0.Vb1.t34 GNDA 0.019434f
C859 two_stage_opamp_dummy_magic_21_0.Vb1.t22 GNDA 0.019434f
C860 two_stage_opamp_dummy_magic_21_0.Vb1.t31 GNDA 0.019434f
C861 two_stage_opamp_dummy_magic_21_0.Vb1.t19 GNDA 0.019434f
C862 two_stage_opamp_dummy_magic_21_0.Vb1.t16 GNDA 0.019434f
C863 two_stage_opamp_dummy_magic_21_0.Vb1.t20 GNDA 0.019434f
C864 two_stage_opamp_dummy_magic_21_0.Vb1.t29 GNDA 0.019434f
C865 two_stage_opamp_dummy_magic_21_0.Vb1.t18 GNDA 0.019434f
C866 two_stage_opamp_dummy_magic_21_0.Vb1.t23 GNDA 0.019434f
C867 two_stage_opamp_dummy_magic_21_0.Vb1.t32 GNDA 0.019434f
C868 two_stage_opamp_dummy_magic_21_0.Vb1.t21 GNDA 0.019434f
C869 two_stage_opamp_dummy_magic_21_0.Vb1.t30 GNDA 0.019434f
C870 two_stage_opamp_dummy_magic_21_0.Vb1.t26 GNDA 0.019434f
C871 two_stage_opamp_dummy_magic_21_0.Vb1.t15 GNDA 0.019434f
C872 two_stage_opamp_dummy_magic_21_0.Vb1.t25 GNDA 0.019434f
C873 two_stage_opamp_dummy_magic_21_0.Vb1.t14 GNDA 0.019434f
C874 two_stage_opamp_dummy_magic_21_0.Vb1.t17 GNDA 0.019434f
C875 two_stage_opamp_dummy_magic_21_0.Vb1.t27 GNDA 0.025206f
C876 two_stage_opamp_dummy_magic_21_0.Vb1.n16 GNDA 0.027407f
C877 two_stage_opamp_dummy_magic_21_0.Vb1.n17 GNDA 0.018486f
C878 two_stage_opamp_dummy_magic_21_0.Vb1.n18 GNDA 0.018486f
C879 two_stage_opamp_dummy_magic_21_0.Vb1.n19 GNDA 0.018486f
C880 two_stage_opamp_dummy_magic_21_0.Vb1.n20 GNDA 0.018486f
C881 two_stage_opamp_dummy_magic_21_0.Vb1.n21 GNDA 0.018486f
C882 two_stage_opamp_dummy_magic_21_0.Vb1.n22 GNDA 0.018486f
C883 two_stage_opamp_dummy_magic_21_0.Vb1.n23 GNDA 0.018486f
C884 two_stage_opamp_dummy_magic_21_0.Vb1.n24 GNDA 0.143303f
C885 two_stage_opamp_dummy_magic_21_0.Vb1.t28 GNDA 0.019434f
C886 two_stage_opamp_dummy_magic_21_0.Vb1.n25 GNDA 0.143303f
C887 two_stage_opamp_dummy_magic_21_0.Vb1.n26 GNDA 0.018486f
C888 two_stage_opamp_dummy_magic_21_0.Vb1.n27 GNDA 0.018486f
C889 two_stage_opamp_dummy_magic_21_0.Vb1.n28 GNDA 0.018486f
C890 two_stage_opamp_dummy_magic_21_0.Vb1.n29 GNDA 0.018486f
C891 two_stage_opamp_dummy_magic_21_0.Vb1.n30 GNDA 0.018486f
C892 two_stage_opamp_dummy_magic_21_0.Vb1.n31 GNDA 0.018486f
C893 two_stage_opamp_dummy_magic_21_0.Vb1.n32 GNDA 0.018486f
C894 two_stage_opamp_dummy_magic_21_0.Vb1.n33 GNDA 0.018486f
C895 two_stage_opamp_dummy_magic_21_0.Vb1.n34 GNDA 0.032945f
C896 two_stage_opamp_dummy_magic_21_0.Vb1.n35 GNDA 1.12646f
C897 bgr_0.VB1_CUR_BIAS GNDA 0.68969f
C898 two_stage_opamp_dummy_magic_21_0.X.t22 GNDA 0.038289f
C899 two_stage_opamp_dummy_magic_21_0.X.t1 GNDA 0.038289f
C900 two_stage_opamp_dummy_magic_21_0.X.n0 GNDA 0.083312f
C901 two_stage_opamp_dummy_magic_21_0.X.n1 GNDA 0.259463f
C902 two_stage_opamp_dummy_magic_21_0.X.n2 GNDA 0.138415f
C903 two_stage_opamp_dummy_magic_21_0.X.n3 GNDA 0.138415f
C904 two_stage_opamp_dummy_magic_21_0.X.t19 GNDA 0.038289f
C905 two_stage_opamp_dummy_magic_21_0.X.t16 GNDA 0.038289f
C906 two_stage_opamp_dummy_magic_21_0.X.n4 GNDA 0.083312f
C907 two_stage_opamp_dummy_magic_21_0.X.n5 GNDA 0.331023f
C908 two_stage_opamp_dummy_magic_21_0.X.t2 GNDA 0.038289f
C909 two_stage_opamp_dummy_magic_21_0.X.t4 GNDA 0.038289f
C910 two_stage_opamp_dummy_magic_21_0.X.n6 GNDA 0.083312f
C911 two_stage_opamp_dummy_magic_21_0.X.n7 GNDA 0.317681f
C912 two_stage_opamp_dummy_magic_21_0.X.n8 GNDA 0.146421f
C913 two_stage_opamp_dummy_magic_21_0.X.n9 GNDA 0.085527f
C914 two_stage_opamp_dummy_magic_21_0.X.t24 GNDA 0.038289f
C915 two_stage_opamp_dummy_magic_21_0.X.t20 GNDA 0.038289f
C916 two_stage_opamp_dummy_magic_21_0.X.n10 GNDA 0.083312f
C917 two_stage_opamp_dummy_magic_21_0.X.n11 GNDA 0.331023f
C918 two_stage_opamp_dummy_magic_21_0.X.t0 GNDA 0.038289f
C919 two_stage_opamp_dummy_magic_21_0.X.t21 GNDA 0.038289f
C920 two_stage_opamp_dummy_magic_21_0.X.n12 GNDA 0.083312f
C921 two_stage_opamp_dummy_magic_21_0.X.n13 GNDA 0.317681f
C922 two_stage_opamp_dummy_magic_21_0.X.n14 GNDA 0.146421f
C923 two_stage_opamp_dummy_magic_21_0.X.n15 GNDA 0.085527f
C924 two_stage_opamp_dummy_magic_21_0.X.t23 GNDA 0.038289f
C925 two_stage_opamp_dummy_magic_21_0.X.t15 GNDA 0.038289f
C926 two_stage_opamp_dummy_magic_21_0.X.n16 GNDA 0.083312f
C927 two_stage_opamp_dummy_magic_21_0.X.n17 GNDA 0.317681f
C928 two_stage_opamp_dummy_magic_21_0.X.n18 GNDA 0.081429f
C929 two_stage_opamp_dummy_magic_21_0.X.n19 GNDA 0.076577f
C930 two_stage_opamp_dummy_magic_21_0.X.n20 GNDA 0.145807f
C931 two_stage_opamp_dummy_magic_21_0.X.t18 GNDA 1.22341f
C932 two_stage_opamp_dummy_magic_21_0.X.t50 GNDA 0.16847f
C933 two_stage_opamp_dummy_magic_21_0.X.t38 GNDA 0.16847f
C934 two_stage_opamp_dummy_magic_21_0.X.t53 GNDA 0.16847f
C935 two_stage_opamp_dummy_magic_21_0.X.t40 GNDA 0.16847f
C936 two_stage_opamp_dummy_magic_21_0.X.t26 GNDA 0.16847f
C937 two_stage_opamp_dummy_magic_21_0.X.t39 GNDA 0.16847f
C938 two_stage_opamp_dummy_magic_21_0.X.t25 GNDA 0.179433f
C939 two_stage_opamp_dummy_magic_21_0.X.n21 GNDA 0.142193f
C940 two_stage_opamp_dummy_magic_21_0.X.n22 GNDA 0.080406f
C941 two_stage_opamp_dummy_magic_21_0.X.n23 GNDA 0.080406f
C942 two_stage_opamp_dummy_magic_21_0.X.n24 GNDA 0.080406f
C943 two_stage_opamp_dummy_magic_21_0.X.n25 GNDA 0.080406f
C944 two_stage_opamp_dummy_magic_21_0.X.n26 GNDA 0.07227f
C945 two_stage_opamp_dummy_magic_21_0.X.t35 GNDA 0.16847f
C946 two_stage_opamp_dummy_magic_21_0.X.t48 GNDA 0.16847f
C947 two_stage_opamp_dummy_magic_21_0.X.t33 GNDA 0.179433f
C948 two_stage_opamp_dummy_magic_21_0.X.n27 GNDA 0.142193f
C949 two_stage_opamp_dummy_magic_21_0.X.n28 GNDA 0.07227f
C950 two_stage_opamp_dummy_magic_21_0.X.n29 GNDA 0.036557f
C951 two_stage_opamp_dummy_magic_21_0.X.n30 GNDA 1.2754f
C952 two_stage_opamp_dummy_magic_21_0.X.t17 GNDA 0.08934f
C953 two_stage_opamp_dummy_magic_21_0.X.t7 GNDA 0.08934f
C954 two_stage_opamp_dummy_magic_21_0.X.n31 GNDA 0.182755f
C955 two_stage_opamp_dummy_magic_21_0.X.n32 GNDA 0.497099f
C956 two_stage_opamp_dummy_magic_21_0.X.n33 GNDA 0.096905f
C957 two_stage_opamp_dummy_magic_21_0.X.n34 GNDA 0.16531f
C958 two_stage_opamp_dummy_magic_21_0.X.t12 GNDA 0.08934f
C959 two_stage_opamp_dummy_magic_21_0.X.t3 GNDA 0.08934f
C960 two_stage_opamp_dummy_magic_21_0.X.n35 GNDA 0.182755f
C961 two_stage_opamp_dummy_magic_21_0.X.n36 GNDA 0.591707f
C962 two_stage_opamp_dummy_magic_21_0.X.t10 GNDA 0.08934f
C963 two_stage_opamp_dummy_magic_21_0.X.t9 GNDA 0.08934f
C964 two_stage_opamp_dummy_magic_21_0.X.n37 GNDA 0.182755f
C965 two_stage_opamp_dummy_magic_21_0.X.n38 GNDA 0.575548f
C966 two_stage_opamp_dummy_magic_21_0.X.n39 GNDA 0.16531f
C967 two_stage_opamp_dummy_magic_21_0.X.n40 GNDA 0.096905f
C968 two_stage_opamp_dummy_magic_21_0.X.t14 GNDA 0.08934f
C969 two_stage_opamp_dummy_magic_21_0.X.t6 GNDA 0.08934f
C970 two_stage_opamp_dummy_magic_21_0.X.n41 GNDA 0.182755f
C971 two_stage_opamp_dummy_magic_21_0.X.n42 GNDA 0.575548f
C972 two_stage_opamp_dummy_magic_21_0.X.n43 GNDA 0.096905f
C973 two_stage_opamp_dummy_magic_21_0.X.t8 GNDA 0.08934f
C974 two_stage_opamp_dummy_magic_21_0.X.t11 GNDA 0.08934f
C975 two_stage_opamp_dummy_magic_21_0.X.n44 GNDA 0.182755f
C976 two_stage_opamp_dummy_magic_21_0.X.n45 GNDA 0.575548f
C977 two_stage_opamp_dummy_magic_21_0.X.n46 GNDA 0.096905f
C978 two_stage_opamp_dummy_magic_21_0.X.n47 GNDA 0.16531f
C979 two_stage_opamp_dummy_magic_21_0.X.t5 GNDA 0.08934f
C980 two_stage_opamp_dummy_magic_21_0.X.t13 GNDA 0.08934f
C981 two_stage_opamp_dummy_magic_21_0.X.n48 GNDA 0.182755f
C982 two_stage_opamp_dummy_magic_21_0.X.n49 GNDA 0.575548f
C983 two_stage_opamp_dummy_magic_21_0.X.n50 GNDA 0.150696f
C984 two_stage_opamp_dummy_magic_21_0.X.n51 GNDA 0.491162f
C985 two_stage_opamp_dummy_magic_21_0.X.t31 GNDA 0.053604f
C986 two_stage_opamp_dummy_magic_21_0.X.t46 GNDA 0.065091f
C987 two_stage_opamp_dummy_magic_21_0.X.n52 GNDA 0.056954f
C988 two_stage_opamp_dummy_magic_21_0.X.t47 GNDA 0.053604f
C989 two_stage_opamp_dummy_magic_21_0.X.t32 GNDA 0.053604f
C990 two_stage_opamp_dummy_magic_21_0.X.t44 GNDA 0.053604f
C991 two_stage_opamp_dummy_magic_21_0.X.t29 GNDA 0.053604f
C992 two_stage_opamp_dummy_magic_21_0.X.t42 GNDA 0.053604f
C993 two_stage_opamp_dummy_magic_21_0.X.t27 GNDA 0.053604f
C994 two_stage_opamp_dummy_magic_21_0.X.t41 GNDA 0.053604f
C995 two_stage_opamp_dummy_magic_21_0.X.t54 GNDA 0.065091f
C996 two_stage_opamp_dummy_magic_21_0.X.n53 GNDA 0.065091f
C997 two_stage_opamp_dummy_magic_21_0.X.n54 GNDA 0.042118f
C998 two_stage_opamp_dummy_magic_21_0.X.n55 GNDA 0.042118f
C999 two_stage_opamp_dummy_magic_21_0.X.n56 GNDA 0.042118f
C1000 two_stage_opamp_dummy_magic_21_0.X.n57 GNDA 0.042118f
C1001 two_stage_opamp_dummy_magic_21_0.X.n58 GNDA 0.042118f
C1002 two_stage_opamp_dummy_magic_21_0.X.n59 GNDA 0.033981f
C1003 two_stage_opamp_dummy_magic_21_0.X.n60 GNDA 0.021431f
C1004 two_stage_opamp_dummy_magic_21_0.X.t36 GNDA 0.082321f
C1005 two_stage_opamp_dummy_magic_21_0.X.t51 GNDA 0.093585f
C1006 two_stage_opamp_dummy_magic_21_0.X.n61 GNDA 0.076321f
C1007 two_stage_opamp_dummy_magic_21_0.X.t52 GNDA 0.082321f
C1008 two_stage_opamp_dummy_magic_21_0.X.t37 GNDA 0.082321f
C1009 two_stage_opamp_dummy_magic_21_0.X.t49 GNDA 0.082321f
C1010 two_stage_opamp_dummy_magic_21_0.X.t34 GNDA 0.082321f
C1011 two_stage_opamp_dummy_magic_21_0.X.t45 GNDA 0.082321f
C1012 two_stage_opamp_dummy_magic_21_0.X.t30 GNDA 0.082321f
C1013 two_stage_opamp_dummy_magic_21_0.X.t43 GNDA 0.082321f
C1014 two_stage_opamp_dummy_magic_21_0.X.t28 GNDA 0.093585f
C1015 two_stage_opamp_dummy_magic_21_0.X.n62 GNDA 0.084458f
C1016 two_stage_opamp_dummy_magic_21_0.X.n63 GNDA 0.05169f
C1017 two_stage_opamp_dummy_magic_21_0.X.n64 GNDA 0.05169f
C1018 two_stage_opamp_dummy_magic_21_0.X.n65 GNDA 0.05169f
C1019 two_stage_opamp_dummy_magic_21_0.X.n66 GNDA 0.05169f
C1020 two_stage_opamp_dummy_magic_21_0.X.n67 GNDA 0.05169f
C1021 two_stage_opamp_dummy_magic_21_0.X.n68 GNDA 0.043554f
C1022 two_stage_opamp_dummy_magic_21_0.X.n69 GNDA 0.021431f
C1023 two_stage_opamp_dummy_magic_21_0.X.n70 GNDA 0.092553f
C1024 two_stage_opamp_dummy_magic_21_0.X.n71 GNDA 1.05185f
C1025 two_stage_opamp_dummy_magic_21_0.X.n72 GNDA 0.412424f
C1026 two_stage_opamp_dummy_magic_21_0.X.n73 GNDA 0.199954f
C1027 two_stage_opamp_dummy_magic_21_0.V_err_p.n0 GNDA 0.381408f
C1028 two_stage_opamp_dummy_magic_21_0.V_err_p.n1 GNDA 0.241974f
C1029 two_stage_opamp_dummy_magic_21_0.V_err_p.n2 GNDA 0.397193f
C1030 two_stage_opamp_dummy_magic_21_0.V_err_p.n3 GNDA 0.457146f
C1031 two_stage_opamp_dummy_magic_21_0.V_err_p.n4 GNDA 0.388376f
C1032 two_stage_opamp_dummy_magic_21_0.V_err_p.t21 GNDA 0.023181f
C1033 two_stage_opamp_dummy_magic_21_0.V_err_p.t10 GNDA 0.023181f
C1034 two_stage_opamp_dummy_magic_21_0.V_err_p.t13 GNDA 0.023181f
C1035 two_stage_opamp_dummy_magic_21_0.V_err_p.n5 GNDA 0.047234f
C1036 two_stage_opamp_dummy_magic_21_0.V_err_p.n6 GNDA 0.348058f
C1037 two_stage_opamp_dummy_magic_21_0.V_err_p.t3 GNDA 0.023181f
C1038 two_stage_opamp_dummy_magic_21_0.V_err_p.t2 GNDA 0.023181f
C1039 two_stage_opamp_dummy_magic_21_0.V_err_p.n7 GNDA 0.047234f
C1040 two_stage_opamp_dummy_magic_21_0.V_err_p.t20 GNDA 0.023181f
C1041 two_stage_opamp_dummy_magic_21_0.V_err_p.t1 GNDA 0.023181f
C1042 two_stage_opamp_dummy_magic_21_0.V_err_p.n8 GNDA 0.047234f
C1043 two_stage_opamp_dummy_magic_21_0.V_err_p.n9 GNDA 0.392203f
C1044 two_stage_opamp_dummy_magic_21_0.V_err_p.n10 GNDA 0.243876f
C1045 two_stage_opamp_dummy_magic_21_0.V_err_p.n11 GNDA 0.38098f
C1046 two_stage_opamp_dummy_magic_21_0.V_err_p.t17 GNDA 0.023181f
C1047 two_stage_opamp_dummy_magic_21_0.V_err_p.t19 GNDA 0.023181f
C1048 two_stage_opamp_dummy_magic_21_0.V_err_p.n12 GNDA 0.047234f
C1049 two_stage_opamp_dummy_magic_21_0.V_err_p.n13 GNDA 0.392203f
C1050 two_stage_opamp_dummy_magic_21_0.V_err_p.n14 GNDA 0.370407f
C1051 two_stage_opamp_dummy_magic_21_0.V_err_p.t14 GNDA 0.023181f
C1052 two_stage_opamp_dummy_magic_21_0.V_err_p.t5 GNDA 0.023181f
C1053 two_stage_opamp_dummy_magic_21_0.V_err_p.n15 GNDA 0.047234f
C1054 two_stage_opamp_dummy_magic_21_0.V_err_p.n16 GNDA 0.324373f
C1055 two_stage_opamp_dummy_magic_21_0.V_err_p.n17 GNDA 0.38098f
C1056 two_stage_opamp_dummy_magic_21_0.V_err_p.t16 GNDA 0.023181f
C1057 two_stage_opamp_dummy_magic_21_0.V_err_p.t4 GNDA 0.023181f
C1058 two_stage_opamp_dummy_magic_21_0.V_err_p.n18 GNDA 0.047234f
C1059 two_stage_opamp_dummy_magic_21_0.V_err_p.n19 GNDA 0.324373f
C1060 two_stage_opamp_dummy_magic_21_0.V_err_p.n20 GNDA 0.249186f
C1061 two_stage_opamp_dummy_magic_21_0.V_err_p.n21 GNDA 0.249186f
C1062 two_stage_opamp_dummy_magic_21_0.V_err_p.t18 GNDA 0.023181f
C1063 two_stage_opamp_dummy_magic_21_0.V_err_p.t12 GNDA 0.023181f
C1064 two_stage_opamp_dummy_magic_21_0.V_err_p.n22 GNDA 0.047234f
C1065 two_stage_opamp_dummy_magic_21_0.V_err_p.n23 GNDA 0.324373f
C1066 two_stage_opamp_dummy_magic_21_0.V_err_p.n24 GNDA 0.243876f
C1067 two_stage_opamp_dummy_magic_21_0.V_err_p.n25 GNDA 0.367618f
C1068 two_stage_opamp_dummy_magic_21_0.V_err_p.t9 GNDA 0.023181f
C1069 two_stage_opamp_dummy_magic_21_0.V_err_p.t6 GNDA 0.023181f
C1070 two_stage_opamp_dummy_magic_21_0.V_err_p.n26 GNDA 0.047234f
C1071 two_stage_opamp_dummy_magic_21_0.V_err_p.t15 GNDA 0.023181f
C1072 two_stage_opamp_dummy_magic_21_0.V_err_p.t7 GNDA 0.023181f
C1073 two_stage_opamp_dummy_magic_21_0.V_err_p.n27 GNDA 0.047234f
C1074 two_stage_opamp_dummy_magic_21_0.V_err_p.n28 GNDA 0.324373f
C1075 two_stage_opamp_dummy_magic_21_0.V_err_p.t8 GNDA 0.023181f
C1076 two_stage_opamp_dummy_magic_21_0.V_err_p.t0 GNDA 0.023181f
C1077 two_stage_opamp_dummy_magic_21_0.V_err_p.n29 GNDA 0.047234f
C1078 two_stage_opamp_dummy_magic_21_0.V_err_p.n30 GNDA 0.324373f
C1079 two_stage_opamp_dummy_magic_21_0.V_err_p.n31 GNDA 0.239531f
C1080 two_stage_opamp_dummy_magic_21_0.V_err_p.n32 GNDA 0.324373f
C1081 two_stage_opamp_dummy_magic_21_0.V_err_p.n33 GNDA 0.047234f
C1082 two_stage_opamp_dummy_magic_21_0.V_err_p.t11 GNDA 0.023181f
C1083 two_stage_opamp_dummy_magic_21_0.VD4.t25 GNDA 0.060801f
C1084 two_stage_opamp_dummy_magic_21_0.VD4.t9 GNDA 0.060801f
C1085 two_stage_opamp_dummy_magic_21_0.VD4.n0 GNDA 0.154331f
C1086 two_stage_opamp_dummy_magic_21_0.VD4.n1 GNDA 0.431096f
C1087 two_stage_opamp_dummy_magic_21_0.VD4.t0 GNDA 0.106612f
C1088 two_stage_opamp_dummy_magic_21_0.VD4.t5 GNDA 0.216278f
C1089 two_stage_opamp_dummy_magic_21_0.VD4.t17 GNDA 0.060801f
C1090 two_stage_opamp_dummy_magic_21_0.VD4.t21 GNDA 0.060801f
C1091 two_stage_opamp_dummy_magic_21_0.VD4.n2 GNDA 0.154331f
C1092 two_stage_opamp_dummy_magic_21_0.VD4.n3 GNDA 0.431096f
C1093 two_stage_opamp_dummy_magic_21_0.VD4.t11 GNDA 0.060801f
C1094 two_stage_opamp_dummy_magic_21_0.VD4.t13 GNDA 0.060801f
C1095 two_stage_opamp_dummy_magic_21_0.VD4.n4 GNDA 0.154331f
C1096 two_stage_opamp_dummy_magic_21_0.VD4.n5 GNDA 0.431096f
C1097 two_stage_opamp_dummy_magic_21_0.VD4.t23 GNDA 0.060801f
C1098 two_stage_opamp_dummy_magic_21_0.VD4.t7 GNDA 0.060801f
C1099 two_stage_opamp_dummy_magic_21_0.VD4.n6 GNDA 0.154331f
C1100 two_stage_opamp_dummy_magic_21_0.VD4.n7 GNDA 0.431096f
C1101 two_stage_opamp_dummy_magic_21_0.VD4.t15 GNDA 0.060801f
C1102 two_stage_opamp_dummy_magic_21_0.VD4.t19 GNDA 0.060801f
C1103 two_stage_opamp_dummy_magic_21_0.VD4.n8 GNDA 0.154331f
C1104 two_stage_opamp_dummy_magic_21_0.VD4.n9 GNDA 0.481515f
C1105 two_stage_opamp_dummy_magic_21_0.VD4.t3 GNDA 0.106612f
C1106 two_stage_opamp_dummy_magic_21_0.VD4.n10 GNDA 0.316782f
C1107 two_stage_opamp_dummy_magic_21_0.VD4.n11 GNDA 0.627403f
C1108 two_stage_opamp_dummy_magic_21_0.VD4.t4 GNDA 0.518263f
C1109 two_stage_opamp_dummy_magic_21_0.VD4.t14 GNDA 0.406498f
C1110 two_stage_opamp_dummy_magic_21_0.VD4.t18 GNDA 0.406498f
C1111 two_stage_opamp_dummy_magic_21_0.VD4.t22 GNDA 0.406498f
C1112 two_stage_opamp_dummy_magic_21_0.VD4.t6 GNDA 0.406498f
C1113 two_stage_opamp_dummy_magic_21_0.VD4.t10 GNDA 0.406498f
C1114 two_stage_opamp_dummy_magic_21_0.VD4.t12 GNDA 0.406498f
C1115 two_stage_opamp_dummy_magic_21_0.VD4.t16 GNDA 0.406498f
C1116 two_stage_opamp_dummy_magic_21_0.VD4.t20 GNDA 0.406498f
C1117 two_stage_opamp_dummy_magic_21_0.VD4.t24 GNDA 0.406498f
C1118 two_stage_opamp_dummy_magic_21_0.VD4.t8 GNDA 0.406498f
C1119 two_stage_opamp_dummy_magic_21_0.VD4.t1 GNDA 0.518263f
C1120 two_stage_opamp_dummy_magic_21_0.VD4.t2 GNDA 0.216278f
C1121 two_stage_opamp_dummy_magic_21_0.VD4.n12 GNDA 0.627403f
C1122 two_stage_opamp_dummy_magic_21_0.VD4.n13 GNDA 0.311031f
C1123 two_stage_opamp_dummy_magic_21_0.VD4.n14 GNDA 0.102448f
C1124 two_stage_opamp_dummy_magic_21_0.VD4.n15 GNDA 0.065949f
C1125 two_stage_opamp_dummy_magic_21_0.VD4.n16 GNDA 0.065949f
C1126 two_stage_opamp_dummy_magic_21_0.VD4.t35 GNDA 0.060801f
C1127 two_stage_opamp_dummy_magic_21_0.VD4.t37 GNDA 0.060801f
C1128 two_stage_opamp_dummy_magic_21_0.VD4.n17 GNDA 0.124375f
C1129 two_stage_opamp_dummy_magic_21_0.VD4.n18 GNDA 0.402689f
C1130 two_stage_opamp_dummy_magic_21_0.VD4.n19 GNDA 0.112503f
C1131 two_stage_opamp_dummy_magic_21_0.VD4.t28 GNDA 0.060801f
C1132 two_stage_opamp_dummy_magic_21_0.VD4.t32 GNDA 0.060801f
C1133 two_stage_opamp_dummy_magic_21_0.VD4.n20 GNDA 0.124375f
C1134 two_stage_opamp_dummy_magic_21_0.VD4.n21 GNDA 0.391692f
C1135 two_stage_opamp_dummy_magic_21_0.VD4.n22 GNDA 0.112503f
C1136 two_stage_opamp_dummy_magic_21_0.VD4.t27 GNDA 0.060801f
C1137 two_stage_opamp_dummy_magic_21_0.VD4.t30 GNDA 0.060801f
C1138 two_stage_opamp_dummy_magic_21_0.VD4.n23 GNDA 0.124375f
C1139 two_stage_opamp_dummy_magic_21_0.VD4.n24 GNDA 0.391692f
C1140 two_stage_opamp_dummy_magic_21_0.VD4.n25 GNDA 0.065949f
C1141 two_stage_opamp_dummy_magic_21_0.VD4.n26 GNDA 0.065949f
C1142 two_stage_opamp_dummy_magic_21_0.VD4.t34 GNDA 0.060801f
C1143 two_stage_opamp_dummy_magic_21_0.VD4.t26 GNDA 0.060801f
C1144 two_stage_opamp_dummy_magic_21_0.VD4.n27 GNDA 0.124375f
C1145 two_stage_opamp_dummy_magic_21_0.VD4.n28 GNDA 0.391692f
C1146 two_stage_opamp_dummy_magic_21_0.VD4.n29 GNDA 0.065949f
C1147 two_stage_opamp_dummy_magic_21_0.VD4.t33 GNDA 0.060801f
C1148 two_stage_opamp_dummy_magic_21_0.VD4.t31 GNDA 0.060801f
C1149 two_stage_opamp_dummy_magic_21_0.VD4.n30 GNDA 0.124375f
C1150 two_stage_opamp_dummy_magic_21_0.VD4.n31 GNDA 0.391692f
C1151 two_stage_opamp_dummy_magic_21_0.VD4.n32 GNDA 0.112503f
C1152 two_stage_opamp_dummy_magic_21_0.VD4.t36 GNDA 0.060801f
C1153 two_stage_opamp_dummy_magic_21_0.VD4.t29 GNDA 0.060801f
C1154 two_stage_opamp_dummy_magic_21_0.VD4.n33 GNDA 0.124375f
C1155 two_stage_opamp_dummy_magic_21_0.VD4.n34 GNDA 0.39719f
C1156 two_stage_opamp_dummy_magic_21_0.VD4.n35 GNDA 0.183347f
C1157 two_stage_opamp_dummy_magic_21_0.Vb2.t1 GNDA 0.028992f
C1158 two_stage_opamp_dummy_magic_21_0.Vb2.t10 GNDA 0.028992f
C1159 two_stage_opamp_dummy_magic_21_0.Vb2.n0 GNDA 0.061566f
C1160 two_stage_opamp_dummy_magic_21_0.Vb2.t0 GNDA 0.054119f
C1161 two_stage_opamp_dummy_magic_21_0.Vb2.n1 GNDA 0.250607f
C1162 two_stage_opamp_dummy_magic_21_0.Vb2.t13 GNDA 0.032501f
C1163 two_stage_opamp_dummy_magic_21_0.Vb2.n2 GNDA 0.124773f
C1164 two_stage_opamp_dummy_magic_21_0.Vb2.t18 GNDA 0.041003f
C1165 two_stage_opamp_dummy_magic_21_0.Vb2.t31 GNDA 0.041003f
C1166 two_stage_opamp_dummy_magic_21_0.Vb2.t25 GNDA 0.041003f
C1167 two_stage_opamp_dummy_magic_21_0.Vb2.t28 GNDA 0.041003f
C1168 two_stage_opamp_dummy_magic_21_0.Vb2.t22 GNDA 0.047317f
C1169 two_stage_opamp_dummy_magic_21_0.Vb2.n3 GNDA 0.038416f
C1170 two_stage_opamp_dummy_magic_21_0.Vb2.n4 GNDA 0.023607f
C1171 two_stage_opamp_dummy_magic_21_0.Vb2.n5 GNDA 0.023607f
C1172 two_stage_opamp_dummy_magic_21_0.Vb2.n6 GNDA 0.020699f
C1173 two_stage_opamp_dummy_magic_21_0.Vb2.t20 GNDA 0.041003f
C1174 two_stage_opamp_dummy_magic_21_0.Vb2.t23 GNDA 0.041003f
C1175 two_stage_opamp_dummy_magic_21_0.Vb2.t21 GNDA 0.041003f
C1176 two_stage_opamp_dummy_magic_21_0.Vb2.t26 GNDA 0.041003f
C1177 two_stage_opamp_dummy_magic_21_0.Vb2.t32 GNDA 0.047317f
C1178 two_stage_opamp_dummy_magic_21_0.Vb2.n7 GNDA 0.038416f
C1179 two_stage_opamp_dummy_magic_21_0.Vb2.n8 GNDA 0.023607f
C1180 two_stage_opamp_dummy_magic_21_0.Vb2.n9 GNDA 0.023607f
C1181 two_stage_opamp_dummy_magic_21_0.Vb2.n10 GNDA 0.020699f
C1182 two_stage_opamp_dummy_magic_21_0.Vb2.n11 GNDA 0.015341f
C1183 two_stage_opamp_dummy_magic_21_0.Vb2.t19 GNDA 0.041003f
C1184 two_stage_opamp_dummy_magic_21_0.Vb2.t16 GNDA 0.041003f
C1185 two_stage_opamp_dummy_magic_21_0.Vb2.t14 GNDA 0.041003f
C1186 two_stage_opamp_dummy_magic_21_0.Vb2.t11 GNDA 0.041003f
C1187 two_stage_opamp_dummy_magic_21_0.Vb2.t29 GNDA 0.047317f
C1188 two_stage_opamp_dummy_magic_21_0.Vb2.n12 GNDA 0.038416f
C1189 two_stage_opamp_dummy_magic_21_0.Vb2.n13 GNDA 0.023607f
C1190 two_stage_opamp_dummy_magic_21_0.Vb2.n14 GNDA 0.023607f
C1191 two_stage_opamp_dummy_magic_21_0.Vb2.n15 GNDA 0.020699f
C1192 two_stage_opamp_dummy_magic_21_0.Vb2.t24 GNDA 0.041003f
C1193 two_stage_opamp_dummy_magic_21_0.Vb2.t30 GNDA 0.041003f
C1194 two_stage_opamp_dummy_magic_21_0.Vb2.t12 GNDA 0.041003f
C1195 two_stage_opamp_dummy_magic_21_0.Vb2.t15 GNDA 0.041003f
C1196 two_stage_opamp_dummy_magic_21_0.Vb2.t17 GNDA 0.047317f
C1197 two_stage_opamp_dummy_magic_21_0.Vb2.n16 GNDA 0.038416f
C1198 two_stage_opamp_dummy_magic_21_0.Vb2.n17 GNDA 0.023607f
C1199 two_stage_opamp_dummy_magic_21_0.Vb2.n18 GNDA 0.023607f
C1200 two_stage_opamp_dummy_magic_21_0.Vb2.n19 GNDA 0.020699f
C1201 two_stage_opamp_dummy_magic_21_0.Vb2.n20 GNDA 0.015116f
C1202 two_stage_opamp_dummy_magic_21_0.Vb2.n21 GNDA 0.329492f
C1203 two_stage_opamp_dummy_magic_21_0.Vb2.n22 GNDA 0.153664f
C1204 two_stage_opamp_dummy_magic_21_0.Vb2.t27 GNDA 0.053285f
C1205 two_stage_opamp_dummy_magic_21_0.Vb2.n23 GNDA 0.680954f
C1206 two_stage_opamp_dummy_magic_21_0.Vb2.n24 GNDA 0.02739f
C1207 two_stage_opamp_dummy_magic_21_0.Vb2.n25 GNDA 0.746366f
C1208 two_stage_opamp_dummy_magic_21_0.Vb2.n26 GNDA 0.02739f
C1209 two_stage_opamp_dummy_magic_21_0.Vb2.n27 GNDA 0.192118f
C1210 two_stage_opamp_dummy_magic_21_0.Vb2.n28 GNDA 0.02822f
C1211 two_stage_opamp_dummy_magic_21_0.Vb2.n29 GNDA 0.284835f
C1212 two_stage_opamp_dummy_magic_21_0.Vb2.n30 GNDA 0.02739f
C1213 two_stage_opamp_dummy_magic_21_0.V_source.t15 GNDA 0.038168f
C1214 two_stage_opamp_dummy_magic_21_0.V_source.t33 GNDA 0.022901f
C1215 two_stage_opamp_dummy_magic_21_0.V_source.t39 GNDA 0.022901f
C1216 two_stage_opamp_dummy_magic_21_0.V_source.n0 GNDA 0.049829f
C1217 two_stage_opamp_dummy_magic_21_0.V_source.n1 GNDA 0.153174f
C1218 two_stage_opamp_dummy_magic_21_0.V_source.n2 GNDA 0.051155f
C1219 two_stage_opamp_dummy_magic_21_0.V_source.t34 GNDA 0.022901f
C1220 two_stage_opamp_dummy_magic_21_0.V_source.t40 GNDA 0.022901f
C1221 two_stage_opamp_dummy_magic_21_0.V_source.n3 GNDA 0.049829f
C1222 two_stage_opamp_dummy_magic_21_0.V_source.n4 GNDA 0.200044f
C1223 two_stage_opamp_dummy_magic_21_0.V_source.n5 GNDA 0.087575f
C1224 two_stage_opamp_dummy_magic_21_0.V_source.t32 GNDA 0.022901f
C1225 two_stage_opamp_dummy_magic_21_0.V_source.t1 GNDA 0.022901f
C1226 two_stage_opamp_dummy_magic_21_0.V_source.n6 GNDA 0.049829f
C1227 two_stage_opamp_dummy_magic_21_0.V_source.n7 GNDA 0.192055f
C1228 two_stage_opamp_dummy_magic_21_0.V_source.n8 GNDA 0.083262f
C1229 two_stage_opamp_dummy_magic_21_0.V_source.t6 GNDA 0.022901f
C1230 two_stage_opamp_dummy_magic_21_0.V_source.t27 GNDA 0.022901f
C1231 two_stage_opamp_dummy_magic_21_0.V_source.n9 GNDA 0.049829f
C1232 two_stage_opamp_dummy_magic_21_0.V_source.n10 GNDA 0.192055f
C1233 two_stage_opamp_dummy_magic_21_0.V_source.n11 GNDA 0.048946f
C1234 two_stage_opamp_dummy_magic_21_0.V_source.n12 GNDA 0.083262f
C1235 two_stage_opamp_dummy_magic_21_0.V_source.t7 GNDA 0.022901f
C1236 two_stage_opamp_dummy_magic_21_0.V_source.t5 GNDA 0.022901f
C1237 two_stage_opamp_dummy_magic_21_0.V_source.n13 GNDA 0.049829f
C1238 two_stage_opamp_dummy_magic_21_0.V_source.n14 GNDA 0.192055f
C1239 two_stage_opamp_dummy_magic_21_0.V_source.n15 GNDA 0.051155f
C1240 two_stage_opamp_dummy_magic_21_0.V_source.n16 GNDA 0.051155f
C1241 two_stage_opamp_dummy_magic_21_0.V_source.n17 GNDA 0.083262f
C1242 two_stage_opamp_dummy_magic_21_0.V_source.t30 GNDA 0.022901f
C1243 two_stage_opamp_dummy_magic_21_0.V_source.t36 GNDA 0.022901f
C1244 two_stage_opamp_dummy_magic_21_0.V_source.n18 GNDA 0.049829f
C1245 two_stage_opamp_dummy_magic_21_0.V_source.n19 GNDA 0.200044f
C1246 two_stage_opamp_dummy_magic_21_0.V_source.t3 GNDA 0.022901f
C1247 two_stage_opamp_dummy_magic_21_0.V_source.t38 GNDA 0.022901f
C1248 two_stage_opamp_dummy_magic_21_0.V_source.n20 GNDA 0.049829f
C1249 two_stage_opamp_dummy_magic_21_0.V_source.n21 GNDA 0.192055f
C1250 two_stage_opamp_dummy_magic_21_0.V_source.n22 GNDA 0.087575f
C1251 two_stage_opamp_dummy_magic_21_0.V_source.n23 GNDA 0.051155f
C1252 two_stage_opamp_dummy_magic_21_0.V_source.t0 GNDA 0.022901f
C1253 two_stage_opamp_dummy_magic_21_0.V_source.t28 GNDA 0.022901f
C1254 two_stage_opamp_dummy_magic_21_0.V_source.n24 GNDA 0.049829f
C1255 two_stage_opamp_dummy_magic_21_0.V_source.n25 GNDA 0.192055f
C1256 two_stage_opamp_dummy_magic_21_0.V_source.n26 GNDA 0.048946f
C1257 two_stage_opamp_dummy_magic_21_0.V_source.t2 GNDA 0.022901f
C1258 two_stage_opamp_dummy_magic_21_0.V_source.t29 GNDA 0.022901f
C1259 two_stage_opamp_dummy_magic_21_0.V_source.n27 GNDA 0.049829f
C1260 two_stage_opamp_dummy_magic_21_0.V_source.n28 GNDA 0.192055f
C1261 two_stage_opamp_dummy_magic_21_0.V_source.n29 GNDA 0.083262f
C1262 two_stage_opamp_dummy_magic_21_0.V_source.t31 GNDA 0.022901f
C1263 two_stage_opamp_dummy_magic_21_0.V_source.t37 GNDA 0.022901f
C1264 two_stage_opamp_dummy_magic_21_0.V_source.n30 GNDA 0.049829f
C1265 two_stage_opamp_dummy_magic_21_0.V_source.n31 GNDA 0.195998f
C1266 two_stage_opamp_dummy_magic_21_0.V_source.n32 GNDA 0.125964f
C1267 two_stage_opamp_dummy_magic_21_0.V_source.n33 GNDA 0.120611f
C1268 two_stage_opamp_dummy_magic_21_0.V_source.n34 GNDA 0.087586f
C1269 two_stage_opamp_dummy_magic_21_0.V_source.n35 GNDA 0.099442f
C1270 two_stage_opamp_dummy_magic_21_0.V_source.t4 GNDA 0.079851f
C1271 two_stage_opamp_dummy_magic_21_0.V_source.n36 GNDA 0.096361f
C1272 two_stage_opamp_dummy_magic_21_0.V_source.n37 GNDA 0.05567f
C1273 two_stage_opamp_dummy_magic_21_0.V_source.t35 GNDA 0.038168f
C1274 two_stage_opamp_dummy_magic_21_0.V_source.t8 GNDA 0.038168f
C1275 two_stage_opamp_dummy_magic_21_0.V_source.n38 GNDA 0.081597f
C1276 two_stage_opamp_dummy_magic_21_0.V_source.n39 GNDA 0.294282f
C1277 two_stage_opamp_dummy_magic_21_0.V_source.t25 GNDA 0.038168f
C1278 two_stage_opamp_dummy_magic_21_0.V_source.t19 GNDA 0.038168f
C1279 two_stage_opamp_dummy_magic_21_0.V_source.n40 GNDA 0.081597f
C1280 two_stage_opamp_dummy_magic_21_0.V_source.n41 GNDA 0.285878f
C1281 two_stage_opamp_dummy_magic_21_0.V_source.n42 GNDA 0.090055f
C1282 two_stage_opamp_dummy_magic_21_0.V_source.n43 GNDA 0.045802f
C1283 two_stage_opamp_dummy_magic_21_0.V_source.n44 GNDA 0.052428f
C1284 two_stage_opamp_dummy_magic_21_0.V_source.n45 GNDA 0.096361f
C1285 two_stage_opamp_dummy_magic_21_0.V_source.t12 GNDA 0.038168f
C1286 two_stage_opamp_dummy_magic_21_0.V_source.t18 GNDA 0.038168f
C1287 two_stage_opamp_dummy_magic_21_0.V_source.n46 GNDA 0.081597f
C1288 two_stage_opamp_dummy_magic_21_0.V_source.n47 GNDA 0.294282f
C1289 two_stage_opamp_dummy_magic_21_0.V_source.t14 GNDA 0.038168f
C1290 two_stage_opamp_dummy_magic_21_0.V_source.t22 GNDA 0.038168f
C1291 two_stage_opamp_dummy_magic_21_0.V_source.n48 GNDA 0.081597f
C1292 two_stage_opamp_dummy_magic_21_0.V_source.n49 GNDA 0.285878f
C1293 two_stage_opamp_dummy_magic_21_0.V_source.n50 GNDA 0.090055f
C1294 two_stage_opamp_dummy_magic_21_0.V_source.n51 GNDA 0.052428f
C1295 two_stage_opamp_dummy_magic_21_0.V_source.t16 GNDA 0.038168f
C1296 two_stage_opamp_dummy_magic_21_0.V_source.t24 GNDA 0.038168f
C1297 two_stage_opamp_dummy_magic_21_0.V_source.n52 GNDA 0.081597f
C1298 two_stage_opamp_dummy_magic_21_0.V_source.n53 GNDA 0.285878f
C1299 two_stage_opamp_dummy_magic_21_0.V_source.n54 GNDA 0.05567f
C1300 two_stage_opamp_dummy_magic_21_0.V_source.t20 GNDA 0.038168f
C1301 two_stage_opamp_dummy_magic_21_0.V_source.t10 GNDA 0.038168f
C1302 two_stage_opamp_dummy_magic_21_0.V_source.n55 GNDA 0.081597f
C1303 two_stage_opamp_dummy_magic_21_0.V_source.n56 GNDA 0.285878f
C1304 two_stage_opamp_dummy_magic_21_0.V_source.n57 GNDA 0.05567f
C1305 two_stage_opamp_dummy_magic_21_0.V_source.n58 GNDA 0.05567f
C1306 two_stage_opamp_dummy_magic_21_0.V_source.t17 GNDA 0.038168f
C1307 two_stage_opamp_dummy_magic_21_0.V_source.t9 GNDA 0.038168f
C1308 two_stage_opamp_dummy_magic_21_0.V_source.n59 GNDA 0.081597f
C1309 two_stage_opamp_dummy_magic_21_0.V_source.n60 GNDA 0.285878f
C1310 two_stage_opamp_dummy_magic_21_0.V_source.n61 GNDA 0.052428f
C1311 two_stage_opamp_dummy_magic_21_0.V_source.t21 GNDA 0.038168f
C1312 two_stage_opamp_dummy_magic_21_0.V_source.t11 GNDA 0.038168f
C1313 two_stage_opamp_dummy_magic_21_0.V_source.n62 GNDA 0.081597f
C1314 two_stage_opamp_dummy_magic_21_0.V_source.n63 GNDA 0.285878f
C1315 two_stage_opamp_dummy_magic_21_0.V_source.n64 GNDA 0.052428f
C1316 two_stage_opamp_dummy_magic_21_0.V_source.n65 GNDA 0.052428f
C1317 two_stage_opamp_dummy_magic_21_0.V_source.t23 GNDA 0.038168f
C1318 two_stage_opamp_dummy_magic_21_0.V_source.t13 GNDA 0.038168f
C1319 two_stage_opamp_dummy_magic_21_0.V_source.n66 GNDA 0.081597f
C1320 two_stage_opamp_dummy_magic_21_0.V_source.n67 GNDA 0.285878f
C1321 two_stage_opamp_dummy_magic_21_0.V_source.n68 GNDA 0.05567f
C1322 two_stage_opamp_dummy_magic_21_0.V_source.n69 GNDA 0.045802f
C1323 two_stage_opamp_dummy_magic_21_0.V_source.n70 GNDA 0.258117f
C1324 two_stage_opamp_dummy_magic_21_0.V_source.n71 GNDA 0.185859f
C1325 two_stage_opamp_dummy_magic_21_0.V_source.n72 GNDA 0.081597f
C1326 two_stage_opamp_dummy_magic_21_0.V_source.t26 GNDA 0.038168f
C1327 bgr_0.cap_res2.t7 GNDA 0.358376f
C1328 bgr_0.cap_res2.t13 GNDA 0.359675f
C1329 bgr_0.cap_res2.t15 GNDA 0.340442f
C1330 bgr_0.cap_res2.t1 GNDA 0.358376f
C1331 bgr_0.cap_res2.t6 GNDA 0.359675f
C1332 bgr_0.cap_res2.t9 GNDA 0.340442f
C1333 bgr_0.cap_res2.t5 GNDA 0.358376f
C1334 bgr_0.cap_res2.t11 GNDA 0.359675f
C1335 bgr_0.cap_res2.t14 GNDA 0.340442f
C1336 bgr_0.cap_res2.t20 GNDA 0.358376f
C1337 bgr_0.cap_res2.t4 GNDA 0.359675f
C1338 bgr_0.cap_res2.t8 GNDA 0.340442f
C1339 bgr_0.cap_res2.t16 GNDA 0.358376f
C1340 bgr_0.cap_res2.t19 GNDA 0.359675f
C1341 bgr_0.cap_res2.t2 GNDA 0.340442f
C1342 bgr_0.cap_res2.n0 GNDA 0.24022f
C1343 bgr_0.cap_res2.t3 GNDA 0.1913f
C1344 bgr_0.cap_res2.n1 GNDA 0.260644f
C1345 bgr_0.cap_res2.t10 GNDA 0.1913f
C1346 bgr_0.cap_res2.n2 GNDA 0.260644f
C1347 bgr_0.cap_res2.t17 GNDA 0.1913f
C1348 bgr_0.cap_res2.n3 GNDA 0.260644f
C1349 bgr_0.cap_res2.t12 GNDA 0.1913f
C1350 bgr_0.cap_res2.n4 GNDA 0.260644f
C1351 bgr_0.cap_res2.t18 GNDA 0.373116f
C1352 bgr_0.cap_res2.t0 GNDA 0.086426f
C1353 bgr_0.1st_Vout_2.n0 GNDA 0.569806f
C1354 bgr_0.1st_Vout_2.n1 GNDA 0.252461f
C1355 bgr_0.1st_Vout_2.n2 GNDA 1.43086f
C1356 bgr_0.1st_Vout_2.n3 GNDA 0.104399f
C1357 bgr_0.1st_Vout_2.n4 GNDA 1.45767f
C1358 bgr_0.1st_Vout_2.t33 GNDA 0.017308f
C1359 bgr_0.1st_Vout_2.t28 GNDA 0.288462f
C1360 bgr_0.1st_Vout_2.t17 GNDA 0.293375f
C1361 bgr_0.1st_Vout_2.t12 GNDA 0.288462f
C1362 bgr_0.1st_Vout_2.t32 GNDA 0.288462f
C1363 bgr_0.1st_Vout_2.t35 GNDA 0.293375f
C1364 bgr_0.1st_Vout_2.t11 GNDA 0.293375f
C1365 bgr_0.1st_Vout_2.t31 GNDA 0.288462f
C1366 bgr_0.1st_Vout_2.t23 GNDA 0.288462f
C1367 bgr_0.1st_Vout_2.t26 GNDA 0.293375f
C1368 bgr_0.1st_Vout_2.t30 GNDA 0.293375f
C1369 bgr_0.1st_Vout_2.t22 GNDA 0.288462f
C1370 bgr_0.1st_Vout_2.t15 GNDA 0.288462f
C1371 bgr_0.1st_Vout_2.t19 GNDA 0.293375f
C1372 bgr_0.1st_Vout_2.t36 GNDA 0.293375f
C1373 bgr_0.1st_Vout_2.t29 GNDA 0.288462f
C1374 bgr_0.1st_Vout_2.t21 GNDA 0.288462f
C1375 bgr_0.1st_Vout_2.t25 GNDA 0.293375f
C1376 bgr_0.1st_Vout_2.t18 GNDA 0.293375f
C1377 bgr_0.1st_Vout_2.t14 GNDA 0.288462f
C1378 bgr_0.1st_Vout_2.t20 GNDA 0.288462f
C1379 bgr_0.1st_Vout_2.t34 GNDA 0.018845f
C1380 bgr_0.1st_Vout_2.n5 GNDA 0.018179f
C1381 bgr_0.1st_Vout_2.t27 GNDA 0.010986f
C1382 bgr_0.1st_Vout_2.t16 GNDA 0.010986f
C1383 bgr_0.1st_Vout_2.n6 GNDA 0.024439f
C1384 bgr_0.1st_Vout_2.n7 GNDA 0.010417f
C1385 bgr_0.1st_Vout_2.t3 GNDA 0.015189f
C1386 bgr_0.1st_Vout_2.n8 GNDA 0.157567f
C1387 bgr_0.1st_Vout_2.n10 GNDA 0.017425f
C1388 bgr_0.1st_Vout_2.t24 GNDA 0.010986f
C1389 bgr_0.1st_Vout_2.t13 GNDA 0.010986f
C1390 bgr_0.1st_Vout_2.n11 GNDA 0.024439f
C1391 bgr_0.1st_Vout_2.n12 GNDA 0.138311f
C1392 bgr_0.1st_Vout_2.n13 GNDA 0.018179f
C1393 bgr_0.1st_Vout_1.n0 GNDA 0.538712f
C1394 bgr_0.1st_Vout_1.n1 GNDA 0.236313f
C1395 bgr_0.1st_Vout_1.n2 GNDA 0.973284f
C1396 bgr_0.1st_Vout_1.n3 GNDA 0.907198f
C1397 bgr_0.1st_Vout_1.n4 GNDA 0.891647f
C1398 bgr_0.1st_Vout_1.t11 GNDA 0.358463f
C1399 bgr_0.1st_Vout_1.t15 GNDA 0.35246f
C1400 bgr_0.1st_Vout_1.t29 GNDA 0.358463f
C1401 bgr_0.1st_Vout_1.t35 GNDA 0.35246f
C1402 bgr_0.1st_Vout_1.t31 GNDA 0.358463f
C1403 bgr_0.1st_Vout_1.t34 GNDA 0.35246f
C1404 bgr_0.1st_Vout_1.t20 GNDA 0.358463f
C1405 bgr_0.1st_Vout_1.t28 GNDA 0.35246f
C1406 bgr_0.1st_Vout_1.t24 GNDA 0.358463f
C1407 bgr_0.1st_Vout_1.t27 GNDA 0.35246f
C1408 bgr_0.1st_Vout_1.t14 GNDA 0.358463f
C1409 bgr_0.1st_Vout_1.t19 GNDA 0.35246f
C1410 bgr_0.1st_Vout_1.t30 GNDA 0.358463f
C1411 bgr_0.1st_Vout_1.t33 GNDA 0.35246f
C1412 bgr_0.1st_Vout_1.t18 GNDA 0.358463f
C1413 bgr_0.1st_Vout_1.t26 GNDA 0.35246f
C1414 bgr_0.1st_Vout_1.t23 GNDA 0.358463f
C1415 bgr_0.1st_Vout_1.t25 GNDA 0.35246f
C1416 bgr_0.1st_Vout_1.t17 GNDA 0.35246f
C1417 bgr_0.1st_Vout_1.t12 GNDA 0.35246f
C1418 bgr_0.1st_Vout_1.t21 GNDA 0.023025f
C1419 bgr_0.1st_Vout_1.n5 GNDA 0.715456f
C1420 bgr_0.1st_Vout_1.n6 GNDA 0.022212f
C1421 bgr_0.1st_Vout_1.n7 GNDA 0.104674f
C1422 bgr_0.1st_Vout_1.t36 GNDA 0.013423f
C1423 bgr_0.1st_Vout_1.t16 GNDA 0.013423f
C1424 bgr_0.1st_Vout_1.n8 GNDA 0.029862f
C1425 bgr_0.1st_Vout_1.n9 GNDA 0.082514f
C1426 bgr_0.1st_Vout_1.t7 GNDA 0.018559f
C1427 bgr_0.1st_Vout_1.n10 GNDA 0.012728f
C1428 bgr_0.1st_Vout_1.n11 GNDA 0.192525f
C1429 bgr_0.1st_Vout_1.n12 GNDA 0.011517f
C1430 bgr_0.1st_Vout_1.n13 GNDA 0.048842f
C1431 bgr_0.1st_Vout_1.n14 GNDA 0.021291f
C1432 bgr_0.1st_Vout_1.n15 GNDA 0.078719f
C1433 bgr_0.1st_Vout_1.n16 GNDA 0.038771f
C1434 bgr_0.1st_Vout_1.t32 GNDA 0.013423f
C1435 bgr_0.1st_Vout_1.t22 GNDA 0.013423f
C1436 bgr_0.1st_Vout_1.n17 GNDA 0.029862f
C1437 bgr_0.1st_Vout_1.n18 GNDA 0.082514f
C1438 bgr_0.1st_Vout_1.n19 GNDA 0.022212f
C1439 bgr_0.1st_Vout_1.n20 GNDA 0.104674f
C1440 bgr_0.1st_Vout_1.t13 GNDA 0.021069f
C1441 bgr_0.V_mir1.t11 GNDA 0.019293f
C1442 bgr_0.V_mir1.t4 GNDA 0.02939f
C1443 bgr_0.V_mir1.t8 GNDA 0.023151f
C1444 bgr_0.V_mir1.t18 GNDA 0.023151f
C1445 bgr_0.V_mir1.t20 GNDA 0.037369f
C1446 bgr_0.V_mir1.n0 GNDA 0.041731f
C1447 bgr_0.V_mir1.n1 GNDA 0.028507f
C1448 bgr_0.V_mir1.n2 GNDA 0.044354f
C1449 bgr_0.V_mir1.t5 GNDA 0.019293f
C1450 bgr_0.V_mir1.t9 GNDA 0.019293f
C1451 bgr_0.V_mir1.n3 GNDA 0.044166f
C1452 bgr_0.V_mir1.n4 GNDA 0.109943f
C1453 bgr_0.V_mir1.n5 GNDA 0.025223f
C1454 bgr_0.V_mir1.t0 GNDA 0.041163f
C1455 bgr_0.V_mir1.n6 GNDA 0.027381f
C1456 bgr_0.V_mir1.n7 GNDA 0.451535f
C1457 bgr_0.V_mir1.n8 GNDA 0.146338f
C1458 bgr_0.V_mir1.t6 GNDA 0.02939f
C1459 bgr_0.V_mir1.t12 GNDA 0.023151f
C1460 bgr_0.V_mir1.t17 GNDA 0.023151f
C1461 bgr_0.V_mir1.t21 GNDA 0.037369f
C1462 bgr_0.V_mir1.n9 GNDA 0.041731f
C1463 bgr_0.V_mir1.n10 GNDA 0.028507f
C1464 bgr_0.V_mir1.n11 GNDA 0.044354f
C1465 bgr_0.V_mir1.t7 GNDA 0.019293f
C1466 bgr_0.V_mir1.t13 GNDA 0.019293f
C1467 bgr_0.V_mir1.n12 GNDA 0.044166f
C1468 bgr_0.V_mir1.n13 GNDA 0.085095f
C1469 bgr_0.V_mir1.n14 GNDA 0.051125f
C1470 bgr_0.V_mir1.n15 GNDA 0.381359f
C1471 bgr_0.V_mir1.t10 GNDA 0.02939f
C1472 bgr_0.V_mir1.t14 GNDA 0.023151f
C1473 bgr_0.V_mir1.t22 GNDA 0.023151f
C1474 bgr_0.V_mir1.t19 GNDA 0.037369f
C1475 bgr_0.V_mir1.n16 GNDA 0.041731f
C1476 bgr_0.V_mir1.n17 GNDA 0.028507f
C1477 bgr_0.V_mir1.n18 GNDA 0.044354f
C1478 bgr_0.V_mir1.n19 GNDA 0.111042f
C1479 bgr_0.V_mir1.n20 GNDA 0.044166f
C1480 bgr_0.V_mir1.t15 GNDA 0.019293f
C1481 bgr_0.Vin+.t7 GNDA 0.010696f
C1482 bgr_0.Vin+.t8 GNDA 0.025367f
C1483 bgr_0.Vin+.t9 GNDA 0.01649f
C1484 bgr_0.Vin+.n0 GNDA 0.054406f
C1485 bgr_0.Vin+.t6 GNDA 0.01649f
C1486 bgr_0.Vin+.n1 GNDA 0.042338f
C1487 bgr_0.Vin+.t10 GNDA 0.01649f
C1488 bgr_0.Vin+.n2 GNDA 0.042909f
C1489 bgr_0.Vin+.n3 GNDA 0.130793f
C1490 bgr_0.Vin+.t2 GNDA 0.05348f
C1491 bgr_0.Vin+.t1 GNDA 0.05348f
C1492 bgr_0.Vin+.n4 GNDA 0.17668f
C1493 bgr_0.Vin+.n5 GNDA 1.27851f
C1494 bgr_0.Vin+.t0 GNDA 0.05348f
C1495 bgr_0.Vin+.t3 GNDA 0.05348f
C1496 bgr_0.Vin+.n6 GNDA 0.17668f
C1497 bgr_0.Vin+.n7 GNDA 1.06526f
C1498 bgr_0.Vin+.t5 GNDA 0.232527f
C1499 bgr_0.Vin+.n8 GNDA 1.7265f
C1500 bgr_0.Vin+.t4 GNDA 0.173951f
C1501 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t3 GNDA 0.01464f
C1502 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t16 GNDA 0.01464f
C1503 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n0 GNDA 0.036714f
C1504 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t4 GNDA 0.01464f
C1505 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t1 GNDA 0.01464f
C1506 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n1 GNDA 0.03652f
C1507 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n2 GNDA 0.324652f
C1508 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t15 GNDA 0.01464f
C1509 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t2 GNDA 0.01464f
C1510 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n3 GNDA 0.02928f
C1511 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n4 GNDA 0.05443f
C1512 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t0 GNDA 0.187219f
C1513 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n5 GNDA 0.046248f
C1514 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n6 GNDA 0.081804f
C1515 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t9 GNDA 0.02928f
C1516 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t5 GNDA 0.02928f
C1517 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n7 GNDA 0.059867f
C1518 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n8 GNDA 0.20109f
C1519 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t8 GNDA 0.02928f
C1520 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t14 GNDA 0.02928f
C1521 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n9 GNDA 0.059867f
C1522 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n10 GNDA 0.193651f
C1523 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n11 GNDA 0.078635f
C1524 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n12 GNDA 0.046248f
C1525 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t12 GNDA 0.02928f
C1526 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t7 GNDA 0.02928f
C1527 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n13 GNDA 0.059867f
C1528 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n14 GNDA 0.193651f
C1529 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n15 GNDA 0.047939f
C1530 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t11 GNDA 0.02928f
C1531 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t6 GNDA 0.02928f
C1532 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n16 GNDA 0.059867f
C1533 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n17 GNDA 0.193651f
C1534 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n18 GNDA 0.081804f
C1535 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t10 GNDA 0.02928f
C1536 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.t13 GNDA 0.02928f
C1537 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n19 GNDA 0.059867f
C1538 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n20 GNDA 0.197477f
C1539 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n21 GNDA 0.119373f
C1540 two_stage_opamp_dummy_magic_21_0.V_CMFB_S3.n22 GNDA 1.32714f
C1541 bgr_0.V_CMFB_S3 GNDA 0.84249f
C1542 two_stage_opamp_dummy_magic_21_0.Y.t6 GNDA 0.037911f
C1543 two_stage_opamp_dummy_magic_21_0.Y.t5 GNDA 0.037911f
C1544 two_stage_opamp_dummy_magic_21_0.Y.n0 GNDA 0.082489f
C1545 two_stage_opamp_dummy_magic_21_0.Y.n1 GNDA 0.256901f
C1546 two_stage_opamp_dummy_magic_21_0.Y.n2 GNDA 0.080625f
C1547 two_stage_opamp_dummy_magic_21_0.Y.t1 GNDA 0.037911f
C1548 two_stage_opamp_dummy_magic_21_0.Y.t19 GNDA 0.037911f
C1549 two_stage_opamp_dummy_magic_21_0.Y.n3 GNDA 0.082489f
C1550 two_stage_opamp_dummy_magic_21_0.Y.n4 GNDA 0.327754f
C1551 two_stage_opamp_dummy_magic_21_0.Y.t18 GNDA 0.037911f
C1552 two_stage_opamp_dummy_magic_21_0.Y.t22 GNDA 0.037911f
C1553 two_stage_opamp_dummy_magic_21_0.Y.n5 GNDA 0.082489f
C1554 two_stage_opamp_dummy_magic_21_0.Y.n6 GNDA 0.327754f
C1555 two_stage_opamp_dummy_magic_21_0.Y.n7 GNDA 0.137048f
C1556 two_stage_opamp_dummy_magic_21_0.Y.t4 GNDA 0.037911f
C1557 two_stage_opamp_dummy_magic_21_0.Y.t23 GNDA 0.037911f
C1558 two_stage_opamp_dummy_magic_21_0.Y.n8 GNDA 0.082489f
C1559 two_stage_opamp_dummy_magic_21_0.Y.n9 GNDA 0.314545f
C1560 two_stage_opamp_dummy_magic_21_0.Y.n10 GNDA 0.144975f
C1561 two_stage_opamp_dummy_magic_21_0.Y.t20 GNDA 0.037911f
C1562 two_stage_opamp_dummy_magic_21_0.Y.t0 GNDA 0.037911f
C1563 two_stage_opamp_dummy_magic_21_0.Y.n11 GNDA 0.082489f
C1564 two_stage_opamp_dummy_magic_21_0.Y.n12 GNDA 0.314545f
C1565 two_stage_opamp_dummy_magic_21_0.Y.n13 GNDA 0.084683f
C1566 two_stage_opamp_dummy_magic_21_0.Y.n14 GNDA 0.084683f
C1567 two_stage_opamp_dummy_magic_21_0.Y.n15 GNDA 0.144975f
C1568 two_stage_opamp_dummy_magic_21_0.Y.t12 GNDA 0.037911f
C1569 two_stage_opamp_dummy_magic_21_0.Y.t10 GNDA 0.037911f
C1570 two_stage_opamp_dummy_magic_21_0.Y.n16 GNDA 0.082489f
C1571 two_stage_opamp_dummy_magic_21_0.Y.n17 GNDA 0.314545f
C1572 two_stage_opamp_dummy_magic_21_0.Y.n18 GNDA 0.137048f
C1573 two_stage_opamp_dummy_magic_21_0.Y.n19 GNDA 0.075821f
C1574 two_stage_opamp_dummy_magic_21_0.Y.n20 GNDA 0.3074f
C1575 two_stage_opamp_dummy_magic_21_0.Y.t8 GNDA 0.088458f
C1576 two_stage_opamp_dummy_magic_21_0.Y.t13 GNDA 0.088458f
C1577 two_stage_opamp_dummy_magic_21_0.Y.n21 GNDA 0.180951f
C1578 two_stage_opamp_dummy_magic_21_0.Y.n22 GNDA 0.492191f
C1579 two_stage_opamp_dummy_magic_21_0.Y.n23 GNDA 0.095948f
C1580 two_stage_opamp_dummy_magic_21_0.Y.n24 GNDA 0.163678f
C1581 two_stage_opamp_dummy_magic_21_0.Y.t11 GNDA 0.088458f
C1582 two_stage_opamp_dummy_magic_21_0.Y.t2 GNDA 0.088458f
C1583 two_stage_opamp_dummy_magic_21_0.Y.n25 GNDA 0.180951f
C1584 two_stage_opamp_dummy_magic_21_0.Y.n26 GNDA 0.585864f
C1585 two_stage_opamp_dummy_magic_21_0.Y.t16 GNDA 0.088458f
C1586 two_stage_opamp_dummy_magic_21_0.Y.t7 GNDA 0.088458f
C1587 two_stage_opamp_dummy_magic_21_0.Y.n27 GNDA 0.180951f
C1588 two_stage_opamp_dummy_magic_21_0.Y.n28 GNDA 0.569865f
C1589 two_stage_opamp_dummy_magic_21_0.Y.n29 GNDA 0.163678f
C1590 two_stage_opamp_dummy_magic_21_0.Y.n30 GNDA 0.095948f
C1591 two_stage_opamp_dummy_magic_21_0.Y.t9 GNDA 0.088458f
C1592 two_stage_opamp_dummy_magic_21_0.Y.t14 GNDA 0.088458f
C1593 two_stage_opamp_dummy_magic_21_0.Y.n31 GNDA 0.180951f
C1594 two_stage_opamp_dummy_magic_21_0.Y.n32 GNDA 0.569865f
C1595 two_stage_opamp_dummy_magic_21_0.Y.n33 GNDA 0.095948f
C1596 two_stage_opamp_dummy_magic_21_0.Y.t15 GNDA 0.088458f
C1597 two_stage_opamp_dummy_magic_21_0.Y.t17 GNDA 0.088458f
C1598 two_stage_opamp_dummy_magic_21_0.Y.n34 GNDA 0.180951f
C1599 two_stage_opamp_dummy_magic_21_0.Y.n35 GNDA 0.569865f
C1600 two_stage_opamp_dummy_magic_21_0.Y.n36 GNDA 0.095948f
C1601 two_stage_opamp_dummy_magic_21_0.Y.n37 GNDA 0.163678f
C1602 two_stage_opamp_dummy_magic_21_0.Y.t24 GNDA 0.088458f
C1603 two_stage_opamp_dummy_magic_21_0.Y.t3 GNDA 0.088458f
C1604 two_stage_opamp_dummy_magic_21_0.Y.n38 GNDA 0.180951f
C1605 two_stage_opamp_dummy_magic_21_0.Y.n39 GNDA 0.569865f
C1606 two_stage_opamp_dummy_magic_21_0.Y.n40 GNDA 0.149208f
C1607 two_stage_opamp_dummy_magic_21_0.Y.n41 GNDA 0.48498f
C1608 two_stage_opamp_dummy_magic_21_0.Y.t41 GNDA 0.053075f
C1609 two_stage_opamp_dummy_magic_21_0.Y.t25 GNDA 0.053075f
C1610 two_stage_opamp_dummy_magic_21_0.Y.t32 GNDA 0.053075f
C1611 two_stage_opamp_dummy_magic_21_0.Y.t50 GNDA 0.053075f
C1612 two_stage_opamp_dummy_magic_21_0.Y.t34 GNDA 0.053075f
C1613 two_stage_opamp_dummy_magic_21_0.Y.t51 GNDA 0.053075f
C1614 two_stage_opamp_dummy_magic_21_0.Y.t37 GNDA 0.053075f
C1615 two_stage_opamp_dummy_magic_21_0.Y.t30 GNDA 0.064448f
C1616 two_stage_opamp_dummy_magic_21_0.Y.n42 GNDA 0.064448f
C1617 two_stage_opamp_dummy_magic_21_0.Y.n43 GNDA 0.041702f
C1618 two_stage_opamp_dummy_magic_21_0.Y.n44 GNDA 0.041702f
C1619 two_stage_opamp_dummy_magic_21_0.Y.n45 GNDA 0.041702f
C1620 two_stage_opamp_dummy_magic_21_0.Y.n46 GNDA 0.041702f
C1621 two_stage_opamp_dummy_magic_21_0.Y.n47 GNDA 0.041702f
C1622 two_stage_opamp_dummy_magic_21_0.Y.n48 GNDA 0.033646f
C1623 two_stage_opamp_dummy_magic_21_0.Y.t53 GNDA 0.053075f
C1624 two_stage_opamp_dummy_magic_21_0.Y.t38 GNDA 0.064448f
C1625 two_stage_opamp_dummy_magic_21_0.Y.n49 GNDA 0.056392f
C1626 two_stage_opamp_dummy_magic_21_0.Y.n50 GNDA 0.021219f
C1627 two_stage_opamp_dummy_magic_21_0.Y.t46 GNDA 0.081508f
C1628 two_stage_opamp_dummy_magic_21_0.Y.t29 GNDA 0.081508f
C1629 two_stage_opamp_dummy_magic_21_0.Y.t36 GNDA 0.081508f
C1630 two_stage_opamp_dummy_magic_21_0.Y.t52 GNDA 0.081508f
C1631 two_stage_opamp_dummy_magic_21_0.Y.t40 GNDA 0.081508f
C1632 two_stage_opamp_dummy_magic_21_0.Y.t54 GNDA 0.081508f
C1633 two_stage_opamp_dummy_magic_21_0.Y.t43 GNDA 0.081508f
C1634 two_stage_opamp_dummy_magic_21_0.Y.t35 GNDA 0.092661f
C1635 two_stage_opamp_dummy_magic_21_0.Y.n51 GNDA 0.083624f
C1636 two_stage_opamp_dummy_magic_21_0.Y.n52 GNDA 0.05118f
C1637 two_stage_opamp_dummy_magic_21_0.Y.n53 GNDA 0.05118f
C1638 two_stage_opamp_dummy_magic_21_0.Y.n54 GNDA 0.05118f
C1639 two_stage_opamp_dummy_magic_21_0.Y.n55 GNDA 0.05118f
C1640 two_stage_opamp_dummy_magic_21_0.Y.n56 GNDA 0.05118f
C1641 two_stage_opamp_dummy_magic_21_0.Y.n57 GNDA 0.043123f
C1642 two_stage_opamp_dummy_magic_21_0.Y.t27 GNDA 0.081508f
C1643 two_stage_opamp_dummy_magic_21_0.Y.t44 GNDA 0.092661f
C1644 two_stage_opamp_dummy_magic_21_0.Y.n58 GNDA 0.075568f
C1645 two_stage_opamp_dummy_magic_21_0.Y.n59 GNDA 0.021219f
C1646 two_stage_opamp_dummy_magic_21_0.Y.n60 GNDA 0.091639f
C1647 two_stage_opamp_dummy_magic_21_0.Y.n61 GNDA 1.04027f
C1648 two_stage_opamp_dummy_magic_21_0.Y.n62 GNDA 0.450882f
C1649 two_stage_opamp_dummy_magic_21_0.Y.t28 GNDA 0.166807f
C1650 two_stage_opamp_dummy_magic_21_0.Y.t47 GNDA 0.166807f
C1651 two_stage_opamp_dummy_magic_21_0.Y.t39 GNDA 0.177661f
C1652 two_stage_opamp_dummy_magic_21_0.Y.n63 GNDA 0.140789f
C1653 two_stage_opamp_dummy_magic_21_0.Y.n64 GNDA 0.071557f
C1654 two_stage_opamp_dummy_magic_21_0.Y.t45 GNDA 0.166807f
C1655 two_stage_opamp_dummy_magic_21_0.Y.t26 GNDA 0.166807f
C1656 two_stage_opamp_dummy_magic_21_0.Y.t42 GNDA 0.166807f
C1657 two_stage_opamp_dummy_magic_21_0.Y.t33 GNDA 0.166807f
C1658 two_stage_opamp_dummy_magic_21_0.Y.t49 GNDA 0.166807f
C1659 two_stage_opamp_dummy_magic_21_0.Y.t31 GNDA 0.166807f
C1660 two_stage_opamp_dummy_magic_21_0.Y.t48 GNDA 0.177661f
C1661 two_stage_opamp_dummy_magic_21_0.Y.n65 GNDA 0.140789f
C1662 two_stage_opamp_dummy_magic_21_0.Y.n66 GNDA 0.079613f
C1663 two_stage_opamp_dummy_magic_21_0.Y.n67 GNDA 0.079613f
C1664 two_stage_opamp_dummy_magic_21_0.Y.n68 GNDA 0.079613f
C1665 two_stage_opamp_dummy_magic_21_0.Y.n69 GNDA 0.079613f
C1666 two_stage_opamp_dummy_magic_21_0.Y.n70 GNDA 0.071557f
C1667 two_stage_opamp_dummy_magic_21_0.Y.n71 GNDA 0.036197f
C1668 two_stage_opamp_dummy_magic_21_0.Y.n72 GNDA 1.26467f
C1669 two_stage_opamp_dummy_magic_21_0.Y.t21 GNDA 1.21199f
C1670 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t21 GNDA 0.014491f
C1671 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t10 GNDA 0.014491f
C1672 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t16 GNDA 0.014491f
C1673 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t9 GNDA 0.014491f
C1674 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t15 GNDA 0.014491f
C1675 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t12 GNDA 0.014491f
C1676 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t17 GNDA 0.014491f
C1677 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t13 GNDA 0.014491f
C1678 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t7 GNDA 0.014491f
C1679 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t8 GNDA 0.044454f
C1680 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n0 GNDA 0.06039f
C1681 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n1 GNDA 0.048586f
C1682 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n2 GNDA 0.048586f
C1683 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n3 GNDA 0.28612f
C1684 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n4 GNDA 0.28612f
C1685 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n5 GNDA 0.048586f
C1686 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n6 GNDA 0.048586f
C1687 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n7 GNDA 0.048586f
C1688 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n8 GNDA 0.07225f
C1689 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t6 GNDA 0.359564f
C1690 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t18 GNDA 0.056228f
C1691 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t11 GNDA 0.021026f
C1692 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n9 GNDA 0.065948f
C1693 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t20 GNDA 0.021026f
C1694 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n10 GNDA 0.053985f
C1695 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t14 GNDA 0.021026f
C1696 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n11 GNDA 0.053985f
C1697 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t19 GNDA 0.021026f
C1698 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n12 GNDA 0.093575f
C1699 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n13 GNDA 1.87082f
C1700 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t5 GNDA 0.068191f
C1701 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t2 GNDA 0.068191f
C1702 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n14 GNDA 0.240167f
C1703 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t3 GNDA 0.068191f
C1704 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t1 GNDA 0.068191f
C1705 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n15 GNDA 0.22851f
C1706 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n16 GNDA 1.0679f
C1707 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t0 GNDA 0.068191f
C1708 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.t4 GNDA 0.068191f
C1709 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n17 GNDA 0.22851f
C1710 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n18 GNDA 0.763632f
C1711 two_stage_opamp_dummy_magic_21_0.V_err_amp_ref.n19 GNDA 1.56767f
C1712 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t1 GNDA 0.343734f
C1713 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t75 GNDA 0.344881f
C1714 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t37 GNDA 0.185242f
C1715 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n0 GNDA 0.197802f
C1716 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t36 GNDA 0.343734f
C1717 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t119 GNDA 0.344881f
C1718 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t74 GNDA 0.185242f
C1719 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n1 GNDA 0.216311f
C1720 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t22 GNDA 0.343734f
C1721 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t97 GNDA 0.344881f
C1722 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t59 GNDA 0.185242f
C1723 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n2 GNDA 0.216311f
C1724 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t54 GNDA 0.343734f
C1725 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t130 GNDA 0.344881f
C1726 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t93 GNDA 0.185242f
C1727 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n3 GNDA 0.216311f
C1728 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t91 GNDA 0.343734f
C1729 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t42 GNDA 0.344881f
C1730 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t135 GNDA 0.36339f
C1731 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t30 GNDA 0.36339f
C1732 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t129 GNDA 0.185242f
C1733 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n4 GNDA 0.216311f
C1734 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t69 GNDA 0.343734f
C1735 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t94 GNDA 0.344881f
C1736 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t115 GNDA 0.36339f
C1737 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t13 GNDA 0.36339f
C1738 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t111 GNDA 0.185242f
C1739 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n5 GNDA 0.216311f
C1740 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t116 GNDA 0.344881f
C1741 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t137 GNDA 0.346131f
C1742 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t71 GNDA 0.344881f
C1743 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t99 GNDA 0.347585f
C1744 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t60 GNDA 0.378048f
C1745 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t122 GNDA 0.344881f
C1746 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t104 GNDA 0.346131f
C1747 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t20 GNDA 0.344881f
C1748 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t35 GNDA 0.346131f
C1749 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t86 GNDA 0.344881f
C1750 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t67 GNDA 0.346131f
C1751 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t120 GNDA 0.344881f
C1752 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t5 GNDA 0.346131f
C1753 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t61 GNDA 0.344881f
C1754 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t113 GNDA 0.346131f
C1755 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t90 GNDA 0.344881f
C1756 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t38 GNDA 0.346131f
C1757 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t101 GNDA 0.344881f
C1758 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t15 GNDA 0.346131f
C1759 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t127 GNDA 0.344881f
C1760 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t76 GNDA 0.346131f
C1761 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t65 GNDA 0.344881f
C1762 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t117 GNDA 0.346131f
C1763 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t98 GNDA 0.344881f
C1764 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t47 GNDA 0.346131f
C1765 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t107 GNDA 0.344881f
C1766 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t21 GNDA 0.346131f
C1767 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t136 GNDA 0.344881f
C1768 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t84 GNDA 0.346131f
C1769 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t8 GNDA 0.344881f
C1770 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t57 GNDA 0.346131f
C1771 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t34 GNDA 0.344881f
C1772 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t123 GNDA 0.346131f
C1773 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t112 GNDA 0.344881f
C1774 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t23 GNDA 0.346131f
C1775 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t4 GNDA 0.344881f
C1776 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t89 GNDA 0.346131f
C1777 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t14 GNDA 0.344881f
C1778 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t62 GNDA 0.346131f
C1779 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t40 GNDA 0.344881f
C1780 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t126 GNDA 0.346131f
C1781 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t51 GNDA 0.344881f
C1782 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t103 GNDA 0.346131f
C1783 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t79 GNDA 0.344881f
C1784 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t29 GNDA 0.346131f
C1785 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t87 GNDA 0.344881f
C1786 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t2 GNDA 0.346131f
C1787 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t121 GNDA 0.344881f
C1788 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t70 GNDA 0.346131f
C1789 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t56 GNDA 0.344881f
C1790 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t109 GNDA 0.346131f
C1791 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t85 GNDA 0.344881f
C1792 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t33 GNDA 0.346131f
C1793 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t95 GNDA 0.344881f
C1794 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t9 GNDA 0.346131f
C1795 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t124 GNDA 0.344881f
C1796 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t73 GNDA 0.346131f
C1797 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t132 GNDA 0.344881f
C1798 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t43 GNDA 0.346131f
C1799 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t27 GNDA 0.344881f
C1800 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t118 GNDA 0.346131f
C1801 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t6 GNDA 0.344881f
C1802 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t68 GNDA 0.36179f
C1803 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t92 GNDA 0.344881f
C1804 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t105 GNDA 0.185242f
C1805 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n6 GNDA 0.198255f
C1806 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t133 GNDA 0.344881f
C1807 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t19 GNDA 0.185242f
C1808 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n7 GNDA 0.196656f
C1809 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t82 GNDA 0.344881f
C1810 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t50 GNDA 0.185242f
C1811 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n8 GNDA 0.196656f
C1812 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t31 GNDA 0.344881f
C1813 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t81 GNDA 0.185242f
C1814 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n9 GNDA 0.196656f
C1815 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t72 GNDA 0.344881f
C1816 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t131 GNDA 0.185242f
C1817 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n10 GNDA 0.196656f
C1818 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t26 GNDA 0.344881f
C1819 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t28 GNDA 0.185242f
C1820 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n11 GNDA 0.196656f
C1821 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t114 GNDA 0.344881f
C1822 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t66 GNDA 0.185242f
C1823 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n12 GNDA 0.196656f
C1824 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t64 GNDA 0.344881f
C1825 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t102 GNDA 0.185242f
C1826 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n13 GNDA 0.196656f
C1827 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t108 GNDA 0.344881f
C1828 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t16 GNDA 0.185242f
C1829 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n14 GNDA 0.196656f
C1830 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t128 GNDA 0.344881f
C1831 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t77 GNDA 0.346131f
C1832 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t48 GNDA 0.344881f
C1833 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t7 GNDA 0.346131f
C1834 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t55 GNDA 0.166734f
C1835 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n15 GNDA 0.215061f
C1836 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t46 GNDA 0.184096f
C1837 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n16 GNDA 0.23357f
C1838 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t78 GNDA 0.184096f
C1839 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n17 GNDA 0.250829f
C1840 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t39 GNDA 0.184096f
C1841 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n18 GNDA 0.250829f
C1842 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t3 GNDA 0.184096f
C1843 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n19 GNDA 0.250829f
C1844 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t32 GNDA 0.184096f
C1845 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n20 GNDA 0.250829f
C1846 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t134 GNDA 0.184096f
C1847 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n21 GNDA 0.250829f
C1848 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t96 GNDA 0.184096f
C1849 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n22 GNDA 0.250829f
C1850 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t58 GNDA 0.184096f
C1851 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n23 GNDA 0.250829f
C1852 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t88 GNDA 0.184096f
C1853 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n24 GNDA 0.250829f
C1854 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t53 GNDA 0.184096f
C1855 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n25 GNDA 0.250829f
C1856 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t17 GNDA 0.184096f
C1857 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n26 GNDA 0.250829f
C1858 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t45 GNDA 0.184096f
C1859 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n27 GNDA 0.250829f
C1860 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t11 GNDA 0.184096f
C1861 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n28 GNDA 0.250829f
C1862 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t106 GNDA 0.184096f
C1863 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n29 GNDA 0.250829f
C1864 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t0 GNDA 0.184096f
C1865 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n30 GNDA 0.250829f
C1866 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t100 GNDA 0.184096f
C1867 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n31 GNDA 0.23357f
C1868 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t24 GNDA 0.343734f
C1869 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t63 GNDA 0.166734f
C1870 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n32 GNDA 0.216311f
C1871 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t41 GNDA 0.343734f
C1872 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t80 GNDA 0.166734f
C1873 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n33 GNDA 0.216311f
C1874 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t10 GNDA 0.343734f
C1875 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t25 GNDA 0.344881f
C1876 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t52 GNDA 0.36339f
C1877 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t83 GNDA 0.36339f
C1878 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t44 GNDA 0.185242f
C1879 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n34 GNDA 0.216311f
C1880 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t110 GNDA 0.343734f
C1881 two_stage_opamp_dummy_magic_21_0.cap_res_Y.n35 GNDA 0.216311f
C1882 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t12 GNDA 0.185242f
C1883 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t49 GNDA 0.36339f
C1884 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t18 GNDA 0.36339f
C1885 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t125 GNDA 0.434792f
C1886 two_stage_opamp_dummy_magic_21_0.cap_res_Y.t138 GNDA 0.291879f
C1887 VOUT+.n0 GNDA 0.084549f
C1888 VOUT+.t16 GNDA 0.05596f
C1889 VOUT+.t13 GNDA 0.05596f
C1890 VOUT+.n1 GNDA 0.120236f
C1891 VOUT+.n2 GNDA 0.33616f
C1892 VOUT+.t11 GNDA 0.05596f
C1893 VOUT+.t10 GNDA 0.05596f
C1894 VOUT+.n3 GNDA 0.120236f
C1895 VOUT+.n4 GNDA 0.323898f
C1896 VOUT+.n5 GNDA 0.117363f
C1897 VOUT+.t12 GNDA 0.05596f
C1898 VOUT+.t15 GNDA 0.05596f
C1899 VOUT+.n6 GNDA 0.120236f
C1900 VOUT+.n7 GNDA 0.330029f
C1901 VOUT+.n8 GNDA 0.060929f
C1902 VOUT+.t9 GNDA 0.092521f
C1903 VOUT+.n9 GNDA 0.113841f
C1904 VOUT+.t0 GNDA 0.047965f
C1905 VOUT+.t5 GNDA 0.047965f
C1906 VOUT+.n10 GNDA 0.098281f
C1907 VOUT+.n11 GNDA 0.251135f
C1908 VOUT+.t18 GNDA 0.047965f
C1909 VOUT+.t4 GNDA 0.047965f
C1910 VOUT+.n12 GNDA 0.098281f
C1911 VOUT+.n13 GNDA 0.292558f
C1912 VOUT+.n14 GNDA 0.034573f
C1913 VOUT+.n15 GNDA 0.060993f
C1914 VOUT+.t1 GNDA 0.047965f
C1915 VOUT+.t17 GNDA 0.047965f
C1916 VOUT+.n16 GNDA 0.098281f
C1917 VOUT+.n17 GNDA 0.292558f
C1918 VOUT+.n18 GNDA 0.060993f
C1919 VOUT+.t2 GNDA 0.047965f
C1920 VOUT+.t3 GNDA 0.047965f
C1921 VOUT+.n19 GNDA 0.098281f
C1922 VOUT+.n20 GNDA 0.287445f
C1923 VOUT+.n21 GNDA 0.060993f
C1924 VOUT+.t8 GNDA 0.047965f
C1925 VOUT+.t6 GNDA 0.047965f
C1926 VOUT+.n22 GNDA 0.098281f
C1927 VOUT+.n23 GNDA 0.287445f
C1928 VOUT+.n24 GNDA 0.034573f
C1929 VOUT+.n25 GNDA 0.034573f
C1930 VOUT+.t14 GNDA 0.047965f
C1931 VOUT+.t7 GNDA 0.047965f
C1932 VOUT+.n26 GNDA 0.098281f
C1933 VOUT+.n27 GNDA 0.287445f
C1934 VOUT+.n28 GNDA 0.034573f
C1935 VOUT+.n29 GNDA 0.050403f
C1936 VOUT+.n30 GNDA 0.200224f
C1937 VOUT+.t101 GNDA 0.319769f
C1938 VOUT+.t108 GNDA 0.325216f
C1939 VOUT+.t149 GNDA 0.319769f
C1940 VOUT+.n31 GNDA 0.214395f
C1941 VOUT+.n32 GNDA 0.139899f
C1942 VOUT+.t48 GNDA 0.324534f
C1943 VOUT+.t92 GNDA 0.324534f
C1944 VOUT+.t42 GNDA 0.324534f
C1945 VOUT+.t130 GNDA 0.324534f
C1946 VOUT+.t84 GNDA 0.324534f
C1947 VOUT+.t125 GNDA 0.324534f
C1948 VOUT+.t74 GNDA 0.324534f
C1949 VOUT+.t23 GNDA 0.324534f
C1950 VOUT+.t64 GNDA 0.324534f
C1951 VOUT+.t150 GNDA 0.324534f
C1952 VOUT+.t88 GNDA 0.319769f
C1953 VOUT+.n33 GNDA 0.215077f
C1954 VOUT+.t51 GNDA 0.319769f
C1955 VOUT+.n34 GNDA 0.275033f
C1956 VOUT+.t137 GNDA 0.319769f
C1957 VOUT+.n35 GNDA 0.275033f
C1958 VOUT+.t106 GNDA 0.319769f
C1959 VOUT+.n36 GNDA 0.275033f
C1960 VOUT+.t75 GNDA 0.319769f
C1961 VOUT+.n37 GNDA 0.275033f
C1962 VOUT+.t25 GNDA 0.319769f
C1963 VOUT+.n38 GNDA 0.275033f
C1964 VOUT+.t128 GNDA 0.319769f
C1965 VOUT+.n39 GNDA 0.275033f
C1966 VOUT+.t90 GNDA 0.319769f
C1967 VOUT+.n40 GNDA 0.275033f
C1968 VOUT+.t54 GNDA 0.319769f
C1969 VOUT+.n41 GNDA 0.275033f
C1970 VOUT+.t140 GNDA 0.319769f
C1971 VOUT+.n42 GNDA 0.275033f
C1972 VOUT+.t110 GNDA 0.319769f
C1973 VOUT+.t28 GNDA 0.325216f
C1974 VOUT+.t79 GNDA 0.319769f
C1975 VOUT+.n43 GNDA 0.214395f
C1976 VOUT+.n44 GNDA 0.259812f
C1977 VOUT+.t24 GNDA 0.325216f
C1978 VOUT+.t113 GNDA 0.319769f
C1979 VOUT+.n45 GNDA 0.214395f
C1980 VOUT+.t78 GNDA 0.319769f
C1981 VOUT+.t129 GNDA 0.325216f
C1982 VOUT+.t38 GNDA 0.319769f
C1983 VOUT+.n46 GNDA 0.214395f
C1984 VOUT+.n47 GNDA 0.259812f
C1985 VOUT+.t61 GNDA 0.325216f
C1986 VOUT+.t147 GNDA 0.319769f
C1987 VOUT+.n48 GNDA 0.214395f
C1988 VOUT+.t117 GNDA 0.319769f
C1989 VOUT+.t32 GNDA 0.325216f
C1990 VOUT+.t83 GNDA 0.319769f
C1991 VOUT+.n49 GNDA 0.214395f
C1992 VOUT+.n50 GNDA 0.259812f
C1993 VOUT+.t100 GNDA 0.325216f
C1994 VOUT+.t47 GNDA 0.319769f
C1995 VOUT+.n51 GNDA 0.214395f
C1996 VOUT+.t153 GNDA 0.319769f
C1997 VOUT+.t71 GNDA 0.325216f
C1998 VOUT+.t123 GNDA 0.319769f
C1999 VOUT+.n52 GNDA 0.214395f
C2000 VOUT+.n53 GNDA 0.259812f
C2001 VOUT+.t69 GNDA 0.325216f
C2002 VOUT+.t154 GNDA 0.319769f
C2003 VOUT+.n54 GNDA 0.214395f
C2004 VOUT+.t124 GNDA 0.319769f
C2005 VOUT+.t35 GNDA 0.325216f
C2006 VOUT+.t86 GNDA 0.319769f
C2007 VOUT+.n55 GNDA 0.214395f
C2008 VOUT+.n56 GNDA 0.259812f
C2009 VOUT+.t96 GNDA 0.319769f
C2010 VOUT+.t85 GNDA 0.325216f
C2011 VOUT+.t57 GNDA 0.319769f
C2012 VOUT+.n57 GNDA 0.214395f
C2013 VOUT+.n58 GNDA 0.139899f
C2014 VOUT+.t132 GNDA 0.324534f
C2015 VOUT+.t115 GNDA 0.324534f
C2016 VOUT+.t131 GNDA 0.325216f
C2017 VOUT+.t104 GNDA 0.319769f
C2018 VOUT+.n59 GNDA 0.214395f
C2019 VOUT+.t73 GNDA 0.319769f
C2020 VOUT+.n60 GNDA 0.134903f
C2021 VOUT+.t146 GNDA 0.324534f
C2022 VOUT+.t31 GNDA 0.325216f
C2023 VOUT+.t138 GNDA 0.319769f
C2024 VOUT+.n61 GNDA 0.214395f
C2025 VOUT+.t107 GNDA 0.319769f
C2026 VOUT+.n62 GNDA 0.134903f
C2027 VOUT+.t46 GNDA 0.324534f
C2028 VOUT+.t62 GNDA 0.325216f
C2029 VOUT+.t41 GNDA 0.319769f
C2030 VOUT+.n63 GNDA 0.214395f
C2031 VOUT+.t143 GNDA 0.319769f
C2032 VOUT+.n64 GNDA 0.134903f
C2033 VOUT+.t87 GNDA 0.324534f
C2034 VOUT+.t114 GNDA 0.325216f
C2035 VOUT+.t21 GNDA 0.319769f
C2036 VOUT+.n65 GNDA 0.214395f
C2037 VOUT+.t126 GNDA 0.319769f
C2038 VOUT+.n66 GNDA 0.134903f
C2039 VOUT+.t65 GNDA 0.324534f
C2040 VOUT+.t26 GNDA 0.324801f
C2041 VOUT+.t102 GNDA 0.324534f
C2042 VOUT+.t59 GNDA 0.324801f
C2043 VOUT+.t134 GNDA 0.324534f
C2044 VOUT+.t37 GNDA 0.324801f
C2045 VOUT+.t120 GNDA 0.324534f
C2046 VOUT+.t81 GNDA 0.324801f
C2047 VOUT+.t155 GNDA 0.324534f
C2048 VOUT+.t119 GNDA 0.319769f
C2049 VOUT+.n67 GNDA 0.353941f
C2050 VOUT+.t82 GNDA 0.319769f
C2051 VOUT+.n68 GNDA 0.413897f
C2052 VOUT+.t97 GNDA 0.319769f
C2053 VOUT+.n69 GNDA 0.413897f
C2054 VOUT+.t63 GNDA 0.319769f
C2055 VOUT+.n70 GNDA 0.413897f
C2056 VOUT+.t27 GNDA 0.319769f
C2057 VOUT+.n71 GNDA 0.339987f
C2058 VOUT+.t45 GNDA 0.319769f
C2059 VOUT+.n72 GNDA 0.339987f
C2060 VOUT+.t144 GNDA 0.319769f
C2061 VOUT+.n73 GNDA 0.339987f
C2062 VOUT+.t112 GNDA 0.319769f
C2063 VOUT+.n74 GNDA 0.339987f
C2064 VOUT+.t76 GNDA 0.319769f
C2065 VOUT+.n75 GNDA 0.275033f
C2066 VOUT+.t93 GNDA 0.319769f
C2067 VOUT+.n76 GNDA 0.275033f
C2068 VOUT+.t56 GNDA 0.319769f
C2069 VOUT+.t40 GNDA 0.325216f
C2070 VOUT+.t19 GNDA 0.319769f
C2071 VOUT+.n77 GNDA 0.214395f
C2072 VOUT+.n78 GNDA 0.259812f
C2073 VOUT+.t34 GNDA 0.325216f
C2074 VOUT+.t52 GNDA 0.319769f
C2075 VOUT+.n79 GNDA 0.214395f
C2076 VOUT+.t156 GNDA 0.319769f
C2077 VOUT+.t136 GNDA 0.325216f
C2078 VOUT+.t121 GNDA 0.319769f
C2079 VOUT+.n80 GNDA 0.214395f
C2080 VOUT+.n81 GNDA 0.259812f
C2081 VOUT+.t70 GNDA 0.325216f
C2082 VOUT+.t89 GNDA 0.319769f
C2083 VOUT+.n82 GNDA 0.214395f
C2084 VOUT+.t50 GNDA 0.319769f
C2085 VOUT+.t36 GNDA 0.325216f
C2086 VOUT+.t151 GNDA 0.319769f
C2087 VOUT+.n83 GNDA 0.214395f
C2088 VOUT+.n84 GNDA 0.259812f
C2089 VOUT+.t95 GNDA 0.325216f
C2090 VOUT+.t43 GNDA 0.319769f
C2091 VOUT+.n85 GNDA 0.214395f
C2092 VOUT+.t145 GNDA 0.319769f
C2093 VOUT+.t66 GNDA 0.325216f
C2094 VOUT+.t118 GNDA 0.319769f
C2095 VOUT+.n86 GNDA 0.214395f
C2096 VOUT+.n87 GNDA 0.259812f
C2097 VOUT+.t55 GNDA 0.325216f
C2098 VOUT+.t141 GNDA 0.319769f
C2099 VOUT+.n88 GNDA 0.214395f
C2100 VOUT+.t111 GNDA 0.319769f
C2101 VOUT+.t29 GNDA 0.325216f
C2102 VOUT+.t80 GNDA 0.319769f
C2103 VOUT+.n89 GNDA 0.214395f
C2104 VOUT+.n90 GNDA 0.259812f
C2105 VOUT+.t91 GNDA 0.325216f
C2106 VOUT+.t39 GNDA 0.319769f
C2107 VOUT+.n91 GNDA 0.214395f
C2108 VOUT+.t139 GNDA 0.319769f
C2109 VOUT+.t58 GNDA 0.325216f
C2110 VOUT+.t109 GNDA 0.319769f
C2111 VOUT+.n92 GNDA 0.214395f
C2112 VOUT+.n93 GNDA 0.259812f
C2113 VOUT+.t49 GNDA 0.325216f
C2114 VOUT+.t135 GNDA 0.319769f
C2115 VOUT+.n94 GNDA 0.214395f
C2116 VOUT+.t103 GNDA 0.319769f
C2117 VOUT+.t20 GNDA 0.325216f
C2118 VOUT+.t72 GNDA 0.319769f
C2119 VOUT+.n95 GNDA 0.214395f
C2120 VOUT+.n96 GNDA 0.259812f
C2121 VOUT+.t148 GNDA 0.325216f
C2122 VOUT+.t99 GNDA 0.319769f
C2123 VOUT+.n97 GNDA 0.214395f
C2124 VOUT+.t68 GNDA 0.319769f
C2125 VOUT+.t122 GNDA 0.325216f
C2126 VOUT+.t33 GNDA 0.319769f
C2127 VOUT+.n98 GNDA 0.214395f
C2128 VOUT+.n99 GNDA 0.259812f
C2129 VOUT+.t44 GNDA 0.325216f
C2130 VOUT+.t133 GNDA 0.319769f
C2131 VOUT+.n100 GNDA 0.214395f
C2132 VOUT+.t98 GNDA 0.319769f
C2133 VOUT+.t152 GNDA 0.325216f
C2134 VOUT+.t67 GNDA 0.319769f
C2135 VOUT+.n101 GNDA 0.214395f
C2136 VOUT+.n102 GNDA 0.259812f
C2137 VOUT+.t142 GNDA 0.325216f
C2138 VOUT+.t94 GNDA 0.319769f
C2139 VOUT+.n103 GNDA 0.214395f
C2140 VOUT+.t60 GNDA 0.319769f
C2141 VOUT+.t116 GNDA 0.325216f
C2142 VOUT+.t30 GNDA 0.319769f
C2143 VOUT+.n104 GNDA 0.214395f
C2144 VOUT+.n105 GNDA 0.259812f
C2145 VOUT+.t77 GNDA 0.325216f
C2146 VOUT+.t127 GNDA 0.319769f
C2147 VOUT+.n106 GNDA 0.214395f
C2148 VOUT+.t22 GNDA 0.319769f
C2149 VOUT+.n107 GNDA 0.259812f
C2150 VOUT+.t53 GNDA 0.319769f
C2151 VOUT+.n108 GNDA 0.139899f
C2152 VOUT+.t105 GNDA 0.319769f
C2153 VOUT+.n109 GNDA 0.254294f
C2154 VOUT+.n110 GNDA 0.313998f
C2155 two_stage_opamp_dummy_magic_21_0.VD2.n0 GNDA 0.483909f
C2156 two_stage_opamp_dummy_magic_21_0.VD2.n1 GNDA 0.099935f
C2157 two_stage_opamp_dummy_magic_21_0.VD2.n2 GNDA 0.167505f
C2158 two_stage_opamp_dummy_magic_21_0.VD2.t3 GNDA 0.053331f
C2159 two_stage_opamp_dummy_magic_21_0.VD2.t9 GNDA 0.053331f
C2160 two_stage_opamp_dummy_magic_21_0.VD2.n3 GNDA 0.116042f
C2161 two_stage_opamp_dummy_magic_21_0.VD2.n4 GNDA 0.192793f
C2162 two_stage_opamp_dummy_magic_21_0.VD2.t10 GNDA 0.053331f
C2163 two_stage_opamp_dummy_magic_21_0.VD2.t4 GNDA 0.053331f
C2164 two_stage_opamp_dummy_magic_21_0.VD2.n5 GNDA 0.116042f
C2165 two_stage_opamp_dummy_magic_21_0.VD2.n6 GNDA 0.461069f
C2166 two_stage_opamp_dummy_magic_21_0.VD2.t20 GNDA 0.053331f
C2167 two_stage_opamp_dummy_magic_21_0.VD2.t7 GNDA 0.053331f
C2168 two_stage_opamp_dummy_magic_21_0.VD2.n7 GNDA 0.116042f
C2169 two_stage_opamp_dummy_magic_21_0.VD2.n8 GNDA 0.461069f
C2170 two_stage_opamp_dummy_magic_21_0.VD2.t21 GNDA 0.053331f
C2171 two_stage_opamp_dummy_magic_21_0.VD2.t19 GNDA 0.053331f
C2172 two_stage_opamp_dummy_magic_21_0.VD2.n9 GNDA 0.116042f
C2173 two_stage_opamp_dummy_magic_21_0.VD2.n10 GNDA 0.442486f
C2174 two_stage_opamp_dummy_magic_21_0.VD2.n11 GNDA 0.203944f
C2175 two_stage_opamp_dummy_magic_21_0.VD2.n12 GNDA 0.119128f
C2176 two_stage_opamp_dummy_magic_21_0.VD2.n13 GNDA 0.203944f
C2177 two_stage_opamp_dummy_magic_21_0.VD2.t8 GNDA 0.053331f
C2178 two_stage_opamp_dummy_magic_21_0.VD2.t11 GNDA 0.053331f
C2179 two_stage_opamp_dummy_magic_21_0.VD2.n14 GNDA 0.116042f
C2180 two_stage_opamp_dummy_magic_21_0.VD2.n15 GNDA 0.442486f
C2181 two_stage_opamp_dummy_magic_21_0.VD2.n16 GNDA 0.192793f
C2182 two_stage_opamp_dummy_magic_21_0.VD2.n17 GNDA 0.106662f
C2183 two_stage_opamp_dummy_magic_21_0.VD2.n18 GNDA 0.205342f
C2184 two_stage_opamp_dummy_magic_21_0.VD2.t14 GNDA 0.053331f
C2185 two_stage_opamp_dummy_magic_21_0.VD2.t13 GNDA 0.053331f
C2186 two_stage_opamp_dummy_magic_21_0.VD2.n19 GNDA 0.116042f
C2187 two_stage_opamp_dummy_magic_21_0.VD2.n20 GNDA 0.465721f
C2188 two_stage_opamp_dummy_magic_21_0.VD2.n21 GNDA 0.205342f
C2189 two_stage_opamp_dummy_magic_21_0.VD2.t17 GNDA 0.053331f
C2190 two_stage_opamp_dummy_magic_21_0.VD2.t1 GNDA 0.053331f
C2191 two_stage_opamp_dummy_magic_21_0.VD2.n22 GNDA 0.116042f
C2192 two_stage_opamp_dummy_magic_21_0.VD2.n23 GNDA 0.447102f
C2193 two_stage_opamp_dummy_magic_21_0.VD2.n24 GNDA 0.192793f
C2194 two_stage_opamp_dummy_magic_21_0.VD2.t6 GNDA 0.053331f
C2195 two_stage_opamp_dummy_magic_21_0.VD2.t0 GNDA 0.053331f
C2196 two_stage_opamp_dummy_magic_21_0.VD2.n25 GNDA 0.116042f
C2197 two_stage_opamp_dummy_magic_21_0.VD2.n26 GNDA 0.447102f
C2198 two_stage_opamp_dummy_magic_21_0.VD2.n27 GNDA 0.113419f
C2199 two_stage_opamp_dummy_magic_21_0.VD2.t16 GNDA 0.053331f
C2200 two_stage_opamp_dummy_magic_21_0.VD2.t15 GNDA 0.053331f
C2201 two_stage_opamp_dummy_magic_21_0.VD2.n28 GNDA 0.116042f
C2202 two_stage_opamp_dummy_magic_21_0.VD2.n29 GNDA 0.465721f
C2203 two_stage_opamp_dummy_magic_21_0.VD2.t18 GNDA 0.053331f
C2204 two_stage_opamp_dummy_magic_21_0.VD2.t12 GNDA 0.053331f
C2205 two_stage_opamp_dummy_magic_21_0.VD2.n30 GNDA 0.116042f
C2206 two_stage_opamp_dummy_magic_21_0.VD2.n31 GNDA 0.447102f
C2207 two_stage_opamp_dummy_magic_21_0.VD2.n32 GNDA 0.192793f
C2208 two_stage_opamp_dummy_magic_21_0.VD2.n33 GNDA 0.113419f
C2209 two_stage_opamp_dummy_magic_21_0.VD2.t5 GNDA 0.053331f
C2210 two_stage_opamp_dummy_magic_21_0.VD2.t2 GNDA 0.053331f
C2211 two_stage_opamp_dummy_magic_21_0.VD2.n34 GNDA 0.116042f
C2212 two_stage_opamp_dummy_magic_21_0.VD2.n35 GNDA 0.447102f
C2213 VOUT-.t11 GNDA 0.047974f
C2214 VOUT-.t0 GNDA 0.047974f
C2215 VOUT-.n0 GNDA 0.098299f
C2216 VOUT-.n1 GNDA 0.251182f
C2217 VOUT-.n2 GNDA 0.034579f
C2218 VOUT-.n3 GNDA 0.061004f
C2219 VOUT-.t15 GNDA 0.047974f
C2220 VOUT-.t3 GNDA 0.047974f
C2221 VOUT-.n4 GNDA 0.098299f
C2222 VOUT-.n5 GNDA 0.292612f
C2223 VOUT-.t5 GNDA 0.047974f
C2224 VOUT-.t18 GNDA 0.047974f
C2225 VOUT-.n6 GNDA 0.098299f
C2226 VOUT-.n7 GNDA 0.287497f
C2227 VOUT-.n8 GNDA 0.061004f
C2228 VOUT-.n9 GNDA 0.034579f
C2229 VOUT-.t1 GNDA 0.047974f
C2230 VOUT-.t17 GNDA 0.047974f
C2231 VOUT-.n10 GNDA 0.098299f
C2232 VOUT-.n11 GNDA 0.287497f
C2233 VOUT-.n12 GNDA 0.034579f
C2234 VOUT-.t12 GNDA 0.047974f
C2235 VOUT-.t2 GNDA 0.047974f
C2236 VOUT-.n13 GNDA 0.098299f
C2237 VOUT-.n14 GNDA 0.287497f
C2238 VOUT-.n15 GNDA 0.034579f
C2239 VOUT-.n16 GNDA 0.061004f
C2240 VOUT-.t4 GNDA 0.047974f
C2241 VOUT-.t16 GNDA 0.047974f
C2242 VOUT-.n17 GNDA 0.098299f
C2243 VOUT-.n18 GNDA 0.292612f
C2244 VOUT-.n19 GNDA 0.050412f
C2245 VOUT-.n20 GNDA 0.199838f
C2246 VOUT-.t117 GNDA 0.325275f
C2247 VOUT-.t25 GNDA 0.319828f
C2248 VOUT-.n21 GNDA 0.214434f
C2249 VOUT-.t124 GNDA 0.319828f
C2250 VOUT-.n22 GNDA 0.139925f
C2251 VOUT-.t72 GNDA 0.325275f
C2252 VOUT-.t38 GNDA 0.319828f
C2253 VOUT-.n23 GNDA 0.214434f
C2254 VOUT-.t127 GNDA 0.319828f
C2255 VOUT-.t34 GNDA 0.324593f
C2256 VOUT-.t86 GNDA 0.324593f
C2257 VOUT-.t42 GNDA 0.324593f
C2258 VOUT-.t96 GNDA 0.324593f
C2259 VOUT-.t143 GNDA 0.324593f
C2260 VOUT-.t106 GNDA 0.324593f
C2261 VOUT-.t154 GNDA 0.324593f
C2262 VOUT-.t64 GNDA 0.324593f
C2263 VOUT-.t116 GNDA 0.324593f
C2264 VOUT-.t73 GNDA 0.324593f
C2265 VOUT-.t149 GNDA 0.319828f
C2266 VOUT-.n24 GNDA 0.215116f
C2267 VOUT-.t58 GNDA 0.319828f
C2268 VOUT-.n25 GNDA 0.275084f
C2269 VOUT-.t97 GNDA 0.319828f
C2270 VOUT-.n26 GNDA 0.275084f
C2271 VOUT-.t131 GNDA 0.319828f
C2272 VOUT-.n27 GNDA 0.275084f
C2273 VOUT-.t24 GNDA 0.319828f
C2274 VOUT-.n28 GNDA 0.275084f
C2275 VOUT-.t75 GNDA 0.319828f
C2276 VOUT-.n29 GNDA 0.275084f
C2277 VOUT-.t113 GNDA 0.319828f
C2278 VOUT-.n30 GNDA 0.275084f
C2279 VOUT-.t144 GNDA 0.319828f
C2280 VOUT-.n31 GNDA 0.275084f
C2281 VOUT-.t54 GNDA 0.319828f
C2282 VOUT-.n32 GNDA 0.275084f
C2283 VOUT-.t94 GNDA 0.319828f
C2284 VOUT-.n33 GNDA 0.275084f
C2285 VOUT-.n34 GNDA 0.25986f
C2286 VOUT-.t37 GNDA 0.325275f
C2287 VOUT-.t142 GNDA 0.319828f
C2288 VOUT-.n35 GNDA 0.214434f
C2289 VOUT-.t93 GNDA 0.319828f
C2290 VOUT-.t20 GNDA 0.325275f
C2291 VOUT-.t57 GNDA 0.319828f
C2292 VOUT-.n36 GNDA 0.214434f
C2293 VOUT-.n37 GNDA 0.25986f
C2294 VOUT-.t79 GNDA 0.325275f
C2295 VOUT-.t41 GNDA 0.319828f
C2296 VOUT-.n38 GNDA 0.214434f
C2297 VOUT-.t133 GNDA 0.319828f
C2298 VOUT-.t60 GNDA 0.325275f
C2299 VOUT-.t100 GNDA 0.319828f
C2300 VOUT-.n39 GNDA 0.214434f
C2301 VOUT-.n40 GNDA 0.25986f
C2302 VOUT-.t121 GNDA 0.325275f
C2303 VOUT-.t83 GNDA 0.319828f
C2304 VOUT-.n41 GNDA 0.214434f
C2305 VOUT-.t31 GNDA 0.319828f
C2306 VOUT-.t104 GNDA 0.325275f
C2307 VOUT-.t137 GNDA 0.319828f
C2308 VOUT-.n42 GNDA 0.214434f
C2309 VOUT-.n43 GNDA 0.25986f
C2310 VOUT-.t84 GNDA 0.325275f
C2311 VOUT-.t49 GNDA 0.319828f
C2312 VOUT-.n44 GNDA 0.214434f
C2313 VOUT-.t138 GNDA 0.319828f
C2314 VOUT-.t66 GNDA 0.325275f
C2315 VOUT-.t103 GNDA 0.319828f
C2316 VOUT-.n45 GNDA 0.214434f
C2317 VOUT-.n46 GNDA 0.25986f
C2318 VOUT-.t108 GNDA 0.325275f
C2319 VOUT-.t69 GNDA 0.319828f
C2320 VOUT-.n47 GNDA 0.214434f
C2321 VOUT-.t90 GNDA 0.319828f
C2322 VOUT-.n48 GNDA 0.139925f
C2323 VOUT-.t67 GNDA 0.325275f
C2324 VOUT-.t30 GNDA 0.319828f
C2325 VOUT-.n49 GNDA 0.214434f
C2326 VOUT-.t51 GNDA 0.319828f
C2327 VOUT-.t53 GNDA 0.324593f
C2328 VOUT-.t156 GNDA 0.324593f
C2329 VOUT-.t44 GNDA 0.325275f
C2330 VOUT-.t136 GNDA 0.319828f
C2331 VOUT-.n50 GNDA 0.214434f
C2332 VOUT-.t101 GNDA 0.319828f
C2333 VOUT-.n51 GNDA 0.134927f
C2334 VOUT-.t36 GNDA 0.324593f
C2335 VOUT-.t151 GNDA 0.325275f
C2336 VOUT-.t98 GNDA 0.319828f
C2337 VOUT-.n52 GNDA 0.214434f
C2338 VOUT-.t59 GNDA 0.319828f
C2339 VOUT-.n53 GNDA 0.134927f
C2340 VOUT-.t140 GNDA 0.324593f
C2341 VOUT-.t118 GNDA 0.325275f
C2342 VOUT-.t56 GNDA 0.319828f
C2343 VOUT-.n54 GNDA 0.214434f
C2344 VOUT-.t21 GNDA 0.319828f
C2345 VOUT-.n55 GNDA 0.134927f
C2346 VOUT-.t105 GNDA 0.324593f
C2347 VOUT-.t65 GNDA 0.325275f
C2348 VOUT-.t80 GNDA 0.319828f
C2349 VOUT-.n56 GNDA 0.214434f
C2350 VOUT-.t43 GNDA 0.319828f
C2351 VOUT-.n57 GNDA 0.134927f
C2352 VOUT-.t125 GNDA 0.324593f
C2353 VOUT-.t145 GNDA 0.324861f
C2354 VOUT-.t87 GNDA 0.324593f
C2355 VOUT-.t110 GNDA 0.324861f
C2356 VOUT-.t50 GNDA 0.324593f
C2357 VOUT-.t70 GNDA 0.324861f
C2358 VOUT-.t150 GNDA 0.324593f
C2359 VOUT-.t95 GNDA 0.324861f
C2360 VOUT-.t32 GNDA 0.324593f
C2361 VOUT-.t134 GNDA 0.319828f
C2362 VOUT-.n58 GNDA 0.354006f
C2363 VOUT-.t111 GNDA 0.319828f
C2364 VOUT-.n59 GNDA 0.413973f
C2365 VOUT-.t147 GNDA 0.319828f
C2366 VOUT-.n60 GNDA 0.413973f
C2367 VOUT-.t45 GNDA 0.319828f
C2368 VOUT-.n61 GNDA 0.413973f
C2369 VOUT-.t85 GNDA 0.319828f
C2370 VOUT-.n62 GNDA 0.340049f
C2371 VOUT-.t61 GNDA 0.319828f
C2372 VOUT-.n63 GNDA 0.340049f
C2373 VOUT-.t102 GNDA 0.319828f
C2374 VOUT-.n64 GNDA 0.340049f
C2375 VOUT-.t139 GNDA 0.319828f
C2376 VOUT-.n65 GNDA 0.340049f
C2377 VOUT-.t119 GNDA 0.319828f
C2378 VOUT-.n66 GNDA 0.275084f
C2379 VOUT-.t155 GNDA 0.319828f
C2380 VOUT-.n67 GNDA 0.275084f
C2381 VOUT-.n68 GNDA 0.25986f
C2382 VOUT-.t27 GNDA 0.325275f
C2383 VOUT-.t130 GNDA 0.319828f
C2384 VOUT-.n69 GNDA 0.214434f
C2385 VOUT-.t152 GNDA 0.319828f
C2386 VOUT-.t76 GNDA 0.325275f
C2387 VOUT-.t115 GNDA 0.319828f
C2388 VOUT-.n70 GNDA 0.214434f
C2389 VOUT-.n71 GNDA 0.25986f
C2390 VOUT-.t62 GNDA 0.325275f
C2391 VOUT-.t23 GNDA 0.319828f
C2392 VOUT-.n72 GNDA 0.214434f
C2393 VOUT-.t47 GNDA 0.319828f
C2394 VOUT-.t112 GNDA 0.325275f
C2395 VOUT-.t148 GNDA 0.319828f
C2396 VOUT-.n73 GNDA 0.214434f
C2397 VOUT-.n74 GNDA 0.25986f
C2398 VOUT-.t114 GNDA 0.325275f
C2399 VOUT-.t78 GNDA 0.319828f
C2400 VOUT-.n75 GNDA 0.214434f
C2401 VOUT-.t26 GNDA 0.319828f
C2402 VOUT-.t99 GNDA 0.325275f
C2403 VOUT-.t132 GNDA 0.319828f
C2404 VOUT-.n76 GNDA 0.214434f
C2405 VOUT-.n77 GNDA 0.25986f
C2406 VOUT-.t74 GNDA 0.325275f
C2407 VOUT-.t39 GNDA 0.319828f
C2408 VOUT-.n78 GNDA 0.214434f
C2409 VOUT-.t128 GNDA 0.319828f
C2410 VOUT-.t55 GNDA 0.325275f
C2411 VOUT-.t92 GNDA 0.319828f
C2412 VOUT-.n79 GNDA 0.214434f
C2413 VOUT-.n80 GNDA 0.25986f
C2414 VOUT-.t109 GNDA 0.325275f
C2415 VOUT-.t71 GNDA 0.319828f
C2416 VOUT-.n81 GNDA 0.214434f
C2417 VOUT-.t19 GNDA 0.319828f
C2418 VOUT-.t91 GNDA 0.325275f
C2419 VOUT-.t126 GNDA 0.319828f
C2420 VOUT-.n82 GNDA 0.214434f
C2421 VOUT-.n83 GNDA 0.25986f
C2422 VOUT-.t68 GNDA 0.325275f
C2423 VOUT-.t33 GNDA 0.319828f
C2424 VOUT-.n84 GNDA 0.214434f
C2425 VOUT-.t122 GNDA 0.319828f
C2426 VOUT-.t52 GNDA 0.325275f
C2427 VOUT-.t88 GNDA 0.319828f
C2428 VOUT-.n85 GNDA 0.214434f
C2429 VOUT-.n86 GNDA 0.25986f
C2430 VOUT-.t29 GNDA 0.325275f
C2431 VOUT-.t135 GNDA 0.319828f
C2432 VOUT-.n87 GNDA 0.214434f
C2433 VOUT-.t82 GNDA 0.319828f
C2434 VOUT-.t153 GNDA 0.325275f
C2435 VOUT-.t48 GNDA 0.319828f
C2436 VOUT-.n88 GNDA 0.214434f
C2437 VOUT-.n89 GNDA 0.25986f
C2438 VOUT-.t63 GNDA 0.325275f
C2439 VOUT-.t28 GNDA 0.319828f
C2440 VOUT-.n90 GNDA 0.214434f
C2441 VOUT-.t120 GNDA 0.319828f
C2442 VOUT-.t46 GNDA 0.325275f
C2443 VOUT-.t81 GNDA 0.319828f
C2444 VOUT-.n91 GNDA 0.214434f
C2445 VOUT-.n92 GNDA 0.25986f
C2446 VOUT-.t22 GNDA 0.325275f
C2447 VOUT-.t129 GNDA 0.319828f
C2448 VOUT-.n93 GNDA 0.214434f
C2449 VOUT-.t77 GNDA 0.319828f
C2450 VOUT-.t146 GNDA 0.325275f
C2451 VOUT-.t40 GNDA 0.319828f
C2452 VOUT-.n94 GNDA 0.214434f
C2453 VOUT-.n95 GNDA 0.25986f
C2454 VOUT-.t123 GNDA 0.325275f
C2455 VOUT-.t89 GNDA 0.319828f
C2456 VOUT-.n96 GNDA 0.214434f
C2457 VOUT-.t35 GNDA 0.319828f
C2458 VOUT-.n97 GNDA 0.25986f
C2459 VOUT-.t141 GNDA 0.319828f
C2460 VOUT-.n98 GNDA 0.139925f
C2461 VOUT-.t107 GNDA 0.319828f
C2462 VOUT-.n99 GNDA 0.254341f
C2463 VOUT-.n100 GNDA 0.313661f
C2464 VOUT-.n101 GNDA 0.084665f
C2465 VOUT-.t9 GNDA 0.05597f
C2466 VOUT-.t13 GNDA 0.05597f
C2467 VOUT-.n102 GNDA 0.120258f
C2468 VOUT-.n103 GNDA 0.336222f
C2469 VOUT-.t8 GNDA 0.05597f
C2470 VOUT-.t7 GNDA 0.05597f
C2471 VOUT-.n104 GNDA 0.120258f
C2472 VOUT-.n105 GNDA 0.323957f
C2473 VOUT-.n106 GNDA 0.117384f
C2474 VOUT-.t14 GNDA 0.05597f
C2475 VOUT-.t6 GNDA 0.05597f
C2476 VOUT-.n107 GNDA 0.120258f
C2477 VOUT-.n108 GNDA 0.328894f
C2478 VOUT-.n109 GNDA 0.056732f
C2479 VOUT-.t10 GNDA 0.092493f
C2480 VOUT-.n110 GNDA 0.109206f
C2481 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t1 GNDA 0.125517f
C2482 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t3 GNDA 0.340499f
C2483 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t6 GNDA 0.313782f
C2484 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t9 GNDA 0.313782f
C2485 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t5 GNDA 0.37241f
C2486 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n0 GNDA 0.196704f
C2487 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n1 GNDA 0.124569f
C2488 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n2 GNDA 0.118809f
C2489 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n3 GNDA 0.608541f
C2490 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t2 GNDA 0.365905f
C2491 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t4 GNDA 0.313782f
C2492 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t8 GNDA 0.37241f
C2493 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n4 GNDA 0.195093f
C2494 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t7 GNDA 0.317627f
C2495 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n5 GNDA 0.210094f
C2496 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.n6 GNDA 0.585951f
C2497 two_stage_opamp_dummy_magic_21_0.V_b_2nd_stage.t0 GNDA 0.124526f
C2498 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t7 GNDA 0.011263f
C2499 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t3 GNDA 0.011263f
C2500 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n0 GNDA 0.028194f
C2501 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t5 GNDA 0.011263f
C2502 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t4 GNDA 0.011263f
C2503 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n1 GNDA 0.028194f
C2504 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t1 GNDA 0.011263f
C2505 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t2 GNDA 0.011263f
C2506 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n2 GNDA 0.028042f
C2507 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n3 GNDA 0.190415f
C2508 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n4 GNDA 0.159941f
C2509 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t11 GNDA 0.011263f
C2510 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t6 GNDA 0.011263f
C2511 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n5 GNDA 0.022525f
C2512 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n6 GNDA 0.039991f
C2513 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t0 GNDA 0.016894f
C2514 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t10 GNDA 0.016894f
C2515 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n7 GNDA 0.039235f
C2516 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t31 GNDA 0.029987f
C2517 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t22 GNDA 0.029987f
C2518 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t28 GNDA 0.029987f
C2519 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t18 GNDA 0.029987f
C2520 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t26 GNDA 0.029987f
C2521 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t16 GNDA 0.029987f
C2522 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t24 GNDA 0.029987f
C2523 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t13 GNDA 0.029987f
C2524 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t20 GNDA 0.029987f
C2525 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t14 GNDA 0.034999f
C2526 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n8 GNDA 0.032999f
C2527 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n9 GNDA 0.020695f
C2528 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n10 GNDA 0.020695f
C2529 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n11 GNDA 0.020695f
C2530 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n12 GNDA 0.020695f
C2531 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n13 GNDA 0.020695f
C2532 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n14 GNDA 0.020695f
C2533 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n15 GNDA 0.020695f
C2534 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n16 GNDA 0.018493f
C2535 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t19 GNDA 0.029987f
C2536 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t29 GNDA 0.029987f
C2537 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t23 GNDA 0.029987f
C2538 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t15 GNDA 0.029987f
C2539 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t25 GNDA 0.029987f
C2540 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t17 GNDA 0.029987f
C2541 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t27 GNDA 0.029987f
C2542 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t21 GNDA 0.029987f
C2543 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t30 GNDA 0.029987f
C2544 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t12 GNDA 0.034999f
C2545 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n17 GNDA 0.032999f
C2546 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n18 GNDA 0.020695f
C2547 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n19 GNDA 0.020695f
C2548 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n20 GNDA 0.020695f
C2549 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n21 GNDA 0.020695f
C2550 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n22 GNDA 0.020695f
C2551 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n23 GNDA 0.020695f
C2552 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n24 GNDA 0.020695f
C2553 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n25 GNDA 0.018493f
C2554 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n26 GNDA 0.015655f
C2555 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n27 GNDA 0.236254f
C2556 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t9 GNDA 0.016894f
C2557 two_stage_opamp_dummy_magic_21_0.V_tail_gate.t8 GNDA 0.016894f
C2558 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n28 GNDA 0.036759f
C2559 two_stage_opamp_dummy_magic_21_0.V_tail_gate.n29 GNDA 0.166086f
C2560 two_stage_opamp_dummy_magic_21_0.err_amp_out.n0 GNDA 0.012844f
C2561 two_stage_opamp_dummy_magic_21_0.err_amp_out.n1 GNDA 0.012527f
C2562 two_stage_opamp_dummy_magic_21_0.err_amp_out.n2 GNDA 0.325317f
C2563 two_stage_opamp_dummy_magic_21_0.err_amp_out.n3 GNDA 0.012527f
C2564 two_stage_opamp_dummy_magic_21_0.err_amp_out.n4 GNDA 0.095072f
C2565 two_stage_opamp_dummy_magic_21_0.err_amp_out.t12 GNDA 0.054088f
C2566 two_stage_opamp_dummy_magic_21_0.err_amp_out.n5 GNDA 0.012001f
C2567 two_stage_opamp_dummy_magic_21_0.err_amp_out.n6 GNDA 0.124861f
C2568 two_stage_opamp_dummy_magic_21_0.err_amp_out.n7 GNDA 0.012001f
C2569 two_stage_opamp_dummy_magic_21_0.err_amp_out.n8 GNDA 0.10815f
C2570 two_stage_opamp_dummy_magic_21_0.err_amp_out.n9 GNDA 0.095072f
C2571 two_stage_opamp_dummy_magic_21_0.err_amp_out.n10 GNDA 0.719147f
C2572 two_stage_opamp_dummy_magic_21_0.err_amp_out.n11 GNDA 0.012001f
C2573 two_stage_opamp_dummy_magic_21_0.err_amp_out.n12 GNDA 0.10815f
C2574 two_stage_opamp_dummy_magic_21_0.err_amp_out.n13 GNDA 0.057175f
C2575 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n0 GNDA 0.408216f
C2576 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n1 GNDA 0.318908f
C2577 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n2 GNDA 0.362794f
C2578 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t9 GNDA 0.014742f
C2579 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t14 GNDA 0.014742f
C2580 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t5 GNDA 0.014742f
C2581 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n3 GNDA 0.031178f
C2582 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n4 GNDA 0.293793f
C2583 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t6 GNDA 0.012162f
C2584 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t17 GNDA 0.012162f
C2585 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t19 GNDA 0.012162f
C2586 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t12 GNDA 0.012162f
C2587 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t8 GNDA 0.012162f
C2588 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t21 GNDA 0.012162f
C2589 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t18 GNDA 0.012162f
C2590 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t4 GNDA 0.026351f
C2591 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n5 GNDA 0.041093f
C2592 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n6 GNDA 0.032064f
C2593 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n7 GNDA 0.028584f
C2594 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n8 GNDA 0.04506f
C2595 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n9 GNDA 0.028584f
C2596 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n10 GNDA 0.032064f
C2597 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n11 GNDA 0.032064f
C2598 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n12 GNDA 0.028584f
C2599 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t10 GNDA 0.012162f
C2600 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t20 GNDA 0.026351f
C2601 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n13 GNDA 0.037614f
C2602 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n14 GNDA 0.04506f
C2603 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t0 GNDA 0.014742f
C2604 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t3 GNDA 0.014742f
C2605 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n15 GNDA 0.030038f
C2606 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t2 GNDA 0.014742f
C2607 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t16 GNDA 0.014742f
C2608 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n16 GNDA 0.030038f
C2609 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n17 GNDA 0.249418f
C2610 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n18 GNDA 0.316023f
C2611 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t1 GNDA 0.014742f
C2612 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t15 GNDA 0.014742f
C2613 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n19 GNDA 0.030038f
C2614 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n20 GNDA 0.249418f
C2615 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n21 GNDA 0.320943f
C2616 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n22 GNDA 0.239385f
C2617 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n23 GNDA 0.23177f
C2618 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t7 GNDA 0.014742f
C2619 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t11 GNDA 0.014742f
C2620 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n24 GNDA 0.031178f
C2621 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n25 GNDA 0.348011f
C2622 two_stage_opamp_dummy_magic_21_0.err_amp_mir.n26 GNDA 0.031178f
C2623 two_stage_opamp_dummy_magic_21_0.err_amp_mir.t13 GNDA 0.014742f
C2624 bgr_0.V_TOP.t24 GNDA 0.095448f
C2625 bgr_0.V_TOP.t33 GNDA 0.095448f
C2626 bgr_0.V_TOP.t39 GNDA 0.095448f
C2627 bgr_0.V_TOP.t16 GNDA 0.095448f
C2628 bgr_0.V_TOP.t15 GNDA 0.095448f
C2629 bgr_0.V_TOP.t28 GNDA 0.095448f
C2630 bgr_0.V_TOP.t38 GNDA 0.095448f
C2631 bgr_0.V_TOP.t14 GNDA 0.095448f
C2632 bgr_0.V_TOP.t27 GNDA 0.095448f
C2633 bgr_0.V_TOP.t26 GNDA 0.095448f
C2634 bgr_0.V_TOP.t37 GNDA 0.095448f
C2635 bgr_0.V_TOP.t46 GNDA 0.095448f
C2636 bgr_0.V_TOP.t18 GNDA 0.095448f
C2637 bgr_0.V_TOP.t30 GNDA 0.095448f
C2638 bgr_0.V_TOP.t29 GNDA 0.124774f
C2639 bgr_0.V_TOP.n0 GNDA 0.069758f
C2640 bgr_0.V_TOP.n1 GNDA 0.050905f
C2641 bgr_0.V_TOP.n2 GNDA 0.050905f
C2642 bgr_0.V_TOP.n3 GNDA 0.050905f
C2643 bgr_0.V_TOP.n4 GNDA 0.050905f
C2644 bgr_0.V_TOP.n5 GNDA 0.04747f
C2645 bgr_0.V_TOP.t9 GNDA 0.122745f
C2646 bgr_0.V_TOP.t40 GNDA 0.36361f
C2647 bgr_0.V_TOP.t31 GNDA 0.369803f
C2648 bgr_0.V_TOP.t35 GNDA 0.36361f
C2649 bgr_0.V_TOP.n6 GNDA 0.243789f
C2650 bgr_0.V_TOP.t32 GNDA 0.36361f
C2651 bgr_0.V_TOP.t22 GNDA 0.369803f
C2652 bgr_0.V_TOP.n7 GNDA 0.311966f
C2653 bgr_0.V_TOP.t20 GNDA 0.369803f
C2654 bgr_0.V_TOP.t25 GNDA 0.36361f
C2655 bgr_0.V_TOP.n8 GNDA 0.243789f
C2656 bgr_0.V_TOP.t21 GNDA 0.36361f
C2657 bgr_0.V_TOP.t45 GNDA 0.369803f
C2658 bgr_0.V_TOP.n9 GNDA 0.380142f
C2659 bgr_0.V_TOP.t42 GNDA 0.369803f
C2660 bgr_0.V_TOP.t49 GNDA 0.36361f
C2661 bgr_0.V_TOP.n10 GNDA 0.243789f
C2662 bgr_0.V_TOP.t44 GNDA 0.36361f
C2663 bgr_0.V_TOP.t36 GNDA 0.369803f
C2664 bgr_0.V_TOP.n11 GNDA 0.380142f
C2665 bgr_0.V_TOP.t17 GNDA 0.369803f
C2666 bgr_0.V_TOP.t23 GNDA 0.36361f
C2667 bgr_0.V_TOP.n12 GNDA 0.243789f
C2668 bgr_0.V_TOP.t19 GNDA 0.36361f
C2669 bgr_0.V_TOP.t43 GNDA 0.369803f
C2670 bgr_0.V_TOP.n13 GNDA 0.380142f
C2671 bgr_0.V_TOP.t34 GNDA 0.369803f
C2672 bgr_0.V_TOP.t41 GNDA 0.36361f
C2673 bgr_0.V_TOP.n14 GNDA 0.311966f
C2674 bgr_0.V_TOP.t47 GNDA 0.36361f
C2675 bgr_0.V_TOP.n15 GNDA 0.159079f
C2676 bgr_0.V_TOP.n16 GNDA 0.544408f
C2677 bgr_0.V_TOP.t1 GNDA 0.102288f
C2678 bgr_0.V_TOP.n17 GNDA 0.724299f
C2679 bgr_0.V_TOP.n18 GNDA 0.022634f
C2680 bgr_0.V_TOP.n19 GNDA 0.414649f
C2681 bgr_0.V_TOP.n20 GNDA 0.021924f
C2682 bgr_0.V_TOP.n21 GNDA 0.022786f
C2683 bgr_0.V_TOP.n22 GNDA 0.022634f
C2684 bgr_0.V_TOP.n23 GNDA 0.209756f
C2685 bgr_0.V_TOP.n24 GNDA 0.127416f
C2686 bgr_0.V_TOP.n25 GNDA 0.072722f
C2687 bgr_0.V_TOP.n26 GNDA 0.022634f
C2688 bgr_0.V_TOP.n27 GNDA 0.125537f
C2689 bgr_0.V_TOP.n28 GNDA 0.022634f
C2690 bgr_0.V_TOP.n29 GNDA 0.124344f
C2691 bgr_0.V_TOP.n30 GNDA 0.273328f
C2692 bgr_0.V_TOP.n31 GNDA 0.019234f
C2693 bgr_0.V_TOP.n32 GNDA 0.04747f
C2694 bgr_0.V_TOP.n33 GNDA 0.050905f
C2695 bgr_0.V_TOP.n34 GNDA 0.050905f
C2696 bgr_0.V_TOP.n35 GNDA 0.050905f
C2697 bgr_0.V_TOP.n36 GNDA 0.050905f
C2698 bgr_0.V_TOP.n37 GNDA 0.050905f
C2699 bgr_0.V_TOP.n38 GNDA 0.050905f
C2700 bgr_0.V_TOP.n39 GNDA 0.04747f
C2701 bgr_0.V_TOP.t48 GNDA 0.109989f
C2702 VDDA.t282 GNDA 0.033583f
C2703 VDDA.t290 GNDA 0.033583f
C2704 VDDA.n0 GNDA 0.071315f
C2705 VDDA.t312 GNDA 0.033583f
C2706 VDDA.t274 GNDA 0.033583f
C2707 VDDA.n1 GNDA 0.085242f
C2708 VDDA.n2 GNDA 0.238109f
C2709 VDDA.t334 GNDA 0.058886f
C2710 VDDA.t387 GNDA 0.119458f
C2711 VDDA.t310 GNDA 0.033583f
C2712 VDDA.t306 GNDA 0.033583f
C2713 VDDA.n3 GNDA 0.085242f
C2714 VDDA.n4 GNDA 0.265957f
C2715 VDDA.t385 GNDA 0.058886f
C2716 VDDA.n5 GNDA 0.17497f
C2717 VDDA.n6 GNDA 0.346536f
C2718 VDDA.t386 GNDA 0.286254f
C2719 VDDA.t309 GNDA 0.224523f
C2720 VDDA.t305 GNDA 0.224523f
C2721 VDDA.t311 GNDA 0.224523f
C2722 VDDA.t273 GNDA 0.224523f
C2723 VDDA.t281 GNDA 0.224523f
C2724 VDDA.t289 GNDA 0.224523f
C2725 VDDA.t283 GNDA 0.224523f
C2726 VDDA.t307 GNDA 0.224523f
C2727 VDDA.t313 GNDA 0.224523f
C2728 VDDA.t275 GNDA 0.224523f
C2729 VDDA.t335 GNDA 0.289995f
C2730 VDDA.t336 GNDA 0.119458f
C2731 VDDA.n7 GNDA 0.361505f
C2732 VDDA.n8 GNDA 0.17497f
C2733 VDDA.t314 GNDA 0.033583f
C2734 VDDA.t276 GNDA 0.033583f
C2735 VDDA.n9 GNDA 0.085242f
C2736 VDDA.n10 GNDA 0.265957f
C2737 VDDA.t284 GNDA 0.033583f
C2738 VDDA.t308 GNDA 0.033583f
C2739 VDDA.n11 GNDA 0.085242f
C2740 VDDA.n12 GNDA 0.238109f
C2741 VDDA.n13 GNDA 0.030704f
C2742 VDDA.n14 GNDA 0.264461f
C2743 VDDA.t317 GNDA 0.028785f
C2744 VDDA.t467 GNDA 0.028785f
C2745 VDDA.n15 GNDA 0.09864f
C2746 VDDA.t235 GNDA 0.028785f
C2747 VDDA.t199 GNDA 0.028785f
C2748 VDDA.n16 GNDA 0.095271f
C2749 VDDA.n17 GNDA 0.365478f
C2750 VDDA.t20 GNDA 0.028785f
C2751 VDDA.t455 GNDA 0.028785f
C2752 VDDA.n18 GNDA 0.095271f
C2753 VDDA.n19 GNDA 0.187782f
C2754 VDDA.t443 GNDA 0.028785f
C2755 VDDA.t157 GNDA 0.028785f
C2756 VDDA.n20 GNDA 0.095271f
C2757 VDDA.n21 GNDA 0.187782f
C2758 VDDA.t468 GNDA 0.028785f
C2759 VDDA.t150 GNDA 0.028785f
C2760 VDDA.n22 GNDA 0.095271f
C2761 VDDA.n23 GNDA 0.187782f
C2762 VDDA.t191 GNDA 0.028785f
C2763 VDDA.t318 GNDA 0.028785f
C2764 VDDA.n24 GNDA 0.095271f
C2765 VDDA.n25 GNDA 0.275108f
C2766 VDDA.t382 GNDA 0.028028f
C2767 VDDA.n26 GNDA 0.146554f
C2768 VDDA.t384 GNDA 0.068464f
C2769 VDDA.n27 GNDA 0.210326f
C2770 VDDA.t383 GNDA 0.170563f
C2771 VDDA.t454 GNDA 0.126654f
C2772 VDDA.t192 GNDA 0.126654f
C2773 VDDA.t457 GNDA 0.126654f
C2774 VDDA.t178 GNDA 0.126654f
C2775 VDDA.t181 GNDA 0.126654f
C2776 VDDA.t198 GNDA 0.126654f
C2777 VDDA.t466 GNDA 0.126654f
C2778 VDDA.t0 GNDA 0.126654f
C2779 VDDA.t456 GNDA 0.126654f
C2780 VDDA.t197 GNDA 0.126654f
C2781 VDDA.t395 GNDA 0.170563f
C2782 VDDA.t396 GNDA 0.068464f
C2783 VDDA.n28 GNDA 0.210326f
C2784 VDDA.t394 GNDA 0.028028f
C2785 VDDA.n29 GNDA 0.111929f
C2786 VDDA.n30 GNDA 0.149323f
C2787 VDDA.n31 GNDA 0.178378f
C2788 VDDA.t379 GNDA 0.013638f
C2789 VDDA.n32 GNDA 0.120653f
C2790 VDDA.t381 GNDA 0.017482f
C2791 VDDA.n33 GNDA 0.054499f
C2792 VDDA.t380 GNDA 0.071842f
C2793 VDDA.t48 GNDA 0.047495f
C2794 VDDA.t438 GNDA 0.047495f
C2795 VDDA.t112 GNDA 0.047495f
C2796 VDDA.t204 GNDA 0.047495f
C2797 VDDA.t1 GNDA 0.047495f
C2798 VDDA.t439 GNDA 0.047495f
C2799 VDDA.t207 GNDA 0.047495f
C2800 VDDA.t442 GNDA 0.047495f
C2801 VDDA.t186 GNDA 0.047495f
C2802 VDDA.t208 GNDA 0.047495f
C2803 VDDA.t362 GNDA 0.071842f
C2804 VDDA.t363 GNDA 0.017482f
C2805 VDDA.n34 GNDA 0.054499f
C2806 VDDA.t361 GNDA 0.013638f
C2807 VDDA.n35 GNDA 0.086142f
C2808 VDDA.n36 GNDA 0.171686f
C2809 VDDA.n37 GNDA 0.102504f
C2810 VDDA.t22 GNDA 0.05757f
C2811 VDDA.t183 GNDA 0.05757f
C2812 VDDA.n38 GNDA 0.171518f
C2813 VDDA.n39 GNDA 0.351889f
C2814 VDDA.t351 GNDA 0.202604f
C2815 VDDA.t81 GNDA 0.05757f
C2816 VDDA.t212 GNDA 0.05757f
C2817 VDDA.n40 GNDA 0.171518f
C2818 VDDA.n41 GNDA 0.351889f
C2819 VDDA.t445 GNDA 0.05757f
C2820 VDDA.t226 GNDA 0.05757f
C2821 VDDA.n42 GNDA 0.171518f
C2822 VDDA.n43 GNDA 0.351889f
C2823 VDDA.t463 GNDA 0.05757f
C2824 VDDA.t73 GNDA 0.05757f
C2825 VDDA.n44 GNDA 0.171518f
C2826 VDDA.n45 GNDA 0.351889f
C2827 VDDA.t180 GNDA 0.05757f
C2828 VDDA.t196 GNDA 0.05757f
C2829 VDDA.n46 GNDA 0.171518f
C2830 VDDA.n47 GNDA 0.372527f
C2831 VDDA.t349 GNDA 0.069848f
C2832 VDDA.n48 GNDA 0.159504f
C2833 VDDA.n49 GNDA 0.677725f
C2834 VDDA.t350 GNDA 0.438944f
C2835 VDDA.t179 GNDA 0.337744f
C2836 VDDA.t195 GNDA 0.337744f
C2837 VDDA.t462 GNDA 0.337744f
C2838 VDDA.t72 GNDA 0.337744f
C2839 VDDA.t444 GNDA 0.337744f
C2840 VDDA.t225 GNDA 0.337744f
C2841 VDDA.t80 GNDA 0.337744f
C2842 VDDA.t211 GNDA 0.337744f
C2843 VDDA.t21 GNDA 0.337744f
C2844 VDDA.t182 GNDA 0.337744f
C2845 VDDA.t365 GNDA 0.438944f
C2846 VDDA.t366 GNDA 0.202604f
C2847 VDDA.n50 GNDA 0.677725f
C2848 VDDA.t364 GNDA 0.069848f
C2849 VDDA.n51 GNDA 0.15706f
C2850 VDDA.n52 GNDA 0.033156f
C2851 VDDA.n53 GNDA 0.0103f
C2852 VDDA.n54 GNDA 0.093806f
C2853 VDDA.t419 GNDA 0.013662f
C2854 VDDA.t415 GNDA 0.017482f
C2855 VDDA.n55 GNDA 0.0103f
C2856 VDDA.n56 GNDA 0.093806f
C2857 VDDA.n57 GNDA 0.0103f
C2858 VDDA.n58 GNDA 0.093806f
C2859 VDDA.n59 GNDA 0.0103f
C2860 VDDA.n60 GNDA 0.093806f
C2861 VDDA.n61 GNDA 0.0103f
C2862 VDDA.n62 GNDA 0.093806f
C2863 VDDA.n63 GNDA 0.0103f
C2864 VDDA.n64 GNDA 0.093806f
C2865 VDDA.n65 GNDA 0.0103f
C2866 VDDA.n66 GNDA 0.093806f
C2867 VDDA.n67 GNDA 0.0103f
C2868 VDDA.n68 GNDA 0.093806f
C2869 VDDA.n69 GNDA 0.0103f
C2870 VDDA.n70 GNDA 0.093806f
C2871 VDDA.n71 GNDA 0.0103f
C2872 VDDA.n72 GNDA 0.116516f
C2873 VDDA.t413 GNDA 0.013662f
C2874 VDDA.n73 GNDA 0.090282f
C2875 VDDA.n74 GNDA 0.054122f
C2876 VDDA.t414 GNDA 0.071842f
C2877 VDDA.t236 GNDA 0.047495f
C2878 VDDA.t247 GNDA 0.047495f
C2879 VDDA.t3 GNDA 0.047495f
C2880 VDDA.t29 GNDA 0.047495f
C2881 VDDA.t193 GNDA 0.047495f
C2882 VDDA.t139 GNDA 0.047495f
C2883 VDDA.t448 GNDA 0.047495f
C2884 VDDA.t27 GNDA 0.047495f
C2885 VDDA.t205 GNDA 0.047495f
C2886 VDDA.t172 GNDA 0.047495f
C2887 VDDA.t446 GNDA 0.047495f
C2888 VDDA.t105 GNDA 0.047495f
C2889 VDDA.t245 GNDA 0.047495f
C2890 VDDA.t123 GNDA 0.047495f
C2891 VDDA.t243 GNDA 0.047495f
C2892 VDDA.t13 GNDA 0.047495f
C2893 VDDA.t15 GNDA 0.047495f
C2894 VDDA.t450 GNDA 0.047495f
C2895 VDDA.t108 GNDA 0.047495f
C2896 VDDA.t11 GNDA 0.047495f
C2897 VDDA.t420 GNDA 0.071842f
C2898 VDDA.t421 GNDA 0.017482f
C2899 VDDA.n75 GNDA 0.054122f
C2900 VDDA.n76 GNDA 0.087748f
C2901 VDDA.n77 GNDA 0.071299f
C2902 VDDA.n78 GNDA 0.071483f
C2903 VDDA.n79 GNDA 0.190006f
C2904 VDDA.n80 GNDA 0.245655f
C2905 VDDA.t278 GNDA 0.033583f
C2906 VDDA.t286 GNDA 0.033583f
C2907 VDDA.n81 GNDA 0.071315f
C2908 VDDA.t296 GNDA 0.033583f
C2909 VDDA.t302 GNDA 0.033583f
C2910 VDDA.n82 GNDA 0.085242f
C2911 VDDA.n83 GNDA 0.238109f
C2912 VDDA.t410 GNDA 0.058886f
C2913 VDDA.t342 GNDA 0.119458f
C2914 VDDA.t292 GNDA 0.033583f
C2915 VDDA.t300 GNDA 0.033583f
C2916 VDDA.n84 GNDA 0.085242f
C2917 VDDA.n85 GNDA 0.265957f
C2918 VDDA.t340 GNDA 0.058886f
C2919 VDDA.n86 GNDA 0.17497f
C2920 VDDA.n87 GNDA 0.346536f
C2921 VDDA.t341 GNDA 0.286254f
C2922 VDDA.t291 GNDA 0.224523f
C2923 VDDA.t299 GNDA 0.224523f
C2924 VDDA.t295 GNDA 0.224523f
C2925 VDDA.t301 GNDA 0.224523f
C2926 VDDA.t277 GNDA 0.224523f
C2927 VDDA.t285 GNDA 0.224523f
C2928 VDDA.t293 GNDA 0.224523f
C2929 VDDA.t287 GNDA 0.224523f
C2930 VDDA.t297 GNDA 0.224523f
C2931 VDDA.t303 GNDA 0.224523f
C2932 VDDA.t411 GNDA 0.286254f
C2933 VDDA.t412 GNDA 0.119458f
C2934 VDDA.n88 GNDA 0.346536f
C2935 VDDA.n89 GNDA 0.17497f
C2936 VDDA.t298 GNDA 0.033583f
C2937 VDDA.t304 GNDA 0.033583f
C2938 VDDA.n90 GNDA 0.085242f
C2939 VDDA.n91 GNDA 0.265957f
C2940 VDDA.t294 GNDA 0.033583f
C2941 VDDA.t288 GNDA 0.033583f
C2942 VDDA.n92 GNDA 0.085242f
C2943 VDDA.n93 GNDA 0.238109f
C2944 VDDA.n94 GNDA 0.030704f
C2945 VDDA.n95 GNDA 0.264461f
C2946 VDDA.t138 GNDA 0.028785f
C2947 VDDA.t316 GNDA 0.028785f
C2948 VDDA.n96 GNDA 0.09864f
C2949 VDDA.t2 GNDA 0.028785f
C2950 VDDA.t136 GNDA 0.028785f
C2951 VDDA.n97 GNDA 0.095271f
C2952 VDDA.n98 GNDA 0.365478f
C2953 VDDA.t43 GNDA 0.028785f
C2954 VDDA.t89 GNDA 0.028785f
C2955 VDDA.n99 GNDA 0.095271f
C2956 VDDA.n100 GNDA 0.187782f
C2957 VDDA.t36 GNDA 0.028785f
C2958 VDDA.t217 GNDA 0.028785f
C2959 VDDA.n101 GNDA 0.095271f
C2960 VDDA.n102 GNDA 0.187782f
C2961 VDDA.t145 GNDA 0.028785f
C2962 VDDA.t45 GNDA 0.028785f
C2963 VDDA.n103 GNDA 0.095271f
C2964 VDDA.n104 GNDA 0.187782f
C2965 VDDA.t315 GNDA 0.028785f
C2966 VDDA.t86 GNDA 0.028785f
C2967 VDDA.n105 GNDA 0.095271f
C2968 VDDA.n106 GNDA 0.275108f
C2969 VDDA.t343 GNDA 0.028028f
C2970 VDDA.n107 GNDA 0.146554f
C2971 VDDA.t345 GNDA 0.068464f
C2972 VDDA.n108 GNDA 0.210326f
C2973 VDDA.t344 GNDA 0.170563f
C2974 VDDA.t8 GNDA 0.126654f
C2975 VDDA.t218 GNDA 0.126654f
C2976 VDDA.t133 GNDA 0.126654f
C2977 VDDA.t137 GNDA 0.126654f
C2978 VDDA.t132 GNDA 0.126654f
C2979 VDDA.t219 GNDA 0.126654f
C2980 VDDA.t91 GNDA 0.126654f
C2981 VDDA.t90 GNDA 0.126654f
C2982 VDDA.t44 GNDA 0.126654f
C2983 VDDA.t31 GNDA 0.126654f
C2984 VDDA.t329 GNDA 0.170563f
C2985 VDDA.t330 GNDA 0.068464f
C2986 VDDA.n109 GNDA 0.210326f
C2987 VDDA.t328 GNDA 0.028028f
C2988 VDDA.n110 GNDA 0.111929f
C2989 VDDA.n111 GNDA 0.149323f
C2990 VDDA.n112 GNDA 0.178378f
C2991 VDDA.t358 GNDA 0.013638f
C2992 VDDA.n113 GNDA 0.120653f
C2993 VDDA.t360 GNDA 0.017482f
C2994 VDDA.n114 GNDA 0.054499f
C2995 VDDA.t359 GNDA 0.071842f
C2996 VDDA.t107 GNDA 0.047495f
C2997 VDDA.t440 GNDA 0.047495f
C2998 VDDA.t209 GNDA 0.047495f
C2999 VDDA.t17 GNDA 0.047495f
C3000 VDDA.t92 GNDA 0.047495f
C3001 VDDA.t441 GNDA 0.047495f
C3002 VDDA.t210 GNDA 0.047495f
C3003 VDDA.t100 GNDA 0.047495f
C3004 VDDA.t99 GNDA 0.047495f
C3005 VDDA.t127 GNDA 0.047495f
C3006 VDDA.t374 GNDA 0.071842f
C3007 VDDA.t375 GNDA 0.017482f
C3008 VDDA.n115 GNDA 0.054499f
C3009 VDDA.t373 GNDA 0.013638f
C3010 VDDA.n116 GNDA 0.086142f
C3011 VDDA.n117 GNDA 0.170995f
C3012 VDDA.n118 GNDA 0.102236f
C3013 VDDA.t83 GNDA 0.05757f
C3014 VDDA.t10 GNDA 0.05757f
C3015 VDDA.n119 GNDA 0.171518f
C3016 VDDA.n120 GNDA 0.351889f
C3017 VDDA.t321 GNDA 0.202604f
C3018 VDDA.t85 GNDA 0.05757f
C3019 VDDA.t221 GNDA 0.05757f
C3020 VDDA.n121 GNDA 0.171518f
C3021 VDDA.n122 GNDA 0.351889f
C3022 VDDA.t135 GNDA 0.05757f
C3023 VDDA.t144 GNDA 0.05757f
C3024 VDDA.n123 GNDA 0.171518f
C3025 VDDA.n124 GNDA 0.351889f
C3026 VDDA.t88 GNDA 0.05757f
C3027 VDDA.t35 GNDA 0.05757f
C3028 VDDA.n125 GNDA 0.171518f
C3029 VDDA.n126 GNDA 0.351889f
C3030 VDDA.t47 GNDA 0.05757f
C3031 VDDA.t33 GNDA 0.05757f
C3032 VDDA.n127 GNDA 0.171518f
C3033 VDDA.n128 GNDA 0.372527f
C3034 VDDA.t319 GNDA 0.069848f
C3035 VDDA.n129 GNDA 0.159504f
C3036 VDDA.n130 GNDA 0.677725f
C3037 VDDA.t320 GNDA 0.438944f
C3038 VDDA.t32 GNDA 0.337744f
C3039 VDDA.t46 GNDA 0.337744f
C3040 VDDA.t34 GNDA 0.337744f
C3041 VDDA.t87 GNDA 0.337744f
C3042 VDDA.t143 GNDA 0.337744f
C3043 VDDA.t134 GNDA 0.337744f
C3044 VDDA.t220 GNDA 0.337744f
C3045 VDDA.t84 GNDA 0.337744f
C3046 VDDA.t9 GNDA 0.337744f
C3047 VDDA.t82 GNDA 0.337744f
C3048 VDDA.t417 GNDA 0.438944f
C3049 VDDA.t418 GNDA 0.202604f
C3050 VDDA.n131 GNDA 0.677725f
C3051 VDDA.t416 GNDA 0.069848f
C3052 VDDA.n132 GNDA 0.15706f
C3053 VDDA.n133 GNDA 0.054822f
C3054 VDDA.n134 GNDA 0.193768f
C3055 VDDA.n135 GNDA 0.245176f
C3056 VDDA.n136 GNDA 0.239695f
C3057 VDDA.t175 GNDA 0.017271f
C3058 VDDA.t408 GNDA 0.017271f
C3059 VDDA.n137 GNDA 0.039065f
C3060 VDDA.n138 GNDA 0.155764f
C3061 VDDA.t400 GNDA 0.036095f
C3062 VDDA.t409 GNDA 0.062339f
C3063 VDDA.t406 GNDA 0.036095f
C3064 VDDA.n139 GNDA 0.095558f
C3065 VDDA.n140 GNDA 0.187693f
C3066 VDDA.t407 GNDA 0.167099f
C3067 VDDA.t174 GNDA 0.126654f
C3068 VDDA.t401 GNDA 0.167099f
C3069 VDDA.t402 GNDA 0.062339f
C3070 VDDA.n141 GNDA 0.187693f
C3071 VDDA.n142 GNDA 0.094649f
C3072 VDDA.n143 GNDA 0.054768f
C3073 VDDA.n144 GNDA 0.097493f
C3074 VDDA.n145 GNDA 0.240959f
C3075 VDDA.t346 GNDA 0.05947f
C3076 VDDA.t280 GNDA 0.033583f
C3077 VDDA.n146 GNDA 0.084362f
C3078 VDDA.t430 GNDA 0.15304f
C3079 VDDA.t428 GNDA 0.05947f
C3080 VDDA.n147 GNDA 0.125613f
C3081 VDDA.n148 GNDA 0.382089f
C3082 VDDA.t429 GNDA 0.286254f
C3083 VDDA.t279 GNDA 0.224523f
C3084 VDDA.t347 GNDA 0.286254f
C3085 VDDA.t348 GNDA 0.119458f
C3086 VDDA.n149 GNDA 0.382089f
C3087 VDDA.n150 GNDA 0.124704f
C3088 VDDA.n151 GNDA 0.054768f
C3089 VDDA.n152 GNDA 0.257238f
C3090 VDDA.n153 GNDA 5.30183f
C3091 VDDA.t148 GNDA 0.53636f
C3092 VDDA.t190 GNDA 0.538304f
C3093 VDDA.t229 GNDA 0.509519f
C3094 VDDA.t58 GNDA 0.53636f
C3095 VDDA.t115 GNDA 0.538304f
C3096 VDDA.t70 GNDA 0.509519f
C3097 VDDA.t69 GNDA 0.53636f
C3098 VDDA.t224 GNDA 0.538304f
C3099 VDDA.t49 GNDA 0.509519f
C3100 VDDA.t437 GNDA 0.53636f
C3101 VDDA.t118 GNDA 0.538304f
C3102 VDDA.t187 GNDA 0.509519f
C3103 VDDA.t233 GNDA 0.53636f
C3104 VDDA.t230 GNDA 0.538304f
C3105 VDDA.t114 GNDA 0.509519f
C3106 VDDA.n154 GNDA 0.359523f
C3107 VDDA.t234 GNDA 0.286307f
C3108 VDDA.n155 GNDA 0.390091f
C3109 VDDA.t113 GNDA 0.286307f
C3110 VDDA.n156 GNDA 0.390091f
C3111 VDDA.t71 GNDA 0.286307f
C3112 VDDA.n157 GNDA 0.390091f
C3113 VDDA.t436 GNDA 0.286307f
C3114 VDDA.n158 GNDA 0.390091f
C3115 VDDA.t149 GNDA 0.501562f
C3116 VDDA.n159 GNDA 4.46716f
C3117 VDDA.t469 GNDA 1.06077f
C3118 VDDA.t471 GNDA 1.13057f
C3119 VDDA.t472 GNDA 1.13013f
C3120 VDDA.t470 GNDA 1.08759f
C3121 VDDA.n160 GNDA 0.757073f
C3122 VDDA.n161 GNDA 0.371783f
C3123 VDDA.n162 GNDA 0.540415f
C3124 VDDA.n163 GNDA 0.986463f
C3125 VDDA.n164 GNDA 0.024133f
C3126 VDDA.n165 GNDA 0.097723f
C3127 VDDA.n166 GNDA 0.040579f
C3128 VDDA.t378 GNDA 0.033375f
C3129 VDDA.n168 GNDA 0.040579f
C3130 VDDA.n169 GNDA 0.024133f
C3131 VDDA.n170 GNDA 0.097723f
C3132 VDDA.t357 GNDA 0.033608f
C3133 VDDA.n171 GNDA 0.040579f
C3134 VDDA.n172 GNDA 0.024133f
C3135 VDDA.n173 GNDA 0.097723f
C3136 VDDA.n174 GNDA 0.024133f
C3137 VDDA.n175 GNDA 0.097723f
C3138 VDDA.n176 GNDA 0.024133f
C3139 VDDA.n177 GNDA 0.097723f
C3140 VDDA.n178 GNDA 0.024133f
C3141 VDDA.n179 GNDA 0.097723f
C3142 VDDA.n180 GNDA 0.024133f
C3143 VDDA.n181 GNDA 0.097723f
C3144 VDDA.n182 GNDA 0.024133f
C3145 VDDA.n183 GNDA 0.097723f
C3146 VDDA.n184 GNDA 0.024133f
C3147 VDDA.n185 GNDA 0.097723f
C3148 VDDA.n186 GNDA 0.024133f
C3149 VDDA.n187 GNDA 0.140434f
C3150 VDDA.n188 GNDA 0.037206f
C3151 VDDA.t331 GNDA 0.03542f
C3152 VDDA.t333 GNDA 0.033375f
C3153 VDDA.n189 GNDA 0.063974f
C3154 VDDA.n190 GNDA 0.097246f
C3155 VDDA.t332 GNDA 0.120603f
C3156 VDDA.t251 GNDA 0.080598f
C3157 VDDA.t59 GNDA 0.080598f
C3158 VDDA.t452 GNDA 0.080598f
C3159 VDDA.t261 GNDA 0.080598f
C3160 VDDA.t460 GNDA 0.080598f
C3161 VDDA.t265 GNDA 0.080598f
C3162 VDDA.t255 GNDA 0.080598f
C3163 VDDA.t95 GNDA 0.080598f
C3164 VDDA.t176 GNDA 0.080598f
C3165 VDDA.t18 GNDA 0.080598f
C3166 VDDA.t259 GNDA 0.080598f
C3167 VDDA.t249 GNDA 0.080598f
C3168 VDDA.t253 GNDA 0.080598f
C3169 VDDA.t155 GNDA 0.080598f
C3170 VDDA.t101 GNDA 0.080598f
C3171 VDDA.t41 GNDA 0.080598f
C3172 VDDA.t263 GNDA 0.080598f
C3173 VDDA.t257 GNDA 0.080598f
C3174 VDDA.t356 GNDA 0.122941f
C3175 VDDA.n191 GNDA 0.175052f
C3176 VDDA.t355 GNDA 0.023751f
C3177 VDDA.n192 GNDA 0.039251f
C3178 VDDA.n193 GNDA 0.071474f
C3179 VDDA.n194 GNDA 0.024133f
C3180 VDDA.n195 GNDA 0.097723f
C3181 VDDA.n196 GNDA 0.024133f
C3182 VDDA.n197 GNDA 0.097723f
C3183 VDDA.n198 GNDA 0.024133f
C3184 VDDA.n199 GNDA 0.097723f
C3185 VDDA.n200 GNDA 0.024133f
C3186 VDDA.n201 GNDA 0.097723f
C3187 VDDA.n202 GNDA 0.024133f
C3188 VDDA.n203 GNDA 0.097723f
C3189 VDDA.n204 GNDA 0.024133f
C3190 VDDA.n205 GNDA 0.097723f
C3191 VDDA.n206 GNDA 0.024133f
C3192 VDDA.n207 GNDA 0.097723f
C3193 VDDA.n208 GNDA 0.024133f
C3194 VDDA.n209 GNDA 0.097723f
C3195 VDDA.n210 GNDA 0.071474f
C3196 VDDA.n211 GNDA 0.035309f
C3197 VDDA.t391 GNDA 0.03542f
C3198 VDDA.t393 GNDA 0.033375f
C3199 VDDA.n212 GNDA 0.063974f
C3200 VDDA.n213 GNDA 0.097246f
C3201 VDDA.t392 GNDA 0.120603f
C3202 VDDA.t65 GNDA 0.080598f
C3203 VDDA.t6 GNDA 0.080598f
C3204 VDDA.t141 GNDA 0.080598f
C3205 VDDA.t162 GNDA 0.080598f
C3206 VDDA.t160 GNDA 0.080598f
C3207 VDDA.t166 GNDA 0.080598f
C3208 VDDA.t93 GNDA 0.080598f
C3209 VDDA.t110 GNDA 0.080598f
C3210 VDDA.t269 GNDA 0.080598f
C3211 VDDA.t241 GNDA 0.080598f
C3212 VDDA.t271 GNDA 0.080598f
C3213 VDDA.t153 GNDA 0.080598f
C3214 VDDA.t168 GNDA 0.080598f
C3215 VDDA.t170 GNDA 0.080598f
C3216 VDDA.t239 GNDA 0.080598f
C3217 VDDA.t202 GNDA 0.080598f
C3218 VDDA.t267 GNDA 0.080598f
C3219 VDDA.t67 GNDA 0.080598f
C3220 VDDA.t377 GNDA 0.099575f
C3221 VDDA.n214 GNDA 0.118274f
C3222 VDDA.n215 GNDA 0.064232f
C3223 VDDA.t376 GNDA 0.035402f
C3224 VDDA.n216 GNDA 0.035309f
C3225 VDDA.n217 GNDA 0.165644f
C3226 VDDA.n218 GNDA 0.319374f
C3227 VDDA.t117 GNDA 0.028785f
C3228 VDDA.t223 GNDA 0.028785f
C3229 VDDA.n219 GNDA 0.095097f
C3230 VDDA.n220 GNDA 0.12271f
C3231 VDDA.n221 GNDA 0.013706f
C3232 VDDA.n222 GNDA 0.01919f
C3233 VDDA.n225 GNDA 0.01919f
C3234 VDDA.n226 GNDA 0.01919f
C3235 VDDA.n227 GNDA 0.033381f
C3236 VDDA.n228 GNDA 0.01919f
C3237 VDDA.n229 GNDA 0.01919f
C3238 VDDA.n230 GNDA 0.01919f
C3239 VDDA.n231 GNDA 0.033583f
C3240 VDDA.t352 GNDA 0.137259f
C3241 VDDA.t388 GNDA 0.01819f
C3242 VDDA.n232 GNDA 0.047135f
C3243 VDDA.t433 GNDA 0.038309f
C3244 VDDA.t390 GNDA 0.033608f
C3245 VDDA.n233 GNDA 0.168132f
C3246 VDDA.t389 GNDA 0.116428f
C3247 VDDA.t238 GNDA 0.073881f
C3248 VDDA.t5 GNDA 0.073881f
C3249 VDDA.t432 GNDA 0.118992f
C3250 VDDA.n234 GNDA 0.176089f
C3251 VDDA.t431 GNDA 0.01819f
C3252 VDDA.n235 GNDA 0.046776f
C3253 VDDA.n236 GNDA 0.14071f
C3254 VDDA.t147 GNDA 0.028785f
C3255 VDDA.t228 GNDA 0.028785f
C3256 VDDA.n237 GNDA 0.095097f
C3257 VDDA.n238 GNDA 0.12271f
C3258 VDDA.t55 GNDA 0.028785f
C3259 VDDA.t57 GNDA 0.028785f
C3260 VDDA.n239 GNDA 0.095097f
C3261 VDDA.n240 GNDA 0.12271f
C3262 VDDA.t53 GNDA 0.028785f
C3263 VDDA.t77 GNDA 0.028785f
C3264 VDDA.n241 GNDA 0.095097f
C3265 VDDA.n242 GNDA 0.12271f
C3266 VDDA.t75 GNDA 0.028785f
C3267 VDDA.t122 GNDA 0.028785f
C3268 VDDA.n243 GNDA 0.095097f
C3269 VDDA.n244 GNDA 0.12271f
C3270 VDDA.t51 GNDA 0.028785f
C3271 VDDA.t120 GNDA 0.028785f
C3272 VDDA.n245 GNDA 0.095097f
C3273 VDDA.n246 GNDA 0.12271f
C3274 VDDA.t435 GNDA 0.028785f
C3275 VDDA.t189 GNDA 0.028785f
C3276 VDDA.n247 GNDA 0.095097f
C3277 VDDA.n248 GNDA 0.12271f
C3278 VDDA.t79 GNDA 0.028785f
C3279 VDDA.t232 GNDA 0.028785f
C3280 VDDA.n249 GNDA 0.095097f
C3281 VDDA.n250 GNDA 0.12271f
C3282 VDDA.n251 GNDA 0.065517f
C3283 VDDA.n252 GNDA 0.051261f
C3284 VDDA.n253 GNDA 0.038058f
C3285 VDDA.n254 GNDA 0.013706f
C3286 VDDA.n255 GNDA 0.033381f
C3287 VDDA.n256 GNDA 0.033583f
C3288 VDDA.n257 GNDA 0.033583f
C3289 VDDA.n258 GNDA 0.033583f
C3290 VDDA.n259 GNDA 0.048609f
C3291 VDDA.n260 GNDA 0.020196f
C3292 VDDA.n261 GNDA 0.26914f
C3293 VDDA.t353 GNDA 0.285451f
C3294 VDDA.t78 GNDA 0.293607f
C3295 VDDA.t231 GNDA 0.293607f
C3296 VDDA.t434 GNDA 0.293607f
C3297 VDDA.t188 GNDA 0.293607f
C3298 VDDA.t50 GNDA 0.293607f
C3299 VDDA.t119 GNDA 0.293607f
C3300 VDDA.t74 GNDA 0.293607f
C3301 VDDA.t121 GNDA 0.293607f
C3302 VDDA.t52 GNDA 0.293607f
C3303 VDDA.t76 GNDA 0.293607f
C3304 VDDA.t54 GNDA 0.293607f
C3305 VDDA.t56 GNDA 0.293607f
C3306 VDDA.t146 GNDA 0.293607f
C3307 VDDA.t227 GNDA 0.293607f
C3308 VDDA.t116 GNDA 0.293607f
C3309 VDDA.t222 GNDA 0.293607f
C3310 VDDA.t323 GNDA 0.285451f
C3311 VDDA.n263 GNDA 0.01919f
C3312 VDDA.n264 GNDA 0.01919f
C3313 VDDA.n265 GNDA 0.033583f
C3314 VDDA.n266 GNDA 0.033381f
C3315 VDDA.n267 GNDA 0.033583f
C3316 VDDA.n268 GNDA 0.01919f
C3317 VDDA.n269 GNDA 0.033583f
C3318 VDDA.n270 GNDA 0.033583f
C3319 VDDA.n271 GNDA 0.033381f
C3320 VDDA.n272 GNDA 0.053032f
C3321 VDDA.n273 GNDA 0.015773f
C3322 VDDA.n274 GNDA 0.26914f
C3323 VDDA.n275 GNDA 0.01919f
C3324 VDDA.n276 GNDA 0.038058f
C3325 VDDA.t322 GNDA 0.137259f
C3326 VDDA.n277 GNDA 0.051261f
C3327 VDDA.n278 GNDA 0.075592f
C3328 VDDA.t370 GNDA 0.017719f
C3329 VDDA.n279 GNDA 0.037863f
C3330 VDDA.t369 GNDA 0.033608f
C3331 VDDA.t372 GNDA 0.033608f
C3332 VDDA.n280 GNDA 0.167186f
C3333 VDDA.t371 GNDA 0.116428f
C3334 VDDA.t37 GNDA 0.073881f
C3335 VDDA.t103 GNDA 0.073881f
C3336 VDDA.t368 GNDA 0.116428f
C3337 VDDA.n281 GNDA 0.167186f
C3338 VDDA.t367 GNDA 0.017719f
C3339 VDDA.n282 GNDA 0.037863f
C3340 VDDA.n283 GNDA 0.091075f
C3341 VDDA.n284 GNDA 0.023141f
C3342 VDDA.n285 GNDA 0.081253f
C3343 VDDA.n286 GNDA 0.188662f
C3344 VDDA.n287 GNDA 0.260576f
C3345 VDDA.n288 GNDA 0.023935f
C3346 VDDA.n289 GNDA 0.084489f
C3347 VDDA.t424 GNDA 0.034982f
C3348 VDDA.t339 GNDA 0.034982f
C3349 VDDA.t337 GNDA 0.018896f
C3350 VDDA.n290 GNDA 0.02389f
C3351 VDDA.n291 GNDA 0.084533f
C3352 VDDA.t425 GNDA 0.018896f
C3353 VDDA.n292 GNDA 0.023945f
C3354 VDDA.n293 GNDA 0.084479f
C3355 VDDA.t327 GNDA 0.035f
C3356 VDDA.t405 GNDA 0.035f
C3357 VDDA.t403 GNDA 0.018896f
C3358 VDDA.n294 GNDA 0.023945f
C3359 VDDA.n295 GNDA 0.115624f
C3360 VDDA.n296 GNDA 0.040132f
C3361 VDDA.n297 GNDA 0.099877f
C3362 VDDA.t404 GNDA 0.105258f
C3363 VDDA.t25 GNDA 0.073881f
C3364 VDDA.t164 GNDA 0.073881f
C3365 VDDA.t97 GNDA 0.073881f
C3366 VDDA.t61 GNDA 0.073881f
C3367 VDDA.t326 GNDA 0.105258f
C3368 VDDA.n298 GNDA 0.099877f
C3369 VDDA.t325 GNDA 0.019495f
C3370 VDDA.n299 GNDA 0.039462f
C3371 VDDA.n300 GNDA 0.058321f
C3372 VDDA.n301 GNDA 0.02389f
C3373 VDDA.n302 GNDA 0.084533f
C3374 VDDA.n303 GNDA 0.02389f
C3375 VDDA.n304 GNDA 0.084533f
C3376 VDDA.n305 GNDA 0.02389f
C3377 VDDA.n306 GNDA 0.084533f
C3378 VDDA.n307 GNDA 0.02389f
C3379 VDDA.n308 GNDA 0.084533f
C3380 VDDA.n309 GNDA 0.058321f
C3381 VDDA.n310 GNDA 0.037331f
C3382 VDDA.t427 GNDA 0.03354f
C3383 VDDA.n311 GNDA 0.1026f
C3384 VDDA.t426 GNDA 0.105527f
C3385 VDDA.t458 GNDA 0.073881f
C3386 VDDA.t215 GNDA 0.073881f
C3387 VDDA.t130 GNDA 0.073881f
C3388 VDDA.t464 GNDA 0.073881f
C3389 VDDA.t213 GNDA 0.073881f
C3390 VDDA.t63 GNDA 0.073881f
C3391 VDDA.t128 GNDA 0.073881f
C3392 VDDA.t200 GNDA 0.073881f
C3393 VDDA.t184 GNDA 0.073881f
C3394 VDDA.t151 GNDA 0.073881f
C3395 VDDA.t398 GNDA 0.105527f
C3396 VDDA.t399 GNDA 0.03354f
C3397 VDDA.n312 GNDA 0.1026f
C3398 VDDA.t397 GNDA 0.018896f
C3399 VDDA.n313 GNDA 0.037331f
C3400 VDDA.n314 GNDA 0.058321f
C3401 VDDA.n315 GNDA 0.023935f
C3402 VDDA.n316 GNDA 0.084489f
C3403 VDDA.n317 GNDA 0.058321f
C3404 VDDA.n318 GNDA 0.038862f
C3405 VDDA.n319 GNDA 0.099896f
C3406 VDDA.t338 GNDA 0.105258f
C3407 VDDA.t39 GNDA 0.073881f
C3408 VDDA.t158 GNDA 0.073881f
C3409 VDDA.t23 GNDA 0.073881f
C3410 VDDA.t125 GNDA 0.073881f
C3411 VDDA.t423 GNDA 0.105258f
C3412 VDDA.n320 GNDA 0.099896f
C3413 VDDA.t422 GNDA 0.018896f
C3414 VDDA.n321 GNDA 0.038862f
C3415 VDDA.n322 GNDA 0.194031f
C3416 VDDA.n323 GNDA 0.226522f
C3417 VDDA.n324 GNDA 1.0799f
C3418 two_stage_opamp_dummy_magic_21_0.Vb3.t5 GNDA 0.012854f
C3419 two_stage_opamp_dummy_magic_21_0.Vb3.t3 GNDA 0.012854f
C3420 two_stage_opamp_dummy_magic_21_0.Vb3.n0 GNDA 0.041405f
C3421 two_stage_opamp_dummy_magic_21_0.Vb3.t7 GNDA 0.012854f
C3422 two_stage_opamp_dummy_magic_21_0.Vb3.t2 GNDA 0.012854f
C3423 two_stage_opamp_dummy_magic_21_0.Vb3.n1 GNDA 0.041405f
C3424 two_stage_opamp_dummy_magic_21_0.Vb3.n2 GNDA 0.228264f
C3425 two_stage_opamp_dummy_magic_21_0.Vb3.t4 GNDA 0.012854f
C3426 two_stage_opamp_dummy_magic_21_0.Vb3.t6 GNDA 0.012854f
C3427 two_stage_opamp_dummy_magic_21_0.Vb3.n3 GNDA 0.038825f
C3428 two_stage_opamp_dummy_magic_21_0.Vb3.n4 GNDA 0.69137f
C3429 two_stage_opamp_dummy_magic_21_0.Vb3.t0 GNDA 0.04499f
C3430 two_stage_opamp_dummy_magic_21_0.Vb3.t1 GNDA 0.04499f
C3431 two_stage_opamp_dummy_magic_21_0.Vb3.n5 GNDA 0.124115f
C3432 two_stage_opamp_dummy_magic_21_0.Vb3.t20 GNDA 0.063629f
C3433 two_stage_opamp_dummy_magic_21_0.Vb3.t23 GNDA 0.063629f
C3434 two_stage_opamp_dummy_magic_21_0.Vb3.t11 GNDA 0.063629f
C3435 two_stage_opamp_dummy_magic_21_0.Vb3.t8 GNDA 0.063629f
C3436 two_stage_opamp_dummy_magic_21_0.Vb3.t27 GNDA 0.073427f
C3437 two_stage_opamp_dummy_magic_21_0.Vb3.n6 GNDA 0.059615f
C3438 two_stage_opamp_dummy_magic_21_0.Vb3.n7 GNDA 0.036635f
C3439 two_stage_opamp_dummy_magic_21_0.Vb3.n8 GNDA 0.036635f
C3440 two_stage_opamp_dummy_magic_21_0.Vb3.n9 GNDA 0.032121f
C3441 two_stage_opamp_dummy_magic_21_0.Vb3.t24 GNDA 0.063629f
C3442 two_stage_opamp_dummy_magic_21_0.Vb3.t28 GNDA 0.063629f
C3443 two_stage_opamp_dummy_magic_21_0.Vb3.t9 GNDA 0.063629f
C3444 two_stage_opamp_dummy_magic_21_0.Vb3.t12 GNDA 0.063629f
C3445 two_stage_opamp_dummy_magic_21_0.Vb3.t10 GNDA 0.073427f
C3446 two_stage_opamp_dummy_magic_21_0.Vb3.n10 GNDA 0.059615f
C3447 two_stage_opamp_dummy_magic_21_0.Vb3.n11 GNDA 0.036635f
C3448 two_stage_opamp_dummy_magic_21_0.Vb3.n12 GNDA 0.036635f
C3449 two_stage_opamp_dummy_magic_21_0.Vb3.n13 GNDA 0.032121f
C3450 two_stage_opamp_dummy_magic_21_0.Vb3.n14 GNDA 0.032418f
C3451 two_stage_opamp_dummy_magic_21_0.Vb3.t22 GNDA 0.063629f
C3452 two_stage_opamp_dummy_magic_21_0.Vb3.t18 GNDA 0.063629f
C3453 two_stage_opamp_dummy_magic_21_0.Vb3.t21 GNDA 0.063629f
C3454 two_stage_opamp_dummy_magic_21_0.Vb3.t16 GNDA 0.063629f
C3455 two_stage_opamp_dummy_magic_21_0.Vb3.t13 GNDA 0.073427f
C3456 two_stage_opamp_dummy_magic_21_0.Vb3.n15 GNDA 0.059615f
C3457 two_stage_opamp_dummy_magic_21_0.Vb3.n16 GNDA 0.036635f
C3458 two_stage_opamp_dummy_magic_21_0.Vb3.n17 GNDA 0.036635f
C3459 two_stage_opamp_dummy_magic_21_0.Vb3.n18 GNDA 0.032121f
C3460 two_stage_opamp_dummy_magic_21_0.Vb3.t26 GNDA 0.063629f
C3461 two_stage_opamp_dummy_magic_21_0.Vb3.t14 GNDA 0.063629f
C3462 two_stage_opamp_dummy_magic_21_0.Vb3.t17 GNDA 0.063629f
C3463 two_stage_opamp_dummy_magic_21_0.Vb3.t15 GNDA 0.063629f
C3464 two_stage_opamp_dummy_magic_21_0.Vb3.t19 GNDA 0.073427f
C3465 two_stage_opamp_dummy_magic_21_0.Vb3.n19 GNDA 0.059615f
C3466 two_stage_opamp_dummy_magic_21_0.Vb3.n20 GNDA 0.036635f
C3467 two_stage_opamp_dummy_magic_21_0.Vb3.n21 GNDA 0.036635f
C3468 two_stage_opamp_dummy_magic_21_0.Vb3.n22 GNDA 0.032121f
C3469 two_stage_opamp_dummy_magic_21_0.Vb3.n23 GNDA 0.033008f
C3470 two_stage_opamp_dummy_magic_21_0.Vb3.n24 GNDA 1.08304f
C3471 two_stage_opamp_dummy_magic_21_0.Vb3.t25 GNDA 0.08312f
C3472 two_stage_opamp_dummy_magic_21_0.Vb3.n25 GNDA 0.29203f
C3473 two_stage_opamp_dummy_magic_21_0.Vb3.n26 GNDA 0.941369f
C3474 bgr_0.VB3_CUR_BIAS GNDA 1.43074f
C3475 bgr_0.NFET_GATE_10uA.t1 GNDA 0.01496f
C3476 bgr_0.NFET_GATE_10uA.t3 GNDA 0.01496f
C3477 bgr_0.NFET_GATE_10uA.n0 GNDA 0.042091f
C3478 bgr_0.NFET_GATE_10uA.t18 GNDA 0.014586f
C3479 bgr_0.NFET_GATE_10uA.t6 GNDA 0.014586f
C3480 bgr_0.NFET_GATE_10uA.t14 GNDA 0.014586f
C3481 bgr_0.NFET_GATE_10uA.t19 GNDA 0.014586f
C3482 bgr_0.NFET_GATE_10uA.t5 GNDA 0.014586f
C3483 bgr_0.NFET_GATE_10uA.t13 GNDA 0.014586f
C3484 bgr_0.NFET_GATE_10uA.t12 GNDA 0.021563f
C3485 bgr_0.NFET_GATE_10uA.n1 GNDA 0.026685f
C3486 bgr_0.NFET_GATE_10uA.n2 GNDA 0.019075f
C3487 bgr_0.NFET_GATE_10uA.n3 GNDA 0.016149f
C3488 bgr_0.NFET_GATE_10uA.t15 GNDA 0.014586f
C3489 bgr_0.NFET_GATE_10uA.t8 GNDA 0.014586f
C3490 bgr_0.NFET_GATE_10uA.t21 GNDA 0.014586f
C3491 bgr_0.NFET_GATE_10uA.t16 GNDA 0.021563f
C3492 bgr_0.NFET_GATE_10uA.n4 GNDA 0.026685f
C3493 bgr_0.NFET_GATE_10uA.n5 GNDA 0.019075f
C3494 bgr_0.NFET_GATE_10uA.n6 GNDA 0.016149f
C3495 bgr_0.NFET_GATE_10uA.t20 GNDA 0.014586f
C3496 bgr_0.NFET_GATE_10uA.t7 GNDA 0.021563f
C3497 bgr_0.NFET_GATE_10uA.n7 GNDA 0.02376f
C3498 bgr_0.NFET_GATE_10uA.n8 GNDA 0.026114f
C3499 bgr_0.NFET_GATE_10uA.t11 GNDA 0.014586f
C3500 bgr_0.NFET_GATE_10uA.t22 GNDA 0.021563f
C3501 bgr_0.NFET_GATE_10uA.n9 GNDA 0.02376f
C3502 bgr_0.NFET_GATE_10uA.t9 GNDA 0.014586f
C3503 bgr_0.NFET_GATE_10uA.t17 GNDA 0.014586f
C3504 bgr_0.NFET_GATE_10uA.t23 GNDA 0.014586f
C3505 bgr_0.NFET_GATE_10uA.t10 GNDA 0.021563f
C3506 bgr_0.NFET_GATE_10uA.n10 GNDA 0.026685f
C3507 bgr_0.NFET_GATE_10uA.n11 GNDA 0.019075f
C3508 bgr_0.NFET_GATE_10uA.n12 GNDA 0.016149f
C3509 bgr_0.NFET_GATE_10uA.n13 GNDA 0.026114f
C3510 bgr_0.NFET_GATE_10uA.n14 GNDA 0.605807f
C3511 bgr_0.NFET_GATE_10uA.n15 GNDA 0.022264f
C3512 bgr_0.NFET_GATE_10uA.n16 GNDA 0.016149f
C3513 bgr_0.NFET_GATE_10uA.n17 GNDA 0.019075f
C3514 bgr_0.NFET_GATE_10uA.n18 GNDA 0.026685f
C3515 bgr_0.NFET_GATE_10uA.t2 GNDA 0.034164f
C3516 bgr_0.NFET_GATE_10uA.n19 GNDA 0.327308f
C3517 bgr_0.NFET_GATE_10uA.t0 GNDA 0.01496f
C3518 bgr_0.NFET_GATE_10uA.t4 GNDA 0.01496f
C3519 bgr_0.NFET_GATE_10uA.n20 GNDA 0.088541f
.ends

