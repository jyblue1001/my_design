* PEX produced on Thu May  8 07:57:57 AM CEST 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from low_voltage_BGR_dummy_magic.ext - technology: sky130A

.subckt low_voltage_BGR_dummy_magic VDDA V_OUT GNDA
X0 GNDA.t17 a_4938_4530.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X1 VDDA.t47 V_TOP.t9 Vin-.t6 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X2 VDDA.t46 V_TOP.t10 V_OUT.t6 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X3 V_mirror.t7 V_mirror.t6 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X4 GNDA.t9 a_4938_4770.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X5 VDDA.t45 V_TOP.t11 Vin-.t4 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X6 1st_Vout.t3 V_mirror.t14 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X7 GNDA.t22 GNDA.t32 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X8 GNDA.t22 GNDA.t33 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X9 V_OUT.t2 VDDA.t31 VDDA.t32 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.6
X10 GNDA.t2 start_up.t0 start_up.t1 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=10
X11 Vin+.t5 V_TOP.t12 VDDA.t44 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X12 Vin-.t1 start_up.t3 V_TOP.t3 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X13 VDDA.t43 V_TOP.t13 start_up.t2 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X14 Vin-.t5 V_TOP.t14 VDDA.t41 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X15 GNDA.t31 GNDA.t29 V_mirror.t9 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.6
X16 V_TOP.t7 V_TOP.t6 GNDA.t14 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=4
X17 VDDA.t3 V_mirror.t4 V_mirror.t5 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X18 V_mirror.t11 Vin-.t7 V_p.t7 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X19 VDDA.t30 VDDA.t29 V_TOP.t4 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.6
X20 1st_Vout.t5 Vin+.t6 V_p.t3 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X21 V_TOP.t2 1st_Vout.t8 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X22 Vin+.t0 a_4938_3210.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X23 VDDA.t40 V_TOP.t15 Vin+.t4 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X24 1st_Vout.t2 V_mirror.t15 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X25 V_p.t6 Vin-.t8 V_mirror.t12 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X26 V_OUT.t0 a_4938_2970.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X27 VDDA.t28 VDDA.t26 V_OUT.t1 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.6
X28 VDDA.t13 1st_Vout.t9 V_TOP.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X29 a_3410_3330.t1 a_4938_3210.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X30 V_OUT.t5 V_TOP.t16 VDDA.t39 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X31 VDDA.t5 V_mirror.t2 V_mirror.t3 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X32 Vin-.t3 V_TOP.t17 VDDA.t38 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X33 a_3410_3450.t1 a_4938_3810.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X34 a_3410_3450.t0 a_4938_3090.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X35 Vin-.t0 a_4938_3090.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X36 VDDA.t37 V_TOP.t18 V_OUT.t4 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X37 GNDA.t27 GNDA.t26 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X38 VDDA.t36 V_TOP.t19 Vin+.t3 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X39 a_3410_3330.t0 a_4938_3930.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X40 a_3410_3570.t0 a_4938_2970.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X41 V_mirror.t10 Vin-.t9 V_p.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X42 a_3410_3570.t1 a_4938_3690.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X43 a_3410_4410.t1 a_4938_3690.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t0 Vin+.t1 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X45 V_p.t2 Vin+.t7 1st_Vout.t4 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X46 GNDA.t7 V_p.t8 V_p.t9 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=4
X47 V_mirror.t1 V_mirror.t0 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X48 V_p.t4 Vin-.t10 V_mirror.t13 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X49 GNDA.t22 GNDA.t25 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X50 GNDA.t22 GNDA.t21 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X51 a_3410_4410.t0 a_4938_4530.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X52 a_3410_4170.t0 a_4938_3930.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X53 V_TOP.t8 1st_Vout.t10 VDDA.t48 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X54 V_p.t1 Vin+.t8 1st_Vout.t7 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X55 GNDA.t27 GNDA.t28 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X56 GNDA.t24 GNDA.t23 Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X57 a_3410_4290.t0 a_4938_4650.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X58 VDDA.t18 V_mirror.t16 1st_Vout.t1 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X59 V_mirror.t8 GNDA.t18 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.6
X60 Vin+.t2 V_TOP.t20 VDDA.t35 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X61 a_3410_4290.t1 a_4938_3810.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X62 VDDA.t22 1st_Vout.t11 V_TOP.t5 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X63 1st_Vout.t6 Vin+.t9 V_p.t0 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X64 GNDA.t34 a_4938_4650.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X65 V_OUT.t3 V_TOP.t21 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X66 VDDA.t9 V_mirror.t17 1st_Vout.t0 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X67 a_3410_4170.t1 a_4938_4770.t1 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X68 V_TOP.t0 VDDA.t23 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.6
R0 GNDA.n1004 GNDA.n964 50274.2
R1 GNDA.n939 GNDA.n595 2115.21
R2 GNDA.n940 GNDA.n939 2079.51
R3 GNDA.n1557 GNDA.t27 1668.97
R4 GNDA.t27 GNDA.n1556 1633.27
R5 GNDA.n1582 GNDA.n1581 1600.21
R6 GNDA.n529 GNDA.n528 1497.38
R7 GNDA.n964 GNDA.t3 1259.74
R8 GNDA.n1353 GNDA.n1352 1214.72
R9 GNDA.n1352 GNDA.n1351 1214.72
R10 GNDA.n1351 GNDA.n1067 1214.72
R11 GNDA.n1269 GNDA.n1067 1214.72
R12 GNDA.n1269 GNDA.n24 1214.72
R13 GNDA.n1283 GNDA.n25 1214.72
R14 GNDA.n1283 GNDA.n1246 1214.72
R15 GNDA.n1289 GNDA.n1246 1214.72
R16 GNDA.n1290 GNDA.n1289 1214.72
R17 GNDA.n1290 GNDA.n26 1214.72
R18 GNDA.t19 GNDA.n964 1001.38
R19 GNDA.t22 GNDA.n22 949.682
R20 GNDA.n1607 GNDA.t22 949.682
R21 GNDA.t22 GNDA.n25 823.313
R22 GNDA.n962 GNDA.n581 803.245
R23 GNDA.n957 GNDA.n581 803.245
R24 GNDA.n957 GNDA.n956 803.245
R25 GNDA.n956 GNDA.n955 803.245
R26 GNDA.n955 GNDA.n578 803.245
R27 GNDA.n948 GNDA.n577 803.245
R28 GNDA.n948 GNDA.n947 803.245
R29 GNDA.n947 GNDA.n946 803.245
R30 GNDA.n946 GNDA.n590 803.245
R31 GNDA.n940 GNDA.n590 803.245
R32 GNDA.n608 GNDA.n595 803.245
R33 GNDA.n730 GNDA.n608 803.245
R34 GNDA.n731 GNDA.n730 803.245
R35 GNDA.n732 GNDA.n731 803.245
R36 GNDA.n732 GNDA.n602 803.245
R37 GNDA.n745 GNDA.n603 803.245
R38 GNDA.n739 GNDA.n603 803.245
R39 GNDA.n739 GNDA.n738 803.245
R40 GNDA.n738 GNDA.n65 803.245
R41 GNDA.n1556 GNDA.n65 803.245
R42 GNDA.n1558 GNDA.n1557 803.245
R43 GNDA.n1558 GNDA.n58 803.245
R44 GNDA.n1565 GNDA.n58 803.245
R45 GNDA.n1566 GNDA.n1565 803.245
R46 GNDA.n1567 GNDA.n1566 803.245
R47 GNDA.n1573 GNDA.n54 803.245
R48 GNDA.n1574 GNDA.n1573 803.245
R49 GNDA.n1575 GNDA.n1574 803.245
R50 GNDA.n1575 GNDA.n50 803.245
R51 GNDA.n1581 GNDA.n50 803.245
R52 GNDA.n1002 GNDA.n1001 686.717
R53 GNDA.n1011 GNDA.n1010 669.307
R54 GNDA.t22 GNDA.n21 623.755
R55 GNDA.t22 GNDA.n1606 623.755
R56 GNDA.n882 GNDA.n580 593.867
R57 GNDA.n110 GNDA.n109 588.271
R58 GNDA.n1005 GNDA.n1004 585.003
R59 GNDA.n971 GNDA.n969 585
R60 GNDA.n998 GNDA.n968 585
R61 GNDA.n1003 GNDA.n968 585
R62 GNDA.n997 GNDA.n996 585
R63 GNDA.n995 GNDA.n994 585
R64 GNDA.n993 GNDA.n976 585
R65 GNDA.n989 GNDA.n988 585
R66 GNDA.n985 GNDA.n967 585
R67 GNDA.n1003 GNDA.n967 585
R68 GNDA.n1388 GNDA.n1387 585
R69 GNDA.n107 GNDA.n106 585
R70 GNDA.n1456 GNDA.n1455 585
R71 GNDA.n1458 GNDA.n105 585
R72 GNDA.n1461 GNDA.n1460 585
R73 GNDA.n102 GNDA.n101 585
R74 GNDA.n1471 GNDA.n1470 585
R75 GNDA.n1473 GNDA.n100 585
R76 GNDA.n1476 GNDA.n1475 585
R77 GNDA.n97 GNDA.n93 585
R78 GNDA.n1487 GNDA.n1486 585
R79 GNDA.n1489 GNDA.n92 585
R80 GNDA.n885 GNDA.n884 585
R81 GNDA.n880 GNDA.n879 585
R82 GNDA.n880 GNDA.n576 585
R83 GNDA.n878 GNDA.n759 585
R84 GNDA.n876 GNDA.n875 585
R85 GNDA.n873 GNDA.n872 585
R86 GNDA.n791 GNDA.n763 585
R87 GNDA.n795 GNDA.n794 585
R88 GNDA.n797 GNDA.n790 585
R89 GNDA.n800 GNDA.n799 585
R90 GNDA.n786 GNDA.n785 585
R91 GNDA.n810 GNDA.n809 585
R92 GNDA.n812 GNDA.n782 585
R93 GNDA.n815 GNDA.n814 585
R94 GNDA.n783 GNDA.n582 585
R95 GNDA.n594 GNDA.n593 585
R96 GNDA.n915 GNDA.n912 585
R97 GNDA.n917 GNDA.n916 585
R98 GNDA.n918 GNDA.n911 585
R99 GNDA.n920 GNDA.n919 585
R100 GNDA.n922 GNDA.n909 585
R101 GNDA.n924 GNDA.n923 585
R102 GNDA.n925 GNDA.n908 585
R103 GNDA.n927 GNDA.n926 585
R104 GNDA.n929 GNDA.n906 585
R105 GNDA.n931 GNDA.n930 585
R106 GNDA.n932 GNDA.n749 585
R107 GNDA.n905 GNDA.n748 585
R108 GNDA.n748 GNDA.n747 585
R109 GNDA.n904 GNDA.n903 585
R110 GNDA.n903 GNDA.n902 585
R111 GNDA.n751 GNDA.n750 585
R112 GNDA.n901 GNDA.n751 585
R113 GNDA.n899 GNDA.n898 585
R114 GNDA.n900 GNDA.n899 585
R115 GNDA.n897 GNDA.n753 585
R116 GNDA.n753 GNDA.n752 585
R117 GNDA.n896 GNDA.n895 585
R118 GNDA.n895 GNDA.n894 585
R119 GNDA.n755 GNDA.n754 585
R120 GNDA.n893 GNDA.n755 585
R121 GNDA.n891 GNDA.n890 585
R122 GNDA.n892 GNDA.n891 585
R123 GNDA.n889 GNDA.n757 585
R124 GNDA.n757 GNDA.n756 585
R125 GNDA.n888 GNDA.n887 585
R126 GNDA.n887 GNDA.n886 585
R127 GNDA.n937 GNDA.n936 585
R128 GNDA.n938 GNDA.n937 585
R129 GNDA.n1525 GNDA.n1524 585
R130 GNDA.n1522 GNDA.n80 585
R131 GNDA.n1521 GNDA.n81 585
R132 GNDA.n1519 GNDA.n1518 585
R133 GNDA.n83 GNDA.n82 585
R134 GNDA.n1510 GNDA.n1509 585
R135 GNDA.n1507 GNDA.n85 585
R136 GNDA.n1505 GNDA.n1504 585
R137 GNDA.n87 GNDA.n86 585
R138 GNDA.n1498 GNDA.n1497 585
R139 GNDA.n1495 GNDA.n89 585
R140 GNDA.n1493 GNDA.n1492 585
R141 GNDA.n934 GNDA.n933 585
R142 GNDA.n933 GNDA.n31 585
R143 GNDA.n75 GNDA.n74 585
R144 GNDA.n74 GNDA.n62 585
R145 GNDA.n1526 GNDA.n1525 585
R146 GNDA.n1514 GNDA.n80 585
R147 GNDA.n1515 GNDA.n81 585
R148 GNDA.n1518 GNDA.n1517 585
R149 GNDA.n1513 GNDA.n83 585
R150 GNDA.n1511 GNDA.n1510 585
R151 GNDA.n85 GNDA.n84 585
R152 GNDA.n1504 GNDA.n1503 585
R153 GNDA.n1501 GNDA.n87 585
R154 GNDA.n1499 GNDA.n1498 585
R155 GNDA.n89 GNDA.n88 585
R156 GNDA.n1492 GNDA.n1491 585
R157 GNDA.n690 GNDA.n689 585
R158 GNDA.n693 GNDA.n692 585
R159 GNDA.n695 GNDA.n694 585
R160 GNDA.n699 GNDA.n698 585
R161 GNDA.n697 GNDA.n616 585
R162 GNDA.n706 GNDA.n705 585
R163 GNDA.n708 GNDA.n707 585
R164 GNDA.n712 GNDA.n711 585
R165 GNDA.n710 GNDA.n612 585
R166 GNDA.n719 GNDA.n718 585
R167 GNDA.n721 GNDA.n720 585
R168 GNDA.n724 GNDA.n723 585
R169 GNDA.n1553 GNDA.n67 585
R170 GNDA.n1552 GNDA.n1551 585
R171 GNDA.n1549 GNDA.n69 585
R172 GNDA.n1547 GNDA.n1546 585
R173 GNDA.n1545 GNDA.n70 585
R174 GNDA.n1544 GNDA.n1543 585
R175 GNDA.n1541 GNDA.n71 585
R176 GNDA.n1539 GNDA.n1538 585
R177 GNDA.n1537 GNDA.n72 585
R178 GNDA.n1536 GNDA.n1535 585
R179 GNDA.n1533 GNDA.n73 585
R180 GNDA.n1531 GNDA.n1530 585
R181 GNDA.n942 GNDA.n941 585
R182 GNDA.n941 GNDA.n940 585
R183 GNDA.n943 GNDA.n591 585
R184 GNDA.n591 GNDA.n590 585
R185 GNDA.n945 GNDA.n944 585
R186 GNDA.n946 GNDA.n945 585
R187 GNDA.n592 GNDA.n589 585
R188 GNDA.n947 GNDA.n589 585
R189 GNDA.n949 GNDA.n588 585
R190 GNDA.n949 GNDA.n948 585
R191 GNDA.n951 GNDA.n950 585
R192 GNDA.n950 GNDA.n577 585
R193 GNDA.n952 GNDA.n586 585
R194 GNDA.n586 GNDA.n578 585
R195 GNDA.n954 GNDA.n953 585
R196 GNDA.n955 GNDA.n954 585
R197 GNDA.n587 GNDA.n584 585
R198 GNDA.n956 GNDA.n584 585
R199 GNDA.n958 GNDA.n585 585
R200 GNDA.n958 GNDA.n957 585
R201 GNDA.n959 GNDA.n581 585
R202 GNDA.n962 GNDA.n961 585
R203 GNDA.n1555 GNDA.n1554 585
R204 GNDA.n1556 GNDA.n1555 585
R205 GNDA.n68 GNDA.n66 585
R206 GNDA.n66 GNDA.n65 585
R207 GNDA.n737 GNDA.n736 585
R208 GNDA.n738 GNDA.n737 585
R209 GNDA.n741 GNDA.n740 585
R210 GNDA.n740 GNDA.n739 585
R211 GNDA.n742 GNDA.n605 585
R212 GNDA.n605 GNDA.n603 585
R213 GNDA.n744 GNDA.n743 585
R214 GNDA.n745 GNDA.n744 585
R215 GNDA.n735 GNDA.n604 585
R216 GNDA.n604 GNDA.n602 585
R217 GNDA.n734 GNDA.n733 585
R218 GNDA.n733 GNDA.n732 585
R219 GNDA.n607 GNDA.n606 585
R220 GNDA.n731 GNDA.n607 585
R221 GNDA.n729 GNDA.n728 585
R222 GNDA.n730 GNDA.n729 585
R223 GNDA.n609 GNDA.n608 585
R224 GNDA.n725 GNDA.n595 585
R225 GNDA.n1580 GNDA.n1579 585
R226 GNDA.n1581 GNDA.n1580 585
R227 GNDA.n1578 GNDA.n51 585
R228 GNDA.n51 GNDA.n50 585
R229 GNDA.n1577 GNDA.n1576 585
R230 GNDA.n1576 GNDA.n1575 585
R231 GNDA.n53 GNDA.n52 585
R232 GNDA.n1574 GNDA.n53 585
R233 GNDA.n1572 GNDA.n1571 585
R234 GNDA.n1573 GNDA.n1572 585
R235 GNDA.n1570 GNDA.n55 585
R236 GNDA.n55 GNDA.n54 585
R237 GNDA.n1569 GNDA.n1568 585
R238 GNDA.n1568 GNDA.n1567 585
R239 GNDA.n57 GNDA.n56 585
R240 GNDA.n1566 GNDA.n57 585
R241 GNDA.n1564 GNDA.n1563 585
R242 GNDA.n1565 GNDA.n1564 585
R243 GNDA.n1562 GNDA.n59 585
R244 GNDA.n59 GNDA.n58 585
R245 GNDA.n49 GNDA.n48 585
R246 GNDA.n1582 GNDA.n49 585
R247 GNDA.n1585 GNDA.n1584 585
R248 GNDA.n1584 GNDA.n1583 585
R249 GNDA.n1586 GNDA.n47 585
R250 GNDA.n47 GNDA.n46 585
R251 GNDA.n1588 GNDA.n1587 585
R252 GNDA.n1589 GNDA.n1588 585
R253 GNDA.n45 GNDA.n44 585
R254 GNDA.n1590 GNDA.n45 585
R255 GNDA.n1593 GNDA.n1592 585
R256 GNDA.n1592 GNDA.n1591 585
R257 GNDA.n1594 GNDA.n43 585
R258 GNDA.n43 GNDA.n42 585
R259 GNDA.n1596 GNDA.n1595 585
R260 GNDA.n1597 GNDA.n1596 585
R261 GNDA.n40 GNDA.n39 585
R262 GNDA.n1598 GNDA.n40 585
R263 GNDA.n1601 GNDA.n1600 585
R264 GNDA.n1600 GNDA.n1599 585
R265 GNDA.n1602 GNDA.n37 585
R266 GNDA.n41 GNDA.n37 585
R267 GNDA.n1604 GNDA.n1603 585
R268 GNDA.n1604 GNDA.n36 585
R269 GNDA.n551 GNDA.n355 585
R270 GNDA.n355 GNDA.n22 585
R271 GNDA.n550 GNDA.n549 585
R272 GNDA.n549 GNDA.n548 585
R273 GNDA.n360 GNDA.n359 585
R274 GNDA.n547 GNDA.n360 585
R275 GNDA.n545 GNDA.n544 585
R276 GNDA.n546 GNDA.n545 585
R277 GNDA.n543 GNDA.n362 585
R278 GNDA.n362 GNDA.n361 585
R279 GNDA.n542 GNDA.n541 585
R280 GNDA.n541 GNDA.n18 585
R281 GNDA.n540 GNDA.n363 585
R282 GNDA.n540 GNDA.n19 585
R283 GNDA.n539 GNDA.n365 585
R284 GNDA.n539 GNDA.n538 585
R285 GNDA.n533 GNDA.n364 585
R286 GNDA.n537 GNDA.n364 585
R287 GNDA.n535 GNDA.n534 585
R288 GNDA.n536 GNDA.n535 585
R289 GNDA.n532 GNDA.n367 585
R290 GNDA.n367 GNDA.n366 585
R291 GNDA.n531 GNDA.n530 585
R292 GNDA.n530 GNDA.n529 585
R293 GNDA.n503 GNDA.n381 585
R294 GNDA.n501 GNDA.n500 585
R295 GNDA.n388 GNDA.n386 585
R296 GNDA.n469 GNDA.n467 585
R297 GNDA.n476 GNDA.n475 585
R298 GNDA.n478 GNDA.n465 585
R299 GNDA.n481 GNDA.n480 585
R300 GNDA.n463 GNDA.n462 585
R301 GNDA.n488 GNDA.n487 585
R302 GNDA.n490 GNDA.n410 585
R303 GNDA.n493 GNDA.n492 585
R304 GNDA.n333 GNDA.n330 585
R305 GNDA.n385 GNDA.n384 585
R306 GNDA.n383 GNDA.n382 585
R307 GNDA.n508 GNDA.n379 585
R308 GNDA.n379 GNDA.n378 585
R309 GNDA.n510 GNDA.n509 585
R310 GNDA.n511 GNDA.n510 585
R311 GNDA.n377 GNDA.n376 585
R312 GNDA.n512 GNDA.n377 585
R313 GNDA.n515 GNDA.n514 585
R314 GNDA.n514 GNDA.n513 585
R315 GNDA.n516 GNDA.n375 585
R316 GNDA.n375 GNDA.n374 585
R317 GNDA.n518 GNDA.n517 585
R318 GNDA.n519 GNDA.n518 585
R319 GNDA.n373 GNDA.n372 585
R320 GNDA.n520 GNDA.n373 585
R321 GNDA.n523 GNDA.n522 585
R322 GNDA.n522 GNDA.n521 585
R323 GNDA.n524 GNDA.n371 585
R324 GNDA.n371 GNDA.n370 585
R325 GNDA.n526 GNDA.n525 585
R326 GNDA.n527 GNDA.n526 585
R327 GNDA.n506 GNDA.n505 585
R328 GNDA.n505 GNDA.n15 585
R329 GNDA.n369 GNDA.n368 585
R330 GNDA.n528 GNDA.n369 585
R331 GNDA.n280 GNDA.n279 585
R332 GNDA.n151 GNDA.n29 585
R333 GNDA.n276 GNDA.n275 585
R334 GNDA.n275 GNDA.n31 585
R335 GNDA.n273 GNDA.n152 585
R336 GNDA.n271 GNDA.n270 585
R337 GNDA.n155 GNDA.n153 585
R338 GNDA.n236 GNDA.n234 585
R339 GNDA.n243 GNDA.n242 585
R340 GNDA.n245 GNDA.n232 585
R341 GNDA.n248 GNDA.n247 585
R342 GNDA.n230 GNDA.n229 585
R343 GNDA.n255 GNDA.n254 585
R344 GNDA.n257 GNDA.n177 585
R345 GNDA.n263 GNDA.n262 585
R346 GNDA.n260 GNDA.n259 585
R347 GNDA.n301 GNDA.n300 585
R348 GNDA.n300 GNDA.n299 585
R349 GNDA.n143 GNDA.n142 585
R350 GNDA.n298 GNDA.n143 585
R351 GNDA.n296 GNDA.n295 585
R352 GNDA.n297 GNDA.n296 585
R353 GNDA.n294 GNDA.n145 585
R354 GNDA.n145 GNDA.n144 585
R355 GNDA.n293 GNDA.n292 585
R356 GNDA.n292 GNDA.n291 585
R357 GNDA.n286 GNDA.n146 585
R358 GNDA.n290 GNDA.n146 585
R359 GNDA.n288 GNDA.n287 585
R360 GNDA.n289 GNDA.n288 585
R361 GNDA.n285 GNDA.n148 585
R362 GNDA.n148 GNDA.n147 585
R363 GNDA.n284 GNDA.n283 585
R364 GNDA.n283 GNDA.n282 585
R365 GNDA.n150 GNDA.n149 585
R366 GNDA.n281 GNDA.n150 585
R367 GNDA.n302 GNDA.n141 585
R368 GNDA.n141 GNDA.n16 585
R369 GNDA.n326 GNDA.n132 585
R370 GNDA.n325 GNDA.n324 585
R371 GNDA.n322 GNDA.n136 585
R372 GNDA.n320 GNDA.n319 585
R373 GNDA.n318 GNDA.n137 585
R374 GNDA.n317 GNDA.n316 585
R375 GNDA.n314 GNDA.n138 585
R376 GNDA.n312 GNDA.n311 585
R377 GNDA.n310 GNDA.n139 585
R378 GNDA.n309 GNDA.n308 585
R379 GNDA.n306 GNDA.n140 585
R380 GNDA.n304 GNDA.n303 585
R381 GNDA.n1528 GNDA.n1527 585
R382 GNDA.n1527 GNDA.n26 585
R383 GNDA.n78 GNDA.n77 585
R384 GNDA.n1290 GNDA.n78 585
R385 GNDA.n1288 GNDA.n1287 585
R386 GNDA.n1289 GNDA.n1288 585
R387 GNDA.n1286 GNDA.n1247 585
R388 GNDA.n1247 GNDA.n1246 585
R389 GNDA.n1285 GNDA.n1284 585
R390 GNDA.n1284 GNDA.n1283 585
R391 GNDA.n1249 GNDA.n1248 585
R392 GNDA.n1249 GNDA.n25 585
R393 GNDA.n1266 GNDA.n1261 585
R394 GNDA.n1261 GNDA.n24 585
R395 GNDA.n1268 GNDA.n1267 585
R396 GNDA.n1269 GNDA.n1268 585
R397 GNDA.n1265 GNDA.n1260 585
R398 GNDA.n1260 GNDA.n1067 585
R399 GNDA.n1264 GNDA.n1066 585
R400 GNDA.n1351 GNDA.n1066 585
R401 GNDA.n1263 GNDA.n1065 585
R402 GNDA.n1352 GNDA.n1065 585
R403 GNDA.n1262 GNDA.n328 585
R404 GNDA.n1353 GNDA.n328 585
R405 GNDA.n1362 GNDA.n135 585
R406 GNDA.n133 GNDA.n130 585
R407 GNDA.n1367 GNDA.n129 585
R408 GNDA.n1368 GNDA.n127 585
R409 GNDA.n1369 GNDA.n126 585
R410 GNDA.n124 GNDA.n121 585
R411 GNDA.n1374 GNDA.n120 585
R412 GNDA.n1375 GNDA.n118 585
R413 GNDA.n1376 GNDA.n117 585
R414 GNDA.n113 GNDA.n112 585
R415 GNDA.n1382 GNDA.n1381 585
R416 GNDA.n1384 GNDA.n111 585
R417 GNDA.n110 GNDA.n31 585
R418 GNDA.n1361 GNDA.n1360 585
R419 GNDA.n1360 GNDA.n1359 585
R420 GNDA.n1363 GNDA.n1362 585
R421 GNDA.n1365 GNDA.n130 585
R422 GNDA.n1367 GNDA.n1366 585
R423 GNDA.n1368 GNDA.n123 585
R424 GNDA.n1370 GNDA.n1369 585
R425 GNDA.n1372 GNDA.n121 585
R426 GNDA.n1374 GNDA.n1373 585
R427 GNDA.n1375 GNDA.n115 585
R428 GNDA.n1377 GNDA.n1376 585
R429 GNDA.n1379 GNDA.n113 585
R430 GNDA.n1381 GNDA.n1380 585
R431 GNDA.n258 GNDA.n111 585
R432 GNDA.n1041 GNDA.n358 585
R433 GNDA.n356 GNDA.n353 585
R434 GNDA.n1046 GNDA.n352 585
R435 GNDA.n1047 GNDA.n350 585
R436 GNDA.n1048 GNDA.n349 585
R437 GNDA.n347 GNDA.n344 585
R438 GNDA.n1053 GNDA.n343 585
R439 GNDA.n1054 GNDA.n341 585
R440 GNDA.n1055 GNDA.n340 585
R441 GNDA.n338 GNDA.n334 585
R442 GNDA.n337 GNDA.n332 585
R443 GNDA.n1062 GNDA.n331 585
R444 GNDA.n1358 GNDA.n1357 585
R445 GNDA.n1359 GNDA.n1358 585
R446 GNDA.n1040 GNDA.n1039 585
R447 GNDA.n1039 GNDA.n21 585
R448 GNDA.n1042 GNDA.n1041 585
R449 GNDA.n1044 GNDA.n353 585
R450 GNDA.n1046 GNDA.n1045 585
R451 GNDA.n1047 GNDA.n346 585
R452 GNDA.n1049 GNDA.n1048 585
R453 GNDA.n1051 GNDA.n344 585
R454 GNDA.n1053 GNDA.n1052 585
R455 GNDA.n1054 GNDA.n335 585
R456 GNDA.n1056 GNDA.n1055 585
R457 GNDA.n1058 GNDA.n334 585
R458 GNDA.n1059 GNDA.n332 585
R459 GNDA.n1062 GNDA.n1061 585
R460 GNDA.n1355 GNDA.n1354 585
R461 GNDA.n1354 GNDA.n1353 585
R462 GNDA.n1069 GNDA.n1064 585
R463 GNDA.n1352 GNDA.n1064 585
R464 GNDA.n1350 GNDA.n1349 585
R465 GNDA.n1351 GNDA.n1350 585
R466 GNDA.n1071 GNDA.n1068 585
R467 GNDA.n1068 GNDA.n1067 585
R468 GNDA.n1270 GNDA.n1259 585
R469 GNDA.n1270 GNDA.n1269 585
R470 GNDA.n1272 GNDA.n1271 585
R471 GNDA.n1271 GNDA.n24 585
R472 GNDA.n1273 GNDA.n1250 585
R473 GNDA.n1250 GNDA.n25 585
R474 GNDA.n1282 GNDA.n1281 585
R475 GNDA.n1283 GNDA.n1282 585
R476 GNDA.n1254 GNDA.n1251 585
R477 GNDA.n1251 GNDA.n1246 585
R478 GNDA.n1093 GNDA.n1091 585
R479 GNDA.n1289 GNDA.n1093 585
R480 GNDA.n1292 GNDA.n1291 585
R481 GNDA.n1291 GNDA.n1290 585
R482 GNDA.n1245 GNDA.n1244 585
R483 GNDA.n1245 GNDA.n26 585
R484 GNDA.n1214 GNDA.n1095 585
R485 GNDA.n1212 GNDA.n1211 585
R486 GNDA.n1098 GNDA.n1096 585
R487 GNDA.n1179 GNDA.n1177 585
R488 GNDA.n1186 GNDA.n1185 585
R489 GNDA.n1188 GNDA.n1175 585
R490 GNDA.n1191 GNDA.n1190 585
R491 GNDA.n1173 GNDA.n1172 585
R492 GNDA.n1198 GNDA.n1197 585
R493 GNDA.n1200 GNDA.n1120 585
R494 GNDA.n1204 GNDA.n1203 585
R495 GNDA.n1201 GNDA.n60 585
R496 GNDA.n1559 GNDA.n1558 585
R497 GNDA.n1557 GNDA.n61 585
R498 GNDA.n1610 GNDA.n9 585
R499 GNDA.n1611 GNDA.n8 585
R500 GNDA.n1612 GNDA.n7 585
R501 GNDA.n32 GNDA.n3 585
R502 GNDA.n1617 GNDA.n2 585
R503 GNDA.n1228 GNDA.n1 585
R504 GNDA.n1234 GNDA.n1230 585
R505 GNDA.n1235 GNDA.n1226 585
R506 GNDA.n1236 GNDA.n1225 585
R507 GNDA.n1223 GNDA.n1220 585
R508 GNDA.n1241 GNDA.n1219 585
R509 GNDA.n1242 GNDA.n1217 585
R510 GNDA.n1215 GNDA.n76 585
R511 GNDA.n1215 GNDA.n62 585
R512 GNDA.n1605 GNDA.n10 585
R513 GNDA.n1606 GNDA.n1605 585
R514 GNDA.n1610 GNDA.n1609 585
R515 GNDA.n1611 GNDA.n6 585
R516 GNDA.n1613 GNDA.n1612 585
R517 GNDA.n1615 GNDA.n3 585
R518 GNDA.n1617 GNDA.n1616 585
R519 GNDA.n1232 GNDA.n1 585
R520 GNDA.n1234 GNDA.n1233 585
R521 GNDA.n1235 GNDA.n1222 585
R522 GNDA.n1237 GNDA.n1236 585
R523 GNDA.n1239 GNDA.n1220 585
R524 GNDA.n1241 GNDA.n1240 585
R525 GNDA.n1242 GNDA.n1094 585
R526 GNDA.n1608 GNDA.n13 585
R527 GNDA.n1608 GNDA.n1607 585
R528 GNDA.n1016 GNDA.n12 585
R529 GNDA.n14 GNDA.n12 585
R530 GNDA.n1018 GNDA.n1017 585
R531 GNDA.n1020 GNDA.n1018 585
R532 GNDA.n1023 GNDA.n1022 585
R533 GNDA.n1022 GNDA.n1021 585
R534 GNDA.n1024 GNDA.n559 585
R535 GNDA.n1019 GNDA.n559 585
R536 GNDA.n1026 GNDA.n1025 585
R537 GNDA.n1026 GNDA.n28 585
R538 GNDA.n1027 GNDA.n558 585
R539 GNDA.n1028 GNDA.n1027 585
R540 GNDA.n1031 GNDA.n1030 585
R541 GNDA.n1030 GNDA.n1029 585
R542 GNDA.n1032 GNDA.n556 585
R543 GNDA.n556 GNDA.n555 585
R544 GNDA.n1034 GNDA.n1033 585
R545 GNDA.n1035 GNDA.n1034 585
R546 GNDA.n557 GNDA.n553 585
R547 GNDA.n1036 GNDA.n553 585
R548 GNDA.n1038 GNDA.n554 585
R549 GNDA.n1038 GNDA.n1037 585
R550 GNDA.n1012 GNDA.n560 585
R551 GNDA.n1014 GNDA.n1013 585
R552 GNDA.n1013 GNDA.n27 585
R553 GNDA.n939 GNDA.n579 582.98
R554 GNDA.n939 GNDA.n746 578.723
R555 GNDA.n1353 GNDA.t22 512.884
R556 GNDA.n529 GNDA.n366 505.748
R557 GNDA.n536 GNDA.n366 505.748
R558 GNDA.n537 GNDA.n536 505.748
R559 GNDA.n538 GNDA.n537 505.748
R560 GNDA.n538 GNDA.n19 505.748
R561 GNDA.n361 GNDA.n18 505.748
R562 GNDA.n546 GNDA.n361 505.748
R563 GNDA.n547 GNDA.n546 505.748
R564 GNDA.n548 GNDA.n547 505.748
R565 GNDA.n548 GNDA.n22 505.748
R566 GNDA.n1037 GNDA.n21 505.748
R567 GNDA.n1037 GNDA.n1036 505.748
R568 GNDA.n1036 GNDA.n1035 505.748
R569 GNDA.n1035 GNDA.n555 505.748
R570 GNDA.n1029 GNDA.n555 505.748
R571 GNDA.n1029 GNDA.n1028 505.748
R572 GNDA.n1019 GNDA.n28 505.748
R573 GNDA.n1021 GNDA.n1019 505.748
R574 GNDA.n1021 GNDA.n1020 505.748
R575 GNDA.n1020 GNDA.n14 505.748
R576 GNDA.n1607 GNDA.n14 505.748
R577 GNDA.n1606 GNDA.n36 505.748
R578 GNDA.n41 GNDA.n36 505.748
R579 GNDA.n1599 GNDA.n41 505.748
R580 GNDA.n1599 GNDA.n1598 505.748
R581 GNDA.n1598 GNDA.n1597 505.748
R582 GNDA.n1597 GNDA.n42 505.748
R583 GNDA.n1591 GNDA.n1590 505.748
R584 GNDA.n1590 GNDA.n1589 505.748
R585 GNDA.n1589 GNDA.n46 505.748
R586 GNDA.n1583 GNDA.n46 505.748
R587 GNDA.n1583 GNDA.n1582 505.748
R588 GNDA.t24 GNDA.n577 419.474
R589 GNDA.t27 GNDA.n745 419.474
R590 GNDA.n54 GNDA.t27 419.474
R591 GNDA.n384 GNDA.n15 410.342
R592 GNDA.t22 GNDA.n24 391.411
R593 GNDA.n299 GNDA.n16 390.029
R594 GNDA.n528 GNDA.n527 390.029
R595 GNDA.t24 GNDA.n578 383.774
R596 GNDA.t27 GNDA.n602 383.774
R597 GNDA.n1567 GNDA.t27 383.774
R598 GNDA.n280 GNDA.n29 365.651
R599 GNDA.n281 GNDA.n280 365.651
R600 GNDA.n282 GNDA.n281 365.651
R601 GNDA.n282 GNDA.n147 365.651
R602 GNDA.n289 GNDA.n147 365.651
R603 GNDA.n291 GNDA.n290 365.651
R604 GNDA.n291 GNDA.n144 365.651
R605 GNDA.n297 GNDA.n144 365.651
R606 GNDA.n298 GNDA.n297 365.651
R607 GNDA.n299 GNDA.n298 365.651
R608 GNDA.n384 GNDA.n383 365.651
R609 GNDA.n383 GNDA.n378 365.651
R610 GNDA.n511 GNDA.n378 365.651
R611 GNDA.n512 GNDA.n511 365.651
R612 GNDA.n513 GNDA.n512 365.651
R613 GNDA.n519 GNDA.n374 365.651
R614 GNDA.n520 GNDA.n519 365.651
R615 GNDA.n521 GNDA.n520 365.651
R616 GNDA.n521 GNDA.n370 365.651
R617 GNDA.n527 GNDA.n370 365.651
R618 GNDA.t22 GNDA.n16 353.464
R619 GNDA.t22 GNDA.n15 349.401
R620 GNDA.t22 GNDA.n18 342.784
R621 GNDA.t22 GNDA.n28 342.784
R622 GNDA.n1591 GNDA.t27 342.784
R623 GNDA.n1001 GNDA.n970 335
R624 GNDA.n987 GNDA.n985 335
R625 GNDA.n746 GNDA.t27 327.661
R626 GNDA.n64 GNDA.t27 172.876
R627 GNDA.t24 GNDA.n579 323.404
R628 GNDA.t27 GNDA.n63 172.615
R629 GNDA.n1004 GNDA.t30 303.449
R630 GNDA.t30 GNDA.t4 303.449
R631 GNDA.t15 GNDA.t8 303.449
R632 GNDA.t8 GNDA.t10 303.449
R633 GNDA.t12 GNDA.t0 303.449
R634 GNDA.t0 GNDA.t11 303.449
R635 GNDA.t5 GNDA.t19 303.449
R636 GNDA.t4 GNDA.t13 273.103
R637 GNDA.t6 GNDA.t5 273.103
R638 GNDA.n1000 GNDA.n999 267.865
R639 GNDA.n991 GNDA.n990 267.865
R640 GNDA.n1154 GNDA.n1109 258.334
R641 GNDA.n1312 GNDA.n1084 258.334
R642 GNDA.n444 GNDA.n399 258.334
R643 GNDA.n656 GNDA.n634 258.334
R644 GNDA.n1418 GNDA.n1400 258.334
R645 GNDA.n835 GNDA.n775 258.334
R646 GNDA.n211 GNDA.n166 258.334
R647 GNDA.n1245 GNDA.n1094 257.466
R648 GNDA.n1201 GNDA.n61 257.466
R649 GNDA.n725 GNDA.n724 257.466
R650 GNDA.n1491 GNDA.n1489 257.466
R651 GNDA.n961 GNDA.n582 257.466
R652 GNDA.n1061 GNDA.n333 257.466
R653 GNDA.n260 GNDA.n258 257.466
R654 GNDA.n960 GNDA.n583 254.444
R655 GNDA.n1386 GNDA.n31 254.34
R656 GNDA.n1457 GNDA.n31 254.34
R657 GNDA.n1459 GNDA.n31 254.34
R658 GNDA.n1472 GNDA.n31 254.34
R659 GNDA.n1474 GNDA.n31 254.34
R660 GNDA.n1488 GNDA.n31 254.34
R661 GNDA.n883 GNDA.n758 254.34
R662 GNDA.n874 GNDA.n576 254.34
R663 GNDA.n762 GNDA.n576 254.34
R664 GNDA.n796 GNDA.n576 254.34
R665 GNDA.n798 GNDA.n576 254.34
R666 GNDA.n811 GNDA.n576 254.34
R667 GNDA.n813 GNDA.n576 254.34
R668 GNDA.n914 GNDA.n579 254.34
R669 GNDA.n913 GNDA.n579 254.34
R670 GNDA.n921 GNDA.n579 254.34
R671 GNDA.n910 GNDA.n579 254.34
R672 GNDA.n928 GNDA.n579 254.34
R673 GNDA.n907 GNDA.n579 254.34
R674 GNDA.n1523 GNDA.n35 254.34
R675 GNDA.n1520 GNDA.n35 254.34
R676 GNDA.n1508 GNDA.n35 254.34
R677 GNDA.n1506 GNDA.n35 254.34
R678 GNDA.n1496 GNDA.n35 254.34
R679 GNDA.n1494 GNDA.n35 254.34
R680 GNDA.n79 GNDA.n5 254.34
R681 GNDA.n1516 GNDA.n5 254.34
R682 GNDA.n1512 GNDA.n5 254.34
R683 GNDA.n1502 GNDA.n5 254.34
R684 GNDA.n1500 GNDA.n5 254.34
R685 GNDA.n1490 GNDA.n5 254.34
R686 GNDA.n746 GNDA.n601 254.34
R687 GNDA.n746 GNDA.n600 254.34
R688 GNDA.n746 GNDA.n599 254.34
R689 GNDA.n746 GNDA.n598 254.34
R690 GNDA.n746 GNDA.n597 254.34
R691 GNDA.n746 GNDA.n596 254.34
R692 GNDA.n1550 GNDA.n63 254.34
R693 GNDA.n1548 GNDA.n63 254.34
R694 GNDA.n1542 GNDA.n63 254.34
R695 GNDA.n1540 GNDA.n63 254.34
R696 GNDA.n1534 GNDA.n63 254.34
R697 GNDA.n1532 GNDA.n63 254.34
R698 GNDA.n727 GNDA.n726 254.34
R699 GNDA.n502 GNDA.n17 254.34
R700 GNDA.n466 GNDA.n17 254.34
R701 GNDA.n477 GNDA.n17 254.34
R702 GNDA.n479 GNDA.n17 254.34
R703 GNDA.n489 GNDA.n17 254.34
R704 GNDA.n491 GNDA.n17 254.34
R705 GNDA.n507 GNDA.n380 254.34
R706 GNDA.n278 GNDA.n277 254.34
R707 GNDA.n272 GNDA.n31 254.34
R708 GNDA.n233 GNDA.n31 254.34
R709 GNDA.n244 GNDA.n31 254.34
R710 GNDA.n246 GNDA.n31 254.34
R711 GNDA.n256 GNDA.n31 254.34
R712 GNDA.n261 GNDA.n31 254.34
R713 GNDA.n323 GNDA.n30 254.34
R714 GNDA.n321 GNDA.n30 254.34
R715 GNDA.n315 GNDA.n30 254.34
R716 GNDA.n313 GNDA.n30 254.34
R717 GNDA.n307 GNDA.n30 254.34
R718 GNDA.n305 GNDA.n30 254.34
R719 GNDA.n134 GNDA.n23 254.34
R720 GNDA.n128 GNDA.n23 254.34
R721 GNDA.n125 GNDA.n23 254.34
R722 GNDA.n119 GNDA.n23 254.34
R723 GNDA.n116 GNDA.n23 254.34
R724 GNDA.n1383 GNDA.n23 254.34
R725 GNDA.n1364 GNDA.n20 254.34
R726 GNDA.n131 GNDA.n20 254.34
R727 GNDA.n1371 GNDA.n20 254.34
R728 GNDA.n122 GNDA.n20 254.34
R729 GNDA.n1378 GNDA.n20 254.34
R730 GNDA.n114 GNDA.n20 254.34
R731 GNDA.n357 GNDA.n23 254.34
R732 GNDA.n351 GNDA.n23 254.34
R733 GNDA.n348 GNDA.n23 254.34
R734 GNDA.n342 GNDA.n23 254.34
R735 GNDA.n339 GNDA.n23 254.34
R736 GNDA.n336 GNDA.n23 254.34
R737 GNDA.n1043 GNDA.n20 254.34
R738 GNDA.n354 GNDA.n20 254.34
R739 GNDA.n1050 GNDA.n20 254.34
R740 GNDA.n345 GNDA.n20 254.34
R741 GNDA.n1057 GNDA.n20 254.34
R742 GNDA.n1060 GNDA.n20 254.34
R743 GNDA.n1213 GNDA.n64 254.34
R744 GNDA.n1176 GNDA.n64 254.34
R745 GNDA.n1187 GNDA.n64 254.34
R746 GNDA.n1189 GNDA.n64 254.34
R747 GNDA.n1199 GNDA.n64 254.34
R748 GNDA.n1202 GNDA.n64 254.34
R749 GNDA.n1561 GNDA.n1560 254.34
R750 GNDA.n35 GNDA.n34 254.34
R751 GNDA.n35 GNDA.n33 254.34
R752 GNDA.n1227 GNDA.n35 254.34
R753 GNDA.n1229 GNDA.n35 254.34
R754 GNDA.n1224 GNDA.n35 254.34
R755 GNDA.n1218 GNDA.n35 254.34
R756 GNDA.n11 GNDA.n5 254.34
R757 GNDA.n1614 GNDA.n5 254.34
R758 GNDA.n5 GNDA.n4 254.34
R759 GNDA.n1231 GNDA.n5 254.34
R760 GNDA.n1238 GNDA.n5 254.34
R761 GNDA.n1221 GNDA.n5 254.34
R762 GNDA.n1609 GNDA.n1608 251.614
R763 GNDA.n1580 GNDA.n49 251.614
R764 GNDA.n1555 GNDA.n67 251.614
R765 GNDA.n1527 GNDA.n1526 251.614
R766 GNDA.n941 GNDA.n594 251.614
R767 GNDA.n1042 GNDA.n355 251.614
R768 GNDA.n1363 GNDA.n132 251.614
R769 GNDA.n1011 GNDA.n27 250.349
R770 GNDA.n969 GNDA.n968 246.25
R771 GNDA.n996 GNDA.n968 246.25
R772 GNDA.n994 GNDA.n993 246.25
R773 GNDA.n988 GNDA.n967 246.25
R774 GNDA.n1007 GNDA.t18 245.133
R775 GNDA.n1003 GNDA.n1002 241.643
R776 GNDA.n1003 GNDA.n965 241.643
R777 GNDA.n1003 GNDA.n966 241.643
R778 GNDA.t24 GNDA.n962 214.2
R779 GNDA.n1013 GNDA.n1012 197
R780 GNDA.n331 GNDA.n329 195.049
R781 GNDA.n1217 GNDA.n1216 195.049
R782 GNDA.n1493 GNDA.n90 195.049
R783 GNDA.n1385 GNDA.n1384 195.049
R784 GNDA.n882 GNDA.n881 195.049
R785 GNDA.n504 GNDA.n385 195.049
R786 GNDA.n274 GNDA.n151 195.049
R787 GNDA.n573 GNDA.t29 192.167
R788 GNDA.n290 GNDA.t22 190.952
R789 GNDA.t22 GNDA.n374 190.952
R790 GNDA.n1039 GNDA.n358 187.249
R791 GNDA.n1605 GNDA.n9 187.249
R792 GNDA.n1524 GNDA.n74 187.249
R793 GNDA.n1360 GNDA.n135 187.249
R794 GNDA.n937 GNDA.n748 187.249
R795 GNDA.n526 GNDA.n369 187.249
R796 GNDA.n300 GNDA.n141 187.249
R797 GNDA.n573 GNDA.t31 185.257
R798 GNDA.n1156 GNDA.n1109 185
R799 GNDA.t28 GNDA.n1109 185
R800 GNDA.n1158 GNDA.n1157 185
R801 GNDA.n1160 GNDA.n1159 185
R802 GNDA.n1162 GNDA.n1161 185
R803 GNDA.n1164 GNDA.n1163 185
R804 GNDA.n1166 GNDA.n1165 185
R805 GNDA.n1168 GNDA.n1167 185
R806 GNDA.n1169 GNDA.n1114 185
R807 GNDA.t28 GNDA.n1114 185
R808 GNDA.n1170 GNDA.n1118 185
R809 GNDA.n1155 GNDA.n1154 185
R810 GNDA.n1153 GNDA.n1152 185
R811 GNDA.n1151 GNDA.n1150 185
R812 GNDA.n1149 GNDA.n1148 185
R813 GNDA.n1147 GNDA.n1146 185
R814 GNDA.n1145 GNDA.n1144 185
R815 GNDA.n1143 GNDA.n1142 185
R816 GNDA.n1141 GNDA.n1140 185
R817 GNDA.n1139 GNDA.n1138 185
R818 GNDA.n1137 GNDA.n1136 185
R819 GNDA.n1135 GNDA.n1134 185
R820 GNDA.n1133 GNDA.n1132 185
R821 GNDA.n1131 GNDA.n1130 185
R822 GNDA.n1129 GNDA.n1128 185
R823 GNDA.n1127 GNDA.n1126 185
R824 GNDA.n1125 GNDA.n1124 185
R825 GNDA.n1123 GNDA.n1122 185
R826 GNDA.n1121 GNDA.n1099 185
R827 GNDA.n1310 GNDA.n1084 185
R828 GNDA.n1084 GNDA.t33 185
R829 GNDA.n1309 GNDA.n1308 185
R830 GNDA.n1306 GNDA.n1085 185
R831 GNDA.n1305 GNDA.n1086 185
R832 GNDA.n1303 GNDA.n1302 185
R833 GNDA.n1301 GNDA.n1087 185
R834 GNDA.n1300 GNDA.n1299 185
R835 GNDA.n1297 GNDA.n1088 185
R836 GNDA.n1297 GNDA.t33 185
R837 GNDA.n1296 GNDA.n1089 185
R838 GNDA.n1312 GNDA.n1311 185
R839 GNDA.n1314 GNDA.n1082 185
R840 GNDA.n1316 GNDA.n1315 185
R841 GNDA.n1317 GNDA.n1081 185
R842 GNDA.n1319 GNDA.n1318 185
R843 GNDA.n1321 GNDA.n1079 185
R844 GNDA.n1323 GNDA.n1322 185
R845 GNDA.n1324 GNDA.n1078 185
R846 GNDA.n1326 GNDA.n1325 185
R847 GNDA.n1328 GNDA.n1077 185
R848 GNDA.n1330 GNDA.n1329 185
R849 GNDA.n1332 GNDA.n1331 185
R850 GNDA.n1335 GNDA.n1334 185
R851 GNDA.n1336 GNDA.n1075 185
R852 GNDA.n1338 GNDA.n1337 185
R853 GNDA.n1340 GNDA.n1074 185
R854 GNDA.n1342 GNDA.n1341 185
R855 GNDA.n1344 GNDA.n1343 185
R856 GNDA.n446 GNDA.n399 185
R857 GNDA.t32 GNDA.n399 185
R858 GNDA.n448 GNDA.n447 185
R859 GNDA.n450 GNDA.n449 185
R860 GNDA.n452 GNDA.n451 185
R861 GNDA.n454 GNDA.n453 185
R862 GNDA.n456 GNDA.n455 185
R863 GNDA.n458 GNDA.n457 185
R864 GNDA.n459 GNDA.n404 185
R865 GNDA.t32 GNDA.n404 185
R866 GNDA.n460 GNDA.n408 185
R867 GNDA.n445 GNDA.n444 185
R868 GNDA.n443 GNDA.n442 185
R869 GNDA.n441 GNDA.n440 185
R870 GNDA.n439 GNDA.n438 185
R871 GNDA.n437 GNDA.n436 185
R872 GNDA.n435 GNDA.n434 185
R873 GNDA.n433 GNDA.n432 185
R874 GNDA.n431 GNDA.n430 185
R875 GNDA.n429 GNDA.n428 185
R876 GNDA.n427 GNDA.n426 185
R877 GNDA.n425 GNDA.n424 185
R878 GNDA.n423 GNDA.n422 185
R879 GNDA.n421 GNDA.n420 185
R880 GNDA.n419 GNDA.n418 185
R881 GNDA.n417 GNDA.n416 185
R882 GNDA.n415 GNDA.n414 185
R883 GNDA.n413 GNDA.n412 185
R884 GNDA.n411 GNDA.n389 185
R885 GNDA.n654 GNDA.n634 185
R886 GNDA.n634 GNDA.t26 185
R887 GNDA.n653 GNDA.n652 185
R888 GNDA.n650 GNDA.n635 185
R889 GNDA.n649 GNDA.n636 185
R890 GNDA.n647 GNDA.n646 185
R891 GNDA.n645 GNDA.n637 185
R892 GNDA.n644 GNDA.n643 185
R893 GNDA.n641 GNDA.n638 185
R894 GNDA.n641 GNDA.t26 185
R895 GNDA.n640 GNDA.n610 185
R896 GNDA.n656 GNDA.n655 185
R897 GNDA.n658 GNDA.n632 185
R898 GNDA.n660 GNDA.n659 185
R899 GNDA.n661 GNDA.n631 185
R900 GNDA.n663 GNDA.n662 185
R901 GNDA.n665 GNDA.n629 185
R902 GNDA.n667 GNDA.n666 185
R903 GNDA.n668 GNDA.n628 185
R904 GNDA.n670 GNDA.n669 185
R905 GNDA.n672 GNDA.n627 185
R906 GNDA.n675 GNDA.n674 185
R907 GNDA.n676 GNDA.n626 185
R908 GNDA.n678 GNDA.n677 185
R909 GNDA.n680 GNDA.n625 185
R910 GNDA.n682 GNDA.n681 185
R911 GNDA.n684 GNDA.n683 185
R912 GNDA.n685 GNDA.n621 185
R913 GNDA.n688 GNDA.n687 185
R914 GNDA.n1416 GNDA.n1400 185
R915 GNDA.n1400 GNDA.t21 185
R916 GNDA.n1415 GNDA.n1414 185
R917 GNDA.n1412 GNDA.n1401 185
R918 GNDA.n1411 GNDA.n1402 185
R919 GNDA.n1409 GNDA.n1408 185
R920 GNDA.n1407 GNDA.n1403 185
R921 GNDA.n1406 GNDA.n1405 185
R922 GNDA.n96 GNDA.n95 185
R923 GNDA.t21 GNDA.n96 185
R924 GNDA.n1484 GNDA.n1483 185
R925 GNDA.n1418 GNDA.n1417 185
R926 GNDA.n1420 GNDA.n1398 185
R927 GNDA.n1422 GNDA.n1421 185
R928 GNDA.n1423 GNDA.n1397 185
R929 GNDA.n1425 GNDA.n1424 185
R930 GNDA.n1427 GNDA.n1395 185
R931 GNDA.n1429 GNDA.n1428 185
R932 GNDA.n1430 GNDA.n1394 185
R933 GNDA.n1432 GNDA.n1431 185
R934 GNDA.n1434 GNDA.n1393 185
R935 GNDA.n1436 GNDA.n1435 185
R936 GNDA.n1438 GNDA.n1437 185
R937 GNDA.n1441 GNDA.n1440 185
R938 GNDA.n1442 GNDA.n1391 185
R939 GNDA.n1444 GNDA.n1443 185
R940 GNDA.n1446 GNDA.n1390 185
R941 GNDA.n1448 GNDA.n1447 185
R942 GNDA.n1450 GNDA.n1449 185
R943 GNDA.n1453 GNDA.n1452 185
R944 GNDA.n1454 GNDA.n104 185
R945 GNDA.n1463 GNDA.n1462 185
R946 GNDA.n1465 GNDA.n103 185
R947 GNDA.n1468 GNDA.n1467 185
R948 GNDA.n1469 GNDA.n99 185
R949 GNDA.n1478 GNDA.n1477 185
R950 GNDA.n1480 GNDA.n98 185
R951 GNDA.n1481 GNDA.n94 185
R952 GNDA.n999 GNDA.n998 185
R953 GNDA.n997 GNDA.n972 185
R954 GNDA.n995 GNDA.n992 185
R955 GNDA.n991 GNDA.n976 185
R956 GNDA.n971 GNDA.n970 185
R957 GNDA.n998 GNDA.n973 185
R958 GNDA.n997 GNDA.n974 185
R959 GNDA.n995 GNDA.n975 185
R960 GNDA.n986 GNDA.n976 185
R961 GNDA.n989 GNDA.n987 185
R962 GNDA.n833 GNDA.n775 185
R963 GNDA.n775 GNDA.t23 185
R964 GNDA.n832 GNDA.n831 185
R965 GNDA.n829 GNDA.n776 185
R966 GNDA.n828 GNDA.n777 185
R967 GNDA.n826 GNDA.n825 185
R968 GNDA.n824 GNDA.n778 185
R969 GNDA.n823 GNDA.n822 185
R970 GNDA.n820 GNDA.n779 185
R971 GNDA.n820 GNDA.t23 185
R972 GNDA.n819 GNDA.n780 185
R973 GNDA.n835 GNDA.n834 185
R974 GNDA.n837 GNDA.n773 185
R975 GNDA.n839 GNDA.n838 185
R976 GNDA.n840 GNDA.n772 185
R977 GNDA.n842 GNDA.n841 185
R978 GNDA.n844 GNDA.n770 185
R979 GNDA.n846 GNDA.n845 185
R980 GNDA.n847 GNDA.n769 185
R981 GNDA.n849 GNDA.n848 185
R982 GNDA.n851 GNDA.n768 185
R983 GNDA.n854 GNDA.n853 185
R984 GNDA.n855 GNDA.n767 185
R985 GNDA.n857 GNDA.n856 185
R986 GNDA.n859 GNDA.n766 185
R987 GNDA.n862 GNDA.n861 185
R988 GNDA.n863 GNDA.n765 185
R989 GNDA.n865 GNDA.n864 185
R990 GNDA.n867 GNDA.n760 185
R991 GNDA.n868 GNDA.n761 185
R992 GNDA.n871 GNDA.n870 185
R993 GNDA.n792 GNDA.n764 185
R994 GNDA.n793 GNDA.n789 185
R995 GNDA.n802 GNDA.n801 185
R996 GNDA.n804 GNDA.n787 185
R997 GNDA.n807 GNDA.n806 185
R998 GNDA.n808 GNDA.n781 185
R999 GNDA.n817 GNDA.n816 185
R1000 GNDA.n623 GNDA.n620 185
R1001 GNDA.n696 GNDA.n619 185
R1002 GNDA.n701 GNDA.n700 185
R1003 GNDA.n704 GNDA.n703 185
R1004 GNDA.n618 GNDA.n615 185
R1005 GNDA.n709 GNDA.n614 185
R1006 GNDA.n714 GNDA.n713 185
R1007 GNDA.n717 GNDA.n716 185
R1008 GNDA.n613 GNDA.n611 185
R1009 GNDA.n499 GNDA.n498 185
R1010 GNDA.n468 GNDA.n390 185
R1011 GNDA.n471 GNDA.n470 185
R1012 GNDA.n474 GNDA.n473 185
R1013 GNDA.n472 GNDA.n464 185
R1014 GNDA.n483 GNDA.n482 185
R1015 GNDA.n485 GNDA.n484 185
R1016 GNDA.n486 GNDA.n409 185
R1017 GNDA.n495 GNDA.n494 185
R1018 GNDA.n213 GNDA.n166 185
R1019 GNDA.t25 GNDA.n166 185
R1020 GNDA.n215 GNDA.n214 185
R1021 GNDA.n217 GNDA.n216 185
R1022 GNDA.n219 GNDA.n218 185
R1023 GNDA.n221 GNDA.n220 185
R1024 GNDA.n223 GNDA.n222 185
R1025 GNDA.n225 GNDA.n224 185
R1026 GNDA.n226 GNDA.n171 185
R1027 GNDA.t25 GNDA.n171 185
R1028 GNDA.n227 GNDA.n175 185
R1029 GNDA.n212 GNDA.n211 185
R1030 GNDA.n210 GNDA.n209 185
R1031 GNDA.n208 GNDA.n207 185
R1032 GNDA.n206 GNDA.n205 185
R1033 GNDA.n204 GNDA.n203 185
R1034 GNDA.n202 GNDA.n201 185
R1035 GNDA.n200 GNDA.n199 185
R1036 GNDA.n198 GNDA.n197 185
R1037 GNDA.n196 GNDA.n195 185
R1038 GNDA.n194 GNDA.n193 185
R1039 GNDA.n192 GNDA.n191 185
R1040 GNDA.n190 GNDA.n189 185
R1041 GNDA.n188 GNDA.n187 185
R1042 GNDA.n186 GNDA.n185 185
R1043 GNDA.n184 GNDA.n183 185
R1044 GNDA.n182 GNDA.n181 185
R1045 GNDA.n180 GNDA.n179 185
R1046 GNDA.n178 GNDA.n156 185
R1047 GNDA.n269 GNDA.n268 185
R1048 GNDA.n235 GNDA.n157 185
R1049 GNDA.n238 GNDA.n237 185
R1050 GNDA.n241 GNDA.n240 185
R1051 GNDA.n239 GNDA.n231 185
R1052 GNDA.n250 GNDA.n249 185
R1053 GNDA.n252 GNDA.n251 185
R1054 GNDA.n253 GNDA.n176 185
R1055 GNDA.n265 GNDA.n264 185
R1056 GNDA.n1345 GNDA.n1070 185
R1057 GNDA.n1348 GNDA.n1347 185
R1058 GNDA.n1258 GNDA.n1072 185
R1059 GNDA.n1257 GNDA.n1256 185
R1060 GNDA.n1275 GNDA.n1274 185
R1061 GNDA.n1277 GNDA.n1252 185
R1062 GNDA.n1280 GNDA.n1279 185
R1063 GNDA.n1253 GNDA.n1090 185
R1064 GNDA.n1294 GNDA.n1293 185
R1065 GNDA.n1210 GNDA.n1209 185
R1066 GNDA.n1178 GNDA.n1100 185
R1067 GNDA.n1181 GNDA.n1180 185
R1068 GNDA.n1184 GNDA.n1183 185
R1069 GNDA.n1182 GNDA.n1174 185
R1070 GNDA.n1193 GNDA.n1192 185
R1071 GNDA.n1195 GNDA.n1194 185
R1072 GNDA.n1196 GNDA.n1119 185
R1073 GNDA.n1206 GNDA.n1205 185
R1074 GNDA.n1038 GNDA.n553 175.546
R1075 GNDA.n1034 GNDA.n553 175.546
R1076 GNDA.n1034 GNDA.n556 175.546
R1077 GNDA.n1030 GNDA.n556 175.546
R1078 GNDA.n1030 GNDA.n1027 175.546
R1079 GNDA.n1027 GNDA.n1026 175.546
R1080 GNDA.n1026 GNDA.n559 175.546
R1081 GNDA.n1022 GNDA.n559 175.546
R1082 GNDA.n1022 GNDA.n1018 175.546
R1083 GNDA.n1018 GNDA.n12 175.546
R1084 GNDA.n1608 GNDA.n12 175.546
R1085 GNDA.n1240 GNDA.n1239 175.546
R1086 GNDA.n1237 GNDA.n1222 175.546
R1087 GNDA.n1233 GNDA.n1232 175.546
R1088 GNDA.n1616 GNDA.n1615 175.546
R1089 GNDA.n1613 GNDA.n6 175.546
R1090 GNDA.n1354 GNDA.n1064 175.546
R1091 GNDA.n1350 GNDA.n1064 175.546
R1092 GNDA.n1350 GNDA.n1068 175.546
R1093 GNDA.n1270 GNDA.n1068 175.546
R1094 GNDA.n1271 GNDA.n1270 175.546
R1095 GNDA.n1271 GNDA.n1250 175.546
R1096 GNDA.n1282 GNDA.n1250 175.546
R1097 GNDA.n1282 GNDA.n1251 175.546
R1098 GNDA.n1251 GNDA.n1093 175.546
R1099 GNDA.n1291 GNDA.n1093 175.546
R1100 GNDA.n1291 GNDA.n1245 175.546
R1101 GNDA.n338 GNDA.n337 175.546
R1102 GNDA.n341 GNDA.n340 175.546
R1103 GNDA.n347 GNDA.n343 175.546
R1104 GNDA.n350 GNDA.n349 175.546
R1105 GNDA.n356 GNDA.n352 175.546
R1106 GNDA.n1212 GNDA.n1096 175.546
R1107 GNDA.n1186 GNDA.n1177 175.546
R1108 GNDA.n1190 GNDA.n1188 175.546
R1109 GNDA.n1198 GNDA.n1172 175.546
R1110 GNDA.n1203 GNDA.n1200 175.546
R1111 GNDA.n1223 GNDA.n1219 175.546
R1112 GNDA.n1226 GNDA.n1225 175.546
R1113 GNDA.n1230 GNDA.n1228 175.546
R1114 GNDA.n32 GNDA.n2 175.546
R1115 GNDA.n8 GNDA.n7 175.546
R1116 GNDA.n1604 GNDA.n37 175.546
R1117 GNDA.n1600 GNDA.n37 175.546
R1118 GNDA.n1600 GNDA.n40 175.546
R1119 GNDA.n1596 GNDA.n40 175.546
R1120 GNDA.n1596 GNDA.n43 175.546
R1121 GNDA.n1592 GNDA.n43 175.546
R1122 GNDA.n1592 GNDA.n45 175.546
R1123 GNDA.n1588 GNDA.n45 175.546
R1124 GNDA.n1588 GNDA.n47 175.546
R1125 GNDA.n1584 GNDA.n47 175.546
R1126 GNDA.n1584 GNDA.n49 175.546
R1127 GNDA.n1559 GNDA.n59 175.546
R1128 GNDA.n1564 GNDA.n59 175.546
R1129 GNDA.n1564 GNDA.n57 175.546
R1130 GNDA.n1568 GNDA.n57 175.546
R1131 GNDA.n1568 GNDA.n55 175.546
R1132 GNDA.n1572 GNDA.n55 175.546
R1133 GNDA.n1572 GNDA.n53 175.546
R1134 GNDA.n1576 GNDA.n53 175.546
R1135 GNDA.n1576 GNDA.n51 175.546
R1136 GNDA.n1580 GNDA.n51 175.546
R1137 GNDA.n1535 GNDA.n1533 175.546
R1138 GNDA.n1539 GNDA.n72 175.546
R1139 GNDA.n1543 GNDA.n1541 175.546
R1140 GNDA.n1547 GNDA.n70 175.546
R1141 GNDA.n1551 GNDA.n1549 175.546
R1142 GNDA.n729 GNDA.n609 175.546
R1143 GNDA.n729 GNDA.n607 175.546
R1144 GNDA.n733 GNDA.n607 175.546
R1145 GNDA.n733 GNDA.n604 175.546
R1146 GNDA.n744 GNDA.n604 175.546
R1147 GNDA.n744 GNDA.n605 175.546
R1148 GNDA.n740 GNDA.n605 175.546
R1149 GNDA.n740 GNDA.n737 175.546
R1150 GNDA.n737 GNDA.n66 175.546
R1151 GNDA.n1555 GNDA.n66 175.546
R1152 GNDA.n694 GNDA.n693 175.546
R1153 GNDA.n698 GNDA.n697 175.546
R1154 GNDA.n707 GNDA.n706 175.546
R1155 GNDA.n711 GNDA.n710 175.546
R1156 GNDA.n720 GNDA.n719 175.546
R1157 GNDA.n1497 GNDA.n1495 175.546
R1158 GNDA.n1505 GNDA.n86 175.546
R1159 GNDA.n1509 GNDA.n1507 175.546
R1160 GNDA.n1519 GNDA.n82 175.546
R1161 GNDA.n1522 GNDA.n1521 175.546
R1162 GNDA.n1382 GNDA.n112 175.546
R1163 GNDA.n118 GNDA.n117 175.546
R1164 GNDA.n124 GNDA.n120 175.546
R1165 GNDA.n127 GNDA.n126 175.546
R1166 GNDA.n133 GNDA.n129 175.546
R1167 GNDA.n1065 GNDA.n328 175.546
R1168 GNDA.n1066 GNDA.n1065 175.546
R1169 GNDA.n1260 GNDA.n1066 175.546
R1170 GNDA.n1268 GNDA.n1260 175.546
R1171 GNDA.n1268 GNDA.n1261 175.546
R1172 GNDA.n1261 GNDA.n1249 175.546
R1173 GNDA.n1284 GNDA.n1249 175.546
R1174 GNDA.n1284 GNDA.n1247 175.546
R1175 GNDA.n1288 GNDA.n1247 175.546
R1176 GNDA.n1288 GNDA.n78 175.546
R1177 GNDA.n1527 GNDA.n78 175.546
R1178 GNDA.n1499 GNDA.n88 175.546
R1179 GNDA.n1503 GNDA.n1501 175.546
R1180 GNDA.n1511 GNDA.n84 175.546
R1181 GNDA.n1517 GNDA.n1513 175.546
R1182 GNDA.n1515 GNDA.n1514 175.546
R1183 GNDA.n1456 GNDA.n106 175.546
R1184 GNDA.n1460 GNDA.n1458 175.546
R1185 GNDA.n1471 GNDA.n101 175.546
R1186 GNDA.n1475 GNDA.n1473 175.546
R1187 GNDA.n1487 GNDA.n93 175.546
R1188 GNDA.n930 GNDA.n929 175.546
R1189 GNDA.n927 GNDA.n908 175.546
R1190 GNDA.n923 GNDA.n922 175.546
R1191 GNDA.n920 GNDA.n911 175.546
R1192 GNDA.n916 GNDA.n915 175.546
R1193 GNDA.n959 GNDA.n958 175.546
R1194 GNDA.n958 GNDA.n584 175.546
R1195 GNDA.n954 GNDA.n584 175.546
R1196 GNDA.n954 GNDA.n586 175.546
R1197 GNDA.n950 GNDA.n586 175.546
R1198 GNDA.n950 GNDA.n949 175.546
R1199 GNDA.n949 GNDA.n589 175.546
R1200 GNDA.n945 GNDA.n589 175.546
R1201 GNDA.n945 GNDA.n591 175.546
R1202 GNDA.n941 GNDA.n591 175.546
R1203 GNDA.n875 GNDA.n873 175.546
R1204 GNDA.n795 GNDA.n791 175.546
R1205 GNDA.n799 GNDA.n797 175.546
R1206 GNDA.n810 GNDA.n785 175.546
R1207 GNDA.n814 GNDA.n812 175.546
R1208 GNDA.n887 GNDA.n884 175.546
R1209 GNDA.n887 GNDA.n757 175.546
R1210 GNDA.n891 GNDA.n757 175.546
R1211 GNDA.n891 GNDA.n755 175.546
R1212 GNDA.n895 GNDA.n755 175.546
R1213 GNDA.n895 GNDA.n753 175.546
R1214 GNDA.n899 GNDA.n753 175.546
R1215 GNDA.n899 GNDA.n751 175.546
R1216 GNDA.n903 GNDA.n751 175.546
R1217 GNDA.n903 GNDA.n748 175.546
R1218 GNDA.n382 GNDA.n379 175.546
R1219 GNDA.n510 GNDA.n379 175.546
R1220 GNDA.n510 GNDA.n377 175.546
R1221 GNDA.n514 GNDA.n377 175.546
R1222 GNDA.n514 GNDA.n375 175.546
R1223 GNDA.n518 GNDA.n375 175.546
R1224 GNDA.n518 GNDA.n373 175.546
R1225 GNDA.n522 GNDA.n373 175.546
R1226 GNDA.n522 GNDA.n371 175.546
R1227 GNDA.n526 GNDA.n371 175.546
R1228 GNDA.n501 GNDA.n386 175.546
R1229 GNDA.n476 GNDA.n467 175.546
R1230 GNDA.n480 GNDA.n478 175.546
R1231 GNDA.n488 GNDA.n462 175.546
R1232 GNDA.n492 GNDA.n490 175.546
R1233 GNDA.n1059 GNDA.n1058 175.546
R1234 GNDA.n1056 GNDA.n335 175.546
R1235 GNDA.n1052 GNDA.n1051 175.546
R1236 GNDA.n1049 GNDA.n346 175.546
R1237 GNDA.n1045 GNDA.n1044 175.546
R1238 GNDA.n530 GNDA.n367 175.546
R1239 GNDA.n535 GNDA.n367 175.546
R1240 GNDA.n535 GNDA.n364 175.546
R1241 GNDA.n539 GNDA.n364 175.546
R1242 GNDA.n540 GNDA.n539 175.546
R1243 GNDA.n541 GNDA.n540 175.546
R1244 GNDA.n541 GNDA.n362 175.546
R1245 GNDA.n545 GNDA.n362 175.546
R1246 GNDA.n545 GNDA.n360 175.546
R1247 GNDA.n549 GNDA.n360 175.546
R1248 GNDA.n549 GNDA.n355 175.546
R1249 GNDA.n308 GNDA.n306 175.546
R1250 GNDA.n312 GNDA.n139 175.546
R1251 GNDA.n316 GNDA.n314 175.546
R1252 GNDA.n320 GNDA.n137 175.546
R1253 GNDA.n324 GNDA.n322 175.546
R1254 GNDA.n1380 GNDA.n1379 175.546
R1255 GNDA.n1377 GNDA.n115 175.546
R1256 GNDA.n1373 GNDA.n1372 175.546
R1257 GNDA.n1370 GNDA.n123 175.546
R1258 GNDA.n1366 GNDA.n1365 175.546
R1259 GNDA.n271 GNDA.n153 175.546
R1260 GNDA.n243 GNDA.n234 175.546
R1261 GNDA.n247 GNDA.n245 175.546
R1262 GNDA.n255 GNDA.n229 175.546
R1263 GNDA.n262 GNDA.n257 175.546
R1264 GNDA.n279 GNDA.n150 175.546
R1265 GNDA.n283 GNDA.n150 175.546
R1266 GNDA.n283 GNDA.n148 175.546
R1267 GNDA.n288 GNDA.n148 175.546
R1268 GNDA.n288 GNDA.n146 175.546
R1269 GNDA.n292 GNDA.n146 175.546
R1270 GNDA.n292 GNDA.n145 175.546
R1271 GNDA.n296 GNDA.n145 175.546
R1272 GNDA.n296 GNDA.n143 175.546
R1273 GNDA.n300 GNDA.n143 175.546
R1274 GNDA.t22 GNDA.n289 174.701
R1275 GNDA.n513 GNDA.t22 174.701
R1276 GNDA.t22 GNDA.n17 172.876
R1277 GNDA.t22 GNDA.n30 172.615
R1278 GNDA.n1209 GNDA.n1099 163.333
R1279 GNDA.n1345 GNDA.n1344 163.333
R1280 GNDA.n498 GNDA.n389 163.333
R1281 GNDA.n687 GNDA.n623 163.333
R1282 GNDA.n1452 GNDA.n1450 163.333
R1283 GNDA.n868 GNDA.n867 163.333
R1284 GNDA.n268 GNDA.n156 163.333
R1285 GNDA.t22 GNDA.n19 162.964
R1286 GNDA.t27 GNDA.n42 162.964
R1287 GNDA.n0 GNDA.n23 22.8229
R1288 GNDA.t22 GNDA.n35 161.738
R1289 GNDA.n567 GNDA.t9 160.534
R1290 GNDA.n566 GNDA.t34 159.927
R1291 GNDA.n939 GNDA.n938 158.506
R1292 GNDA.n939 GNDA.n31 157.35
R1293 GNDA.t10 GNDA.n1003 151.725
R1294 GNDA.n565 GNDA.t17 150.327
R1295 GNDA.n1180 GNDA.n1100 150
R1296 GNDA.n1183 GNDA.n1182 150
R1297 GNDA.n1194 GNDA.n1193 150
R1298 GNDA.n1206 GNDA.n1119 150
R1299 GNDA.n1124 GNDA.n1123 150
R1300 GNDA.n1128 GNDA.n1127 150
R1301 GNDA.n1132 GNDA.n1131 150
R1302 GNDA.n1136 GNDA.n1135 150
R1303 GNDA.n1140 GNDA.n1139 150
R1304 GNDA.n1144 GNDA.n1143 150
R1305 GNDA.n1148 GNDA.n1147 150
R1306 GNDA.n1152 GNDA.n1151 150
R1307 GNDA.n1118 GNDA.n1114 150
R1308 GNDA.n1167 GNDA.n1114 150
R1309 GNDA.n1165 GNDA.n1164 150
R1310 GNDA.n1161 GNDA.n1160 150
R1311 GNDA.n1157 GNDA.n1109 150
R1312 GNDA.n1347 GNDA.n1072 150
R1313 GNDA.n1275 GNDA.n1256 150
R1314 GNDA.n1279 GNDA.n1277 150
R1315 GNDA.n1294 GNDA.n1090 150
R1316 GNDA.n1341 GNDA.n1340 150
R1317 GNDA.n1338 GNDA.n1075 150
R1318 GNDA.n1334 GNDA.n1332 150
R1319 GNDA.n1329 GNDA.n1328 150
R1320 GNDA.n1326 GNDA.n1078 150
R1321 GNDA.n1322 GNDA.n1321 150
R1322 GNDA.n1319 GNDA.n1081 150
R1323 GNDA.n1315 GNDA.n1314 150
R1324 GNDA.n1297 GNDA.n1296 150
R1325 GNDA.n1299 GNDA.n1297 150
R1326 GNDA.n1303 GNDA.n1087 150
R1327 GNDA.n1306 GNDA.n1305 150
R1328 GNDA.n1308 GNDA.n1084 150
R1329 GNDA.n470 GNDA.n390 150
R1330 GNDA.n473 GNDA.n472 150
R1331 GNDA.n484 GNDA.n483 150
R1332 GNDA.n495 GNDA.n409 150
R1333 GNDA.n414 GNDA.n413 150
R1334 GNDA.n418 GNDA.n417 150
R1335 GNDA.n422 GNDA.n421 150
R1336 GNDA.n426 GNDA.n425 150
R1337 GNDA.n430 GNDA.n429 150
R1338 GNDA.n434 GNDA.n433 150
R1339 GNDA.n438 GNDA.n437 150
R1340 GNDA.n442 GNDA.n441 150
R1341 GNDA.n408 GNDA.n404 150
R1342 GNDA.n457 GNDA.n404 150
R1343 GNDA.n455 GNDA.n454 150
R1344 GNDA.n451 GNDA.n450 150
R1345 GNDA.n447 GNDA.n399 150
R1346 GNDA.n701 GNDA.n619 150
R1347 GNDA.n703 GNDA.n618 150
R1348 GNDA.n714 GNDA.n614 150
R1349 GNDA.n716 GNDA.n613 150
R1350 GNDA.n685 GNDA.n684 150
R1351 GNDA.n681 GNDA.n680 150
R1352 GNDA.n678 GNDA.n626 150
R1353 GNDA.n674 GNDA.n672 150
R1354 GNDA.n670 GNDA.n628 150
R1355 GNDA.n666 GNDA.n665 150
R1356 GNDA.n663 GNDA.n631 150
R1357 GNDA.n659 GNDA.n658 150
R1358 GNDA.n641 GNDA.n640 150
R1359 GNDA.n643 GNDA.n641 150
R1360 GNDA.n647 GNDA.n637 150
R1361 GNDA.n650 GNDA.n649 150
R1362 GNDA.n652 GNDA.n634 150
R1363 GNDA.n1463 GNDA.n104 150
R1364 GNDA.n1467 GNDA.n1465 150
R1365 GNDA.n1478 GNDA.n99 150
R1366 GNDA.n1481 GNDA.n1480 150
R1367 GNDA.n1447 GNDA.n1446 150
R1368 GNDA.n1444 GNDA.n1391 150
R1369 GNDA.n1440 GNDA.n1438 150
R1370 GNDA.n1435 GNDA.n1434 150
R1371 GNDA.n1432 GNDA.n1394 150
R1372 GNDA.n1428 GNDA.n1427 150
R1373 GNDA.n1425 GNDA.n1397 150
R1374 GNDA.n1421 GNDA.n1420 150
R1375 GNDA.n1483 GNDA.n96 150
R1376 GNDA.n1405 GNDA.n96 150
R1377 GNDA.n1409 GNDA.n1403 150
R1378 GNDA.n1412 GNDA.n1411 150
R1379 GNDA.n1414 GNDA.n1400 150
R1380 GNDA.n973 GNDA.n970 150
R1381 GNDA.n974 GNDA.n973 150
R1382 GNDA.n986 GNDA.n975 150
R1383 GNDA.n987 GNDA.n986 150
R1384 GNDA.n999 GNDA.n972 150
R1385 GNDA.n992 GNDA.n991 150
R1386 GNDA.n870 GNDA.n764 150
R1387 GNDA.n802 GNDA.n789 150
R1388 GNDA.n806 GNDA.n804 150
R1389 GNDA.n817 GNDA.n781 150
R1390 GNDA.n865 GNDA.n765 150
R1391 GNDA.n861 GNDA.n859 150
R1392 GNDA.n857 GNDA.n767 150
R1393 GNDA.n853 GNDA.n851 150
R1394 GNDA.n849 GNDA.n769 150
R1395 GNDA.n845 GNDA.n844 150
R1396 GNDA.n842 GNDA.n772 150
R1397 GNDA.n838 GNDA.n837 150
R1398 GNDA.n820 GNDA.n819 150
R1399 GNDA.n822 GNDA.n820 150
R1400 GNDA.n826 GNDA.n778 150
R1401 GNDA.n829 GNDA.n828 150
R1402 GNDA.n831 GNDA.n775 150
R1403 GNDA.n237 GNDA.n157 150
R1404 GNDA.n240 GNDA.n239 150
R1405 GNDA.n251 GNDA.n250 150
R1406 GNDA.n265 GNDA.n176 150
R1407 GNDA.n181 GNDA.n180 150
R1408 GNDA.n185 GNDA.n184 150
R1409 GNDA.n189 GNDA.n188 150
R1410 GNDA.n193 GNDA.n192 150
R1411 GNDA.n197 GNDA.n196 150
R1412 GNDA.n201 GNDA.n200 150
R1413 GNDA.n205 GNDA.n204 150
R1414 GNDA.n209 GNDA.n208 150
R1415 GNDA.n175 GNDA.n171 150
R1416 GNDA.n224 GNDA.n171 150
R1417 GNDA.n222 GNDA.n221 150
R1418 GNDA.n218 GNDA.n217 150
R1419 GNDA.n214 GNDA.n166 150
R1420 GNDA.n1005 GNDA.t2 135.69
R1421 GNDA.n1007 GNDA.t20 130
R1422 GNDA.n1039 GNDA.n1038 126.782
R1423 GNDA.n1605 GNDA.n1604 126.782
R1424 GNDA.n1531 GNDA.n74 126.782
R1425 GNDA.n1360 GNDA.n328 126.782
R1426 GNDA.n937 GNDA.n749 126.782
R1427 GNDA.n530 GNDA.n369 126.782
R1428 GNDA.n304 GNDA.n141 126.782
R1429 GNDA.n1354 GNDA.n329 124.832
R1430 GNDA.n1216 GNDA.n1214 124.832
R1431 GNDA.n689 GNDA.n90 124.832
R1432 GNDA.n1387 GNDA.n1385 124.832
R1433 GNDA.n881 GNDA.n759 124.832
R1434 GNDA.n504 GNDA.n503 124.832
R1435 GNDA.n274 GNDA.n273 124.832
R1436 GNDA.t1 GNDA.t12 121.379
R1437 GNDA.t22 GNDA.n27 112.388
R1438 GNDA.n938 GNDA.n747 111.07
R1439 GNDA.n886 GNDA.n885 104.129
R1440 GNDA.n886 GNDA.n756 104.129
R1441 GNDA.n892 GNDA.n756 104.129
R1442 GNDA.n893 GNDA.n892 104.129
R1443 GNDA.n894 GNDA.n752 104.129
R1444 GNDA.n900 GNDA.n752 104.129
R1445 GNDA.n901 GNDA.n900 104.129
R1446 GNDA.n902 GNDA.n901 104.129
R1447 GNDA.n902 GNDA.n747 104.129
R1448 GNDA.n996 GNDA.n965 101.718
R1449 GNDA.n993 GNDA.n966 101.718
R1450 GNDA.n1002 GNDA.n969 101.718
R1451 GNDA.n994 GNDA.n965 101.718
R1452 GNDA.n988 GNDA.n966 101.718
R1453 GNDA.t22 GNDA.n29 97.5074
R1454 GNDA.n0 GNDA.t22 51.5983
R1455 GNDA.t27 GNDA.n62 95.5728
R1456 GNDA.t22 GNDA.n31 89.0881
R1457 GNDA.n1012 GNDA.n1011 84.306
R1458 GNDA.t22 GNDA.n26 80.9821
R1459 GNDA.n1240 GNDA.n1221 76.3222
R1460 GNDA.n1238 GNDA.n1237 76.3222
R1461 GNDA.n1233 GNDA.n1231 76.3222
R1462 GNDA.n1616 GNDA.n4 76.3222
R1463 GNDA.n1614 GNDA.n1613 76.3222
R1464 GNDA.n1609 GNDA.n11 76.3222
R1465 GNDA.n337 GNDA.n336 76.3222
R1466 GNDA.n340 GNDA.n339 76.3222
R1467 GNDA.n343 GNDA.n342 76.3222
R1468 GNDA.n349 GNDA.n348 76.3222
R1469 GNDA.n352 GNDA.n351 76.3222
R1470 GNDA.n358 GNDA.n357 76.3222
R1471 GNDA.n1214 GNDA.n1213 76.3222
R1472 GNDA.n1176 GNDA.n1096 76.3222
R1473 GNDA.n1187 GNDA.n1186 76.3222
R1474 GNDA.n1190 GNDA.n1189 76.3222
R1475 GNDA.n1199 GNDA.n1198 76.3222
R1476 GNDA.n1203 GNDA.n1202 76.3222
R1477 GNDA.n1218 GNDA.n1217 76.3222
R1478 GNDA.n1224 GNDA.n1223 76.3222
R1479 GNDA.n1229 GNDA.n1226 76.3222
R1480 GNDA.n1228 GNDA.n1227 76.3222
R1481 GNDA.n33 GNDA.n32 76.3222
R1482 GNDA.n34 GNDA.n9 76.3222
R1483 GNDA.n1560 GNDA.n1559 76.3222
R1484 GNDA.n1533 GNDA.n1532 76.3222
R1485 GNDA.n1534 GNDA.n72 76.3222
R1486 GNDA.n1541 GNDA.n1540 76.3222
R1487 GNDA.n1542 GNDA.n70 76.3222
R1488 GNDA.n1549 GNDA.n1548 76.3222
R1489 GNDA.n1550 GNDA.n67 76.3222
R1490 GNDA.n726 GNDA.n725 76.3222
R1491 GNDA.n689 GNDA.n601 76.3222
R1492 GNDA.n694 GNDA.n600 76.3222
R1493 GNDA.n697 GNDA.n599 76.3222
R1494 GNDA.n707 GNDA.n598 76.3222
R1495 GNDA.n710 GNDA.n597 76.3222
R1496 GNDA.n720 GNDA.n596 76.3222
R1497 GNDA.n1494 GNDA.n1493 76.3222
R1498 GNDA.n1497 GNDA.n1496 76.3222
R1499 GNDA.n1506 GNDA.n1505 76.3222
R1500 GNDA.n1509 GNDA.n1508 76.3222
R1501 GNDA.n1520 GNDA.n1519 76.3222
R1502 GNDA.n1523 GNDA.n1522 76.3222
R1503 GNDA.n1383 GNDA.n1382 76.3222
R1504 GNDA.n117 GNDA.n116 76.3222
R1505 GNDA.n120 GNDA.n119 76.3222
R1506 GNDA.n126 GNDA.n125 76.3222
R1507 GNDA.n129 GNDA.n128 76.3222
R1508 GNDA.n135 GNDA.n134 76.3222
R1509 GNDA.n1490 GNDA.n88 76.3222
R1510 GNDA.n1501 GNDA.n1500 76.3222
R1511 GNDA.n1502 GNDA.n84 76.3222
R1512 GNDA.n1513 GNDA.n1512 76.3222
R1513 GNDA.n1516 GNDA.n1515 76.3222
R1514 GNDA.n1526 GNDA.n79 76.3222
R1515 GNDA.n1387 GNDA.n1386 76.3222
R1516 GNDA.n1457 GNDA.n1456 76.3222
R1517 GNDA.n1460 GNDA.n1459 76.3222
R1518 GNDA.n1472 GNDA.n1471 76.3222
R1519 GNDA.n1475 GNDA.n1474 76.3222
R1520 GNDA.n1488 GNDA.n1487 76.3222
R1521 GNDA.n1386 GNDA.n106 76.3222
R1522 GNDA.n1458 GNDA.n1457 76.3222
R1523 GNDA.n1459 GNDA.n101 76.3222
R1524 GNDA.n1473 GNDA.n1472 76.3222
R1525 GNDA.n1474 GNDA.n93 76.3222
R1526 GNDA.n1489 GNDA.n1488 76.3222
R1527 GNDA.n930 GNDA.n907 76.3222
R1528 GNDA.n928 GNDA.n927 76.3222
R1529 GNDA.n923 GNDA.n910 76.3222
R1530 GNDA.n921 GNDA.n920 76.3222
R1531 GNDA.n916 GNDA.n913 76.3222
R1532 GNDA.n914 GNDA.n594 76.3222
R1533 GNDA.n960 GNDA.n959 76.3222
R1534 GNDA.n874 GNDA.n759 76.3222
R1535 GNDA.n873 GNDA.n762 76.3222
R1536 GNDA.n796 GNDA.n795 76.3222
R1537 GNDA.n799 GNDA.n798 76.3222
R1538 GNDA.n811 GNDA.n810 76.3222
R1539 GNDA.n814 GNDA.n813 76.3222
R1540 GNDA.n884 GNDA.n883 76.3222
R1541 GNDA.n883 GNDA.n882 76.3222
R1542 GNDA.n875 GNDA.n874 76.3222
R1543 GNDA.n791 GNDA.n762 76.3222
R1544 GNDA.n797 GNDA.n796 76.3222
R1545 GNDA.n798 GNDA.n785 76.3222
R1546 GNDA.n812 GNDA.n811 76.3222
R1547 GNDA.n813 GNDA.n582 76.3222
R1548 GNDA.n915 GNDA.n914 76.3222
R1549 GNDA.n913 GNDA.n911 76.3222
R1550 GNDA.n922 GNDA.n921 76.3222
R1551 GNDA.n910 GNDA.n908 76.3222
R1552 GNDA.n929 GNDA.n928 76.3222
R1553 GNDA.n907 GNDA.n749 76.3222
R1554 GNDA.n1524 GNDA.n1523 76.3222
R1555 GNDA.n1521 GNDA.n1520 76.3222
R1556 GNDA.n1508 GNDA.n82 76.3222
R1557 GNDA.n1507 GNDA.n1506 76.3222
R1558 GNDA.n1496 GNDA.n86 76.3222
R1559 GNDA.n1495 GNDA.n1494 76.3222
R1560 GNDA.n1514 GNDA.n79 76.3222
R1561 GNDA.n1517 GNDA.n1516 76.3222
R1562 GNDA.n1512 GNDA.n1511 76.3222
R1563 GNDA.n1503 GNDA.n1502 76.3222
R1564 GNDA.n1500 GNDA.n1499 76.3222
R1565 GNDA.n1491 GNDA.n1490 76.3222
R1566 GNDA.n693 GNDA.n601 76.3222
R1567 GNDA.n698 GNDA.n600 76.3222
R1568 GNDA.n706 GNDA.n599 76.3222
R1569 GNDA.n711 GNDA.n598 76.3222
R1570 GNDA.n719 GNDA.n597 76.3222
R1571 GNDA.n724 GNDA.n596 76.3222
R1572 GNDA.n1551 GNDA.n1550 76.3222
R1573 GNDA.n1548 GNDA.n1547 76.3222
R1574 GNDA.n1543 GNDA.n1542 76.3222
R1575 GNDA.n1540 GNDA.n1539 76.3222
R1576 GNDA.n1535 GNDA.n1534 76.3222
R1577 GNDA.n1532 GNDA.n1531 76.3222
R1578 GNDA.n961 GNDA.n960 76.3222
R1579 GNDA.n726 GNDA.n609 76.3222
R1580 GNDA.n385 GNDA.n380 76.3222
R1581 GNDA.n503 GNDA.n502 76.3222
R1582 GNDA.n466 GNDA.n386 76.3222
R1583 GNDA.n477 GNDA.n476 76.3222
R1584 GNDA.n480 GNDA.n479 76.3222
R1585 GNDA.n489 GNDA.n488 76.3222
R1586 GNDA.n492 GNDA.n491 76.3222
R1587 GNDA.n1060 GNDA.n1059 76.3222
R1588 GNDA.n1057 GNDA.n1056 76.3222
R1589 GNDA.n1052 GNDA.n345 76.3222
R1590 GNDA.n1050 GNDA.n1049 76.3222
R1591 GNDA.n1045 GNDA.n354 76.3222
R1592 GNDA.n1043 GNDA.n1042 76.3222
R1593 GNDA.n502 GNDA.n501 76.3222
R1594 GNDA.n467 GNDA.n466 76.3222
R1595 GNDA.n478 GNDA.n477 76.3222
R1596 GNDA.n479 GNDA.n462 76.3222
R1597 GNDA.n490 GNDA.n489 76.3222
R1598 GNDA.n491 GNDA.n333 76.3222
R1599 GNDA.n382 GNDA.n380 76.3222
R1600 GNDA.n306 GNDA.n305 76.3222
R1601 GNDA.n307 GNDA.n139 76.3222
R1602 GNDA.n314 GNDA.n313 76.3222
R1603 GNDA.n315 GNDA.n137 76.3222
R1604 GNDA.n322 GNDA.n321 76.3222
R1605 GNDA.n323 GNDA.n132 76.3222
R1606 GNDA.n1380 GNDA.n114 76.3222
R1607 GNDA.n1378 GNDA.n1377 76.3222
R1608 GNDA.n1373 GNDA.n122 76.3222
R1609 GNDA.n1371 GNDA.n1370 76.3222
R1610 GNDA.n1366 GNDA.n131 76.3222
R1611 GNDA.n1364 GNDA.n1363 76.3222
R1612 GNDA.n273 GNDA.n272 76.3222
R1613 GNDA.n233 GNDA.n153 76.3222
R1614 GNDA.n244 GNDA.n243 76.3222
R1615 GNDA.n247 GNDA.n246 76.3222
R1616 GNDA.n256 GNDA.n255 76.3222
R1617 GNDA.n262 GNDA.n261 76.3222
R1618 GNDA.n279 GNDA.n278 76.3222
R1619 GNDA.n278 GNDA.n151 76.3222
R1620 GNDA.n272 GNDA.n271 76.3222
R1621 GNDA.n234 GNDA.n233 76.3222
R1622 GNDA.n245 GNDA.n244 76.3222
R1623 GNDA.n246 GNDA.n229 76.3222
R1624 GNDA.n257 GNDA.n256 76.3222
R1625 GNDA.n261 GNDA.n260 76.3222
R1626 GNDA.n324 GNDA.n323 76.3222
R1627 GNDA.n321 GNDA.n320 76.3222
R1628 GNDA.n316 GNDA.n315 76.3222
R1629 GNDA.n313 GNDA.n312 76.3222
R1630 GNDA.n308 GNDA.n307 76.3222
R1631 GNDA.n305 GNDA.n304 76.3222
R1632 GNDA.n134 GNDA.n133 76.3222
R1633 GNDA.n128 GNDA.n127 76.3222
R1634 GNDA.n125 GNDA.n124 76.3222
R1635 GNDA.n119 GNDA.n118 76.3222
R1636 GNDA.n116 GNDA.n112 76.3222
R1637 GNDA.n1384 GNDA.n1383 76.3222
R1638 GNDA.n1365 GNDA.n1364 76.3222
R1639 GNDA.n131 GNDA.n123 76.3222
R1640 GNDA.n1372 GNDA.n1371 76.3222
R1641 GNDA.n122 GNDA.n115 76.3222
R1642 GNDA.n1379 GNDA.n1378 76.3222
R1643 GNDA.n258 GNDA.n114 76.3222
R1644 GNDA.n357 GNDA.n356 76.3222
R1645 GNDA.n351 GNDA.n350 76.3222
R1646 GNDA.n348 GNDA.n347 76.3222
R1647 GNDA.n342 GNDA.n341 76.3222
R1648 GNDA.n339 GNDA.n338 76.3222
R1649 GNDA.n336 GNDA.n331 76.3222
R1650 GNDA.n1044 GNDA.n1043 76.3222
R1651 GNDA.n354 GNDA.n346 76.3222
R1652 GNDA.n1051 GNDA.n1050 76.3222
R1653 GNDA.n345 GNDA.n335 76.3222
R1654 GNDA.n1058 GNDA.n1057 76.3222
R1655 GNDA.n1061 GNDA.n1060 76.3222
R1656 GNDA.n1213 GNDA.n1212 76.3222
R1657 GNDA.n1177 GNDA.n1176 76.3222
R1658 GNDA.n1188 GNDA.n1187 76.3222
R1659 GNDA.n1189 GNDA.n1172 76.3222
R1660 GNDA.n1200 GNDA.n1199 76.3222
R1661 GNDA.n1202 GNDA.n1201 76.3222
R1662 GNDA.n1560 GNDA.n61 76.3222
R1663 GNDA.n34 GNDA.n8 76.3222
R1664 GNDA.n33 GNDA.n7 76.3222
R1665 GNDA.n1227 GNDA.n2 76.3222
R1666 GNDA.n1230 GNDA.n1229 76.3222
R1667 GNDA.n1225 GNDA.n1224 76.3222
R1668 GNDA.n1219 GNDA.n1218 76.3222
R1669 GNDA.n11 GNDA.n6 76.3222
R1670 GNDA.n1615 GNDA.n1614 76.3222
R1671 GNDA.n1232 GNDA.n4 76.3222
R1672 GNDA.n1231 GNDA.n1222 76.3222
R1673 GNDA.n1239 GNDA.n1238 76.3222
R1674 GNDA.n1221 GNDA.n1094 76.3222
R1675 GNDA.t7 GNDA.n974 75.0005
R1676 GNDA.n975 GNDA.t7 75.0005
R1677 GNDA.t14 GNDA.n972 75.0005
R1678 GNDA.n992 GNDA.t14 75.0005
R1679 GNDA.t22 GNDA.n20 74.7579
R1680 GNDA.t22 GNDA.n5 74.7579
R1681 GNDA.n1207 GNDA.n1206 74.5978
R1682 GNDA.n1207 GNDA.n1118 74.5978
R1683 GNDA.n1295 GNDA.n1294 74.5978
R1684 GNDA.n1296 GNDA.n1295 74.5978
R1685 GNDA.n496 GNDA.n495 74.5978
R1686 GNDA.n496 GNDA.n408 74.5978
R1687 GNDA.n639 GNDA.n613 74.5978
R1688 GNDA.n640 GNDA.n639 74.5978
R1689 GNDA.n1482 GNDA.n1481 74.5978
R1690 GNDA.n1483 GNDA.n1482 74.5978
R1691 GNDA.n818 GNDA.n817 74.5978
R1692 GNDA.n819 GNDA.n818 74.5978
R1693 GNDA.n266 GNDA.n265 74.5978
R1694 GNDA.n266 GNDA.n175 74.5978
R1695 GNDA.n885 GNDA.t16 70.5764
R1696 GNDA.n1136 GNDA.n1108 69.3109
R1697 GNDA.n1139 GNDA.n1108 69.3109
R1698 GNDA.n1328 GNDA.n1327 69.3109
R1699 GNDA.n1327 GNDA.n1326 69.3109
R1700 GNDA.n426 GNDA.n398 69.3109
R1701 GNDA.n429 GNDA.n398 69.3109
R1702 GNDA.n672 GNDA.n671 69.3109
R1703 GNDA.n671 GNDA.n670 69.3109
R1704 GNDA.n1434 GNDA.n1433 69.3109
R1705 GNDA.n1433 GNDA.n1432 69.3109
R1706 GNDA.n851 GNDA.n850 69.3109
R1707 GNDA.n850 GNDA.n849 69.3109
R1708 GNDA.n193 GNDA.n165 69.3109
R1709 GNDA.n196 GNDA.n165 69.3109
R1710 GNDA.t28 GNDA.n1107 65.8183
R1711 GNDA.t28 GNDA.n1105 65.8183
R1712 GNDA.t28 GNDA.n1103 65.8183
R1713 GNDA.t28 GNDA.n1110 65.8183
R1714 GNDA.t28 GNDA.n1111 65.8183
R1715 GNDA.t28 GNDA.n1112 65.8183
R1716 GNDA.t28 GNDA.n1113 65.8183
R1717 GNDA.t28 GNDA.n1106 65.8183
R1718 GNDA.t28 GNDA.n1104 65.8183
R1719 GNDA.t28 GNDA.n1102 65.8183
R1720 GNDA.t28 GNDA.n1101 65.8183
R1721 GNDA.n1307 GNDA.t33 65.8183
R1722 GNDA.n1304 GNDA.t33 65.8183
R1723 GNDA.n1298 GNDA.t33 65.8183
R1724 GNDA.n1313 GNDA.t33 65.8183
R1725 GNDA.n1083 GNDA.t33 65.8183
R1726 GNDA.n1320 GNDA.t33 65.8183
R1727 GNDA.n1080 GNDA.t33 65.8183
R1728 GNDA.n1076 GNDA.t33 65.8183
R1729 GNDA.n1333 GNDA.t33 65.8183
R1730 GNDA.n1339 GNDA.t33 65.8183
R1731 GNDA.n1073 GNDA.t33 65.8183
R1732 GNDA.t32 GNDA.n397 65.8183
R1733 GNDA.t32 GNDA.n395 65.8183
R1734 GNDA.t32 GNDA.n393 65.8183
R1735 GNDA.t32 GNDA.n400 65.8183
R1736 GNDA.t32 GNDA.n401 65.8183
R1737 GNDA.t32 GNDA.n402 65.8183
R1738 GNDA.t32 GNDA.n403 65.8183
R1739 GNDA.t32 GNDA.n396 65.8183
R1740 GNDA.t32 GNDA.n394 65.8183
R1741 GNDA.t32 GNDA.n392 65.8183
R1742 GNDA.t32 GNDA.n391 65.8183
R1743 GNDA.n651 GNDA.t26 65.8183
R1744 GNDA.n648 GNDA.t26 65.8183
R1745 GNDA.n642 GNDA.t26 65.8183
R1746 GNDA.n657 GNDA.t26 65.8183
R1747 GNDA.n633 GNDA.t26 65.8183
R1748 GNDA.n664 GNDA.t26 65.8183
R1749 GNDA.n630 GNDA.t26 65.8183
R1750 GNDA.n673 GNDA.t26 65.8183
R1751 GNDA.n679 GNDA.t26 65.8183
R1752 GNDA.n624 GNDA.t26 65.8183
R1753 GNDA.n686 GNDA.t26 65.8183
R1754 GNDA.n1413 GNDA.t21 65.8183
R1755 GNDA.n1410 GNDA.t21 65.8183
R1756 GNDA.n1404 GNDA.t21 65.8183
R1757 GNDA.n1419 GNDA.t21 65.8183
R1758 GNDA.n1399 GNDA.t21 65.8183
R1759 GNDA.n1426 GNDA.t21 65.8183
R1760 GNDA.n1396 GNDA.t21 65.8183
R1761 GNDA.n1392 GNDA.t21 65.8183
R1762 GNDA.n1439 GNDA.t21 65.8183
R1763 GNDA.n1445 GNDA.t21 65.8183
R1764 GNDA.n108 GNDA.t21 65.8183
R1765 GNDA.n1451 GNDA.t21 65.8183
R1766 GNDA.n1464 GNDA.t21 65.8183
R1767 GNDA.n1466 GNDA.t21 65.8183
R1768 GNDA.n1479 GNDA.t21 65.8183
R1769 GNDA.n830 GNDA.t23 65.8183
R1770 GNDA.n827 GNDA.t23 65.8183
R1771 GNDA.n821 GNDA.t23 65.8183
R1772 GNDA.n836 GNDA.t23 65.8183
R1773 GNDA.n774 GNDA.t23 65.8183
R1774 GNDA.n843 GNDA.t23 65.8183
R1775 GNDA.n771 GNDA.t23 65.8183
R1776 GNDA.n852 GNDA.t23 65.8183
R1777 GNDA.n858 GNDA.t23 65.8183
R1778 GNDA.n860 GNDA.t23 65.8183
R1779 GNDA.n866 GNDA.t23 65.8183
R1780 GNDA.n869 GNDA.t23 65.8183
R1781 GNDA.n788 GNDA.t23 65.8183
R1782 GNDA.n803 GNDA.t23 65.8183
R1783 GNDA.n805 GNDA.t23 65.8183
R1784 GNDA.n622 GNDA.t26 65.8183
R1785 GNDA.n702 GNDA.t26 65.8183
R1786 GNDA.n617 GNDA.t26 65.8183
R1787 GNDA.n715 GNDA.t26 65.8183
R1788 GNDA.n497 GNDA.t32 65.8183
R1789 GNDA.t32 GNDA.n405 65.8183
R1790 GNDA.t32 GNDA.n406 65.8183
R1791 GNDA.t32 GNDA.n407 65.8183
R1792 GNDA.t25 GNDA.n164 65.8183
R1793 GNDA.t25 GNDA.n162 65.8183
R1794 GNDA.t25 GNDA.n160 65.8183
R1795 GNDA.t25 GNDA.n167 65.8183
R1796 GNDA.t25 GNDA.n168 65.8183
R1797 GNDA.t25 GNDA.n169 65.8183
R1798 GNDA.t25 GNDA.n170 65.8183
R1799 GNDA.t25 GNDA.n163 65.8183
R1800 GNDA.t25 GNDA.n161 65.8183
R1801 GNDA.t25 GNDA.n159 65.8183
R1802 GNDA.t25 GNDA.n158 65.8183
R1803 GNDA.n267 GNDA.t25 65.8183
R1804 GNDA.t25 GNDA.n172 65.8183
R1805 GNDA.t25 GNDA.n173 65.8183
R1806 GNDA.t25 GNDA.n174 65.8183
R1807 GNDA.n1346 GNDA.t33 65.8183
R1808 GNDA.n1255 GNDA.t33 65.8183
R1809 GNDA.n1276 GNDA.t33 65.8183
R1810 GNDA.n1278 GNDA.t33 65.8183
R1811 GNDA.n1208 GNDA.t28 65.8183
R1812 GNDA.t28 GNDA.n1115 65.8183
R1813 GNDA.t28 GNDA.n1116 65.8183
R1814 GNDA.t28 GNDA.n1117 65.8183
R1815 GNDA.t28 GNDA.n1108 57.8461
R1816 GNDA.n1327 GNDA.t33 57.8461
R1817 GNDA.t32 GNDA.n398 57.8461
R1818 GNDA.n671 GNDA.t26 57.8461
R1819 GNDA.n1433 GNDA.t21 57.8461
R1820 GNDA.n850 GNDA.t23 57.8461
R1821 GNDA.t25 GNDA.n165 57.8461
R1822 GNDA.n1482 GNDA.t21 55.2026
R1823 GNDA.n818 GNDA.t23 55.2026
R1824 GNDA.n639 GNDA.t26 55.2026
R1825 GNDA.t32 GNDA.n496 55.2026
R1826 GNDA.t25 GNDA.n266 55.2026
R1827 GNDA.n1295 GNDA.t33 55.2026
R1828 GNDA.t28 GNDA.n1207 55.2026
R1829 GNDA.n894 GNDA.t24 54.3786
R1830 GNDA.n1209 GNDA.n1208 53.3664
R1831 GNDA.n1180 GNDA.n1115 53.3664
R1832 GNDA.n1182 GNDA.n1116 53.3664
R1833 GNDA.n1194 GNDA.n1117 53.3664
R1834 GNDA.n1101 GNDA.n1099 53.3664
R1835 GNDA.n1124 GNDA.n1102 53.3664
R1836 GNDA.n1128 GNDA.n1104 53.3664
R1837 GNDA.n1132 GNDA.n1106 53.3664
R1838 GNDA.n1143 GNDA.n1113 53.3664
R1839 GNDA.n1147 GNDA.n1112 53.3664
R1840 GNDA.n1151 GNDA.n1111 53.3664
R1841 GNDA.n1154 GNDA.n1110 53.3664
R1842 GNDA.n1167 GNDA.n1103 53.3664
R1843 GNDA.n1164 GNDA.n1105 53.3664
R1844 GNDA.n1160 GNDA.n1107 53.3664
R1845 GNDA.n1157 GNDA.n1107 53.3664
R1846 GNDA.n1161 GNDA.n1105 53.3664
R1847 GNDA.n1165 GNDA.n1103 53.3664
R1848 GNDA.n1152 GNDA.n1110 53.3664
R1849 GNDA.n1148 GNDA.n1111 53.3664
R1850 GNDA.n1144 GNDA.n1112 53.3664
R1851 GNDA.n1140 GNDA.n1113 53.3664
R1852 GNDA.n1135 GNDA.n1106 53.3664
R1853 GNDA.n1131 GNDA.n1104 53.3664
R1854 GNDA.n1127 GNDA.n1102 53.3664
R1855 GNDA.n1123 GNDA.n1101 53.3664
R1856 GNDA.n1346 GNDA.n1345 53.3664
R1857 GNDA.n1255 GNDA.n1072 53.3664
R1858 GNDA.n1276 GNDA.n1275 53.3664
R1859 GNDA.n1279 GNDA.n1278 53.3664
R1860 GNDA.n1344 GNDA.n1073 53.3664
R1861 GNDA.n1340 GNDA.n1339 53.3664
R1862 GNDA.n1333 GNDA.n1075 53.3664
R1863 GNDA.n1332 GNDA.n1076 53.3664
R1864 GNDA.n1322 GNDA.n1080 53.3664
R1865 GNDA.n1320 GNDA.n1319 53.3664
R1866 GNDA.n1315 GNDA.n1083 53.3664
R1867 GNDA.n1313 GNDA.n1312 53.3664
R1868 GNDA.n1299 GNDA.n1298 53.3664
R1869 GNDA.n1304 GNDA.n1303 53.3664
R1870 GNDA.n1307 GNDA.n1306 53.3664
R1871 GNDA.n1308 GNDA.n1307 53.3664
R1872 GNDA.n1305 GNDA.n1304 53.3664
R1873 GNDA.n1298 GNDA.n1087 53.3664
R1874 GNDA.n1314 GNDA.n1313 53.3664
R1875 GNDA.n1083 GNDA.n1081 53.3664
R1876 GNDA.n1321 GNDA.n1320 53.3664
R1877 GNDA.n1080 GNDA.n1078 53.3664
R1878 GNDA.n1329 GNDA.n1076 53.3664
R1879 GNDA.n1334 GNDA.n1333 53.3664
R1880 GNDA.n1339 GNDA.n1338 53.3664
R1881 GNDA.n1341 GNDA.n1073 53.3664
R1882 GNDA.n498 GNDA.n497 53.3664
R1883 GNDA.n470 GNDA.n405 53.3664
R1884 GNDA.n472 GNDA.n406 53.3664
R1885 GNDA.n484 GNDA.n407 53.3664
R1886 GNDA.n391 GNDA.n389 53.3664
R1887 GNDA.n414 GNDA.n392 53.3664
R1888 GNDA.n418 GNDA.n394 53.3664
R1889 GNDA.n422 GNDA.n396 53.3664
R1890 GNDA.n433 GNDA.n403 53.3664
R1891 GNDA.n437 GNDA.n402 53.3664
R1892 GNDA.n441 GNDA.n401 53.3664
R1893 GNDA.n444 GNDA.n400 53.3664
R1894 GNDA.n457 GNDA.n393 53.3664
R1895 GNDA.n454 GNDA.n395 53.3664
R1896 GNDA.n450 GNDA.n397 53.3664
R1897 GNDA.n447 GNDA.n397 53.3664
R1898 GNDA.n451 GNDA.n395 53.3664
R1899 GNDA.n455 GNDA.n393 53.3664
R1900 GNDA.n442 GNDA.n400 53.3664
R1901 GNDA.n438 GNDA.n401 53.3664
R1902 GNDA.n434 GNDA.n402 53.3664
R1903 GNDA.n430 GNDA.n403 53.3664
R1904 GNDA.n425 GNDA.n396 53.3664
R1905 GNDA.n421 GNDA.n394 53.3664
R1906 GNDA.n417 GNDA.n392 53.3664
R1907 GNDA.n413 GNDA.n391 53.3664
R1908 GNDA.n623 GNDA.n622 53.3664
R1909 GNDA.n702 GNDA.n701 53.3664
R1910 GNDA.n618 GNDA.n617 53.3664
R1911 GNDA.n715 GNDA.n714 53.3664
R1912 GNDA.n687 GNDA.n686 53.3664
R1913 GNDA.n684 GNDA.n624 53.3664
R1914 GNDA.n680 GNDA.n679 53.3664
R1915 GNDA.n673 GNDA.n626 53.3664
R1916 GNDA.n666 GNDA.n630 53.3664
R1917 GNDA.n664 GNDA.n663 53.3664
R1918 GNDA.n659 GNDA.n633 53.3664
R1919 GNDA.n657 GNDA.n656 53.3664
R1920 GNDA.n643 GNDA.n642 53.3664
R1921 GNDA.n648 GNDA.n647 53.3664
R1922 GNDA.n651 GNDA.n650 53.3664
R1923 GNDA.n652 GNDA.n651 53.3664
R1924 GNDA.n649 GNDA.n648 53.3664
R1925 GNDA.n642 GNDA.n637 53.3664
R1926 GNDA.n658 GNDA.n657 53.3664
R1927 GNDA.n633 GNDA.n631 53.3664
R1928 GNDA.n665 GNDA.n664 53.3664
R1929 GNDA.n630 GNDA.n628 53.3664
R1930 GNDA.n674 GNDA.n673 53.3664
R1931 GNDA.n679 GNDA.n678 53.3664
R1932 GNDA.n681 GNDA.n624 53.3664
R1933 GNDA.n686 GNDA.n685 53.3664
R1934 GNDA.n1452 GNDA.n1451 53.3664
R1935 GNDA.n1464 GNDA.n1463 53.3664
R1936 GNDA.n1467 GNDA.n1466 53.3664
R1937 GNDA.n1479 GNDA.n1478 53.3664
R1938 GNDA.n1450 GNDA.n108 53.3664
R1939 GNDA.n1446 GNDA.n1445 53.3664
R1940 GNDA.n1439 GNDA.n1391 53.3664
R1941 GNDA.n1438 GNDA.n1392 53.3664
R1942 GNDA.n1428 GNDA.n1396 53.3664
R1943 GNDA.n1426 GNDA.n1425 53.3664
R1944 GNDA.n1421 GNDA.n1399 53.3664
R1945 GNDA.n1419 GNDA.n1418 53.3664
R1946 GNDA.n1405 GNDA.n1404 53.3664
R1947 GNDA.n1410 GNDA.n1409 53.3664
R1948 GNDA.n1413 GNDA.n1412 53.3664
R1949 GNDA.n1414 GNDA.n1413 53.3664
R1950 GNDA.n1411 GNDA.n1410 53.3664
R1951 GNDA.n1404 GNDA.n1403 53.3664
R1952 GNDA.n1420 GNDA.n1419 53.3664
R1953 GNDA.n1399 GNDA.n1397 53.3664
R1954 GNDA.n1427 GNDA.n1426 53.3664
R1955 GNDA.n1396 GNDA.n1394 53.3664
R1956 GNDA.n1435 GNDA.n1392 53.3664
R1957 GNDA.n1440 GNDA.n1439 53.3664
R1958 GNDA.n1445 GNDA.n1444 53.3664
R1959 GNDA.n1447 GNDA.n108 53.3664
R1960 GNDA.n1451 GNDA.n104 53.3664
R1961 GNDA.n1465 GNDA.n1464 53.3664
R1962 GNDA.n1466 GNDA.n99 53.3664
R1963 GNDA.n1480 GNDA.n1479 53.3664
R1964 GNDA.n869 GNDA.n868 53.3664
R1965 GNDA.n788 GNDA.n764 53.3664
R1966 GNDA.n803 GNDA.n802 53.3664
R1967 GNDA.n806 GNDA.n805 53.3664
R1968 GNDA.n867 GNDA.n866 53.3664
R1969 GNDA.n860 GNDA.n765 53.3664
R1970 GNDA.n859 GNDA.n858 53.3664
R1971 GNDA.n852 GNDA.n767 53.3664
R1972 GNDA.n845 GNDA.n771 53.3664
R1973 GNDA.n843 GNDA.n842 53.3664
R1974 GNDA.n838 GNDA.n774 53.3664
R1975 GNDA.n836 GNDA.n835 53.3664
R1976 GNDA.n822 GNDA.n821 53.3664
R1977 GNDA.n827 GNDA.n826 53.3664
R1978 GNDA.n830 GNDA.n829 53.3664
R1979 GNDA.n831 GNDA.n830 53.3664
R1980 GNDA.n828 GNDA.n827 53.3664
R1981 GNDA.n821 GNDA.n778 53.3664
R1982 GNDA.n837 GNDA.n836 53.3664
R1983 GNDA.n774 GNDA.n772 53.3664
R1984 GNDA.n844 GNDA.n843 53.3664
R1985 GNDA.n771 GNDA.n769 53.3664
R1986 GNDA.n853 GNDA.n852 53.3664
R1987 GNDA.n858 GNDA.n857 53.3664
R1988 GNDA.n861 GNDA.n860 53.3664
R1989 GNDA.n866 GNDA.n865 53.3664
R1990 GNDA.n870 GNDA.n869 53.3664
R1991 GNDA.n789 GNDA.n788 53.3664
R1992 GNDA.n804 GNDA.n803 53.3664
R1993 GNDA.n805 GNDA.n781 53.3664
R1994 GNDA.n622 GNDA.n619 53.3664
R1995 GNDA.n703 GNDA.n702 53.3664
R1996 GNDA.n617 GNDA.n614 53.3664
R1997 GNDA.n716 GNDA.n715 53.3664
R1998 GNDA.n497 GNDA.n390 53.3664
R1999 GNDA.n473 GNDA.n405 53.3664
R2000 GNDA.n483 GNDA.n406 53.3664
R2001 GNDA.n409 GNDA.n407 53.3664
R2002 GNDA.n268 GNDA.n267 53.3664
R2003 GNDA.n237 GNDA.n172 53.3664
R2004 GNDA.n239 GNDA.n173 53.3664
R2005 GNDA.n251 GNDA.n174 53.3664
R2006 GNDA.n158 GNDA.n156 53.3664
R2007 GNDA.n181 GNDA.n159 53.3664
R2008 GNDA.n185 GNDA.n161 53.3664
R2009 GNDA.n189 GNDA.n163 53.3664
R2010 GNDA.n200 GNDA.n170 53.3664
R2011 GNDA.n204 GNDA.n169 53.3664
R2012 GNDA.n208 GNDA.n168 53.3664
R2013 GNDA.n211 GNDA.n167 53.3664
R2014 GNDA.n224 GNDA.n160 53.3664
R2015 GNDA.n221 GNDA.n162 53.3664
R2016 GNDA.n217 GNDA.n164 53.3664
R2017 GNDA.n214 GNDA.n164 53.3664
R2018 GNDA.n218 GNDA.n162 53.3664
R2019 GNDA.n222 GNDA.n160 53.3664
R2020 GNDA.n209 GNDA.n167 53.3664
R2021 GNDA.n205 GNDA.n168 53.3664
R2022 GNDA.n201 GNDA.n169 53.3664
R2023 GNDA.n197 GNDA.n170 53.3664
R2024 GNDA.n192 GNDA.n163 53.3664
R2025 GNDA.n188 GNDA.n161 53.3664
R2026 GNDA.n184 GNDA.n159 53.3664
R2027 GNDA.n180 GNDA.n158 53.3664
R2028 GNDA.n267 GNDA.n157 53.3664
R2029 GNDA.n240 GNDA.n172 53.3664
R2030 GNDA.n250 GNDA.n173 53.3664
R2031 GNDA.n176 GNDA.n174 53.3664
R2032 GNDA.n1347 GNDA.n1346 53.3664
R2033 GNDA.n1256 GNDA.n1255 53.3664
R2034 GNDA.n1277 GNDA.n1276 53.3664
R2035 GNDA.n1278 GNDA.n1090 53.3664
R2036 GNDA.n1208 GNDA.n1100 53.3664
R2037 GNDA.n1183 GNDA.n1115 53.3664
R2038 GNDA.n1193 GNDA.n1116 53.3664
R2039 GNDA.n1119 GNDA.n1117 53.3664
R2040 GNDA.n1028 GNDA.n27 50.5752
R2041 GNDA.t24 GNDA.n893 49.7507
R2042 GNDA.n1359 GNDA.n0 13.4867
R2043 GNDA.n62 GNDA.n35 42.2728
R2044 GNDA.n1008 GNDA.n1007 38.9537
R2045 GNDA.t3 GNDA.n963 38.5425
R2046 GNDA.n963 GNDA.t24 37.0972
R2047 GNDA.n935 GNDA.n934 32.7993
R2048 GNDA.t13 GNDA.t15 30.3453
R2049 GNDA.n1003 GNDA.t1 30.3453
R2050 GNDA.t11 GNDA.t6 30.3453
R2051 GNDA.n1006 GNDA.n1005 28.6501
R2052 GNDA.n1156 GNDA.n1155 27.5561
R2053 GNDA.n1311 GNDA.n1310 27.5561
R2054 GNDA.n446 GNDA.n445 27.5561
R2055 GNDA.n655 GNDA.n654 27.5561
R2056 GNDA.n1417 GNDA.n1416 27.5561
R2057 GNDA.n834 GNDA.n833 27.5561
R2058 GNDA.n213 GNDA.n212 27.5561
R2059 GNDA.n1138 GNDA.n1137 23.6449
R2060 GNDA.n1325 GNDA.n1077 23.6449
R2061 GNDA.n428 GNDA.n427 23.6449
R2062 GNDA.n669 GNDA.n627 23.6449
R2063 GNDA.n1431 GNDA.n1393 23.6449
R2064 GNDA.n848 GNDA.n768 23.6449
R2065 GNDA.n195 GNDA.n194 23.6449
R2066 GNDA.n574 GNDA.n573 20.9605
R2067 GNDA.n1010 GNDA.n1009 17.4917
R2068 GNDA.n1579 GNDA.n48 17.0672
R2069 GNDA.n942 GNDA.n593 17.0672
R2070 GNDA.n1554 GNDA.n1553 17.0672
R2071 GNDA.n1015 GNDA.n1014 16.9605
R2072 GNDA.n1170 GNDA.n1169 16.0005
R2073 GNDA.n1169 GNDA.n1168 16.0005
R2074 GNDA.n1168 GNDA.n1166 16.0005
R2075 GNDA.n1166 GNDA.n1163 16.0005
R2076 GNDA.n1163 GNDA.n1162 16.0005
R2077 GNDA.n1162 GNDA.n1159 16.0005
R2078 GNDA.n1159 GNDA.n1158 16.0005
R2079 GNDA.n1158 GNDA.n1156 16.0005
R2080 GNDA.n1141 GNDA.n1138 16.0005
R2081 GNDA.n1142 GNDA.n1141 16.0005
R2082 GNDA.n1145 GNDA.n1142 16.0005
R2083 GNDA.n1146 GNDA.n1145 16.0005
R2084 GNDA.n1149 GNDA.n1146 16.0005
R2085 GNDA.n1150 GNDA.n1149 16.0005
R2086 GNDA.n1153 GNDA.n1150 16.0005
R2087 GNDA.n1155 GNDA.n1153 16.0005
R2088 GNDA.n1122 GNDA.n1121 16.0005
R2089 GNDA.n1125 GNDA.n1122 16.0005
R2090 GNDA.n1126 GNDA.n1125 16.0005
R2091 GNDA.n1129 GNDA.n1126 16.0005
R2092 GNDA.n1130 GNDA.n1129 16.0005
R2093 GNDA.n1134 GNDA.n1133 16.0005
R2094 GNDA.n1137 GNDA.n1134 16.0005
R2095 GNDA.n1089 GNDA.n1088 16.0005
R2096 GNDA.n1300 GNDA.n1088 16.0005
R2097 GNDA.n1301 GNDA.n1300 16.0005
R2098 GNDA.n1302 GNDA.n1301 16.0005
R2099 GNDA.n1302 GNDA.n1086 16.0005
R2100 GNDA.n1086 GNDA.n1085 16.0005
R2101 GNDA.n1309 GNDA.n1085 16.0005
R2102 GNDA.n1310 GNDA.n1309 16.0005
R2103 GNDA.n1325 GNDA.n1324 16.0005
R2104 GNDA.n1324 GNDA.n1323 16.0005
R2105 GNDA.n1323 GNDA.n1079 16.0005
R2106 GNDA.n1318 GNDA.n1079 16.0005
R2107 GNDA.n1318 GNDA.n1317 16.0005
R2108 GNDA.n1317 GNDA.n1316 16.0005
R2109 GNDA.n1316 GNDA.n1082 16.0005
R2110 GNDA.n1311 GNDA.n1082 16.0005
R2111 GNDA.n1343 GNDA.n1342 16.0005
R2112 GNDA.n1342 GNDA.n1074 16.0005
R2113 GNDA.n1337 GNDA.n1074 16.0005
R2114 GNDA.n1337 GNDA.n1336 16.0005
R2115 GNDA.n1336 GNDA.n1335 16.0005
R2116 GNDA.n1331 GNDA.n1330 16.0005
R2117 GNDA.n1330 GNDA.n1077 16.0005
R2118 GNDA.n460 GNDA.n459 16.0005
R2119 GNDA.n459 GNDA.n458 16.0005
R2120 GNDA.n458 GNDA.n456 16.0005
R2121 GNDA.n456 GNDA.n453 16.0005
R2122 GNDA.n453 GNDA.n452 16.0005
R2123 GNDA.n452 GNDA.n449 16.0005
R2124 GNDA.n449 GNDA.n448 16.0005
R2125 GNDA.n448 GNDA.n446 16.0005
R2126 GNDA.n431 GNDA.n428 16.0005
R2127 GNDA.n432 GNDA.n431 16.0005
R2128 GNDA.n435 GNDA.n432 16.0005
R2129 GNDA.n436 GNDA.n435 16.0005
R2130 GNDA.n439 GNDA.n436 16.0005
R2131 GNDA.n440 GNDA.n439 16.0005
R2132 GNDA.n443 GNDA.n440 16.0005
R2133 GNDA.n445 GNDA.n443 16.0005
R2134 GNDA.n412 GNDA.n411 16.0005
R2135 GNDA.n415 GNDA.n412 16.0005
R2136 GNDA.n416 GNDA.n415 16.0005
R2137 GNDA.n419 GNDA.n416 16.0005
R2138 GNDA.n420 GNDA.n419 16.0005
R2139 GNDA.n424 GNDA.n423 16.0005
R2140 GNDA.n427 GNDA.n424 16.0005
R2141 GNDA.n638 GNDA.n610 16.0005
R2142 GNDA.n644 GNDA.n638 16.0005
R2143 GNDA.n645 GNDA.n644 16.0005
R2144 GNDA.n646 GNDA.n645 16.0005
R2145 GNDA.n646 GNDA.n636 16.0005
R2146 GNDA.n636 GNDA.n635 16.0005
R2147 GNDA.n653 GNDA.n635 16.0005
R2148 GNDA.n654 GNDA.n653 16.0005
R2149 GNDA.n669 GNDA.n668 16.0005
R2150 GNDA.n668 GNDA.n667 16.0005
R2151 GNDA.n667 GNDA.n629 16.0005
R2152 GNDA.n662 GNDA.n629 16.0005
R2153 GNDA.n662 GNDA.n661 16.0005
R2154 GNDA.n661 GNDA.n660 16.0005
R2155 GNDA.n660 GNDA.n632 16.0005
R2156 GNDA.n655 GNDA.n632 16.0005
R2157 GNDA.n688 GNDA.n621 16.0005
R2158 GNDA.n683 GNDA.n621 16.0005
R2159 GNDA.n683 GNDA.n682 16.0005
R2160 GNDA.n682 GNDA.n625 16.0005
R2161 GNDA.n677 GNDA.n625 16.0005
R2162 GNDA.n676 GNDA.n675 16.0005
R2163 GNDA.n675 GNDA.n627 16.0005
R2164 GNDA.n1484 GNDA.n95 16.0005
R2165 GNDA.n1406 GNDA.n95 16.0005
R2166 GNDA.n1407 GNDA.n1406 16.0005
R2167 GNDA.n1408 GNDA.n1407 16.0005
R2168 GNDA.n1408 GNDA.n1402 16.0005
R2169 GNDA.n1402 GNDA.n1401 16.0005
R2170 GNDA.n1415 GNDA.n1401 16.0005
R2171 GNDA.n1416 GNDA.n1415 16.0005
R2172 GNDA.n1431 GNDA.n1430 16.0005
R2173 GNDA.n1430 GNDA.n1429 16.0005
R2174 GNDA.n1429 GNDA.n1395 16.0005
R2175 GNDA.n1424 GNDA.n1395 16.0005
R2176 GNDA.n1424 GNDA.n1423 16.0005
R2177 GNDA.n1423 GNDA.n1422 16.0005
R2178 GNDA.n1422 GNDA.n1398 16.0005
R2179 GNDA.n1417 GNDA.n1398 16.0005
R2180 GNDA.n1449 GNDA.n1448 16.0005
R2181 GNDA.n1448 GNDA.n1390 16.0005
R2182 GNDA.n1443 GNDA.n1390 16.0005
R2183 GNDA.n1443 GNDA.n1442 16.0005
R2184 GNDA.n1442 GNDA.n1441 16.0005
R2185 GNDA.n1437 GNDA.n1436 16.0005
R2186 GNDA.n1436 GNDA.n1393 16.0005
R2187 GNDA.n780 GNDA.n779 16.0005
R2188 GNDA.n823 GNDA.n779 16.0005
R2189 GNDA.n824 GNDA.n823 16.0005
R2190 GNDA.n825 GNDA.n824 16.0005
R2191 GNDA.n825 GNDA.n777 16.0005
R2192 GNDA.n777 GNDA.n776 16.0005
R2193 GNDA.n832 GNDA.n776 16.0005
R2194 GNDA.n833 GNDA.n832 16.0005
R2195 GNDA.n848 GNDA.n847 16.0005
R2196 GNDA.n847 GNDA.n846 16.0005
R2197 GNDA.n846 GNDA.n770 16.0005
R2198 GNDA.n841 GNDA.n770 16.0005
R2199 GNDA.n841 GNDA.n840 16.0005
R2200 GNDA.n840 GNDA.n839 16.0005
R2201 GNDA.n839 GNDA.n773 16.0005
R2202 GNDA.n834 GNDA.n773 16.0005
R2203 GNDA.n864 GNDA.n760 16.0005
R2204 GNDA.n864 GNDA.n863 16.0005
R2205 GNDA.n863 GNDA.n862 16.0005
R2206 GNDA.n862 GNDA.n766 16.0005
R2207 GNDA.n856 GNDA.n766 16.0005
R2208 GNDA.n855 GNDA.n854 16.0005
R2209 GNDA.n854 GNDA.n768 16.0005
R2210 GNDA.n227 GNDA.n226 16.0005
R2211 GNDA.n226 GNDA.n225 16.0005
R2212 GNDA.n225 GNDA.n223 16.0005
R2213 GNDA.n223 GNDA.n220 16.0005
R2214 GNDA.n220 GNDA.n219 16.0005
R2215 GNDA.n219 GNDA.n216 16.0005
R2216 GNDA.n216 GNDA.n215 16.0005
R2217 GNDA.n215 GNDA.n213 16.0005
R2218 GNDA.n198 GNDA.n195 16.0005
R2219 GNDA.n199 GNDA.n198 16.0005
R2220 GNDA.n202 GNDA.n199 16.0005
R2221 GNDA.n203 GNDA.n202 16.0005
R2222 GNDA.n206 GNDA.n203 16.0005
R2223 GNDA.n207 GNDA.n206 16.0005
R2224 GNDA.n210 GNDA.n207 16.0005
R2225 GNDA.n212 GNDA.n210 16.0005
R2226 GNDA.n179 GNDA.n178 16.0005
R2227 GNDA.n182 GNDA.n179 16.0005
R2228 GNDA.n183 GNDA.n182 16.0005
R2229 GNDA.n186 GNDA.n183 16.0005
R2230 GNDA.n187 GNDA.n186 16.0005
R2231 GNDA.n191 GNDA.n190 16.0005
R2232 GNDA.n194 GNDA.n191 16.0005
R2233 GNDA.n1014 GNDA.n560 16.0005
R2234 GNDA.n1010 GNDA.n560 16.0005
R2235 GNDA.n1529 GNDA.n76 15.5383
R2236 GNDA.n1357 GNDA.n327 15.5383
R2237 GNDA.t16 GNDA.n580 13.9723
R2238 GNDA.n980 GNDA.n977 13.6307
R2239 GNDA.n963 GNDA.n576 13.4881
R2240 GNDA.n1133 GNDA 12.9783
R2241 GNDA.n1331 GNDA 12.9783
R2242 GNDA.n423 GNDA 12.9783
R2243 GNDA GNDA.n676 12.9783
R2244 GNDA.n1437 GNDA 12.9783
R2245 GNDA GNDA.n855 12.9783
R2246 GNDA.n190 GNDA 12.9783
R2247 GNDA.n983 GNDA.n982 12.8005
R2248 GNDA.n984 GNDA.n983 12.8005
R2249 GNDA.n525 GNDA.n368 12.4126
R2250 GNDA.n302 GNDA.n301 12.4126
R2251 GNDA.n1603 GNDA.n1602 11.6369
R2252 GNDA.n1602 GNDA.n1601 11.6369
R2253 GNDA.n1601 GNDA.n39 11.6369
R2254 GNDA.n1595 GNDA.n39 11.6369
R2255 GNDA.n1595 GNDA.n1594 11.6369
R2256 GNDA.n1594 GNDA.n1593 11.6369
R2257 GNDA.n1593 GNDA.n44 11.6369
R2258 GNDA.n1587 GNDA.n44 11.6369
R2259 GNDA.n1587 GNDA.n1586 11.6369
R2260 GNDA.n1586 GNDA.n1585 11.6369
R2261 GNDA.n1585 GNDA.n48 11.6369
R2262 GNDA.n1563 GNDA.n1562 11.6369
R2263 GNDA.n1563 GNDA.n56 11.6369
R2264 GNDA.n1569 GNDA.n56 11.6369
R2265 GNDA.n1570 GNDA.n1569 11.6369
R2266 GNDA.n1571 GNDA.n1570 11.6369
R2267 GNDA.n1571 GNDA.n52 11.6369
R2268 GNDA.n1577 GNDA.n52 11.6369
R2269 GNDA.n1578 GNDA.n1577 11.6369
R2270 GNDA.n1579 GNDA.n1578 11.6369
R2271 GNDA.n587 GNDA.n585 11.6369
R2272 GNDA.n953 GNDA.n587 11.6369
R2273 GNDA.n953 GNDA.n952 11.6369
R2274 GNDA.n952 GNDA.n951 11.6369
R2275 GNDA.n951 GNDA.n588 11.6369
R2276 GNDA.n592 GNDA.n588 11.6369
R2277 GNDA.n944 GNDA.n592 11.6369
R2278 GNDA.n944 GNDA.n943 11.6369
R2279 GNDA.n943 GNDA.n942 11.6369
R2280 GNDA.n932 GNDA.n931 11.6369
R2281 GNDA.n931 GNDA.n906 11.6369
R2282 GNDA.n926 GNDA.n906 11.6369
R2283 GNDA.n926 GNDA.n925 11.6369
R2284 GNDA.n925 GNDA.n924 11.6369
R2285 GNDA.n924 GNDA.n909 11.6369
R2286 GNDA.n919 GNDA.n909 11.6369
R2287 GNDA.n919 GNDA.n918 11.6369
R2288 GNDA.n918 GNDA.n917 11.6369
R2289 GNDA.n917 GNDA.n912 11.6369
R2290 GNDA.n912 GNDA.n593 11.6369
R2291 GNDA.n728 GNDA.n606 11.6369
R2292 GNDA.n734 GNDA.n606 11.6369
R2293 GNDA.n735 GNDA.n734 11.6369
R2294 GNDA.n743 GNDA.n735 11.6369
R2295 GNDA.n743 GNDA.n742 11.6369
R2296 GNDA.n742 GNDA.n741 11.6369
R2297 GNDA.n741 GNDA.n736 11.6369
R2298 GNDA.n736 GNDA.n68 11.6369
R2299 GNDA.n1554 GNDA.n68 11.6369
R2300 GNDA.n1530 GNDA.n73 11.6369
R2301 GNDA.n1536 GNDA.n73 11.6369
R2302 GNDA.n1537 GNDA.n1536 11.6369
R2303 GNDA.n1538 GNDA.n1537 11.6369
R2304 GNDA.n1538 GNDA.n71 11.6369
R2305 GNDA.n1544 GNDA.n71 11.6369
R2306 GNDA.n1545 GNDA.n1544 11.6369
R2307 GNDA.n1546 GNDA.n1545 11.6369
R2308 GNDA.n1546 GNDA.n69 11.6369
R2309 GNDA.n1552 GNDA.n69 11.6369
R2310 GNDA.n1553 GNDA.n1552 11.6369
R2311 GNDA.n532 GNDA.n531 11.6369
R2312 GNDA.n534 GNDA.n532 11.6369
R2313 GNDA.n534 GNDA.n533 11.6369
R2314 GNDA.n533 GNDA.n365 11.6369
R2315 GNDA.n365 GNDA.n363 11.6369
R2316 GNDA.n542 GNDA.n363 11.6369
R2317 GNDA.n543 GNDA.n542 11.6369
R2318 GNDA.n544 GNDA.n543 11.6369
R2319 GNDA.n544 GNDA.n359 11.6369
R2320 GNDA.n550 GNDA.n359 11.6369
R2321 GNDA.n551 GNDA.n550 11.6369
R2322 GNDA.n509 GNDA.n508 11.6369
R2323 GNDA.n509 GNDA.n376 11.6369
R2324 GNDA.n515 GNDA.n376 11.6369
R2325 GNDA.n516 GNDA.n515 11.6369
R2326 GNDA.n517 GNDA.n372 11.6369
R2327 GNDA.n523 GNDA.n372 11.6369
R2328 GNDA.n524 GNDA.n523 11.6369
R2329 GNDA.n525 GNDA.n524 11.6369
R2330 GNDA.n284 GNDA.n149 11.6369
R2331 GNDA.n285 GNDA.n284 11.6369
R2332 GNDA.n287 GNDA.n285 11.6369
R2333 GNDA.n287 GNDA.n286 11.6369
R2334 GNDA.n294 GNDA.n293 11.6369
R2335 GNDA.n295 GNDA.n294 11.6369
R2336 GNDA.n295 GNDA.n142 11.6369
R2337 GNDA.n301 GNDA.n142 11.6369
R2338 GNDA.n303 GNDA.n140 11.6369
R2339 GNDA.n309 GNDA.n140 11.6369
R2340 GNDA.n310 GNDA.n309 11.6369
R2341 GNDA.n311 GNDA.n310 11.6369
R2342 GNDA.n311 GNDA.n138 11.6369
R2343 GNDA.n317 GNDA.n138 11.6369
R2344 GNDA.n318 GNDA.n317 11.6369
R2345 GNDA.n319 GNDA.n318 11.6369
R2346 GNDA.n319 GNDA.n136 11.6369
R2347 GNDA.n325 GNDA.n136 11.6369
R2348 GNDA.n326 GNDA.n325 11.6369
R2349 GNDA.n1263 GNDA.n1262 11.6369
R2350 GNDA.n1264 GNDA.n1263 11.6369
R2351 GNDA.n1265 GNDA.n1264 11.6369
R2352 GNDA.n1267 GNDA.n1265 11.6369
R2353 GNDA.n1267 GNDA.n1266 11.6369
R2354 GNDA.n1266 GNDA.n1248 11.6369
R2355 GNDA.n1285 GNDA.n1248 11.6369
R2356 GNDA.n1286 GNDA.n1285 11.6369
R2357 GNDA.n1287 GNDA.n1286 11.6369
R2358 GNDA.n1287 GNDA.n77 11.6369
R2359 GNDA.n1528 GNDA.n77 11.6369
R2360 GNDA.n557 GNDA.n554 11.6369
R2361 GNDA.n1033 GNDA.n557 11.6369
R2362 GNDA.n1033 GNDA.n1032 11.6369
R2363 GNDA.n1032 GNDA.n1031 11.6369
R2364 GNDA.n1031 GNDA.n558 11.6369
R2365 GNDA.n1025 GNDA.n1024 11.6369
R2366 GNDA.n1024 GNDA.n1023 11.6369
R2367 GNDA.n1023 GNDA.n1017 11.6369
R2368 GNDA.n1017 GNDA.n1016 11.6369
R2369 GNDA.n1016 GNDA.n13 11.6369
R2370 GNDA.t24 GNDA.n580 11.5635
R2371 GNDA.n508 GNDA.n507 11.3514
R2372 GNDA.n277 GNDA.n149 11.3514
R2373 GNDA.n1562 GNDA.n1561 11.249
R2374 GNDA.n585 GNDA.n583 11.249
R2375 GNDA.n728 GNDA.n727 11.249
R2376 GNDA.n1025 GNDA.n1015 10.4732
R2377 GNDA.n517 GNDA 10.3439
R2378 GNDA.n293 GNDA 10.3439
R2379 GNDA.n979 GNDA.n575 9.723
R2380 GNDA.n982 GNDA.n981 9.3005
R2381 GNDA.n983 GNDA.n978 9.3005
R2382 GNDA.n531 GNDA.n368 8.79242
R2383 GNDA.n303 GNDA.n302 8.79242
R2384 GNDA.n1603 GNDA.n38 8.53383
R2385 GNDA.n935 GNDA.n932 8.53383
R2386 GNDA.n1530 GNDA.n1529 8.53383
R2387 GNDA.n1262 GNDA.n327 8.53383
R2388 GNDA.n554 GNDA.n552 8.53383
R2389 GNDA.n888 GNDA.n758 8.41193
R2390 GNDA.n1171 GNDA.n1170 8.35606
R2391 GNDA.n1092 GNDA.n1089 8.35606
R2392 GNDA.n461 GNDA.n460 8.35606
R2393 GNDA.n722 GNDA.n610 8.35606
R2394 GNDA.n1485 GNDA.n1484 8.35606
R2395 GNDA.n784 GNDA.n780 8.35606
R2396 GNDA.n228 GNDA.n227 8.35606
R2397 GNDA.n574 GNDA.n572 7.93895
R2398 GNDA.n1009 GNDA.n1008 7.70747
R2399 GNDA.n936 GNDA.n905 7.02221
R2400 GNDA.n889 GNDA.n888 6.58336
R2401 GNDA.n890 GNDA.n889 6.58336
R2402 GNDA.n890 GNDA.n754 6.58336
R2403 GNDA.n896 GNDA.n754 6.58336
R2404 GNDA.n898 GNDA.n897 6.58336
R2405 GNDA.n898 GNDA.n750 6.58336
R2406 GNDA.n904 GNDA.n750 6.58336
R2407 GNDA.n905 GNDA.n904 6.58336
R2408 GNDA.n1009 GNDA.n561 6.36092
R2409 GNDA.n897 GNDA 5.85193
R2410 GNDA.n998 GNDA.n971 5.81868
R2411 GNDA.n998 GNDA.n997 5.81868
R2412 GNDA.n997 GNDA.n995 5.81868
R2413 GNDA.n995 GNDA.n976 5.81868
R2414 GNDA.n989 GNDA.n976 5.81868
R2415 GNDA.n1008 GNDA.n1006 5.21178
R2416 GNDA.n879 GNDA.n878 4.6085
R2417 GNDA.n506 GNDA.n381 4.6085
R2418 GNDA.n276 GNDA.n152 4.6085
R2419 GNDA.n1525 GNDA.n75 4.55161
R2420 GNDA.n1362 GNDA.n1361 4.55161
R2421 GNDA.n1041 GNDA.n1040 4.55161
R2422 GNDA.n1610 GNDA.n10 4.55161
R2423 GNDA.n979 GNDA.n978 4.5005
R2424 GNDA.n565 GNDA.n563 4.5005
R2425 GNDA.n566 GNDA.n564 4.5005
R2426 GNDA.n568 GNDA.n567 4.5005
R2427 GNDA.n552 GNDA.n551 4.39646
R2428 GNDA.n327 GNDA.n326 4.39646
R2429 GNDA.n1529 GNDA.n1528 4.39646
R2430 GNDA.n38 GNDA.n13 4.39646
R2431 GNDA.n727 GNDA.n723 4.3013
R2432 GNDA.n1561 GNDA.n60 4.3013
R2433 GNDA.n984 GNDA.n977 4.26767
R2434 GNDA.n982 GNDA.n977 4.26767
R2435 GNDA.n1492 GNDA.n89 4.26717
R2436 GNDA.n1498 GNDA.n89 4.26717
R2437 GNDA.n1498 GNDA.n87 4.26717
R2438 GNDA.n1504 GNDA.n87 4.26717
R2439 GNDA.n1504 GNDA.n85 4.26717
R2440 GNDA.n1510 GNDA.n85 4.26717
R2441 GNDA.n1518 GNDA.n83 4.26717
R2442 GNDA.n1518 GNDA.n81 4.26717
R2443 GNDA.n81 GNDA.n80 4.26717
R2444 GNDA.n1525 GNDA.n80 4.26717
R2445 GNDA.n1381 GNDA.n111 4.26717
R2446 GNDA.n1381 GNDA.n113 4.26717
R2447 GNDA.n1376 GNDA.n113 4.26717
R2448 GNDA.n1376 GNDA.n1375 4.26717
R2449 GNDA.n1375 GNDA.n1374 4.26717
R2450 GNDA.n1374 GNDA.n121 4.26717
R2451 GNDA.n1369 GNDA.n1368 4.26717
R2452 GNDA.n1368 GNDA.n1367 4.26717
R2453 GNDA.n1367 GNDA.n130 4.26717
R2454 GNDA.n1362 GNDA.n130 4.26717
R2455 GNDA.n1062 GNDA.n332 4.26717
R2456 GNDA.n334 GNDA.n332 4.26717
R2457 GNDA.n1055 GNDA.n334 4.26717
R2458 GNDA.n1055 GNDA.n1054 4.26717
R2459 GNDA.n1054 GNDA.n1053 4.26717
R2460 GNDA.n1053 GNDA.n344 4.26717
R2461 GNDA.n1048 GNDA.n1047 4.26717
R2462 GNDA.n1047 GNDA.n1046 4.26717
R2463 GNDA.n1046 GNDA.n353 4.26717
R2464 GNDA.n1041 GNDA.n353 4.26717
R2465 GNDA.n1242 GNDA.n1241 4.26717
R2466 GNDA.n1241 GNDA.n1220 4.26717
R2467 GNDA.n1236 GNDA.n1220 4.26717
R2468 GNDA.n1236 GNDA.n1235 4.26717
R2469 GNDA.n1235 GNDA.n1234 4.26717
R2470 GNDA.n1234 GNDA.n1 4.26717
R2471 GNDA.n1617 GNDA.n3 4.26717
R2472 GNDA.n1612 GNDA.n3 4.26717
R2473 GNDA.n1612 GNDA.n1611 4.26717
R2474 GNDA.n1611 GNDA.n1610 4.26717
R2475 GNDA.n783 GNDA.n583 4.1989
R2476 GNDA GNDA.n83 3.79309
R2477 GNDA.n1369 GNDA 3.79309
R2478 GNDA.n1048 GNDA 3.79309
R2479 GNDA GNDA.n1617 3.79309
R2480 GNDA.n1001 GNDA.n1000 3.70778
R2481 GNDA.n990 GNDA.n985 3.70778
R2482 GNDA.n1455 GNDA.n1453 3.5845
R2483 GNDA.n1454 GNDA.n105 3.5845
R2484 GNDA.n1462 GNDA.n1461 3.5845
R2485 GNDA.n103 GNDA.n102 3.5845
R2486 GNDA.n1470 GNDA.n1468 3.5845
R2487 GNDA.n1469 GNDA.n100 3.5845
R2488 GNDA.n1477 GNDA.n1476 3.5845
R2489 GNDA.n98 GNDA.n97 3.5845
R2490 GNDA.n1486 GNDA.n94 3.5845
R2491 GNDA.n872 GNDA.n761 3.5845
R2492 GNDA.n871 GNDA.n763 3.5845
R2493 GNDA.n794 GNDA.n792 3.5845
R2494 GNDA.n793 GNDA.n790 3.5845
R2495 GNDA.n801 GNDA.n800 3.5845
R2496 GNDA.n787 GNDA.n786 3.5845
R2497 GNDA.n809 GNDA.n807 3.5845
R2498 GNDA.n808 GNDA.n782 3.5845
R2499 GNDA.n816 GNDA.n815 3.5845
R2500 GNDA.n695 GNDA.n620 3.5845
R2501 GNDA.n699 GNDA.n696 3.5845
R2502 GNDA.n700 GNDA.n616 3.5845
R2503 GNDA.n705 GNDA.n704 3.5845
R2504 GNDA.n708 GNDA.n615 3.5845
R2505 GNDA.n712 GNDA.n709 3.5845
R2506 GNDA.n713 GNDA.n612 3.5845
R2507 GNDA.n718 GNDA.n717 3.5845
R2508 GNDA.n721 GNDA.n611 3.5845
R2509 GNDA.n499 GNDA.n388 3.5845
R2510 GNDA.n469 GNDA.n468 3.5845
R2511 GNDA.n475 GNDA.n471 3.5845
R2512 GNDA.n474 GNDA.n465 3.5845
R2513 GNDA.n481 GNDA.n464 3.5845
R2514 GNDA.n482 GNDA.n463 3.5845
R2515 GNDA.n487 GNDA.n485 3.5845
R2516 GNDA.n486 GNDA.n410 3.5845
R2517 GNDA.n494 GNDA.n493 3.5845
R2518 GNDA.n269 GNDA.n155 3.5845
R2519 GNDA.n236 GNDA.n235 3.5845
R2520 GNDA.n242 GNDA.n238 3.5845
R2521 GNDA.n241 GNDA.n232 3.5845
R2522 GNDA.n248 GNDA.n231 3.5845
R2523 GNDA.n249 GNDA.n230 3.5845
R2524 GNDA.n254 GNDA.n252 3.5845
R2525 GNDA.n253 GNDA.n177 3.5845
R2526 GNDA.n264 GNDA.n263 3.5845
R2527 GNDA.n1349 GNDA.n1070 3.5845
R2528 GNDA.n1348 GNDA.n1071 3.5845
R2529 GNDA.n1259 GNDA.n1258 3.5845
R2530 GNDA.n1272 GNDA.n1257 3.5845
R2531 GNDA.n1274 GNDA.n1273 3.5845
R2532 GNDA.n1281 GNDA.n1252 3.5845
R2533 GNDA.n1280 GNDA.n1254 3.5845
R2534 GNDA.n1253 GNDA.n1091 3.5845
R2535 GNDA.n1293 GNDA.n1292 3.5845
R2536 GNDA.n1210 GNDA.n1098 3.5845
R2537 GNDA.n1179 GNDA.n1178 3.5845
R2538 GNDA.n1185 GNDA.n1181 3.5845
R2539 GNDA.n1184 GNDA.n1175 3.5845
R2540 GNDA.n1191 GNDA.n1174 3.5845
R2541 GNDA.n1192 GNDA.n1173 3.5845
R2542 GNDA.n1197 GNDA.n1195 3.5845
R2543 GNDA.n1196 GNDA.n1120 3.5845
R2544 GNDA.n1205 GNDA.n1204 3.5845
R2545 GNDA.n571 GNDA.n563 3.4105
R2546 GNDA.n570 GNDA.n564 3.4105
R2547 GNDA.n569 GNDA.n568 3.4105
R2548 GNDA.n572 GNDA.n571 3.4105
R2549 GNDA.n570 GNDA.n562 3.4105
R2550 GNDA.n569 GNDA.n561 3.4105
R2551 GNDA.n1388 GNDA.n109 3.3797
R2552 GNDA.n1485 GNDA.n92 3.3797
R2553 GNDA.n784 GNDA.n783 3.3797
R2554 GNDA.n690 GNDA.n91 3.3797
R2555 GNDA.n723 GNDA.n722 3.3797
R2556 GNDA.n461 GNDA.n330 3.3797
R2557 GNDA.n259 GNDA.n228 3.3797
R2558 GNDA.n1356 GNDA.n1355 3.3797
R2559 GNDA.n1244 GNDA.n1092 3.3797
R2560 GNDA.n1243 GNDA.n1095 3.3797
R2561 GNDA.n1171 GNDA.n60 3.3797
R2562 GNDA.n934 GNDA.n91 3.27161
R2563 GNDA.n1357 GNDA.n1356 3.27161
R2564 GNDA.n1243 GNDA.n76 3.27161
R2565 GNDA.n1130 GNDA 3.02272
R2566 GNDA.n1335 GNDA 3.02272
R2567 GNDA.n420 GNDA 3.02272
R2568 GNDA.n677 GNDA 3.02272
R2569 GNDA.n1441 GNDA 3.02272
R2570 GNDA.n856 GNDA 3.02272
R2571 GNDA.n187 GNDA 3.02272
R2572 GNDA.n1389 GNDA.n107 2.8677
R2573 GNDA.n877 GNDA.n876 2.8677
R2574 GNDA.n692 GNDA.n691 2.8677
R2575 GNDA.n500 GNDA.n387 2.8677
R2576 GNDA.n270 GNDA.n154 2.8677
R2577 GNDA.n1069 GNDA.n1063 2.8677
R2578 GNDA.n1211 GNDA.n1097 2.8677
R2579 GNDA.n980 GNDA.n979 2.376
R2580 GNDA.n985 GNDA.n984 2.32777
R2581 GNDA.n1121 GNDA.n1097 2.31161
R2582 GNDA.n1343 GNDA.n1063 2.31161
R2583 GNDA.n411 GNDA.n387 2.31161
R2584 GNDA.n691 GNDA.n688 2.31161
R2585 GNDA.n1449 GNDA.n1389 2.31161
R2586 GNDA.n877 GNDA.n760 2.31161
R2587 GNDA.n178 GNDA.n154 2.31161
R2588 GNDA.n1000 GNDA.n971 2.04803
R2589 GNDA.n990 GNDA.n989 2.04803
R2590 GNDA.n1358 GNDA.n329 1.951
R2591 GNDA.n1216 GNDA.n1215 1.951
R2592 GNDA.n933 GNDA.n90 1.951
R2593 GNDA.n1385 GNDA.n110 1.951
R2594 GNDA.n881 GNDA.n880 1.951
R2595 GNDA.n505 GNDA.n504 1.951
R2596 GNDA.n275 GNDA.n274 1.951
R2597 GNDA.n1389 GNDA.n1388 1.7413
R2598 GNDA.n92 GNDA.n91 1.7413
R2599 GNDA.n878 GNDA.n877 1.7413
R2600 GNDA.n691 GNDA.n690 1.7413
R2601 GNDA.n387 GNDA.n381 1.7413
R2602 GNDA.n1356 GNDA.n330 1.7413
R2603 GNDA.n154 GNDA.n152 1.7413
R2604 GNDA.n259 GNDA.n109 1.7413
R2605 GNDA.n1355 GNDA.n1063 1.7413
R2606 GNDA.n1244 GNDA.n1243 1.7413
R2607 GNDA.n1097 GNDA.n1095 1.7413
R2608 GNDA.n1492 GNDA.n91 1.51754
R2609 GNDA.n111 GNDA.n109 1.51754
R2610 GNDA.n1356 GNDA.n1062 1.51754
R2611 GNDA.n1243 GNDA.n1242 1.51754
R2612 GNDA GNDA.n516 1.29343
R2613 GNDA.n286 GNDA 1.29343
R2614 GNDA.n1486 GNDA.n1485 1.2293
R2615 GNDA.n815 GNDA.n784 1.2293
R2616 GNDA.n722 GNDA.n721 1.2293
R2617 GNDA.n493 GNDA.n461 1.2293
R2618 GNDA.n263 GNDA.n228 1.2293
R2619 GNDA.n1292 GNDA.n1092 1.2293
R2620 GNDA.n1204 GNDA.n1171 1.2293
R2621 GNDA.n879 GNDA.n758 1.1781
R2622 GNDA.n507 GNDA.n506 1.1781
R2623 GNDA.n277 GNDA.n276 1.1781
R2624 GNDA.n1015 GNDA.n558 1.16414
R2625 GNDA.n1453 GNDA.n107 1.0245
R2626 GNDA.n1455 GNDA.n1454 1.0245
R2627 GNDA.n1462 GNDA.n105 1.0245
R2628 GNDA.n1461 GNDA.n103 1.0245
R2629 GNDA.n1468 GNDA.n102 1.0245
R2630 GNDA.n1470 GNDA.n1469 1.0245
R2631 GNDA.n1477 GNDA.n100 1.0245
R2632 GNDA.n1476 GNDA.n98 1.0245
R2633 GNDA.n97 GNDA.n94 1.0245
R2634 GNDA.n876 GNDA.n761 1.0245
R2635 GNDA.n872 GNDA.n871 1.0245
R2636 GNDA.n792 GNDA.n763 1.0245
R2637 GNDA.n794 GNDA.n793 1.0245
R2638 GNDA.n801 GNDA.n790 1.0245
R2639 GNDA.n800 GNDA.n787 1.0245
R2640 GNDA.n807 GNDA.n786 1.0245
R2641 GNDA.n809 GNDA.n808 1.0245
R2642 GNDA.n816 GNDA.n782 1.0245
R2643 GNDA.n692 GNDA.n620 1.0245
R2644 GNDA.n696 GNDA.n695 1.0245
R2645 GNDA.n700 GNDA.n699 1.0245
R2646 GNDA.n704 GNDA.n616 1.0245
R2647 GNDA.n705 GNDA.n615 1.0245
R2648 GNDA.n709 GNDA.n708 1.0245
R2649 GNDA.n713 GNDA.n712 1.0245
R2650 GNDA.n717 GNDA.n612 1.0245
R2651 GNDA.n718 GNDA.n611 1.0245
R2652 GNDA.n500 GNDA.n499 1.0245
R2653 GNDA.n468 GNDA.n388 1.0245
R2654 GNDA.n471 GNDA.n469 1.0245
R2655 GNDA.n475 GNDA.n474 1.0245
R2656 GNDA.n465 GNDA.n464 1.0245
R2657 GNDA.n482 GNDA.n481 1.0245
R2658 GNDA.n485 GNDA.n463 1.0245
R2659 GNDA.n487 GNDA.n486 1.0245
R2660 GNDA.n494 GNDA.n410 1.0245
R2661 GNDA.n270 GNDA.n269 1.0245
R2662 GNDA.n235 GNDA.n155 1.0245
R2663 GNDA.n238 GNDA.n236 1.0245
R2664 GNDA.n242 GNDA.n241 1.0245
R2665 GNDA.n232 GNDA.n231 1.0245
R2666 GNDA.n249 GNDA.n248 1.0245
R2667 GNDA.n252 GNDA.n230 1.0245
R2668 GNDA.n254 GNDA.n253 1.0245
R2669 GNDA.n264 GNDA.n177 1.0245
R2670 GNDA.n1070 GNDA.n1069 1.0245
R2671 GNDA.n1349 GNDA.n1348 1.0245
R2672 GNDA.n1258 GNDA.n1071 1.0245
R2673 GNDA.n1259 GNDA.n1257 1.0245
R2674 GNDA.n1274 GNDA.n1272 1.0245
R2675 GNDA.n1273 GNDA.n1252 1.0245
R2676 GNDA.n1281 GNDA.n1280 1.0245
R2677 GNDA.n1254 GNDA.n1253 1.0245
R2678 GNDA.n1293 GNDA.n1091 1.0245
R2679 GNDA.n1211 GNDA.n1210 1.0245
R2680 GNDA.n1178 GNDA.n1098 1.0245
R2681 GNDA.n1181 GNDA.n1179 1.0245
R2682 GNDA.n1185 GNDA.n1184 1.0245
R2683 GNDA.n1175 GNDA.n1174 1.0245
R2684 GNDA.n1192 GNDA.n1191 1.0245
R2685 GNDA.n1195 GNDA.n1173 1.0245
R2686 GNDA.n1197 GNDA.n1196 1.0245
R2687 GNDA.n1205 GNDA.n1120 1.0245
R2688 GNDA GNDA.n896 0.731929
R2689 GNDA.n1510 GNDA 0.474574
R2690 GNDA GNDA.n121 0.474574
R2691 GNDA GNDA.n344 0.474574
R2692 GNDA GNDA.n1 0.474574
R2693 GNDA GNDA.n574 0.417625
R2694 GNDA.n575 GNDA 0.264875
R2695 GNDA.n1006 GNDA.n575 0.170875
R2696 GNDA.n936 GNDA.n935 0.146786
R2697 GNDA.n981 GNDA.n978 0.1255
R2698 GNDA.n566 GNDA.n565 0.1255
R2699 GNDA.n567 GNDA.n566 0.1255
R2700 GNDA.n564 GNDA.n563 0.1255
R2701 GNDA.n568 GNDA.n564 0.1255
R2702 GNDA.n1529 GNDA.n75 0.0953148
R2703 GNDA.n1361 GNDA.n327 0.0953148
R2704 GNDA.n1040 GNDA.n552 0.0953148
R2705 GNDA.n38 GNDA.n10 0.0953148
R2706 GNDA.n981 GNDA.n980 0.0618108
R2707 GNDA.n571 GNDA.n570 0.0475
R2708 GNDA.n570 GNDA.n569 0.0475
R2709 GNDA.n572 GNDA.n562 0.0475
R2710 GNDA.n562 GNDA.n561 0.0475
R2711 a_4938_4530.t0 a_4938_4530.t1 483.048
R2712 V_TOP.n18 V_TOP.t13 750.967
R2713 V_TOP.n7 V_TOP.t18 404.88
R2714 V_TOP.n2 V_TOP.n0 276.313
R2715 V_TOP.n2 V_TOP.n1 272.688
R2716 V_TOP.n5 V_TOP.n3 268.188
R2717 V_TOP.n8 V_TOP.n7 244.214
R2718 V_TOP.n9 V_TOP.n8 244.214
R2719 V_TOP.n10 V_TOP.n9 244.214
R2720 V_TOP.n11 V_TOP.n10 244.214
R2721 V_TOP.n12 V_TOP.n11 244.214
R2722 V_TOP.n13 V_TOP.n12 244.214
R2723 V_TOP.n14 V_TOP.n13 244.214
R2724 V_TOP.n15 V_TOP.n14 244.214
R2725 V_TOP.n16 V_TOP.n15 244.214
R2726 V_TOP.n17 V_TOP.n16 224.052
R2727 V_TOP.t3 V_TOP.n19 221.411
R2728 V_TOP.n18 V_TOP.n17 181.601
R2729 V_TOP.n4 V_TOP.t7 161.034
R2730 V_TOP.n7 V_TOP.t12 160.667
R2731 V_TOP.n8 V_TOP.t19 160.667
R2732 V_TOP.n9 V_TOP.t14 160.667
R2733 V_TOP.n10 V_TOP.t9 160.667
R2734 V_TOP.n11 V_TOP.t16 160.667
R2735 V_TOP.n12 V_TOP.t10 160.667
R2736 V_TOP.n13 V_TOP.t17 160.667
R2737 V_TOP.n14 V_TOP.t11 160.667
R2738 V_TOP.n15 V_TOP.t20 160.667
R2739 V_TOP.n16 V_TOP.t15 160.667
R2740 V_TOP.n17 V_TOP.t21 160.667
R2741 V_TOP.n4 V_TOP.t6 109.861
R2742 V_TOP.n19 V_TOP.n18 84.24
R2743 V_TOP.n19 V_TOP.n6 61.4838
R2744 V_TOP.n5 V_TOP.n4 21.4255
R2745 V_TOP.n3 V_TOP.t4 19.7005
R2746 V_TOP.n3 V_TOP.t8 19.7005
R2747 V_TOP.n1 V_TOP.t5 19.7005
R2748 V_TOP.n1 V_TOP.t2 19.7005
R2749 V_TOP.n0 V_TOP.t1 19.7005
R2750 V_TOP.n0 V_TOP.t0 19.7005
R2751 V_TOP.n6 V_TOP.n5 4.5005
R2752 V_TOP.n6 V_TOP.n2 3.6255
R2753 Vin-.n8 Vin-.t1 460.144
R2754 Vin-.n13 Vin-.t8 205.968
R2755 Vin-.n8 Vin-.t9 205.968
R2756 Vin-.n11 Vin-.n10 205.946
R2757 Vin-.n15 Vin-.t0 175.276
R2758 Vin-.n10 Vin-.n9 165.8
R2759 Vin-.n12 Vin-.n11 165.8
R2760 Vin-.n7 Vin-.n5 156.615
R2761 Vin-.n7 Vin-.n6 154.24
R2762 Vin-.n1 Vin-.n0 83.5719
R2763 Vin-.n22 Vin-.n21 83.5719
R2764 Vin-.n20 Vin-.n19 83.5719
R2765 Vin-.n25 Vin-.n1 73.682
R2766 Vin-.n20 Vin-.n4 73.3165
R2767 Vin-.n11 Vin-.t7 40.1672
R2768 Vin-.n10 Vin-.t10 40.1672
R2769 Vin-.n21 Vin-.n20 26.074
R2770 Vin-.t2 Vin-.n1 25.7843
R2771 Vin-.n16 Vin-.n15 15.4
R2772 Vin-.n14 Vin-.n7 12.6255
R2773 Vin-.n6 Vin-.t6 9.8505
R2774 Vin-.n6 Vin-.t5 9.8505
R2775 Vin-.n5 Vin-.t4 9.8505
R2776 Vin-.n5 Vin-.t3 9.8505
R2777 Vin-.n14 Vin-.n13 7.59425
R2778 Vin-.n16 Vin-.n4 2.19742
R2779 Vin-.n9 Vin-.n8 1.7505
R2780 Vin-.n13 Vin-.n12 1.7505
R2781 Vin-.n24 Vin-.n23 1.5505
R2782 Vin-.n3 Vin-.n2 1.5505
R2783 Vin-.n18 Vin-.n17 1.5505
R2784 Vin-.n15 Vin-.n14 1.53175
R2785 Vin-.n18 Vin-.n4 1.19225
R2786 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6.Emitter Vin-.n25 1.07742
R2787 Vin-.n23 Vin-.n22 1.07024
R2788 Vin-.n19 Vin-.n18 0.959578
R2789 Vin-.n19 Vin-.n3 0.885803
R2790 Vin-.n22 Vin-.n3 0.77514
R2791 Vin-.n25 Vin-.n24 0.763532
R2792 Vin-.n23 Vin-.n0 0.590702
R2793 Vin-.n12 Vin-.n9 0.5005
R2794 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6.Emitter Vin-.n0 0.498483
R2795 Vin-.n21 Vin-.t2 0.290206
R2796 Vin-.n17 Vin-.n16 0.0183571
R2797 Vin-.n17 Vin-.n2 0.0183571
R2798 Vin-.n24 Vin-.n2 0.0183571
R2799 VDDA.n51 VDDA.n35 587.407
R2800 VDDA.n45 VDDA.n39 587.407
R2801 VDDA.n80 VDDA.n4 587.407
R2802 VDDA.n84 VDDA.n83 587.407
R2803 VDDA.n92 VDDA.n80 585
R2804 VDDA.n91 VDDA.n81 585
R2805 VDDA.n90 VDDA.n82 585
R2806 VDDA.n87 VDDA.n83 585
R2807 VDDA.n49 VDDA.n35 585
R2808 VDDA.n48 VDDA.n47 585
R2809 VDDA.n46 VDDA.n38 585
R2810 VDDA.n45 VDDA.n44 585
R2811 VDDA.t30 VDDA.n11 464.281
R2812 VDDA.n17 VDDA.t30 464.281
R2813 VDDA.n75 VDDA.t25 464.281
R2814 VDDA.t25 VDDA.n74 464.281
R2815 VDDA.n97 VDDA.t31 328.668
R2816 VDDA.n34 VDDA.t26 328.668
R2817 VDDA.n0 VDDA.t43 298.221
R2818 VDDA.n70 VDDA.t23 248.333
R2819 VDDA.n57 VDDA.t29 248.333
R2820 VDDA.n47 VDDA.n35 246.25
R2821 VDDA.n46 VDDA.n45 246.25
R2822 VDDA.n81 VDDA.n80 246.25
R2823 VDDA.n83 VDDA.n82 246.25
R2824 VDDA.n74 VDDA.n9 243.698
R2825 VDDA.n21 VDDA.n17 243.698
R2826 VDDA.n96 VDDA.n95 238.367
R2827 VDDA.n77 VDDA.n76 238.367
R2828 VDDA.n56 VDDA.n55 238.367
R2829 VDDA.n59 VDDA.n58 205.488
R2830 VDDA.n61 VDDA.n60 205.488
R2831 VDDA.n63 VDDA.n62 205.488
R2832 VDDA.n65 VDDA.n64 205.488
R2833 VDDA.n67 VDDA.n66 205.488
R2834 VDDA.n69 VDDA.n68 205.488
R2835 VDDA.n84 VDDA.n8 190.333
R2836 VDDA.n39 VDDA.n16 190.333
R2837 VDDA.n18 VDDA.n12 185
R2838 VDDA.n20 VDDA.n19 185
R2839 VDDA.n71 VDDA.n10 185
R2840 VDDA.n73 VDDA.n72 185
R2841 VDDA.n79 VDDA.n5 185
R2842 VDDA.n93 VDDA.n92 185
R2843 VDDA.n94 VDDA.n93 185
R2844 VDDA.n91 VDDA.n78 185
R2845 VDDA.n90 VDDA.n89 185
R2846 VDDA.n88 VDDA.n87 185
R2847 VDDA.n86 VDDA.n85 185
R2848 VDDA.n94 VDDA.n8 185
R2849 VDDA.n53 VDDA.n52 185
R2850 VDDA.n54 VDDA.n53 185
R2851 VDDA.n50 VDDA.n22 185
R2852 VDDA.n49 VDDA.n36 185
R2853 VDDA.n48 VDDA.n37 185
R2854 VDDA.n40 VDDA.n38 185
R2855 VDDA.n44 VDDA.n41 185
R2856 VDDA.n43 VDDA.n42 185
R2857 VDDA.n54 VDDA.n16 185
R2858 VDDA.n3 VDDA.n2 154.242
R2859 VDDA.n24 VDDA.n23 154.242
R2860 VDDA.n26 VDDA.n25 154.242
R2861 VDDA.n28 VDDA.n27 154.242
R2862 VDDA.n30 VDDA.n29 154.242
R2863 VDDA.n32 VDDA.n31 154.242
R2864 VDDA.n93 VDDA.n5 150
R2865 VDDA.n93 VDDA.n78 150
R2866 VDDA.n89 VDDA.n88 150
R2867 VDDA.n85 VDDA.n8 150
R2868 VDDA.n72 VDDA.n10 150
R2869 VDDA.n20 VDDA.n12 150
R2870 VDDA.n53 VDDA.n22 150
R2871 VDDA.n37 VDDA.n36 150
R2872 VDDA.n41 VDDA.n40 150
R2873 VDDA.n42 VDDA.n16 150
R2874 VDDA.t16 VDDA.t42 138.082
R2875 VDDA.n47 VDDA.t28 123.126
R2876 VDDA.t28 VDDA.n46 123.126
R2877 VDDA.t32 VDDA.n81 123.126
R2878 VDDA.n82 VDDA.t32 123.126
R2879 VDDA.t27 VDDA.t33 110.466
R2880 VDDA.t33 VDDA.t2 110.466
R2881 VDDA.t2 VDDA.t10 110.466
R2882 VDDA.t10 VDDA.t8 110.466
R2883 VDDA.t8 VDDA.t6 110.466
R2884 VDDA.t6 VDDA.t21 110.466
R2885 VDDA.t21 VDDA.t14 110.466
R2886 VDDA.t14 VDDA.t17 110.466
R2887 VDDA.t17 VDDA.t0 110.466
R2888 VDDA.t0 VDDA.t4 110.466
R2889 VDDA.t4 VDDA.t19 110.466
R2890 VDDA.t19 VDDA.t12 110.466
R2891 VDDA.t12 VDDA.t24 110.466
R2892 VDDA.n54 VDDA.t16 107.704
R2893 VDDA.n54 VDDA.t27 99.4191
R2894 VDDA.n94 VDDA.t24 99.4191
R2895 VDDA.n55 VDDA.n54 65.8183
R2896 VDDA.n54 VDDA.n21 65.8183
R2897 VDDA.n94 VDDA.n77 65.8183
R2898 VDDA.n94 VDDA.n9 65.8183
R2899 VDDA.n95 VDDA.n94 65.8183
R2900 VDDA.n94 VDDA.n6 65.8183
R2901 VDDA.n94 VDDA.n7 65.8183
R2902 VDDA.n54 VDDA.n13 65.8183
R2903 VDDA.n54 VDDA.n14 65.8183
R2904 VDDA.n54 VDDA.n15 65.8183
R2905 VDDA.n78 VDDA.n6 53.3664
R2906 VDDA.n88 VDDA.n7 53.3664
R2907 VDDA.n72 VDDA.n9 53.3664
R2908 VDDA.n21 VDDA.n20 53.3664
R2909 VDDA.n55 VDDA.n12 53.3664
R2910 VDDA.n77 VDDA.n10 53.3664
R2911 VDDA.n95 VDDA.n5 53.3664
R2912 VDDA.n89 VDDA.n6 53.3664
R2913 VDDA.n85 VDDA.n7 53.3664
R2914 VDDA.n22 VDDA.n13 53.3664
R2915 VDDA.n37 VDDA.n14 53.3664
R2916 VDDA.n41 VDDA.n15 53.3664
R2917 VDDA.n36 VDDA.n13 53.3664
R2918 VDDA.n40 VDDA.n14 53.3664
R2919 VDDA.n42 VDDA.n15 53.3664
R2920 VDDA.n99 VDDA.n98 23.3792
R2921 VDDA.n58 VDDA.t48 19.7005
R2922 VDDA.n58 VDDA.t3 19.7005
R2923 VDDA.n60 VDDA.t11 19.7005
R2924 VDDA.n60 VDDA.t9 19.7005
R2925 VDDA.n62 VDDA.t7 19.7005
R2926 VDDA.n62 VDDA.t22 19.7005
R2927 VDDA.n64 VDDA.t15 19.7005
R2928 VDDA.n64 VDDA.t18 19.7005
R2929 VDDA.n66 VDDA.t1 19.7005
R2930 VDDA.n66 VDDA.t5 19.7005
R2931 VDDA.n68 VDDA.t20 19.7005
R2932 VDDA.n68 VDDA.t13 19.7005
R2933 VDDA.n97 VDDA.n96 16.4576
R2934 VDDA.n76 VDDA.n70 16.4576
R2935 VDDA.n57 VDDA.n56 16.4576
R2936 VDDA.n52 VDDA.n34 16.4576
R2937 VDDA VDDA.n99 15.2934
R2938 VDDA.n70 VDDA.n69 14.9255
R2939 VDDA.n59 VDDA.n57 14.9255
R2940 VDDA.n34 VDDA.n33 13.8005
R2941 VDDA.n98 VDDA.n97 13.8005
R2942 VDDA.n99 VDDA.n1 11.8918
R2943 VDDA.n2 VDDA.t44 9.8505
R2944 VDDA.n2 VDDA.t37 9.8505
R2945 VDDA.n23 VDDA.t41 9.8505
R2946 VDDA.n23 VDDA.t36 9.8505
R2947 VDDA.n25 VDDA.t39 9.8505
R2948 VDDA.n25 VDDA.t47 9.8505
R2949 VDDA.n27 VDDA.t38 9.8505
R2950 VDDA.n27 VDDA.t46 9.8505
R2951 VDDA.n29 VDDA.t35 9.8505
R2952 VDDA.n29 VDDA.t45 9.8505
R2953 VDDA.n31 VDDA.t34 9.8505
R2954 VDDA.n31 VDDA.t40 9.8505
R2955 VDDA.n92 VDDA.n79 9.14336
R2956 VDDA.n92 VDDA.n91 9.14336
R2957 VDDA.n91 VDDA.n90 9.14336
R2958 VDDA.n90 VDDA.n87 9.14336
R2959 VDDA.n87 VDDA.n86 9.14336
R2960 VDDA.n73 VDDA.n71 9.14336
R2961 VDDA.n19 VDDA.n18 9.14336
R2962 VDDA.n50 VDDA.n49 9.14336
R2963 VDDA.n49 VDDA.n48 9.14336
R2964 VDDA.n48 VDDA.n38 9.14336
R2965 VDDA.n44 VDDA.n38 9.14336
R2966 VDDA.n44 VDDA.n43 9.14336
R2967 VDDA.n33 VDDA.n1 6.12925
R2968 VDDA.n52 VDDA.n51 5.33286
R2969 VDDA.n96 VDDA.n4 5.33286
R2970 VDDA.n76 VDDA.n75 5.33286
R2971 VDDA.n56 VDDA.n11 5.33286
R2972 VDDA.n79 VDDA.n4 3.75335
R2973 VDDA.n86 VDDA.n84 3.75335
R2974 VDDA.n75 VDDA.n71 3.75335
R2975 VDDA.n74 VDDA.n73 3.75335
R2976 VDDA.n18 VDDA.n11 3.75335
R2977 VDDA.n19 VDDA.n17 3.75335
R2978 VDDA.n51 VDDA.n50 3.75335
R2979 VDDA.n43 VDDA.n39 3.75335
R2980 VDDA.n69 VDDA.n67 1.1255
R2981 VDDA.n67 VDDA.n65 1.1255
R2982 VDDA.n65 VDDA.n63 1.1255
R2983 VDDA.n63 VDDA.n61 1.1255
R2984 VDDA.n61 VDDA.n59 1.1255
R2985 VDDA.n33 VDDA.n32 1.1255
R2986 VDDA.n32 VDDA.n30 1.1255
R2987 VDDA.n30 VDDA.n28 1.1255
R2988 VDDA.n28 VDDA.n26 1.1255
R2989 VDDA.n26 VDDA.n24 1.1255
R2990 VDDA.n24 VDDA.n3 1.1255
R2991 VDDA.n98 VDDA.n3 1.1255
R2992 VDDA VDDA.n0 0.958125
R2993 VDDA.n1 VDDA.n0 0.729
R2994 V_OUT.n3 V_OUT.n0 215.465
R2995 V_OUT.n2 V_OUT.n1 211.84
R2996 V_OUT.n2 V_OUT.t0 174.102
R2997 V_OUT.n5 V_OUT.n3 160.59
R2998 V_OUT V_OUT.n5 100.555
R2999 V_OUT.n5 V_OUT.n4 51.2504
R3000 V_OUT.n4 V_OUT.t6 9.8505
R3001 V_OUT.n4 V_OUT.t5 9.8505
R3002 V_OUT.n1 V_OUT.t4 9.8505
R3003 V_OUT.n1 V_OUT.t2 9.8505
R3004 V_OUT.n0 V_OUT.t1 9.8505
R3005 V_OUT.n0 V_OUT.t3 9.8505
R3006 V_OUT.n3 V_OUT.n2 3.6255
R3007 V_mirror.n9 V_mirror.t16 324.548
R3008 V_mirror.n4 V_mirror.t15 324.548
R3009 V_mirror.n10 V_mirror.n9 244.214
R3010 V_mirror.n5 V_mirror.n4 244.214
R3011 V_mirror.n2 V_mirror.n0 195.852
R3012 V_mirror.n7 V_mirror.n3 194.888
R3013 V_mirror.n12 V_mirror.n8 194.888
R3014 V_mirror.n2 V_mirror.n1 193.477
R3015 V_mirror.n15 V_mirror.n14 188.977
R3016 V_mirror.n11 V_mirror.t6 157.453
R3017 V_mirror.n6 V_mirror.t4 157.453
R3018 V_mirror.n7 V_mirror.n6 152
R3019 V_mirror.n12 V_mirror.n11 152
R3020 V_mirror.n9 V_mirror.t14 80.3338
R3021 V_mirror.n10 V_mirror.t2 80.3338
R3022 V_mirror.n4 V_mirror.t17 80.3338
R3023 V_mirror.n5 V_mirror.t0 80.3338
R3024 V_mirror.n11 V_mirror.n10 77.1205
R3025 V_mirror.n6 V_mirror.n5 77.1205
R3026 V_mirror.n1 V_mirror.t13 24.0005
R3027 V_mirror.n1 V_mirror.t11 24.0005
R3028 V_mirror.n0 V_mirror.t9 24.0005
R3029 V_mirror.n0 V_mirror.t10 24.0005
R3030 V_mirror.n14 V_mirror.t12 24.0005
R3031 V_mirror.n14 V_mirror.t8 24.0005
R3032 V_mirror.n13 V_mirror.n7 23.1755
R3033 V_mirror.n3 V_mirror.t5 19.7005
R3034 V_mirror.n3 V_mirror.t1 19.7005
R3035 V_mirror.n8 V_mirror.t3 19.7005
R3036 V_mirror.n8 V_mirror.t7 19.7005
R3037 V_mirror.n13 V_mirror.n12 9.3005
R3038 V_mirror V_mirror.n15 4.5005
R3039 V_mirror V_mirror.n2 2.3755
R3040 V_mirror.n15 V_mirror.n13 0.8755
R3041 a_4938_4770.t0 a_4938_4770.t1 258.591
R3042 1st_Vout.n8 1st_Vout.t9 419.377
R3043 1st_Vout.n7 1st_Vout.t10 419.377
R3044 1st_Vout.n1 1st_Vout.n0 100.352
R3045 1st_Vout.n9 1st_Vout.n8 237.488
R3046 1st_Vout.n6 1st_Vout.n2 232.988
R3047 1st_Vout.n5 1st_Vout.n4 171.553
R3048 1st_Vout.n5 1st_Vout.n3 160.178
R3049 1st_Vout.n1 1st_Vout.t11 165.934
R3050 1st_Vout.n1 1st_Vout.t8 165.934
R3051 1st_Vout.n4 1st_Vout.t4 24.0005
R3052 1st_Vout.n4 1st_Vout.t6 24.0005
R3053 1st_Vout.n3 1st_Vout.t7 24.0005
R3054 1st_Vout.n3 1st_Vout.t5 24.0005
R3055 1st_Vout.n2 1st_Vout.t0 19.7005
R3056 1st_Vout.n2 1st_Vout.t2 19.7005
R3057 1st_Vout.n9 1st_Vout.t1 19.7005
R3058 1st_Vout.t3 1st_Vout.n9 19.7005
R3059 1st_Vout.n7 1st_Vout.n6 4.5005
R3060 1st_Vout.n8 1st_Vout.n0 1.313
R3061 1st_Vout.n6 1st_Vout.n5 0.8755
R3062 1st_Vout.n0 1st_Vout.n7 0.813
R3063 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t0 158.431
R3064 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n15 83.5719
R3065 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n12 83.5719
R3066 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n21 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n11 83.5719
R3067 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n29 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n28 83.5719
R3068 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n9 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n7 83.5719
R3069 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n34 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n6 83.5719
R3070 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n48 83.5719
R3071 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n45 83.5719
R3072 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n44 83.5719
R3073 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n61 83.5719
R3074 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n40 83.5719
R3075 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n39 83.5719
R3076 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n84 83.5719
R3077 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n85 83.5719
R3078 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n88 83.5719
R3079 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n0 83.5719
R3080 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n79 83.5719
R3081 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n76 83.5719
R3082 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n13 73.682
R3083 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n46 73.682
R3084 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n86 73.682
R3085 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n23 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n11 73.3165
R3086 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n36 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n6 73.3165
R3087 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n44 73.3165
R3088 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n39 73.3165
R3089 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n84 73.3165
R3090 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n4 73.3165
R3091 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n28 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n27 73.19
R3092 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n60 73.19
R3093 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n1 73.19
R3094 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n11 26.074
R3095 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n9 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n6 26.074
R3096 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n44 26.074
R3097 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n39 26.074
R3098 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n84 26.074
R3099 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n77 26.074
R3100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t1 25.7843
R3101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n28 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t4 25.7843
R3102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t5 25.7843
R3103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t2 25.7843
R3104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t6 25.7843
R3105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n78 25.7843
R3106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n27 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n25 2.36206
R3107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n58 2.36206
R3108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n1 2.36206
R3109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n24 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n23 2.19742
R3110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n37 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n36 2.19742
R3111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n56 2.19742
R3112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n69 2.19742
R3113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n96 2.19742
R3114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n4 2.19742
R3115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n26 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n8 1.5505
R3116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n31 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n30 1.5505
R3117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n33 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n32 1.5505
R3118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n35 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n5 1.5505
R3119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n18 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n17 1.5505
R3120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n20 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n19 1.5505
R3121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n10 1.5505
R3122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n41 1.5505
R3123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n63 1.5505
R3124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n65 1.5505
R3125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n38 1.5505
R3126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n50 1.5505
R3127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n52 1.5505
R3128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n43 1.5505
R3129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n99 1.5505
R3130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n81 1.5505
R3131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n2 1.5505
R3132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n74 1.5505
R3133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n90 1.5505
R3134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n92 1.5505
R3135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n83 1.5505
R3136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n37 1.26871
R3137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n23 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n22 1.19225
R3138 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n36 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n35 1.19225
R3139 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n55 1.19225
R3140 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n68 1.19225
R3141 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n95 1.19225
R3142 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n4 1.19225
R3143 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n13 1.07742
R3144 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n46 1.07742
R3145 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n86 1.07742
R3146 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n17 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n12 1.07024
R3147 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n30 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n7 1.07024
R3148 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n45 1.07024
R3149 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n40 1.07024
R3150 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n85 1.07024
R3151 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n80 1.07024
R3152 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n27 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n26 1.0237
R3153 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n59 1.0237
R3154 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n1 1.0237
R3155 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n21 0.959578
R3156 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n35 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n34 0.959578
R3157 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n54 0.959578
R3158 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n67 0.959578
R3159 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n94 0.959578
R3160 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n75 0.959578
R3161 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n21 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n20 0.885803
R3162 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n34 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n33 0.885803
R3163 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n53 0.885803
R3164 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n66 0.885803
R3165 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n93 0.885803
R3166 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n3 0.885803
R3167 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n20 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n12 0.77514
R3168 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n33 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n7 0.77514
R3169 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n45 0.77514
R3170 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n40 0.77514
R3171 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n85 0.77514
R3172 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n3 0.77514
R3173 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n18 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n13 0.763532
R3174 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n46 0.763532
R3175 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n86 0.763532
R3176 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n26 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.756696
R3177 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.756696
R3178 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n100 0.756696
R3179 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n17 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n16 0.590702
R3180 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n30 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n29 0.590702
R3181 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n49 0.590702
R3182 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n62 0.590702
R3183 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n89 0.590702
R3184 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n0 0.590702
R3185 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n72 0.590143
R3186 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n71 0.554071
R3187 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.498483
R3188 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n29 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.498483
R3189 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.498483
R3190 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.498483
R3191 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.498483
R3192 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n0 0.498483
R3193 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n14 0.290206
R3194 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n9 0.290206
R3195 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t5 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n47 0.290206
R3196 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n42 0.290206
R3197 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t6 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n87 0.290206
R3198 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.t3 0.290206
R3199 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n25 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n24 0.154071
R3200 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n57 0.154071
R3201 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n97 0.154071
R3202 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n70 0.0901429
R3203 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n37 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n5 0.0183571
R3204 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n32 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n5 0.0183571
R3205 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n32 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n31 0.0183571
R3206 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n31 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n8 0.0183571
R3207 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n25 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n8 0.0183571
R3208 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n24 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n10 0.0183571
R3209 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n19 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n10 0.0183571
R3210 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n19 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n18 0.0183571
R3211 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n38 0.0183571
R3212 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n38 0.0183571
R3213 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n64 0.0183571
R3214 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n41 0.0183571
R3215 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n41 0.0183571
R3216 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n43 0.0183571
R3217 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n43 0.0183571
R3218 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n51 0.0183571
R3219 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n73 0.0183571
R3220 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n2 0.0183571
R3221 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n2 0.0183571
R3222 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n82 0.0183571
R3223 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n98 0.0183571
R3224 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n83 0.0183571
R3225 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n83 0.0183571
R3226 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter.n91 0.0183571
R3227 start_up.n1 start_up.t3 776.592
R3228 start_up.t2 start_up.n2 500.086
R3229 start_up.t2 start_up.n2 461.389
R3230 start_up.n0 start_up.t1 268.95
R3231 start_up.n1 start_up.n0 148.969
R3232 start_up.n2 start_up.n1 49.6698
R3233 start_up.n0 start_up.t0 14.4499
R3234 Vin+.n2 Vin+.n0 187.791
R3235 Vin+.n2 Vin+.n1 183.041
R3236 Vin+.t0 Vin+.n7 177.677
R3237 Vin+.n6 Vin+.n4 168.175
R3238 Vin+.n6 Vin+.n5 165.8
R3239 Vin+.n3 Vin+.t1 159.726
R3240 Vin+.n5 Vin+.t9 119.43
R3241 Vin+.n5 Vin+.t7 119.43
R3242 Vin+.n4 Vin+.t6 119.43
R3243 Vin+.n4 Vin+.t8 119.43
R3244 Vin+.n1 Vin+.t3 9.8505
R3245 Vin+.n1 Vin+.t5 9.8505
R3246 Vin+.n0 Vin+.t4 9.8505
R3247 Vin+.n0 Vin+.t2 9.8505
R3248 Vin+.n3 Vin+.n2 8.6255
R3249 Vin+.n7 Vin+.n6 8.188
R3250 Vin+.n7 Vin+.n3 3.09425
R3251 V_p.n11 V_p.t9 196.089
R3252 V_p.n1 V_p.n5 169.001
R3253 V_p.n1 V_p.n6 167.876
R3254 V_p.n0 V_p.n2 154.077
R3255 V_p.n7 V_p.n4 154.077
R3256 V_p.n10 V_p.n3 152
R3257 V_p.n11 V_p.n10 89.2066
R3258 V_p.n9 V_p.n8 68.85
R3259 V_p.n8 V_p.n7 45.1025
R3260 V_p.n8 V_p.n3 26.8309
R3261 V_p.n9 V_p.t8 24.1005
R3262 V_p.n2 V_p.t0 24.0005
R3263 V_p.n2 V_p.t6 24.0005
R3264 V_p.n4 V_p.t7 24.0005
R3265 V_p.n4 V_p.t2 24.0005
R3266 V_p.n5 V_p.t5 24.0005
R3267 V_p.n5 V_p.t1 24.0005
R3268 V_p.n6 V_p.t3 24.0005
R3269 V_p.n6 V_p.t4 24.0005
R3270 V_p.n12 V_p.n11 19.0351
R3271 V_p.n10 V_p.n9 17.5278
R3272 V_p.n1 V_p.n0 14.9255
R3273 V_p.n7 V_p.n1 14.9255
R3274 V_p V_p.n0 12.8005
R3275 V_p.n12 V_p.n3 6.4005
R3276 V_p V_p.n12 6.4005
R3277 a_4938_3210.t0 a_4938_3210.t1 258.591
R3278 a_4938_2970.t0 a_4938_2970.t1 483.048
R3279 a_3410_3330.t0 a_3410_3330.t1 483.048
R3280 a_3410_3450.t0 a_3410_3450.t1 376.99
R3281 a_4938_3810.t0 a_4938_3810.t1 415.39
R3282 a_4938_3090.t0 a_4938_3090.t1 376.99
R3283 a_4938_3930.t0 a_4938_3930.t1 280.534
R3284 a_3410_3570.t0 a_3410_3570.t1 258.591
R3285 a_4938_3690.t0 a_4938_3690.t1 521.448
R3286 a_3410_4410.t0 a_3410_4410.t1 258.591
R3287 a_3410_4170.t0 a_3410_4170.t1 483.048
R3288 a_3410_4290.t0 a_3410_4290.t1 376.99
R3289 a_4938_4650.t0 a_4938_4650.t1 376.99
C0 VDDA V_OUT 2.78133f
C1 V_mirror V_p 0.138864f
C2 VDDA V_p 0.027153f
C3 VDDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter 0.069333f
C4 VDDA V_mirror 1.72554f
C5 V_OUT GNDA 1.826189f
C6 VDDA GNDA 44.76623f
C7 V_p GNDA 2.34007f
C8 V_mirror GNDA 1.89738f
C9 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5.Emitter GNDA 11.8561f
C10 Vin+.t4 GNDA 0.064698f
C11 Vin+.t2 GNDA 0.064698f
C12 Vin+.n0 GNDA 0.257812f
C13 Vin+.t3 GNDA 0.064698f
C14 Vin+.t5 GNDA 0.064698f
C15 Vin+.n1 GNDA 0.250566f
C16 Vin+.n2 GNDA 0.70129f
C17 Vin+.t1 GNDA 0.159367f
C18 Vin+.n3 GNDA 0.567461f
C19 Vin+.t8 GNDA 0.0888f
C20 Vin+.t6 GNDA 0.0888f
C21 Vin+.n4 GNDA 0.069752f
C22 Vin+.t7 GNDA 0.0888f
C23 Vin+.t9 GNDA 0.0888f
C24 Vin+.n5 GNDA 0.067874f
C25 Vin+.n6 GNDA 0.421232f
C26 Vin+.n7 GNDA 0.97459f
C27 Vin+.t0 GNDA 0.216063f
C28 V_OUT.t1 GNDA 0.099964f
C29 V_OUT.t3 GNDA 0.099964f
C30 V_OUT.n0 GNDA 0.416226f
C31 V_OUT.t0 GNDA 0.357326f
C32 V_OUT.t4 GNDA 0.099964f
C33 V_OUT.t2 GNDA 0.099964f
C34 V_OUT.n1 GNDA 0.409535f
C35 V_OUT.n2 GNDA 1.82908f
C36 V_OUT.n3 GNDA 0.861714f
C37 V_OUT.t6 GNDA 0.099964f
C38 V_OUT.t5 GNDA 0.099964f
C39 V_OUT.n4 GNDA 0.199928f
C40 V_OUT.n5 GNDA 0.22287f
C41 VDDA.t43 GNDA 0.018318f
C42 VDDA.n0 GNDA 0.107843f
C43 VDDA.n1 GNDA 0.355239f
C44 VDDA.n2 GNDA 0.034575f
C45 VDDA.n3 GNDA 0.032759f
C46 VDDA.t31 GNDA 0.051643f
C47 VDDA.t24 GNDA 0.19577f
C48 VDDA.t23 GNDA 0.028665f
C49 VDDA.t29 GNDA 0.028603f
C50 VDDA.t42 GNDA 0.267896f
C51 VDDA.t16 GNDA 0.229257f
C52 VDDA.t12 GNDA 0.206074f
C53 VDDA.t19 GNDA 0.206074f
C54 VDDA.t4 GNDA 0.206074f
C55 VDDA.t0 GNDA 0.206074f
C56 VDDA.t17 GNDA 0.206074f
C57 VDDA.t14 GNDA 0.206074f
C58 VDDA.t21 GNDA 0.206074f
C59 VDDA.t6 GNDA 0.206074f
C60 VDDA.t8 GNDA 0.206074f
C61 VDDA.t10 GNDA 0.206074f
C62 VDDA.t2 GNDA 0.206074f
C63 VDDA.t33 GNDA 0.206074f
C64 VDDA.t27 GNDA 0.19577f
C65 VDDA.t30 GNDA 0.012635f
C66 VDDA.n17 GNDA 0.011669f
C67 VDDA.t26 GNDA 0.051643f
C68 VDDA.n23 GNDA 0.034575f
C69 VDDA.n24 GNDA 0.032759f
C70 VDDA.n25 GNDA 0.034575f
C71 VDDA.n26 GNDA 0.032759f
C72 VDDA.n27 GNDA 0.034575f
C73 VDDA.n28 GNDA 0.032759f
C74 VDDA.n29 GNDA 0.034575f
C75 VDDA.n30 GNDA 0.032759f
C76 VDDA.n31 GNDA 0.034575f
C77 VDDA.n32 GNDA 0.032759f
C78 VDDA.n33 GNDA 0.027862f
C79 VDDA.n34 GNDA 0.021493f
C80 VDDA.n39 GNDA 0.01214f
C81 VDDA.n54 GNDA 0.193194f
C82 VDDA.n56 GNDA 0.010041f
C83 VDDA.n57 GNDA 0.015593f
C84 VDDA.n58 GNDA 0.013997f
C85 VDDA.n59 GNDA 0.038853f
C86 VDDA.n60 GNDA 0.013997f
C87 VDDA.n61 GNDA 0.029375f
C88 VDDA.n62 GNDA 0.013997f
C89 VDDA.n63 GNDA 0.029375f
C90 VDDA.n64 GNDA 0.013997f
C91 VDDA.n65 GNDA 0.029375f
C92 VDDA.n66 GNDA 0.013997f
C93 VDDA.n67 GNDA 0.029375f
C94 VDDA.n68 GNDA 0.013997f
C95 VDDA.n69 GNDA 0.038853f
C96 VDDA.n70 GNDA 0.01649f
C97 VDDA.n74 GNDA 0.011669f
C98 VDDA.t25 GNDA 0.012635f
C99 VDDA.n76 GNDA 0.010041f
C100 VDDA.n84 GNDA 0.01214f
C101 VDDA.n94 GNDA 0.175163f
C102 VDDA.n96 GNDA 0.010041f
C103 VDDA.n97 GNDA 0.021493f
C104 VDDA.n98 GNDA 0.097987f
C105 VDDA.n99 GNDA 0.864337f
C106 Vin-.n0 GNDA 0.047608f
C107 Vin-.n1 GNDA 0.325376f
C108 Vin-.n2 GNDA 0.162777f
C109 Vin-.n3 GNDA 0.072622f
C110 Vin-.n4 GNDA 0.330576f
C111 Vin-.t4 GNDA 0.037206f
C112 Vin-.t3 GNDA 0.037206f
C113 Vin-.n5 GNDA 0.136197f
C114 Vin-.t6 GNDA 0.037206f
C115 Vin-.t5 GNDA 0.037206f
C116 Vin-.n6 GNDA 0.134212f
C117 Vin-.n7 GNDA 0.391595f
C118 Vin-.t1 GNDA 0.101166f
C119 Vin-.t9 GNDA 0.063261f
C120 Vin-.n8 GNDA 0.284839f
C121 Vin-.n9 GNDA 0.07277f
C122 Vin-.t7 GNDA 0.033486f
C123 Vin-.t10 GNDA 0.033486f
C124 Vin-.n10 GNDA 0.041639f
C125 Vin-.n11 GNDA 0.041639f
C126 Vin-.n12 GNDA 0.07277f
C127 Vin-.t8 GNDA 0.063261f
C128 Vin-.n13 GNDA 0.153586f
C129 Vin-.n14 GNDA 0.192224f
C130 Vin-.t0 GNDA 0.115957f
C131 Vin-.n15 GNDA 0.565395f
C132 Vin-.n16 GNDA 1.05108f
C133 Vin-.n17 GNDA 0.162777f
C134 Vin-.n18 GNDA 0.105859f
C135 Vin-.n19 GNDA 0.080691f
C136 Vin-.n20 GNDA 0.323119f
C137 Vin-.t2 GNDA 0.071157f
C138 Vin-.n21 GNDA 0.071948f
C139 Vin-.n22 GNDA 0.080691f
C140 Vin-.n23 GNDA 0.072622f
C141 Vin-.n24 GNDA 0.631116f
C142 Vin-.n25 GNDA 0.379166f
C143 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6.Emitter GNDA 0.084511f
C144 V_TOP.t1 GNDA 0.013008f
C145 V_TOP.t0 GNDA 0.013008f
C146 V_TOP.n0 GNDA 0.048818f
C147 V_TOP.t5 GNDA 0.013008f
C148 V_TOP.t2 GNDA 0.013008f
C149 V_TOP.n1 GNDA 0.047513f
C150 V_TOP.n2 GNDA 0.234076f
C151 V_TOP.t4 GNDA 0.013008f
C152 V_TOP.t8 GNDA 0.013008f
C153 V_TOP.n3 GNDA 0.046629f
C154 V_TOP.t7 GNDA 0.087254f
C155 V_TOP.t6 GNDA 1.066f
C156 V_TOP.n4 GNDA 0.310646f
C157 V_TOP.n5 GNDA 0.134354f
C158 V_TOP.n6 GNDA 0.116934f
C159 V_TOP.t13 GNDA 0.023383f
C160 V_TOP.t21 GNDA 0.11122f
C161 V_TOP.t15 GNDA 0.11122f
C162 V_TOP.t20 GNDA 0.11122f
C163 V_TOP.t11 GNDA 0.11122f
C164 V_TOP.t17 GNDA 0.11122f
C165 V_TOP.t10 GNDA 0.11122f
C166 V_TOP.t16 GNDA 0.11122f
C167 V_TOP.t9 GNDA 0.11122f
C168 V_TOP.t14 GNDA 0.11122f
C169 V_TOP.t19 GNDA 0.11122f
C170 V_TOP.t12 GNDA 0.11122f
C171 V_TOP.t18 GNDA 0.14182f
C172 V_TOP.n7 GNDA 0.072815f
C173 V_TOP.n8 GNDA 0.052683f
C174 V_TOP.n9 GNDA 0.052683f
C175 V_TOP.n10 GNDA 0.052683f
C176 V_TOP.n11 GNDA 0.052683f
C177 V_TOP.n12 GNDA 0.052683f
C178 V_TOP.n13 GNDA 0.052683f
C179 V_TOP.n14 GNDA 0.052683f
C180 V_TOP.n15 GNDA 0.052683f
C181 V_TOP.n16 GNDA 0.052238f
C182 V_TOP.n17 GNDA 0.067442f
C183 V_TOP.n18 GNDA 0.14944f
C184 V_TOP.n19 GNDA 0.043484f
C185 V_TOP.t3 GNDA 0.034232f
.ends

