* PEX produced on Mon Feb  3 03:10:48 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from charge_pump_full_magic.ext - technology: sky130A

.subckt charge_pump_full_magic VDDA V_OUT GNDA UP_PFD DOWN_PFD I_IN
X0 GNDA DOWN_PFD a_1870_3900# GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 GNDA I_IN a_0_4990# GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X2 VDDA a_1710_3900# V_OUT VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X3 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out charge_pump_full_5_0.opamp_cell_0.p_right GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X4 a_2870_3900# a_2580_3900# sky130_fd_pr__cap_mim_m3_1 l=2.6 w=2.6
X5 a_1710_3900# a_1420_3900# sky130_fd_pr__cap_mim_m3_1 l=6 w=4.2
X6 charge_pump_full_5_0.opamp_cell_0.v_common_p charge_pump_full_5_0.opamp_cell_0.p_bias VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X7 a_1130_3900# a_840_3900# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X8 a_2870_3900# a_2580_3900# I_IN GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X9 V_OUT a_1710_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X10 V_OUT a_1710_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X11 a_0_4990# I_IN GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X12 charge_pump_full_5_0.opamp_cell_0.v_common_p a_0_4990# charge_pump_full_5_0.opamp_cell_0.p_right VDDA sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X13 VDDA a_1710_3900# V_OUT VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X14 charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.n_left VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X15 a_1710_3900# a_1420_3900# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X16 charge_pump_full_5_0.opamp_cell_0.p_left charge_pump_full_5_0.opamp_cell_0.p_left GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X17 charge_pump_full_5_0.opamp_cell_0.n_right a_8046_2450# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X18 a_0_4990# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X19 charge_pump_full_5_0.opamp_cell_0.v_common_n a_0_4990# charge_pump_full_5_0.opamp_cell_0.n_right GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X20 V_OUT a_1710_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X21 a_840_3900# UP_PFD VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X22 a_2580_3900# a_2290_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X23 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out a_5120_2450# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X24 VDDA charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.n_right VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X25 charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.opamp_cell_0.n_bias GNDA GNDA sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X26 VDDA charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out a_0_4990# VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X27 I_IN I_IN GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X28 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.p_bias VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X29 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out charge_pump_full_5_0.opamp_cell_0.n_right VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X30 charge_pump_full_5_0.opamp_cell_0.n_right a_0_4990# charge_pump_full_5_0.opamp_cell_0.v_common_n GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X31 V_OUT a_2870_3900# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X32 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.n_bias GNDA sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X33 VDDA a_1710_3900# V_OUT VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X34 charge_pump_full_5_0.opamp_cell_0.v_common_p charge_pump_full_5_0.opamp_cell_0.p_bias VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X35 a_1710_3900# a_1130_3900# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X36 GNDA charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.opamp_cell_0.n_bias GNDA sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X37 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.p_bias VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X38 GNDA I_IN I_IN GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X39 GNDA charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.opamp_cell_0.v_common_n GNDA sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X40 a_840_3900# UP_PFD GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X41 a_2580_3900# a_2290_3900# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X42 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out charge_pump_full_5_0.opamp_cell_0.p_right GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X43 GNDA a_2870_3900# V_OUT GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X44 VDDA charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.p_bias VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X45 charge_pump_full_5_0.opamp_cell_0.p_right a_0_4990# charge_pump_full_5_0.opamp_cell_0.v_common_p VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X46 I_IN I_IN GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X47 VDDA charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out a_0_4990# VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X48 a_0_4990# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X49 VDDA charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.v_common_p VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X50 GNDA charge_pump_full_5_0.opamp_cell_0.p_left charge_pump_full_5_0.opamp_cell_0.p_right GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X51 GNDA V_OUT sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X52 GNDA a_15082_6070# sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X53 V_OUT a_15082_6070# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X54 GNDA I_IN I_IN GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X55 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out a_8046_2450# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X56 a_0_4990# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X57 a_1420_3900# a_1130_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X58 V_OUT a_1710_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X59 a_2290_3900# GNDA a_1870_3900# VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X60 charge_pump_full_5_0.opamp_cell_0.v_common_p V_OUT charge_pump_full_5_0.opamp_cell_0.p_left VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X61 VDDA charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out a_0_4990# VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X62 charge_pump_full_5_0.opamp_cell_0.n_right charge_pump_full_5_0.opamp_cell_0.n_left VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X63 a_1710_3900# a_1130_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X64 VDDA charge_pump_full_5_0.opamp_cell_0.n_right charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X65 charge_pump_full_5_0.opamp_cell_0.p_right charge_pump_full_5_0.opamp_cell_0.p_left GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X66 VDDA a_1710_3900# V_OUT VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X67 VDDA DOWN_PFD a_1870_3900# VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X68 charge_pump_full_5_0.opamp_cell_0.v_common_n V_OUT charge_pump_full_5_0.opamp_cell_0.n_left GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X69 a_0_4990# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X70 charge_pump_full_5_0.opamp_cell_0.p_left V_OUT charge_pump_full_5_0.opamp_cell_0.v_common_p VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X71 VDDA charge_pump_full_5_0.opamp_cell_0.n_right charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X72 GNDA charge_pump_full_5_0.opamp_cell_0.p_right charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X73 a_5120_2450# charge_pump_full_5_0.opamp_cell_0.p_right GNDA sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X74 a_1130_3900# a_840_3900# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X75 a_2870_3900# a_2290_3900# I_IN VDDA sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X76 VDDA charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.n_left VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X77 GNDA I_IN a_0_4990# GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X78 V_OUT a_2870_3900# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X79 a_1420_3900# a_1130_3900# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X80 GNDA charge_pump_full_5_0.opamp_cell_0.p_left charge_pump_full_5_0.opamp_cell_0.p_left GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X81 GNDA charge_pump_full_5_0.opamp_cell_0.p_right charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X82 a_2290_3900# VDDA a_1870_3900# GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X83 GNDA a_2870_3900# V_OUT GNDA sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X84 VDDA charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out a_0_4990# VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X85 VDDA charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.p_bias VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X86 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out charge_pump_full_5_0.opamp_cell_0.n_right VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X87 charge_pump_full_5_0.opamp_cell_0.n_left V_OUT charge_pump_full_5_0.opamp_cell_0.v_common_n GNDA sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X88 a_0_4990# I_IN GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X89 VDDA charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.v_common_p VDDA sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X90 a_2870_3900# a_2290_3900# GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X91 charge_pump_full_5_0.opamp_cell_0.v_common_n charge_pump_full_5_0.opamp_cell_0.n_bias GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
C0 charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.opamp_cell_0.p_bias 0.148683f
C1 a_0_4990# charge_pump_full_5_0.opamp_cell_0.p_right 0.17573f
C2 charge_pump_full_5_0.opamp_cell_0.p_left charge_pump_full_5_0.opamp_cell_0.p_bias 0.090982f
C3 DOWN_PFD a_0_4990# 0.130956f
C4 a_840_3900# a_0_4990# 0.06669f
C5 a_1420_3900# a_0_4990# 0.100664f
C6 DOWN_PFD a_1870_3900# 0.068964f
C7 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out charge_pump_full_5_0.opamp_cell_0.n_right 0.565978f
C8 charge_pump_full_5_0.opamp_cell_0.n_left a_0_4990# 0.098351f
C9 V_OUT charge_pump_full_5_0.opamp_cell_0.p_right 0.249338f
C10 charge_pump_full_5_0.opamp_cell_0.v_common_n charge_pump_full_5_0.opamp_cell_0.n_left 0.096235f
C11 V_OUT a_2870_3900# 0.313706f
C12 a_8046_2450# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.187394f
C13 charge_pump_full_5_0.opamp_cell_0.v_common_p charge_pump_full_5_0.opamp_cell_0.n_right 0.019186f
C14 a_1420_3900# V_OUT 0.203398f
C15 V_OUT charge_pump_full_5_0.opamp_cell_0.n_left 0.047975f
C16 a_1710_3900# a_0_4990# 0.083727f
C17 I_IN a_0_4990# 0.453001f
C18 a_1710_3900# a_1870_3900# 0.252612f
C19 charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.157586f
C20 a_1710_3900# V_OUT 0.56786f
C21 VDDA a_2580_3900# 0.361352f
C22 a_1130_3900# a_2290_3900# 0.047593f
C23 charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.p_right 0.072353f
C24 DOWN_PFD a_840_3900# 0.016162f
C25 a_5120_2450# charge_pump_full_5_0.opamp_cell_0.p_right 0.027587f
C26 DOWN_PFD a_1420_3900# 0.010851f
C27 a_1420_3900# a_2870_3900# 0.010789f
C28 a_1130_3900# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.18867f
C29 a_1420_3900# a_5120_2450# 0.100687f
C30 charge_pump_full_5_0.opamp_cell_0.p_left charge_pump_full_5_0.opamp_cell_0.v_common_p 0.174112f
C31 VDDA charge_pump_full_5_0.opamp_cell_0.n_right 0.73301f
C32 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.091153f
C33 DOWN_PFD a_1710_3900# 0.014109f
C34 a_1710_3900# a_2870_3900# 1.53843f
C35 I_IN DOWN_PFD 0.218332f
C36 a_1420_3900# a_1710_3900# 1.84668f
C37 I_IN a_2870_3900# 0.257967f
C38 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.v_common_p 0.608314f
C39 VDDA UP_PFD 0.20974f
C40 VDDA charge_pump_full_5_0.opamp_cell_0.p_left 0.129595f
C41 I_IN a_1710_3900# 0.037077f
C42 a_0_4990# a_2580_3900# 0.035849f
C43 VDDA a_1130_3900# 1.86766f
C44 VDDA charge_pump_full_5_0.opamp_cell_0.p_bias 4.59302f
C45 V_OUT a_2580_3900# 0.231008f
C46 a_0_4990# charge_pump_full_5_0.opamp_cell_0.n_right 0.016449f
C47 charge_pump_full_5_0.opamp_cell_0.v_common_n charge_pump_full_5_0.opamp_cell_0.n_right 0.10809f
C48 a_8046_2450# V_OUT 0.564385f
C49 a_2870_3900# a_2580_3900# 1.71852f
C50 a_1420_3900# a_2580_3900# 0.151144f
C51 VDDA a_2290_3900# 0.828477f
C52 charge_pump_full_5_0.opamp_cell_0.n_bias a_0_4990# 0.042036f
C53 UP_PFD a_0_4990# 0.041114f
C54 charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.opamp_cell_0.v_common_n 0.286889f
C55 charge_pump_full_5_0.opamp_cell_0.p_right charge_pump_full_5_0.opamp_cell_0.n_right 0.602936f
C56 charge_pump_full_5_0.opamp_cell_0.p_left a_0_4990# 0.103108f
C57 VDDA charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 4.62038f
C58 a_1130_3900# a_0_4990# 0.06808f
C59 charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.n_right 0.188651f
C60 a_1710_3900# a_2580_3900# 0.041266f
C61 V_OUT charge_pump_full_5_0.opamp_cell_0.p_left 0.182006f
C62 VDDA charge_pump_full_5_0.opamp_cell_0.v_common_p 2.01449f
C63 I_IN a_2580_3900# 0.29494f
C64 charge_pump_full_5_0.opamp_cell_0.p_bias a_0_4990# 0.141466f
C65 a_8046_2450# a_5120_2450# 0.371805f
C66 charge_pump_full_5_0.opamp_cell_0.n_bias charge_pump_full_5_0.opamp_cell_0.p_right 0.114142f
C67 V_OUT charge_pump_full_5_0.opamp_cell_0.p_bias 0.17648f
C68 charge_pump_full_5_0.opamp_cell_0.p_left charge_pump_full_5_0.opamp_cell_0.p_right 0.123547f
C69 DOWN_PFD UP_PFD 0.0436f
C70 a_840_3900# UP_PFD 0.065398f
C71 DOWN_PFD a_1130_3900# 0.058317f
C72 a_840_3900# a_1130_3900# 0.103876f
C73 a_1130_3900# a_1420_3900# 0.212799f
C74 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.p_right 0.016838f
C75 a_1870_3900# a_2290_3900# 0.253578f
C76 a_0_4990# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.623646f
C77 charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.p_bias 0.025924f
C78 a_5120_2450# charge_pump_full_5_0.opamp_cell_0.p_bias 0.020761f
C79 charge_pump_full_5_0.opamp_cell_0.v_common_n charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.057403f
C80 a_1130_3900# a_1710_3900# 0.193792f
C81 a_0_4990# charge_pump_full_5_0.opamp_cell_0.v_common_p 0.062421f
C82 V_OUT charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.180404f
C83 V_OUT charge_pump_full_5_0.opamp_cell_0.v_common_p 0.070614f
C84 a_2870_3900# a_2290_3900# 0.106599f
C85 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out charge_pump_full_5_0.opamp_cell_0.p_right 0.389947f
C86 a_1420_3900# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 1.84716f
C87 charge_pump_full_5_0.opamp_cell_0.p_right charge_pump_full_5_0.opamp_cell_0.v_common_p 0.170357f
C88 charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.048528f
C89 a_5120_2450# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.468482f
C90 V_OUT a_15082_6070# 2.20249f
C91 VDDA a_0_4990# 3.43501f
C92 VDDA a_1870_3900# 0.683927f
C93 a_1710_3900# a_2290_3900# 0.053508f
C94 I_IN a_2290_3900# 0.117646f
C95 charge_pump_full_5_0.opamp_cell_0.n_left charge_pump_full_5_0.opamp_cell_0.v_common_p 0.085408f
C96 VDDA V_OUT 3.31676f
C97 a_8046_2450# charge_pump_full_5_0.opamp_cell_0.n_right 0.028293f
C98 a_1710_3900# charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out 0.742675f
C99 VDDA charge_pump_full_5_0.opamp_cell_0.p_right 0.154177f
C100 DOWN_PFD VDDA 0.096195f
C101 VDDA a_2870_3900# 0.497611f
C102 VDDA a_840_3900# 0.575947f
C103 VDDA a_1420_3900# 2.25464f
C104 VDDA charge_pump_full_5_0.opamp_cell_0.n_left 0.829877f
C105 charge_pump_full_5_0.opamp_cell_0.p_bias charge_pump_full_5_0.opamp_cell_0.n_right 0.011765f
C106 charge_pump_full_5_0.opamp_cell_0.v_common_n a_0_4990# 0.164393f
C107 VDDA a_1710_3900# 4.22066f
C108 a_0_4990# a_1870_3900# 0.010789f
C109 I_IN VDDA 0.19824f
C110 V_OUT a_0_4990# 0.460948f
C111 V_OUT charge_pump_full_5_0.opamp_cell_0.v_common_n 0.029566f
C112 a_2580_3900# a_2290_3900# 0.229502f
C113 I_IN GNDA 5.01709f
C114 DOWN_PFD GNDA 1.4812f
C115 UP_PFD GNDA 0.660505f
C116 V_OUT GNDA 24.163f
C117 VDDA GNDA 24.7686f
C118 a_8046_2450# GNDA 3.33383f
C119 a_5120_2450# GNDA 3.32008f
C120 charge_pump_full_5_0.opamp_cell_0.n_bias GNDA 4.14103f
C121 charge_pump_full_5_0.opamp_cell_0.v_common_n GNDA 1.23735f
C122 charge_pump_full_5_0.opamp_cell_0.p_right GNDA 3.50336f
C123 charge_pump_full_5_0.opamp_cell_0.p_left GNDA 1.06547f
C124 charge_pump_full_5_0.opamp_cell_0.n_right GNDA 2.33883f
C125 charge_pump_full_5_0.opamp_cell_0.n_left GNDA 0.460695f
C126 charge_pump_full_5_0.opamp_cell_0.v_common_p GNDA 0.046438f
C127 charge_pump_full_5_0.opamp_cell_0.p_bias GNDA 3.28171f
C128 a_2870_3900# GNDA 3.50986f
C129 a_2580_3900# GNDA 3.23767f
C130 a_1870_3900# GNDA 0.560184f
C131 a_2290_3900# GNDA 1.39218f
C132 a_1420_3900# GNDA 2.58292f
C133 a_840_3900# GNDA 0.522028f
C134 a_1130_3900# GNDA 0.744855f
C135 a_1710_3900# GNDA 2.00507f
C136 charge_pump_full_5_0.charge_pump_cell_0.OPAMP_out GNDA 5.95931f
C137 a_0_4990# GNDA 9.052549f
C138 a_15082_6070# GNDA 62.2621f
.ends

