magic
tech sky130A
timestamp 1738241744
<< nwell >>
rect 8750 1770 10680 2355
<< pwell >>
rect 9430 1670 9445 1675
rect 8925 1540 10240 1665
rect 9490 1535 10240 1540
rect 9490 1530 9855 1535
rect 9490 1470 9655 1530
rect 9770 1495 9855 1530
rect 9770 1480 9820 1495
rect 9840 1480 9855 1495
rect 9770 1470 9855 1480
rect 9800 1465 9840 1470
rect 9850 1440 9890 1465
<< nmos >>
rect 8995 1560 9010 1660
rect 9140 1560 9155 1660
rect 9285 1560 9300 1660
rect 9430 1560 9445 1660
rect 9575 1560 9590 1660
rect 9720 1560 9735 1660
rect 9865 1560 9880 1660
rect 10010 1560 10025 1660
rect 10155 1560 10170 1660
rect 8840 1305 8900 1405
rect 8950 1305 9010 1405
rect 9060 1305 9120 1405
rect 9170 1305 9230 1405
rect 9500 1305 9560 1405
rect 9610 1305 9670 1405
rect 9720 1305 9780 1405
rect 9830 1305 9890 1405
rect 10220 1305 10280 1405
rect 10330 1305 10390 1405
rect 10440 1305 10500 1405
rect 10550 1305 10610 1405
<< pmos >>
rect 8820 2235 8880 2335
rect 8930 2235 8990 2335
rect 9040 2235 9100 2335
rect 9150 2235 9210 2335
rect 9260 2235 9320 2335
rect 9370 2235 9430 2335
rect 9480 2235 9540 2335
rect 9590 2235 9650 2335
rect 9780 2235 9840 2335
rect 9890 2235 9950 2335
rect 10000 2235 10060 2335
rect 10110 2235 10170 2335
rect 10220 2235 10280 2335
rect 10330 2235 10390 2335
rect 10440 2235 10500 2335
rect 10550 2235 10610 2335
rect 8995 1790 9010 1990
rect 9140 1790 9155 1990
rect 9285 1790 9300 1990
rect 9430 1790 9445 1990
rect 9575 1790 9590 1990
rect 9720 1790 9735 1990
rect 9865 1790 9880 1990
rect 10010 1790 10025 1990
rect 10155 1790 10170 1990
<< ndiff >>
rect 8945 1645 8995 1660
rect 8945 1575 8960 1645
rect 8980 1575 8995 1645
rect 8945 1560 8995 1575
rect 9010 1645 9060 1660
rect 9010 1575 9025 1645
rect 9045 1575 9060 1645
rect 9010 1560 9060 1575
rect 9090 1645 9140 1660
rect 9090 1575 9105 1645
rect 9125 1575 9140 1645
rect 9090 1560 9140 1575
rect 9155 1645 9205 1660
rect 9155 1575 9170 1645
rect 9190 1575 9205 1645
rect 9155 1560 9205 1575
rect 9235 1645 9285 1660
rect 9235 1575 9250 1645
rect 9270 1575 9285 1645
rect 9235 1560 9285 1575
rect 9300 1645 9350 1660
rect 9300 1575 9315 1645
rect 9335 1575 9350 1645
rect 9300 1560 9350 1575
rect 9380 1645 9430 1660
rect 9380 1575 9395 1645
rect 9415 1575 9430 1645
rect 9380 1560 9430 1575
rect 9445 1645 9495 1660
rect 9445 1575 9460 1645
rect 9480 1575 9495 1645
rect 9445 1560 9495 1575
rect 9525 1645 9575 1660
rect 9525 1575 9540 1645
rect 9560 1575 9575 1645
rect 9525 1560 9575 1575
rect 9590 1645 9640 1660
rect 9590 1575 9605 1645
rect 9625 1575 9640 1645
rect 9590 1560 9640 1575
rect 9670 1645 9720 1660
rect 9670 1575 9685 1645
rect 9705 1575 9720 1645
rect 9670 1560 9720 1575
rect 9735 1645 9785 1660
rect 9735 1575 9750 1645
rect 9770 1575 9785 1645
rect 9735 1560 9785 1575
rect 9815 1645 9865 1660
rect 9815 1575 9830 1645
rect 9850 1575 9865 1645
rect 9815 1560 9865 1575
rect 9880 1645 9930 1660
rect 9880 1575 9895 1645
rect 9915 1575 9930 1645
rect 9880 1560 9930 1575
rect 9960 1645 10010 1660
rect 9960 1575 9975 1645
rect 9995 1575 10010 1645
rect 9960 1560 10010 1575
rect 10025 1645 10075 1660
rect 10025 1575 10040 1645
rect 10060 1575 10075 1645
rect 10025 1560 10075 1575
rect 10105 1645 10155 1660
rect 10105 1575 10120 1645
rect 10140 1575 10155 1645
rect 10105 1560 10155 1575
rect 10170 1645 10220 1660
rect 10170 1575 10185 1645
rect 10205 1575 10220 1645
rect 10170 1560 10220 1575
rect 8790 1390 8840 1405
rect 8790 1320 8805 1390
rect 8825 1320 8840 1390
rect 8790 1305 8840 1320
rect 8900 1390 8950 1405
rect 8900 1320 8915 1390
rect 8935 1320 8950 1390
rect 8900 1305 8950 1320
rect 9010 1390 9060 1405
rect 9010 1320 9025 1390
rect 9045 1320 9060 1390
rect 9010 1305 9060 1320
rect 9120 1390 9170 1405
rect 9120 1320 9135 1390
rect 9155 1320 9170 1390
rect 9120 1305 9170 1320
rect 9230 1390 9280 1405
rect 9230 1320 9245 1390
rect 9265 1320 9280 1390
rect 9230 1305 9280 1320
rect 9450 1390 9500 1405
rect 9450 1320 9465 1390
rect 9485 1320 9500 1390
rect 9450 1305 9500 1320
rect 9560 1390 9610 1405
rect 9560 1320 9575 1390
rect 9595 1320 9610 1390
rect 9560 1305 9610 1320
rect 9670 1390 9720 1405
rect 9670 1320 9685 1390
rect 9705 1320 9720 1390
rect 9670 1305 9720 1320
rect 9780 1390 9830 1405
rect 9780 1320 9795 1390
rect 9815 1320 9830 1390
rect 9780 1305 9830 1320
rect 9890 1390 9940 1405
rect 9890 1320 9905 1390
rect 9925 1320 9940 1390
rect 9890 1305 9940 1320
rect 10170 1390 10220 1405
rect 10170 1320 10185 1390
rect 10205 1320 10220 1390
rect 10170 1305 10220 1320
rect 10280 1390 10330 1405
rect 10280 1320 10295 1390
rect 10315 1320 10330 1390
rect 10280 1305 10330 1320
rect 10390 1390 10440 1405
rect 10390 1320 10405 1390
rect 10425 1320 10440 1390
rect 10390 1305 10440 1320
rect 10500 1390 10550 1405
rect 10500 1320 10515 1390
rect 10535 1320 10550 1390
rect 10500 1305 10550 1320
rect 10610 1390 10660 1405
rect 10610 1320 10625 1390
rect 10645 1320 10660 1390
rect 10610 1305 10660 1320
<< pdiff >>
rect 8770 2320 8820 2335
rect 8770 2250 8785 2320
rect 8805 2250 8820 2320
rect 8770 2235 8820 2250
rect 8880 2320 8930 2335
rect 8880 2250 8895 2320
rect 8915 2250 8930 2320
rect 8880 2235 8930 2250
rect 8990 2320 9040 2335
rect 8990 2250 9005 2320
rect 9025 2250 9040 2320
rect 8990 2235 9040 2250
rect 9100 2320 9150 2335
rect 9100 2250 9115 2320
rect 9135 2250 9150 2320
rect 9100 2235 9150 2250
rect 9210 2320 9260 2335
rect 9210 2250 9225 2320
rect 9245 2250 9260 2320
rect 9210 2235 9260 2250
rect 9320 2320 9370 2335
rect 9320 2250 9335 2320
rect 9355 2250 9370 2320
rect 9320 2235 9370 2250
rect 9430 2320 9480 2335
rect 9430 2250 9445 2320
rect 9465 2250 9480 2320
rect 9430 2235 9480 2250
rect 9540 2320 9590 2335
rect 9540 2250 9555 2320
rect 9575 2250 9590 2320
rect 9540 2235 9590 2250
rect 9650 2320 9700 2335
rect 9650 2250 9665 2320
rect 9685 2250 9700 2320
rect 9650 2235 9700 2250
rect 9730 2320 9780 2335
rect 9730 2250 9745 2320
rect 9765 2250 9780 2320
rect 9730 2235 9780 2250
rect 9840 2320 9890 2335
rect 9840 2250 9855 2320
rect 9875 2250 9890 2320
rect 9840 2235 9890 2250
rect 9950 2320 10000 2335
rect 9950 2250 9965 2320
rect 9985 2250 10000 2320
rect 9950 2235 10000 2250
rect 10060 2320 10110 2335
rect 10060 2250 10075 2320
rect 10095 2250 10110 2320
rect 10060 2235 10110 2250
rect 10170 2320 10220 2335
rect 10170 2250 10185 2320
rect 10205 2250 10220 2320
rect 10170 2235 10220 2250
rect 10280 2320 10330 2335
rect 10280 2250 10295 2320
rect 10315 2250 10330 2320
rect 10280 2235 10330 2250
rect 10390 2320 10440 2335
rect 10390 2250 10405 2320
rect 10425 2250 10440 2320
rect 10390 2235 10440 2250
rect 10500 2320 10550 2335
rect 10500 2250 10515 2320
rect 10535 2250 10550 2320
rect 10500 2235 10550 2250
rect 10610 2320 10660 2335
rect 10610 2250 10625 2320
rect 10645 2250 10660 2320
rect 10610 2235 10660 2250
rect 8945 1975 8995 1990
rect 8945 1805 8960 1975
rect 8980 1805 8995 1975
rect 8945 1790 8995 1805
rect 9010 1975 9060 1990
rect 9010 1805 9025 1975
rect 9045 1805 9060 1975
rect 9010 1790 9060 1805
rect 9090 1975 9140 1990
rect 9090 1805 9105 1975
rect 9125 1805 9140 1975
rect 9090 1790 9140 1805
rect 9155 1975 9205 1990
rect 9155 1805 9170 1975
rect 9190 1805 9205 1975
rect 9155 1790 9205 1805
rect 9235 1975 9285 1990
rect 9235 1805 9250 1975
rect 9270 1805 9285 1975
rect 9235 1790 9285 1805
rect 9300 1975 9350 1990
rect 9300 1805 9315 1975
rect 9335 1805 9350 1975
rect 9300 1790 9350 1805
rect 9380 1975 9430 1990
rect 9380 1805 9395 1975
rect 9415 1805 9430 1975
rect 9380 1790 9430 1805
rect 9445 1975 9495 1990
rect 9445 1805 9460 1975
rect 9480 1805 9495 1975
rect 9445 1790 9495 1805
rect 9525 1975 9575 1990
rect 9525 1805 9540 1975
rect 9560 1805 9575 1975
rect 9525 1790 9575 1805
rect 9590 1975 9640 1990
rect 9590 1805 9605 1975
rect 9625 1805 9640 1975
rect 9590 1790 9640 1805
rect 9670 1975 9720 1990
rect 9670 1805 9685 1975
rect 9705 1805 9720 1975
rect 9670 1790 9720 1805
rect 9735 1975 9785 1990
rect 9735 1805 9750 1975
rect 9770 1805 9785 1975
rect 9735 1790 9785 1805
rect 9815 1975 9865 1990
rect 9815 1805 9830 1975
rect 9850 1805 9865 1975
rect 9815 1790 9865 1805
rect 9880 1975 9930 1990
rect 9880 1805 9895 1975
rect 9915 1805 9930 1975
rect 9880 1790 9930 1805
rect 9960 1975 10010 1990
rect 9960 1805 9975 1975
rect 9995 1805 10010 1975
rect 9960 1790 10010 1805
rect 10025 1975 10075 1990
rect 10025 1805 10040 1975
rect 10060 1805 10075 1975
rect 10025 1790 10075 1805
rect 10105 1975 10155 1990
rect 10105 1805 10120 1975
rect 10140 1805 10155 1975
rect 10105 1790 10155 1805
rect 10170 1975 10220 1990
rect 10170 1805 10185 1975
rect 10205 1805 10220 1975
rect 10170 1790 10220 1805
<< ndiffc >>
rect 8960 1575 8980 1645
rect 9025 1575 9045 1645
rect 9105 1575 9125 1645
rect 9170 1575 9190 1645
rect 9250 1575 9270 1645
rect 9315 1575 9335 1645
rect 9395 1575 9415 1645
rect 9460 1575 9480 1645
rect 9540 1575 9560 1645
rect 9605 1575 9625 1645
rect 9685 1575 9705 1645
rect 9750 1575 9770 1645
rect 9830 1575 9850 1645
rect 9895 1575 9915 1645
rect 9975 1575 9995 1645
rect 10040 1575 10060 1645
rect 10120 1575 10140 1645
rect 10185 1575 10205 1645
rect 8805 1320 8825 1390
rect 8915 1320 8935 1390
rect 9025 1320 9045 1390
rect 9135 1320 9155 1390
rect 9245 1320 9265 1390
rect 9465 1320 9485 1390
rect 9575 1320 9595 1390
rect 9685 1320 9705 1390
rect 9795 1320 9815 1390
rect 9905 1320 9925 1390
rect 10185 1320 10205 1390
rect 10295 1320 10315 1390
rect 10405 1320 10425 1390
rect 10515 1320 10535 1390
rect 10625 1320 10645 1390
<< pdiffc >>
rect 8785 2250 8805 2320
rect 8895 2250 8915 2320
rect 9005 2250 9025 2320
rect 9115 2250 9135 2320
rect 9225 2250 9245 2320
rect 9335 2250 9355 2320
rect 9445 2250 9465 2320
rect 9555 2250 9575 2320
rect 9665 2250 9685 2320
rect 9745 2250 9765 2320
rect 9855 2250 9875 2320
rect 9965 2250 9985 2320
rect 10075 2250 10095 2320
rect 10185 2250 10205 2320
rect 10295 2250 10315 2320
rect 10405 2250 10425 2320
rect 10515 2250 10535 2320
rect 10625 2250 10645 2320
rect 8960 1805 8980 1975
rect 9025 1805 9045 1975
rect 9105 1805 9125 1975
rect 9170 1805 9190 1975
rect 9250 1805 9270 1975
rect 9315 1805 9335 1975
rect 9395 1805 9415 1975
rect 9460 1805 9480 1975
rect 9540 1805 9560 1975
rect 9605 1805 9625 1975
rect 9685 1805 9705 1975
rect 9750 1805 9770 1975
rect 9830 1805 9850 1975
rect 9895 1805 9915 1975
rect 9975 1805 9995 1975
rect 10040 1805 10060 1975
rect 10120 1805 10140 1975
rect 10185 1805 10205 1975
<< psubdiff >>
rect 10250 1645 10300 1660
rect 10250 1575 10265 1645
rect 10285 1575 10300 1645
rect 10250 1560 10300 1575
<< nsubdiff >>
rect 10250 1975 10300 1990
rect 10250 1805 10265 1975
rect 10285 1805 10300 1975
rect 10250 1790 10300 1805
<< psubdiffcont >>
rect 10265 1575 10285 1645
<< nsubdiffcont >>
rect 10265 1805 10285 1975
<< poly >>
rect 8820 2335 8880 2350
rect 8930 2335 8990 2350
rect 9040 2335 9100 2350
rect 9150 2335 9210 2350
rect 9260 2335 9320 2350
rect 9370 2335 9430 2350
rect 9480 2335 9540 2350
rect 9590 2335 9650 2350
rect 9780 2335 9840 2350
rect 9890 2335 9950 2350
rect 10000 2335 10060 2350
rect 10110 2335 10170 2350
rect 10220 2335 10280 2350
rect 10330 2335 10390 2350
rect 10440 2335 10500 2350
rect 10550 2335 10610 2350
rect 8820 2225 8880 2235
rect 8930 2225 8990 2235
rect 9040 2225 9100 2235
rect 9150 2225 9210 2235
rect 9260 2225 9320 2235
rect 9370 2225 9430 2235
rect 9480 2225 9540 2235
rect 9590 2225 9650 2235
rect 8820 2205 9650 2225
rect 9780 2225 9840 2235
rect 9890 2225 9950 2235
rect 10000 2225 10060 2235
rect 10110 2225 10170 2235
rect 10220 2225 10280 2235
rect 10330 2225 10390 2235
rect 10440 2225 10500 2235
rect 10550 2225 10610 2235
rect 9780 2210 10610 2225
rect 10635 2210 10675 2220
rect 9400 2120 9415 2205
rect 9385 2110 9425 2120
rect 9385 2090 9395 2110
rect 9415 2090 9425 2110
rect 9385 2080 9425 2090
rect 9285 2040 10170 2055
rect 10345 2045 10360 2210
rect 10635 2190 10645 2210
rect 10665 2190 10675 2210
rect 10635 2180 10675 2190
rect 8995 1990 9010 2005
rect 9140 1990 9155 2005
rect 9285 1990 9300 2040
rect 9430 1990 9445 2005
rect 9575 1990 9590 2005
rect 9720 1990 9735 2005
rect 9865 1990 9880 2005
rect 10010 1990 10025 2005
rect 10155 1990 10170 2040
rect 10330 2035 10370 2045
rect 10330 2015 10340 2035
rect 10360 2015 10370 2035
rect 10330 2005 10370 2015
rect 10635 1815 10650 2180
rect 10635 1800 10885 1815
rect 8995 1735 9010 1790
rect 9140 1750 9155 1790
rect 9285 1750 9300 1790
rect 9430 1775 9445 1790
rect 8630 1720 9010 1735
rect 8995 1660 9010 1720
rect 9115 1740 9155 1750
rect 9115 1720 9125 1740
rect 9145 1720 9155 1740
rect 9115 1710 9155 1720
rect 9260 1740 9300 1750
rect 9260 1720 9270 1740
rect 9290 1720 9300 1740
rect 9325 1765 9445 1775
rect 9325 1745 9335 1765
rect 9355 1760 9445 1765
rect 9355 1745 9365 1760
rect 9325 1735 9365 1745
rect 9260 1710 9300 1720
rect 9140 1660 9155 1710
rect 9285 1685 9300 1710
rect 9285 1670 9445 1685
rect 9285 1660 9300 1670
rect 9430 1660 9445 1670
rect 9575 1660 9590 1790
rect 9720 1780 9735 1790
rect 9640 1765 9735 1780
rect 9760 1765 9800 1775
rect 9865 1765 9880 1790
rect 10010 1765 10025 1790
rect 10155 1775 10170 1790
rect 9640 1715 9655 1765
rect 9760 1745 9770 1765
rect 9790 1750 10135 1765
rect 9790 1745 9800 1750
rect 9760 1740 9800 1745
rect 9615 1705 9655 1715
rect 9800 1710 9840 1715
rect 9615 1685 9625 1705
rect 9645 1685 9655 1705
rect 9615 1675 9655 1685
rect 9720 1705 9840 1710
rect 9720 1695 9810 1705
rect 9720 1660 9735 1695
rect 9800 1685 9810 1695
rect 9830 1685 9840 1705
rect 9800 1675 9840 1685
rect 9865 1660 9880 1750
rect 10120 1730 10135 1750
rect 10120 1715 10170 1730
rect 9905 1700 9945 1710
rect 9905 1680 9915 1700
rect 9935 1685 9945 1700
rect 9935 1680 10025 1685
rect 9905 1670 10025 1680
rect 10010 1660 10025 1670
rect 10155 1660 10170 1715
rect 10345 1705 10385 1715
rect 10345 1685 10355 1705
rect 10375 1685 10385 1705
rect 10345 1675 10385 1685
rect 8995 1545 9010 1560
rect 9140 1545 9155 1560
rect 9285 1545 9300 1560
rect 9430 1545 9445 1560
rect 9575 1520 9590 1560
rect 9720 1545 9735 1560
rect 8630 1505 9590 1520
rect 9865 1480 9880 1560
rect 10010 1545 10025 1560
rect 10010 1535 10065 1545
rect 10010 1515 10035 1535
rect 10055 1515 10065 1535
rect 10010 1505 10065 1515
rect 10155 1480 10170 1560
rect 9800 1470 9840 1480
rect 8795 1450 8835 1460
rect 8795 1430 8805 1450
rect 8825 1440 8835 1450
rect 9015 1450 9055 1460
rect 9015 1440 9025 1450
rect 8825 1430 9025 1440
rect 9045 1440 9055 1450
rect 9235 1450 9275 1460
rect 9235 1440 9245 1450
rect 9045 1430 9245 1440
rect 9265 1440 9275 1450
rect 9800 1450 9810 1470
rect 9830 1450 9840 1470
rect 9865 1465 10170 1480
rect 9800 1440 9840 1450
rect 9265 1430 9890 1440
rect 10370 1430 10385 1675
rect 10635 1455 10650 1800
rect 10635 1445 10675 1455
rect 8795 1415 9890 1430
rect 8840 1405 8900 1415
rect 8950 1405 9010 1415
rect 9060 1405 9120 1415
rect 9170 1405 9230 1415
rect 9500 1405 9560 1415
rect 9610 1405 9670 1415
rect 9720 1405 9780 1415
rect 9830 1405 9890 1415
rect 10220 1415 10610 1430
rect 10635 1425 10645 1445
rect 10665 1425 10675 1445
rect 10635 1415 10675 1425
rect 10220 1405 10280 1415
rect 10330 1405 10390 1415
rect 10440 1405 10500 1415
rect 10550 1405 10610 1415
rect 8840 1290 8900 1305
rect 8950 1290 9010 1305
rect 9060 1290 9120 1305
rect 9170 1290 9230 1305
rect 9500 1290 9560 1305
rect 9610 1290 9670 1305
rect 9720 1290 9780 1305
rect 9830 1290 9890 1305
rect 10220 1290 10280 1305
rect 10330 1290 10390 1305
rect 10440 1290 10500 1305
rect 10550 1290 10610 1305
<< polycont >>
rect 9395 2090 9415 2110
rect 10645 2190 10665 2210
rect 10340 2015 10360 2035
rect 9125 1720 9145 1740
rect 9270 1720 9290 1740
rect 9335 1745 9355 1765
rect 9770 1745 9790 1765
rect 9625 1685 9645 1705
rect 9810 1685 9830 1705
rect 9915 1680 9935 1700
rect 10355 1685 10375 1705
rect 10035 1515 10055 1535
rect 8805 1430 8825 1450
rect 9025 1430 9045 1450
rect 9245 1430 9265 1450
rect 9810 1450 9830 1470
rect 10645 1425 10665 1445
<< locali >>
rect 8785 2350 9685 2370
rect 8785 2330 8805 2350
rect 9005 2330 9025 2350
rect 9225 2330 9245 2350
rect 9445 2330 9465 2350
rect 9665 2330 9685 2350
rect 9745 2350 10645 2370
rect 9745 2330 9765 2350
rect 9965 2330 9985 2350
rect 10185 2330 10205 2350
rect 10405 2330 10425 2350
rect 10625 2330 10645 2350
rect 8775 2320 8815 2330
rect 8775 2250 8785 2320
rect 8805 2250 8815 2320
rect 8775 2240 8815 2250
rect 8885 2320 8925 2330
rect 8885 2250 8895 2320
rect 8915 2250 8925 2320
rect 8885 2240 8925 2250
rect 8995 2320 9035 2330
rect 8995 2250 9005 2320
rect 9025 2250 9035 2320
rect 8995 2240 9035 2250
rect 9105 2320 9145 2330
rect 9105 2250 9115 2320
rect 9135 2250 9145 2320
rect 9105 2240 9145 2250
rect 9215 2320 9255 2330
rect 9215 2250 9225 2320
rect 9245 2250 9255 2320
rect 9215 2240 9255 2250
rect 9325 2320 9365 2330
rect 9325 2250 9335 2320
rect 9355 2250 9365 2320
rect 9325 2240 9365 2250
rect 9435 2320 9475 2330
rect 9435 2250 9445 2320
rect 9465 2250 9475 2320
rect 9435 2240 9475 2250
rect 9545 2320 9585 2330
rect 9545 2250 9555 2320
rect 9575 2250 9585 2320
rect 9545 2240 9585 2250
rect 9655 2320 9695 2330
rect 9655 2250 9665 2320
rect 9685 2250 9695 2320
rect 9655 2240 9695 2250
rect 9735 2320 9775 2330
rect 9735 2250 9745 2320
rect 9765 2250 9775 2320
rect 9735 2240 9775 2250
rect 9845 2320 9885 2330
rect 9845 2250 9855 2320
rect 9875 2250 9885 2320
rect 9845 2240 9885 2250
rect 9955 2320 9995 2330
rect 9955 2250 9965 2320
rect 9985 2250 9995 2320
rect 9955 2240 9995 2250
rect 10065 2320 10105 2330
rect 10065 2250 10075 2320
rect 10095 2250 10105 2320
rect 10065 2240 10105 2250
rect 10175 2320 10215 2330
rect 10175 2250 10185 2320
rect 10205 2250 10215 2320
rect 10175 2240 10215 2250
rect 10285 2320 10325 2330
rect 10285 2250 10295 2320
rect 10315 2250 10325 2320
rect 10285 2240 10325 2250
rect 10395 2320 10435 2330
rect 10395 2250 10405 2320
rect 10425 2250 10435 2320
rect 10395 2240 10435 2250
rect 10505 2320 10545 2330
rect 10505 2250 10515 2320
rect 10535 2250 10545 2320
rect 10505 2240 10545 2250
rect 10615 2320 10655 2330
rect 10615 2250 10625 2320
rect 10645 2250 10655 2320
rect 10615 2240 10655 2250
rect 8785 2220 8805 2240
rect 9665 2235 9685 2240
rect 8730 2200 8805 2220
rect 10635 2220 10655 2240
rect 10635 2210 10675 2220
rect 8730 1545 8750 2200
rect 10635 2190 10645 2210
rect 10665 2190 10675 2210
rect 10635 2180 10675 2190
rect 9315 2140 10835 2160
rect 9315 1985 9335 2140
rect 9385 2110 9425 2120
rect 9385 2090 9395 2110
rect 9415 2090 9425 2110
rect 9385 2080 9425 2090
rect 9395 1985 9415 2080
rect 10330 2035 10370 2045
rect 10330 2025 10340 2035
rect 9460 2015 10340 2025
rect 10360 2025 10370 2035
rect 10360 2015 10795 2025
rect 9460 2005 10795 2015
rect 9460 1985 9480 2005
rect 10185 1985 10205 2005
rect 8950 1975 8990 1985
rect 8950 1805 8960 1975
rect 8980 1805 8990 1975
rect 8950 1795 8990 1805
rect 9015 1975 9055 1985
rect 9015 1805 9025 1975
rect 9045 1805 9055 1975
rect 9015 1795 9055 1805
rect 9095 1975 9135 1985
rect 9095 1805 9105 1975
rect 9125 1805 9135 1975
rect 9095 1795 9135 1805
rect 9160 1975 9200 1985
rect 9160 1805 9170 1975
rect 9190 1805 9200 1975
rect 9160 1795 9200 1805
rect 9240 1975 9280 1985
rect 9240 1805 9250 1975
rect 9270 1805 9280 1975
rect 9240 1795 9280 1805
rect 9305 1975 9345 1985
rect 9305 1805 9315 1975
rect 9335 1805 9345 1975
rect 9305 1795 9345 1805
rect 9385 1975 9425 1985
rect 9385 1805 9395 1975
rect 9415 1805 9425 1975
rect 9385 1795 9425 1805
rect 9450 1975 9490 1985
rect 9450 1805 9460 1975
rect 9480 1805 9490 1975
rect 9450 1795 9490 1805
rect 9530 1975 9570 1985
rect 9530 1805 9540 1975
rect 9560 1805 9570 1975
rect 9530 1795 9570 1805
rect 9595 1975 9635 1985
rect 9595 1805 9605 1975
rect 9625 1825 9635 1975
rect 9675 1975 9715 1985
rect 9625 1805 9640 1825
rect 9595 1795 9640 1805
rect 9675 1805 9685 1975
rect 9705 1805 9715 1975
rect 9675 1795 9715 1805
rect 9740 1975 9780 1985
rect 9740 1805 9750 1975
rect 9770 1805 9780 1975
rect 9740 1795 9780 1805
rect 9820 1975 9860 1985
rect 9820 1805 9830 1975
rect 9850 1805 9860 1975
rect 9820 1795 9860 1805
rect 9885 1975 9925 1985
rect 9885 1805 9895 1975
rect 9915 1805 9925 1975
rect 9885 1795 9925 1805
rect 9965 1975 10005 1985
rect 9965 1805 9975 1975
rect 9995 1805 10005 1975
rect 9965 1795 10005 1805
rect 10030 1975 10070 1985
rect 10030 1805 10040 1975
rect 10060 1805 10070 1975
rect 10030 1795 10070 1805
rect 10110 1975 10150 1985
rect 10110 1805 10120 1975
rect 10140 1805 10150 1975
rect 10110 1795 10150 1805
rect 10175 1975 10215 1985
rect 10175 1805 10185 1975
rect 10205 1805 10215 1975
rect 10175 1795 10215 1805
rect 10255 1975 10295 1985
rect 10255 1805 10265 1975
rect 10285 1805 10295 1975
rect 10255 1795 10295 1805
rect 9035 1740 9055 1795
rect 9115 1740 9155 1750
rect 9035 1720 9125 1740
rect 9145 1720 9155 1740
rect 9035 1655 9055 1720
rect 9115 1710 9155 1720
rect 9180 1740 9200 1795
rect 9325 1775 9345 1795
rect 9325 1765 9365 1775
rect 9260 1740 9300 1750
rect 9180 1720 9270 1740
rect 9290 1720 9300 1740
rect 9180 1655 9200 1720
rect 9260 1710 9300 1720
rect 9325 1745 9335 1765
rect 9355 1745 9365 1765
rect 9325 1735 9365 1745
rect 9325 1655 9345 1735
rect 9395 1655 9415 1795
rect 9450 1655 9470 1795
rect 9550 1775 9570 1795
rect 9685 1775 9705 1795
rect 9550 1755 9705 1775
rect 9550 1655 9570 1755
rect 9615 1705 9655 1715
rect 9615 1685 9625 1705
rect 9645 1685 9655 1705
rect 9615 1675 9655 1685
rect 9615 1655 9635 1675
rect 9685 1655 9705 1755
rect 9750 1775 9770 1795
rect 9750 1765 9800 1775
rect 9750 1745 9770 1765
rect 9790 1745 9800 1765
rect 9750 1740 9800 1745
rect 9750 1655 9770 1740
rect 9825 1715 9845 1795
rect 9800 1705 9845 1715
rect 9800 1685 9810 1705
rect 9830 1685 9845 1705
rect 9800 1675 9845 1685
rect 9905 1710 9925 1795
rect 9905 1700 9945 1710
rect 9905 1680 9915 1700
rect 9935 1680 9945 1700
rect 9905 1670 9945 1680
rect 9905 1655 9925 1670
rect 9975 1655 9995 1795
rect 10040 1715 10060 1795
rect 10040 1705 10755 1715
rect 10040 1695 10355 1705
rect 10040 1655 10060 1695
rect 10185 1655 10205 1695
rect 10345 1685 10355 1695
rect 10375 1695 10755 1705
rect 10375 1685 10385 1695
rect 10345 1675 10385 1685
rect 8950 1645 8990 1655
rect 8950 1575 8960 1645
rect 8980 1575 8990 1645
rect 8950 1565 8990 1575
rect 9015 1645 9055 1655
rect 9015 1575 9025 1645
rect 9045 1575 9055 1645
rect 9015 1565 9055 1575
rect 9095 1645 9135 1655
rect 9095 1575 9105 1645
rect 9125 1575 9135 1645
rect 9095 1565 9135 1575
rect 9160 1645 9200 1655
rect 9160 1575 9170 1645
rect 9190 1575 9200 1645
rect 9160 1565 9200 1575
rect 9240 1645 9280 1655
rect 9240 1575 9250 1645
rect 9270 1575 9280 1645
rect 9240 1565 9280 1575
rect 9305 1645 9345 1655
rect 9305 1575 9315 1645
rect 9335 1575 9345 1645
rect 9305 1565 9345 1575
rect 9385 1645 9425 1655
rect 9385 1575 9395 1645
rect 9415 1575 9425 1645
rect 9385 1565 9425 1575
rect 9450 1645 9490 1655
rect 9450 1575 9460 1645
rect 9480 1575 9490 1645
rect 9450 1565 9490 1575
rect 9530 1645 9570 1655
rect 9530 1575 9540 1645
rect 9560 1575 9570 1645
rect 9530 1565 9570 1575
rect 9595 1645 9635 1655
rect 9595 1575 9605 1645
rect 9625 1575 9635 1645
rect 9595 1565 9635 1575
rect 9675 1645 9715 1655
rect 9675 1575 9685 1645
rect 9705 1575 9715 1645
rect 9675 1565 9715 1575
rect 9740 1645 9780 1655
rect 9740 1575 9750 1645
rect 9770 1575 9780 1645
rect 9740 1565 9780 1575
rect 9820 1645 9860 1655
rect 9820 1575 9830 1645
rect 9850 1575 9860 1645
rect 9820 1565 9860 1575
rect 9885 1645 9925 1655
rect 9885 1575 9895 1645
rect 9915 1575 9925 1645
rect 9885 1565 9925 1575
rect 9965 1645 10005 1655
rect 9965 1575 9975 1645
rect 9995 1575 10005 1645
rect 9965 1565 10005 1575
rect 10030 1645 10075 1655
rect 10030 1575 10040 1645
rect 10060 1575 10075 1645
rect 10030 1565 10075 1575
rect 10110 1645 10150 1655
rect 10110 1575 10120 1645
rect 10140 1575 10150 1645
rect 10110 1565 10150 1575
rect 10175 1645 10215 1655
rect 10175 1575 10185 1645
rect 10205 1575 10215 1645
rect 10175 1565 10215 1575
rect 10255 1645 10295 1655
rect 10255 1575 10265 1645
rect 10285 1575 10295 1645
rect 10255 1565 10295 1575
rect 8730 1525 9485 1545
rect 9975 1530 9995 1565
rect 8795 1450 8835 1460
rect 8795 1430 8805 1450
rect 8825 1430 8835 1450
rect 8795 1420 8835 1430
rect 9015 1450 9055 1460
rect 9015 1430 9025 1450
rect 9045 1430 9055 1450
rect 9015 1420 9055 1430
rect 9235 1450 9275 1460
rect 9235 1430 9245 1450
rect 9265 1430 9275 1450
rect 9235 1420 9275 1430
rect 8805 1400 8825 1420
rect 9025 1400 9045 1420
rect 9245 1400 9265 1420
rect 9465 1400 9485 1525
rect 9820 1510 9995 1530
rect 10025 1535 10065 1545
rect 10025 1515 10035 1535
rect 10055 1525 10065 1535
rect 10055 1515 10715 1525
rect 9820 1480 9840 1510
rect 10025 1505 10715 1515
rect 9800 1470 9840 1480
rect 9800 1450 9810 1470
rect 9830 1450 9840 1470
rect 9800 1440 9840 1450
rect 10635 1445 10675 1455
rect 10635 1425 10645 1445
rect 10665 1425 10675 1445
rect 10635 1415 10675 1425
rect 9685 1400 9705 1405
rect 10635 1400 10655 1415
rect 8795 1390 8835 1400
rect 8795 1320 8805 1390
rect 8825 1320 8835 1390
rect 8795 1310 8835 1320
rect 8905 1390 8945 1400
rect 8905 1320 8915 1390
rect 8935 1320 8945 1390
rect 8905 1310 8945 1320
rect 9015 1390 9055 1400
rect 9015 1320 9025 1390
rect 9045 1320 9055 1390
rect 9015 1310 9055 1320
rect 9125 1390 9165 1400
rect 9125 1320 9135 1390
rect 9155 1320 9165 1390
rect 9125 1310 9165 1320
rect 9235 1390 9275 1400
rect 9235 1320 9245 1390
rect 9265 1320 9275 1390
rect 9235 1310 9275 1320
rect 9455 1390 9495 1400
rect 9455 1320 9465 1390
rect 9485 1320 9495 1390
rect 9455 1310 9495 1320
rect 9565 1390 9605 1400
rect 9565 1320 9575 1390
rect 9595 1320 9605 1390
rect 9565 1310 9605 1320
rect 9675 1390 9715 1400
rect 9675 1320 9685 1390
rect 9705 1320 9715 1390
rect 9675 1310 9715 1320
rect 9785 1390 9825 1400
rect 9785 1320 9795 1390
rect 9815 1320 9825 1390
rect 9785 1310 9825 1320
rect 9895 1390 9935 1400
rect 9895 1320 9905 1390
rect 9925 1320 9935 1390
rect 9895 1310 9935 1320
rect 10175 1390 10215 1400
rect 10175 1320 10185 1390
rect 10205 1320 10215 1390
rect 10175 1310 10215 1320
rect 10285 1390 10325 1400
rect 10285 1320 10295 1390
rect 10315 1320 10325 1390
rect 10285 1310 10325 1320
rect 10395 1390 10435 1400
rect 10395 1320 10405 1390
rect 10425 1320 10435 1390
rect 10395 1310 10435 1320
rect 10505 1390 10545 1400
rect 10505 1320 10515 1390
rect 10535 1320 10545 1390
rect 10505 1310 10545 1320
rect 10615 1390 10655 1400
rect 10615 1320 10625 1390
rect 10645 1320 10655 1390
rect 10615 1310 10655 1320
rect 8805 1290 8825 1310
rect 9025 1290 9045 1310
rect 9245 1290 9265 1310
rect 8655 1270 9265 1290
rect 9465 1290 9485 1310
rect 9685 1290 9705 1310
rect 9905 1290 9925 1310
rect 9465 1270 9925 1290
rect 10185 1290 10205 1310
rect 10405 1290 10425 1310
rect 10625 1290 10645 1310
rect 10185 1270 10645 1290
rect 10695 930 10715 1505
rect 9465 910 10715 930
rect 9465 770 9490 910
rect 10735 890 10755 1695
rect 9435 760 9490 770
rect 9435 725 9445 760
rect 9480 725 9490 760
rect 9435 715 9490 725
rect 9655 870 10755 890
rect 9655 770 9675 870
rect 10775 850 10795 2005
rect 9965 830 10795 850
rect 9965 770 9985 830
rect 10815 810 10835 2140
rect 9655 760 9710 770
rect 9655 725 9665 760
rect 9700 725 9710 760
rect 9655 715 9710 725
rect 9860 760 9985 770
rect 9860 725 9870 760
rect 9905 750 9985 760
rect 10100 790 10835 810
rect 10100 770 10120 790
rect 10100 760 10295 770
rect 10100 750 10250 760
rect 9905 725 9915 750
rect 9860 715 9915 725
rect 10240 725 10250 750
rect 10285 725 10295 760
rect 10240 715 10295 725
<< viali >>
rect 8895 2250 8915 2320
rect 9115 2250 9135 2320
rect 9335 2250 9355 2320
rect 9555 2250 9575 2320
rect 9855 2250 9875 2320
rect 10075 2250 10095 2320
rect 10295 2250 10315 2320
rect 10515 2250 10535 2320
rect 8960 1805 8980 1975
rect 9105 1805 9125 1975
rect 9250 1805 9270 1975
rect 9605 1805 9625 1975
rect 9830 1805 9850 1975
rect 10120 1805 10140 1975
rect 10265 1805 10285 1975
rect 8960 1575 8980 1645
rect 9105 1575 9125 1645
rect 9250 1575 9270 1645
rect 9605 1575 9625 1645
rect 9830 1575 9850 1645
rect 10120 1575 10140 1645
rect 10265 1575 10285 1645
rect 8915 1320 8935 1390
rect 9135 1320 9155 1390
rect 9575 1320 9595 1390
rect 9795 1320 9815 1390
rect 10295 1320 10315 1390
rect 10515 1320 10535 1390
rect 9445 725 9480 760
rect 9665 725 9700 760
rect 9870 725 9905 760
rect 10250 725 10285 760
<< metal1 >>
rect 8775 2320 10885 2425
rect 8775 2250 8895 2320
rect 8915 2250 9115 2320
rect 9135 2250 9335 2320
rect 9355 2250 9555 2320
rect 9575 2250 9855 2320
rect 9875 2250 10075 2320
rect 10095 2250 10295 2320
rect 10315 2250 10515 2320
rect 10535 2250 10885 2320
rect 8775 1975 10885 2250
rect 8775 1805 8960 1975
rect 8980 1805 9105 1975
rect 9125 1805 9250 1975
rect 9270 1805 9605 1975
rect 9625 1805 9830 1975
rect 9850 1805 10120 1975
rect 10140 1805 10265 1975
rect 10285 1805 10885 1975
rect 8775 1790 10885 1805
rect 8775 1645 10885 1660
rect 8775 1575 8960 1645
rect 8980 1575 9105 1645
rect 9125 1575 9250 1645
rect 9270 1575 9605 1645
rect 9625 1575 9830 1645
rect 9850 1575 10120 1645
rect 10140 1575 10265 1645
rect 10285 1575 10885 1645
rect 8775 1390 10885 1575
rect 8775 1320 8915 1390
rect 8935 1320 9135 1390
rect 9155 1320 9575 1390
rect 9595 1320 9795 1390
rect 9815 1320 10295 1390
rect 10315 1320 10515 1390
rect 10535 1320 10885 1390
rect 8775 1305 10885 1320
rect 9435 760 9490 770
rect 9435 725 9445 760
rect 9480 725 9490 760
rect 9435 715 9490 725
rect 9655 760 9710 770
rect 9655 725 9665 760
rect 9700 725 9710 760
rect 9655 715 9710 725
rect 9860 760 9915 770
rect 9860 725 9870 760
rect 9905 725 9915 760
rect 9860 715 9915 725
rect 10240 760 10295 770
rect 10240 725 10250 760
rect 10285 725 10295 760
rect 10240 715 10295 725
<< via1 >>
rect 9445 725 9480 760
rect 9665 725 9700 760
rect 9870 725 9905 760
rect 10250 725 10285 760
<< metal2 >>
rect 9435 760 9490 770
rect 9435 725 9445 760
rect 9480 725 9490 760
rect 9435 715 9490 725
rect 9655 760 9710 770
rect 9655 725 9665 760
rect 9700 725 9710 760
rect 9655 715 9710 725
rect 9860 760 9915 770
rect 9860 725 9870 760
rect 9905 725 9915 760
rect 9860 715 9915 725
rect 10240 760 10295 770
rect 10240 725 10250 760
rect 10285 725 10295 760
rect 10240 715 10295 725
<< via2 >>
rect 9445 725 9480 760
rect 9665 725 9700 760
rect 9870 725 9905 760
rect 10250 725 10285 760
<< metal3 >>
rect 9435 760 9490 770
rect 9435 725 9445 760
rect 9480 725 9490 760
rect 9435 595 9490 725
rect 9655 760 9710 770
rect 9655 725 9665 760
rect 9700 725 9710 760
rect 9655 715 9710 725
rect 9860 760 9915 770
rect 9860 725 9870 760
rect 9905 725 9915 760
rect 9860 715 9915 725
rect 10240 760 10295 770
rect 10240 725 10250 760
rect 10285 725 10295 760
rect 10240 595 10295 725
rect 9435 305 9725 595
rect 9845 -35 10295 595
<< via3 >>
rect 9665 725 9700 760
rect 9870 725 9905 760
<< mimcap >>
rect 9450 570 9710 580
rect 9450 535 9665 570
rect 9700 535 9710 570
rect 9450 320 9710 535
rect 9860 570 10280 580
rect 9860 535 9870 570
rect 9905 535 10280 570
rect 9860 -20 10280 535
<< mimcapcontact >>
rect 9665 535 9700 570
rect 9870 535 9905 570
<< metal4 >>
rect 9655 760 9710 770
rect 9655 725 9665 760
rect 9700 725 9710 760
rect 9655 570 9710 725
rect 9655 535 9665 570
rect 9700 535 9710 570
rect 9655 525 9710 535
rect 9860 760 9915 770
rect 9860 725 9870 760
rect 9905 725 9915 760
rect 9860 570 9915 725
rect 9860 535 9870 570
rect 9905 535 9915 570
rect 9860 525 9915 535
<< labels >>
flabel poly 8630 1730 8630 1730 7 FreeSans 400 0 -200 0 UP_PFD
flabel poly 8630 1510 8630 1510 7 FreeSans 400 0 -200 0 DOWN_PFD
flabel locali 8655 1280 8655 1280 7 FreeSans 400 0 -200 0 I_IN
flabel locali 9425 2120 9425 2120 2 FreeSans 400 0 120 120 OPAMP_out
<< end >>
