magic
tech sky130A
timestamp 1751624208
<< nwell >>
rect 56075 4295 56435 4595
rect 56750 4295 57110 4850
rect 57420 4295 57780 4890
rect 54885 3575 55785 4155
rect 55935 3575 56835 4155
rect 56965 3575 57865 4155
rect 58015 3575 58915 4155
rect 54885 2615 55725 3445
rect 56205 3165 57595 3445
rect 55995 2710 56835 2990
rect 56965 2705 57805 2990
rect 58075 2615 58915 3445
rect 54885 2055 55725 2485
rect 58075 2055 58915 2485
<< pwell >>
rect 54480 3365 54770 3370
rect 54480 3345 54585 3365
rect 54665 3345 54770 3365
rect 54480 2635 54770 3345
rect 59030 3365 59320 3370
rect 59030 3345 59135 3365
rect 59215 3345 59320 3365
rect 59030 2635 59320 3345
rect 54395 1510 54760 2305
rect 56490 2310 57320 2565
rect 54900 1510 55710 2010
rect 56020 1930 56830 2280
rect 56970 2125 57780 2280
rect 56965 2085 57780 2125
rect 56970 1930 57780 2085
rect 59405 2395 59425 2415
rect 59235 2305 59275 2320
rect 55975 1460 57825 1810
rect 58090 1510 58900 2010
rect 59040 1510 59405 2305
rect 54650 498 54905 1385
rect 54980 520 55730 1430
rect 56150 835 57655 1320
rect 56650 530 57145 795
rect 58070 510 58820 1430
rect 58425 505 58465 510
rect 58900 500 59150 1385
<< nmos >>
rect 56590 2410 56605 2460
rect 56645 2410 56660 2460
rect 56700 2410 56715 2460
rect 56755 2410 56770 2460
rect 56810 2410 56825 2460
rect 56865 2410 56880 2460
rect 56920 2410 56935 2460
rect 56975 2410 56990 2460
rect 57030 2410 57045 2460
rect 57085 2410 57100 2460
rect 57140 2410 57155 2460
rect 57195 2410 57210 2460
rect 54995 1610 55010 1910
rect 55050 1610 55065 1910
rect 55105 1610 55120 1910
rect 55160 1610 55175 1910
rect 55215 1610 55230 1910
rect 55270 1610 55285 1910
rect 55325 1610 55340 1910
rect 55380 1610 55395 1910
rect 55435 1610 55450 1910
rect 55490 1610 55505 1910
rect 55545 1610 55560 1910
rect 55600 1610 55615 1910
rect 56115 2030 56130 2180
rect 56170 2030 56185 2180
rect 56225 2030 56240 2180
rect 56280 2030 56295 2180
rect 56335 2030 56350 2180
rect 56390 2030 56405 2180
rect 56445 2030 56460 2180
rect 56500 2030 56515 2180
rect 56555 2030 56570 2180
rect 56610 2030 56625 2180
rect 56665 2030 56680 2180
rect 56720 2030 56735 2180
rect 57065 2030 57080 2180
rect 57120 2030 57135 2180
rect 57175 2030 57190 2180
rect 57230 2030 57245 2180
rect 57285 2030 57300 2180
rect 57340 2030 57355 2180
rect 57395 2030 57410 2180
rect 57450 2030 57465 2180
rect 57505 2030 57520 2180
rect 57560 2030 57575 2180
rect 57615 2030 57630 2180
rect 57670 2030 57685 2180
rect 56070 1560 56085 1710
rect 56125 1560 56140 1710
rect 56180 1560 56195 1710
rect 56235 1560 56250 1710
rect 56290 1560 56305 1710
rect 56345 1560 56360 1710
rect 56400 1560 56415 1710
rect 56455 1560 56470 1710
rect 56510 1560 56525 1710
rect 56565 1560 56580 1710
rect 56620 1560 56635 1710
rect 56675 1560 56690 1710
rect 56810 1560 56825 1710
rect 56865 1560 56880 1710
rect 56920 1560 56935 1710
rect 56975 1560 56990 1710
rect 57110 1560 57125 1710
rect 57165 1560 57180 1710
rect 57220 1560 57235 1710
rect 57275 1560 57290 1710
rect 57330 1560 57345 1710
rect 57385 1560 57400 1710
rect 57440 1560 57455 1710
rect 57495 1560 57510 1710
rect 57550 1560 57565 1710
rect 57605 1560 57620 1710
rect 57660 1560 57675 1710
rect 57715 1560 57730 1710
rect 58185 1610 58200 1910
rect 58240 1610 58255 1910
rect 58295 1610 58310 1910
rect 58350 1610 58365 1910
rect 58405 1610 58420 1910
rect 58460 1610 58475 1910
rect 58515 1610 58530 1910
rect 58570 1610 58585 1910
rect 58625 1610 58640 1910
rect 58680 1610 58695 1910
rect 58735 1610 58750 1910
rect 58790 1610 58805 1910
rect 55075 620 55135 1320
rect 55175 620 55235 1320
rect 55275 620 55335 1320
rect 55375 620 55435 1320
rect 55475 620 55535 1320
rect 55575 620 55635 1320
rect 56260 955 56275 1205
rect 56315 955 56330 1205
rect 56370 955 56385 1205
rect 56425 955 56440 1205
rect 56480 955 56495 1205
rect 56535 955 56550 1205
rect 56590 955 56605 1205
rect 56645 955 56660 1205
rect 56700 955 56715 1205
rect 56755 955 56770 1205
rect 56810 955 56825 1205
rect 56865 955 56880 1205
rect 56920 955 56935 1205
rect 56975 955 56990 1205
rect 57030 955 57045 1205
rect 57085 955 57100 1205
rect 57140 955 57155 1205
rect 57195 955 57210 1205
rect 57250 955 57265 1205
rect 57305 955 57320 1205
rect 57360 955 57375 1205
rect 57415 955 57430 1205
rect 57470 955 57485 1205
rect 57525 955 57540 1205
rect 56750 590 57040 690
rect 58165 620 58225 1320
rect 58265 620 58325 1320
rect 58365 620 58425 1320
rect 58465 620 58525 1320
rect 58565 620 58625 1320
rect 58665 620 58725 1320
<< pmos >>
rect 56185 4415 56205 4478
rect 56245 4415 56265 4478
rect 56305 4415 56325 4478
rect 56860 4415 56880 4735
rect 56920 4415 56940 4735
rect 56980 4415 57000 4735
rect 57530 4415 57550 4775
rect 57590 4415 57610 4775
rect 57650 4415 57670 4775
rect 54995 3690 55015 4040
rect 55055 3690 55075 4040
rect 55115 3690 55135 4040
rect 55175 3690 55195 4040
rect 55235 3690 55255 4040
rect 55295 3690 55315 4040
rect 55355 3690 55375 4040
rect 55415 3690 55435 4040
rect 55475 3690 55495 4040
rect 55535 3690 55555 4040
rect 55595 3690 55615 4040
rect 55655 3690 55675 4040
rect 56045 3690 56065 4040
rect 56105 3690 56125 4040
rect 56165 3690 56185 4040
rect 56225 3690 56245 4040
rect 56285 3690 56305 4040
rect 56345 3690 56365 4040
rect 56405 3690 56425 4040
rect 56465 3690 56485 4040
rect 56525 3690 56545 4040
rect 56585 3690 56605 4040
rect 56645 3690 56665 4040
rect 56705 3690 56725 4040
rect 57075 3690 57095 4040
rect 57135 3690 57155 4040
rect 57195 3690 57215 4040
rect 57255 3690 57275 4040
rect 57315 3690 57335 4040
rect 57375 3690 57395 4040
rect 57435 3690 57455 4040
rect 57495 3690 57515 4040
rect 57555 3690 57575 4040
rect 57615 3690 57635 4040
rect 57675 3690 57695 4040
rect 57735 3690 57755 4040
rect 58125 3690 58145 4040
rect 58185 3690 58205 4040
rect 58245 3690 58265 4040
rect 58305 3690 58325 4040
rect 58365 3690 58385 4040
rect 58425 3690 58445 4040
rect 58485 3690 58505 4040
rect 58545 3690 58565 4040
rect 58605 3690 58625 4040
rect 58665 3690 58685 4040
rect 58725 3690 58745 4040
rect 58785 3690 58805 4040
rect 54995 2730 55010 3330
rect 55050 2730 55065 3330
rect 55105 2730 55120 3330
rect 55160 2730 55175 3330
rect 55215 2730 55230 3330
rect 55270 2730 55285 3330
rect 55325 2730 55340 3330
rect 55380 2730 55395 3330
rect 55435 2730 55450 3330
rect 55490 2730 55505 3330
rect 55545 2730 55560 3330
rect 55600 2730 55615 3330
rect 56315 3280 56330 3330
rect 56370 3280 56385 3330
rect 56425 3280 56440 3330
rect 56480 3280 56495 3330
rect 56535 3280 56550 3330
rect 56590 3280 56605 3330
rect 56645 3280 56660 3330
rect 56700 3280 56715 3330
rect 56755 3280 56770 3330
rect 56810 3280 56825 3330
rect 56865 3280 56880 3330
rect 56920 3280 56935 3330
rect 56975 3280 56990 3330
rect 57030 3280 57045 3330
rect 57085 3280 57100 3330
rect 57140 3280 57155 3330
rect 57195 3280 57210 3330
rect 57250 3280 57265 3330
rect 57305 3280 57320 3330
rect 57360 3280 57375 3330
rect 57415 3280 57430 3330
rect 57470 3280 57485 3330
rect 56105 2825 56120 2875
rect 56160 2825 56175 2875
rect 56215 2825 56230 2875
rect 56270 2825 56285 2875
rect 56325 2825 56340 2875
rect 56380 2825 56395 2875
rect 56435 2825 56450 2875
rect 56490 2825 56505 2875
rect 56545 2825 56560 2875
rect 56600 2825 56615 2875
rect 56655 2825 56670 2875
rect 56710 2825 56725 2875
rect 57075 2825 57090 2875
rect 57130 2825 57145 2875
rect 57185 2825 57200 2875
rect 57240 2825 57255 2875
rect 57295 2825 57310 2875
rect 57350 2825 57365 2875
rect 57405 2825 57420 2875
rect 57460 2825 57475 2875
rect 57515 2825 57530 2875
rect 57570 2825 57585 2875
rect 57625 2825 57640 2875
rect 57680 2825 57695 2875
rect 58185 2730 58200 3330
rect 58240 2730 58255 3330
rect 58295 2730 58310 3330
rect 58350 2730 58365 3330
rect 58405 2730 58420 3330
rect 58460 2730 58475 3330
rect 58515 2730 58530 3330
rect 58570 2730 58585 3330
rect 58625 2730 58640 3330
rect 58680 2730 58695 3330
rect 58735 2730 58750 3330
rect 58790 2730 58805 3330
rect 54995 2170 55010 2370
rect 55050 2170 55065 2370
rect 55105 2170 55120 2370
rect 55160 2170 55175 2370
rect 55215 2170 55230 2370
rect 55270 2170 55285 2370
rect 55325 2170 55340 2370
rect 55380 2170 55395 2370
rect 55435 2170 55450 2370
rect 55490 2170 55505 2370
rect 55545 2170 55560 2370
rect 55600 2170 55615 2370
rect 58185 2170 58200 2370
rect 58240 2170 58255 2370
rect 58295 2170 58310 2370
rect 58350 2170 58365 2370
rect 58405 2170 58420 2370
rect 58460 2170 58475 2370
rect 58515 2170 58530 2370
rect 58570 2170 58585 2370
rect 58625 2170 58640 2370
rect 58680 2170 58695 2370
rect 58735 2170 58750 2370
rect 58790 2170 58805 2370
<< ndiff >>
rect 56550 2445 56590 2460
rect 56550 2425 56560 2445
rect 56580 2425 56590 2445
rect 56550 2410 56590 2425
rect 56605 2445 56645 2460
rect 56605 2425 56615 2445
rect 56635 2425 56645 2445
rect 56605 2410 56645 2425
rect 56660 2445 56700 2460
rect 56660 2425 56670 2445
rect 56690 2425 56700 2445
rect 56660 2410 56700 2425
rect 56715 2445 56755 2460
rect 56715 2425 56725 2445
rect 56745 2425 56755 2445
rect 56715 2410 56755 2425
rect 56770 2445 56810 2460
rect 56770 2425 56780 2445
rect 56800 2425 56810 2445
rect 56770 2410 56810 2425
rect 56825 2445 56865 2460
rect 56825 2425 56835 2445
rect 56855 2425 56865 2445
rect 56825 2410 56865 2425
rect 56880 2445 56920 2460
rect 56880 2425 56890 2445
rect 56910 2425 56920 2445
rect 56880 2410 56920 2425
rect 56935 2445 56975 2460
rect 56935 2425 56945 2445
rect 56965 2425 56975 2445
rect 56935 2410 56975 2425
rect 56990 2445 57030 2460
rect 56990 2425 57000 2445
rect 57020 2425 57030 2445
rect 56990 2410 57030 2425
rect 57045 2445 57085 2460
rect 57045 2425 57055 2445
rect 57075 2425 57085 2445
rect 57045 2410 57085 2425
rect 57100 2445 57140 2460
rect 57100 2425 57110 2445
rect 57130 2425 57140 2445
rect 57100 2410 57140 2425
rect 57155 2445 57195 2460
rect 57155 2425 57165 2445
rect 57185 2425 57195 2445
rect 57155 2410 57195 2425
rect 57210 2445 57250 2460
rect 57210 2425 57220 2445
rect 57240 2425 57250 2445
rect 57210 2410 57250 2425
rect 54955 1895 54995 1910
rect 54955 1875 54965 1895
rect 54985 1875 54995 1895
rect 54955 1845 54995 1875
rect 54955 1825 54965 1845
rect 54985 1825 54995 1845
rect 54955 1795 54995 1825
rect 54955 1775 54965 1795
rect 54985 1775 54995 1795
rect 54955 1745 54995 1775
rect 54955 1725 54965 1745
rect 54985 1725 54995 1745
rect 54955 1695 54995 1725
rect 54955 1675 54965 1695
rect 54985 1675 54995 1695
rect 54955 1645 54995 1675
rect 54955 1625 54965 1645
rect 54985 1625 54995 1645
rect 54955 1610 54995 1625
rect 55010 1895 55050 1910
rect 55010 1875 55020 1895
rect 55040 1875 55050 1895
rect 55010 1845 55050 1875
rect 55010 1825 55020 1845
rect 55040 1825 55050 1845
rect 55010 1795 55050 1825
rect 55010 1775 55020 1795
rect 55040 1775 55050 1795
rect 55010 1745 55050 1775
rect 55010 1725 55020 1745
rect 55040 1725 55050 1745
rect 55010 1695 55050 1725
rect 55010 1675 55020 1695
rect 55040 1675 55050 1695
rect 55010 1645 55050 1675
rect 55010 1625 55020 1645
rect 55040 1625 55050 1645
rect 55010 1610 55050 1625
rect 55065 1895 55105 1910
rect 55065 1875 55075 1895
rect 55095 1875 55105 1895
rect 55065 1845 55105 1875
rect 55065 1825 55075 1845
rect 55095 1825 55105 1845
rect 55065 1795 55105 1825
rect 55065 1775 55075 1795
rect 55095 1775 55105 1795
rect 55065 1745 55105 1775
rect 55065 1725 55075 1745
rect 55095 1725 55105 1745
rect 55065 1695 55105 1725
rect 55065 1675 55075 1695
rect 55095 1675 55105 1695
rect 55065 1645 55105 1675
rect 55065 1625 55075 1645
rect 55095 1625 55105 1645
rect 55065 1610 55105 1625
rect 55120 1895 55160 1910
rect 55120 1875 55130 1895
rect 55150 1875 55160 1895
rect 55120 1845 55160 1875
rect 55120 1825 55130 1845
rect 55150 1825 55160 1845
rect 55120 1795 55160 1825
rect 55120 1775 55130 1795
rect 55150 1775 55160 1795
rect 55120 1745 55160 1775
rect 55120 1725 55130 1745
rect 55150 1725 55160 1745
rect 55120 1695 55160 1725
rect 55120 1675 55130 1695
rect 55150 1675 55160 1695
rect 55120 1645 55160 1675
rect 55120 1625 55130 1645
rect 55150 1625 55160 1645
rect 55120 1610 55160 1625
rect 55175 1895 55215 1910
rect 55175 1875 55185 1895
rect 55205 1875 55215 1895
rect 55175 1845 55215 1875
rect 55175 1825 55185 1845
rect 55205 1825 55215 1845
rect 55175 1795 55215 1825
rect 55175 1775 55185 1795
rect 55205 1775 55215 1795
rect 55175 1745 55215 1775
rect 55175 1725 55185 1745
rect 55205 1725 55215 1745
rect 55175 1695 55215 1725
rect 55175 1675 55185 1695
rect 55205 1675 55215 1695
rect 55175 1645 55215 1675
rect 55175 1625 55185 1645
rect 55205 1625 55215 1645
rect 55175 1610 55215 1625
rect 55230 1895 55270 1910
rect 55230 1875 55240 1895
rect 55260 1875 55270 1895
rect 55230 1845 55270 1875
rect 55230 1825 55240 1845
rect 55260 1825 55270 1845
rect 55230 1795 55270 1825
rect 55230 1775 55240 1795
rect 55260 1775 55270 1795
rect 55230 1745 55270 1775
rect 55230 1725 55240 1745
rect 55260 1725 55270 1745
rect 55230 1695 55270 1725
rect 55230 1675 55240 1695
rect 55260 1675 55270 1695
rect 55230 1645 55270 1675
rect 55230 1625 55240 1645
rect 55260 1625 55270 1645
rect 55230 1610 55270 1625
rect 55285 1895 55325 1910
rect 55285 1875 55295 1895
rect 55315 1875 55325 1895
rect 55285 1845 55325 1875
rect 55285 1825 55295 1845
rect 55315 1825 55325 1845
rect 55285 1795 55325 1825
rect 55285 1775 55295 1795
rect 55315 1775 55325 1795
rect 55285 1745 55325 1775
rect 55285 1725 55295 1745
rect 55315 1725 55325 1745
rect 55285 1695 55325 1725
rect 55285 1675 55295 1695
rect 55315 1675 55325 1695
rect 55285 1645 55325 1675
rect 55285 1625 55295 1645
rect 55315 1625 55325 1645
rect 55285 1610 55325 1625
rect 55340 1895 55380 1910
rect 55340 1875 55350 1895
rect 55370 1875 55380 1895
rect 55340 1845 55380 1875
rect 55340 1825 55350 1845
rect 55370 1825 55380 1845
rect 55340 1795 55380 1825
rect 55340 1775 55350 1795
rect 55370 1775 55380 1795
rect 55340 1745 55380 1775
rect 55340 1725 55350 1745
rect 55370 1725 55380 1745
rect 55340 1695 55380 1725
rect 55340 1675 55350 1695
rect 55370 1675 55380 1695
rect 55340 1645 55380 1675
rect 55340 1625 55350 1645
rect 55370 1625 55380 1645
rect 55340 1610 55380 1625
rect 55395 1895 55435 1910
rect 55395 1875 55405 1895
rect 55425 1875 55435 1895
rect 55395 1845 55435 1875
rect 55395 1825 55405 1845
rect 55425 1825 55435 1845
rect 55395 1795 55435 1825
rect 55395 1775 55405 1795
rect 55425 1775 55435 1795
rect 55395 1745 55435 1775
rect 55395 1725 55405 1745
rect 55425 1725 55435 1745
rect 55395 1695 55435 1725
rect 55395 1675 55405 1695
rect 55425 1675 55435 1695
rect 55395 1645 55435 1675
rect 55395 1625 55405 1645
rect 55425 1625 55435 1645
rect 55395 1610 55435 1625
rect 55450 1895 55490 1910
rect 55450 1875 55460 1895
rect 55480 1875 55490 1895
rect 55450 1845 55490 1875
rect 55450 1825 55460 1845
rect 55480 1825 55490 1845
rect 55450 1795 55490 1825
rect 55450 1775 55460 1795
rect 55480 1775 55490 1795
rect 55450 1745 55490 1775
rect 55450 1725 55460 1745
rect 55480 1725 55490 1745
rect 55450 1695 55490 1725
rect 55450 1675 55460 1695
rect 55480 1675 55490 1695
rect 55450 1645 55490 1675
rect 55450 1625 55460 1645
rect 55480 1625 55490 1645
rect 55450 1610 55490 1625
rect 55505 1895 55545 1910
rect 55505 1875 55515 1895
rect 55535 1875 55545 1895
rect 55505 1845 55545 1875
rect 55505 1825 55515 1845
rect 55535 1825 55545 1845
rect 55505 1795 55545 1825
rect 55505 1775 55515 1795
rect 55535 1775 55545 1795
rect 55505 1745 55545 1775
rect 55505 1725 55515 1745
rect 55535 1725 55545 1745
rect 55505 1695 55545 1725
rect 55505 1675 55515 1695
rect 55535 1675 55545 1695
rect 55505 1645 55545 1675
rect 55505 1625 55515 1645
rect 55535 1625 55545 1645
rect 55505 1610 55545 1625
rect 55560 1895 55600 1910
rect 55560 1875 55570 1895
rect 55590 1875 55600 1895
rect 55560 1845 55600 1875
rect 55560 1825 55570 1845
rect 55590 1825 55600 1845
rect 55560 1795 55600 1825
rect 55560 1775 55570 1795
rect 55590 1775 55600 1795
rect 55560 1745 55600 1775
rect 55560 1725 55570 1745
rect 55590 1725 55600 1745
rect 55560 1695 55600 1725
rect 55560 1675 55570 1695
rect 55590 1675 55600 1695
rect 55560 1645 55600 1675
rect 55560 1625 55570 1645
rect 55590 1625 55600 1645
rect 55560 1610 55600 1625
rect 55615 1895 55655 1910
rect 55615 1875 55625 1895
rect 55645 1875 55655 1895
rect 55615 1845 55655 1875
rect 55615 1825 55625 1845
rect 55645 1825 55655 1845
rect 55615 1795 55655 1825
rect 55615 1775 55625 1795
rect 55645 1775 55655 1795
rect 55615 1745 55655 1775
rect 55615 1725 55625 1745
rect 55645 1725 55655 1745
rect 55615 1695 55655 1725
rect 55615 1675 55625 1695
rect 55645 1675 55655 1695
rect 55615 1645 55655 1675
rect 55615 1625 55625 1645
rect 55645 1625 55655 1645
rect 55615 1610 55655 1625
rect 56075 2165 56115 2180
rect 56075 2145 56085 2165
rect 56105 2145 56115 2165
rect 56075 2115 56115 2145
rect 56075 2095 56085 2115
rect 56105 2095 56115 2115
rect 56075 2065 56115 2095
rect 56075 2045 56085 2065
rect 56105 2045 56115 2065
rect 56075 2030 56115 2045
rect 56130 2165 56170 2180
rect 56130 2145 56140 2165
rect 56160 2145 56170 2165
rect 56130 2115 56170 2145
rect 56130 2095 56140 2115
rect 56160 2095 56170 2115
rect 56130 2065 56170 2095
rect 56130 2045 56140 2065
rect 56160 2045 56170 2065
rect 56130 2030 56170 2045
rect 56185 2165 56225 2180
rect 56185 2145 56195 2165
rect 56215 2145 56225 2165
rect 56185 2115 56225 2145
rect 56185 2095 56195 2115
rect 56215 2095 56225 2115
rect 56185 2065 56225 2095
rect 56185 2045 56195 2065
rect 56215 2045 56225 2065
rect 56185 2030 56225 2045
rect 56240 2165 56280 2180
rect 56240 2145 56250 2165
rect 56270 2145 56280 2165
rect 56240 2115 56280 2145
rect 56240 2095 56250 2115
rect 56270 2095 56280 2115
rect 56240 2065 56280 2095
rect 56240 2045 56250 2065
rect 56270 2045 56280 2065
rect 56240 2030 56280 2045
rect 56295 2165 56335 2180
rect 56295 2145 56305 2165
rect 56325 2145 56335 2165
rect 56295 2115 56335 2145
rect 56295 2095 56305 2115
rect 56325 2095 56335 2115
rect 56295 2065 56335 2095
rect 56295 2045 56305 2065
rect 56325 2045 56335 2065
rect 56295 2030 56335 2045
rect 56350 2165 56390 2180
rect 56350 2145 56360 2165
rect 56380 2145 56390 2165
rect 56350 2115 56390 2145
rect 56350 2095 56360 2115
rect 56380 2095 56390 2115
rect 56350 2065 56390 2095
rect 56350 2045 56360 2065
rect 56380 2045 56390 2065
rect 56350 2030 56390 2045
rect 56405 2165 56445 2180
rect 56405 2145 56415 2165
rect 56435 2145 56445 2165
rect 56405 2115 56445 2145
rect 56405 2095 56415 2115
rect 56435 2095 56445 2115
rect 56405 2065 56445 2095
rect 56405 2045 56415 2065
rect 56435 2045 56445 2065
rect 56405 2030 56445 2045
rect 56460 2165 56500 2180
rect 56460 2145 56470 2165
rect 56490 2145 56500 2165
rect 56460 2115 56500 2145
rect 56460 2095 56470 2115
rect 56490 2095 56500 2115
rect 56460 2065 56500 2095
rect 56460 2045 56470 2065
rect 56490 2045 56500 2065
rect 56460 2030 56500 2045
rect 56515 2165 56555 2180
rect 56515 2145 56525 2165
rect 56545 2145 56555 2165
rect 56515 2115 56555 2145
rect 56515 2095 56525 2115
rect 56545 2095 56555 2115
rect 56515 2065 56555 2095
rect 56515 2045 56525 2065
rect 56545 2045 56555 2065
rect 56515 2030 56555 2045
rect 56570 2165 56610 2180
rect 56570 2145 56580 2165
rect 56600 2145 56610 2165
rect 56570 2115 56610 2145
rect 56570 2095 56580 2115
rect 56600 2095 56610 2115
rect 56570 2065 56610 2095
rect 56570 2045 56580 2065
rect 56600 2045 56610 2065
rect 56570 2030 56610 2045
rect 56625 2165 56665 2180
rect 56625 2145 56635 2165
rect 56655 2145 56665 2165
rect 56625 2115 56665 2145
rect 56625 2095 56635 2115
rect 56655 2095 56665 2115
rect 56625 2065 56665 2095
rect 56625 2045 56635 2065
rect 56655 2045 56665 2065
rect 56625 2030 56665 2045
rect 56680 2165 56720 2180
rect 56680 2145 56690 2165
rect 56710 2145 56720 2165
rect 56680 2115 56720 2145
rect 56680 2095 56690 2115
rect 56710 2095 56720 2115
rect 56680 2065 56720 2095
rect 56680 2045 56690 2065
rect 56710 2045 56720 2065
rect 56680 2030 56720 2045
rect 56735 2165 56775 2180
rect 56735 2145 56745 2165
rect 56765 2145 56775 2165
rect 56735 2115 56775 2145
rect 56735 2095 56745 2115
rect 56765 2095 56775 2115
rect 56735 2065 56775 2095
rect 56735 2045 56745 2065
rect 56765 2045 56775 2065
rect 56735 2030 56775 2045
rect 57025 2165 57065 2180
rect 57025 2145 57035 2165
rect 57055 2145 57065 2165
rect 57025 2115 57065 2145
rect 57025 2095 57035 2115
rect 57055 2095 57065 2115
rect 57025 2065 57065 2095
rect 57025 2045 57035 2065
rect 57055 2045 57065 2065
rect 57025 2030 57065 2045
rect 57080 2165 57120 2180
rect 57080 2145 57090 2165
rect 57110 2145 57120 2165
rect 57080 2115 57120 2145
rect 57080 2095 57090 2115
rect 57110 2095 57120 2115
rect 57080 2065 57120 2095
rect 57080 2045 57090 2065
rect 57110 2045 57120 2065
rect 57080 2030 57120 2045
rect 57135 2165 57175 2180
rect 57135 2145 57145 2165
rect 57165 2145 57175 2165
rect 57135 2115 57175 2145
rect 57135 2095 57145 2115
rect 57165 2095 57175 2115
rect 57135 2065 57175 2095
rect 57135 2045 57145 2065
rect 57165 2045 57175 2065
rect 57135 2030 57175 2045
rect 57190 2165 57230 2180
rect 57190 2145 57200 2165
rect 57220 2145 57230 2165
rect 57190 2115 57230 2145
rect 57190 2095 57200 2115
rect 57220 2095 57230 2115
rect 57190 2065 57230 2095
rect 57190 2045 57200 2065
rect 57220 2045 57230 2065
rect 57190 2030 57230 2045
rect 57245 2165 57285 2180
rect 57245 2145 57255 2165
rect 57275 2145 57285 2165
rect 57245 2115 57285 2145
rect 57245 2095 57255 2115
rect 57275 2095 57285 2115
rect 57245 2065 57285 2095
rect 57245 2045 57255 2065
rect 57275 2045 57285 2065
rect 57245 2030 57285 2045
rect 57300 2165 57340 2180
rect 57300 2145 57310 2165
rect 57330 2145 57340 2165
rect 57300 2115 57340 2145
rect 57300 2095 57310 2115
rect 57330 2095 57340 2115
rect 57300 2065 57340 2095
rect 57300 2045 57310 2065
rect 57330 2045 57340 2065
rect 57300 2030 57340 2045
rect 57355 2165 57395 2180
rect 57355 2145 57365 2165
rect 57385 2145 57395 2165
rect 57355 2115 57395 2145
rect 57355 2095 57365 2115
rect 57385 2095 57395 2115
rect 57355 2065 57395 2095
rect 57355 2045 57365 2065
rect 57385 2045 57395 2065
rect 57355 2030 57395 2045
rect 57410 2165 57450 2180
rect 57410 2145 57420 2165
rect 57440 2145 57450 2165
rect 57410 2115 57450 2145
rect 57410 2095 57420 2115
rect 57440 2095 57450 2115
rect 57410 2065 57450 2095
rect 57410 2045 57420 2065
rect 57440 2045 57450 2065
rect 57410 2030 57450 2045
rect 57465 2165 57505 2180
rect 57465 2145 57475 2165
rect 57495 2145 57505 2165
rect 57465 2115 57505 2145
rect 57465 2095 57475 2115
rect 57495 2095 57505 2115
rect 57465 2065 57505 2095
rect 57465 2045 57475 2065
rect 57495 2045 57505 2065
rect 57465 2030 57505 2045
rect 57520 2165 57560 2180
rect 57520 2145 57530 2165
rect 57550 2145 57560 2165
rect 57520 2115 57560 2145
rect 57520 2095 57530 2115
rect 57550 2095 57560 2115
rect 57520 2065 57560 2095
rect 57520 2045 57530 2065
rect 57550 2045 57560 2065
rect 57520 2030 57560 2045
rect 57575 2165 57615 2180
rect 57575 2145 57585 2165
rect 57605 2145 57615 2165
rect 57575 2115 57615 2145
rect 57575 2095 57585 2115
rect 57605 2095 57615 2115
rect 57575 2065 57615 2095
rect 57575 2045 57585 2065
rect 57605 2045 57615 2065
rect 57575 2030 57615 2045
rect 57630 2165 57670 2180
rect 57630 2145 57640 2165
rect 57660 2145 57670 2165
rect 57630 2115 57670 2145
rect 57630 2095 57640 2115
rect 57660 2095 57670 2115
rect 57630 2065 57670 2095
rect 57630 2045 57640 2065
rect 57660 2045 57670 2065
rect 57630 2030 57670 2045
rect 57685 2165 57725 2180
rect 57685 2145 57695 2165
rect 57715 2145 57725 2165
rect 57685 2115 57725 2145
rect 57685 2095 57695 2115
rect 57715 2095 57725 2115
rect 57685 2065 57725 2095
rect 57685 2045 57695 2065
rect 57715 2045 57725 2065
rect 57685 2030 57725 2045
rect 56030 1695 56070 1710
rect 56030 1675 56040 1695
rect 56060 1675 56070 1695
rect 56030 1645 56070 1675
rect 56030 1625 56040 1645
rect 56060 1625 56070 1645
rect 56030 1595 56070 1625
rect 56030 1575 56040 1595
rect 56060 1575 56070 1595
rect 56030 1560 56070 1575
rect 56085 1695 56125 1710
rect 56085 1675 56095 1695
rect 56115 1675 56125 1695
rect 56085 1645 56125 1675
rect 56085 1625 56095 1645
rect 56115 1625 56125 1645
rect 56085 1595 56125 1625
rect 56085 1575 56095 1595
rect 56115 1575 56125 1595
rect 56085 1560 56125 1575
rect 56140 1695 56180 1710
rect 56140 1675 56150 1695
rect 56170 1675 56180 1695
rect 56140 1645 56180 1675
rect 56140 1625 56150 1645
rect 56170 1625 56180 1645
rect 56140 1595 56180 1625
rect 56140 1575 56150 1595
rect 56170 1575 56180 1595
rect 56140 1560 56180 1575
rect 56195 1695 56235 1710
rect 56195 1675 56205 1695
rect 56225 1675 56235 1695
rect 56195 1645 56235 1675
rect 56195 1625 56205 1645
rect 56225 1625 56235 1645
rect 56195 1595 56235 1625
rect 56195 1575 56205 1595
rect 56225 1575 56235 1595
rect 56195 1560 56235 1575
rect 56250 1695 56290 1710
rect 56250 1675 56260 1695
rect 56280 1675 56290 1695
rect 56250 1645 56290 1675
rect 56250 1625 56260 1645
rect 56280 1625 56290 1645
rect 56250 1595 56290 1625
rect 56250 1575 56260 1595
rect 56280 1575 56290 1595
rect 56250 1560 56290 1575
rect 56305 1695 56345 1710
rect 56305 1675 56315 1695
rect 56335 1675 56345 1695
rect 56305 1645 56345 1675
rect 56305 1625 56315 1645
rect 56335 1625 56345 1645
rect 56305 1595 56345 1625
rect 56305 1575 56315 1595
rect 56335 1575 56345 1595
rect 56305 1560 56345 1575
rect 56360 1695 56400 1710
rect 56360 1675 56370 1695
rect 56390 1675 56400 1695
rect 56360 1645 56400 1675
rect 56360 1625 56370 1645
rect 56390 1625 56400 1645
rect 56360 1595 56400 1625
rect 56360 1575 56370 1595
rect 56390 1575 56400 1595
rect 56360 1560 56400 1575
rect 56415 1695 56455 1710
rect 56415 1675 56425 1695
rect 56445 1675 56455 1695
rect 56415 1645 56455 1675
rect 56415 1625 56425 1645
rect 56445 1625 56455 1645
rect 56415 1595 56455 1625
rect 56415 1575 56425 1595
rect 56445 1575 56455 1595
rect 56415 1560 56455 1575
rect 56470 1695 56510 1710
rect 56470 1675 56480 1695
rect 56500 1675 56510 1695
rect 56470 1645 56510 1675
rect 56470 1625 56480 1645
rect 56500 1625 56510 1645
rect 56470 1595 56510 1625
rect 56470 1575 56480 1595
rect 56500 1575 56510 1595
rect 56470 1560 56510 1575
rect 56525 1695 56565 1710
rect 56525 1675 56535 1695
rect 56555 1675 56565 1695
rect 56525 1645 56565 1675
rect 56525 1625 56535 1645
rect 56555 1625 56565 1645
rect 56525 1595 56565 1625
rect 56525 1575 56535 1595
rect 56555 1575 56565 1595
rect 56525 1560 56565 1575
rect 56580 1695 56620 1710
rect 56580 1675 56590 1695
rect 56610 1675 56620 1695
rect 56580 1645 56620 1675
rect 56580 1625 56590 1645
rect 56610 1625 56620 1645
rect 56580 1595 56620 1625
rect 56580 1575 56590 1595
rect 56610 1575 56620 1595
rect 56580 1560 56620 1575
rect 56635 1695 56675 1710
rect 56635 1675 56645 1695
rect 56665 1675 56675 1695
rect 56635 1645 56675 1675
rect 56635 1625 56645 1645
rect 56665 1625 56675 1645
rect 56635 1595 56675 1625
rect 56635 1575 56645 1595
rect 56665 1575 56675 1595
rect 56635 1560 56675 1575
rect 56690 1695 56730 1710
rect 56690 1675 56700 1695
rect 56720 1675 56730 1695
rect 56690 1645 56730 1675
rect 56690 1625 56700 1645
rect 56720 1625 56730 1645
rect 56690 1595 56730 1625
rect 56690 1575 56700 1595
rect 56720 1575 56730 1595
rect 56690 1560 56730 1575
rect 56770 1695 56810 1710
rect 56770 1675 56780 1695
rect 56800 1675 56810 1695
rect 56770 1645 56810 1675
rect 56770 1625 56780 1645
rect 56800 1625 56810 1645
rect 56770 1595 56810 1625
rect 56770 1575 56780 1595
rect 56800 1575 56810 1595
rect 56770 1560 56810 1575
rect 56825 1695 56865 1710
rect 56825 1675 56835 1695
rect 56855 1675 56865 1695
rect 56825 1645 56865 1675
rect 56825 1625 56835 1645
rect 56855 1625 56865 1645
rect 56825 1595 56865 1625
rect 56825 1575 56835 1595
rect 56855 1575 56865 1595
rect 56825 1560 56865 1575
rect 56880 1695 56920 1710
rect 56880 1675 56890 1695
rect 56910 1675 56920 1695
rect 56880 1645 56920 1675
rect 56880 1625 56890 1645
rect 56910 1625 56920 1645
rect 56880 1595 56920 1625
rect 56880 1575 56890 1595
rect 56910 1575 56920 1595
rect 56880 1560 56920 1575
rect 56935 1695 56975 1710
rect 56935 1675 56945 1695
rect 56965 1675 56975 1695
rect 56935 1645 56975 1675
rect 56935 1625 56945 1645
rect 56965 1625 56975 1645
rect 56935 1595 56975 1625
rect 56935 1575 56945 1595
rect 56965 1575 56975 1595
rect 56935 1560 56975 1575
rect 56990 1695 57030 1710
rect 56990 1675 57000 1695
rect 57020 1675 57030 1695
rect 56990 1645 57030 1675
rect 56990 1625 57000 1645
rect 57020 1625 57030 1645
rect 56990 1595 57030 1625
rect 56990 1575 57000 1595
rect 57020 1575 57030 1595
rect 56990 1560 57030 1575
rect 57070 1695 57110 1710
rect 57070 1675 57080 1695
rect 57100 1675 57110 1695
rect 57070 1645 57110 1675
rect 57070 1625 57080 1645
rect 57100 1625 57110 1645
rect 57070 1595 57110 1625
rect 57070 1575 57080 1595
rect 57100 1575 57110 1595
rect 57070 1560 57110 1575
rect 57125 1695 57165 1710
rect 57125 1675 57135 1695
rect 57155 1675 57165 1695
rect 57125 1645 57165 1675
rect 57125 1625 57135 1645
rect 57155 1625 57165 1645
rect 57125 1595 57165 1625
rect 57125 1575 57135 1595
rect 57155 1575 57165 1595
rect 57125 1560 57165 1575
rect 57180 1695 57220 1710
rect 57180 1675 57190 1695
rect 57210 1675 57220 1695
rect 57180 1645 57220 1675
rect 57180 1625 57190 1645
rect 57210 1625 57220 1645
rect 57180 1595 57220 1625
rect 57180 1575 57190 1595
rect 57210 1575 57220 1595
rect 57180 1560 57220 1575
rect 57235 1695 57275 1710
rect 57235 1675 57245 1695
rect 57265 1675 57275 1695
rect 57235 1645 57275 1675
rect 57235 1625 57245 1645
rect 57265 1625 57275 1645
rect 57235 1595 57275 1625
rect 57235 1575 57245 1595
rect 57265 1575 57275 1595
rect 57235 1560 57275 1575
rect 57290 1695 57330 1710
rect 57290 1675 57300 1695
rect 57320 1675 57330 1695
rect 57290 1645 57330 1675
rect 57290 1625 57300 1645
rect 57320 1625 57330 1645
rect 57290 1595 57330 1625
rect 57290 1575 57300 1595
rect 57320 1575 57330 1595
rect 57290 1560 57330 1575
rect 57345 1695 57385 1710
rect 57345 1675 57355 1695
rect 57375 1675 57385 1695
rect 57345 1645 57385 1675
rect 57345 1625 57355 1645
rect 57375 1625 57385 1645
rect 57345 1595 57385 1625
rect 57345 1575 57355 1595
rect 57375 1575 57385 1595
rect 57345 1560 57385 1575
rect 57400 1695 57440 1710
rect 57400 1675 57410 1695
rect 57430 1675 57440 1695
rect 57400 1645 57440 1675
rect 57400 1625 57410 1645
rect 57430 1625 57440 1645
rect 57400 1595 57440 1625
rect 57400 1575 57410 1595
rect 57430 1575 57440 1595
rect 57400 1560 57440 1575
rect 57455 1695 57495 1710
rect 57455 1675 57465 1695
rect 57485 1675 57495 1695
rect 57455 1645 57495 1675
rect 57455 1625 57465 1645
rect 57485 1625 57495 1645
rect 57455 1595 57495 1625
rect 57455 1575 57465 1595
rect 57485 1575 57495 1595
rect 57455 1560 57495 1575
rect 57510 1695 57550 1710
rect 57510 1675 57520 1695
rect 57540 1675 57550 1695
rect 57510 1645 57550 1675
rect 57510 1625 57520 1645
rect 57540 1625 57550 1645
rect 57510 1595 57550 1625
rect 57510 1575 57520 1595
rect 57540 1575 57550 1595
rect 57510 1560 57550 1575
rect 57565 1695 57605 1710
rect 57565 1675 57575 1695
rect 57595 1675 57605 1695
rect 57565 1645 57605 1675
rect 57565 1625 57575 1645
rect 57595 1625 57605 1645
rect 57565 1595 57605 1625
rect 57565 1575 57575 1595
rect 57595 1575 57605 1595
rect 57565 1560 57605 1575
rect 57620 1695 57660 1710
rect 57620 1675 57630 1695
rect 57650 1675 57660 1695
rect 57620 1645 57660 1675
rect 57620 1625 57630 1645
rect 57650 1625 57660 1645
rect 57620 1595 57660 1625
rect 57620 1575 57630 1595
rect 57650 1575 57660 1595
rect 57620 1560 57660 1575
rect 57675 1695 57715 1710
rect 57675 1675 57685 1695
rect 57705 1675 57715 1695
rect 57675 1645 57715 1675
rect 57675 1625 57685 1645
rect 57705 1625 57715 1645
rect 57675 1595 57715 1625
rect 57675 1575 57685 1595
rect 57705 1575 57715 1595
rect 57675 1560 57715 1575
rect 57730 1695 57770 1710
rect 57730 1675 57740 1695
rect 57760 1675 57770 1695
rect 57730 1645 57770 1675
rect 57730 1625 57740 1645
rect 57760 1625 57770 1645
rect 57730 1595 57770 1625
rect 57730 1575 57740 1595
rect 57760 1575 57770 1595
rect 57730 1560 57770 1575
rect 58145 1895 58185 1910
rect 58145 1875 58155 1895
rect 58175 1875 58185 1895
rect 58145 1845 58185 1875
rect 58145 1825 58155 1845
rect 58175 1825 58185 1845
rect 58145 1795 58185 1825
rect 58145 1775 58155 1795
rect 58175 1775 58185 1795
rect 58145 1745 58185 1775
rect 58145 1725 58155 1745
rect 58175 1725 58185 1745
rect 58145 1695 58185 1725
rect 58145 1675 58155 1695
rect 58175 1675 58185 1695
rect 58145 1645 58185 1675
rect 58145 1625 58155 1645
rect 58175 1625 58185 1645
rect 58145 1610 58185 1625
rect 58200 1895 58240 1910
rect 58200 1875 58210 1895
rect 58230 1875 58240 1895
rect 58200 1845 58240 1875
rect 58200 1825 58210 1845
rect 58230 1825 58240 1845
rect 58200 1795 58240 1825
rect 58200 1775 58210 1795
rect 58230 1775 58240 1795
rect 58200 1745 58240 1775
rect 58200 1725 58210 1745
rect 58230 1725 58240 1745
rect 58200 1695 58240 1725
rect 58200 1675 58210 1695
rect 58230 1675 58240 1695
rect 58200 1645 58240 1675
rect 58200 1625 58210 1645
rect 58230 1625 58240 1645
rect 58200 1610 58240 1625
rect 58255 1895 58295 1910
rect 58255 1875 58265 1895
rect 58285 1875 58295 1895
rect 58255 1845 58295 1875
rect 58255 1825 58265 1845
rect 58285 1825 58295 1845
rect 58255 1795 58295 1825
rect 58255 1775 58265 1795
rect 58285 1775 58295 1795
rect 58255 1745 58295 1775
rect 58255 1725 58265 1745
rect 58285 1725 58295 1745
rect 58255 1695 58295 1725
rect 58255 1675 58265 1695
rect 58285 1675 58295 1695
rect 58255 1645 58295 1675
rect 58255 1625 58265 1645
rect 58285 1625 58295 1645
rect 58255 1610 58295 1625
rect 58310 1895 58350 1910
rect 58310 1875 58320 1895
rect 58340 1875 58350 1895
rect 58310 1845 58350 1875
rect 58310 1825 58320 1845
rect 58340 1825 58350 1845
rect 58310 1795 58350 1825
rect 58310 1775 58320 1795
rect 58340 1775 58350 1795
rect 58310 1745 58350 1775
rect 58310 1725 58320 1745
rect 58340 1725 58350 1745
rect 58310 1695 58350 1725
rect 58310 1675 58320 1695
rect 58340 1675 58350 1695
rect 58310 1645 58350 1675
rect 58310 1625 58320 1645
rect 58340 1625 58350 1645
rect 58310 1610 58350 1625
rect 58365 1895 58405 1910
rect 58365 1875 58375 1895
rect 58395 1875 58405 1895
rect 58365 1845 58405 1875
rect 58365 1825 58375 1845
rect 58395 1825 58405 1845
rect 58365 1795 58405 1825
rect 58365 1775 58375 1795
rect 58395 1775 58405 1795
rect 58365 1745 58405 1775
rect 58365 1725 58375 1745
rect 58395 1725 58405 1745
rect 58365 1695 58405 1725
rect 58365 1675 58375 1695
rect 58395 1675 58405 1695
rect 58365 1645 58405 1675
rect 58365 1625 58375 1645
rect 58395 1625 58405 1645
rect 58365 1610 58405 1625
rect 58420 1895 58460 1910
rect 58420 1875 58430 1895
rect 58450 1875 58460 1895
rect 58420 1845 58460 1875
rect 58420 1825 58430 1845
rect 58450 1825 58460 1845
rect 58420 1795 58460 1825
rect 58420 1775 58430 1795
rect 58450 1775 58460 1795
rect 58420 1745 58460 1775
rect 58420 1725 58430 1745
rect 58450 1725 58460 1745
rect 58420 1695 58460 1725
rect 58420 1675 58430 1695
rect 58450 1675 58460 1695
rect 58420 1645 58460 1675
rect 58420 1625 58430 1645
rect 58450 1625 58460 1645
rect 58420 1610 58460 1625
rect 58475 1895 58515 1910
rect 58475 1875 58485 1895
rect 58505 1875 58515 1895
rect 58475 1845 58515 1875
rect 58475 1825 58485 1845
rect 58505 1825 58515 1845
rect 58475 1795 58515 1825
rect 58475 1775 58485 1795
rect 58505 1775 58515 1795
rect 58475 1745 58515 1775
rect 58475 1725 58485 1745
rect 58505 1725 58515 1745
rect 58475 1695 58515 1725
rect 58475 1675 58485 1695
rect 58505 1675 58515 1695
rect 58475 1645 58515 1675
rect 58475 1625 58485 1645
rect 58505 1625 58515 1645
rect 58475 1610 58515 1625
rect 58530 1895 58570 1910
rect 58530 1875 58540 1895
rect 58560 1875 58570 1895
rect 58530 1845 58570 1875
rect 58530 1825 58540 1845
rect 58560 1825 58570 1845
rect 58530 1795 58570 1825
rect 58530 1775 58540 1795
rect 58560 1775 58570 1795
rect 58530 1745 58570 1775
rect 58530 1725 58540 1745
rect 58560 1725 58570 1745
rect 58530 1695 58570 1725
rect 58530 1675 58540 1695
rect 58560 1675 58570 1695
rect 58530 1645 58570 1675
rect 58530 1625 58540 1645
rect 58560 1625 58570 1645
rect 58530 1610 58570 1625
rect 58585 1895 58625 1910
rect 58585 1875 58595 1895
rect 58615 1875 58625 1895
rect 58585 1845 58625 1875
rect 58585 1825 58595 1845
rect 58615 1825 58625 1845
rect 58585 1795 58625 1825
rect 58585 1775 58595 1795
rect 58615 1775 58625 1795
rect 58585 1745 58625 1775
rect 58585 1725 58595 1745
rect 58615 1725 58625 1745
rect 58585 1695 58625 1725
rect 58585 1675 58595 1695
rect 58615 1675 58625 1695
rect 58585 1645 58625 1675
rect 58585 1625 58595 1645
rect 58615 1625 58625 1645
rect 58585 1610 58625 1625
rect 58640 1895 58680 1910
rect 58640 1875 58650 1895
rect 58670 1875 58680 1895
rect 58640 1845 58680 1875
rect 58640 1825 58650 1845
rect 58670 1825 58680 1845
rect 58640 1795 58680 1825
rect 58640 1775 58650 1795
rect 58670 1775 58680 1795
rect 58640 1745 58680 1775
rect 58640 1725 58650 1745
rect 58670 1725 58680 1745
rect 58640 1695 58680 1725
rect 58640 1675 58650 1695
rect 58670 1675 58680 1695
rect 58640 1645 58680 1675
rect 58640 1625 58650 1645
rect 58670 1625 58680 1645
rect 58640 1610 58680 1625
rect 58695 1895 58735 1910
rect 58695 1875 58705 1895
rect 58725 1875 58735 1895
rect 58695 1845 58735 1875
rect 58695 1825 58705 1845
rect 58725 1825 58735 1845
rect 58695 1795 58735 1825
rect 58695 1775 58705 1795
rect 58725 1775 58735 1795
rect 58695 1745 58735 1775
rect 58695 1725 58705 1745
rect 58725 1725 58735 1745
rect 58695 1695 58735 1725
rect 58695 1675 58705 1695
rect 58725 1675 58735 1695
rect 58695 1645 58735 1675
rect 58695 1625 58705 1645
rect 58725 1625 58735 1645
rect 58695 1610 58735 1625
rect 58750 1895 58790 1910
rect 58750 1875 58760 1895
rect 58780 1875 58790 1895
rect 58750 1845 58790 1875
rect 58750 1825 58760 1845
rect 58780 1825 58790 1845
rect 58750 1795 58790 1825
rect 58750 1775 58760 1795
rect 58780 1775 58790 1795
rect 58750 1745 58790 1775
rect 58750 1725 58760 1745
rect 58780 1725 58790 1745
rect 58750 1695 58790 1725
rect 58750 1675 58760 1695
rect 58780 1675 58790 1695
rect 58750 1645 58790 1675
rect 58750 1625 58760 1645
rect 58780 1625 58790 1645
rect 58750 1610 58790 1625
rect 58805 1895 58845 1910
rect 58805 1875 58815 1895
rect 58835 1875 58845 1895
rect 58805 1845 58845 1875
rect 58805 1825 58815 1845
rect 58835 1825 58845 1845
rect 58805 1795 58845 1825
rect 58805 1775 58815 1795
rect 58835 1775 58845 1795
rect 58805 1745 58845 1775
rect 58805 1725 58815 1745
rect 58835 1725 58845 1745
rect 58805 1695 58845 1725
rect 58805 1675 58815 1695
rect 58835 1675 58845 1695
rect 58805 1645 58845 1675
rect 58805 1625 58815 1645
rect 58835 1625 58845 1645
rect 58805 1610 58845 1625
rect 55035 1305 55075 1320
rect 55035 1285 55045 1305
rect 55065 1285 55075 1305
rect 55035 1255 55075 1285
rect 55035 1235 55045 1255
rect 55065 1235 55075 1255
rect 55035 1205 55075 1235
rect 55035 1185 55045 1205
rect 55065 1185 55075 1205
rect 55035 1155 55075 1185
rect 55035 1135 55045 1155
rect 55065 1135 55075 1155
rect 55035 1105 55075 1135
rect 55035 1085 55045 1105
rect 55065 1085 55075 1105
rect 55035 1055 55075 1085
rect 55035 1035 55045 1055
rect 55065 1035 55075 1055
rect 55035 1005 55075 1035
rect 55035 985 55045 1005
rect 55065 985 55075 1005
rect 55035 955 55075 985
rect 55035 935 55045 955
rect 55065 935 55075 955
rect 55035 905 55075 935
rect 55035 885 55045 905
rect 55065 885 55075 905
rect 55035 855 55075 885
rect 55035 835 55045 855
rect 55065 835 55075 855
rect 55035 805 55075 835
rect 55035 785 55045 805
rect 55065 785 55075 805
rect 55035 755 55075 785
rect 55035 735 55045 755
rect 55065 735 55075 755
rect 55035 705 55075 735
rect 55035 685 55045 705
rect 55065 685 55075 705
rect 55035 655 55075 685
rect 55035 635 55045 655
rect 55065 635 55075 655
rect 55035 620 55075 635
rect 55135 1305 55175 1320
rect 55135 1285 55145 1305
rect 55165 1285 55175 1305
rect 55135 1255 55175 1285
rect 55135 1235 55145 1255
rect 55165 1235 55175 1255
rect 55135 1205 55175 1235
rect 55135 1185 55145 1205
rect 55165 1185 55175 1205
rect 55135 1155 55175 1185
rect 55135 1135 55145 1155
rect 55165 1135 55175 1155
rect 55135 1105 55175 1135
rect 55135 1085 55145 1105
rect 55165 1085 55175 1105
rect 55135 1055 55175 1085
rect 55135 1035 55145 1055
rect 55165 1035 55175 1055
rect 55135 1005 55175 1035
rect 55135 985 55145 1005
rect 55165 985 55175 1005
rect 55135 955 55175 985
rect 55135 935 55145 955
rect 55165 935 55175 955
rect 55135 905 55175 935
rect 55135 885 55145 905
rect 55165 885 55175 905
rect 55135 855 55175 885
rect 55135 835 55145 855
rect 55165 835 55175 855
rect 55135 805 55175 835
rect 55135 785 55145 805
rect 55165 785 55175 805
rect 55135 755 55175 785
rect 55135 735 55145 755
rect 55165 735 55175 755
rect 55135 705 55175 735
rect 55135 685 55145 705
rect 55165 685 55175 705
rect 55135 655 55175 685
rect 55135 635 55145 655
rect 55165 635 55175 655
rect 55135 620 55175 635
rect 55235 1305 55275 1320
rect 55235 1285 55245 1305
rect 55265 1285 55275 1305
rect 55235 1255 55275 1285
rect 55235 1235 55245 1255
rect 55265 1235 55275 1255
rect 55235 1205 55275 1235
rect 55235 1185 55245 1205
rect 55265 1185 55275 1205
rect 55235 1155 55275 1185
rect 55235 1135 55245 1155
rect 55265 1135 55275 1155
rect 55235 1105 55275 1135
rect 55235 1085 55245 1105
rect 55265 1085 55275 1105
rect 55235 1055 55275 1085
rect 55235 1035 55245 1055
rect 55265 1035 55275 1055
rect 55235 1005 55275 1035
rect 55235 985 55245 1005
rect 55265 985 55275 1005
rect 55235 955 55275 985
rect 55235 935 55245 955
rect 55265 935 55275 955
rect 55235 905 55275 935
rect 55235 885 55245 905
rect 55265 885 55275 905
rect 55235 855 55275 885
rect 55235 835 55245 855
rect 55265 835 55275 855
rect 55235 805 55275 835
rect 55235 785 55245 805
rect 55265 785 55275 805
rect 55235 755 55275 785
rect 55235 735 55245 755
rect 55265 735 55275 755
rect 55235 705 55275 735
rect 55235 685 55245 705
rect 55265 685 55275 705
rect 55235 655 55275 685
rect 55235 635 55245 655
rect 55265 635 55275 655
rect 55235 620 55275 635
rect 55335 1305 55375 1320
rect 55335 1285 55345 1305
rect 55365 1285 55375 1305
rect 55335 1255 55375 1285
rect 55335 1235 55345 1255
rect 55365 1235 55375 1255
rect 55335 1205 55375 1235
rect 55335 1185 55345 1205
rect 55365 1185 55375 1205
rect 55335 1155 55375 1185
rect 55335 1135 55345 1155
rect 55365 1135 55375 1155
rect 55335 1105 55375 1135
rect 55335 1085 55345 1105
rect 55365 1085 55375 1105
rect 55335 1055 55375 1085
rect 55335 1035 55345 1055
rect 55365 1035 55375 1055
rect 55335 1005 55375 1035
rect 55335 985 55345 1005
rect 55365 985 55375 1005
rect 55335 955 55375 985
rect 55335 935 55345 955
rect 55365 935 55375 955
rect 55335 905 55375 935
rect 55335 885 55345 905
rect 55365 885 55375 905
rect 55335 855 55375 885
rect 55335 835 55345 855
rect 55365 835 55375 855
rect 55335 805 55375 835
rect 55335 785 55345 805
rect 55365 785 55375 805
rect 55335 755 55375 785
rect 55335 735 55345 755
rect 55365 735 55375 755
rect 55335 705 55375 735
rect 55335 685 55345 705
rect 55365 685 55375 705
rect 55335 655 55375 685
rect 55335 635 55345 655
rect 55365 635 55375 655
rect 55335 620 55375 635
rect 55435 1305 55475 1320
rect 55435 1285 55445 1305
rect 55465 1285 55475 1305
rect 55435 1255 55475 1285
rect 55435 1235 55445 1255
rect 55465 1235 55475 1255
rect 55435 1205 55475 1235
rect 55435 1185 55445 1205
rect 55465 1185 55475 1205
rect 55435 1155 55475 1185
rect 55435 1135 55445 1155
rect 55465 1135 55475 1155
rect 55435 1105 55475 1135
rect 55435 1085 55445 1105
rect 55465 1085 55475 1105
rect 55435 1055 55475 1085
rect 55435 1035 55445 1055
rect 55465 1035 55475 1055
rect 55435 1005 55475 1035
rect 55435 985 55445 1005
rect 55465 985 55475 1005
rect 55435 955 55475 985
rect 55435 935 55445 955
rect 55465 935 55475 955
rect 55435 905 55475 935
rect 55435 885 55445 905
rect 55465 885 55475 905
rect 55435 855 55475 885
rect 55435 835 55445 855
rect 55465 835 55475 855
rect 55435 805 55475 835
rect 55435 785 55445 805
rect 55465 785 55475 805
rect 55435 755 55475 785
rect 55435 735 55445 755
rect 55465 735 55475 755
rect 55435 705 55475 735
rect 55435 685 55445 705
rect 55465 685 55475 705
rect 55435 655 55475 685
rect 55435 635 55445 655
rect 55465 635 55475 655
rect 55435 620 55475 635
rect 55535 1305 55575 1320
rect 55535 1285 55545 1305
rect 55565 1285 55575 1305
rect 55535 1255 55575 1285
rect 55535 1235 55545 1255
rect 55565 1235 55575 1255
rect 55535 1205 55575 1235
rect 55535 1185 55545 1205
rect 55565 1185 55575 1205
rect 55535 1155 55575 1185
rect 55535 1135 55545 1155
rect 55565 1135 55575 1155
rect 55535 1105 55575 1135
rect 55535 1085 55545 1105
rect 55565 1085 55575 1105
rect 55535 1055 55575 1085
rect 55535 1035 55545 1055
rect 55565 1035 55575 1055
rect 55535 1005 55575 1035
rect 55535 985 55545 1005
rect 55565 985 55575 1005
rect 55535 955 55575 985
rect 55535 935 55545 955
rect 55565 935 55575 955
rect 55535 905 55575 935
rect 55535 885 55545 905
rect 55565 885 55575 905
rect 55535 855 55575 885
rect 55535 835 55545 855
rect 55565 835 55575 855
rect 55535 805 55575 835
rect 55535 785 55545 805
rect 55565 785 55575 805
rect 55535 755 55575 785
rect 55535 735 55545 755
rect 55565 735 55575 755
rect 55535 705 55575 735
rect 55535 685 55545 705
rect 55565 685 55575 705
rect 55535 655 55575 685
rect 55535 635 55545 655
rect 55565 635 55575 655
rect 55535 620 55575 635
rect 55635 1305 55675 1320
rect 55635 1285 55645 1305
rect 55665 1285 55675 1305
rect 55635 1255 55675 1285
rect 55635 1235 55645 1255
rect 55665 1235 55675 1255
rect 55635 1205 55675 1235
rect 55635 1185 55645 1205
rect 55665 1185 55675 1205
rect 55635 1155 55675 1185
rect 55635 1135 55645 1155
rect 55665 1135 55675 1155
rect 55635 1105 55675 1135
rect 55635 1085 55645 1105
rect 55665 1085 55675 1105
rect 55635 1055 55675 1085
rect 55635 1035 55645 1055
rect 55665 1035 55675 1055
rect 55635 1005 55675 1035
rect 55635 985 55645 1005
rect 55665 985 55675 1005
rect 55635 955 55675 985
rect 55635 935 55645 955
rect 55665 935 55675 955
rect 55635 905 55675 935
rect 55635 885 55645 905
rect 55665 885 55675 905
rect 55635 855 55675 885
rect 55635 835 55645 855
rect 55665 835 55675 855
rect 55635 805 55675 835
rect 55635 785 55645 805
rect 55665 785 55675 805
rect 55635 755 55675 785
rect 55635 735 55645 755
rect 55665 735 55675 755
rect 55635 705 55675 735
rect 55635 685 55645 705
rect 55665 685 55675 705
rect 55635 655 55675 685
rect 55635 635 55645 655
rect 55665 635 55675 655
rect 55635 620 55675 635
rect 56220 1190 56260 1205
rect 56220 1170 56230 1190
rect 56250 1170 56260 1190
rect 56220 1140 56260 1170
rect 56220 1120 56230 1140
rect 56250 1120 56260 1140
rect 56220 1090 56260 1120
rect 56220 1070 56230 1090
rect 56250 1070 56260 1090
rect 56220 1040 56260 1070
rect 56220 1020 56230 1040
rect 56250 1020 56260 1040
rect 56220 990 56260 1020
rect 56220 970 56230 990
rect 56250 970 56260 990
rect 56220 955 56260 970
rect 56275 1190 56315 1205
rect 56275 1170 56285 1190
rect 56305 1170 56315 1190
rect 56275 1140 56315 1170
rect 56275 1120 56285 1140
rect 56305 1120 56315 1140
rect 56275 1090 56315 1120
rect 56275 1070 56285 1090
rect 56305 1070 56315 1090
rect 56275 1040 56315 1070
rect 56275 1020 56285 1040
rect 56305 1020 56315 1040
rect 56275 990 56315 1020
rect 56275 970 56285 990
rect 56305 970 56315 990
rect 56275 955 56315 970
rect 56330 1190 56370 1205
rect 56330 1170 56340 1190
rect 56360 1170 56370 1190
rect 56330 1140 56370 1170
rect 56330 1120 56340 1140
rect 56360 1120 56370 1140
rect 56330 1090 56370 1120
rect 56330 1070 56340 1090
rect 56360 1070 56370 1090
rect 56330 1040 56370 1070
rect 56330 1020 56340 1040
rect 56360 1020 56370 1040
rect 56330 990 56370 1020
rect 56330 970 56340 990
rect 56360 970 56370 990
rect 56330 955 56370 970
rect 56385 1190 56425 1205
rect 56385 1170 56395 1190
rect 56415 1170 56425 1190
rect 56385 1140 56425 1170
rect 56385 1120 56395 1140
rect 56415 1120 56425 1140
rect 56385 1090 56425 1120
rect 56385 1070 56395 1090
rect 56415 1070 56425 1090
rect 56385 1040 56425 1070
rect 56385 1020 56395 1040
rect 56415 1020 56425 1040
rect 56385 990 56425 1020
rect 56385 970 56395 990
rect 56415 970 56425 990
rect 56385 955 56425 970
rect 56440 1190 56480 1205
rect 56440 1170 56450 1190
rect 56470 1170 56480 1190
rect 56440 1140 56480 1170
rect 56440 1120 56450 1140
rect 56470 1120 56480 1140
rect 56440 1090 56480 1120
rect 56440 1070 56450 1090
rect 56470 1070 56480 1090
rect 56440 1040 56480 1070
rect 56440 1020 56450 1040
rect 56470 1020 56480 1040
rect 56440 990 56480 1020
rect 56440 970 56450 990
rect 56470 970 56480 990
rect 56440 955 56480 970
rect 56495 1190 56535 1205
rect 56495 1170 56505 1190
rect 56525 1170 56535 1190
rect 56495 1140 56535 1170
rect 56495 1120 56505 1140
rect 56525 1120 56535 1140
rect 56495 1090 56535 1120
rect 56495 1070 56505 1090
rect 56525 1070 56535 1090
rect 56495 1040 56535 1070
rect 56495 1020 56505 1040
rect 56525 1020 56535 1040
rect 56495 990 56535 1020
rect 56495 970 56505 990
rect 56525 970 56535 990
rect 56495 955 56535 970
rect 56550 1190 56590 1205
rect 56550 1170 56560 1190
rect 56580 1170 56590 1190
rect 56550 1140 56590 1170
rect 56550 1120 56560 1140
rect 56580 1120 56590 1140
rect 56550 1090 56590 1120
rect 56550 1070 56560 1090
rect 56580 1070 56590 1090
rect 56550 1040 56590 1070
rect 56550 1020 56560 1040
rect 56580 1020 56590 1040
rect 56550 990 56590 1020
rect 56550 970 56560 990
rect 56580 970 56590 990
rect 56550 955 56590 970
rect 56605 1190 56645 1205
rect 56605 1170 56615 1190
rect 56635 1170 56645 1190
rect 56605 1140 56645 1170
rect 56605 1120 56615 1140
rect 56635 1120 56645 1140
rect 56605 1090 56645 1120
rect 56605 1070 56615 1090
rect 56635 1070 56645 1090
rect 56605 1040 56645 1070
rect 56605 1020 56615 1040
rect 56635 1020 56645 1040
rect 56605 990 56645 1020
rect 56605 970 56615 990
rect 56635 970 56645 990
rect 56605 955 56645 970
rect 56660 1190 56700 1205
rect 56660 1170 56670 1190
rect 56690 1170 56700 1190
rect 56660 1140 56700 1170
rect 56660 1120 56670 1140
rect 56690 1120 56700 1140
rect 56660 1090 56700 1120
rect 56660 1070 56670 1090
rect 56690 1070 56700 1090
rect 56660 1040 56700 1070
rect 56660 1020 56670 1040
rect 56690 1020 56700 1040
rect 56660 990 56700 1020
rect 56660 970 56670 990
rect 56690 970 56700 990
rect 56660 955 56700 970
rect 56715 1190 56755 1205
rect 56715 1170 56725 1190
rect 56745 1170 56755 1190
rect 56715 1140 56755 1170
rect 56715 1120 56725 1140
rect 56745 1120 56755 1140
rect 56715 1090 56755 1120
rect 56715 1070 56725 1090
rect 56745 1070 56755 1090
rect 56715 1040 56755 1070
rect 56715 1020 56725 1040
rect 56745 1020 56755 1040
rect 56715 990 56755 1020
rect 56715 970 56725 990
rect 56745 970 56755 990
rect 56715 955 56755 970
rect 56770 1190 56810 1205
rect 56770 1170 56780 1190
rect 56800 1170 56810 1190
rect 56770 1140 56810 1170
rect 56770 1120 56780 1140
rect 56800 1120 56810 1140
rect 56770 1090 56810 1120
rect 56770 1070 56780 1090
rect 56800 1070 56810 1090
rect 56770 1040 56810 1070
rect 56770 1020 56780 1040
rect 56800 1020 56810 1040
rect 56770 990 56810 1020
rect 56770 970 56780 990
rect 56800 970 56810 990
rect 56770 955 56810 970
rect 56825 1190 56865 1205
rect 56825 1170 56835 1190
rect 56855 1170 56865 1190
rect 56825 1140 56865 1170
rect 56825 1120 56835 1140
rect 56855 1120 56865 1140
rect 56825 1090 56865 1120
rect 56825 1070 56835 1090
rect 56855 1070 56865 1090
rect 56825 1040 56865 1070
rect 56825 1020 56835 1040
rect 56855 1020 56865 1040
rect 56825 990 56865 1020
rect 56825 970 56835 990
rect 56855 970 56865 990
rect 56825 955 56865 970
rect 56880 1190 56920 1205
rect 56880 1170 56890 1190
rect 56910 1170 56920 1190
rect 56880 1140 56920 1170
rect 56880 1120 56890 1140
rect 56910 1120 56920 1140
rect 56880 1090 56920 1120
rect 56880 1070 56890 1090
rect 56910 1070 56920 1090
rect 56880 1040 56920 1070
rect 56880 1020 56890 1040
rect 56910 1020 56920 1040
rect 56880 990 56920 1020
rect 56880 970 56890 990
rect 56910 970 56920 990
rect 56880 955 56920 970
rect 56935 1190 56975 1205
rect 56935 1170 56945 1190
rect 56965 1170 56975 1190
rect 56935 1140 56975 1170
rect 56935 1120 56945 1140
rect 56965 1120 56975 1140
rect 56935 1090 56975 1120
rect 56935 1070 56945 1090
rect 56965 1070 56975 1090
rect 56935 1040 56975 1070
rect 56935 1020 56945 1040
rect 56965 1020 56975 1040
rect 56935 990 56975 1020
rect 56935 970 56945 990
rect 56965 970 56975 990
rect 56935 955 56975 970
rect 56990 1190 57030 1205
rect 56990 1170 57000 1190
rect 57020 1170 57030 1190
rect 56990 1140 57030 1170
rect 56990 1120 57000 1140
rect 57020 1120 57030 1140
rect 56990 1090 57030 1120
rect 56990 1070 57000 1090
rect 57020 1070 57030 1090
rect 56990 1040 57030 1070
rect 56990 1020 57000 1040
rect 57020 1020 57030 1040
rect 56990 990 57030 1020
rect 56990 970 57000 990
rect 57020 970 57030 990
rect 56990 955 57030 970
rect 57045 1190 57085 1205
rect 57045 1170 57055 1190
rect 57075 1170 57085 1190
rect 57045 1140 57085 1170
rect 57045 1120 57055 1140
rect 57075 1120 57085 1140
rect 57045 1090 57085 1120
rect 57045 1070 57055 1090
rect 57075 1070 57085 1090
rect 57045 1040 57085 1070
rect 57045 1020 57055 1040
rect 57075 1020 57085 1040
rect 57045 990 57085 1020
rect 57045 970 57055 990
rect 57075 970 57085 990
rect 57045 955 57085 970
rect 57100 1190 57140 1205
rect 57100 1170 57110 1190
rect 57130 1170 57140 1190
rect 57100 1140 57140 1170
rect 57100 1120 57110 1140
rect 57130 1120 57140 1140
rect 57100 1090 57140 1120
rect 57100 1070 57110 1090
rect 57130 1070 57140 1090
rect 57100 1040 57140 1070
rect 57100 1020 57110 1040
rect 57130 1020 57140 1040
rect 57100 990 57140 1020
rect 57100 970 57110 990
rect 57130 970 57140 990
rect 57100 955 57140 970
rect 57155 1190 57195 1205
rect 57155 1170 57165 1190
rect 57185 1170 57195 1190
rect 57155 1140 57195 1170
rect 57155 1120 57165 1140
rect 57185 1120 57195 1140
rect 57155 1090 57195 1120
rect 57155 1070 57165 1090
rect 57185 1070 57195 1090
rect 57155 1040 57195 1070
rect 57155 1020 57165 1040
rect 57185 1020 57195 1040
rect 57155 990 57195 1020
rect 57155 970 57165 990
rect 57185 970 57195 990
rect 57155 955 57195 970
rect 57210 1190 57250 1205
rect 57210 1170 57220 1190
rect 57240 1170 57250 1190
rect 57210 1140 57250 1170
rect 57210 1120 57220 1140
rect 57240 1120 57250 1140
rect 57210 1090 57250 1120
rect 57210 1070 57220 1090
rect 57240 1070 57250 1090
rect 57210 1040 57250 1070
rect 57210 1020 57220 1040
rect 57240 1020 57250 1040
rect 57210 990 57250 1020
rect 57210 970 57220 990
rect 57240 970 57250 990
rect 57210 955 57250 970
rect 57265 1190 57305 1205
rect 57265 1170 57275 1190
rect 57295 1170 57305 1190
rect 57265 1140 57305 1170
rect 57265 1120 57275 1140
rect 57295 1120 57305 1140
rect 57265 1090 57305 1120
rect 57265 1070 57275 1090
rect 57295 1070 57305 1090
rect 57265 1040 57305 1070
rect 57265 1020 57275 1040
rect 57295 1020 57305 1040
rect 57265 990 57305 1020
rect 57265 970 57275 990
rect 57295 970 57305 990
rect 57265 955 57305 970
rect 57320 1190 57360 1205
rect 57320 1170 57330 1190
rect 57350 1170 57360 1190
rect 57320 1140 57360 1170
rect 57320 1120 57330 1140
rect 57350 1120 57360 1140
rect 57320 1090 57360 1120
rect 57320 1070 57330 1090
rect 57350 1070 57360 1090
rect 57320 1040 57360 1070
rect 57320 1020 57330 1040
rect 57350 1020 57360 1040
rect 57320 990 57360 1020
rect 57320 970 57330 990
rect 57350 970 57360 990
rect 57320 955 57360 970
rect 57375 1190 57415 1205
rect 57375 1170 57385 1190
rect 57405 1170 57415 1190
rect 57375 1140 57415 1170
rect 57375 1120 57385 1140
rect 57405 1120 57415 1140
rect 57375 1090 57415 1120
rect 57375 1070 57385 1090
rect 57405 1070 57415 1090
rect 57375 1040 57415 1070
rect 57375 1020 57385 1040
rect 57405 1020 57415 1040
rect 57375 990 57415 1020
rect 57375 970 57385 990
rect 57405 970 57415 990
rect 57375 955 57415 970
rect 57430 1190 57470 1205
rect 57430 1170 57440 1190
rect 57460 1170 57470 1190
rect 57430 1140 57470 1170
rect 57430 1120 57440 1140
rect 57460 1120 57470 1140
rect 57430 1090 57470 1120
rect 57430 1070 57440 1090
rect 57460 1070 57470 1090
rect 57430 1040 57470 1070
rect 57430 1020 57440 1040
rect 57460 1020 57470 1040
rect 57430 990 57470 1020
rect 57430 970 57440 990
rect 57460 970 57470 990
rect 57430 955 57470 970
rect 57485 1190 57525 1205
rect 57485 1170 57495 1190
rect 57515 1170 57525 1190
rect 57485 1140 57525 1170
rect 57485 1120 57495 1140
rect 57515 1120 57525 1140
rect 57485 1090 57525 1120
rect 57485 1070 57495 1090
rect 57515 1070 57525 1090
rect 57485 1040 57525 1070
rect 57485 1020 57495 1040
rect 57515 1020 57525 1040
rect 57485 990 57525 1020
rect 57485 970 57495 990
rect 57515 970 57525 990
rect 57485 955 57525 970
rect 57540 1190 57580 1205
rect 57540 1170 57550 1190
rect 57570 1170 57580 1190
rect 57540 1140 57580 1170
rect 57540 1120 57550 1140
rect 57570 1120 57580 1140
rect 57540 1090 57580 1120
rect 57540 1070 57550 1090
rect 57570 1070 57580 1090
rect 57540 1040 57580 1070
rect 57540 1020 57550 1040
rect 57570 1020 57580 1040
rect 57540 990 57580 1020
rect 57540 970 57550 990
rect 57570 970 57580 990
rect 57540 955 57580 970
rect 56710 675 56750 690
rect 56710 655 56720 675
rect 56740 655 56750 675
rect 56710 625 56750 655
rect 56710 605 56720 625
rect 56740 605 56750 625
rect 56710 590 56750 605
rect 57040 675 57080 690
rect 57040 655 57050 675
rect 57070 655 57080 675
rect 57040 625 57080 655
rect 57040 605 57050 625
rect 57070 605 57080 625
rect 57040 590 57080 605
rect 58125 1305 58165 1320
rect 58125 1285 58135 1305
rect 58155 1285 58165 1305
rect 58125 1255 58165 1285
rect 58125 1235 58135 1255
rect 58155 1235 58165 1255
rect 58125 1205 58165 1235
rect 58125 1185 58135 1205
rect 58155 1185 58165 1205
rect 58125 1155 58165 1185
rect 58125 1135 58135 1155
rect 58155 1135 58165 1155
rect 58125 1105 58165 1135
rect 58125 1085 58135 1105
rect 58155 1085 58165 1105
rect 58125 1055 58165 1085
rect 58125 1035 58135 1055
rect 58155 1035 58165 1055
rect 58125 1005 58165 1035
rect 58125 985 58135 1005
rect 58155 985 58165 1005
rect 58125 955 58165 985
rect 58125 935 58135 955
rect 58155 935 58165 955
rect 58125 905 58165 935
rect 58125 885 58135 905
rect 58155 885 58165 905
rect 58125 855 58165 885
rect 58125 835 58135 855
rect 58155 835 58165 855
rect 58125 805 58165 835
rect 58125 785 58135 805
rect 58155 785 58165 805
rect 58125 755 58165 785
rect 58125 735 58135 755
rect 58155 735 58165 755
rect 58125 705 58165 735
rect 58125 685 58135 705
rect 58155 685 58165 705
rect 58125 655 58165 685
rect 58125 635 58135 655
rect 58155 635 58165 655
rect 58125 620 58165 635
rect 58225 1305 58265 1320
rect 58225 1285 58235 1305
rect 58255 1285 58265 1305
rect 58225 1255 58265 1285
rect 58225 1235 58235 1255
rect 58255 1235 58265 1255
rect 58225 1205 58265 1235
rect 58225 1185 58235 1205
rect 58255 1185 58265 1205
rect 58225 1155 58265 1185
rect 58225 1135 58235 1155
rect 58255 1135 58265 1155
rect 58225 1105 58265 1135
rect 58225 1085 58235 1105
rect 58255 1085 58265 1105
rect 58225 1055 58265 1085
rect 58225 1035 58235 1055
rect 58255 1035 58265 1055
rect 58225 1005 58265 1035
rect 58225 985 58235 1005
rect 58255 985 58265 1005
rect 58225 955 58265 985
rect 58225 935 58235 955
rect 58255 935 58265 955
rect 58225 905 58265 935
rect 58225 885 58235 905
rect 58255 885 58265 905
rect 58225 855 58265 885
rect 58225 835 58235 855
rect 58255 835 58265 855
rect 58225 805 58265 835
rect 58225 785 58235 805
rect 58255 785 58265 805
rect 58225 755 58265 785
rect 58225 735 58235 755
rect 58255 735 58265 755
rect 58225 705 58265 735
rect 58225 685 58235 705
rect 58255 685 58265 705
rect 58225 655 58265 685
rect 58225 635 58235 655
rect 58255 635 58265 655
rect 58225 620 58265 635
rect 58325 1305 58365 1320
rect 58325 1285 58335 1305
rect 58355 1285 58365 1305
rect 58325 1255 58365 1285
rect 58325 1235 58335 1255
rect 58355 1235 58365 1255
rect 58325 1205 58365 1235
rect 58325 1185 58335 1205
rect 58355 1185 58365 1205
rect 58325 1155 58365 1185
rect 58325 1135 58335 1155
rect 58355 1135 58365 1155
rect 58325 1105 58365 1135
rect 58325 1085 58335 1105
rect 58355 1085 58365 1105
rect 58325 1055 58365 1085
rect 58325 1035 58335 1055
rect 58355 1035 58365 1055
rect 58325 1005 58365 1035
rect 58325 985 58335 1005
rect 58355 985 58365 1005
rect 58325 955 58365 985
rect 58325 935 58335 955
rect 58355 935 58365 955
rect 58325 905 58365 935
rect 58325 885 58335 905
rect 58355 885 58365 905
rect 58325 855 58365 885
rect 58325 835 58335 855
rect 58355 835 58365 855
rect 58325 805 58365 835
rect 58325 785 58335 805
rect 58355 785 58365 805
rect 58325 755 58365 785
rect 58325 735 58335 755
rect 58355 735 58365 755
rect 58325 705 58365 735
rect 58325 685 58335 705
rect 58355 685 58365 705
rect 58325 655 58365 685
rect 58325 635 58335 655
rect 58355 635 58365 655
rect 58325 620 58365 635
rect 58425 1305 58465 1320
rect 58425 1285 58435 1305
rect 58455 1285 58465 1305
rect 58425 1255 58465 1285
rect 58425 1235 58435 1255
rect 58455 1235 58465 1255
rect 58425 1205 58465 1235
rect 58425 1185 58435 1205
rect 58455 1185 58465 1205
rect 58425 1155 58465 1185
rect 58425 1135 58435 1155
rect 58455 1135 58465 1155
rect 58425 1105 58465 1135
rect 58425 1085 58435 1105
rect 58455 1085 58465 1105
rect 58425 1055 58465 1085
rect 58425 1035 58435 1055
rect 58455 1035 58465 1055
rect 58425 1005 58465 1035
rect 58425 985 58435 1005
rect 58455 985 58465 1005
rect 58425 955 58465 985
rect 58425 935 58435 955
rect 58455 935 58465 955
rect 58425 905 58465 935
rect 58425 885 58435 905
rect 58455 885 58465 905
rect 58425 855 58465 885
rect 58425 835 58435 855
rect 58455 835 58465 855
rect 58425 805 58465 835
rect 58425 785 58435 805
rect 58455 785 58465 805
rect 58425 755 58465 785
rect 58425 735 58435 755
rect 58455 735 58465 755
rect 58425 705 58465 735
rect 58425 685 58435 705
rect 58455 685 58465 705
rect 58425 655 58465 685
rect 58425 635 58435 655
rect 58455 635 58465 655
rect 58425 620 58465 635
rect 58525 1305 58565 1320
rect 58525 1285 58535 1305
rect 58555 1285 58565 1305
rect 58525 1255 58565 1285
rect 58525 1235 58535 1255
rect 58555 1235 58565 1255
rect 58525 1205 58565 1235
rect 58525 1185 58535 1205
rect 58555 1185 58565 1205
rect 58525 1155 58565 1185
rect 58525 1135 58535 1155
rect 58555 1135 58565 1155
rect 58525 1105 58565 1135
rect 58525 1085 58535 1105
rect 58555 1085 58565 1105
rect 58525 1055 58565 1085
rect 58525 1035 58535 1055
rect 58555 1035 58565 1055
rect 58525 1005 58565 1035
rect 58525 985 58535 1005
rect 58555 985 58565 1005
rect 58525 955 58565 985
rect 58525 935 58535 955
rect 58555 935 58565 955
rect 58525 905 58565 935
rect 58525 885 58535 905
rect 58555 885 58565 905
rect 58525 855 58565 885
rect 58525 835 58535 855
rect 58555 835 58565 855
rect 58525 805 58565 835
rect 58525 785 58535 805
rect 58555 785 58565 805
rect 58525 755 58565 785
rect 58525 735 58535 755
rect 58555 735 58565 755
rect 58525 705 58565 735
rect 58525 685 58535 705
rect 58555 685 58565 705
rect 58525 655 58565 685
rect 58525 635 58535 655
rect 58555 635 58565 655
rect 58525 620 58565 635
rect 58625 1305 58665 1320
rect 58625 1285 58635 1305
rect 58655 1285 58665 1305
rect 58625 1255 58665 1285
rect 58625 1235 58635 1255
rect 58655 1235 58665 1255
rect 58625 1205 58665 1235
rect 58625 1185 58635 1205
rect 58655 1185 58665 1205
rect 58625 1155 58665 1185
rect 58625 1135 58635 1155
rect 58655 1135 58665 1155
rect 58625 1105 58665 1135
rect 58625 1085 58635 1105
rect 58655 1085 58665 1105
rect 58625 1055 58665 1085
rect 58625 1035 58635 1055
rect 58655 1035 58665 1055
rect 58625 1005 58665 1035
rect 58625 985 58635 1005
rect 58655 985 58665 1005
rect 58625 955 58665 985
rect 58625 935 58635 955
rect 58655 935 58665 955
rect 58625 905 58665 935
rect 58625 885 58635 905
rect 58655 885 58665 905
rect 58625 855 58665 885
rect 58625 835 58635 855
rect 58655 835 58665 855
rect 58625 805 58665 835
rect 58625 785 58635 805
rect 58655 785 58665 805
rect 58625 755 58665 785
rect 58625 735 58635 755
rect 58655 735 58665 755
rect 58625 705 58665 735
rect 58625 685 58635 705
rect 58655 685 58665 705
rect 58625 655 58665 685
rect 58625 635 58635 655
rect 58655 635 58665 655
rect 58625 620 58665 635
rect 58725 1305 58765 1320
rect 58725 1285 58735 1305
rect 58755 1285 58765 1305
rect 58725 1255 58765 1285
rect 58725 1235 58735 1255
rect 58755 1235 58765 1255
rect 58725 1205 58765 1235
rect 58725 1185 58735 1205
rect 58755 1185 58765 1205
rect 58725 1155 58765 1185
rect 58725 1135 58735 1155
rect 58755 1135 58765 1155
rect 58725 1105 58765 1135
rect 58725 1085 58735 1105
rect 58755 1085 58765 1105
rect 58725 1055 58765 1085
rect 58725 1035 58735 1055
rect 58755 1035 58765 1055
rect 58725 1005 58765 1035
rect 58725 985 58735 1005
rect 58755 985 58765 1005
rect 58725 955 58765 985
rect 58725 935 58735 955
rect 58755 935 58765 955
rect 58725 905 58765 935
rect 58725 885 58735 905
rect 58755 885 58765 905
rect 58725 855 58765 885
rect 58725 835 58735 855
rect 58755 835 58765 855
rect 58725 805 58765 835
rect 58725 785 58735 805
rect 58755 785 58765 805
rect 58725 755 58765 785
rect 58725 735 58735 755
rect 58755 735 58765 755
rect 58725 705 58765 735
rect 58725 685 58735 705
rect 58755 685 58765 705
rect 58725 655 58765 685
rect 58725 635 58735 655
rect 58755 635 58765 655
rect 58725 620 58765 635
<< pdiff >>
rect 56145 4450 56185 4478
rect 56145 4430 56155 4450
rect 56175 4430 56185 4450
rect 56145 4415 56185 4430
rect 56205 4450 56245 4478
rect 56205 4430 56215 4450
rect 56235 4430 56245 4450
rect 56205 4415 56245 4430
rect 56265 4450 56305 4478
rect 56265 4430 56275 4450
rect 56295 4430 56305 4450
rect 56265 4415 56305 4430
rect 56325 4450 56365 4478
rect 56325 4430 56335 4450
rect 56355 4430 56365 4450
rect 56325 4415 56365 4430
rect 56820 4705 56860 4735
rect 56820 4435 56830 4705
rect 56850 4435 56860 4705
rect 56820 4415 56860 4435
rect 56880 4705 56920 4735
rect 56880 4435 56890 4705
rect 56910 4435 56920 4705
rect 56880 4415 56920 4435
rect 56940 4705 56980 4735
rect 56940 4435 56950 4705
rect 56970 4435 56980 4705
rect 56940 4415 56980 4435
rect 57000 4705 57040 4735
rect 57000 4435 57010 4705
rect 57030 4435 57040 4705
rect 57000 4415 57040 4435
rect 57490 4745 57530 4775
rect 57490 4435 57500 4745
rect 57520 4435 57530 4745
rect 57490 4415 57530 4435
rect 57550 4745 57590 4775
rect 57550 4435 57560 4745
rect 57580 4435 57590 4745
rect 57550 4415 57590 4435
rect 57610 4745 57650 4775
rect 57610 4435 57620 4745
rect 57640 4435 57650 4745
rect 57610 4415 57650 4435
rect 57670 4745 57710 4775
rect 57670 4435 57680 4745
rect 57700 4435 57710 4745
rect 57670 4415 57710 4435
rect 54955 4025 54995 4040
rect 54955 4005 54965 4025
rect 54985 4005 54995 4025
rect 54955 3975 54995 4005
rect 54955 3955 54965 3975
rect 54985 3955 54995 3975
rect 54955 3925 54995 3955
rect 54955 3905 54965 3925
rect 54985 3905 54995 3925
rect 54955 3875 54995 3905
rect 54955 3855 54965 3875
rect 54985 3855 54995 3875
rect 54955 3825 54995 3855
rect 54955 3805 54965 3825
rect 54985 3805 54995 3825
rect 54955 3775 54995 3805
rect 54955 3755 54965 3775
rect 54985 3755 54995 3775
rect 54955 3725 54995 3755
rect 54955 3705 54965 3725
rect 54985 3705 54995 3725
rect 54955 3690 54995 3705
rect 55015 4025 55055 4040
rect 55015 4005 55025 4025
rect 55045 4005 55055 4025
rect 55015 3975 55055 4005
rect 55015 3955 55025 3975
rect 55045 3955 55055 3975
rect 55015 3925 55055 3955
rect 55015 3905 55025 3925
rect 55045 3905 55055 3925
rect 55015 3875 55055 3905
rect 55015 3855 55025 3875
rect 55045 3855 55055 3875
rect 55015 3825 55055 3855
rect 55015 3805 55025 3825
rect 55045 3805 55055 3825
rect 55015 3775 55055 3805
rect 55015 3755 55025 3775
rect 55045 3755 55055 3775
rect 55015 3725 55055 3755
rect 55015 3705 55025 3725
rect 55045 3705 55055 3725
rect 55015 3690 55055 3705
rect 55075 4025 55115 4040
rect 55075 4005 55085 4025
rect 55105 4005 55115 4025
rect 55075 3975 55115 4005
rect 55075 3955 55085 3975
rect 55105 3955 55115 3975
rect 55075 3925 55115 3955
rect 55075 3905 55085 3925
rect 55105 3905 55115 3925
rect 55075 3875 55115 3905
rect 55075 3855 55085 3875
rect 55105 3855 55115 3875
rect 55075 3825 55115 3855
rect 55075 3805 55085 3825
rect 55105 3805 55115 3825
rect 55075 3775 55115 3805
rect 55075 3755 55085 3775
rect 55105 3755 55115 3775
rect 55075 3725 55115 3755
rect 55075 3705 55085 3725
rect 55105 3705 55115 3725
rect 55075 3690 55115 3705
rect 55135 4025 55175 4040
rect 55135 4005 55145 4025
rect 55165 4005 55175 4025
rect 55135 3975 55175 4005
rect 55135 3955 55145 3975
rect 55165 3955 55175 3975
rect 55135 3925 55175 3955
rect 55135 3905 55145 3925
rect 55165 3905 55175 3925
rect 55135 3875 55175 3905
rect 55135 3855 55145 3875
rect 55165 3855 55175 3875
rect 55135 3825 55175 3855
rect 55135 3805 55145 3825
rect 55165 3805 55175 3825
rect 55135 3775 55175 3805
rect 55135 3755 55145 3775
rect 55165 3755 55175 3775
rect 55135 3725 55175 3755
rect 55135 3705 55145 3725
rect 55165 3705 55175 3725
rect 55135 3690 55175 3705
rect 55195 4025 55235 4040
rect 55195 4005 55205 4025
rect 55225 4005 55235 4025
rect 55195 3975 55235 4005
rect 55195 3955 55205 3975
rect 55225 3955 55235 3975
rect 55195 3925 55235 3955
rect 55195 3905 55205 3925
rect 55225 3905 55235 3925
rect 55195 3875 55235 3905
rect 55195 3855 55205 3875
rect 55225 3855 55235 3875
rect 55195 3825 55235 3855
rect 55195 3805 55205 3825
rect 55225 3805 55235 3825
rect 55195 3775 55235 3805
rect 55195 3755 55205 3775
rect 55225 3755 55235 3775
rect 55195 3725 55235 3755
rect 55195 3705 55205 3725
rect 55225 3705 55235 3725
rect 55195 3690 55235 3705
rect 55255 4025 55295 4040
rect 55255 4005 55265 4025
rect 55285 4005 55295 4025
rect 55255 3975 55295 4005
rect 55255 3955 55265 3975
rect 55285 3955 55295 3975
rect 55255 3925 55295 3955
rect 55255 3905 55265 3925
rect 55285 3905 55295 3925
rect 55255 3875 55295 3905
rect 55255 3855 55265 3875
rect 55285 3855 55295 3875
rect 55255 3825 55295 3855
rect 55255 3805 55265 3825
rect 55285 3805 55295 3825
rect 55255 3775 55295 3805
rect 55255 3755 55265 3775
rect 55285 3755 55295 3775
rect 55255 3725 55295 3755
rect 55255 3705 55265 3725
rect 55285 3705 55295 3725
rect 55255 3690 55295 3705
rect 55315 4025 55355 4040
rect 55315 4005 55325 4025
rect 55345 4005 55355 4025
rect 55315 3975 55355 4005
rect 55315 3955 55325 3975
rect 55345 3955 55355 3975
rect 55315 3925 55355 3955
rect 55315 3905 55325 3925
rect 55345 3905 55355 3925
rect 55315 3875 55355 3905
rect 55315 3855 55325 3875
rect 55345 3855 55355 3875
rect 55315 3825 55355 3855
rect 55315 3805 55325 3825
rect 55345 3805 55355 3825
rect 55315 3775 55355 3805
rect 55315 3755 55325 3775
rect 55345 3755 55355 3775
rect 55315 3725 55355 3755
rect 55315 3705 55325 3725
rect 55345 3705 55355 3725
rect 55315 3690 55355 3705
rect 55375 4025 55415 4040
rect 55375 4005 55385 4025
rect 55405 4005 55415 4025
rect 55375 3975 55415 4005
rect 55375 3955 55385 3975
rect 55405 3955 55415 3975
rect 55375 3925 55415 3955
rect 55375 3905 55385 3925
rect 55405 3905 55415 3925
rect 55375 3875 55415 3905
rect 55375 3855 55385 3875
rect 55405 3855 55415 3875
rect 55375 3825 55415 3855
rect 55375 3805 55385 3825
rect 55405 3805 55415 3825
rect 55375 3775 55415 3805
rect 55375 3755 55385 3775
rect 55405 3755 55415 3775
rect 55375 3725 55415 3755
rect 55375 3705 55385 3725
rect 55405 3705 55415 3725
rect 55375 3690 55415 3705
rect 55435 4025 55475 4040
rect 55435 4005 55445 4025
rect 55465 4005 55475 4025
rect 55435 3975 55475 4005
rect 55435 3955 55445 3975
rect 55465 3955 55475 3975
rect 55435 3925 55475 3955
rect 55435 3905 55445 3925
rect 55465 3905 55475 3925
rect 55435 3875 55475 3905
rect 55435 3855 55445 3875
rect 55465 3855 55475 3875
rect 55435 3825 55475 3855
rect 55435 3805 55445 3825
rect 55465 3805 55475 3825
rect 55435 3775 55475 3805
rect 55435 3755 55445 3775
rect 55465 3755 55475 3775
rect 55435 3725 55475 3755
rect 55435 3705 55445 3725
rect 55465 3705 55475 3725
rect 55435 3690 55475 3705
rect 55495 4025 55535 4040
rect 55495 4005 55505 4025
rect 55525 4005 55535 4025
rect 55495 3975 55535 4005
rect 55495 3955 55505 3975
rect 55525 3955 55535 3975
rect 55495 3925 55535 3955
rect 55495 3905 55505 3925
rect 55525 3905 55535 3925
rect 55495 3875 55535 3905
rect 55495 3855 55505 3875
rect 55525 3855 55535 3875
rect 55495 3825 55535 3855
rect 55495 3805 55505 3825
rect 55525 3805 55535 3825
rect 55495 3775 55535 3805
rect 55495 3755 55505 3775
rect 55525 3755 55535 3775
rect 55495 3725 55535 3755
rect 55495 3705 55505 3725
rect 55525 3705 55535 3725
rect 55495 3690 55535 3705
rect 55555 4025 55595 4040
rect 55555 4005 55565 4025
rect 55585 4005 55595 4025
rect 55555 3975 55595 4005
rect 55555 3955 55565 3975
rect 55585 3955 55595 3975
rect 55555 3925 55595 3955
rect 55555 3905 55565 3925
rect 55585 3905 55595 3925
rect 55555 3875 55595 3905
rect 55555 3855 55565 3875
rect 55585 3855 55595 3875
rect 55555 3825 55595 3855
rect 55555 3805 55565 3825
rect 55585 3805 55595 3825
rect 55555 3775 55595 3805
rect 55555 3755 55565 3775
rect 55585 3755 55595 3775
rect 55555 3725 55595 3755
rect 55555 3705 55565 3725
rect 55585 3705 55595 3725
rect 55555 3690 55595 3705
rect 55615 4025 55655 4040
rect 55615 4005 55625 4025
rect 55645 4005 55655 4025
rect 55615 3975 55655 4005
rect 55615 3955 55625 3975
rect 55645 3955 55655 3975
rect 55615 3925 55655 3955
rect 55615 3905 55625 3925
rect 55645 3905 55655 3925
rect 55615 3875 55655 3905
rect 55615 3855 55625 3875
rect 55645 3855 55655 3875
rect 55615 3825 55655 3855
rect 55615 3805 55625 3825
rect 55645 3805 55655 3825
rect 55615 3775 55655 3805
rect 55615 3755 55625 3775
rect 55645 3755 55655 3775
rect 55615 3725 55655 3755
rect 55615 3705 55625 3725
rect 55645 3705 55655 3725
rect 55615 3690 55655 3705
rect 55675 4025 55715 4040
rect 55675 4005 55685 4025
rect 55705 4005 55715 4025
rect 55675 3975 55715 4005
rect 55675 3955 55685 3975
rect 55705 3955 55715 3975
rect 55675 3925 55715 3955
rect 55675 3905 55685 3925
rect 55705 3905 55715 3925
rect 55675 3875 55715 3905
rect 55675 3855 55685 3875
rect 55705 3855 55715 3875
rect 55675 3825 55715 3855
rect 55675 3805 55685 3825
rect 55705 3805 55715 3825
rect 55675 3775 55715 3805
rect 55675 3755 55685 3775
rect 55705 3755 55715 3775
rect 55675 3725 55715 3755
rect 55675 3705 55685 3725
rect 55705 3705 55715 3725
rect 55675 3690 55715 3705
rect 56005 4025 56045 4040
rect 56005 4005 56015 4025
rect 56035 4005 56045 4025
rect 56005 3975 56045 4005
rect 56005 3955 56015 3975
rect 56035 3955 56045 3975
rect 56005 3925 56045 3955
rect 56005 3905 56015 3925
rect 56035 3905 56045 3925
rect 56005 3875 56045 3905
rect 56005 3855 56015 3875
rect 56035 3855 56045 3875
rect 56005 3825 56045 3855
rect 56005 3805 56015 3825
rect 56035 3805 56045 3825
rect 56005 3775 56045 3805
rect 56005 3755 56015 3775
rect 56035 3755 56045 3775
rect 56005 3725 56045 3755
rect 56005 3705 56015 3725
rect 56035 3705 56045 3725
rect 56005 3690 56045 3705
rect 56065 4025 56105 4040
rect 56065 4005 56075 4025
rect 56095 4005 56105 4025
rect 56065 3975 56105 4005
rect 56065 3955 56075 3975
rect 56095 3955 56105 3975
rect 56065 3925 56105 3955
rect 56065 3905 56075 3925
rect 56095 3905 56105 3925
rect 56065 3875 56105 3905
rect 56065 3855 56075 3875
rect 56095 3855 56105 3875
rect 56065 3825 56105 3855
rect 56065 3805 56075 3825
rect 56095 3805 56105 3825
rect 56065 3775 56105 3805
rect 56065 3755 56075 3775
rect 56095 3755 56105 3775
rect 56065 3725 56105 3755
rect 56065 3705 56075 3725
rect 56095 3705 56105 3725
rect 56065 3690 56105 3705
rect 56125 4025 56165 4040
rect 56125 4005 56135 4025
rect 56155 4005 56165 4025
rect 56125 3975 56165 4005
rect 56125 3955 56135 3975
rect 56155 3955 56165 3975
rect 56125 3925 56165 3955
rect 56125 3905 56135 3925
rect 56155 3905 56165 3925
rect 56125 3875 56165 3905
rect 56125 3855 56135 3875
rect 56155 3855 56165 3875
rect 56125 3825 56165 3855
rect 56125 3805 56135 3825
rect 56155 3805 56165 3825
rect 56125 3775 56165 3805
rect 56125 3755 56135 3775
rect 56155 3755 56165 3775
rect 56125 3725 56165 3755
rect 56125 3705 56135 3725
rect 56155 3705 56165 3725
rect 56125 3690 56165 3705
rect 56185 4025 56225 4040
rect 56185 4005 56195 4025
rect 56215 4005 56225 4025
rect 56185 3975 56225 4005
rect 56185 3955 56195 3975
rect 56215 3955 56225 3975
rect 56185 3925 56225 3955
rect 56185 3905 56195 3925
rect 56215 3905 56225 3925
rect 56185 3875 56225 3905
rect 56185 3855 56195 3875
rect 56215 3855 56225 3875
rect 56185 3825 56225 3855
rect 56185 3805 56195 3825
rect 56215 3805 56225 3825
rect 56185 3775 56225 3805
rect 56185 3755 56195 3775
rect 56215 3755 56225 3775
rect 56185 3725 56225 3755
rect 56185 3705 56195 3725
rect 56215 3705 56225 3725
rect 56185 3690 56225 3705
rect 56245 4025 56285 4040
rect 56245 4005 56255 4025
rect 56275 4005 56285 4025
rect 56245 3975 56285 4005
rect 56245 3955 56255 3975
rect 56275 3955 56285 3975
rect 56245 3925 56285 3955
rect 56245 3905 56255 3925
rect 56275 3905 56285 3925
rect 56245 3875 56285 3905
rect 56245 3855 56255 3875
rect 56275 3855 56285 3875
rect 56245 3825 56285 3855
rect 56245 3805 56255 3825
rect 56275 3805 56285 3825
rect 56245 3775 56285 3805
rect 56245 3755 56255 3775
rect 56275 3755 56285 3775
rect 56245 3725 56285 3755
rect 56245 3705 56255 3725
rect 56275 3705 56285 3725
rect 56245 3690 56285 3705
rect 56305 4025 56345 4040
rect 56305 4005 56315 4025
rect 56335 4005 56345 4025
rect 56305 3975 56345 4005
rect 56305 3955 56315 3975
rect 56335 3955 56345 3975
rect 56305 3925 56345 3955
rect 56305 3905 56315 3925
rect 56335 3905 56345 3925
rect 56305 3875 56345 3905
rect 56305 3855 56315 3875
rect 56335 3855 56345 3875
rect 56305 3825 56345 3855
rect 56305 3805 56315 3825
rect 56335 3805 56345 3825
rect 56305 3775 56345 3805
rect 56305 3755 56315 3775
rect 56335 3755 56345 3775
rect 56305 3725 56345 3755
rect 56305 3705 56315 3725
rect 56335 3705 56345 3725
rect 56305 3690 56345 3705
rect 56365 4025 56405 4040
rect 56365 4005 56375 4025
rect 56395 4005 56405 4025
rect 56365 3975 56405 4005
rect 56365 3955 56375 3975
rect 56395 3955 56405 3975
rect 56365 3925 56405 3955
rect 56365 3905 56375 3925
rect 56395 3905 56405 3925
rect 56365 3875 56405 3905
rect 56365 3855 56375 3875
rect 56395 3855 56405 3875
rect 56365 3825 56405 3855
rect 56365 3805 56375 3825
rect 56395 3805 56405 3825
rect 56365 3775 56405 3805
rect 56365 3755 56375 3775
rect 56395 3755 56405 3775
rect 56365 3725 56405 3755
rect 56365 3705 56375 3725
rect 56395 3705 56405 3725
rect 56365 3690 56405 3705
rect 56425 4025 56465 4040
rect 56425 4005 56435 4025
rect 56455 4005 56465 4025
rect 56425 3975 56465 4005
rect 56425 3955 56435 3975
rect 56455 3955 56465 3975
rect 56425 3925 56465 3955
rect 56425 3905 56435 3925
rect 56455 3905 56465 3925
rect 56425 3875 56465 3905
rect 56425 3855 56435 3875
rect 56455 3855 56465 3875
rect 56425 3825 56465 3855
rect 56425 3805 56435 3825
rect 56455 3805 56465 3825
rect 56425 3775 56465 3805
rect 56425 3755 56435 3775
rect 56455 3755 56465 3775
rect 56425 3725 56465 3755
rect 56425 3705 56435 3725
rect 56455 3705 56465 3725
rect 56425 3690 56465 3705
rect 56485 4025 56525 4040
rect 56485 4005 56495 4025
rect 56515 4005 56525 4025
rect 56485 3975 56525 4005
rect 56485 3955 56495 3975
rect 56515 3955 56525 3975
rect 56485 3925 56525 3955
rect 56485 3905 56495 3925
rect 56515 3905 56525 3925
rect 56485 3875 56525 3905
rect 56485 3855 56495 3875
rect 56515 3855 56525 3875
rect 56485 3825 56525 3855
rect 56485 3805 56495 3825
rect 56515 3805 56525 3825
rect 56485 3775 56525 3805
rect 56485 3755 56495 3775
rect 56515 3755 56525 3775
rect 56485 3725 56525 3755
rect 56485 3705 56495 3725
rect 56515 3705 56525 3725
rect 56485 3690 56525 3705
rect 56545 4025 56585 4040
rect 56545 4005 56555 4025
rect 56575 4005 56585 4025
rect 56545 3975 56585 4005
rect 56545 3955 56555 3975
rect 56575 3955 56585 3975
rect 56545 3925 56585 3955
rect 56545 3905 56555 3925
rect 56575 3905 56585 3925
rect 56545 3875 56585 3905
rect 56545 3855 56555 3875
rect 56575 3855 56585 3875
rect 56545 3825 56585 3855
rect 56545 3805 56555 3825
rect 56575 3805 56585 3825
rect 56545 3775 56585 3805
rect 56545 3755 56555 3775
rect 56575 3755 56585 3775
rect 56545 3725 56585 3755
rect 56545 3705 56555 3725
rect 56575 3705 56585 3725
rect 56545 3690 56585 3705
rect 56605 4025 56645 4040
rect 56605 4005 56615 4025
rect 56635 4005 56645 4025
rect 56605 3975 56645 4005
rect 56605 3955 56615 3975
rect 56635 3955 56645 3975
rect 56605 3925 56645 3955
rect 56605 3905 56615 3925
rect 56635 3905 56645 3925
rect 56605 3875 56645 3905
rect 56605 3855 56615 3875
rect 56635 3855 56645 3875
rect 56605 3825 56645 3855
rect 56605 3805 56615 3825
rect 56635 3805 56645 3825
rect 56605 3775 56645 3805
rect 56605 3755 56615 3775
rect 56635 3755 56645 3775
rect 56605 3725 56645 3755
rect 56605 3705 56615 3725
rect 56635 3705 56645 3725
rect 56605 3690 56645 3705
rect 56665 4025 56705 4040
rect 56665 4005 56675 4025
rect 56695 4005 56705 4025
rect 56665 3975 56705 4005
rect 56665 3955 56675 3975
rect 56695 3955 56705 3975
rect 56665 3925 56705 3955
rect 56665 3905 56675 3925
rect 56695 3905 56705 3925
rect 56665 3875 56705 3905
rect 56665 3855 56675 3875
rect 56695 3855 56705 3875
rect 56665 3825 56705 3855
rect 56665 3805 56675 3825
rect 56695 3805 56705 3825
rect 56665 3775 56705 3805
rect 56665 3755 56675 3775
rect 56695 3755 56705 3775
rect 56665 3725 56705 3755
rect 56665 3705 56675 3725
rect 56695 3705 56705 3725
rect 56665 3690 56705 3705
rect 56725 4025 56765 4040
rect 56725 4005 56735 4025
rect 56755 4005 56765 4025
rect 56725 3975 56765 4005
rect 56725 3955 56735 3975
rect 56755 3955 56765 3975
rect 56725 3925 56765 3955
rect 56725 3905 56735 3925
rect 56755 3905 56765 3925
rect 56725 3875 56765 3905
rect 56725 3855 56735 3875
rect 56755 3855 56765 3875
rect 56725 3825 56765 3855
rect 56725 3805 56735 3825
rect 56755 3805 56765 3825
rect 56725 3775 56765 3805
rect 56725 3755 56735 3775
rect 56755 3755 56765 3775
rect 56725 3725 56765 3755
rect 56725 3705 56735 3725
rect 56755 3705 56765 3725
rect 56725 3690 56765 3705
rect 57035 4025 57075 4040
rect 57035 4005 57045 4025
rect 57065 4005 57075 4025
rect 57035 3975 57075 4005
rect 57035 3955 57045 3975
rect 57065 3955 57075 3975
rect 57035 3925 57075 3955
rect 57035 3905 57045 3925
rect 57065 3905 57075 3925
rect 57035 3875 57075 3905
rect 57035 3855 57045 3875
rect 57065 3855 57075 3875
rect 57035 3825 57075 3855
rect 57035 3805 57045 3825
rect 57065 3805 57075 3825
rect 57035 3775 57075 3805
rect 57035 3755 57045 3775
rect 57065 3755 57075 3775
rect 57035 3725 57075 3755
rect 57035 3705 57045 3725
rect 57065 3705 57075 3725
rect 57035 3690 57075 3705
rect 57095 4025 57135 4040
rect 57095 4005 57105 4025
rect 57125 4005 57135 4025
rect 57095 3975 57135 4005
rect 57095 3955 57105 3975
rect 57125 3955 57135 3975
rect 57095 3925 57135 3955
rect 57095 3905 57105 3925
rect 57125 3905 57135 3925
rect 57095 3875 57135 3905
rect 57095 3855 57105 3875
rect 57125 3855 57135 3875
rect 57095 3825 57135 3855
rect 57095 3805 57105 3825
rect 57125 3805 57135 3825
rect 57095 3775 57135 3805
rect 57095 3755 57105 3775
rect 57125 3755 57135 3775
rect 57095 3725 57135 3755
rect 57095 3705 57105 3725
rect 57125 3705 57135 3725
rect 57095 3690 57135 3705
rect 57155 4025 57195 4040
rect 57155 4005 57165 4025
rect 57185 4005 57195 4025
rect 57155 3975 57195 4005
rect 57155 3955 57165 3975
rect 57185 3955 57195 3975
rect 57155 3925 57195 3955
rect 57155 3905 57165 3925
rect 57185 3905 57195 3925
rect 57155 3875 57195 3905
rect 57155 3855 57165 3875
rect 57185 3855 57195 3875
rect 57155 3825 57195 3855
rect 57155 3805 57165 3825
rect 57185 3805 57195 3825
rect 57155 3775 57195 3805
rect 57155 3755 57165 3775
rect 57185 3755 57195 3775
rect 57155 3725 57195 3755
rect 57155 3705 57165 3725
rect 57185 3705 57195 3725
rect 57155 3690 57195 3705
rect 57215 4025 57255 4040
rect 57215 4005 57225 4025
rect 57245 4005 57255 4025
rect 57215 3975 57255 4005
rect 57215 3955 57225 3975
rect 57245 3955 57255 3975
rect 57215 3925 57255 3955
rect 57215 3905 57225 3925
rect 57245 3905 57255 3925
rect 57215 3875 57255 3905
rect 57215 3855 57225 3875
rect 57245 3855 57255 3875
rect 57215 3825 57255 3855
rect 57215 3805 57225 3825
rect 57245 3805 57255 3825
rect 57215 3775 57255 3805
rect 57215 3755 57225 3775
rect 57245 3755 57255 3775
rect 57215 3725 57255 3755
rect 57215 3705 57225 3725
rect 57245 3705 57255 3725
rect 57215 3690 57255 3705
rect 57275 4025 57315 4040
rect 57275 4005 57285 4025
rect 57305 4005 57315 4025
rect 57275 3975 57315 4005
rect 57275 3955 57285 3975
rect 57305 3955 57315 3975
rect 57275 3925 57315 3955
rect 57275 3905 57285 3925
rect 57305 3905 57315 3925
rect 57275 3875 57315 3905
rect 57275 3855 57285 3875
rect 57305 3855 57315 3875
rect 57275 3825 57315 3855
rect 57275 3805 57285 3825
rect 57305 3805 57315 3825
rect 57275 3775 57315 3805
rect 57275 3755 57285 3775
rect 57305 3755 57315 3775
rect 57275 3725 57315 3755
rect 57275 3705 57285 3725
rect 57305 3705 57315 3725
rect 57275 3690 57315 3705
rect 57335 4025 57375 4040
rect 57335 4005 57345 4025
rect 57365 4005 57375 4025
rect 57335 3975 57375 4005
rect 57335 3955 57345 3975
rect 57365 3955 57375 3975
rect 57335 3925 57375 3955
rect 57335 3905 57345 3925
rect 57365 3905 57375 3925
rect 57335 3875 57375 3905
rect 57335 3855 57345 3875
rect 57365 3855 57375 3875
rect 57335 3825 57375 3855
rect 57335 3805 57345 3825
rect 57365 3805 57375 3825
rect 57335 3775 57375 3805
rect 57335 3755 57345 3775
rect 57365 3755 57375 3775
rect 57335 3725 57375 3755
rect 57335 3705 57345 3725
rect 57365 3705 57375 3725
rect 57335 3690 57375 3705
rect 57395 4025 57435 4040
rect 57395 4005 57405 4025
rect 57425 4005 57435 4025
rect 57395 3975 57435 4005
rect 57395 3955 57405 3975
rect 57425 3955 57435 3975
rect 57395 3925 57435 3955
rect 57395 3905 57405 3925
rect 57425 3905 57435 3925
rect 57395 3875 57435 3905
rect 57395 3855 57405 3875
rect 57425 3855 57435 3875
rect 57395 3825 57435 3855
rect 57395 3805 57405 3825
rect 57425 3805 57435 3825
rect 57395 3775 57435 3805
rect 57395 3755 57405 3775
rect 57425 3755 57435 3775
rect 57395 3725 57435 3755
rect 57395 3705 57405 3725
rect 57425 3705 57435 3725
rect 57395 3690 57435 3705
rect 57455 4025 57495 4040
rect 57455 4005 57465 4025
rect 57485 4005 57495 4025
rect 57455 3975 57495 4005
rect 57455 3955 57465 3975
rect 57485 3955 57495 3975
rect 57455 3925 57495 3955
rect 57455 3905 57465 3925
rect 57485 3905 57495 3925
rect 57455 3875 57495 3905
rect 57455 3855 57465 3875
rect 57485 3855 57495 3875
rect 57455 3825 57495 3855
rect 57455 3805 57465 3825
rect 57485 3805 57495 3825
rect 57455 3775 57495 3805
rect 57455 3755 57465 3775
rect 57485 3755 57495 3775
rect 57455 3725 57495 3755
rect 57455 3705 57465 3725
rect 57485 3705 57495 3725
rect 57455 3690 57495 3705
rect 57515 4025 57555 4040
rect 57515 4005 57525 4025
rect 57545 4005 57555 4025
rect 57515 3975 57555 4005
rect 57515 3955 57525 3975
rect 57545 3955 57555 3975
rect 57515 3925 57555 3955
rect 57515 3905 57525 3925
rect 57545 3905 57555 3925
rect 57515 3875 57555 3905
rect 57515 3855 57525 3875
rect 57545 3855 57555 3875
rect 57515 3825 57555 3855
rect 57515 3805 57525 3825
rect 57545 3805 57555 3825
rect 57515 3775 57555 3805
rect 57515 3755 57525 3775
rect 57545 3755 57555 3775
rect 57515 3725 57555 3755
rect 57515 3705 57525 3725
rect 57545 3705 57555 3725
rect 57515 3690 57555 3705
rect 57575 4025 57615 4040
rect 57575 4005 57585 4025
rect 57605 4005 57615 4025
rect 57575 3975 57615 4005
rect 57575 3955 57585 3975
rect 57605 3955 57615 3975
rect 57575 3925 57615 3955
rect 57575 3905 57585 3925
rect 57605 3905 57615 3925
rect 57575 3875 57615 3905
rect 57575 3855 57585 3875
rect 57605 3855 57615 3875
rect 57575 3825 57615 3855
rect 57575 3805 57585 3825
rect 57605 3805 57615 3825
rect 57575 3775 57615 3805
rect 57575 3755 57585 3775
rect 57605 3755 57615 3775
rect 57575 3725 57615 3755
rect 57575 3705 57585 3725
rect 57605 3705 57615 3725
rect 57575 3690 57615 3705
rect 57635 4025 57675 4040
rect 57635 4005 57645 4025
rect 57665 4005 57675 4025
rect 57635 3975 57675 4005
rect 57635 3955 57645 3975
rect 57665 3955 57675 3975
rect 57635 3925 57675 3955
rect 57635 3905 57645 3925
rect 57665 3905 57675 3925
rect 57635 3875 57675 3905
rect 57635 3855 57645 3875
rect 57665 3855 57675 3875
rect 57635 3825 57675 3855
rect 57635 3805 57645 3825
rect 57665 3805 57675 3825
rect 57635 3775 57675 3805
rect 57635 3755 57645 3775
rect 57665 3755 57675 3775
rect 57635 3725 57675 3755
rect 57635 3705 57645 3725
rect 57665 3705 57675 3725
rect 57635 3690 57675 3705
rect 57695 4025 57735 4040
rect 57695 4005 57705 4025
rect 57725 4005 57735 4025
rect 57695 3975 57735 4005
rect 57695 3955 57705 3975
rect 57725 3955 57735 3975
rect 57695 3925 57735 3955
rect 57695 3905 57705 3925
rect 57725 3905 57735 3925
rect 57695 3875 57735 3905
rect 57695 3855 57705 3875
rect 57725 3855 57735 3875
rect 57695 3825 57735 3855
rect 57695 3805 57705 3825
rect 57725 3805 57735 3825
rect 57695 3775 57735 3805
rect 57695 3755 57705 3775
rect 57725 3755 57735 3775
rect 57695 3725 57735 3755
rect 57695 3705 57705 3725
rect 57725 3705 57735 3725
rect 57695 3690 57735 3705
rect 57755 4025 57795 4040
rect 57755 4005 57765 4025
rect 57785 4005 57795 4025
rect 57755 3975 57795 4005
rect 57755 3955 57765 3975
rect 57785 3955 57795 3975
rect 57755 3925 57795 3955
rect 57755 3905 57765 3925
rect 57785 3905 57795 3925
rect 57755 3875 57795 3905
rect 57755 3855 57765 3875
rect 57785 3855 57795 3875
rect 57755 3825 57795 3855
rect 57755 3805 57765 3825
rect 57785 3805 57795 3825
rect 57755 3775 57795 3805
rect 57755 3755 57765 3775
rect 57785 3755 57795 3775
rect 57755 3725 57795 3755
rect 57755 3705 57765 3725
rect 57785 3705 57795 3725
rect 57755 3690 57795 3705
rect 58085 4025 58125 4040
rect 58085 4005 58095 4025
rect 58115 4005 58125 4025
rect 58085 3975 58125 4005
rect 58085 3955 58095 3975
rect 58115 3955 58125 3975
rect 58085 3925 58125 3955
rect 58085 3905 58095 3925
rect 58115 3905 58125 3925
rect 58085 3875 58125 3905
rect 58085 3855 58095 3875
rect 58115 3855 58125 3875
rect 58085 3825 58125 3855
rect 58085 3805 58095 3825
rect 58115 3805 58125 3825
rect 58085 3775 58125 3805
rect 58085 3755 58095 3775
rect 58115 3755 58125 3775
rect 58085 3725 58125 3755
rect 58085 3705 58095 3725
rect 58115 3705 58125 3725
rect 58085 3690 58125 3705
rect 58145 4025 58185 4040
rect 58145 4005 58155 4025
rect 58175 4005 58185 4025
rect 58145 3975 58185 4005
rect 58145 3955 58155 3975
rect 58175 3955 58185 3975
rect 58145 3925 58185 3955
rect 58145 3905 58155 3925
rect 58175 3905 58185 3925
rect 58145 3875 58185 3905
rect 58145 3855 58155 3875
rect 58175 3855 58185 3875
rect 58145 3825 58185 3855
rect 58145 3805 58155 3825
rect 58175 3805 58185 3825
rect 58145 3775 58185 3805
rect 58145 3755 58155 3775
rect 58175 3755 58185 3775
rect 58145 3725 58185 3755
rect 58145 3705 58155 3725
rect 58175 3705 58185 3725
rect 58145 3690 58185 3705
rect 58205 4025 58245 4040
rect 58205 4005 58215 4025
rect 58235 4005 58245 4025
rect 58205 3975 58245 4005
rect 58205 3955 58215 3975
rect 58235 3955 58245 3975
rect 58205 3925 58245 3955
rect 58205 3905 58215 3925
rect 58235 3905 58245 3925
rect 58205 3875 58245 3905
rect 58205 3855 58215 3875
rect 58235 3855 58245 3875
rect 58205 3825 58245 3855
rect 58205 3805 58215 3825
rect 58235 3805 58245 3825
rect 58205 3775 58245 3805
rect 58205 3755 58215 3775
rect 58235 3755 58245 3775
rect 58205 3725 58245 3755
rect 58205 3705 58215 3725
rect 58235 3705 58245 3725
rect 58205 3690 58245 3705
rect 58265 4025 58305 4040
rect 58265 4005 58275 4025
rect 58295 4005 58305 4025
rect 58265 3975 58305 4005
rect 58265 3955 58275 3975
rect 58295 3955 58305 3975
rect 58265 3925 58305 3955
rect 58265 3905 58275 3925
rect 58295 3905 58305 3925
rect 58265 3875 58305 3905
rect 58265 3855 58275 3875
rect 58295 3855 58305 3875
rect 58265 3825 58305 3855
rect 58265 3805 58275 3825
rect 58295 3805 58305 3825
rect 58265 3775 58305 3805
rect 58265 3755 58275 3775
rect 58295 3755 58305 3775
rect 58265 3725 58305 3755
rect 58265 3705 58275 3725
rect 58295 3705 58305 3725
rect 58265 3690 58305 3705
rect 58325 4025 58365 4040
rect 58325 4005 58335 4025
rect 58355 4005 58365 4025
rect 58325 3975 58365 4005
rect 58325 3955 58335 3975
rect 58355 3955 58365 3975
rect 58325 3925 58365 3955
rect 58325 3905 58335 3925
rect 58355 3905 58365 3925
rect 58325 3875 58365 3905
rect 58325 3855 58335 3875
rect 58355 3855 58365 3875
rect 58325 3825 58365 3855
rect 58325 3805 58335 3825
rect 58355 3805 58365 3825
rect 58325 3775 58365 3805
rect 58325 3755 58335 3775
rect 58355 3755 58365 3775
rect 58325 3725 58365 3755
rect 58325 3705 58335 3725
rect 58355 3705 58365 3725
rect 58325 3690 58365 3705
rect 58385 4025 58425 4040
rect 58385 4005 58395 4025
rect 58415 4005 58425 4025
rect 58385 3975 58425 4005
rect 58385 3955 58395 3975
rect 58415 3955 58425 3975
rect 58385 3925 58425 3955
rect 58385 3905 58395 3925
rect 58415 3905 58425 3925
rect 58385 3875 58425 3905
rect 58385 3855 58395 3875
rect 58415 3855 58425 3875
rect 58385 3825 58425 3855
rect 58385 3805 58395 3825
rect 58415 3805 58425 3825
rect 58385 3775 58425 3805
rect 58385 3755 58395 3775
rect 58415 3755 58425 3775
rect 58385 3725 58425 3755
rect 58385 3705 58395 3725
rect 58415 3705 58425 3725
rect 58385 3690 58425 3705
rect 58445 4025 58485 4040
rect 58445 4005 58455 4025
rect 58475 4005 58485 4025
rect 58445 3975 58485 4005
rect 58445 3955 58455 3975
rect 58475 3955 58485 3975
rect 58445 3925 58485 3955
rect 58445 3905 58455 3925
rect 58475 3905 58485 3925
rect 58445 3875 58485 3905
rect 58445 3855 58455 3875
rect 58475 3855 58485 3875
rect 58445 3825 58485 3855
rect 58445 3805 58455 3825
rect 58475 3805 58485 3825
rect 58445 3775 58485 3805
rect 58445 3755 58455 3775
rect 58475 3755 58485 3775
rect 58445 3725 58485 3755
rect 58445 3705 58455 3725
rect 58475 3705 58485 3725
rect 58445 3690 58485 3705
rect 58505 4025 58545 4040
rect 58505 4005 58515 4025
rect 58535 4005 58545 4025
rect 58505 3975 58545 4005
rect 58505 3955 58515 3975
rect 58535 3955 58545 3975
rect 58505 3925 58545 3955
rect 58505 3905 58515 3925
rect 58535 3905 58545 3925
rect 58505 3875 58545 3905
rect 58505 3855 58515 3875
rect 58535 3855 58545 3875
rect 58505 3825 58545 3855
rect 58505 3805 58515 3825
rect 58535 3805 58545 3825
rect 58505 3775 58545 3805
rect 58505 3755 58515 3775
rect 58535 3755 58545 3775
rect 58505 3725 58545 3755
rect 58505 3705 58515 3725
rect 58535 3705 58545 3725
rect 58505 3690 58545 3705
rect 58565 4025 58605 4040
rect 58565 4005 58575 4025
rect 58595 4005 58605 4025
rect 58565 3975 58605 4005
rect 58565 3955 58575 3975
rect 58595 3955 58605 3975
rect 58565 3925 58605 3955
rect 58565 3905 58575 3925
rect 58595 3905 58605 3925
rect 58565 3875 58605 3905
rect 58565 3855 58575 3875
rect 58595 3855 58605 3875
rect 58565 3825 58605 3855
rect 58565 3805 58575 3825
rect 58595 3805 58605 3825
rect 58565 3775 58605 3805
rect 58565 3755 58575 3775
rect 58595 3755 58605 3775
rect 58565 3725 58605 3755
rect 58565 3705 58575 3725
rect 58595 3705 58605 3725
rect 58565 3690 58605 3705
rect 58625 4025 58665 4040
rect 58625 4005 58635 4025
rect 58655 4005 58665 4025
rect 58625 3975 58665 4005
rect 58625 3955 58635 3975
rect 58655 3955 58665 3975
rect 58625 3925 58665 3955
rect 58625 3905 58635 3925
rect 58655 3905 58665 3925
rect 58625 3875 58665 3905
rect 58625 3855 58635 3875
rect 58655 3855 58665 3875
rect 58625 3825 58665 3855
rect 58625 3805 58635 3825
rect 58655 3805 58665 3825
rect 58625 3775 58665 3805
rect 58625 3755 58635 3775
rect 58655 3755 58665 3775
rect 58625 3725 58665 3755
rect 58625 3705 58635 3725
rect 58655 3705 58665 3725
rect 58625 3690 58665 3705
rect 58685 4025 58725 4040
rect 58685 4005 58695 4025
rect 58715 4005 58725 4025
rect 58685 3975 58725 4005
rect 58685 3955 58695 3975
rect 58715 3955 58725 3975
rect 58685 3925 58725 3955
rect 58685 3905 58695 3925
rect 58715 3905 58725 3925
rect 58685 3875 58725 3905
rect 58685 3855 58695 3875
rect 58715 3855 58725 3875
rect 58685 3825 58725 3855
rect 58685 3805 58695 3825
rect 58715 3805 58725 3825
rect 58685 3775 58725 3805
rect 58685 3755 58695 3775
rect 58715 3755 58725 3775
rect 58685 3725 58725 3755
rect 58685 3705 58695 3725
rect 58715 3705 58725 3725
rect 58685 3690 58725 3705
rect 58745 4025 58785 4040
rect 58745 4005 58755 4025
rect 58775 4005 58785 4025
rect 58745 3975 58785 4005
rect 58745 3955 58755 3975
rect 58775 3955 58785 3975
rect 58745 3925 58785 3955
rect 58745 3905 58755 3925
rect 58775 3905 58785 3925
rect 58745 3875 58785 3905
rect 58745 3855 58755 3875
rect 58775 3855 58785 3875
rect 58745 3825 58785 3855
rect 58745 3805 58755 3825
rect 58775 3805 58785 3825
rect 58745 3775 58785 3805
rect 58745 3755 58755 3775
rect 58775 3755 58785 3775
rect 58745 3725 58785 3755
rect 58745 3705 58755 3725
rect 58775 3705 58785 3725
rect 58745 3690 58785 3705
rect 58805 4025 58845 4040
rect 58805 4005 58815 4025
rect 58835 4005 58845 4025
rect 58805 3975 58845 4005
rect 58805 3955 58815 3975
rect 58835 3955 58845 3975
rect 58805 3925 58845 3955
rect 58805 3905 58815 3925
rect 58835 3905 58845 3925
rect 58805 3875 58845 3905
rect 58805 3855 58815 3875
rect 58835 3855 58845 3875
rect 58805 3825 58845 3855
rect 58805 3805 58815 3825
rect 58835 3805 58845 3825
rect 58805 3775 58845 3805
rect 58805 3755 58815 3775
rect 58835 3755 58845 3775
rect 58805 3725 58845 3755
rect 58805 3705 58815 3725
rect 58835 3705 58845 3725
rect 58805 3690 58845 3705
rect 54955 3315 54995 3330
rect 54955 3295 54965 3315
rect 54985 3295 54995 3315
rect 54955 3265 54995 3295
rect 54955 3245 54965 3265
rect 54985 3245 54995 3265
rect 54955 3215 54995 3245
rect 54955 3195 54965 3215
rect 54985 3195 54995 3215
rect 54955 3165 54995 3195
rect 54955 3145 54965 3165
rect 54985 3145 54995 3165
rect 54955 3115 54995 3145
rect 54955 3095 54965 3115
rect 54985 3095 54995 3115
rect 54955 3065 54995 3095
rect 54955 3045 54965 3065
rect 54985 3045 54995 3065
rect 54955 3015 54995 3045
rect 54955 2995 54965 3015
rect 54985 2995 54995 3015
rect 54955 2965 54995 2995
rect 54955 2945 54965 2965
rect 54985 2945 54995 2965
rect 54955 2915 54995 2945
rect 54955 2895 54965 2915
rect 54985 2895 54995 2915
rect 54955 2865 54995 2895
rect 54955 2845 54965 2865
rect 54985 2845 54995 2865
rect 54955 2815 54995 2845
rect 54955 2795 54965 2815
rect 54985 2795 54995 2815
rect 54955 2765 54995 2795
rect 54955 2745 54965 2765
rect 54985 2745 54995 2765
rect 54955 2730 54995 2745
rect 55010 3315 55050 3330
rect 55010 3295 55020 3315
rect 55040 3295 55050 3315
rect 55010 3265 55050 3295
rect 55010 3245 55020 3265
rect 55040 3245 55050 3265
rect 55010 3215 55050 3245
rect 55010 3195 55020 3215
rect 55040 3195 55050 3215
rect 55010 3165 55050 3195
rect 55010 3145 55020 3165
rect 55040 3145 55050 3165
rect 55010 3115 55050 3145
rect 55010 3095 55020 3115
rect 55040 3095 55050 3115
rect 55010 3065 55050 3095
rect 55010 3045 55020 3065
rect 55040 3045 55050 3065
rect 55010 3015 55050 3045
rect 55010 2995 55020 3015
rect 55040 2995 55050 3015
rect 55010 2965 55050 2995
rect 55010 2945 55020 2965
rect 55040 2945 55050 2965
rect 55010 2915 55050 2945
rect 55010 2895 55020 2915
rect 55040 2895 55050 2915
rect 55010 2865 55050 2895
rect 55010 2845 55020 2865
rect 55040 2845 55050 2865
rect 55010 2815 55050 2845
rect 55010 2795 55020 2815
rect 55040 2795 55050 2815
rect 55010 2765 55050 2795
rect 55010 2745 55020 2765
rect 55040 2745 55050 2765
rect 55010 2730 55050 2745
rect 55065 3315 55105 3330
rect 55065 3295 55075 3315
rect 55095 3295 55105 3315
rect 55065 3265 55105 3295
rect 55065 3245 55075 3265
rect 55095 3245 55105 3265
rect 55065 3215 55105 3245
rect 55065 3195 55075 3215
rect 55095 3195 55105 3215
rect 55065 3165 55105 3195
rect 55065 3145 55075 3165
rect 55095 3145 55105 3165
rect 55065 3115 55105 3145
rect 55065 3095 55075 3115
rect 55095 3095 55105 3115
rect 55065 3065 55105 3095
rect 55065 3045 55075 3065
rect 55095 3045 55105 3065
rect 55065 3015 55105 3045
rect 55065 2995 55075 3015
rect 55095 2995 55105 3015
rect 55065 2965 55105 2995
rect 55065 2945 55075 2965
rect 55095 2945 55105 2965
rect 55065 2915 55105 2945
rect 55065 2895 55075 2915
rect 55095 2895 55105 2915
rect 55065 2865 55105 2895
rect 55065 2845 55075 2865
rect 55095 2845 55105 2865
rect 55065 2815 55105 2845
rect 55065 2795 55075 2815
rect 55095 2795 55105 2815
rect 55065 2765 55105 2795
rect 55065 2745 55075 2765
rect 55095 2745 55105 2765
rect 55065 2730 55105 2745
rect 55120 3315 55160 3330
rect 55120 3295 55130 3315
rect 55150 3295 55160 3315
rect 55120 3265 55160 3295
rect 55120 3245 55130 3265
rect 55150 3245 55160 3265
rect 55120 3215 55160 3245
rect 55120 3195 55130 3215
rect 55150 3195 55160 3215
rect 55120 3165 55160 3195
rect 55120 3145 55130 3165
rect 55150 3145 55160 3165
rect 55120 3115 55160 3145
rect 55120 3095 55130 3115
rect 55150 3095 55160 3115
rect 55120 3065 55160 3095
rect 55120 3045 55130 3065
rect 55150 3045 55160 3065
rect 55120 3015 55160 3045
rect 55120 2995 55130 3015
rect 55150 2995 55160 3015
rect 55120 2965 55160 2995
rect 55120 2945 55130 2965
rect 55150 2945 55160 2965
rect 55120 2915 55160 2945
rect 55120 2895 55130 2915
rect 55150 2895 55160 2915
rect 55120 2865 55160 2895
rect 55120 2845 55130 2865
rect 55150 2845 55160 2865
rect 55120 2815 55160 2845
rect 55120 2795 55130 2815
rect 55150 2795 55160 2815
rect 55120 2765 55160 2795
rect 55120 2745 55130 2765
rect 55150 2745 55160 2765
rect 55120 2730 55160 2745
rect 55175 3315 55215 3330
rect 55175 3295 55185 3315
rect 55205 3295 55215 3315
rect 55175 3265 55215 3295
rect 55175 3245 55185 3265
rect 55205 3245 55215 3265
rect 55175 3215 55215 3245
rect 55175 3195 55185 3215
rect 55205 3195 55215 3215
rect 55175 3165 55215 3195
rect 55175 3145 55185 3165
rect 55205 3145 55215 3165
rect 55175 3115 55215 3145
rect 55175 3095 55185 3115
rect 55205 3095 55215 3115
rect 55175 3065 55215 3095
rect 55175 3045 55185 3065
rect 55205 3045 55215 3065
rect 55175 3015 55215 3045
rect 55175 2995 55185 3015
rect 55205 2995 55215 3015
rect 55175 2965 55215 2995
rect 55175 2945 55185 2965
rect 55205 2945 55215 2965
rect 55175 2915 55215 2945
rect 55175 2895 55185 2915
rect 55205 2895 55215 2915
rect 55175 2865 55215 2895
rect 55175 2845 55185 2865
rect 55205 2845 55215 2865
rect 55175 2815 55215 2845
rect 55175 2795 55185 2815
rect 55205 2795 55215 2815
rect 55175 2765 55215 2795
rect 55175 2745 55185 2765
rect 55205 2745 55215 2765
rect 55175 2730 55215 2745
rect 55230 3315 55270 3330
rect 55230 3295 55240 3315
rect 55260 3295 55270 3315
rect 55230 3265 55270 3295
rect 55230 3245 55240 3265
rect 55260 3245 55270 3265
rect 55230 3215 55270 3245
rect 55230 3195 55240 3215
rect 55260 3195 55270 3215
rect 55230 3165 55270 3195
rect 55230 3145 55240 3165
rect 55260 3145 55270 3165
rect 55230 3115 55270 3145
rect 55230 3095 55240 3115
rect 55260 3095 55270 3115
rect 55230 3065 55270 3095
rect 55230 3045 55240 3065
rect 55260 3045 55270 3065
rect 55230 3015 55270 3045
rect 55230 2995 55240 3015
rect 55260 2995 55270 3015
rect 55230 2965 55270 2995
rect 55230 2945 55240 2965
rect 55260 2945 55270 2965
rect 55230 2915 55270 2945
rect 55230 2895 55240 2915
rect 55260 2895 55270 2915
rect 55230 2865 55270 2895
rect 55230 2845 55240 2865
rect 55260 2845 55270 2865
rect 55230 2815 55270 2845
rect 55230 2795 55240 2815
rect 55260 2795 55270 2815
rect 55230 2765 55270 2795
rect 55230 2745 55240 2765
rect 55260 2745 55270 2765
rect 55230 2730 55270 2745
rect 55285 3315 55325 3330
rect 55285 3295 55295 3315
rect 55315 3295 55325 3315
rect 55285 3265 55325 3295
rect 55285 3245 55295 3265
rect 55315 3245 55325 3265
rect 55285 3215 55325 3245
rect 55285 3195 55295 3215
rect 55315 3195 55325 3215
rect 55285 3165 55325 3195
rect 55285 3145 55295 3165
rect 55315 3145 55325 3165
rect 55285 3115 55325 3145
rect 55285 3095 55295 3115
rect 55315 3095 55325 3115
rect 55285 3065 55325 3095
rect 55285 3045 55295 3065
rect 55315 3045 55325 3065
rect 55285 3015 55325 3045
rect 55285 2995 55295 3015
rect 55315 2995 55325 3015
rect 55285 2965 55325 2995
rect 55285 2945 55295 2965
rect 55315 2945 55325 2965
rect 55285 2915 55325 2945
rect 55285 2895 55295 2915
rect 55315 2895 55325 2915
rect 55285 2865 55325 2895
rect 55285 2845 55295 2865
rect 55315 2845 55325 2865
rect 55285 2815 55325 2845
rect 55285 2795 55295 2815
rect 55315 2795 55325 2815
rect 55285 2765 55325 2795
rect 55285 2745 55295 2765
rect 55315 2745 55325 2765
rect 55285 2730 55325 2745
rect 55340 3315 55380 3330
rect 55340 3295 55350 3315
rect 55370 3295 55380 3315
rect 55340 3265 55380 3295
rect 55340 3245 55350 3265
rect 55370 3245 55380 3265
rect 55340 3215 55380 3245
rect 55340 3195 55350 3215
rect 55370 3195 55380 3215
rect 55340 3165 55380 3195
rect 55340 3145 55350 3165
rect 55370 3145 55380 3165
rect 55340 3115 55380 3145
rect 55340 3095 55350 3115
rect 55370 3095 55380 3115
rect 55340 3065 55380 3095
rect 55340 3045 55350 3065
rect 55370 3045 55380 3065
rect 55340 3015 55380 3045
rect 55340 2995 55350 3015
rect 55370 2995 55380 3015
rect 55340 2965 55380 2995
rect 55340 2945 55350 2965
rect 55370 2945 55380 2965
rect 55340 2915 55380 2945
rect 55340 2895 55350 2915
rect 55370 2895 55380 2915
rect 55340 2865 55380 2895
rect 55340 2845 55350 2865
rect 55370 2845 55380 2865
rect 55340 2815 55380 2845
rect 55340 2795 55350 2815
rect 55370 2795 55380 2815
rect 55340 2765 55380 2795
rect 55340 2745 55350 2765
rect 55370 2745 55380 2765
rect 55340 2730 55380 2745
rect 55395 3315 55435 3330
rect 55395 3295 55405 3315
rect 55425 3295 55435 3315
rect 55395 3265 55435 3295
rect 55395 3245 55405 3265
rect 55425 3245 55435 3265
rect 55395 3215 55435 3245
rect 55395 3195 55405 3215
rect 55425 3195 55435 3215
rect 55395 3165 55435 3195
rect 55395 3145 55405 3165
rect 55425 3145 55435 3165
rect 55395 3115 55435 3145
rect 55395 3095 55405 3115
rect 55425 3095 55435 3115
rect 55395 3065 55435 3095
rect 55395 3045 55405 3065
rect 55425 3045 55435 3065
rect 55395 3015 55435 3045
rect 55395 2995 55405 3015
rect 55425 2995 55435 3015
rect 55395 2965 55435 2995
rect 55395 2945 55405 2965
rect 55425 2945 55435 2965
rect 55395 2915 55435 2945
rect 55395 2895 55405 2915
rect 55425 2895 55435 2915
rect 55395 2865 55435 2895
rect 55395 2845 55405 2865
rect 55425 2845 55435 2865
rect 55395 2815 55435 2845
rect 55395 2795 55405 2815
rect 55425 2795 55435 2815
rect 55395 2765 55435 2795
rect 55395 2745 55405 2765
rect 55425 2745 55435 2765
rect 55395 2730 55435 2745
rect 55450 3315 55490 3330
rect 55450 3295 55460 3315
rect 55480 3295 55490 3315
rect 55450 3265 55490 3295
rect 55450 3245 55460 3265
rect 55480 3245 55490 3265
rect 55450 3215 55490 3245
rect 55450 3195 55460 3215
rect 55480 3195 55490 3215
rect 55450 3165 55490 3195
rect 55450 3145 55460 3165
rect 55480 3145 55490 3165
rect 55450 3115 55490 3145
rect 55450 3095 55460 3115
rect 55480 3095 55490 3115
rect 55450 3065 55490 3095
rect 55450 3045 55460 3065
rect 55480 3045 55490 3065
rect 55450 3015 55490 3045
rect 55450 2995 55460 3015
rect 55480 2995 55490 3015
rect 55450 2965 55490 2995
rect 55450 2945 55460 2965
rect 55480 2945 55490 2965
rect 55450 2915 55490 2945
rect 55450 2895 55460 2915
rect 55480 2895 55490 2915
rect 55450 2865 55490 2895
rect 55450 2845 55460 2865
rect 55480 2845 55490 2865
rect 55450 2815 55490 2845
rect 55450 2795 55460 2815
rect 55480 2795 55490 2815
rect 55450 2765 55490 2795
rect 55450 2745 55460 2765
rect 55480 2745 55490 2765
rect 55450 2730 55490 2745
rect 55505 3315 55545 3330
rect 55505 3295 55515 3315
rect 55535 3295 55545 3315
rect 55505 3265 55545 3295
rect 55505 3245 55515 3265
rect 55535 3245 55545 3265
rect 55505 3215 55545 3245
rect 55505 3195 55515 3215
rect 55535 3195 55545 3215
rect 55505 3165 55545 3195
rect 55505 3145 55515 3165
rect 55535 3145 55545 3165
rect 55505 3115 55545 3145
rect 55505 3095 55515 3115
rect 55535 3095 55545 3115
rect 55505 3065 55545 3095
rect 55505 3045 55515 3065
rect 55535 3045 55545 3065
rect 55505 3015 55545 3045
rect 55505 2995 55515 3015
rect 55535 2995 55545 3015
rect 55505 2965 55545 2995
rect 55505 2945 55515 2965
rect 55535 2945 55545 2965
rect 55505 2915 55545 2945
rect 55505 2895 55515 2915
rect 55535 2895 55545 2915
rect 55505 2865 55545 2895
rect 55505 2845 55515 2865
rect 55535 2845 55545 2865
rect 55505 2815 55545 2845
rect 55505 2795 55515 2815
rect 55535 2795 55545 2815
rect 55505 2765 55545 2795
rect 55505 2745 55515 2765
rect 55535 2745 55545 2765
rect 55505 2730 55545 2745
rect 55560 3315 55600 3330
rect 55560 3295 55570 3315
rect 55590 3295 55600 3315
rect 55560 3265 55600 3295
rect 55560 3245 55570 3265
rect 55590 3245 55600 3265
rect 55560 3215 55600 3245
rect 55560 3195 55570 3215
rect 55590 3195 55600 3215
rect 55560 3165 55600 3195
rect 55560 3145 55570 3165
rect 55590 3145 55600 3165
rect 55560 3115 55600 3145
rect 55560 3095 55570 3115
rect 55590 3095 55600 3115
rect 55560 3065 55600 3095
rect 55560 3045 55570 3065
rect 55590 3045 55600 3065
rect 55560 3015 55600 3045
rect 55560 2995 55570 3015
rect 55590 2995 55600 3015
rect 55560 2965 55600 2995
rect 55560 2945 55570 2965
rect 55590 2945 55600 2965
rect 55560 2915 55600 2945
rect 55560 2895 55570 2915
rect 55590 2895 55600 2915
rect 55560 2865 55600 2895
rect 55560 2845 55570 2865
rect 55590 2845 55600 2865
rect 55560 2815 55600 2845
rect 55560 2795 55570 2815
rect 55590 2795 55600 2815
rect 55560 2765 55600 2795
rect 55560 2745 55570 2765
rect 55590 2745 55600 2765
rect 55560 2730 55600 2745
rect 55615 3315 55655 3330
rect 55615 3295 55625 3315
rect 55645 3295 55655 3315
rect 55615 3265 55655 3295
rect 55615 3245 55625 3265
rect 55645 3245 55655 3265
rect 55615 3215 55655 3245
rect 55615 3195 55625 3215
rect 55645 3195 55655 3215
rect 55615 3165 55655 3195
rect 55615 3145 55625 3165
rect 55645 3145 55655 3165
rect 55615 3115 55655 3145
rect 55615 3095 55625 3115
rect 55645 3095 55655 3115
rect 55615 3065 55655 3095
rect 55615 3045 55625 3065
rect 55645 3045 55655 3065
rect 55615 3015 55655 3045
rect 55615 2995 55625 3015
rect 55645 2995 55655 3015
rect 55615 2965 55655 2995
rect 55615 2945 55625 2965
rect 55645 2945 55655 2965
rect 55615 2915 55655 2945
rect 55615 2895 55625 2915
rect 55645 2895 55655 2915
rect 55615 2865 55655 2895
rect 55615 2845 55625 2865
rect 55645 2845 55655 2865
rect 55615 2815 55655 2845
rect 55615 2795 55625 2815
rect 55645 2795 55655 2815
rect 55615 2765 55655 2795
rect 55615 2745 55625 2765
rect 55645 2745 55655 2765
rect 55615 2730 55655 2745
rect 56275 3315 56315 3330
rect 56275 3295 56285 3315
rect 56305 3295 56315 3315
rect 56275 3280 56315 3295
rect 56330 3315 56370 3330
rect 56330 3295 56340 3315
rect 56360 3295 56370 3315
rect 56330 3280 56370 3295
rect 56385 3315 56425 3330
rect 56385 3295 56395 3315
rect 56415 3295 56425 3315
rect 56385 3280 56425 3295
rect 56440 3315 56480 3330
rect 56440 3295 56450 3315
rect 56470 3295 56480 3315
rect 56440 3280 56480 3295
rect 56495 3315 56535 3330
rect 56495 3295 56505 3315
rect 56525 3295 56535 3315
rect 56495 3280 56535 3295
rect 56550 3315 56590 3330
rect 56550 3295 56560 3315
rect 56580 3295 56590 3315
rect 56550 3280 56590 3295
rect 56605 3315 56645 3330
rect 56605 3295 56615 3315
rect 56635 3295 56645 3315
rect 56605 3280 56645 3295
rect 56660 3315 56700 3330
rect 56660 3295 56670 3315
rect 56690 3295 56700 3315
rect 56660 3280 56700 3295
rect 56715 3315 56755 3330
rect 56715 3295 56725 3315
rect 56745 3295 56755 3315
rect 56715 3280 56755 3295
rect 56770 3315 56810 3330
rect 56770 3295 56780 3315
rect 56800 3295 56810 3315
rect 56770 3280 56810 3295
rect 56825 3315 56865 3330
rect 56825 3295 56835 3315
rect 56855 3295 56865 3315
rect 56825 3280 56865 3295
rect 56880 3315 56920 3330
rect 56880 3295 56890 3315
rect 56910 3295 56920 3315
rect 56880 3280 56920 3295
rect 56935 3315 56975 3330
rect 56935 3295 56945 3315
rect 56965 3295 56975 3315
rect 56935 3280 56975 3295
rect 56990 3315 57030 3330
rect 56990 3295 57000 3315
rect 57020 3295 57030 3315
rect 56990 3280 57030 3295
rect 57045 3315 57085 3330
rect 57045 3295 57055 3315
rect 57075 3295 57085 3315
rect 57045 3280 57085 3295
rect 57100 3315 57140 3330
rect 57100 3295 57110 3315
rect 57130 3295 57140 3315
rect 57100 3280 57140 3295
rect 57155 3315 57195 3330
rect 57155 3295 57165 3315
rect 57185 3295 57195 3315
rect 57155 3280 57195 3295
rect 57210 3315 57250 3330
rect 57210 3295 57220 3315
rect 57240 3295 57250 3315
rect 57210 3280 57250 3295
rect 57265 3315 57305 3330
rect 57265 3295 57275 3315
rect 57295 3295 57305 3315
rect 57265 3280 57305 3295
rect 57320 3315 57360 3330
rect 57320 3295 57330 3315
rect 57350 3295 57360 3315
rect 57320 3280 57360 3295
rect 57375 3315 57415 3330
rect 57375 3295 57385 3315
rect 57405 3295 57415 3315
rect 57375 3280 57415 3295
rect 57430 3315 57470 3330
rect 57430 3295 57440 3315
rect 57460 3295 57470 3315
rect 57430 3280 57470 3295
rect 57485 3315 57525 3330
rect 57485 3295 57495 3315
rect 57515 3295 57525 3315
rect 57485 3280 57525 3295
rect 56065 2860 56105 2875
rect 56065 2840 56075 2860
rect 56095 2840 56105 2860
rect 56065 2825 56105 2840
rect 56120 2860 56160 2875
rect 56120 2840 56130 2860
rect 56150 2840 56160 2860
rect 56120 2825 56160 2840
rect 56175 2860 56215 2875
rect 56175 2840 56185 2860
rect 56205 2840 56215 2860
rect 56175 2825 56215 2840
rect 56230 2860 56270 2875
rect 56230 2840 56240 2860
rect 56260 2840 56270 2860
rect 56230 2825 56270 2840
rect 56285 2860 56325 2875
rect 56285 2840 56295 2860
rect 56315 2840 56325 2860
rect 56285 2825 56325 2840
rect 56340 2860 56380 2875
rect 56340 2840 56350 2860
rect 56370 2840 56380 2860
rect 56340 2825 56380 2840
rect 56395 2860 56435 2875
rect 56395 2840 56405 2860
rect 56425 2840 56435 2860
rect 56395 2825 56435 2840
rect 56450 2860 56490 2875
rect 56450 2840 56460 2860
rect 56480 2840 56490 2860
rect 56450 2825 56490 2840
rect 56505 2860 56545 2875
rect 56505 2840 56515 2860
rect 56535 2840 56545 2860
rect 56505 2825 56545 2840
rect 56560 2860 56600 2875
rect 56560 2840 56570 2860
rect 56590 2840 56600 2860
rect 56560 2825 56600 2840
rect 56615 2860 56655 2875
rect 56615 2840 56625 2860
rect 56645 2840 56655 2860
rect 56615 2825 56655 2840
rect 56670 2860 56710 2875
rect 56670 2840 56680 2860
rect 56700 2840 56710 2860
rect 56670 2825 56710 2840
rect 56725 2860 56765 2875
rect 56725 2840 56735 2860
rect 56755 2840 56765 2860
rect 56725 2825 56765 2840
rect 57035 2860 57075 2875
rect 57035 2840 57045 2860
rect 57065 2840 57075 2860
rect 57035 2825 57075 2840
rect 57090 2860 57130 2875
rect 57090 2840 57100 2860
rect 57120 2840 57130 2860
rect 57090 2825 57130 2840
rect 57145 2860 57185 2875
rect 57145 2840 57155 2860
rect 57175 2840 57185 2860
rect 57145 2825 57185 2840
rect 57200 2860 57240 2875
rect 57200 2840 57210 2860
rect 57230 2840 57240 2860
rect 57200 2825 57240 2840
rect 57255 2860 57295 2875
rect 57255 2840 57265 2860
rect 57285 2840 57295 2860
rect 57255 2825 57295 2840
rect 57310 2860 57350 2875
rect 57310 2840 57320 2860
rect 57340 2840 57350 2860
rect 57310 2825 57350 2840
rect 57365 2860 57405 2875
rect 57365 2840 57375 2860
rect 57395 2840 57405 2860
rect 57365 2825 57405 2840
rect 57420 2860 57460 2875
rect 57420 2840 57430 2860
rect 57450 2840 57460 2860
rect 57420 2825 57460 2840
rect 57475 2860 57515 2875
rect 57475 2840 57485 2860
rect 57505 2840 57515 2860
rect 57475 2825 57515 2840
rect 57530 2860 57570 2875
rect 57530 2840 57540 2860
rect 57560 2840 57570 2860
rect 57530 2825 57570 2840
rect 57585 2860 57625 2875
rect 57585 2840 57595 2860
rect 57615 2840 57625 2860
rect 57585 2825 57625 2840
rect 57640 2860 57680 2875
rect 57640 2840 57650 2860
rect 57670 2840 57680 2860
rect 57640 2825 57680 2840
rect 57695 2860 57735 2875
rect 57695 2840 57705 2860
rect 57725 2840 57735 2860
rect 57695 2825 57735 2840
rect 58145 3315 58185 3330
rect 58145 3295 58155 3315
rect 58175 3295 58185 3315
rect 58145 3265 58185 3295
rect 58145 3245 58155 3265
rect 58175 3245 58185 3265
rect 58145 3215 58185 3245
rect 58145 3195 58155 3215
rect 58175 3195 58185 3215
rect 58145 3165 58185 3195
rect 58145 3145 58155 3165
rect 58175 3145 58185 3165
rect 58145 3115 58185 3145
rect 58145 3095 58155 3115
rect 58175 3095 58185 3115
rect 58145 3065 58185 3095
rect 58145 3045 58155 3065
rect 58175 3045 58185 3065
rect 58145 3015 58185 3045
rect 58145 2995 58155 3015
rect 58175 2995 58185 3015
rect 58145 2965 58185 2995
rect 58145 2945 58155 2965
rect 58175 2945 58185 2965
rect 58145 2915 58185 2945
rect 58145 2895 58155 2915
rect 58175 2895 58185 2915
rect 58145 2865 58185 2895
rect 58145 2845 58155 2865
rect 58175 2845 58185 2865
rect 58145 2815 58185 2845
rect 58145 2795 58155 2815
rect 58175 2795 58185 2815
rect 58145 2765 58185 2795
rect 58145 2745 58155 2765
rect 58175 2745 58185 2765
rect 58145 2730 58185 2745
rect 58200 3315 58240 3330
rect 58200 3295 58210 3315
rect 58230 3295 58240 3315
rect 58200 3265 58240 3295
rect 58200 3245 58210 3265
rect 58230 3245 58240 3265
rect 58200 3215 58240 3245
rect 58200 3195 58210 3215
rect 58230 3195 58240 3215
rect 58200 3165 58240 3195
rect 58200 3145 58210 3165
rect 58230 3145 58240 3165
rect 58200 3115 58240 3145
rect 58200 3095 58210 3115
rect 58230 3095 58240 3115
rect 58200 3065 58240 3095
rect 58200 3045 58210 3065
rect 58230 3045 58240 3065
rect 58200 3015 58240 3045
rect 58200 2995 58210 3015
rect 58230 2995 58240 3015
rect 58200 2965 58240 2995
rect 58200 2945 58210 2965
rect 58230 2945 58240 2965
rect 58200 2915 58240 2945
rect 58200 2895 58210 2915
rect 58230 2895 58240 2915
rect 58200 2865 58240 2895
rect 58200 2845 58210 2865
rect 58230 2845 58240 2865
rect 58200 2815 58240 2845
rect 58200 2795 58210 2815
rect 58230 2795 58240 2815
rect 58200 2765 58240 2795
rect 58200 2745 58210 2765
rect 58230 2745 58240 2765
rect 58200 2730 58240 2745
rect 58255 3315 58295 3330
rect 58255 3295 58265 3315
rect 58285 3295 58295 3315
rect 58255 3265 58295 3295
rect 58255 3245 58265 3265
rect 58285 3245 58295 3265
rect 58255 3215 58295 3245
rect 58255 3195 58265 3215
rect 58285 3195 58295 3215
rect 58255 3165 58295 3195
rect 58255 3145 58265 3165
rect 58285 3145 58295 3165
rect 58255 3115 58295 3145
rect 58255 3095 58265 3115
rect 58285 3095 58295 3115
rect 58255 3065 58295 3095
rect 58255 3045 58265 3065
rect 58285 3045 58295 3065
rect 58255 3015 58295 3045
rect 58255 2995 58265 3015
rect 58285 2995 58295 3015
rect 58255 2965 58295 2995
rect 58255 2945 58265 2965
rect 58285 2945 58295 2965
rect 58255 2915 58295 2945
rect 58255 2895 58265 2915
rect 58285 2895 58295 2915
rect 58255 2865 58295 2895
rect 58255 2845 58265 2865
rect 58285 2845 58295 2865
rect 58255 2815 58295 2845
rect 58255 2795 58265 2815
rect 58285 2795 58295 2815
rect 58255 2765 58295 2795
rect 58255 2745 58265 2765
rect 58285 2745 58295 2765
rect 58255 2730 58295 2745
rect 58310 3315 58350 3330
rect 58310 3295 58320 3315
rect 58340 3295 58350 3315
rect 58310 3265 58350 3295
rect 58310 3245 58320 3265
rect 58340 3245 58350 3265
rect 58310 3215 58350 3245
rect 58310 3195 58320 3215
rect 58340 3195 58350 3215
rect 58310 3165 58350 3195
rect 58310 3145 58320 3165
rect 58340 3145 58350 3165
rect 58310 3115 58350 3145
rect 58310 3095 58320 3115
rect 58340 3095 58350 3115
rect 58310 3065 58350 3095
rect 58310 3045 58320 3065
rect 58340 3045 58350 3065
rect 58310 3015 58350 3045
rect 58310 2995 58320 3015
rect 58340 2995 58350 3015
rect 58310 2965 58350 2995
rect 58310 2945 58320 2965
rect 58340 2945 58350 2965
rect 58310 2915 58350 2945
rect 58310 2895 58320 2915
rect 58340 2895 58350 2915
rect 58310 2865 58350 2895
rect 58310 2845 58320 2865
rect 58340 2845 58350 2865
rect 58310 2815 58350 2845
rect 58310 2795 58320 2815
rect 58340 2795 58350 2815
rect 58310 2765 58350 2795
rect 58310 2745 58320 2765
rect 58340 2745 58350 2765
rect 58310 2730 58350 2745
rect 58365 3315 58405 3330
rect 58365 3295 58375 3315
rect 58395 3295 58405 3315
rect 58365 3265 58405 3295
rect 58365 3245 58375 3265
rect 58395 3245 58405 3265
rect 58365 3215 58405 3245
rect 58365 3195 58375 3215
rect 58395 3195 58405 3215
rect 58365 3165 58405 3195
rect 58365 3145 58375 3165
rect 58395 3145 58405 3165
rect 58365 3115 58405 3145
rect 58365 3095 58375 3115
rect 58395 3095 58405 3115
rect 58365 3065 58405 3095
rect 58365 3045 58375 3065
rect 58395 3045 58405 3065
rect 58365 3015 58405 3045
rect 58365 2995 58375 3015
rect 58395 2995 58405 3015
rect 58365 2965 58405 2995
rect 58365 2945 58375 2965
rect 58395 2945 58405 2965
rect 58365 2915 58405 2945
rect 58365 2895 58375 2915
rect 58395 2895 58405 2915
rect 58365 2865 58405 2895
rect 58365 2845 58375 2865
rect 58395 2845 58405 2865
rect 58365 2815 58405 2845
rect 58365 2795 58375 2815
rect 58395 2795 58405 2815
rect 58365 2765 58405 2795
rect 58365 2745 58375 2765
rect 58395 2745 58405 2765
rect 58365 2730 58405 2745
rect 58420 3315 58460 3330
rect 58420 3295 58430 3315
rect 58450 3295 58460 3315
rect 58420 3265 58460 3295
rect 58420 3245 58430 3265
rect 58450 3245 58460 3265
rect 58420 3215 58460 3245
rect 58420 3195 58430 3215
rect 58450 3195 58460 3215
rect 58420 3165 58460 3195
rect 58420 3145 58430 3165
rect 58450 3145 58460 3165
rect 58420 3115 58460 3145
rect 58420 3095 58430 3115
rect 58450 3095 58460 3115
rect 58420 3065 58460 3095
rect 58420 3045 58430 3065
rect 58450 3045 58460 3065
rect 58420 3015 58460 3045
rect 58420 2995 58430 3015
rect 58450 2995 58460 3015
rect 58420 2965 58460 2995
rect 58420 2945 58430 2965
rect 58450 2945 58460 2965
rect 58420 2915 58460 2945
rect 58420 2895 58430 2915
rect 58450 2895 58460 2915
rect 58420 2865 58460 2895
rect 58420 2845 58430 2865
rect 58450 2845 58460 2865
rect 58420 2815 58460 2845
rect 58420 2795 58430 2815
rect 58450 2795 58460 2815
rect 58420 2765 58460 2795
rect 58420 2745 58430 2765
rect 58450 2745 58460 2765
rect 58420 2730 58460 2745
rect 58475 3315 58515 3330
rect 58475 3295 58485 3315
rect 58505 3295 58515 3315
rect 58475 3265 58515 3295
rect 58475 3245 58485 3265
rect 58505 3245 58515 3265
rect 58475 3215 58515 3245
rect 58475 3195 58485 3215
rect 58505 3195 58515 3215
rect 58475 3165 58515 3195
rect 58475 3145 58485 3165
rect 58505 3145 58515 3165
rect 58475 3115 58515 3145
rect 58475 3095 58485 3115
rect 58505 3095 58515 3115
rect 58475 3065 58515 3095
rect 58475 3045 58485 3065
rect 58505 3045 58515 3065
rect 58475 3015 58515 3045
rect 58475 2995 58485 3015
rect 58505 2995 58515 3015
rect 58475 2965 58515 2995
rect 58475 2945 58485 2965
rect 58505 2945 58515 2965
rect 58475 2915 58515 2945
rect 58475 2895 58485 2915
rect 58505 2895 58515 2915
rect 58475 2865 58515 2895
rect 58475 2845 58485 2865
rect 58505 2845 58515 2865
rect 58475 2815 58515 2845
rect 58475 2795 58485 2815
rect 58505 2795 58515 2815
rect 58475 2765 58515 2795
rect 58475 2745 58485 2765
rect 58505 2745 58515 2765
rect 58475 2730 58515 2745
rect 58530 3315 58570 3330
rect 58530 3295 58540 3315
rect 58560 3295 58570 3315
rect 58530 3265 58570 3295
rect 58530 3245 58540 3265
rect 58560 3245 58570 3265
rect 58530 3215 58570 3245
rect 58530 3195 58540 3215
rect 58560 3195 58570 3215
rect 58530 3165 58570 3195
rect 58530 3145 58540 3165
rect 58560 3145 58570 3165
rect 58530 3115 58570 3145
rect 58530 3095 58540 3115
rect 58560 3095 58570 3115
rect 58530 3065 58570 3095
rect 58530 3045 58540 3065
rect 58560 3045 58570 3065
rect 58530 3015 58570 3045
rect 58530 2995 58540 3015
rect 58560 2995 58570 3015
rect 58530 2965 58570 2995
rect 58530 2945 58540 2965
rect 58560 2945 58570 2965
rect 58530 2915 58570 2945
rect 58530 2895 58540 2915
rect 58560 2895 58570 2915
rect 58530 2865 58570 2895
rect 58530 2845 58540 2865
rect 58560 2845 58570 2865
rect 58530 2815 58570 2845
rect 58530 2795 58540 2815
rect 58560 2795 58570 2815
rect 58530 2765 58570 2795
rect 58530 2745 58540 2765
rect 58560 2745 58570 2765
rect 58530 2730 58570 2745
rect 58585 3315 58625 3330
rect 58585 3295 58595 3315
rect 58615 3295 58625 3315
rect 58585 3265 58625 3295
rect 58585 3245 58595 3265
rect 58615 3245 58625 3265
rect 58585 3215 58625 3245
rect 58585 3195 58595 3215
rect 58615 3195 58625 3215
rect 58585 3165 58625 3195
rect 58585 3145 58595 3165
rect 58615 3145 58625 3165
rect 58585 3115 58625 3145
rect 58585 3095 58595 3115
rect 58615 3095 58625 3115
rect 58585 3065 58625 3095
rect 58585 3045 58595 3065
rect 58615 3045 58625 3065
rect 58585 3015 58625 3045
rect 58585 2995 58595 3015
rect 58615 2995 58625 3015
rect 58585 2965 58625 2995
rect 58585 2945 58595 2965
rect 58615 2945 58625 2965
rect 58585 2915 58625 2945
rect 58585 2895 58595 2915
rect 58615 2895 58625 2915
rect 58585 2865 58625 2895
rect 58585 2845 58595 2865
rect 58615 2845 58625 2865
rect 58585 2815 58625 2845
rect 58585 2795 58595 2815
rect 58615 2795 58625 2815
rect 58585 2765 58625 2795
rect 58585 2745 58595 2765
rect 58615 2745 58625 2765
rect 58585 2730 58625 2745
rect 58640 3315 58680 3330
rect 58640 3295 58650 3315
rect 58670 3295 58680 3315
rect 58640 3265 58680 3295
rect 58640 3245 58650 3265
rect 58670 3245 58680 3265
rect 58640 3215 58680 3245
rect 58640 3195 58650 3215
rect 58670 3195 58680 3215
rect 58640 3165 58680 3195
rect 58640 3145 58650 3165
rect 58670 3145 58680 3165
rect 58640 3115 58680 3145
rect 58640 3095 58650 3115
rect 58670 3095 58680 3115
rect 58640 3065 58680 3095
rect 58640 3045 58650 3065
rect 58670 3045 58680 3065
rect 58640 3015 58680 3045
rect 58640 2995 58650 3015
rect 58670 2995 58680 3015
rect 58640 2965 58680 2995
rect 58640 2945 58650 2965
rect 58670 2945 58680 2965
rect 58640 2915 58680 2945
rect 58640 2895 58650 2915
rect 58670 2895 58680 2915
rect 58640 2865 58680 2895
rect 58640 2845 58650 2865
rect 58670 2845 58680 2865
rect 58640 2815 58680 2845
rect 58640 2795 58650 2815
rect 58670 2795 58680 2815
rect 58640 2765 58680 2795
rect 58640 2745 58650 2765
rect 58670 2745 58680 2765
rect 58640 2730 58680 2745
rect 58695 3315 58735 3330
rect 58695 3295 58705 3315
rect 58725 3295 58735 3315
rect 58695 3265 58735 3295
rect 58695 3245 58705 3265
rect 58725 3245 58735 3265
rect 58695 3215 58735 3245
rect 58695 3195 58705 3215
rect 58725 3195 58735 3215
rect 58695 3165 58735 3195
rect 58695 3145 58705 3165
rect 58725 3145 58735 3165
rect 58695 3115 58735 3145
rect 58695 3095 58705 3115
rect 58725 3095 58735 3115
rect 58695 3065 58735 3095
rect 58695 3045 58705 3065
rect 58725 3045 58735 3065
rect 58695 3015 58735 3045
rect 58695 2995 58705 3015
rect 58725 2995 58735 3015
rect 58695 2965 58735 2995
rect 58695 2945 58705 2965
rect 58725 2945 58735 2965
rect 58695 2915 58735 2945
rect 58695 2895 58705 2915
rect 58725 2895 58735 2915
rect 58695 2865 58735 2895
rect 58695 2845 58705 2865
rect 58725 2845 58735 2865
rect 58695 2815 58735 2845
rect 58695 2795 58705 2815
rect 58725 2795 58735 2815
rect 58695 2765 58735 2795
rect 58695 2745 58705 2765
rect 58725 2745 58735 2765
rect 58695 2730 58735 2745
rect 58750 3315 58790 3330
rect 58750 3295 58760 3315
rect 58780 3295 58790 3315
rect 58750 3265 58790 3295
rect 58750 3245 58760 3265
rect 58780 3245 58790 3265
rect 58750 3215 58790 3245
rect 58750 3195 58760 3215
rect 58780 3195 58790 3215
rect 58750 3165 58790 3195
rect 58750 3145 58760 3165
rect 58780 3145 58790 3165
rect 58750 3115 58790 3145
rect 58750 3095 58760 3115
rect 58780 3095 58790 3115
rect 58750 3065 58790 3095
rect 58750 3045 58760 3065
rect 58780 3045 58790 3065
rect 58750 3015 58790 3045
rect 58750 2995 58760 3015
rect 58780 2995 58790 3015
rect 58750 2965 58790 2995
rect 58750 2945 58760 2965
rect 58780 2945 58790 2965
rect 58750 2915 58790 2945
rect 58750 2895 58760 2915
rect 58780 2895 58790 2915
rect 58750 2865 58790 2895
rect 58750 2845 58760 2865
rect 58780 2845 58790 2865
rect 58750 2815 58790 2845
rect 58750 2795 58760 2815
rect 58780 2795 58790 2815
rect 58750 2765 58790 2795
rect 58750 2745 58760 2765
rect 58780 2745 58790 2765
rect 58750 2730 58790 2745
rect 58805 3315 58845 3330
rect 58805 3295 58815 3315
rect 58835 3295 58845 3315
rect 58805 3265 58845 3295
rect 58805 3245 58815 3265
rect 58835 3245 58845 3265
rect 58805 3215 58845 3245
rect 58805 3195 58815 3215
rect 58835 3195 58845 3215
rect 58805 3165 58845 3195
rect 58805 3145 58815 3165
rect 58835 3145 58845 3165
rect 58805 3115 58845 3145
rect 58805 3095 58815 3115
rect 58835 3095 58845 3115
rect 58805 3065 58845 3095
rect 58805 3045 58815 3065
rect 58835 3045 58845 3065
rect 58805 3015 58845 3045
rect 58805 2995 58815 3015
rect 58835 2995 58845 3015
rect 58805 2965 58845 2995
rect 58805 2945 58815 2965
rect 58835 2945 58845 2965
rect 58805 2915 58845 2945
rect 58805 2895 58815 2915
rect 58835 2895 58845 2915
rect 58805 2865 58845 2895
rect 58805 2845 58815 2865
rect 58835 2845 58845 2865
rect 58805 2815 58845 2845
rect 58805 2795 58815 2815
rect 58835 2795 58845 2815
rect 58805 2765 58845 2795
rect 58805 2745 58815 2765
rect 58835 2745 58845 2765
rect 58805 2730 58845 2745
rect 54955 2355 54995 2370
rect 54955 2335 54965 2355
rect 54985 2335 54995 2355
rect 54955 2305 54995 2335
rect 54955 2285 54965 2305
rect 54985 2285 54995 2305
rect 54955 2255 54995 2285
rect 54955 2235 54965 2255
rect 54985 2235 54995 2255
rect 54955 2205 54995 2235
rect 54955 2185 54965 2205
rect 54985 2185 54995 2205
rect 54955 2170 54995 2185
rect 55010 2355 55050 2370
rect 55010 2335 55020 2355
rect 55040 2335 55050 2355
rect 55010 2305 55050 2335
rect 55010 2285 55020 2305
rect 55040 2285 55050 2305
rect 55010 2255 55050 2285
rect 55010 2235 55020 2255
rect 55040 2235 55050 2255
rect 55010 2205 55050 2235
rect 55010 2185 55020 2205
rect 55040 2185 55050 2205
rect 55010 2170 55050 2185
rect 55065 2355 55105 2370
rect 55065 2335 55075 2355
rect 55095 2335 55105 2355
rect 55065 2305 55105 2335
rect 55065 2285 55075 2305
rect 55095 2285 55105 2305
rect 55065 2255 55105 2285
rect 55065 2235 55075 2255
rect 55095 2235 55105 2255
rect 55065 2205 55105 2235
rect 55065 2185 55075 2205
rect 55095 2185 55105 2205
rect 55065 2170 55105 2185
rect 55120 2355 55160 2370
rect 55120 2335 55130 2355
rect 55150 2335 55160 2355
rect 55120 2305 55160 2335
rect 55120 2285 55130 2305
rect 55150 2285 55160 2305
rect 55120 2255 55160 2285
rect 55120 2235 55130 2255
rect 55150 2235 55160 2255
rect 55120 2205 55160 2235
rect 55120 2185 55130 2205
rect 55150 2185 55160 2205
rect 55120 2170 55160 2185
rect 55175 2355 55215 2370
rect 55175 2335 55185 2355
rect 55205 2335 55215 2355
rect 55175 2305 55215 2335
rect 55175 2285 55185 2305
rect 55205 2285 55215 2305
rect 55175 2255 55215 2285
rect 55175 2235 55185 2255
rect 55205 2235 55215 2255
rect 55175 2205 55215 2235
rect 55175 2185 55185 2205
rect 55205 2185 55215 2205
rect 55175 2170 55215 2185
rect 55230 2355 55270 2370
rect 55230 2335 55240 2355
rect 55260 2335 55270 2355
rect 55230 2305 55270 2335
rect 55230 2285 55240 2305
rect 55260 2285 55270 2305
rect 55230 2255 55270 2285
rect 55230 2235 55240 2255
rect 55260 2235 55270 2255
rect 55230 2205 55270 2235
rect 55230 2185 55240 2205
rect 55260 2185 55270 2205
rect 55230 2170 55270 2185
rect 55285 2355 55325 2370
rect 55285 2335 55295 2355
rect 55315 2335 55325 2355
rect 55285 2305 55325 2335
rect 55285 2285 55295 2305
rect 55315 2285 55325 2305
rect 55285 2255 55325 2285
rect 55285 2235 55295 2255
rect 55315 2235 55325 2255
rect 55285 2205 55325 2235
rect 55285 2185 55295 2205
rect 55315 2185 55325 2205
rect 55285 2170 55325 2185
rect 55340 2355 55380 2370
rect 55340 2335 55350 2355
rect 55370 2335 55380 2355
rect 55340 2305 55380 2335
rect 55340 2285 55350 2305
rect 55370 2285 55380 2305
rect 55340 2255 55380 2285
rect 55340 2235 55350 2255
rect 55370 2235 55380 2255
rect 55340 2205 55380 2235
rect 55340 2185 55350 2205
rect 55370 2185 55380 2205
rect 55340 2170 55380 2185
rect 55395 2355 55435 2370
rect 55395 2335 55405 2355
rect 55425 2335 55435 2355
rect 55395 2305 55435 2335
rect 55395 2285 55405 2305
rect 55425 2285 55435 2305
rect 55395 2255 55435 2285
rect 55395 2235 55405 2255
rect 55425 2235 55435 2255
rect 55395 2205 55435 2235
rect 55395 2185 55405 2205
rect 55425 2185 55435 2205
rect 55395 2170 55435 2185
rect 55450 2355 55490 2370
rect 55450 2335 55460 2355
rect 55480 2335 55490 2355
rect 55450 2305 55490 2335
rect 55450 2285 55460 2305
rect 55480 2285 55490 2305
rect 55450 2255 55490 2285
rect 55450 2235 55460 2255
rect 55480 2235 55490 2255
rect 55450 2205 55490 2235
rect 55450 2185 55460 2205
rect 55480 2185 55490 2205
rect 55450 2170 55490 2185
rect 55505 2355 55545 2370
rect 55505 2335 55515 2355
rect 55535 2335 55545 2355
rect 55505 2305 55545 2335
rect 55505 2285 55515 2305
rect 55535 2285 55545 2305
rect 55505 2255 55545 2285
rect 55505 2235 55515 2255
rect 55535 2235 55545 2255
rect 55505 2205 55545 2235
rect 55505 2185 55515 2205
rect 55535 2185 55545 2205
rect 55505 2170 55545 2185
rect 55560 2355 55600 2370
rect 55560 2335 55570 2355
rect 55590 2335 55600 2355
rect 55560 2305 55600 2335
rect 55560 2285 55570 2305
rect 55590 2285 55600 2305
rect 55560 2255 55600 2285
rect 55560 2235 55570 2255
rect 55590 2235 55600 2255
rect 55560 2205 55600 2235
rect 55560 2185 55570 2205
rect 55590 2185 55600 2205
rect 55560 2170 55600 2185
rect 55615 2355 55655 2370
rect 55615 2335 55625 2355
rect 55645 2335 55655 2355
rect 55615 2305 55655 2335
rect 55615 2285 55625 2305
rect 55645 2285 55655 2305
rect 55615 2255 55655 2285
rect 55615 2235 55625 2255
rect 55645 2235 55655 2255
rect 55615 2205 55655 2235
rect 55615 2185 55625 2205
rect 55645 2185 55655 2205
rect 55615 2170 55655 2185
rect 58145 2355 58185 2370
rect 58145 2335 58155 2355
rect 58175 2335 58185 2355
rect 58145 2305 58185 2335
rect 58145 2285 58155 2305
rect 58175 2285 58185 2305
rect 58145 2255 58185 2285
rect 58145 2235 58155 2255
rect 58175 2235 58185 2255
rect 58145 2205 58185 2235
rect 58145 2185 58155 2205
rect 58175 2185 58185 2205
rect 58145 2170 58185 2185
rect 58200 2355 58240 2370
rect 58200 2335 58210 2355
rect 58230 2335 58240 2355
rect 58200 2305 58240 2335
rect 58200 2285 58210 2305
rect 58230 2285 58240 2305
rect 58200 2255 58240 2285
rect 58200 2235 58210 2255
rect 58230 2235 58240 2255
rect 58200 2205 58240 2235
rect 58200 2185 58210 2205
rect 58230 2185 58240 2205
rect 58200 2170 58240 2185
rect 58255 2355 58295 2370
rect 58255 2335 58265 2355
rect 58285 2335 58295 2355
rect 58255 2305 58295 2335
rect 58255 2285 58265 2305
rect 58285 2285 58295 2305
rect 58255 2255 58295 2285
rect 58255 2235 58265 2255
rect 58285 2235 58295 2255
rect 58255 2205 58295 2235
rect 58255 2185 58265 2205
rect 58285 2185 58295 2205
rect 58255 2170 58295 2185
rect 58310 2355 58350 2370
rect 58310 2335 58320 2355
rect 58340 2335 58350 2355
rect 58310 2305 58350 2335
rect 58310 2285 58320 2305
rect 58340 2285 58350 2305
rect 58310 2255 58350 2285
rect 58310 2235 58320 2255
rect 58340 2235 58350 2255
rect 58310 2205 58350 2235
rect 58310 2185 58320 2205
rect 58340 2185 58350 2205
rect 58310 2170 58350 2185
rect 58365 2355 58405 2370
rect 58365 2335 58375 2355
rect 58395 2335 58405 2355
rect 58365 2305 58405 2335
rect 58365 2285 58375 2305
rect 58395 2285 58405 2305
rect 58365 2255 58405 2285
rect 58365 2235 58375 2255
rect 58395 2235 58405 2255
rect 58365 2205 58405 2235
rect 58365 2185 58375 2205
rect 58395 2185 58405 2205
rect 58365 2170 58405 2185
rect 58420 2355 58460 2370
rect 58420 2335 58430 2355
rect 58450 2335 58460 2355
rect 58420 2305 58460 2335
rect 58420 2285 58430 2305
rect 58450 2285 58460 2305
rect 58420 2255 58460 2285
rect 58420 2235 58430 2255
rect 58450 2235 58460 2255
rect 58420 2205 58460 2235
rect 58420 2185 58430 2205
rect 58450 2185 58460 2205
rect 58420 2170 58460 2185
rect 58475 2355 58515 2370
rect 58475 2335 58485 2355
rect 58505 2335 58515 2355
rect 58475 2305 58515 2335
rect 58475 2285 58485 2305
rect 58505 2285 58515 2305
rect 58475 2255 58515 2285
rect 58475 2235 58485 2255
rect 58505 2235 58515 2255
rect 58475 2205 58515 2235
rect 58475 2185 58485 2205
rect 58505 2185 58515 2205
rect 58475 2170 58515 2185
rect 58530 2355 58570 2370
rect 58530 2335 58540 2355
rect 58560 2335 58570 2355
rect 58530 2305 58570 2335
rect 58530 2285 58540 2305
rect 58560 2285 58570 2305
rect 58530 2255 58570 2285
rect 58530 2235 58540 2255
rect 58560 2235 58570 2255
rect 58530 2205 58570 2235
rect 58530 2185 58540 2205
rect 58560 2185 58570 2205
rect 58530 2170 58570 2185
rect 58585 2355 58625 2370
rect 58585 2335 58595 2355
rect 58615 2335 58625 2355
rect 58585 2305 58625 2335
rect 58585 2285 58595 2305
rect 58615 2285 58625 2305
rect 58585 2255 58625 2285
rect 58585 2235 58595 2255
rect 58615 2235 58625 2255
rect 58585 2205 58625 2235
rect 58585 2185 58595 2205
rect 58615 2185 58625 2205
rect 58585 2170 58625 2185
rect 58640 2355 58680 2370
rect 58640 2335 58650 2355
rect 58670 2335 58680 2355
rect 58640 2305 58680 2335
rect 58640 2285 58650 2305
rect 58670 2285 58680 2305
rect 58640 2255 58680 2285
rect 58640 2235 58650 2255
rect 58670 2235 58680 2255
rect 58640 2205 58680 2235
rect 58640 2185 58650 2205
rect 58670 2185 58680 2205
rect 58640 2170 58680 2185
rect 58695 2355 58735 2370
rect 58695 2335 58705 2355
rect 58725 2335 58735 2355
rect 58695 2305 58735 2335
rect 58695 2285 58705 2305
rect 58725 2285 58735 2305
rect 58695 2255 58735 2285
rect 58695 2235 58705 2255
rect 58725 2235 58735 2255
rect 58695 2205 58735 2235
rect 58695 2185 58705 2205
rect 58725 2185 58735 2205
rect 58695 2170 58735 2185
rect 58750 2355 58790 2370
rect 58750 2335 58760 2355
rect 58780 2335 58790 2355
rect 58750 2305 58790 2335
rect 58750 2285 58760 2305
rect 58780 2285 58790 2305
rect 58750 2255 58790 2285
rect 58750 2235 58760 2255
rect 58780 2235 58790 2255
rect 58750 2205 58790 2235
rect 58750 2185 58760 2205
rect 58780 2185 58790 2205
rect 58750 2170 58790 2185
rect 58805 2355 58845 2370
rect 58805 2335 58815 2355
rect 58835 2335 58845 2355
rect 58805 2305 58845 2335
rect 58805 2285 58815 2305
rect 58835 2285 58845 2305
rect 58805 2255 58845 2285
rect 58805 2235 58815 2255
rect 58835 2235 58845 2255
rect 58805 2205 58845 2235
rect 58805 2185 58815 2205
rect 58835 2185 58845 2205
rect 58805 2170 58845 2185
<< ndiffc >>
rect 56560 2425 56580 2445
rect 56615 2425 56635 2445
rect 56670 2425 56690 2445
rect 56725 2425 56745 2445
rect 56780 2425 56800 2445
rect 56835 2425 56855 2445
rect 56890 2425 56910 2445
rect 56945 2425 56965 2445
rect 57000 2425 57020 2445
rect 57055 2425 57075 2445
rect 57110 2425 57130 2445
rect 57165 2425 57185 2445
rect 57220 2425 57240 2445
rect 54965 1875 54985 1895
rect 54965 1825 54985 1845
rect 54965 1775 54985 1795
rect 54965 1725 54985 1745
rect 54965 1675 54985 1695
rect 54965 1625 54985 1645
rect 55020 1875 55040 1895
rect 55020 1825 55040 1845
rect 55020 1775 55040 1795
rect 55020 1725 55040 1745
rect 55020 1675 55040 1695
rect 55020 1625 55040 1645
rect 55075 1875 55095 1895
rect 55075 1825 55095 1845
rect 55075 1775 55095 1795
rect 55075 1725 55095 1745
rect 55075 1675 55095 1695
rect 55075 1625 55095 1645
rect 55130 1875 55150 1895
rect 55130 1825 55150 1845
rect 55130 1775 55150 1795
rect 55130 1725 55150 1745
rect 55130 1675 55150 1695
rect 55130 1625 55150 1645
rect 55185 1875 55205 1895
rect 55185 1825 55205 1845
rect 55185 1775 55205 1795
rect 55185 1725 55205 1745
rect 55185 1675 55205 1695
rect 55185 1625 55205 1645
rect 55240 1875 55260 1895
rect 55240 1825 55260 1845
rect 55240 1775 55260 1795
rect 55240 1725 55260 1745
rect 55240 1675 55260 1695
rect 55240 1625 55260 1645
rect 55295 1875 55315 1895
rect 55295 1825 55315 1845
rect 55295 1775 55315 1795
rect 55295 1725 55315 1745
rect 55295 1675 55315 1695
rect 55295 1625 55315 1645
rect 55350 1875 55370 1895
rect 55350 1825 55370 1845
rect 55350 1775 55370 1795
rect 55350 1725 55370 1745
rect 55350 1675 55370 1695
rect 55350 1625 55370 1645
rect 55405 1875 55425 1895
rect 55405 1825 55425 1845
rect 55405 1775 55425 1795
rect 55405 1725 55425 1745
rect 55405 1675 55425 1695
rect 55405 1625 55425 1645
rect 55460 1875 55480 1895
rect 55460 1825 55480 1845
rect 55460 1775 55480 1795
rect 55460 1725 55480 1745
rect 55460 1675 55480 1695
rect 55460 1625 55480 1645
rect 55515 1875 55535 1895
rect 55515 1825 55535 1845
rect 55515 1775 55535 1795
rect 55515 1725 55535 1745
rect 55515 1675 55535 1695
rect 55515 1625 55535 1645
rect 55570 1875 55590 1895
rect 55570 1825 55590 1845
rect 55570 1775 55590 1795
rect 55570 1725 55590 1745
rect 55570 1675 55590 1695
rect 55570 1625 55590 1645
rect 55625 1875 55645 1895
rect 55625 1825 55645 1845
rect 55625 1775 55645 1795
rect 55625 1725 55645 1745
rect 55625 1675 55645 1695
rect 55625 1625 55645 1645
rect 56085 2145 56105 2165
rect 56085 2095 56105 2115
rect 56085 2045 56105 2065
rect 56140 2145 56160 2165
rect 56140 2095 56160 2115
rect 56140 2045 56160 2065
rect 56195 2145 56215 2165
rect 56195 2095 56215 2115
rect 56195 2045 56215 2065
rect 56250 2145 56270 2165
rect 56250 2095 56270 2115
rect 56250 2045 56270 2065
rect 56305 2145 56325 2165
rect 56305 2095 56325 2115
rect 56305 2045 56325 2065
rect 56360 2145 56380 2165
rect 56360 2095 56380 2115
rect 56360 2045 56380 2065
rect 56415 2145 56435 2165
rect 56415 2095 56435 2115
rect 56415 2045 56435 2065
rect 56470 2145 56490 2165
rect 56470 2095 56490 2115
rect 56470 2045 56490 2065
rect 56525 2145 56545 2165
rect 56525 2095 56545 2115
rect 56525 2045 56545 2065
rect 56580 2145 56600 2165
rect 56580 2095 56600 2115
rect 56580 2045 56600 2065
rect 56635 2145 56655 2165
rect 56635 2095 56655 2115
rect 56635 2045 56655 2065
rect 56690 2145 56710 2165
rect 56690 2095 56710 2115
rect 56690 2045 56710 2065
rect 56745 2145 56765 2165
rect 56745 2095 56765 2115
rect 56745 2045 56765 2065
rect 57035 2145 57055 2165
rect 57035 2095 57055 2115
rect 57035 2045 57055 2065
rect 57090 2145 57110 2165
rect 57090 2095 57110 2115
rect 57090 2045 57110 2065
rect 57145 2145 57165 2165
rect 57145 2095 57165 2115
rect 57145 2045 57165 2065
rect 57200 2145 57220 2165
rect 57200 2095 57220 2115
rect 57200 2045 57220 2065
rect 57255 2145 57275 2165
rect 57255 2095 57275 2115
rect 57255 2045 57275 2065
rect 57310 2145 57330 2165
rect 57310 2095 57330 2115
rect 57310 2045 57330 2065
rect 57365 2145 57385 2165
rect 57365 2095 57385 2115
rect 57365 2045 57385 2065
rect 57420 2145 57440 2165
rect 57420 2095 57440 2115
rect 57420 2045 57440 2065
rect 57475 2145 57495 2165
rect 57475 2095 57495 2115
rect 57475 2045 57495 2065
rect 57530 2145 57550 2165
rect 57530 2095 57550 2115
rect 57530 2045 57550 2065
rect 57585 2145 57605 2165
rect 57585 2095 57605 2115
rect 57585 2045 57605 2065
rect 57640 2145 57660 2165
rect 57640 2095 57660 2115
rect 57640 2045 57660 2065
rect 57695 2145 57715 2165
rect 57695 2095 57715 2115
rect 57695 2045 57715 2065
rect 56040 1675 56060 1695
rect 56040 1625 56060 1645
rect 56040 1575 56060 1595
rect 56095 1675 56115 1695
rect 56095 1625 56115 1645
rect 56095 1575 56115 1595
rect 56150 1675 56170 1695
rect 56150 1625 56170 1645
rect 56150 1575 56170 1595
rect 56205 1675 56225 1695
rect 56205 1625 56225 1645
rect 56205 1575 56225 1595
rect 56260 1675 56280 1695
rect 56260 1625 56280 1645
rect 56260 1575 56280 1595
rect 56315 1675 56335 1695
rect 56315 1625 56335 1645
rect 56315 1575 56335 1595
rect 56370 1675 56390 1695
rect 56370 1625 56390 1645
rect 56370 1575 56390 1595
rect 56425 1675 56445 1695
rect 56425 1625 56445 1645
rect 56425 1575 56445 1595
rect 56480 1675 56500 1695
rect 56480 1625 56500 1645
rect 56480 1575 56500 1595
rect 56535 1675 56555 1695
rect 56535 1625 56555 1645
rect 56535 1575 56555 1595
rect 56590 1675 56610 1695
rect 56590 1625 56610 1645
rect 56590 1575 56610 1595
rect 56645 1675 56665 1695
rect 56645 1625 56665 1645
rect 56645 1575 56665 1595
rect 56700 1675 56720 1695
rect 56700 1625 56720 1645
rect 56700 1575 56720 1595
rect 56780 1675 56800 1695
rect 56780 1625 56800 1645
rect 56780 1575 56800 1595
rect 56835 1675 56855 1695
rect 56835 1625 56855 1645
rect 56835 1575 56855 1595
rect 56890 1675 56910 1695
rect 56890 1625 56910 1645
rect 56890 1575 56910 1595
rect 56945 1675 56965 1695
rect 56945 1625 56965 1645
rect 56945 1575 56965 1595
rect 57000 1675 57020 1695
rect 57000 1625 57020 1645
rect 57000 1575 57020 1595
rect 57080 1675 57100 1695
rect 57080 1625 57100 1645
rect 57080 1575 57100 1595
rect 57135 1675 57155 1695
rect 57135 1625 57155 1645
rect 57135 1575 57155 1595
rect 57190 1675 57210 1695
rect 57190 1625 57210 1645
rect 57190 1575 57210 1595
rect 57245 1675 57265 1695
rect 57245 1625 57265 1645
rect 57245 1575 57265 1595
rect 57300 1675 57320 1695
rect 57300 1625 57320 1645
rect 57300 1575 57320 1595
rect 57355 1675 57375 1695
rect 57355 1625 57375 1645
rect 57355 1575 57375 1595
rect 57410 1675 57430 1695
rect 57410 1625 57430 1645
rect 57410 1575 57430 1595
rect 57465 1675 57485 1695
rect 57465 1625 57485 1645
rect 57465 1575 57485 1595
rect 57520 1675 57540 1695
rect 57520 1625 57540 1645
rect 57520 1575 57540 1595
rect 57575 1675 57595 1695
rect 57575 1625 57595 1645
rect 57575 1575 57595 1595
rect 57630 1675 57650 1695
rect 57630 1625 57650 1645
rect 57630 1575 57650 1595
rect 57685 1675 57705 1695
rect 57685 1625 57705 1645
rect 57685 1575 57705 1595
rect 57740 1675 57760 1695
rect 57740 1625 57760 1645
rect 57740 1575 57760 1595
rect 58155 1875 58175 1895
rect 58155 1825 58175 1845
rect 58155 1775 58175 1795
rect 58155 1725 58175 1745
rect 58155 1675 58175 1695
rect 58155 1625 58175 1645
rect 58210 1875 58230 1895
rect 58210 1825 58230 1845
rect 58210 1775 58230 1795
rect 58210 1725 58230 1745
rect 58210 1675 58230 1695
rect 58210 1625 58230 1645
rect 58265 1875 58285 1895
rect 58265 1825 58285 1845
rect 58265 1775 58285 1795
rect 58265 1725 58285 1745
rect 58265 1675 58285 1695
rect 58265 1625 58285 1645
rect 58320 1875 58340 1895
rect 58320 1825 58340 1845
rect 58320 1775 58340 1795
rect 58320 1725 58340 1745
rect 58320 1675 58340 1695
rect 58320 1625 58340 1645
rect 58375 1875 58395 1895
rect 58375 1825 58395 1845
rect 58375 1775 58395 1795
rect 58375 1725 58395 1745
rect 58375 1675 58395 1695
rect 58375 1625 58395 1645
rect 58430 1875 58450 1895
rect 58430 1825 58450 1845
rect 58430 1775 58450 1795
rect 58430 1725 58450 1745
rect 58430 1675 58450 1695
rect 58430 1625 58450 1645
rect 58485 1875 58505 1895
rect 58485 1825 58505 1845
rect 58485 1775 58505 1795
rect 58485 1725 58505 1745
rect 58485 1675 58505 1695
rect 58485 1625 58505 1645
rect 58540 1875 58560 1895
rect 58540 1825 58560 1845
rect 58540 1775 58560 1795
rect 58540 1725 58560 1745
rect 58540 1675 58560 1695
rect 58540 1625 58560 1645
rect 58595 1875 58615 1895
rect 58595 1825 58615 1845
rect 58595 1775 58615 1795
rect 58595 1725 58615 1745
rect 58595 1675 58615 1695
rect 58595 1625 58615 1645
rect 58650 1875 58670 1895
rect 58650 1825 58670 1845
rect 58650 1775 58670 1795
rect 58650 1725 58670 1745
rect 58650 1675 58670 1695
rect 58650 1625 58670 1645
rect 58705 1875 58725 1895
rect 58705 1825 58725 1845
rect 58705 1775 58725 1795
rect 58705 1725 58725 1745
rect 58705 1675 58725 1695
rect 58705 1625 58725 1645
rect 58760 1875 58780 1895
rect 58760 1825 58780 1845
rect 58760 1775 58780 1795
rect 58760 1725 58780 1745
rect 58760 1675 58780 1695
rect 58760 1625 58780 1645
rect 58815 1875 58835 1895
rect 58815 1825 58835 1845
rect 58815 1775 58835 1795
rect 58815 1725 58835 1745
rect 58815 1675 58835 1695
rect 58815 1625 58835 1645
rect 55045 1285 55065 1305
rect 55045 1235 55065 1255
rect 55045 1185 55065 1205
rect 55045 1135 55065 1155
rect 55045 1085 55065 1105
rect 55045 1035 55065 1055
rect 55045 985 55065 1005
rect 55045 935 55065 955
rect 55045 885 55065 905
rect 55045 835 55065 855
rect 55045 785 55065 805
rect 55045 735 55065 755
rect 55045 685 55065 705
rect 55045 635 55065 655
rect 55145 1285 55165 1305
rect 55145 1235 55165 1255
rect 55145 1185 55165 1205
rect 55145 1135 55165 1155
rect 55145 1085 55165 1105
rect 55145 1035 55165 1055
rect 55145 985 55165 1005
rect 55145 935 55165 955
rect 55145 885 55165 905
rect 55145 835 55165 855
rect 55145 785 55165 805
rect 55145 735 55165 755
rect 55145 685 55165 705
rect 55145 635 55165 655
rect 55245 1285 55265 1305
rect 55245 1235 55265 1255
rect 55245 1185 55265 1205
rect 55245 1135 55265 1155
rect 55245 1085 55265 1105
rect 55245 1035 55265 1055
rect 55245 985 55265 1005
rect 55245 935 55265 955
rect 55245 885 55265 905
rect 55245 835 55265 855
rect 55245 785 55265 805
rect 55245 735 55265 755
rect 55245 685 55265 705
rect 55245 635 55265 655
rect 55345 1285 55365 1305
rect 55345 1235 55365 1255
rect 55345 1185 55365 1205
rect 55345 1135 55365 1155
rect 55345 1085 55365 1105
rect 55345 1035 55365 1055
rect 55345 985 55365 1005
rect 55345 935 55365 955
rect 55345 885 55365 905
rect 55345 835 55365 855
rect 55345 785 55365 805
rect 55345 735 55365 755
rect 55345 685 55365 705
rect 55345 635 55365 655
rect 55445 1285 55465 1305
rect 55445 1235 55465 1255
rect 55445 1185 55465 1205
rect 55445 1135 55465 1155
rect 55445 1085 55465 1105
rect 55445 1035 55465 1055
rect 55445 985 55465 1005
rect 55445 935 55465 955
rect 55445 885 55465 905
rect 55445 835 55465 855
rect 55445 785 55465 805
rect 55445 735 55465 755
rect 55445 685 55465 705
rect 55445 635 55465 655
rect 55545 1285 55565 1305
rect 55545 1235 55565 1255
rect 55545 1185 55565 1205
rect 55545 1135 55565 1155
rect 55545 1085 55565 1105
rect 55545 1035 55565 1055
rect 55545 985 55565 1005
rect 55545 935 55565 955
rect 55545 885 55565 905
rect 55545 835 55565 855
rect 55545 785 55565 805
rect 55545 735 55565 755
rect 55545 685 55565 705
rect 55545 635 55565 655
rect 55645 1285 55665 1305
rect 55645 1235 55665 1255
rect 55645 1185 55665 1205
rect 55645 1135 55665 1155
rect 55645 1085 55665 1105
rect 55645 1035 55665 1055
rect 55645 985 55665 1005
rect 55645 935 55665 955
rect 55645 885 55665 905
rect 55645 835 55665 855
rect 55645 785 55665 805
rect 55645 735 55665 755
rect 55645 685 55665 705
rect 55645 635 55665 655
rect 56230 1170 56250 1190
rect 56230 1120 56250 1140
rect 56230 1070 56250 1090
rect 56230 1020 56250 1040
rect 56230 970 56250 990
rect 56285 1170 56305 1190
rect 56285 1120 56305 1140
rect 56285 1070 56305 1090
rect 56285 1020 56305 1040
rect 56285 970 56305 990
rect 56340 1170 56360 1190
rect 56340 1120 56360 1140
rect 56340 1070 56360 1090
rect 56340 1020 56360 1040
rect 56340 970 56360 990
rect 56395 1170 56415 1190
rect 56395 1120 56415 1140
rect 56395 1070 56415 1090
rect 56395 1020 56415 1040
rect 56395 970 56415 990
rect 56450 1170 56470 1190
rect 56450 1120 56470 1140
rect 56450 1070 56470 1090
rect 56450 1020 56470 1040
rect 56450 970 56470 990
rect 56505 1170 56525 1190
rect 56505 1120 56525 1140
rect 56505 1070 56525 1090
rect 56505 1020 56525 1040
rect 56505 970 56525 990
rect 56560 1170 56580 1190
rect 56560 1120 56580 1140
rect 56560 1070 56580 1090
rect 56560 1020 56580 1040
rect 56560 970 56580 990
rect 56615 1170 56635 1190
rect 56615 1120 56635 1140
rect 56615 1070 56635 1090
rect 56615 1020 56635 1040
rect 56615 970 56635 990
rect 56670 1170 56690 1190
rect 56670 1120 56690 1140
rect 56670 1070 56690 1090
rect 56670 1020 56690 1040
rect 56670 970 56690 990
rect 56725 1170 56745 1190
rect 56725 1120 56745 1140
rect 56725 1070 56745 1090
rect 56725 1020 56745 1040
rect 56725 970 56745 990
rect 56780 1170 56800 1190
rect 56780 1120 56800 1140
rect 56780 1070 56800 1090
rect 56780 1020 56800 1040
rect 56780 970 56800 990
rect 56835 1170 56855 1190
rect 56835 1120 56855 1140
rect 56835 1070 56855 1090
rect 56835 1020 56855 1040
rect 56835 970 56855 990
rect 56890 1170 56910 1190
rect 56890 1120 56910 1140
rect 56890 1070 56910 1090
rect 56890 1020 56910 1040
rect 56890 970 56910 990
rect 56945 1170 56965 1190
rect 56945 1120 56965 1140
rect 56945 1070 56965 1090
rect 56945 1020 56965 1040
rect 56945 970 56965 990
rect 57000 1170 57020 1190
rect 57000 1120 57020 1140
rect 57000 1070 57020 1090
rect 57000 1020 57020 1040
rect 57000 970 57020 990
rect 57055 1170 57075 1190
rect 57055 1120 57075 1140
rect 57055 1070 57075 1090
rect 57055 1020 57075 1040
rect 57055 970 57075 990
rect 57110 1170 57130 1190
rect 57110 1120 57130 1140
rect 57110 1070 57130 1090
rect 57110 1020 57130 1040
rect 57110 970 57130 990
rect 57165 1170 57185 1190
rect 57165 1120 57185 1140
rect 57165 1070 57185 1090
rect 57165 1020 57185 1040
rect 57165 970 57185 990
rect 57220 1170 57240 1190
rect 57220 1120 57240 1140
rect 57220 1070 57240 1090
rect 57220 1020 57240 1040
rect 57220 970 57240 990
rect 57275 1170 57295 1190
rect 57275 1120 57295 1140
rect 57275 1070 57295 1090
rect 57275 1020 57295 1040
rect 57275 970 57295 990
rect 57330 1170 57350 1190
rect 57330 1120 57350 1140
rect 57330 1070 57350 1090
rect 57330 1020 57350 1040
rect 57330 970 57350 990
rect 57385 1170 57405 1190
rect 57385 1120 57405 1140
rect 57385 1070 57405 1090
rect 57385 1020 57405 1040
rect 57385 970 57405 990
rect 57440 1170 57460 1190
rect 57440 1120 57460 1140
rect 57440 1070 57460 1090
rect 57440 1020 57460 1040
rect 57440 970 57460 990
rect 57495 1170 57515 1190
rect 57495 1120 57515 1140
rect 57495 1070 57515 1090
rect 57495 1020 57515 1040
rect 57495 970 57515 990
rect 57550 1170 57570 1190
rect 57550 1120 57570 1140
rect 57550 1070 57570 1090
rect 57550 1020 57570 1040
rect 57550 970 57570 990
rect 56720 655 56740 675
rect 56720 605 56740 625
rect 57050 655 57070 675
rect 57050 605 57070 625
rect 58135 1285 58155 1305
rect 58135 1235 58155 1255
rect 58135 1185 58155 1205
rect 58135 1135 58155 1155
rect 58135 1085 58155 1105
rect 58135 1035 58155 1055
rect 58135 985 58155 1005
rect 58135 935 58155 955
rect 58135 885 58155 905
rect 58135 835 58155 855
rect 58135 785 58155 805
rect 58135 735 58155 755
rect 58135 685 58155 705
rect 58135 635 58155 655
rect 58235 1285 58255 1305
rect 58235 1235 58255 1255
rect 58235 1185 58255 1205
rect 58235 1135 58255 1155
rect 58235 1085 58255 1105
rect 58235 1035 58255 1055
rect 58235 985 58255 1005
rect 58235 935 58255 955
rect 58235 885 58255 905
rect 58235 835 58255 855
rect 58235 785 58255 805
rect 58235 735 58255 755
rect 58235 685 58255 705
rect 58235 635 58255 655
rect 58335 1285 58355 1305
rect 58335 1235 58355 1255
rect 58335 1185 58355 1205
rect 58335 1135 58355 1155
rect 58335 1085 58355 1105
rect 58335 1035 58355 1055
rect 58335 985 58355 1005
rect 58335 935 58355 955
rect 58335 885 58355 905
rect 58335 835 58355 855
rect 58335 785 58355 805
rect 58335 735 58355 755
rect 58335 685 58355 705
rect 58335 635 58355 655
rect 58435 1285 58455 1305
rect 58435 1235 58455 1255
rect 58435 1185 58455 1205
rect 58435 1135 58455 1155
rect 58435 1085 58455 1105
rect 58435 1035 58455 1055
rect 58435 985 58455 1005
rect 58435 935 58455 955
rect 58435 885 58455 905
rect 58435 835 58455 855
rect 58435 785 58455 805
rect 58435 735 58455 755
rect 58435 685 58455 705
rect 58435 635 58455 655
rect 58535 1285 58555 1305
rect 58535 1235 58555 1255
rect 58535 1185 58555 1205
rect 58535 1135 58555 1155
rect 58535 1085 58555 1105
rect 58535 1035 58555 1055
rect 58535 985 58555 1005
rect 58535 935 58555 955
rect 58535 885 58555 905
rect 58535 835 58555 855
rect 58535 785 58555 805
rect 58535 735 58555 755
rect 58535 685 58555 705
rect 58535 635 58555 655
rect 58635 1285 58655 1305
rect 58635 1235 58655 1255
rect 58635 1185 58655 1205
rect 58635 1135 58655 1155
rect 58635 1085 58655 1105
rect 58635 1035 58655 1055
rect 58635 985 58655 1005
rect 58635 935 58655 955
rect 58635 885 58655 905
rect 58635 835 58655 855
rect 58635 785 58655 805
rect 58635 735 58655 755
rect 58635 685 58655 705
rect 58635 635 58655 655
rect 58735 1285 58755 1305
rect 58735 1235 58755 1255
rect 58735 1185 58755 1205
rect 58735 1135 58755 1155
rect 58735 1085 58755 1105
rect 58735 1035 58755 1055
rect 58735 985 58755 1005
rect 58735 935 58755 955
rect 58735 885 58755 905
rect 58735 835 58755 855
rect 58735 785 58755 805
rect 58735 735 58755 755
rect 58735 685 58755 705
rect 58735 635 58755 655
<< pdiffc >>
rect 56155 4430 56175 4450
rect 56215 4430 56235 4450
rect 56275 4430 56295 4450
rect 56335 4430 56355 4450
rect 56830 4435 56850 4705
rect 56890 4435 56910 4705
rect 56950 4435 56970 4705
rect 57010 4435 57030 4705
rect 57500 4435 57520 4745
rect 57560 4435 57580 4745
rect 57620 4435 57640 4745
rect 57680 4435 57700 4745
rect 54965 4005 54985 4025
rect 54965 3955 54985 3975
rect 54965 3905 54985 3925
rect 54965 3855 54985 3875
rect 54965 3805 54985 3825
rect 54965 3755 54985 3775
rect 54965 3705 54985 3725
rect 55025 4005 55045 4025
rect 55025 3955 55045 3975
rect 55025 3905 55045 3925
rect 55025 3855 55045 3875
rect 55025 3805 55045 3825
rect 55025 3755 55045 3775
rect 55025 3705 55045 3725
rect 55085 4005 55105 4025
rect 55085 3955 55105 3975
rect 55085 3905 55105 3925
rect 55085 3855 55105 3875
rect 55085 3805 55105 3825
rect 55085 3755 55105 3775
rect 55085 3705 55105 3725
rect 55145 4005 55165 4025
rect 55145 3955 55165 3975
rect 55145 3905 55165 3925
rect 55145 3855 55165 3875
rect 55145 3805 55165 3825
rect 55145 3755 55165 3775
rect 55145 3705 55165 3725
rect 55205 4005 55225 4025
rect 55205 3955 55225 3975
rect 55205 3905 55225 3925
rect 55205 3855 55225 3875
rect 55205 3805 55225 3825
rect 55205 3755 55225 3775
rect 55205 3705 55225 3725
rect 55265 4005 55285 4025
rect 55265 3955 55285 3975
rect 55265 3905 55285 3925
rect 55265 3855 55285 3875
rect 55265 3805 55285 3825
rect 55265 3755 55285 3775
rect 55265 3705 55285 3725
rect 55325 4005 55345 4025
rect 55325 3955 55345 3975
rect 55325 3905 55345 3925
rect 55325 3855 55345 3875
rect 55325 3805 55345 3825
rect 55325 3755 55345 3775
rect 55325 3705 55345 3725
rect 55385 4005 55405 4025
rect 55385 3955 55405 3975
rect 55385 3905 55405 3925
rect 55385 3855 55405 3875
rect 55385 3805 55405 3825
rect 55385 3755 55405 3775
rect 55385 3705 55405 3725
rect 55445 4005 55465 4025
rect 55445 3955 55465 3975
rect 55445 3905 55465 3925
rect 55445 3855 55465 3875
rect 55445 3805 55465 3825
rect 55445 3755 55465 3775
rect 55445 3705 55465 3725
rect 55505 4005 55525 4025
rect 55505 3955 55525 3975
rect 55505 3905 55525 3925
rect 55505 3855 55525 3875
rect 55505 3805 55525 3825
rect 55505 3755 55525 3775
rect 55505 3705 55525 3725
rect 55565 4005 55585 4025
rect 55565 3955 55585 3975
rect 55565 3905 55585 3925
rect 55565 3855 55585 3875
rect 55565 3805 55585 3825
rect 55565 3755 55585 3775
rect 55565 3705 55585 3725
rect 55625 4005 55645 4025
rect 55625 3955 55645 3975
rect 55625 3905 55645 3925
rect 55625 3855 55645 3875
rect 55625 3805 55645 3825
rect 55625 3755 55645 3775
rect 55625 3705 55645 3725
rect 55685 4005 55705 4025
rect 55685 3955 55705 3975
rect 55685 3905 55705 3925
rect 55685 3855 55705 3875
rect 55685 3805 55705 3825
rect 55685 3755 55705 3775
rect 55685 3705 55705 3725
rect 56015 4005 56035 4025
rect 56015 3955 56035 3975
rect 56015 3905 56035 3925
rect 56015 3855 56035 3875
rect 56015 3805 56035 3825
rect 56015 3755 56035 3775
rect 56015 3705 56035 3725
rect 56075 4005 56095 4025
rect 56075 3955 56095 3975
rect 56075 3905 56095 3925
rect 56075 3855 56095 3875
rect 56075 3805 56095 3825
rect 56075 3755 56095 3775
rect 56075 3705 56095 3725
rect 56135 4005 56155 4025
rect 56135 3955 56155 3975
rect 56135 3905 56155 3925
rect 56135 3855 56155 3875
rect 56135 3805 56155 3825
rect 56135 3755 56155 3775
rect 56135 3705 56155 3725
rect 56195 4005 56215 4025
rect 56195 3955 56215 3975
rect 56195 3905 56215 3925
rect 56195 3855 56215 3875
rect 56195 3805 56215 3825
rect 56195 3755 56215 3775
rect 56195 3705 56215 3725
rect 56255 4005 56275 4025
rect 56255 3955 56275 3975
rect 56255 3905 56275 3925
rect 56255 3855 56275 3875
rect 56255 3805 56275 3825
rect 56255 3755 56275 3775
rect 56255 3705 56275 3725
rect 56315 4005 56335 4025
rect 56315 3955 56335 3975
rect 56315 3905 56335 3925
rect 56315 3855 56335 3875
rect 56315 3805 56335 3825
rect 56315 3755 56335 3775
rect 56315 3705 56335 3725
rect 56375 4005 56395 4025
rect 56375 3955 56395 3975
rect 56375 3905 56395 3925
rect 56375 3855 56395 3875
rect 56375 3805 56395 3825
rect 56375 3755 56395 3775
rect 56375 3705 56395 3725
rect 56435 4005 56455 4025
rect 56435 3955 56455 3975
rect 56435 3905 56455 3925
rect 56435 3855 56455 3875
rect 56435 3805 56455 3825
rect 56435 3755 56455 3775
rect 56435 3705 56455 3725
rect 56495 4005 56515 4025
rect 56495 3955 56515 3975
rect 56495 3905 56515 3925
rect 56495 3855 56515 3875
rect 56495 3805 56515 3825
rect 56495 3755 56515 3775
rect 56495 3705 56515 3725
rect 56555 4005 56575 4025
rect 56555 3955 56575 3975
rect 56555 3905 56575 3925
rect 56555 3855 56575 3875
rect 56555 3805 56575 3825
rect 56555 3755 56575 3775
rect 56555 3705 56575 3725
rect 56615 4005 56635 4025
rect 56615 3955 56635 3975
rect 56615 3905 56635 3925
rect 56615 3855 56635 3875
rect 56615 3805 56635 3825
rect 56615 3755 56635 3775
rect 56615 3705 56635 3725
rect 56675 4005 56695 4025
rect 56675 3955 56695 3975
rect 56675 3905 56695 3925
rect 56675 3855 56695 3875
rect 56675 3805 56695 3825
rect 56675 3755 56695 3775
rect 56675 3705 56695 3725
rect 56735 4005 56755 4025
rect 56735 3955 56755 3975
rect 56735 3905 56755 3925
rect 56735 3855 56755 3875
rect 56735 3805 56755 3825
rect 56735 3755 56755 3775
rect 56735 3705 56755 3725
rect 57045 4005 57065 4025
rect 57045 3955 57065 3975
rect 57045 3905 57065 3925
rect 57045 3855 57065 3875
rect 57045 3805 57065 3825
rect 57045 3755 57065 3775
rect 57045 3705 57065 3725
rect 57105 4005 57125 4025
rect 57105 3955 57125 3975
rect 57105 3905 57125 3925
rect 57105 3855 57125 3875
rect 57105 3805 57125 3825
rect 57105 3755 57125 3775
rect 57105 3705 57125 3725
rect 57165 4005 57185 4025
rect 57165 3955 57185 3975
rect 57165 3905 57185 3925
rect 57165 3855 57185 3875
rect 57165 3805 57185 3825
rect 57165 3755 57185 3775
rect 57165 3705 57185 3725
rect 57225 4005 57245 4025
rect 57225 3955 57245 3975
rect 57225 3905 57245 3925
rect 57225 3855 57245 3875
rect 57225 3805 57245 3825
rect 57225 3755 57245 3775
rect 57225 3705 57245 3725
rect 57285 4005 57305 4025
rect 57285 3955 57305 3975
rect 57285 3905 57305 3925
rect 57285 3855 57305 3875
rect 57285 3805 57305 3825
rect 57285 3755 57305 3775
rect 57285 3705 57305 3725
rect 57345 4005 57365 4025
rect 57345 3955 57365 3975
rect 57345 3905 57365 3925
rect 57345 3855 57365 3875
rect 57345 3805 57365 3825
rect 57345 3755 57365 3775
rect 57345 3705 57365 3725
rect 57405 4005 57425 4025
rect 57405 3955 57425 3975
rect 57405 3905 57425 3925
rect 57405 3855 57425 3875
rect 57405 3805 57425 3825
rect 57405 3755 57425 3775
rect 57405 3705 57425 3725
rect 57465 4005 57485 4025
rect 57465 3955 57485 3975
rect 57465 3905 57485 3925
rect 57465 3855 57485 3875
rect 57465 3805 57485 3825
rect 57465 3755 57485 3775
rect 57465 3705 57485 3725
rect 57525 4005 57545 4025
rect 57525 3955 57545 3975
rect 57525 3905 57545 3925
rect 57525 3855 57545 3875
rect 57525 3805 57545 3825
rect 57525 3755 57545 3775
rect 57525 3705 57545 3725
rect 57585 4005 57605 4025
rect 57585 3955 57605 3975
rect 57585 3905 57605 3925
rect 57585 3855 57605 3875
rect 57585 3805 57605 3825
rect 57585 3755 57605 3775
rect 57585 3705 57605 3725
rect 57645 4005 57665 4025
rect 57645 3955 57665 3975
rect 57645 3905 57665 3925
rect 57645 3855 57665 3875
rect 57645 3805 57665 3825
rect 57645 3755 57665 3775
rect 57645 3705 57665 3725
rect 57705 4005 57725 4025
rect 57705 3955 57725 3975
rect 57705 3905 57725 3925
rect 57705 3855 57725 3875
rect 57705 3805 57725 3825
rect 57705 3755 57725 3775
rect 57705 3705 57725 3725
rect 57765 4005 57785 4025
rect 57765 3955 57785 3975
rect 57765 3905 57785 3925
rect 57765 3855 57785 3875
rect 57765 3805 57785 3825
rect 57765 3755 57785 3775
rect 57765 3705 57785 3725
rect 58095 4005 58115 4025
rect 58095 3955 58115 3975
rect 58095 3905 58115 3925
rect 58095 3855 58115 3875
rect 58095 3805 58115 3825
rect 58095 3755 58115 3775
rect 58095 3705 58115 3725
rect 58155 4005 58175 4025
rect 58155 3955 58175 3975
rect 58155 3905 58175 3925
rect 58155 3855 58175 3875
rect 58155 3805 58175 3825
rect 58155 3755 58175 3775
rect 58155 3705 58175 3725
rect 58215 4005 58235 4025
rect 58215 3955 58235 3975
rect 58215 3905 58235 3925
rect 58215 3855 58235 3875
rect 58215 3805 58235 3825
rect 58215 3755 58235 3775
rect 58215 3705 58235 3725
rect 58275 4005 58295 4025
rect 58275 3955 58295 3975
rect 58275 3905 58295 3925
rect 58275 3855 58295 3875
rect 58275 3805 58295 3825
rect 58275 3755 58295 3775
rect 58275 3705 58295 3725
rect 58335 4005 58355 4025
rect 58335 3955 58355 3975
rect 58335 3905 58355 3925
rect 58335 3855 58355 3875
rect 58335 3805 58355 3825
rect 58335 3755 58355 3775
rect 58335 3705 58355 3725
rect 58395 4005 58415 4025
rect 58395 3955 58415 3975
rect 58395 3905 58415 3925
rect 58395 3855 58415 3875
rect 58395 3805 58415 3825
rect 58395 3755 58415 3775
rect 58395 3705 58415 3725
rect 58455 4005 58475 4025
rect 58455 3955 58475 3975
rect 58455 3905 58475 3925
rect 58455 3855 58475 3875
rect 58455 3805 58475 3825
rect 58455 3755 58475 3775
rect 58455 3705 58475 3725
rect 58515 4005 58535 4025
rect 58515 3955 58535 3975
rect 58515 3905 58535 3925
rect 58515 3855 58535 3875
rect 58515 3805 58535 3825
rect 58515 3755 58535 3775
rect 58515 3705 58535 3725
rect 58575 4005 58595 4025
rect 58575 3955 58595 3975
rect 58575 3905 58595 3925
rect 58575 3855 58595 3875
rect 58575 3805 58595 3825
rect 58575 3755 58595 3775
rect 58575 3705 58595 3725
rect 58635 4005 58655 4025
rect 58635 3955 58655 3975
rect 58635 3905 58655 3925
rect 58635 3855 58655 3875
rect 58635 3805 58655 3825
rect 58635 3755 58655 3775
rect 58635 3705 58655 3725
rect 58695 4005 58715 4025
rect 58695 3955 58715 3975
rect 58695 3905 58715 3925
rect 58695 3855 58715 3875
rect 58695 3805 58715 3825
rect 58695 3755 58715 3775
rect 58695 3705 58715 3725
rect 58755 4005 58775 4025
rect 58755 3955 58775 3975
rect 58755 3905 58775 3925
rect 58755 3855 58775 3875
rect 58755 3805 58775 3825
rect 58755 3755 58775 3775
rect 58755 3705 58775 3725
rect 58815 4005 58835 4025
rect 58815 3955 58835 3975
rect 58815 3905 58835 3925
rect 58815 3855 58835 3875
rect 58815 3805 58835 3825
rect 58815 3755 58835 3775
rect 58815 3705 58835 3725
rect 54965 3295 54985 3315
rect 54965 3245 54985 3265
rect 54965 3195 54985 3215
rect 54965 3145 54985 3165
rect 54965 3095 54985 3115
rect 54965 3045 54985 3065
rect 54965 2995 54985 3015
rect 54965 2945 54985 2965
rect 54965 2895 54985 2915
rect 54965 2845 54985 2865
rect 54965 2795 54985 2815
rect 54965 2745 54985 2765
rect 55020 3295 55040 3315
rect 55020 3245 55040 3265
rect 55020 3195 55040 3215
rect 55020 3145 55040 3165
rect 55020 3095 55040 3115
rect 55020 3045 55040 3065
rect 55020 2995 55040 3015
rect 55020 2945 55040 2965
rect 55020 2895 55040 2915
rect 55020 2845 55040 2865
rect 55020 2795 55040 2815
rect 55020 2745 55040 2765
rect 55075 3295 55095 3315
rect 55075 3245 55095 3265
rect 55075 3195 55095 3215
rect 55075 3145 55095 3165
rect 55075 3095 55095 3115
rect 55075 3045 55095 3065
rect 55075 2995 55095 3015
rect 55075 2945 55095 2965
rect 55075 2895 55095 2915
rect 55075 2845 55095 2865
rect 55075 2795 55095 2815
rect 55075 2745 55095 2765
rect 55130 3295 55150 3315
rect 55130 3245 55150 3265
rect 55130 3195 55150 3215
rect 55130 3145 55150 3165
rect 55130 3095 55150 3115
rect 55130 3045 55150 3065
rect 55130 2995 55150 3015
rect 55130 2945 55150 2965
rect 55130 2895 55150 2915
rect 55130 2845 55150 2865
rect 55130 2795 55150 2815
rect 55130 2745 55150 2765
rect 55185 3295 55205 3315
rect 55185 3245 55205 3265
rect 55185 3195 55205 3215
rect 55185 3145 55205 3165
rect 55185 3095 55205 3115
rect 55185 3045 55205 3065
rect 55185 2995 55205 3015
rect 55185 2945 55205 2965
rect 55185 2895 55205 2915
rect 55185 2845 55205 2865
rect 55185 2795 55205 2815
rect 55185 2745 55205 2765
rect 55240 3295 55260 3315
rect 55240 3245 55260 3265
rect 55240 3195 55260 3215
rect 55240 3145 55260 3165
rect 55240 3095 55260 3115
rect 55240 3045 55260 3065
rect 55240 2995 55260 3015
rect 55240 2945 55260 2965
rect 55240 2895 55260 2915
rect 55240 2845 55260 2865
rect 55240 2795 55260 2815
rect 55240 2745 55260 2765
rect 55295 3295 55315 3315
rect 55295 3245 55315 3265
rect 55295 3195 55315 3215
rect 55295 3145 55315 3165
rect 55295 3095 55315 3115
rect 55295 3045 55315 3065
rect 55295 2995 55315 3015
rect 55295 2945 55315 2965
rect 55295 2895 55315 2915
rect 55295 2845 55315 2865
rect 55295 2795 55315 2815
rect 55295 2745 55315 2765
rect 55350 3295 55370 3315
rect 55350 3245 55370 3265
rect 55350 3195 55370 3215
rect 55350 3145 55370 3165
rect 55350 3095 55370 3115
rect 55350 3045 55370 3065
rect 55350 2995 55370 3015
rect 55350 2945 55370 2965
rect 55350 2895 55370 2915
rect 55350 2845 55370 2865
rect 55350 2795 55370 2815
rect 55350 2745 55370 2765
rect 55405 3295 55425 3315
rect 55405 3245 55425 3265
rect 55405 3195 55425 3215
rect 55405 3145 55425 3165
rect 55405 3095 55425 3115
rect 55405 3045 55425 3065
rect 55405 2995 55425 3015
rect 55405 2945 55425 2965
rect 55405 2895 55425 2915
rect 55405 2845 55425 2865
rect 55405 2795 55425 2815
rect 55405 2745 55425 2765
rect 55460 3295 55480 3315
rect 55460 3245 55480 3265
rect 55460 3195 55480 3215
rect 55460 3145 55480 3165
rect 55460 3095 55480 3115
rect 55460 3045 55480 3065
rect 55460 2995 55480 3015
rect 55460 2945 55480 2965
rect 55460 2895 55480 2915
rect 55460 2845 55480 2865
rect 55460 2795 55480 2815
rect 55460 2745 55480 2765
rect 55515 3295 55535 3315
rect 55515 3245 55535 3265
rect 55515 3195 55535 3215
rect 55515 3145 55535 3165
rect 55515 3095 55535 3115
rect 55515 3045 55535 3065
rect 55515 2995 55535 3015
rect 55515 2945 55535 2965
rect 55515 2895 55535 2915
rect 55515 2845 55535 2865
rect 55515 2795 55535 2815
rect 55515 2745 55535 2765
rect 55570 3295 55590 3315
rect 55570 3245 55590 3265
rect 55570 3195 55590 3215
rect 55570 3145 55590 3165
rect 55570 3095 55590 3115
rect 55570 3045 55590 3065
rect 55570 2995 55590 3015
rect 55570 2945 55590 2965
rect 55570 2895 55590 2915
rect 55570 2845 55590 2865
rect 55570 2795 55590 2815
rect 55570 2745 55590 2765
rect 55625 3295 55645 3315
rect 55625 3245 55645 3265
rect 55625 3195 55645 3215
rect 55625 3145 55645 3165
rect 55625 3095 55645 3115
rect 55625 3045 55645 3065
rect 55625 2995 55645 3015
rect 55625 2945 55645 2965
rect 55625 2895 55645 2915
rect 55625 2845 55645 2865
rect 55625 2795 55645 2815
rect 55625 2745 55645 2765
rect 56285 3295 56305 3315
rect 56340 3295 56360 3315
rect 56395 3295 56415 3315
rect 56450 3295 56470 3315
rect 56505 3295 56525 3315
rect 56560 3295 56580 3315
rect 56615 3295 56635 3315
rect 56670 3295 56690 3315
rect 56725 3295 56745 3315
rect 56780 3295 56800 3315
rect 56835 3295 56855 3315
rect 56890 3295 56910 3315
rect 56945 3295 56965 3315
rect 57000 3295 57020 3315
rect 57055 3295 57075 3315
rect 57110 3295 57130 3315
rect 57165 3295 57185 3315
rect 57220 3295 57240 3315
rect 57275 3295 57295 3315
rect 57330 3295 57350 3315
rect 57385 3295 57405 3315
rect 57440 3295 57460 3315
rect 57495 3295 57515 3315
rect 56075 2840 56095 2860
rect 56130 2840 56150 2860
rect 56185 2840 56205 2860
rect 56240 2840 56260 2860
rect 56295 2840 56315 2860
rect 56350 2840 56370 2860
rect 56405 2840 56425 2860
rect 56460 2840 56480 2860
rect 56515 2840 56535 2860
rect 56570 2840 56590 2860
rect 56625 2840 56645 2860
rect 56680 2840 56700 2860
rect 56735 2840 56755 2860
rect 57045 2840 57065 2860
rect 57100 2840 57120 2860
rect 57155 2840 57175 2860
rect 57210 2840 57230 2860
rect 57265 2840 57285 2860
rect 57320 2840 57340 2860
rect 57375 2840 57395 2860
rect 57430 2840 57450 2860
rect 57485 2840 57505 2860
rect 57540 2840 57560 2860
rect 57595 2840 57615 2860
rect 57650 2840 57670 2860
rect 57705 2840 57725 2860
rect 58155 3295 58175 3315
rect 58155 3245 58175 3265
rect 58155 3195 58175 3215
rect 58155 3145 58175 3165
rect 58155 3095 58175 3115
rect 58155 3045 58175 3065
rect 58155 2995 58175 3015
rect 58155 2945 58175 2965
rect 58155 2895 58175 2915
rect 58155 2845 58175 2865
rect 58155 2795 58175 2815
rect 58155 2745 58175 2765
rect 58210 3295 58230 3315
rect 58210 3245 58230 3265
rect 58210 3195 58230 3215
rect 58210 3145 58230 3165
rect 58210 3095 58230 3115
rect 58210 3045 58230 3065
rect 58210 2995 58230 3015
rect 58210 2945 58230 2965
rect 58210 2895 58230 2915
rect 58210 2845 58230 2865
rect 58210 2795 58230 2815
rect 58210 2745 58230 2765
rect 58265 3295 58285 3315
rect 58265 3245 58285 3265
rect 58265 3195 58285 3215
rect 58265 3145 58285 3165
rect 58265 3095 58285 3115
rect 58265 3045 58285 3065
rect 58265 2995 58285 3015
rect 58265 2945 58285 2965
rect 58265 2895 58285 2915
rect 58265 2845 58285 2865
rect 58265 2795 58285 2815
rect 58265 2745 58285 2765
rect 58320 3295 58340 3315
rect 58320 3245 58340 3265
rect 58320 3195 58340 3215
rect 58320 3145 58340 3165
rect 58320 3095 58340 3115
rect 58320 3045 58340 3065
rect 58320 2995 58340 3015
rect 58320 2945 58340 2965
rect 58320 2895 58340 2915
rect 58320 2845 58340 2865
rect 58320 2795 58340 2815
rect 58320 2745 58340 2765
rect 58375 3295 58395 3315
rect 58375 3245 58395 3265
rect 58375 3195 58395 3215
rect 58375 3145 58395 3165
rect 58375 3095 58395 3115
rect 58375 3045 58395 3065
rect 58375 2995 58395 3015
rect 58375 2945 58395 2965
rect 58375 2895 58395 2915
rect 58375 2845 58395 2865
rect 58375 2795 58395 2815
rect 58375 2745 58395 2765
rect 58430 3295 58450 3315
rect 58430 3245 58450 3265
rect 58430 3195 58450 3215
rect 58430 3145 58450 3165
rect 58430 3095 58450 3115
rect 58430 3045 58450 3065
rect 58430 2995 58450 3015
rect 58430 2945 58450 2965
rect 58430 2895 58450 2915
rect 58430 2845 58450 2865
rect 58430 2795 58450 2815
rect 58430 2745 58450 2765
rect 58485 3295 58505 3315
rect 58485 3245 58505 3265
rect 58485 3195 58505 3215
rect 58485 3145 58505 3165
rect 58485 3095 58505 3115
rect 58485 3045 58505 3065
rect 58485 2995 58505 3015
rect 58485 2945 58505 2965
rect 58485 2895 58505 2915
rect 58485 2845 58505 2865
rect 58485 2795 58505 2815
rect 58485 2745 58505 2765
rect 58540 3295 58560 3315
rect 58540 3245 58560 3265
rect 58540 3195 58560 3215
rect 58540 3145 58560 3165
rect 58540 3095 58560 3115
rect 58540 3045 58560 3065
rect 58540 2995 58560 3015
rect 58540 2945 58560 2965
rect 58540 2895 58560 2915
rect 58540 2845 58560 2865
rect 58540 2795 58560 2815
rect 58540 2745 58560 2765
rect 58595 3295 58615 3315
rect 58595 3245 58615 3265
rect 58595 3195 58615 3215
rect 58595 3145 58615 3165
rect 58595 3095 58615 3115
rect 58595 3045 58615 3065
rect 58595 2995 58615 3015
rect 58595 2945 58615 2965
rect 58595 2895 58615 2915
rect 58595 2845 58615 2865
rect 58595 2795 58615 2815
rect 58595 2745 58615 2765
rect 58650 3295 58670 3315
rect 58650 3245 58670 3265
rect 58650 3195 58670 3215
rect 58650 3145 58670 3165
rect 58650 3095 58670 3115
rect 58650 3045 58670 3065
rect 58650 2995 58670 3015
rect 58650 2945 58670 2965
rect 58650 2895 58670 2915
rect 58650 2845 58670 2865
rect 58650 2795 58670 2815
rect 58650 2745 58670 2765
rect 58705 3295 58725 3315
rect 58705 3245 58725 3265
rect 58705 3195 58725 3215
rect 58705 3145 58725 3165
rect 58705 3095 58725 3115
rect 58705 3045 58725 3065
rect 58705 2995 58725 3015
rect 58705 2945 58725 2965
rect 58705 2895 58725 2915
rect 58705 2845 58725 2865
rect 58705 2795 58725 2815
rect 58705 2745 58725 2765
rect 58760 3295 58780 3315
rect 58760 3245 58780 3265
rect 58760 3195 58780 3215
rect 58760 3145 58780 3165
rect 58760 3095 58780 3115
rect 58760 3045 58780 3065
rect 58760 2995 58780 3015
rect 58760 2945 58780 2965
rect 58760 2895 58780 2915
rect 58760 2845 58780 2865
rect 58760 2795 58780 2815
rect 58760 2745 58780 2765
rect 58815 3295 58835 3315
rect 58815 3245 58835 3265
rect 58815 3195 58835 3215
rect 58815 3145 58835 3165
rect 58815 3095 58835 3115
rect 58815 3045 58835 3065
rect 58815 2995 58835 3015
rect 58815 2945 58835 2965
rect 58815 2895 58835 2915
rect 58815 2845 58835 2865
rect 58815 2795 58835 2815
rect 58815 2745 58835 2765
rect 54965 2335 54985 2355
rect 54965 2285 54985 2305
rect 54965 2235 54985 2255
rect 54965 2185 54985 2205
rect 55020 2335 55040 2355
rect 55020 2285 55040 2305
rect 55020 2235 55040 2255
rect 55020 2185 55040 2205
rect 55075 2335 55095 2355
rect 55075 2285 55095 2305
rect 55075 2235 55095 2255
rect 55075 2185 55095 2205
rect 55130 2335 55150 2355
rect 55130 2285 55150 2305
rect 55130 2235 55150 2255
rect 55130 2185 55150 2205
rect 55185 2335 55205 2355
rect 55185 2285 55205 2305
rect 55185 2235 55205 2255
rect 55185 2185 55205 2205
rect 55240 2335 55260 2355
rect 55240 2285 55260 2305
rect 55240 2235 55260 2255
rect 55240 2185 55260 2205
rect 55295 2335 55315 2355
rect 55295 2285 55315 2305
rect 55295 2235 55315 2255
rect 55295 2185 55315 2205
rect 55350 2335 55370 2355
rect 55350 2285 55370 2305
rect 55350 2235 55370 2255
rect 55350 2185 55370 2205
rect 55405 2335 55425 2355
rect 55405 2285 55425 2305
rect 55405 2235 55425 2255
rect 55405 2185 55425 2205
rect 55460 2335 55480 2355
rect 55460 2285 55480 2305
rect 55460 2235 55480 2255
rect 55460 2185 55480 2205
rect 55515 2335 55535 2355
rect 55515 2285 55535 2305
rect 55515 2235 55535 2255
rect 55515 2185 55535 2205
rect 55570 2335 55590 2355
rect 55570 2285 55590 2305
rect 55570 2235 55590 2255
rect 55570 2185 55590 2205
rect 55625 2335 55645 2355
rect 55625 2285 55645 2305
rect 55625 2235 55645 2255
rect 55625 2185 55645 2205
rect 58155 2335 58175 2355
rect 58155 2285 58175 2305
rect 58155 2235 58175 2255
rect 58155 2185 58175 2205
rect 58210 2335 58230 2355
rect 58210 2285 58230 2305
rect 58210 2235 58230 2255
rect 58210 2185 58230 2205
rect 58265 2335 58285 2355
rect 58265 2285 58285 2305
rect 58265 2235 58285 2255
rect 58265 2185 58285 2205
rect 58320 2335 58340 2355
rect 58320 2285 58340 2305
rect 58320 2235 58340 2255
rect 58320 2185 58340 2205
rect 58375 2335 58395 2355
rect 58375 2285 58395 2305
rect 58375 2235 58395 2255
rect 58375 2185 58395 2205
rect 58430 2335 58450 2355
rect 58430 2285 58450 2305
rect 58430 2235 58450 2255
rect 58430 2185 58450 2205
rect 58485 2335 58505 2355
rect 58485 2285 58505 2305
rect 58485 2235 58505 2255
rect 58485 2185 58505 2205
rect 58540 2335 58560 2355
rect 58540 2285 58560 2305
rect 58540 2235 58560 2255
rect 58540 2185 58560 2205
rect 58595 2335 58615 2355
rect 58595 2285 58615 2305
rect 58595 2235 58615 2255
rect 58595 2185 58615 2205
rect 58650 2335 58670 2355
rect 58650 2285 58670 2305
rect 58650 2235 58670 2255
rect 58650 2185 58670 2205
rect 58705 2335 58725 2355
rect 58705 2285 58725 2305
rect 58705 2235 58725 2255
rect 58705 2185 58725 2205
rect 58760 2335 58780 2355
rect 58760 2285 58780 2305
rect 58760 2235 58780 2255
rect 58760 2185 58780 2205
rect 58815 2335 58835 2355
rect 58815 2285 58835 2305
rect 58815 2235 58835 2255
rect 58815 2185 58835 2205
<< psubdiff >>
rect 54485 3345 54765 3365
rect 54485 3040 54505 3345
rect 54485 2660 54505 2945
rect 54745 3040 54765 3345
rect 54745 2660 54765 2945
rect 54485 2640 54585 2660
rect 54665 2640 54765 2660
rect 59035 3345 59315 3365
rect 59035 3040 59055 3345
rect 59035 2660 59055 2945
rect 59295 3040 59315 3345
rect 59295 2660 59315 2945
rect 59035 2640 59135 2660
rect 59215 2640 59315 2660
rect 56500 2535 56860 2555
rect 56940 2535 57300 2555
rect 56500 2465 56520 2535
rect 54400 2280 54535 2300
rect 54615 2280 54755 2300
rect 54400 1945 54420 2280
rect 54400 1535 54420 1865
rect 54735 1945 54755 2280
rect 57280 2465 57300 2535
rect 56500 2335 56520 2385
rect 57280 2335 57300 2385
rect 56500 2315 56860 2335
rect 56940 2315 57300 2335
rect 56025 2255 56825 2275
rect 56025 2145 56045 2255
rect 54735 1535 54755 1865
rect 54400 1515 54535 1535
rect 54615 1515 54755 1535
rect 54905 1985 55265 2005
rect 55345 1985 55705 2005
rect 54905 1800 54925 1985
rect 54905 1535 54925 1720
rect 55685 1800 55705 1985
rect 56025 1955 56045 2065
rect 56805 2145 56825 2255
rect 56805 1955 56825 2065
rect 56025 1935 56825 1955
rect 56975 2255 57775 2275
rect 56975 2145 56995 2255
rect 56975 1955 56995 2065
rect 57755 2145 57775 2255
rect 59235 2300 59275 2320
rect 59045 2280 59185 2300
rect 59265 2280 59400 2300
rect 57755 1955 57775 2065
rect 56975 1935 57775 1955
rect 58095 1985 58455 2005
rect 58535 1985 58895 2005
rect 55685 1535 55705 1720
rect 54905 1515 55265 1535
rect 55345 1515 55705 1535
rect 55980 1785 56860 1805
rect 56940 1785 57820 1805
rect 55980 1675 56000 1785
rect 55980 1485 56000 1595
rect 57800 1675 57820 1785
rect 57800 1485 57820 1595
rect 58095 1800 58115 1985
rect 58095 1535 58115 1720
rect 58875 1800 58895 1985
rect 58875 1535 58895 1720
rect 58095 1515 58455 1535
rect 58535 1515 58895 1535
rect 59045 1945 59065 2280
rect 59045 1535 59065 1865
rect 59380 1945 59400 2280
rect 59380 1535 59400 1865
rect 59045 1515 59185 1535
rect 59265 1515 59400 1535
rect 55980 1465 56860 1485
rect 56940 1465 57820 1485
rect 54985 1395 55315 1415
rect 55395 1395 55725 1415
rect 54660 1340 54735 1360
rect 54815 1340 54895 1360
rect 54660 965 54680 1340
rect 54660 533 54680 885
rect 54875 965 54895 1340
rect 54875 533 54895 885
rect 54660 513 54735 533
rect 54815 513 54895 533
rect 54985 1010 55005 1395
rect 54985 545 55005 930
rect 55705 1010 55725 1395
rect 58075 1395 58405 1415
rect 58485 1395 58815 1415
rect 55705 545 55725 930
rect 56170 1280 56860 1300
rect 56940 1280 57440 1300
rect 57520 1280 57635 1300
rect 56170 1100 56190 1280
rect 56170 875 56190 1020
rect 57615 1100 57635 1280
rect 57615 875 57635 1020
rect 56170 855 56860 875
rect 56940 855 57440 875
rect 57520 855 57635 875
rect 58075 1010 58095 1395
rect 54985 525 55315 545
rect 55395 525 55725 545
rect 56660 765 56865 785
rect 56935 765 57135 785
rect 56660 695 56680 765
rect 57115 695 57135 765
rect 56660 555 56680 615
rect 57115 555 57135 615
rect 56660 535 56865 555
rect 56935 535 57135 555
rect 58075 545 58095 930
rect 58795 1010 58815 1395
rect 58795 545 58815 930
rect 58075 525 58405 545
rect 58485 525 58815 545
rect 58905 1340 58985 1360
rect 59065 1340 59140 1360
rect 58905 965 58925 1340
rect 58905 533 58925 885
rect 59120 965 59140 1340
rect 59120 533 59140 885
rect 58905 513 58985 533
rect 59065 513 59140 533
<< nsubdiff >>
rect 57440 4850 57530 4870
rect 57610 4850 57760 4870
rect 56770 4810 56905 4830
rect 56980 4810 57090 4830
rect 56770 4740 56790 4810
rect 57070 4750 57090 4810
rect 56095 4555 56215 4575
rect 56295 4555 56415 4575
rect 56095 4495 56115 4555
rect 56395 4495 56415 4555
rect 56095 4335 56115 4400
rect 56395 4335 56415 4400
rect 56095 4315 56215 4335
rect 56295 4315 56415 4335
rect 56770 4335 56790 4400
rect 57070 4335 57090 4400
rect 56770 4315 56900 4335
rect 56980 4315 57090 4335
rect 57440 4785 57460 4850
rect 57740 4790 57760 4850
rect 57440 4335 57460 4405
rect 57740 4335 57760 4405
rect 57440 4315 57530 4335
rect 57610 4315 57760 4335
rect 54905 4115 55295 4135
rect 55375 4115 55765 4135
rect 54905 3905 54925 4115
rect 54905 3615 54925 3825
rect 55745 3905 55765 4115
rect 55745 3615 55765 3825
rect 54905 3595 55295 3615
rect 55375 3595 55765 3615
rect 55955 4115 56345 4135
rect 56425 4115 56815 4135
rect 55955 3905 55975 4115
rect 55955 3615 55975 3825
rect 56795 3905 56815 4115
rect 56795 3615 56815 3825
rect 55955 3595 56345 3615
rect 56425 3595 56815 3615
rect 56985 4115 57375 4135
rect 57455 4115 57845 4135
rect 56985 3905 57005 4115
rect 56985 3615 57005 3825
rect 57825 3905 57845 4115
rect 57825 3615 57845 3825
rect 56985 3595 57375 3615
rect 57455 3595 57845 3615
rect 58035 4115 58425 4135
rect 58505 4115 58895 4135
rect 58035 3905 58055 4115
rect 58035 3615 58055 3825
rect 58875 3905 58895 4115
rect 58875 3615 58895 3825
rect 58035 3595 58425 3615
rect 58505 3595 58895 3615
rect 54905 3405 55265 3425
rect 55345 3405 55705 3425
rect 54905 3075 54925 3405
rect 54905 2655 54925 2980
rect 55685 3075 55705 3405
rect 56225 3405 56860 3425
rect 56940 3405 57575 3425
rect 56225 3345 56245 3405
rect 57555 3345 57575 3405
rect 56225 3205 56245 3265
rect 57555 3205 57575 3265
rect 56225 3185 56860 3205
rect 56940 3185 57575 3205
rect 58095 3405 58455 3425
rect 58535 3405 58895 3425
rect 55685 2655 55705 2980
rect 58095 3075 58115 3405
rect 56015 2950 56375 2970
rect 56455 2950 56815 2970
rect 56015 2890 56035 2950
rect 56795 2890 56815 2950
rect 56015 2750 56035 2810
rect 56795 2750 56815 2810
rect 56015 2730 56375 2750
rect 56455 2730 56815 2750
rect 56985 2950 57345 2970
rect 57425 2950 57785 2970
rect 56985 2890 57005 2950
rect 57765 2890 57785 2950
rect 56985 2750 57005 2810
rect 57765 2750 57785 2810
rect 56985 2730 57345 2750
rect 57425 2730 57785 2750
rect 54905 2635 55265 2655
rect 55345 2635 55705 2655
rect 58095 2655 58115 2980
rect 58875 3075 58895 3405
rect 58875 2655 58895 2980
rect 58095 2635 58455 2655
rect 58535 2635 58895 2655
rect 54905 2445 55265 2465
rect 55345 2445 55705 2465
rect 54905 2310 54925 2445
rect 54905 2095 54925 2230
rect 55685 2310 55705 2445
rect 58095 2445 58455 2465
rect 58535 2445 58895 2465
rect 58095 2310 58115 2445
rect 55685 2095 55705 2230
rect 54905 2075 55265 2095
rect 55345 2075 55705 2095
rect 58095 2095 58115 2230
rect 58875 2310 58895 2445
rect 58875 2095 58895 2230
rect 58095 2075 58455 2095
rect 58535 2075 58895 2095
<< psubdiffcont >>
rect 54485 2945 54505 3040
rect 54745 2945 54765 3040
rect 54585 2640 54665 2660
rect 59035 2945 59055 3040
rect 59295 2945 59315 3040
rect 59135 2640 59215 2660
rect 56860 2535 56940 2555
rect 54535 2280 54615 2300
rect 54400 1865 54420 1945
rect 56500 2385 56520 2465
rect 57280 2385 57300 2465
rect 56860 2315 56940 2335
rect 56025 2065 56045 2145
rect 54735 1865 54755 1945
rect 54535 1515 54615 1535
rect 55265 1985 55345 2005
rect 54905 1720 54925 1800
rect 56805 2065 56825 2145
rect 56975 2065 56995 2145
rect 57755 2065 57775 2145
rect 59185 2280 59265 2300
rect 58455 1985 58535 2005
rect 55685 1720 55705 1800
rect 55265 1515 55345 1535
rect 56860 1785 56940 1805
rect 55980 1595 56000 1675
rect 57800 1595 57820 1675
rect 58095 1720 58115 1800
rect 58875 1720 58895 1800
rect 58455 1515 58535 1535
rect 59045 1865 59065 1945
rect 59380 1865 59400 1945
rect 59185 1515 59265 1535
rect 56860 1465 56940 1485
rect 55315 1395 55395 1415
rect 54735 1340 54815 1360
rect 54660 885 54680 965
rect 54875 885 54895 965
rect 54735 513 54815 533
rect 54985 930 55005 1010
rect 58405 1395 58485 1415
rect 55705 930 55725 1010
rect 56860 1280 56940 1300
rect 57440 1280 57520 1300
rect 56170 1020 56190 1100
rect 57615 1020 57635 1100
rect 56860 855 56940 875
rect 57440 855 57520 875
rect 58075 930 58095 1010
rect 55315 525 55395 545
rect 56865 765 56935 785
rect 56660 615 56680 695
rect 57115 615 57135 695
rect 56865 535 56935 555
rect 58795 930 58815 1010
rect 58405 525 58485 545
rect 58985 1340 59065 1360
rect 58905 885 58925 965
rect 59120 885 59140 965
rect 58985 513 59065 533
<< nsubdiffcont >>
rect 57530 4850 57610 4870
rect 56905 4810 56980 4830
rect 56215 4555 56295 4575
rect 56095 4400 56115 4495
rect 56395 4400 56415 4495
rect 56215 4315 56295 4335
rect 56770 4400 56790 4740
rect 57070 4400 57090 4750
rect 56900 4315 56980 4335
rect 57440 4405 57460 4785
rect 57740 4405 57760 4790
rect 57530 4315 57610 4335
rect 55295 4115 55375 4135
rect 54905 3825 54925 3905
rect 55745 3825 55765 3905
rect 55295 3595 55375 3615
rect 56345 4115 56425 4135
rect 55955 3825 55975 3905
rect 56795 3825 56815 3905
rect 56345 3595 56425 3615
rect 57375 4115 57455 4135
rect 56985 3825 57005 3905
rect 57825 3825 57845 3905
rect 57375 3595 57455 3615
rect 58425 4115 58505 4135
rect 58035 3825 58055 3905
rect 58875 3825 58895 3905
rect 58425 3595 58505 3615
rect 55265 3405 55345 3425
rect 54905 2980 54925 3075
rect 56860 3405 56940 3425
rect 56225 3265 56245 3345
rect 57555 3265 57575 3345
rect 56860 3185 56940 3205
rect 58455 3405 58535 3425
rect 55685 2980 55705 3075
rect 58095 2980 58115 3075
rect 56375 2950 56455 2970
rect 56015 2810 56035 2890
rect 56795 2810 56815 2890
rect 56375 2730 56455 2750
rect 57345 2950 57425 2970
rect 56985 2810 57005 2890
rect 57765 2810 57785 2890
rect 57345 2730 57425 2750
rect 55265 2635 55345 2655
rect 58875 2980 58895 3075
rect 58455 2635 58535 2655
rect 55265 2445 55345 2465
rect 54905 2230 54925 2310
rect 58455 2445 58535 2465
rect 55685 2230 55705 2310
rect 55265 2075 55345 2095
rect 58095 2230 58115 2310
rect 58875 2230 58895 2310
rect 58455 2075 58535 2095
<< poly >>
rect 57000 4780 57040 4790
rect 57000 4765 57010 4780
rect 56980 4760 57010 4765
rect 57030 4760 57040 4780
rect 56980 4750 57040 4760
rect 56185 4478 56205 4493
rect 56245 4478 56265 4493
rect 56305 4478 56325 4493
rect 56185 4405 56205 4415
rect 56150 4390 56205 4405
rect 56245 4400 56265 4415
rect 56305 4405 56325 4415
rect 56235 4390 56275 4400
rect 56305 4390 56360 4405
rect 56150 4370 56155 4390
rect 56175 4370 56180 4390
rect 56150 4360 56180 4370
rect 56235 4370 56245 4390
rect 56265 4370 56275 4390
rect 56235 4360 56275 4370
rect 56330 4370 56335 4390
rect 56355 4370 56360 4390
rect 56330 4360 56360 4370
rect 56860 4735 56880 4750
rect 56920 4735 56940 4750
rect 56980 4735 57000 4750
rect 56860 4405 56880 4415
rect 56825 4390 56880 4405
rect 56920 4395 56940 4415
rect 56980 4405 57000 4415
rect 56825 4370 56830 4390
rect 56850 4370 56855 4390
rect 56825 4360 56855 4370
rect 56910 4385 56950 4395
rect 56980 4390 57035 4405
rect 56910 4365 56920 4385
rect 56940 4365 56950 4385
rect 56910 4355 56950 4365
rect 57005 4370 57010 4390
rect 57030 4370 57035 4390
rect 57005 4360 57035 4370
rect 57530 4775 57550 4790
rect 57590 4775 57610 4790
rect 57650 4775 57670 4790
rect 57530 4405 57550 4415
rect 57495 4390 57550 4405
rect 57590 4395 57610 4415
rect 57495 4370 57500 4390
rect 57520 4370 57525 4390
rect 57495 4360 57525 4370
rect 57571 4385 57610 4395
rect 57650 4405 57670 4415
rect 57650 4390 57705 4405
rect 57571 4365 57577 4385
rect 57595 4375 57610 4385
rect 57595 4365 57603 4375
rect 57571 4355 57603 4365
rect 57675 4370 57680 4390
rect 57700 4370 57705 4390
rect 57675 4360 57705 4370
rect 54995 4040 55015 4055
rect 55055 4040 55075 4055
rect 55115 4040 55135 4055
rect 55175 4040 55195 4055
rect 55235 4040 55255 4055
rect 55295 4040 55315 4055
rect 55355 4040 55375 4055
rect 55415 4040 55435 4055
rect 55475 4040 55495 4055
rect 55535 4040 55555 4055
rect 55595 4040 55615 4055
rect 55655 4040 55675 4055
rect 54995 3680 55015 3690
rect 54960 3665 55015 3680
rect 55055 3680 55075 3690
rect 55115 3680 55135 3690
rect 55175 3680 55195 3690
rect 55235 3680 55255 3690
rect 55295 3680 55315 3690
rect 55355 3680 55375 3690
rect 55415 3680 55435 3690
rect 55475 3680 55495 3690
rect 55535 3680 55555 3690
rect 55595 3680 55615 3690
rect 55055 3665 55615 3680
rect 55655 3680 55675 3690
rect 55655 3665 55710 3680
rect 54960 3645 54965 3665
rect 54985 3645 54990 3665
rect 54960 3635 54990 3645
rect 55318 3645 55326 3665
rect 55344 3645 55352 3665
rect 55318 3635 55352 3645
rect 55680 3645 55685 3665
rect 55705 3645 55710 3665
rect 55680 3635 55710 3645
rect 56045 4040 56065 4055
rect 56105 4040 56125 4055
rect 56165 4040 56185 4055
rect 56225 4040 56245 4055
rect 56285 4040 56305 4055
rect 56345 4040 56365 4055
rect 56405 4040 56425 4055
rect 56465 4040 56485 4055
rect 56525 4040 56545 4055
rect 56585 4040 56605 4055
rect 56645 4040 56665 4055
rect 56705 4040 56725 4055
rect 56045 3680 56065 3690
rect 56010 3665 56065 3680
rect 56105 3680 56125 3690
rect 56165 3680 56185 3690
rect 56225 3680 56245 3690
rect 56285 3680 56305 3690
rect 56345 3680 56365 3690
rect 56405 3680 56425 3690
rect 56465 3680 56485 3690
rect 56525 3680 56545 3690
rect 56585 3680 56605 3690
rect 56645 3680 56665 3690
rect 56105 3665 56665 3680
rect 56705 3680 56725 3690
rect 56705 3665 56760 3680
rect 56010 3645 56015 3665
rect 56035 3645 56040 3665
rect 56010 3635 56040 3645
rect 56368 3645 56376 3665
rect 56394 3645 56402 3665
rect 56368 3635 56402 3645
rect 56730 3645 56735 3665
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 57075 4040 57095 4055
rect 57135 4040 57155 4055
rect 57195 4040 57215 4055
rect 57255 4040 57275 4055
rect 57315 4040 57335 4055
rect 57375 4040 57395 4055
rect 57435 4040 57455 4055
rect 57495 4040 57515 4055
rect 57555 4040 57575 4055
rect 57615 4040 57635 4055
rect 57675 4040 57695 4055
rect 57735 4040 57755 4055
rect 57075 3680 57095 3690
rect 57040 3665 57095 3680
rect 57135 3680 57155 3690
rect 57195 3680 57215 3690
rect 57255 3680 57275 3690
rect 57315 3680 57335 3690
rect 57375 3680 57395 3690
rect 57435 3680 57455 3690
rect 57495 3680 57515 3690
rect 57555 3680 57575 3690
rect 57615 3680 57635 3690
rect 57675 3680 57695 3690
rect 57135 3665 57695 3680
rect 57735 3680 57755 3690
rect 57735 3665 57790 3680
rect 57040 3645 57045 3665
rect 57065 3645 57070 3665
rect 57040 3635 57070 3645
rect 57398 3645 57406 3665
rect 57424 3645 57432 3665
rect 57398 3635 57432 3645
rect 57760 3645 57765 3665
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 58125 4040 58145 4055
rect 58185 4040 58205 4055
rect 58245 4040 58265 4055
rect 58305 4040 58325 4055
rect 58365 4040 58385 4055
rect 58425 4040 58445 4055
rect 58485 4040 58505 4055
rect 58545 4040 58565 4055
rect 58605 4040 58625 4055
rect 58665 4040 58685 4055
rect 58725 4040 58745 4055
rect 58785 4040 58805 4055
rect 58125 3680 58145 3690
rect 58090 3665 58145 3680
rect 58185 3680 58205 3690
rect 58245 3680 58265 3690
rect 58305 3680 58325 3690
rect 58365 3680 58385 3690
rect 58425 3680 58445 3690
rect 58485 3680 58505 3690
rect 58545 3680 58565 3690
rect 58605 3680 58625 3690
rect 58665 3680 58685 3690
rect 58725 3680 58745 3690
rect 58185 3665 58745 3680
rect 58785 3680 58805 3690
rect 58785 3665 58840 3680
rect 58090 3645 58095 3665
rect 58115 3645 58120 3665
rect 58090 3635 58120 3645
rect 58448 3645 58456 3665
rect 58474 3645 58482 3665
rect 58448 3635 58482 3645
rect 58810 3645 58815 3665
rect 58835 3645 58840 3665
rect 58810 3635 58840 3645
rect 54995 3330 55010 3345
rect 55050 3330 55065 3345
rect 55105 3330 55120 3345
rect 55160 3330 55175 3345
rect 55215 3330 55230 3345
rect 55270 3330 55285 3345
rect 55325 3330 55340 3345
rect 55380 3330 55395 3345
rect 55435 3330 55450 3345
rect 55490 3330 55505 3345
rect 55545 3330 55560 3345
rect 55600 3330 55615 3345
rect 56315 3330 56330 3345
rect 56370 3330 56385 3345
rect 56425 3330 56440 3345
rect 56480 3330 56495 3345
rect 56535 3330 56550 3345
rect 56590 3330 56605 3345
rect 56645 3330 56660 3345
rect 56700 3330 56715 3345
rect 56755 3330 56770 3345
rect 56810 3330 56825 3345
rect 56865 3330 56880 3345
rect 56920 3330 56935 3345
rect 56975 3330 56990 3345
rect 57030 3330 57045 3345
rect 57085 3330 57100 3345
rect 57140 3330 57155 3345
rect 57195 3330 57210 3345
rect 57250 3330 57265 3345
rect 57305 3330 57320 3345
rect 57360 3330 57375 3345
rect 57415 3330 57430 3345
rect 57470 3330 57485 3345
rect 56315 3270 56330 3280
rect 56280 3255 56330 3270
rect 56370 3270 56385 3280
rect 56425 3270 56440 3280
rect 56480 3270 56495 3280
rect 56535 3270 56550 3280
rect 56590 3270 56605 3280
rect 56645 3270 56660 3280
rect 56700 3270 56715 3280
rect 56755 3270 56770 3280
rect 56810 3270 56825 3280
rect 56865 3270 56880 3280
rect 56920 3270 56935 3280
rect 56975 3270 56990 3280
rect 57030 3270 57045 3280
rect 57085 3270 57100 3280
rect 57140 3270 57155 3280
rect 57195 3270 57210 3280
rect 57250 3270 57265 3280
rect 57305 3270 57320 3280
rect 57360 3270 57375 3280
rect 57415 3270 57430 3280
rect 56370 3255 57430 3270
rect 57470 3270 57485 3280
rect 57470 3255 57520 3270
rect 56280 3235 56285 3255
rect 56305 3235 56310 3255
rect 56280 3225 56310 3235
rect 56497 3235 56505 3255
rect 56525 3235 56533 3255
rect 56497 3225 56533 3235
rect 57490 3235 57495 3255
rect 57515 3235 57520 3255
rect 57490 3225 57520 3235
rect 54995 2720 55010 2730
rect 54960 2705 55010 2720
rect 55050 2720 55065 2730
rect 55105 2720 55120 2730
rect 55160 2720 55175 2730
rect 55215 2720 55230 2730
rect 55270 2720 55285 2730
rect 55325 2720 55340 2730
rect 55380 2720 55395 2730
rect 55435 2720 55450 2730
rect 55490 2720 55505 2730
rect 55545 2720 55560 2730
rect 55050 2705 55560 2720
rect 55600 2720 55615 2730
rect 55600 2705 55650 2720
rect 54960 2685 54965 2705
rect 54985 2685 54990 2705
rect 54960 2675 54990 2685
rect 55178 2685 55186 2705
rect 55204 2685 55212 2705
rect 55178 2675 55212 2685
rect 55620 2685 55625 2705
rect 55645 2685 55650 2705
rect 55620 2675 55650 2685
rect 58185 3330 58200 3345
rect 58240 3330 58255 3345
rect 58295 3330 58310 3345
rect 58350 3330 58365 3345
rect 58405 3330 58420 3345
rect 58460 3330 58475 3345
rect 58515 3330 58530 3345
rect 58570 3330 58585 3345
rect 58625 3330 58640 3345
rect 58680 3330 58695 3345
rect 58735 3330 58750 3345
rect 58790 3330 58805 3345
rect 56145 2920 56175 2930
rect 56145 2900 56150 2920
rect 56170 2900 56175 2920
rect 56345 2920 56375 2930
rect 56345 2900 56350 2920
rect 56370 2900 56375 2920
rect 56560 2920 56600 2930
rect 56560 2900 56570 2920
rect 56590 2900 56600 2920
rect 56145 2890 56175 2900
rect 56105 2875 56120 2890
rect 56160 2875 56175 2890
rect 56215 2875 56230 2890
rect 56270 2875 56285 2890
rect 56325 2885 56395 2900
rect 56325 2875 56340 2885
rect 56380 2875 56395 2885
rect 56435 2875 56450 2890
rect 56490 2875 56505 2890
rect 56545 2885 56615 2900
rect 56545 2875 56560 2885
rect 56600 2875 56615 2885
rect 56655 2875 56670 2890
rect 56710 2875 56725 2890
rect 56105 2815 56120 2825
rect 56070 2800 56120 2815
rect 56160 2810 56175 2825
rect 56215 2815 56230 2825
rect 56270 2815 56285 2825
rect 56215 2810 56285 2815
rect 56325 2810 56340 2825
rect 56380 2810 56395 2825
rect 56435 2815 56450 2825
rect 56490 2815 56505 2825
rect 56435 2810 56505 2815
rect 56545 2810 56560 2825
rect 56600 2810 56615 2825
rect 56655 2810 56670 2825
rect 56215 2800 56304 2810
rect 56435 2800 56524 2810
rect 56070 2780 56075 2800
rect 56095 2780 56100 2800
rect 56070 2770 56100 2780
rect 56272 2780 56278 2800
rect 56295 2780 56304 2800
rect 56272 2770 56304 2780
rect 56492 2780 56498 2800
rect 56515 2780 56524 2800
rect 56492 2770 56524 2780
rect 56636 2800 56670 2810
rect 56710 2815 56725 2825
rect 56710 2800 56760 2815
rect 56636 2780 56645 2800
rect 56662 2780 56670 2800
rect 56636 2770 56670 2780
rect 56730 2780 56735 2800
rect 56755 2780 56760 2800
rect 56730 2770 56760 2780
rect 57113 2920 57143 2930
rect 57113 2900 57118 2920
rect 57138 2900 57143 2920
rect 57310 2920 57350 2930
rect 57310 2900 57320 2920
rect 57340 2900 57350 2920
rect 57530 2920 57570 2930
rect 57530 2900 57540 2920
rect 57560 2900 57570 2920
rect 57113 2890 57145 2900
rect 57075 2875 57090 2890
rect 57130 2875 57145 2890
rect 57185 2875 57200 2890
rect 57240 2875 57255 2890
rect 57295 2885 57365 2900
rect 57295 2875 57310 2885
rect 57350 2875 57365 2885
rect 57405 2875 57420 2890
rect 57460 2875 57475 2890
rect 57515 2885 57585 2900
rect 57515 2875 57530 2885
rect 57570 2875 57585 2885
rect 57625 2875 57640 2890
rect 57680 2875 57695 2890
rect 57075 2815 57090 2825
rect 57040 2800 57090 2815
rect 57130 2810 57145 2825
rect 57185 2815 57200 2825
rect 57240 2815 57255 2825
rect 57185 2810 57255 2815
rect 57295 2810 57310 2825
rect 57350 2810 57365 2825
rect 57405 2815 57420 2825
rect 57460 2815 57475 2825
rect 57405 2810 57475 2815
rect 57515 2810 57530 2825
rect 57570 2810 57585 2825
rect 57625 2810 57640 2825
rect 57185 2800 57274 2810
rect 57405 2800 57494 2810
rect 57040 2780 57045 2800
rect 57065 2780 57070 2800
rect 57040 2770 57070 2780
rect 57242 2780 57248 2800
rect 57265 2780 57274 2800
rect 57242 2770 57274 2780
rect 57462 2780 57468 2800
rect 57485 2780 57494 2800
rect 57462 2770 57494 2780
rect 57606 2800 57640 2810
rect 57680 2815 57695 2825
rect 57680 2800 57730 2815
rect 57606 2780 57615 2800
rect 57632 2780 57640 2800
rect 57606 2770 57640 2780
rect 57700 2780 57705 2800
rect 57725 2780 57730 2800
rect 57700 2770 57730 2780
rect 58185 2720 58200 2730
rect 58150 2705 58200 2720
rect 58240 2720 58255 2730
rect 58295 2720 58310 2730
rect 58350 2720 58365 2730
rect 58405 2720 58420 2730
rect 58460 2720 58475 2730
rect 58515 2720 58530 2730
rect 58570 2720 58585 2730
rect 58625 2720 58640 2730
rect 58680 2720 58695 2730
rect 58735 2720 58750 2730
rect 58240 2705 58750 2720
rect 58790 2720 58805 2730
rect 58790 2705 58840 2720
rect 58150 2685 58155 2705
rect 58175 2685 58180 2705
rect 58150 2675 58180 2685
rect 58588 2685 58596 2705
rect 58614 2685 58622 2705
rect 58588 2675 58622 2685
rect 58810 2685 58815 2705
rect 58835 2685 58840 2705
rect 58810 2675 58840 2685
rect 56555 2505 56585 2515
rect 56555 2485 56560 2505
rect 56580 2485 56585 2505
rect 56715 2505 56755 2515
rect 56715 2485 56725 2505
rect 56745 2485 56755 2505
rect 56935 2505 56975 2515
rect 56935 2485 56945 2505
rect 56965 2485 56975 2505
rect 57215 2505 57245 2515
rect 57215 2485 57220 2505
rect 57240 2485 57245 2505
rect 56555 2470 56605 2485
rect 54995 2370 55010 2385
rect 55050 2370 55065 2385
rect 55105 2370 55120 2385
rect 55160 2370 55175 2385
rect 55215 2370 55230 2385
rect 55270 2370 55285 2385
rect 55325 2370 55340 2385
rect 55380 2370 55395 2385
rect 55435 2370 55450 2385
rect 55490 2370 55505 2385
rect 55545 2370 55560 2385
rect 55600 2370 55615 2385
rect 56590 2460 56605 2470
rect 56645 2470 57155 2485
rect 56645 2460 56660 2470
rect 56700 2460 56715 2470
rect 56755 2460 56770 2470
rect 56810 2460 56825 2470
rect 56865 2460 56880 2470
rect 56920 2460 56935 2470
rect 56975 2460 56990 2470
rect 57030 2460 57045 2470
rect 57085 2460 57100 2470
rect 57140 2460 57155 2470
rect 57195 2470 57245 2485
rect 57195 2460 57210 2470
rect 56590 2395 56605 2410
rect 56645 2395 56660 2410
rect 56700 2395 56715 2410
rect 56755 2395 56770 2410
rect 56810 2395 56825 2410
rect 56865 2395 56880 2410
rect 56920 2395 56935 2410
rect 56975 2395 56990 2410
rect 57030 2395 57045 2410
rect 57085 2395 57100 2410
rect 57140 2395 57155 2410
rect 57195 2395 57210 2410
rect 58185 2370 58200 2385
rect 58240 2370 58255 2385
rect 58295 2370 58310 2385
rect 58350 2370 58365 2385
rect 58405 2370 58420 2385
rect 58460 2370 58475 2385
rect 58515 2370 58530 2385
rect 58570 2370 58585 2385
rect 58625 2370 58640 2385
rect 58680 2370 58695 2385
rect 58735 2370 58750 2385
rect 58790 2370 58805 2385
rect 54995 2160 55010 2170
rect 54960 2145 55010 2160
rect 55050 2160 55065 2170
rect 55105 2160 55120 2170
rect 55160 2160 55175 2170
rect 55215 2160 55230 2170
rect 55270 2160 55285 2170
rect 55325 2160 55340 2170
rect 55380 2160 55395 2170
rect 55435 2160 55450 2170
rect 55490 2160 55505 2170
rect 55545 2160 55560 2170
rect 55050 2145 55560 2160
rect 55600 2160 55615 2170
rect 55600 2145 55650 2160
rect 54960 2125 54965 2145
rect 54985 2125 54990 2145
rect 54960 2115 54990 2125
rect 55453 2125 55461 2145
rect 55479 2125 55487 2145
rect 55453 2115 55487 2125
rect 55620 2125 55625 2145
rect 55645 2125 55650 2145
rect 55620 2115 55650 2125
rect 56080 2225 56110 2235
rect 56080 2205 56085 2225
rect 56105 2205 56110 2225
rect 56410 2225 56440 2235
rect 56410 2205 56415 2225
rect 56435 2205 56440 2225
rect 56740 2225 56770 2235
rect 56740 2205 56745 2225
rect 56765 2205 56770 2225
rect 56080 2190 56130 2205
rect 56115 2180 56130 2190
rect 56170 2190 56680 2205
rect 56170 2180 56185 2190
rect 56225 2180 56240 2190
rect 56280 2180 56295 2190
rect 56335 2180 56350 2190
rect 56390 2180 56405 2190
rect 56445 2180 56460 2190
rect 56500 2180 56515 2190
rect 56555 2180 56570 2190
rect 56610 2180 56625 2190
rect 56665 2180 56680 2190
rect 56720 2190 56770 2205
rect 56720 2180 56735 2190
rect 54960 1955 54990 1965
rect 54960 1935 54965 1955
rect 54985 1935 54990 1955
rect 55453 1955 55487 1965
rect 55453 1935 55461 1955
rect 55479 1935 55487 1955
rect 55620 1955 55650 1965
rect 55620 1935 55625 1955
rect 55645 1935 55650 1955
rect 54960 1920 55010 1935
rect 54995 1910 55010 1920
rect 55050 1920 55560 1935
rect 55050 1910 55065 1920
rect 55105 1910 55120 1920
rect 55160 1910 55175 1920
rect 55215 1910 55230 1920
rect 55270 1910 55285 1920
rect 55325 1910 55340 1920
rect 55380 1910 55395 1920
rect 55435 1910 55450 1920
rect 55490 1910 55505 1920
rect 55545 1910 55560 1920
rect 55600 1920 55650 1935
rect 55600 1910 55615 1920
rect 56115 2015 56130 2030
rect 56170 2015 56185 2030
rect 56225 2015 56240 2030
rect 56280 2015 56295 2030
rect 56335 2015 56350 2030
rect 56390 2015 56405 2030
rect 56445 2015 56460 2030
rect 56500 2015 56515 2030
rect 56555 2015 56570 2030
rect 56610 2015 56625 2030
rect 56665 2015 56680 2030
rect 56720 2015 56735 2030
rect 57030 2225 57060 2235
rect 57030 2205 57035 2225
rect 57055 2205 57060 2225
rect 57360 2225 57390 2235
rect 57360 2205 57365 2225
rect 57385 2205 57390 2225
rect 57690 2225 57720 2235
rect 57690 2205 57695 2225
rect 57715 2205 57720 2225
rect 57030 2190 57080 2205
rect 57065 2180 57080 2190
rect 57120 2190 57630 2205
rect 57120 2180 57135 2190
rect 57175 2180 57190 2190
rect 57230 2180 57245 2190
rect 57285 2180 57300 2190
rect 57340 2180 57355 2190
rect 57395 2180 57410 2190
rect 57450 2180 57465 2190
rect 57505 2180 57520 2190
rect 57560 2180 57575 2190
rect 57615 2180 57630 2190
rect 57670 2190 57720 2205
rect 57670 2180 57685 2190
rect 58185 2160 58200 2170
rect 58150 2145 58200 2160
rect 58240 2160 58255 2170
rect 58295 2160 58310 2170
rect 58350 2160 58365 2170
rect 58405 2160 58420 2170
rect 58460 2160 58475 2170
rect 58515 2160 58530 2170
rect 58570 2160 58585 2170
rect 58625 2160 58640 2170
rect 58680 2160 58695 2170
rect 58735 2160 58750 2170
rect 58240 2145 58750 2160
rect 58790 2160 58805 2170
rect 58790 2145 58840 2160
rect 58150 2125 58155 2145
rect 58175 2125 58180 2145
rect 58150 2115 58180 2125
rect 58313 2125 58321 2145
rect 58339 2125 58347 2145
rect 58313 2115 58347 2125
rect 58810 2125 58815 2145
rect 58835 2125 58840 2145
rect 58810 2115 58840 2125
rect 57065 2015 57080 2030
rect 57120 2015 57135 2030
rect 57175 2015 57190 2030
rect 57230 2015 57245 2030
rect 57285 2015 57300 2030
rect 57340 2015 57355 2030
rect 57395 2015 57410 2030
rect 57450 2015 57465 2030
rect 57505 2015 57520 2030
rect 57560 2015 57575 2030
rect 57615 2015 57630 2030
rect 57670 2015 57685 2030
rect 54995 1595 55010 1610
rect 55050 1595 55065 1610
rect 55105 1595 55120 1610
rect 55160 1595 55175 1610
rect 55215 1595 55230 1610
rect 55270 1595 55285 1610
rect 55325 1595 55340 1610
rect 55380 1595 55395 1610
rect 55435 1595 55450 1610
rect 55490 1595 55505 1610
rect 55545 1595 55560 1610
rect 55600 1595 55615 1610
rect 56035 1755 56065 1765
rect 56035 1735 56040 1755
rect 56060 1735 56065 1755
rect 56237 1755 56269 1765
rect 56237 1735 56243 1755
rect 56260 1735 56269 1755
rect 56457 1755 56489 1765
rect 56457 1735 56463 1755
rect 56480 1735 56489 1755
rect 56035 1720 56085 1735
rect 56180 1725 56269 1735
rect 56400 1725 56489 1735
rect 56601 1755 56635 1765
rect 56601 1735 56610 1755
rect 56627 1735 56635 1755
rect 56695 1755 56725 1765
rect 56695 1735 56700 1755
rect 56720 1735 56725 1755
rect 56601 1725 56635 1735
rect 56070 1710 56085 1720
rect 56125 1710 56140 1725
rect 56180 1720 56250 1725
rect 56180 1710 56195 1720
rect 56235 1710 56250 1720
rect 56290 1710 56305 1725
rect 56345 1710 56360 1725
rect 56400 1720 56470 1725
rect 56400 1710 56415 1720
rect 56455 1710 56470 1720
rect 56510 1710 56525 1725
rect 56565 1710 56580 1725
rect 56620 1710 56635 1725
rect 56675 1720 56725 1735
rect 56775 1755 56805 1765
rect 56775 1735 56780 1755
rect 56800 1735 56805 1755
rect 56867 1755 56899 1765
rect 56867 1740 56873 1755
rect 56865 1735 56873 1740
rect 56890 1735 56899 1755
rect 56995 1755 57025 1765
rect 56995 1735 57000 1755
rect 57020 1735 57025 1755
rect 56775 1720 56825 1735
rect 56675 1710 56690 1720
rect 56810 1710 56825 1720
rect 56865 1725 56899 1735
rect 56865 1710 56880 1725
rect 56920 1710 56935 1725
rect 56975 1720 57025 1735
rect 57075 1755 57105 1765
rect 57075 1735 57080 1755
rect 57100 1735 57105 1755
rect 57277 1755 57309 1765
rect 57277 1735 57283 1755
rect 57300 1735 57309 1755
rect 57497 1755 57529 1765
rect 57497 1735 57503 1755
rect 57520 1735 57529 1755
rect 57075 1720 57125 1735
rect 57220 1725 57309 1735
rect 57440 1725 57529 1735
rect 57641 1755 57675 1765
rect 57641 1735 57650 1755
rect 57667 1735 57675 1755
rect 57735 1755 57765 1765
rect 57735 1735 57740 1755
rect 57760 1735 57765 1755
rect 57641 1725 57675 1735
rect 56975 1710 56990 1720
rect 57110 1710 57125 1720
rect 57165 1710 57180 1725
rect 57220 1720 57290 1725
rect 57220 1710 57235 1720
rect 57275 1710 57290 1720
rect 57330 1710 57345 1725
rect 57385 1710 57400 1725
rect 57440 1720 57510 1725
rect 57440 1710 57455 1720
rect 57495 1710 57510 1720
rect 57550 1710 57565 1725
rect 57605 1710 57620 1725
rect 57660 1710 57675 1725
rect 57715 1720 57765 1735
rect 57715 1710 57730 1720
rect 56070 1545 56085 1560
rect 56125 1545 56140 1560
rect 56180 1545 56195 1560
rect 56235 1545 56250 1560
rect 56290 1550 56305 1560
rect 56345 1550 56360 1560
rect 56106 1535 56140 1545
rect 56290 1535 56360 1550
rect 56400 1545 56415 1560
rect 56455 1545 56470 1560
rect 56510 1550 56525 1560
rect 56565 1550 56580 1560
rect 56510 1535 56580 1550
rect 56620 1545 56635 1560
rect 56675 1545 56690 1560
rect 56810 1545 56825 1560
rect 56865 1545 56880 1560
rect 56920 1545 56935 1560
rect 56975 1545 56990 1560
rect 57110 1545 57125 1560
rect 57165 1545 57180 1560
rect 57220 1545 57235 1560
rect 57275 1545 57290 1560
rect 57330 1550 57345 1560
rect 57385 1550 57400 1560
rect 56920 1535 56954 1545
rect 56106 1515 56112 1535
rect 56129 1515 56138 1535
rect 56106 1505 56138 1515
rect 56305 1515 56315 1535
rect 56335 1515 56345 1535
rect 56305 1505 56345 1515
rect 56525 1515 56535 1535
rect 56555 1515 56565 1535
rect 56525 1505 56565 1515
rect 56922 1515 56928 1535
rect 56945 1515 56954 1535
rect 56922 1505 56954 1515
rect 57146 1535 57180 1545
rect 57330 1535 57400 1550
rect 57440 1545 57455 1560
rect 57495 1545 57510 1560
rect 57550 1550 57565 1560
rect 57605 1550 57620 1560
rect 57550 1535 57620 1550
rect 57660 1545 57675 1560
rect 57715 1545 57730 1560
rect 57146 1515 57152 1535
rect 57169 1515 57178 1535
rect 57146 1505 57178 1515
rect 57345 1515 57355 1535
rect 57375 1515 57385 1535
rect 57345 1505 57385 1515
rect 57565 1515 57575 1535
rect 57595 1515 57605 1535
rect 57565 1505 57605 1515
rect 58150 1955 58180 1965
rect 58150 1935 58155 1955
rect 58175 1935 58180 1955
rect 58313 1955 58347 1965
rect 58313 1935 58321 1955
rect 58339 1935 58347 1955
rect 58810 1955 58840 1965
rect 58810 1935 58815 1955
rect 58835 1935 58840 1955
rect 58150 1920 58200 1935
rect 58185 1910 58200 1920
rect 58240 1920 58750 1935
rect 58240 1910 58255 1920
rect 58295 1910 58310 1920
rect 58350 1910 58365 1920
rect 58405 1910 58420 1920
rect 58460 1910 58475 1920
rect 58515 1910 58530 1920
rect 58570 1910 58585 1920
rect 58625 1910 58640 1920
rect 58680 1910 58695 1920
rect 58735 1910 58750 1920
rect 58790 1920 58840 1935
rect 58790 1910 58805 1920
rect 58185 1595 58200 1610
rect 58240 1595 58255 1610
rect 58295 1595 58310 1610
rect 58350 1595 58365 1610
rect 58405 1595 58420 1610
rect 58460 1595 58475 1610
rect 58515 1595 58530 1610
rect 58570 1595 58585 1610
rect 58625 1595 58640 1610
rect 58680 1595 58695 1610
rect 58735 1595 58750 1610
rect 58790 1595 58805 1610
rect 55040 1365 55070 1375
rect 55040 1345 55045 1365
rect 55065 1345 55070 1365
rect 55438 1365 55472 1375
rect 55438 1345 55446 1365
rect 55464 1345 55472 1365
rect 55640 1365 55670 1375
rect 55640 1345 55645 1365
rect 55665 1345 55670 1365
rect 55040 1330 55135 1345
rect 55075 1320 55135 1330
rect 55175 1330 55535 1345
rect 55175 1320 55235 1330
rect 55275 1320 55335 1330
rect 55375 1320 55435 1330
rect 55475 1320 55535 1330
rect 55575 1330 55670 1345
rect 55575 1320 55635 1330
rect 55075 605 55135 620
rect 55175 605 55235 620
rect 55275 605 55335 620
rect 55375 605 55435 620
rect 55475 605 55535 620
rect 55575 605 55635 620
rect 56830 1250 56860 1260
rect 56830 1230 56835 1250
rect 56855 1230 56860 1250
rect 57470 1250 57504 1260
rect 57470 1230 57479 1250
rect 57499 1230 57504 1250
rect 56260 1205 56275 1220
rect 56315 1215 57375 1230
rect 57470 1220 57504 1230
rect 56315 1205 56330 1215
rect 56370 1205 56385 1215
rect 56425 1205 56440 1215
rect 56480 1205 56495 1215
rect 56535 1205 56550 1215
rect 56590 1205 56605 1215
rect 56645 1205 56660 1215
rect 56700 1205 56715 1215
rect 56755 1205 56770 1215
rect 56810 1205 56825 1215
rect 56865 1205 56880 1215
rect 56920 1205 56935 1215
rect 56975 1205 56990 1215
rect 57030 1205 57045 1215
rect 57085 1205 57100 1215
rect 57140 1205 57155 1215
rect 57195 1205 57210 1215
rect 57250 1205 57265 1215
rect 57305 1205 57320 1215
rect 57360 1205 57375 1215
rect 57415 1205 57430 1220
rect 57470 1205 57485 1220
rect 57525 1205 57540 1220
rect 56260 940 56275 955
rect 56315 940 56330 955
rect 56370 940 56385 955
rect 56425 940 56440 955
rect 56480 940 56495 955
rect 56535 940 56550 955
rect 56590 940 56605 955
rect 56645 940 56660 955
rect 56700 940 56715 955
rect 56755 940 56770 955
rect 56810 940 56825 955
rect 56865 940 56880 955
rect 56920 940 56935 955
rect 56975 940 56990 955
rect 57030 940 57045 955
rect 57085 940 57100 955
rect 57140 940 57155 955
rect 57195 940 57210 955
rect 57250 940 57265 955
rect 57305 940 57320 955
rect 57360 940 57375 955
rect 56210 930 56275 940
rect 56210 910 56220 930
rect 56240 925 56275 930
rect 57415 925 57430 955
rect 57470 940 57485 955
rect 57525 940 57540 955
rect 57525 930 57585 940
rect 57525 925 57555 930
rect 56240 910 56250 925
rect 56210 900 56250 910
rect 57545 910 57555 925
rect 57575 910 57585 930
rect 57545 900 57585 910
rect 58130 1365 58160 1375
rect 58130 1345 58135 1365
rect 58155 1345 58160 1365
rect 58328 1365 58362 1375
rect 58328 1345 58336 1365
rect 58354 1345 58362 1365
rect 58730 1365 58760 1375
rect 58730 1345 58735 1365
rect 58755 1345 58760 1365
rect 58130 1330 58225 1345
rect 58165 1320 58225 1330
rect 58265 1330 58625 1345
rect 58265 1320 58325 1330
rect 58365 1320 58425 1330
rect 58465 1320 58525 1330
rect 58565 1320 58625 1330
rect 58665 1330 58760 1345
rect 58665 1320 58725 1330
rect 56755 735 56795 745
rect 56755 715 56765 735
rect 56785 715 56795 735
rect 56755 705 56795 715
rect 56875 735 56915 745
rect 56875 715 56885 735
rect 56905 715 56915 735
rect 56875 705 56915 715
rect 56995 735 57035 745
rect 56995 715 57005 735
rect 57025 715 57035 735
rect 56995 705 57035 715
rect 56750 690 57040 705
rect 56750 575 57040 590
rect 58165 605 58225 620
rect 58265 605 58325 620
rect 58365 605 58425 620
rect 58465 605 58525 620
rect 58565 605 58625 620
rect 58665 605 58725 620
<< polycont >>
rect 57010 4760 57030 4780
rect 56155 4370 56175 4390
rect 56245 4370 56265 4390
rect 56335 4370 56355 4390
rect 56830 4370 56850 4390
rect 56920 4365 56940 4385
rect 57010 4370 57030 4390
rect 57500 4370 57520 4390
rect 57577 4365 57595 4385
rect 57680 4370 57700 4390
rect 54965 3645 54985 3665
rect 55326 3645 55344 3665
rect 55685 3645 55705 3665
rect 56015 3645 56035 3665
rect 56376 3645 56394 3665
rect 56735 3645 56755 3665
rect 57045 3645 57065 3665
rect 57406 3645 57424 3665
rect 57765 3645 57785 3665
rect 58095 3645 58115 3665
rect 58456 3645 58474 3665
rect 58815 3645 58835 3665
rect 56285 3235 56305 3255
rect 56505 3235 56525 3255
rect 57495 3235 57515 3255
rect 54965 2685 54985 2705
rect 55186 2685 55204 2705
rect 55625 2685 55645 2705
rect 56150 2900 56170 2920
rect 56350 2900 56370 2920
rect 56570 2900 56590 2920
rect 56075 2780 56095 2800
rect 56278 2780 56295 2800
rect 56498 2780 56515 2800
rect 56645 2780 56662 2800
rect 56735 2780 56755 2800
rect 57118 2900 57138 2920
rect 57320 2900 57340 2920
rect 57540 2900 57560 2920
rect 57045 2780 57065 2800
rect 57248 2780 57265 2800
rect 57468 2780 57485 2800
rect 57615 2780 57632 2800
rect 57705 2780 57725 2800
rect 58155 2685 58175 2705
rect 58596 2685 58614 2705
rect 58815 2685 58835 2705
rect 56560 2485 56580 2505
rect 56725 2485 56745 2505
rect 56945 2485 56965 2505
rect 57220 2485 57240 2505
rect 54965 2125 54985 2145
rect 55461 2125 55479 2145
rect 55625 2125 55645 2145
rect 56085 2205 56105 2225
rect 56415 2205 56435 2225
rect 56745 2205 56765 2225
rect 54965 1935 54985 1955
rect 55461 1935 55479 1955
rect 55625 1935 55645 1955
rect 57035 2205 57055 2225
rect 57365 2205 57385 2225
rect 57695 2205 57715 2225
rect 58155 2125 58175 2145
rect 58321 2125 58339 2145
rect 58815 2125 58835 2145
rect 56040 1735 56060 1755
rect 56243 1735 56260 1755
rect 56463 1735 56480 1755
rect 56610 1735 56627 1755
rect 56700 1735 56720 1755
rect 56780 1735 56800 1755
rect 56873 1735 56890 1755
rect 57000 1735 57020 1755
rect 57080 1735 57100 1755
rect 57283 1735 57300 1755
rect 57503 1735 57520 1755
rect 57650 1735 57667 1755
rect 57740 1735 57760 1755
rect 56112 1515 56129 1535
rect 56315 1515 56335 1535
rect 56535 1515 56555 1535
rect 56928 1515 56945 1535
rect 57152 1515 57169 1535
rect 57355 1515 57375 1535
rect 57575 1515 57595 1535
rect 58155 1935 58175 1955
rect 58321 1935 58339 1955
rect 58815 1935 58835 1955
rect 55045 1345 55065 1365
rect 55446 1345 55464 1365
rect 55645 1345 55665 1365
rect 56835 1230 56855 1250
rect 57479 1230 57499 1250
rect 56220 910 56240 930
rect 57555 910 57575 930
rect 58135 1345 58155 1365
rect 58336 1345 58354 1365
rect 58735 1345 58755 1365
rect 56765 715 56785 735
rect 56885 715 56905 735
rect 57005 715 57025 735
<< xpolycontact >>
rect 54554 3065 54695 3285
rect 54554 2720 54695 2940
rect 59105 3065 59246 3285
rect 59105 2720 59246 2940
rect 54470 1989 54505 2209
rect 54470 1600 54505 1820
rect 54530 1989 54565 2209
rect 54530 1600 54565 1820
rect 54590 1989 54625 2209
rect 54590 1600 54625 1820
rect 54650 1989 54685 2209
rect 54650 1600 54685 1820
rect 59115 1979 59150 2199
rect 59115 1600 59150 1820
rect 59175 1979 59210 2199
rect 59175 1600 59210 1820
rect 59235 1979 59270 2199
rect 59235 1600 59270 1820
rect 59295 1979 59330 2199
rect 59295 1600 59330 1820
rect 54730 1050 54765 1270
rect 54730 583 54765 803
rect 54790 1050 54825 1270
rect 54790 583 54825 803
rect 58975 1050 59010 1270
rect 58975 583 59010 803
rect 59035 1050 59070 1270
rect 59035 583 59070 803
<< ppolyres >>
rect 54554 2940 54695 3065
rect 59105 2940 59246 3065
<< xpolyres >>
rect 54470 1820 54505 1989
rect 54530 1820 54565 1989
rect 54590 1820 54625 1989
rect 54650 1820 54685 1989
rect 59115 1820 59150 1979
rect 59175 1820 59210 1979
rect 59235 1820 59270 1979
rect 59295 1820 59330 1979
rect 54730 803 54765 1050
rect 54790 803 54825 1050
rect 58975 803 59010 1050
rect 59035 803 59070 1050
<< locali >>
rect 57440 4850 57530 4870
rect 57610 4850 57760 4870
rect 56770 4810 56905 4830
rect 56980 4810 57090 4830
rect 56770 4740 56790 4810
rect 56820 4780 56860 4790
rect 56820 4760 56830 4780
rect 56850 4760 56860 4780
rect 56820 4750 56860 4760
rect 56887 4780 56913 4790
rect 56887 4760 56890 4780
rect 56910 4760 56913 4780
rect 56887 4750 56913 4760
rect 56940 4780 56980 4790
rect 56940 4760 56950 4780
rect 56970 4760 56980 4780
rect 56940 4750 56980 4760
rect 57000 4780 57040 4790
rect 57000 4760 57010 4780
rect 57030 4760 57040 4780
rect 57000 4750 57040 4760
rect 57070 4750 57090 4810
rect 56095 4555 56215 4575
rect 56295 4555 56415 4575
rect 56095 4495 56115 4555
rect 56145 4525 56185 4535
rect 56145 4505 56155 4525
rect 56175 4505 56185 4525
rect 56145 4495 56185 4505
rect 56205 4525 56245 4535
rect 56205 4505 56215 4525
rect 56235 4505 56245 4525
rect 56205 4495 56245 4505
rect 56325 4525 56365 4535
rect 56325 4505 56335 4525
rect 56355 4505 56365 4525
rect 56325 4495 56365 4505
rect 56395 4495 56415 4555
rect 56155 4473 56175 4495
rect 56215 4473 56235 4495
rect 56335 4473 56355 4495
rect 56095 4335 56115 4400
rect 56150 4450 56180 4473
rect 56150 4430 56155 4450
rect 56175 4430 56180 4450
rect 56150 4390 56180 4430
rect 56210 4450 56240 4473
rect 56210 4430 56215 4450
rect 56235 4430 56240 4450
rect 56210 4420 56240 4430
rect 56270 4450 56300 4473
rect 56270 4430 56275 4450
rect 56295 4430 56300 4450
rect 56270 4420 56300 4430
rect 56330 4450 56360 4473
rect 56330 4430 56335 4450
rect 56355 4430 56360 4450
rect 56275 4400 56295 4420
rect 56150 4370 56155 4390
rect 56175 4370 56180 4390
rect 56150 4360 56180 4370
rect 56235 4390 56295 4400
rect 56235 4370 56245 4390
rect 56265 4380 56295 4390
rect 56330 4390 56360 4430
rect 56265 4370 56275 4380
rect 56235 4360 56275 4370
rect 56330 4370 56335 4390
rect 56355 4370 56360 4390
rect 56330 4360 56360 4370
rect 56155 4335 56175 4360
rect 56335 4335 56355 4360
rect 56395 4335 56415 4400
rect 56095 4315 56215 4335
rect 56295 4315 56415 4335
rect 56830 4730 56850 4750
rect 56890 4730 56910 4750
rect 56950 4730 56970 4750
rect 57010 4730 57030 4750
rect 56770 4335 56790 4400
rect 56825 4705 56855 4730
rect 56825 4435 56830 4705
rect 56850 4435 56855 4705
rect 56825 4390 56855 4435
rect 56885 4705 56915 4730
rect 56885 4435 56890 4705
rect 56910 4435 56915 4705
rect 56885 4420 56915 4435
rect 56945 4705 56975 4730
rect 56945 4435 56950 4705
rect 56970 4435 56975 4705
rect 56945 4420 56975 4435
rect 57005 4705 57035 4730
rect 57005 4435 57010 4705
rect 57030 4435 57035 4705
rect 56825 4370 56830 4390
rect 56850 4370 56855 4390
rect 56825 4360 56855 4370
rect 56910 4385 56950 4395
rect 56910 4365 56920 4385
rect 56940 4365 56950 4385
rect 56830 4335 56850 4360
rect 56910 4355 56950 4365
rect 57005 4390 57035 4435
rect 57005 4370 57010 4390
rect 57030 4370 57035 4390
rect 57005 4360 57035 4370
rect 57010 4335 57030 4360
rect 57070 4335 57090 4400
rect 56770 4315 56900 4335
rect 56980 4315 57090 4335
rect 57440 4785 57460 4850
rect 57490 4820 57530 4830
rect 57490 4800 57500 4820
rect 57520 4800 57530 4820
rect 57490 4790 57530 4800
rect 57550 4820 57590 4830
rect 57550 4800 57560 4820
rect 57580 4800 57590 4820
rect 57550 4790 57590 4800
rect 57670 4820 57710 4830
rect 57670 4800 57680 4820
rect 57700 4800 57710 4820
rect 57670 4790 57710 4800
rect 57740 4790 57760 4850
rect 57500 4770 57520 4790
rect 57560 4770 57580 4790
rect 57680 4770 57700 4790
rect 57440 4335 57460 4405
rect 57495 4745 57525 4770
rect 57495 4435 57500 4745
rect 57520 4435 57525 4745
rect 57495 4390 57525 4435
rect 57555 4745 57585 4770
rect 57555 4435 57560 4745
rect 57580 4435 57585 4745
rect 57555 4420 57585 4435
rect 57615 4745 57645 4770
rect 57615 4435 57620 4745
rect 57640 4435 57645 4745
rect 57615 4420 57645 4435
rect 57675 4745 57705 4770
rect 57675 4435 57680 4745
rect 57700 4435 57705 4745
rect 57620 4400 57640 4420
rect 57495 4370 57500 4390
rect 57520 4370 57525 4390
rect 57495 4360 57525 4370
rect 57571 4385 57603 4395
rect 57571 4365 57577 4385
rect 57595 4365 57603 4385
rect 57500 4335 57520 4360
rect 57571 4355 57603 4365
rect 57620 4390 57650 4400
rect 57620 4370 57625 4390
rect 57645 4370 57650 4390
rect 57620 4360 57650 4370
rect 57675 4390 57705 4435
rect 57675 4370 57680 4390
rect 57700 4370 57705 4390
rect 57675 4360 57705 4370
rect 57680 4335 57700 4360
rect 57740 4335 57760 4405
rect 57440 4315 57530 4335
rect 57610 4315 57760 4335
rect 54905 4115 55295 4135
rect 55375 4115 55765 4135
rect 54905 3905 54925 4115
rect 55325 4095 55345 4115
rect 55075 4085 55115 4095
rect 55075 4065 55085 4085
rect 55105 4065 55115 4085
rect 55075 4055 55115 4065
rect 55195 4085 55235 4095
rect 55195 4065 55205 4085
rect 55225 4065 55235 4085
rect 55195 4055 55235 4065
rect 55315 4085 55355 4095
rect 55315 4065 55325 4085
rect 55345 4065 55355 4085
rect 55315 4055 55355 4065
rect 55435 4085 55475 4095
rect 55435 4065 55445 4085
rect 55465 4065 55475 4085
rect 55435 4055 55475 4065
rect 55555 4085 55595 4095
rect 55555 4065 55565 4085
rect 55585 4065 55595 4085
rect 55555 4055 55595 4065
rect 55085 4035 55105 4055
rect 55205 4035 55225 4055
rect 55325 4035 55345 4055
rect 55445 4035 55465 4055
rect 55565 4035 55585 4055
rect 54905 3615 54925 3825
rect 54960 4025 54990 4035
rect 54960 4005 54965 4025
rect 54985 4005 54990 4025
rect 54960 3975 54990 4005
rect 54960 3955 54965 3975
rect 54985 3955 54990 3975
rect 54960 3925 54990 3955
rect 54960 3905 54965 3925
rect 54985 3905 54990 3925
rect 54960 3875 54990 3905
rect 54960 3855 54965 3875
rect 54985 3855 54990 3875
rect 54960 3825 54990 3855
rect 54960 3805 54965 3825
rect 54985 3805 54990 3825
rect 54960 3775 54990 3805
rect 54960 3755 54965 3775
rect 54985 3755 54990 3775
rect 54960 3725 54990 3755
rect 54960 3705 54965 3725
rect 54985 3705 54990 3725
rect 54960 3665 54990 3705
rect 55020 4025 55050 4035
rect 55020 4005 55025 4025
rect 55045 4005 55050 4025
rect 55020 3975 55050 4005
rect 55020 3955 55025 3975
rect 55045 3955 55050 3975
rect 55020 3925 55050 3955
rect 55020 3905 55025 3925
rect 55045 3905 55050 3925
rect 55020 3875 55050 3905
rect 55020 3855 55025 3875
rect 55045 3855 55050 3875
rect 55020 3825 55050 3855
rect 55020 3805 55025 3825
rect 55045 3805 55050 3825
rect 55020 3775 55050 3805
rect 55020 3755 55025 3775
rect 55045 3755 55050 3775
rect 55020 3725 55050 3755
rect 55020 3705 55025 3725
rect 55045 3705 55050 3725
rect 55020 3695 55050 3705
rect 55080 4025 55110 4035
rect 55080 4005 55085 4025
rect 55105 4005 55110 4025
rect 55080 3975 55110 4005
rect 55080 3955 55085 3975
rect 55105 3955 55110 3975
rect 55080 3925 55110 3955
rect 55080 3905 55085 3925
rect 55105 3905 55110 3925
rect 55080 3875 55110 3905
rect 55080 3855 55085 3875
rect 55105 3855 55110 3875
rect 55080 3825 55110 3855
rect 55080 3805 55085 3825
rect 55105 3805 55110 3825
rect 55080 3775 55110 3805
rect 55080 3755 55085 3775
rect 55105 3755 55110 3775
rect 55080 3725 55110 3755
rect 55080 3705 55085 3725
rect 55105 3705 55110 3725
rect 55080 3695 55110 3705
rect 55140 4025 55170 4035
rect 55140 4005 55145 4025
rect 55165 4005 55170 4025
rect 55140 3975 55170 4005
rect 55140 3955 55145 3975
rect 55165 3955 55170 3975
rect 55140 3925 55170 3955
rect 55140 3905 55145 3925
rect 55165 3905 55170 3925
rect 55140 3875 55170 3905
rect 55140 3855 55145 3875
rect 55165 3855 55170 3875
rect 55140 3825 55170 3855
rect 55140 3805 55145 3825
rect 55165 3805 55170 3825
rect 55140 3775 55170 3805
rect 55140 3755 55145 3775
rect 55165 3755 55170 3775
rect 55140 3725 55170 3755
rect 55140 3705 55145 3725
rect 55165 3705 55170 3725
rect 55140 3695 55170 3705
rect 55200 4025 55230 4035
rect 55200 4005 55205 4025
rect 55225 4005 55230 4025
rect 55200 3975 55230 4005
rect 55200 3955 55205 3975
rect 55225 3955 55230 3975
rect 55200 3925 55230 3955
rect 55200 3905 55205 3925
rect 55225 3905 55230 3925
rect 55200 3875 55230 3905
rect 55200 3855 55205 3875
rect 55225 3855 55230 3875
rect 55200 3825 55230 3855
rect 55200 3805 55205 3825
rect 55225 3805 55230 3825
rect 55200 3775 55230 3805
rect 55200 3755 55205 3775
rect 55225 3755 55230 3775
rect 55200 3725 55230 3755
rect 55200 3705 55205 3725
rect 55225 3705 55230 3725
rect 55200 3695 55230 3705
rect 55260 4025 55290 4035
rect 55260 4005 55265 4025
rect 55285 4005 55290 4025
rect 55260 3975 55290 4005
rect 55260 3955 55265 3975
rect 55285 3955 55290 3975
rect 55260 3925 55290 3955
rect 55260 3905 55265 3925
rect 55285 3905 55290 3925
rect 55260 3875 55290 3905
rect 55260 3855 55265 3875
rect 55285 3855 55290 3875
rect 55260 3825 55290 3855
rect 55260 3805 55265 3825
rect 55285 3805 55290 3825
rect 55260 3775 55290 3805
rect 55260 3755 55265 3775
rect 55285 3755 55290 3775
rect 55260 3725 55290 3755
rect 55260 3705 55265 3725
rect 55285 3705 55290 3725
rect 55260 3695 55290 3705
rect 55320 4025 55350 4035
rect 55320 4005 55325 4025
rect 55345 4005 55350 4025
rect 55320 3975 55350 4005
rect 55320 3955 55325 3975
rect 55345 3955 55350 3975
rect 55320 3925 55350 3955
rect 55320 3905 55325 3925
rect 55345 3905 55350 3925
rect 55320 3875 55350 3905
rect 55320 3855 55325 3875
rect 55345 3855 55350 3875
rect 55320 3825 55350 3855
rect 55320 3805 55325 3825
rect 55345 3805 55350 3825
rect 55320 3775 55350 3805
rect 55320 3755 55325 3775
rect 55345 3755 55350 3775
rect 55320 3725 55350 3755
rect 55320 3705 55325 3725
rect 55345 3705 55350 3725
rect 55320 3695 55350 3705
rect 55380 4025 55410 4035
rect 55380 4005 55385 4025
rect 55405 4005 55410 4025
rect 55380 3975 55410 4005
rect 55380 3955 55385 3975
rect 55405 3955 55410 3975
rect 55380 3925 55410 3955
rect 55380 3905 55385 3925
rect 55405 3905 55410 3925
rect 55380 3875 55410 3905
rect 55380 3855 55385 3875
rect 55405 3855 55410 3875
rect 55380 3825 55410 3855
rect 55380 3805 55385 3825
rect 55405 3805 55410 3825
rect 55380 3775 55410 3805
rect 55380 3755 55385 3775
rect 55405 3755 55410 3775
rect 55380 3725 55410 3755
rect 55380 3705 55385 3725
rect 55405 3705 55410 3725
rect 55380 3695 55410 3705
rect 55440 4025 55470 4035
rect 55440 4005 55445 4025
rect 55465 4005 55470 4025
rect 55440 3975 55470 4005
rect 55440 3955 55445 3975
rect 55465 3955 55470 3975
rect 55440 3925 55470 3955
rect 55440 3905 55445 3925
rect 55465 3905 55470 3925
rect 55440 3875 55470 3905
rect 55440 3855 55445 3875
rect 55465 3855 55470 3875
rect 55440 3825 55470 3855
rect 55440 3805 55445 3825
rect 55465 3805 55470 3825
rect 55440 3775 55470 3805
rect 55440 3755 55445 3775
rect 55465 3755 55470 3775
rect 55440 3725 55470 3755
rect 55440 3705 55445 3725
rect 55465 3705 55470 3725
rect 55440 3695 55470 3705
rect 55500 4025 55530 4035
rect 55500 4005 55505 4025
rect 55525 4005 55530 4025
rect 55500 3975 55530 4005
rect 55500 3955 55505 3975
rect 55525 3955 55530 3975
rect 55500 3925 55530 3955
rect 55500 3905 55505 3925
rect 55525 3905 55530 3925
rect 55500 3875 55530 3905
rect 55500 3855 55505 3875
rect 55525 3855 55530 3875
rect 55500 3825 55530 3855
rect 55500 3805 55505 3825
rect 55525 3805 55530 3825
rect 55500 3775 55530 3805
rect 55500 3755 55505 3775
rect 55525 3755 55530 3775
rect 55500 3725 55530 3755
rect 55500 3705 55505 3725
rect 55525 3705 55530 3725
rect 55500 3695 55530 3705
rect 55560 4025 55590 4035
rect 55560 4005 55565 4025
rect 55585 4005 55590 4025
rect 55560 3975 55590 4005
rect 55560 3955 55565 3975
rect 55585 3955 55590 3975
rect 55560 3925 55590 3955
rect 55560 3905 55565 3925
rect 55585 3905 55590 3925
rect 55560 3875 55590 3905
rect 55560 3855 55565 3875
rect 55585 3855 55590 3875
rect 55560 3825 55590 3855
rect 55560 3805 55565 3825
rect 55585 3805 55590 3825
rect 55560 3775 55590 3805
rect 55560 3755 55565 3775
rect 55585 3755 55590 3775
rect 55560 3725 55590 3755
rect 55560 3705 55565 3725
rect 55585 3705 55590 3725
rect 55560 3695 55590 3705
rect 55620 4025 55650 4035
rect 55620 4005 55625 4025
rect 55645 4005 55650 4025
rect 55620 3975 55650 4005
rect 55620 3955 55625 3975
rect 55645 3955 55650 3975
rect 55620 3925 55650 3955
rect 55620 3905 55625 3925
rect 55645 3905 55650 3925
rect 55620 3875 55650 3905
rect 55620 3855 55625 3875
rect 55645 3855 55650 3875
rect 55620 3825 55650 3855
rect 55620 3805 55625 3825
rect 55645 3805 55650 3825
rect 55620 3775 55650 3805
rect 55620 3755 55625 3775
rect 55645 3755 55650 3775
rect 55620 3725 55650 3755
rect 55620 3705 55625 3725
rect 55645 3705 55650 3725
rect 55620 3695 55650 3705
rect 55680 4025 55710 4035
rect 55680 4005 55685 4025
rect 55705 4005 55710 4025
rect 55680 3975 55710 4005
rect 55680 3955 55685 3975
rect 55705 3955 55710 3975
rect 55680 3925 55710 3955
rect 55680 3905 55685 3925
rect 55705 3905 55710 3925
rect 55680 3875 55710 3905
rect 55680 3855 55685 3875
rect 55705 3855 55710 3875
rect 55680 3825 55710 3855
rect 55680 3805 55685 3825
rect 55705 3805 55710 3825
rect 55680 3775 55710 3805
rect 55680 3755 55685 3775
rect 55705 3755 55710 3775
rect 55680 3725 55710 3755
rect 55680 3705 55685 3725
rect 55705 3705 55710 3725
rect 55025 3675 55045 3695
rect 55145 3675 55165 3695
rect 55265 3675 55285 3695
rect 55385 3675 55405 3695
rect 55505 3675 55525 3695
rect 55625 3675 55645 3695
rect 54960 3645 54965 3665
rect 54985 3645 54990 3665
rect 54960 3635 54990 3645
rect 55015 3665 55055 3675
rect 55015 3645 55025 3665
rect 55045 3645 55055 3665
rect 55015 3635 55055 3645
rect 55135 3665 55175 3675
rect 55135 3645 55145 3665
rect 55165 3645 55175 3665
rect 55135 3635 55175 3645
rect 55255 3665 55295 3675
rect 55255 3645 55265 3665
rect 55285 3645 55295 3665
rect 55255 3635 55295 3645
rect 55318 3665 55352 3675
rect 55318 3645 55326 3665
rect 55344 3645 55352 3665
rect 55318 3635 55352 3645
rect 55375 3665 55415 3675
rect 55375 3645 55385 3665
rect 55405 3645 55415 3665
rect 55375 3635 55415 3645
rect 55495 3665 55535 3675
rect 55495 3645 55505 3665
rect 55525 3645 55535 3665
rect 55495 3635 55535 3645
rect 55615 3665 55655 3675
rect 55615 3645 55625 3665
rect 55645 3645 55655 3665
rect 55615 3635 55655 3645
rect 55680 3665 55710 3705
rect 55680 3645 55685 3665
rect 55705 3645 55710 3665
rect 55680 3635 55710 3645
rect 55745 3905 55765 4115
rect 54965 3615 54985 3635
rect 55685 3615 55705 3635
rect 55745 3615 55765 3825
rect 54905 3595 55295 3615
rect 55375 3595 55765 3615
rect 55955 4115 56345 4135
rect 56425 4115 56815 4135
rect 55955 3905 55975 4115
rect 56125 4085 56165 4095
rect 56125 4065 56135 4085
rect 56155 4065 56165 4085
rect 56125 4055 56165 4065
rect 56245 4085 56285 4095
rect 56245 4065 56255 4085
rect 56275 4065 56285 4085
rect 56245 4055 56285 4065
rect 56365 4085 56405 4095
rect 56365 4065 56375 4085
rect 56395 4065 56405 4085
rect 56365 4055 56405 4065
rect 56485 4085 56525 4095
rect 56485 4065 56495 4085
rect 56515 4065 56525 4085
rect 56485 4055 56525 4065
rect 56605 4085 56645 4095
rect 56605 4065 56615 4085
rect 56635 4065 56645 4085
rect 56605 4055 56645 4065
rect 56135 4035 56155 4055
rect 56255 4035 56275 4055
rect 56375 4035 56395 4055
rect 56495 4035 56515 4055
rect 56615 4035 56635 4055
rect 55955 3615 55975 3825
rect 56010 4025 56040 4035
rect 56010 4005 56015 4025
rect 56035 4005 56040 4025
rect 56010 3975 56040 4005
rect 56010 3955 56015 3975
rect 56035 3955 56040 3975
rect 56010 3925 56040 3955
rect 56010 3905 56015 3925
rect 56035 3905 56040 3925
rect 56010 3875 56040 3905
rect 56010 3855 56015 3875
rect 56035 3855 56040 3875
rect 56010 3825 56040 3855
rect 56010 3805 56015 3825
rect 56035 3805 56040 3825
rect 56010 3775 56040 3805
rect 56010 3755 56015 3775
rect 56035 3755 56040 3775
rect 56010 3725 56040 3755
rect 56010 3705 56015 3725
rect 56035 3705 56040 3725
rect 56010 3665 56040 3705
rect 56070 4025 56100 4035
rect 56070 4005 56075 4025
rect 56095 4005 56100 4025
rect 56070 3975 56100 4005
rect 56070 3955 56075 3975
rect 56095 3955 56100 3975
rect 56070 3925 56100 3955
rect 56070 3905 56075 3925
rect 56095 3905 56100 3925
rect 56070 3875 56100 3905
rect 56070 3855 56075 3875
rect 56095 3855 56100 3875
rect 56070 3825 56100 3855
rect 56070 3805 56075 3825
rect 56095 3805 56100 3825
rect 56070 3775 56100 3805
rect 56070 3755 56075 3775
rect 56095 3755 56100 3775
rect 56070 3725 56100 3755
rect 56070 3705 56075 3725
rect 56095 3705 56100 3725
rect 56070 3695 56100 3705
rect 56130 4025 56160 4035
rect 56130 4005 56135 4025
rect 56155 4005 56160 4025
rect 56130 3975 56160 4005
rect 56130 3955 56135 3975
rect 56155 3955 56160 3975
rect 56130 3925 56160 3955
rect 56130 3905 56135 3925
rect 56155 3905 56160 3925
rect 56130 3875 56160 3905
rect 56130 3855 56135 3875
rect 56155 3855 56160 3875
rect 56130 3825 56160 3855
rect 56130 3805 56135 3825
rect 56155 3805 56160 3825
rect 56130 3775 56160 3805
rect 56130 3755 56135 3775
rect 56155 3755 56160 3775
rect 56130 3725 56160 3755
rect 56130 3705 56135 3725
rect 56155 3705 56160 3725
rect 56130 3695 56160 3705
rect 56190 4025 56220 4035
rect 56190 4005 56195 4025
rect 56215 4005 56220 4025
rect 56190 3975 56220 4005
rect 56190 3955 56195 3975
rect 56215 3955 56220 3975
rect 56190 3925 56220 3955
rect 56190 3905 56195 3925
rect 56215 3905 56220 3925
rect 56190 3875 56220 3905
rect 56190 3855 56195 3875
rect 56215 3855 56220 3875
rect 56190 3825 56220 3855
rect 56190 3805 56195 3825
rect 56215 3805 56220 3825
rect 56190 3775 56220 3805
rect 56190 3755 56195 3775
rect 56215 3755 56220 3775
rect 56190 3725 56220 3755
rect 56190 3705 56195 3725
rect 56215 3705 56220 3725
rect 56190 3695 56220 3705
rect 56250 4025 56280 4035
rect 56250 4005 56255 4025
rect 56275 4005 56280 4025
rect 56250 3975 56280 4005
rect 56250 3955 56255 3975
rect 56275 3955 56280 3975
rect 56250 3925 56280 3955
rect 56250 3905 56255 3925
rect 56275 3905 56280 3925
rect 56250 3875 56280 3905
rect 56250 3855 56255 3875
rect 56275 3855 56280 3875
rect 56250 3825 56280 3855
rect 56250 3805 56255 3825
rect 56275 3805 56280 3825
rect 56250 3775 56280 3805
rect 56250 3755 56255 3775
rect 56275 3755 56280 3775
rect 56250 3725 56280 3755
rect 56250 3705 56255 3725
rect 56275 3705 56280 3725
rect 56250 3695 56280 3705
rect 56310 4025 56340 4035
rect 56310 4005 56315 4025
rect 56335 4005 56340 4025
rect 56310 3975 56340 4005
rect 56310 3955 56315 3975
rect 56335 3955 56340 3975
rect 56310 3925 56340 3955
rect 56310 3905 56315 3925
rect 56335 3905 56340 3925
rect 56310 3875 56340 3905
rect 56310 3855 56315 3875
rect 56335 3855 56340 3875
rect 56310 3825 56340 3855
rect 56310 3805 56315 3825
rect 56335 3805 56340 3825
rect 56310 3775 56340 3805
rect 56310 3755 56315 3775
rect 56335 3755 56340 3775
rect 56310 3725 56340 3755
rect 56310 3705 56315 3725
rect 56335 3705 56340 3725
rect 56310 3695 56340 3705
rect 56370 4025 56400 4035
rect 56370 4005 56375 4025
rect 56395 4005 56400 4025
rect 56370 3975 56400 4005
rect 56370 3955 56375 3975
rect 56395 3955 56400 3975
rect 56370 3925 56400 3955
rect 56370 3905 56375 3925
rect 56395 3905 56400 3925
rect 56370 3875 56400 3905
rect 56370 3855 56375 3875
rect 56395 3855 56400 3875
rect 56370 3825 56400 3855
rect 56370 3805 56375 3825
rect 56395 3805 56400 3825
rect 56370 3775 56400 3805
rect 56370 3755 56375 3775
rect 56395 3755 56400 3775
rect 56370 3725 56400 3755
rect 56370 3705 56375 3725
rect 56395 3705 56400 3725
rect 56370 3695 56400 3705
rect 56430 4025 56460 4035
rect 56430 4005 56435 4025
rect 56455 4005 56460 4025
rect 56430 3975 56460 4005
rect 56430 3955 56435 3975
rect 56455 3955 56460 3975
rect 56430 3925 56460 3955
rect 56430 3905 56435 3925
rect 56455 3905 56460 3925
rect 56430 3875 56460 3905
rect 56430 3855 56435 3875
rect 56455 3855 56460 3875
rect 56430 3825 56460 3855
rect 56430 3805 56435 3825
rect 56455 3805 56460 3825
rect 56430 3775 56460 3805
rect 56430 3755 56435 3775
rect 56455 3755 56460 3775
rect 56430 3725 56460 3755
rect 56430 3705 56435 3725
rect 56455 3705 56460 3725
rect 56430 3695 56460 3705
rect 56490 4025 56520 4035
rect 56490 4005 56495 4025
rect 56515 4005 56520 4025
rect 56490 3975 56520 4005
rect 56490 3955 56495 3975
rect 56515 3955 56520 3975
rect 56490 3925 56520 3955
rect 56490 3905 56495 3925
rect 56515 3905 56520 3925
rect 56490 3875 56520 3905
rect 56490 3855 56495 3875
rect 56515 3855 56520 3875
rect 56490 3825 56520 3855
rect 56490 3805 56495 3825
rect 56515 3805 56520 3825
rect 56490 3775 56520 3805
rect 56490 3755 56495 3775
rect 56515 3755 56520 3775
rect 56490 3725 56520 3755
rect 56490 3705 56495 3725
rect 56515 3705 56520 3725
rect 56490 3695 56520 3705
rect 56550 4025 56580 4035
rect 56550 4005 56555 4025
rect 56575 4005 56580 4025
rect 56550 3975 56580 4005
rect 56550 3955 56555 3975
rect 56575 3955 56580 3975
rect 56550 3925 56580 3955
rect 56550 3905 56555 3925
rect 56575 3905 56580 3925
rect 56550 3875 56580 3905
rect 56550 3855 56555 3875
rect 56575 3855 56580 3875
rect 56550 3825 56580 3855
rect 56550 3805 56555 3825
rect 56575 3805 56580 3825
rect 56550 3775 56580 3805
rect 56550 3755 56555 3775
rect 56575 3755 56580 3775
rect 56550 3725 56580 3755
rect 56550 3705 56555 3725
rect 56575 3705 56580 3725
rect 56550 3695 56580 3705
rect 56610 4025 56640 4035
rect 56610 4005 56615 4025
rect 56635 4005 56640 4025
rect 56610 3975 56640 4005
rect 56610 3955 56615 3975
rect 56635 3955 56640 3975
rect 56610 3925 56640 3955
rect 56610 3905 56615 3925
rect 56635 3905 56640 3925
rect 56610 3875 56640 3905
rect 56610 3855 56615 3875
rect 56635 3855 56640 3875
rect 56610 3825 56640 3855
rect 56610 3805 56615 3825
rect 56635 3805 56640 3825
rect 56610 3775 56640 3805
rect 56610 3755 56615 3775
rect 56635 3755 56640 3775
rect 56610 3725 56640 3755
rect 56610 3705 56615 3725
rect 56635 3705 56640 3725
rect 56610 3695 56640 3705
rect 56670 4025 56700 4035
rect 56670 4005 56675 4025
rect 56695 4005 56700 4025
rect 56670 3975 56700 4005
rect 56670 3955 56675 3975
rect 56695 3955 56700 3975
rect 56670 3925 56700 3955
rect 56670 3905 56675 3925
rect 56695 3905 56700 3925
rect 56670 3875 56700 3905
rect 56670 3855 56675 3875
rect 56695 3855 56700 3875
rect 56670 3825 56700 3855
rect 56670 3805 56675 3825
rect 56695 3805 56700 3825
rect 56670 3775 56700 3805
rect 56670 3755 56675 3775
rect 56695 3755 56700 3775
rect 56670 3725 56700 3755
rect 56670 3705 56675 3725
rect 56695 3705 56700 3725
rect 56670 3695 56700 3705
rect 56730 4025 56760 4035
rect 56730 4005 56735 4025
rect 56755 4005 56760 4025
rect 56730 3975 56760 4005
rect 56730 3955 56735 3975
rect 56755 3955 56760 3975
rect 56730 3925 56760 3955
rect 56730 3905 56735 3925
rect 56755 3905 56760 3925
rect 56730 3875 56760 3905
rect 56730 3855 56735 3875
rect 56755 3855 56760 3875
rect 56730 3825 56760 3855
rect 56730 3805 56735 3825
rect 56755 3805 56760 3825
rect 56730 3775 56760 3805
rect 56730 3755 56735 3775
rect 56755 3755 56760 3775
rect 56730 3725 56760 3755
rect 56730 3705 56735 3725
rect 56755 3705 56760 3725
rect 56075 3675 56095 3695
rect 56195 3675 56215 3695
rect 56315 3675 56335 3695
rect 56435 3675 56455 3695
rect 56555 3675 56575 3695
rect 56675 3675 56695 3695
rect 56010 3645 56015 3665
rect 56035 3645 56040 3665
rect 56010 3635 56040 3645
rect 56065 3665 56105 3675
rect 56065 3645 56075 3665
rect 56095 3645 56105 3665
rect 56065 3635 56105 3645
rect 56185 3665 56225 3675
rect 56185 3645 56195 3665
rect 56215 3645 56225 3665
rect 56185 3635 56225 3645
rect 56305 3665 56345 3675
rect 56305 3645 56315 3665
rect 56335 3645 56345 3665
rect 56305 3635 56345 3645
rect 56368 3665 56402 3675
rect 56368 3645 56376 3665
rect 56394 3645 56402 3665
rect 56368 3635 56402 3645
rect 56425 3665 56465 3675
rect 56425 3645 56435 3665
rect 56455 3645 56465 3665
rect 56425 3635 56465 3645
rect 56545 3665 56585 3675
rect 56545 3645 56555 3665
rect 56575 3645 56585 3665
rect 56545 3635 56585 3645
rect 56665 3665 56705 3675
rect 56665 3645 56675 3665
rect 56695 3645 56705 3665
rect 56665 3635 56705 3645
rect 56730 3665 56760 3705
rect 56730 3645 56735 3665
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 56795 3905 56815 4115
rect 56015 3615 56035 3635
rect 56735 3615 56755 3635
rect 56795 3615 56815 3825
rect 55955 3595 56345 3615
rect 56425 3595 56815 3615
rect 56985 4115 57375 4135
rect 57455 4115 57845 4135
rect 56985 3905 57005 4115
rect 57155 4085 57195 4095
rect 57155 4065 57165 4085
rect 57185 4065 57195 4085
rect 57155 4055 57195 4065
rect 57275 4085 57315 4095
rect 57275 4065 57285 4085
rect 57305 4065 57315 4085
rect 57275 4055 57315 4065
rect 57395 4085 57435 4095
rect 57395 4065 57405 4085
rect 57425 4065 57435 4085
rect 57395 4055 57435 4065
rect 57515 4085 57555 4095
rect 57515 4065 57525 4085
rect 57545 4065 57555 4085
rect 57515 4055 57555 4065
rect 57635 4085 57675 4095
rect 57635 4065 57645 4085
rect 57665 4065 57675 4085
rect 57635 4055 57675 4065
rect 57165 4035 57185 4055
rect 57285 4035 57305 4055
rect 57405 4035 57425 4055
rect 57525 4035 57545 4055
rect 57645 4035 57665 4055
rect 56985 3615 57005 3825
rect 57040 4025 57070 4035
rect 57040 4005 57045 4025
rect 57065 4005 57070 4025
rect 57040 3975 57070 4005
rect 57040 3955 57045 3975
rect 57065 3955 57070 3975
rect 57040 3925 57070 3955
rect 57040 3905 57045 3925
rect 57065 3905 57070 3925
rect 57040 3875 57070 3905
rect 57040 3855 57045 3875
rect 57065 3855 57070 3875
rect 57040 3825 57070 3855
rect 57040 3805 57045 3825
rect 57065 3805 57070 3825
rect 57040 3775 57070 3805
rect 57040 3755 57045 3775
rect 57065 3755 57070 3775
rect 57040 3725 57070 3755
rect 57040 3705 57045 3725
rect 57065 3705 57070 3725
rect 57040 3665 57070 3705
rect 57100 4025 57130 4035
rect 57100 4005 57105 4025
rect 57125 4005 57130 4025
rect 57100 3975 57130 4005
rect 57100 3955 57105 3975
rect 57125 3955 57130 3975
rect 57100 3925 57130 3955
rect 57100 3905 57105 3925
rect 57125 3905 57130 3925
rect 57100 3875 57130 3905
rect 57100 3855 57105 3875
rect 57125 3855 57130 3875
rect 57100 3825 57130 3855
rect 57100 3805 57105 3825
rect 57125 3805 57130 3825
rect 57100 3775 57130 3805
rect 57100 3755 57105 3775
rect 57125 3755 57130 3775
rect 57100 3725 57130 3755
rect 57100 3705 57105 3725
rect 57125 3705 57130 3725
rect 57100 3695 57130 3705
rect 57160 4025 57190 4035
rect 57160 4005 57165 4025
rect 57185 4005 57190 4025
rect 57160 3975 57190 4005
rect 57160 3955 57165 3975
rect 57185 3955 57190 3975
rect 57160 3925 57190 3955
rect 57160 3905 57165 3925
rect 57185 3905 57190 3925
rect 57160 3875 57190 3905
rect 57160 3855 57165 3875
rect 57185 3855 57190 3875
rect 57160 3825 57190 3855
rect 57160 3805 57165 3825
rect 57185 3805 57190 3825
rect 57160 3775 57190 3805
rect 57160 3755 57165 3775
rect 57185 3755 57190 3775
rect 57160 3725 57190 3755
rect 57160 3705 57165 3725
rect 57185 3705 57190 3725
rect 57160 3695 57190 3705
rect 57220 4025 57250 4035
rect 57220 4005 57225 4025
rect 57245 4005 57250 4025
rect 57220 3975 57250 4005
rect 57220 3955 57225 3975
rect 57245 3955 57250 3975
rect 57220 3925 57250 3955
rect 57220 3905 57225 3925
rect 57245 3905 57250 3925
rect 57220 3875 57250 3905
rect 57220 3855 57225 3875
rect 57245 3855 57250 3875
rect 57220 3825 57250 3855
rect 57220 3805 57225 3825
rect 57245 3805 57250 3825
rect 57220 3775 57250 3805
rect 57220 3755 57225 3775
rect 57245 3755 57250 3775
rect 57220 3725 57250 3755
rect 57220 3705 57225 3725
rect 57245 3705 57250 3725
rect 57220 3695 57250 3705
rect 57280 4025 57310 4035
rect 57280 4005 57285 4025
rect 57305 4005 57310 4025
rect 57280 3975 57310 4005
rect 57280 3955 57285 3975
rect 57305 3955 57310 3975
rect 57280 3925 57310 3955
rect 57280 3905 57285 3925
rect 57305 3905 57310 3925
rect 57280 3875 57310 3905
rect 57280 3855 57285 3875
rect 57305 3855 57310 3875
rect 57280 3825 57310 3855
rect 57280 3805 57285 3825
rect 57305 3805 57310 3825
rect 57280 3775 57310 3805
rect 57280 3755 57285 3775
rect 57305 3755 57310 3775
rect 57280 3725 57310 3755
rect 57280 3705 57285 3725
rect 57305 3705 57310 3725
rect 57280 3695 57310 3705
rect 57340 4025 57370 4035
rect 57340 4005 57345 4025
rect 57365 4005 57370 4025
rect 57340 3975 57370 4005
rect 57340 3955 57345 3975
rect 57365 3955 57370 3975
rect 57340 3925 57370 3955
rect 57340 3905 57345 3925
rect 57365 3905 57370 3925
rect 57340 3875 57370 3905
rect 57340 3855 57345 3875
rect 57365 3855 57370 3875
rect 57340 3825 57370 3855
rect 57340 3805 57345 3825
rect 57365 3805 57370 3825
rect 57340 3775 57370 3805
rect 57340 3755 57345 3775
rect 57365 3755 57370 3775
rect 57340 3725 57370 3755
rect 57340 3705 57345 3725
rect 57365 3705 57370 3725
rect 57340 3695 57370 3705
rect 57400 4025 57430 4035
rect 57400 4005 57405 4025
rect 57425 4005 57430 4025
rect 57400 3975 57430 4005
rect 57400 3955 57405 3975
rect 57425 3955 57430 3975
rect 57400 3925 57430 3955
rect 57400 3905 57405 3925
rect 57425 3905 57430 3925
rect 57400 3875 57430 3905
rect 57400 3855 57405 3875
rect 57425 3855 57430 3875
rect 57400 3825 57430 3855
rect 57400 3805 57405 3825
rect 57425 3805 57430 3825
rect 57400 3775 57430 3805
rect 57400 3755 57405 3775
rect 57425 3755 57430 3775
rect 57400 3725 57430 3755
rect 57400 3705 57405 3725
rect 57425 3705 57430 3725
rect 57400 3695 57430 3705
rect 57460 4025 57490 4035
rect 57460 4005 57465 4025
rect 57485 4005 57490 4025
rect 57460 3975 57490 4005
rect 57460 3955 57465 3975
rect 57485 3955 57490 3975
rect 57460 3925 57490 3955
rect 57460 3905 57465 3925
rect 57485 3905 57490 3925
rect 57460 3875 57490 3905
rect 57460 3855 57465 3875
rect 57485 3855 57490 3875
rect 57460 3825 57490 3855
rect 57460 3805 57465 3825
rect 57485 3805 57490 3825
rect 57460 3775 57490 3805
rect 57460 3755 57465 3775
rect 57485 3755 57490 3775
rect 57460 3725 57490 3755
rect 57460 3705 57465 3725
rect 57485 3705 57490 3725
rect 57460 3695 57490 3705
rect 57520 4025 57550 4035
rect 57520 4005 57525 4025
rect 57545 4005 57550 4025
rect 57520 3975 57550 4005
rect 57520 3955 57525 3975
rect 57545 3955 57550 3975
rect 57520 3925 57550 3955
rect 57520 3905 57525 3925
rect 57545 3905 57550 3925
rect 57520 3875 57550 3905
rect 57520 3855 57525 3875
rect 57545 3855 57550 3875
rect 57520 3825 57550 3855
rect 57520 3805 57525 3825
rect 57545 3805 57550 3825
rect 57520 3775 57550 3805
rect 57520 3755 57525 3775
rect 57545 3755 57550 3775
rect 57520 3725 57550 3755
rect 57520 3705 57525 3725
rect 57545 3705 57550 3725
rect 57520 3695 57550 3705
rect 57580 4025 57610 4035
rect 57580 4005 57585 4025
rect 57605 4005 57610 4025
rect 57580 3975 57610 4005
rect 57580 3955 57585 3975
rect 57605 3955 57610 3975
rect 57580 3925 57610 3955
rect 57580 3905 57585 3925
rect 57605 3905 57610 3925
rect 57580 3875 57610 3905
rect 57580 3855 57585 3875
rect 57605 3855 57610 3875
rect 57580 3825 57610 3855
rect 57580 3805 57585 3825
rect 57605 3805 57610 3825
rect 57580 3775 57610 3805
rect 57580 3755 57585 3775
rect 57605 3755 57610 3775
rect 57580 3725 57610 3755
rect 57580 3705 57585 3725
rect 57605 3705 57610 3725
rect 57580 3695 57610 3705
rect 57640 4025 57670 4035
rect 57640 4005 57645 4025
rect 57665 4005 57670 4025
rect 57640 3975 57670 4005
rect 57640 3955 57645 3975
rect 57665 3955 57670 3975
rect 57640 3925 57670 3955
rect 57640 3905 57645 3925
rect 57665 3905 57670 3925
rect 57640 3875 57670 3905
rect 57640 3855 57645 3875
rect 57665 3855 57670 3875
rect 57640 3825 57670 3855
rect 57640 3805 57645 3825
rect 57665 3805 57670 3825
rect 57640 3775 57670 3805
rect 57640 3755 57645 3775
rect 57665 3755 57670 3775
rect 57640 3725 57670 3755
rect 57640 3705 57645 3725
rect 57665 3705 57670 3725
rect 57640 3695 57670 3705
rect 57700 4025 57730 4035
rect 57700 4005 57705 4025
rect 57725 4005 57730 4025
rect 57700 3975 57730 4005
rect 57700 3955 57705 3975
rect 57725 3955 57730 3975
rect 57700 3925 57730 3955
rect 57700 3905 57705 3925
rect 57725 3905 57730 3925
rect 57700 3875 57730 3905
rect 57700 3855 57705 3875
rect 57725 3855 57730 3875
rect 57700 3825 57730 3855
rect 57700 3805 57705 3825
rect 57725 3805 57730 3825
rect 57700 3775 57730 3805
rect 57700 3755 57705 3775
rect 57725 3755 57730 3775
rect 57700 3725 57730 3755
rect 57700 3705 57705 3725
rect 57725 3705 57730 3725
rect 57700 3695 57730 3705
rect 57760 4025 57790 4035
rect 57760 4005 57765 4025
rect 57785 4005 57790 4025
rect 57760 3975 57790 4005
rect 57760 3955 57765 3975
rect 57785 3955 57790 3975
rect 57760 3925 57790 3955
rect 57760 3905 57765 3925
rect 57785 3905 57790 3925
rect 57760 3875 57790 3905
rect 57760 3855 57765 3875
rect 57785 3855 57790 3875
rect 57760 3825 57790 3855
rect 57760 3805 57765 3825
rect 57785 3805 57790 3825
rect 57760 3775 57790 3805
rect 57760 3755 57765 3775
rect 57785 3755 57790 3775
rect 57760 3725 57790 3755
rect 57760 3705 57765 3725
rect 57785 3705 57790 3725
rect 57105 3675 57125 3695
rect 57225 3675 57245 3695
rect 57345 3675 57365 3695
rect 57465 3675 57485 3695
rect 57585 3675 57605 3695
rect 57705 3675 57725 3695
rect 57040 3645 57045 3665
rect 57065 3645 57070 3665
rect 57040 3635 57070 3645
rect 57095 3665 57135 3675
rect 57095 3645 57105 3665
rect 57125 3645 57135 3665
rect 57095 3635 57135 3645
rect 57215 3665 57255 3675
rect 57215 3645 57225 3665
rect 57245 3645 57255 3665
rect 57215 3635 57255 3645
rect 57335 3665 57375 3675
rect 57335 3645 57345 3665
rect 57365 3645 57375 3665
rect 57335 3635 57375 3645
rect 57398 3665 57432 3675
rect 57398 3645 57406 3665
rect 57424 3645 57432 3665
rect 57398 3635 57432 3645
rect 57455 3665 57495 3675
rect 57455 3645 57465 3665
rect 57485 3645 57495 3665
rect 57455 3635 57495 3645
rect 57575 3665 57615 3675
rect 57575 3645 57585 3665
rect 57605 3645 57615 3665
rect 57575 3635 57615 3645
rect 57695 3665 57735 3675
rect 57695 3645 57705 3665
rect 57725 3645 57735 3665
rect 57695 3635 57735 3645
rect 57760 3665 57790 3705
rect 57760 3645 57765 3665
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 57825 3905 57845 4115
rect 57045 3615 57065 3635
rect 57765 3615 57785 3635
rect 57825 3615 57845 3825
rect 56985 3595 57375 3615
rect 57455 3595 57845 3615
rect 58035 4115 58425 4135
rect 58505 4115 58895 4135
rect 58035 3905 58055 4115
rect 58455 4095 58475 4115
rect 58205 4085 58245 4095
rect 58205 4065 58215 4085
rect 58235 4065 58245 4085
rect 58205 4055 58245 4065
rect 58325 4085 58365 4095
rect 58325 4065 58335 4085
rect 58355 4065 58365 4085
rect 58325 4055 58365 4065
rect 58445 4085 58485 4095
rect 58445 4065 58455 4085
rect 58475 4065 58485 4085
rect 58445 4055 58485 4065
rect 58565 4085 58605 4095
rect 58565 4065 58575 4085
rect 58595 4065 58605 4085
rect 58565 4055 58605 4065
rect 58685 4085 58725 4095
rect 58685 4065 58695 4085
rect 58715 4065 58725 4085
rect 58685 4055 58725 4065
rect 58215 4035 58235 4055
rect 58335 4035 58355 4055
rect 58455 4035 58475 4055
rect 58575 4035 58595 4055
rect 58695 4035 58715 4055
rect 58035 3615 58055 3825
rect 58090 4025 58120 4035
rect 58090 4005 58095 4025
rect 58115 4005 58120 4025
rect 58090 3975 58120 4005
rect 58090 3955 58095 3975
rect 58115 3955 58120 3975
rect 58090 3925 58120 3955
rect 58090 3905 58095 3925
rect 58115 3905 58120 3925
rect 58090 3875 58120 3905
rect 58090 3855 58095 3875
rect 58115 3855 58120 3875
rect 58090 3825 58120 3855
rect 58090 3805 58095 3825
rect 58115 3805 58120 3825
rect 58090 3775 58120 3805
rect 58090 3755 58095 3775
rect 58115 3755 58120 3775
rect 58090 3725 58120 3755
rect 58090 3705 58095 3725
rect 58115 3705 58120 3725
rect 58090 3665 58120 3705
rect 58150 4025 58180 4035
rect 58150 4005 58155 4025
rect 58175 4005 58180 4025
rect 58150 3975 58180 4005
rect 58150 3955 58155 3975
rect 58175 3955 58180 3975
rect 58150 3925 58180 3955
rect 58150 3905 58155 3925
rect 58175 3905 58180 3925
rect 58150 3875 58180 3905
rect 58150 3855 58155 3875
rect 58175 3855 58180 3875
rect 58150 3825 58180 3855
rect 58150 3805 58155 3825
rect 58175 3805 58180 3825
rect 58150 3775 58180 3805
rect 58150 3755 58155 3775
rect 58175 3755 58180 3775
rect 58150 3725 58180 3755
rect 58150 3705 58155 3725
rect 58175 3705 58180 3725
rect 58150 3695 58180 3705
rect 58210 4025 58240 4035
rect 58210 4005 58215 4025
rect 58235 4005 58240 4025
rect 58210 3975 58240 4005
rect 58210 3955 58215 3975
rect 58235 3955 58240 3975
rect 58210 3925 58240 3955
rect 58210 3905 58215 3925
rect 58235 3905 58240 3925
rect 58210 3875 58240 3905
rect 58210 3855 58215 3875
rect 58235 3855 58240 3875
rect 58210 3825 58240 3855
rect 58210 3805 58215 3825
rect 58235 3805 58240 3825
rect 58210 3775 58240 3805
rect 58210 3755 58215 3775
rect 58235 3755 58240 3775
rect 58210 3725 58240 3755
rect 58210 3705 58215 3725
rect 58235 3705 58240 3725
rect 58210 3695 58240 3705
rect 58270 4025 58300 4035
rect 58270 4005 58275 4025
rect 58295 4005 58300 4025
rect 58270 3975 58300 4005
rect 58270 3955 58275 3975
rect 58295 3955 58300 3975
rect 58270 3925 58300 3955
rect 58270 3905 58275 3925
rect 58295 3905 58300 3925
rect 58270 3875 58300 3905
rect 58270 3855 58275 3875
rect 58295 3855 58300 3875
rect 58270 3825 58300 3855
rect 58270 3805 58275 3825
rect 58295 3805 58300 3825
rect 58270 3775 58300 3805
rect 58270 3755 58275 3775
rect 58295 3755 58300 3775
rect 58270 3725 58300 3755
rect 58270 3705 58275 3725
rect 58295 3705 58300 3725
rect 58270 3695 58300 3705
rect 58330 4025 58360 4035
rect 58330 4005 58335 4025
rect 58355 4005 58360 4025
rect 58330 3975 58360 4005
rect 58330 3955 58335 3975
rect 58355 3955 58360 3975
rect 58330 3925 58360 3955
rect 58330 3905 58335 3925
rect 58355 3905 58360 3925
rect 58330 3875 58360 3905
rect 58330 3855 58335 3875
rect 58355 3855 58360 3875
rect 58330 3825 58360 3855
rect 58330 3805 58335 3825
rect 58355 3805 58360 3825
rect 58330 3775 58360 3805
rect 58330 3755 58335 3775
rect 58355 3755 58360 3775
rect 58330 3725 58360 3755
rect 58330 3705 58335 3725
rect 58355 3705 58360 3725
rect 58330 3695 58360 3705
rect 58390 4025 58420 4035
rect 58390 4005 58395 4025
rect 58415 4005 58420 4025
rect 58390 3975 58420 4005
rect 58390 3955 58395 3975
rect 58415 3955 58420 3975
rect 58390 3925 58420 3955
rect 58390 3905 58395 3925
rect 58415 3905 58420 3925
rect 58390 3875 58420 3905
rect 58390 3855 58395 3875
rect 58415 3855 58420 3875
rect 58390 3825 58420 3855
rect 58390 3805 58395 3825
rect 58415 3805 58420 3825
rect 58390 3775 58420 3805
rect 58390 3755 58395 3775
rect 58415 3755 58420 3775
rect 58390 3725 58420 3755
rect 58390 3705 58395 3725
rect 58415 3705 58420 3725
rect 58390 3695 58420 3705
rect 58450 4025 58480 4035
rect 58450 4005 58455 4025
rect 58475 4005 58480 4025
rect 58450 3975 58480 4005
rect 58450 3955 58455 3975
rect 58475 3955 58480 3975
rect 58450 3925 58480 3955
rect 58450 3905 58455 3925
rect 58475 3905 58480 3925
rect 58450 3875 58480 3905
rect 58450 3855 58455 3875
rect 58475 3855 58480 3875
rect 58450 3825 58480 3855
rect 58450 3805 58455 3825
rect 58475 3805 58480 3825
rect 58450 3775 58480 3805
rect 58450 3755 58455 3775
rect 58475 3755 58480 3775
rect 58450 3725 58480 3755
rect 58450 3705 58455 3725
rect 58475 3705 58480 3725
rect 58450 3695 58480 3705
rect 58510 4025 58540 4035
rect 58510 4005 58515 4025
rect 58535 4005 58540 4025
rect 58510 3975 58540 4005
rect 58510 3955 58515 3975
rect 58535 3955 58540 3975
rect 58510 3925 58540 3955
rect 58510 3905 58515 3925
rect 58535 3905 58540 3925
rect 58510 3875 58540 3905
rect 58510 3855 58515 3875
rect 58535 3855 58540 3875
rect 58510 3825 58540 3855
rect 58510 3805 58515 3825
rect 58535 3805 58540 3825
rect 58510 3775 58540 3805
rect 58510 3755 58515 3775
rect 58535 3755 58540 3775
rect 58510 3725 58540 3755
rect 58510 3705 58515 3725
rect 58535 3705 58540 3725
rect 58510 3695 58540 3705
rect 58570 4025 58600 4035
rect 58570 4005 58575 4025
rect 58595 4005 58600 4025
rect 58570 3975 58600 4005
rect 58570 3955 58575 3975
rect 58595 3955 58600 3975
rect 58570 3925 58600 3955
rect 58570 3905 58575 3925
rect 58595 3905 58600 3925
rect 58570 3875 58600 3905
rect 58570 3855 58575 3875
rect 58595 3855 58600 3875
rect 58570 3825 58600 3855
rect 58570 3805 58575 3825
rect 58595 3805 58600 3825
rect 58570 3775 58600 3805
rect 58570 3755 58575 3775
rect 58595 3755 58600 3775
rect 58570 3725 58600 3755
rect 58570 3705 58575 3725
rect 58595 3705 58600 3725
rect 58570 3695 58600 3705
rect 58630 4025 58660 4035
rect 58630 4005 58635 4025
rect 58655 4005 58660 4025
rect 58630 3975 58660 4005
rect 58630 3955 58635 3975
rect 58655 3955 58660 3975
rect 58630 3925 58660 3955
rect 58630 3905 58635 3925
rect 58655 3905 58660 3925
rect 58630 3875 58660 3905
rect 58630 3855 58635 3875
rect 58655 3855 58660 3875
rect 58630 3825 58660 3855
rect 58630 3805 58635 3825
rect 58655 3805 58660 3825
rect 58630 3775 58660 3805
rect 58630 3755 58635 3775
rect 58655 3755 58660 3775
rect 58630 3725 58660 3755
rect 58630 3705 58635 3725
rect 58655 3705 58660 3725
rect 58630 3695 58660 3705
rect 58690 4025 58720 4035
rect 58690 4005 58695 4025
rect 58715 4005 58720 4025
rect 58690 3975 58720 4005
rect 58690 3955 58695 3975
rect 58715 3955 58720 3975
rect 58690 3925 58720 3955
rect 58690 3905 58695 3925
rect 58715 3905 58720 3925
rect 58690 3875 58720 3905
rect 58690 3855 58695 3875
rect 58715 3855 58720 3875
rect 58690 3825 58720 3855
rect 58690 3805 58695 3825
rect 58715 3805 58720 3825
rect 58690 3775 58720 3805
rect 58690 3755 58695 3775
rect 58715 3755 58720 3775
rect 58690 3725 58720 3755
rect 58690 3705 58695 3725
rect 58715 3705 58720 3725
rect 58690 3695 58720 3705
rect 58750 4025 58780 4035
rect 58750 4005 58755 4025
rect 58775 4005 58780 4025
rect 58750 3975 58780 4005
rect 58750 3955 58755 3975
rect 58775 3955 58780 3975
rect 58750 3925 58780 3955
rect 58750 3905 58755 3925
rect 58775 3905 58780 3925
rect 58750 3875 58780 3905
rect 58750 3855 58755 3875
rect 58775 3855 58780 3875
rect 58750 3825 58780 3855
rect 58750 3805 58755 3825
rect 58775 3805 58780 3825
rect 58750 3775 58780 3805
rect 58750 3755 58755 3775
rect 58775 3755 58780 3775
rect 58750 3725 58780 3755
rect 58750 3705 58755 3725
rect 58775 3705 58780 3725
rect 58750 3695 58780 3705
rect 58810 4025 58840 4035
rect 58810 4005 58815 4025
rect 58835 4005 58840 4025
rect 58810 3975 58840 4005
rect 58810 3955 58815 3975
rect 58835 3955 58840 3975
rect 58810 3925 58840 3955
rect 58810 3905 58815 3925
rect 58835 3905 58840 3925
rect 58810 3875 58840 3905
rect 58810 3855 58815 3875
rect 58835 3855 58840 3875
rect 58810 3825 58840 3855
rect 58810 3805 58815 3825
rect 58835 3805 58840 3825
rect 58810 3775 58840 3805
rect 58810 3755 58815 3775
rect 58835 3755 58840 3775
rect 58810 3725 58840 3755
rect 58810 3705 58815 3725
rect 58835 3705 58840 3725
rect 58155 3675 58175 3695
rect 58275 3675 58295 3695
rect 58395 3675 58415 3695
rect 58515 3675 58535 3695
rect 58635 3675 58655 3695
rect 58755 3675 58775 3695
rect 58090 3645 58095 3665
rect 58115 3645 58120 3665
rect 58090 3635 58120 3645
rect 58145 3665 58185 3675
rect 58145 3645 58155 3665
rect 58175 3645 58185 3665
rect 58145 3635 58185 3645
rect 58265 3665 58305 3675
rect 58265 3645 58275 3665
rect 58295 3645 58305 3665
rect 58265 3635 58305 3645
rect 58385 3665 58425 3675
rect 58385 3645 58395 3665
rect 58415 3645 58425 3665
rect 58385 3635 58425 3645
rect 58448 3665 58482 3675
rect 58448 3645 58456 3665
rect 58474 3645 58482 3665
rect 58448 3635 58482 3645
rect 58505 3665 58545 3675
rect 58505 3645 58515 3665
rect 58535 3645 58545 3665
rect 58505 3635 58545 3645
rect 58625 3665 58665 3675
rect 58625 3645 58635 3665
rect 58655 3645 58665 3665
rect 58625 3635 58665 3645
rect 58745 3665 58785 3675
rect 58745 3645 58755 3665
rect 58775 3645 58785 3665
rect 58745 3635 58785 3645
rect 58810 3665 58840 3705
rect 58810 3645 58815 3665
rect 58835 3645 58840 3665
rect 58810 3635 58840 3645
rect 58875 3905 58895 4115
rect 58095 3615 58115 3635
rect 58815 3615 58835 3635
rect 58875 3615 58895 3825
rect 58035 3595 58425 3615
rect 58505 3595 58895 3615
rect 54905 3405 55265 3425
rect 55345 3405 55705 3425
rect 54485 3345 54765 3365
rect 54485 3040 54505 3345
rect 54554 3320 54695 3325
rect 54554 3290 54560 3320
rect 54590 3290 54610 3320
rect 54640 3290 54659 3320
rect 54689 3290 54695 3320
rect 54554 3285 54695 3290
rect 54485 2660 54505 2945
rect 54745 3040 54765 3345
rect 54554 2715 54695 2720
rect 54554 2685 54560 2715
rect 54590 2685 54610 2715
rect 54640 2685 54659 2715
rect 54689 2685 54695 2715
rect 54554 2680 54695 2685
rect 54745 2660 54765 2945
rect 54485 2650 54585 2660
rect 54485 2640 54535 2650
rect 54525 2630 54535 2640
rect 54555 2640 54585 2650
rect 54665 2640 54765 2660
rect 54905 3075 54925 3405
rect 54955 3375 54995 3385
rect 54955 3355 54965 3375
rect 54985 3355 54995 3375
rect 54955 3345 54995 3355
rect 55065 3375 55105 3385
rect 55065 3355 55075 3375
rect 55095 3355 55105 3375
rect 55065 3345 55105 3355
rect 55175 3375 55215 3385
rect 55175 3355 55185 3375
rect 55205 3355 55215 3375
rect 55175 3345 55215 3355
rect 55285 3375 55325 3385
rect 55285 3355 55295 3375
rect 55315 3355 55325 3375
rect 55285 3345 55325 3355
rect 55395 3375 55435 3385
rect 55395 3355 55405 3375
rect 55425 3355 55435 3375
rect 55395 3345 55435 3355
rect 55505 3375 55545 3385
rect 55505 3355 55515 3375
rect 55535 3355 55545 3375
rect 55505 3345 55545 3355
rect 55615 3375 55655 3385
rect 55615 3355 55625 3375
rect 55645 3355 55655 3375
rect 55615 3345 55655 3355
rect 54965 3325 54985 3345
rect 55075 3325 55095 3345
rect 55185 3325 55205 3345
rect 55295 3325 55315 3345
rect 55405 3325 55425 3345
rect 55515 3325 55535 3345
rect 55625 3325 55645 3345
rect 54905 2655 54925 2980
rect 54960 3315 54990 3325
rect 54960 3295 54965 3315
rect 54985 3295 54990 3315
rect 54960 3265 54990 3295
rect 54960 3245 54965 3265
rect 54985 3245 54990 3265
rect 54960 3215 54990 3245
rect 54960 3195 54965 3215
rect 54985 3195 54990 3215
rect 54960 3165 54990 3195
rect 54960 3145 54965 3165
rect 54985 3145 54990 3165
rect 54960 3115 54990 3145
rect 54960 3095 54965 3115
rect 54985 3095 54990 3115
rect 54960 3065 54990 3095
rect 54960 3045 54965 3065
rect 54985 3045 54990 3065
rect 54960 3015 54990 3045
rect 54960 2995 54965 3015
rect 54985 2995 54990 3015
rect 54960 2965 54990 2995
rect 54960 2945 54965 2965
rect 54985 2945 54990 2965
rect 54960 2915 54990 2945
rect 54960 2895 54965 2915
rect 54985 2895 54990 2915
rect 54960 2865 54990 2895
rect 54960 2845 54965 2865
rect 54985 2845 54990 2865
rect 54960 2815 54990 2845
rect 54960 2795 54965 2815
rect 54985 2795 54990 2815
rect 54960 2765 54990 2795
rect 54960 2745 54965 2765
rect 54985 2745 54990 2765
rect 54960 2705 54990 2745
rect 55015 3315 55045 3325
rect 55015 3295 55020 3315
rect 55040 3295 55045 3315
rect 55015 3265 55045 3295
rect 55015 3245 55020 3265
rect 55040 3245 55045 3265
rect 55015 3215 55045 3245
rect 55015 3195 55020 3215
rect 55040 3195 55045 3215
rect 55015 3165 55045 3195
rect 55015 3145 55020 3165
rect 55040 3145 55045 3165
rect 55015 3115 55045 3145
rect 55015 3095 55020 3115
rect 55040 3095 55045 3115
rect 55015 3065 55045 3095
rect 55015 3045 55020 3065
rect 55040 3045 55045 3065
rect 55015 3015 55045 3045
rect 55015 2995 55020 3015
rect 55040 2995 55045 3015
rect 55015 2965 55045 2995
rect 55015 2945 55020 2965
rect 55040 2945 55045 2965
rect 55015 2915 55045 2945
rect 55015 2895 55020 2915
rect 55040 2895 55045 2915
rect 55015 2865 55045 2895
rect 55015 2845 55020 2865
rect 55040 2845 55045 2865
rect 55015 2815 55045 2845
rect 55015 2795 55020 2815
rect 55040 2795 55045 2815
rect 55015 2765 55045 2795
rect 55015 2745 55020 2765
rect 55040 2745 55045 2765
rect 55015 2735 55045 2745
rect 55070 3315 55100 3325
rect 55070 3295 55075 3315
rect 55095 3295 55100 3315
rect 55070 3265 55100 3295
rect 55070 3245 55075 3265
rect 55095 3245 55100 3265
rect 55070 3215 55100 3245
rect 55070 3195 55075 3215
rect 55095 3195 55100 3215
rect 55070 3165 55100 3195
rect 55070 3145 55075 3165
rect 55095 3145 55100 3165
rect 55070 3115 55100 3145
rect 55070 3095 55075 3115
rect 55095 3095 55100 3115
rect 55070 3065 55100 3095
rect 55070 3045 55075 3065
rect 55095 3045 55100 3065
rect 55070 3015 55100 3045
rect 55070 2995 55075 3015
rect 55095 2995 55100 3015
rect 55070 2965 55100 2995
rect 55070 2945 55075 2965
rect 55095 2945 55100 2965
rect 55070 2915 55100 2945
rect 55070 2895 55075 2915
rect 55095 2895 55100 2915
rect 55070 2865 55100 2895
rect 55070 2845 55075 2865
rect 55095 2845 55100 2865
rect 55070 2815 55100 2845
rect 55070 2795 55075 2815
rect 55095 2795 55100 2815
rect 55070 2765 55100 2795
rect 55070 2745 55075 2765
rect 55095 2745 55100 2765
rect 55070 2735 55100 2745
rect 55125 3315 55155 3325
rect 55125 3295 55130 3315
rect 55150 3295 55155 3315
rect 55125 3265 55155 3295
rect 55125 3245 55130 3265
rect 55150 3245 55155 3265
rect 55125 3215 55155 3245
rect 55125 3195 55130 3215
rect 55150 3195 55155 3215
rect 55125 3165 55155 3195
rect 55125 3145 55130 3165
rect 55150 3145 55155 3165
rect 55125 3115 55155 3145
rect 55125 3095 55130 3115
rect 55150 3095 55155 3115
rect 55125 3065 55155 3095
rect 55125 3045 55130 3065
rect 55150 3045 55155 3065
rect 55125 3015 55155 3045
rect 55125 2995 55130 3015
rect 55150 2995 55155 3015
rect 55125 2965 55155 2995
rect 55125 2945 55130 2965
rect 55150 2945 55155 2965
rect 55125 2915 55155 2945
rect 55125 2895 55130 2915
rect 55150 2895 55155 2915
rect 55125 2865 55155 2895
rect 55125 2845 55130 2865
rect 55150 2845 55155 2865
rect 55125 2815 55155 2845
rect 55125 2795 55130 2815
rect 55150 2795 55155 2815
rect 55125 2765 55155 2795
rect 55125 2745 55130 2765
rect 55150 2745 55155 2765
rect 55125 2735 55155 2745
rect 55180 3315 55210 3325
rect 55180 3295 55185 3315
rect 55205 3295 55210 3315
rect 55180 3265 55210 3295
rect 55180 3245 55185 3265
rect 55205 3245 55210 3265
rect 55180 3215 55210 3245
rect 55180 3195 55185 3215
rect 55205 3195 55210 3215
rect 55180 3165 55210 3195
rect 55180 3145 55185 3165
rect 55205 3145 55210 3165
rect 55180 3115 55210 3145
rect 55180 3095 55185 3115
rect 55205 3095 55210 3115
rect 55180 3065 55210 3095
rect 55180 3045 55185 3065
rect 55205 3045 55210 3065
rect 55180 3015 55210 3045
rect 55180 2995 55185 3015
rect 55205 2995 55210 3015
rect 55180 2965 55210 2995
rect 55180 2945 55185 2965
rect 55205 2945 55210 2965
rect 55180 2915 55210 2945
rect 55180 2895 55185 2915
rect 55205 2895 55210 2915
rect 55180 2865 55210 2895
rect 55180 2845 55185 2865
rect 55205 2845 55210 2865
rect 55180 2815 55210 2845
rect 55180 2795 55185 2815
rect 55205 2795 55210 2815
rect 55180 2765 55210 2795
rect 55180 2745 55185 2765
rect 55205 2745 55210 2765
rect 55180 2735 55210 2745
rect 55235 3315 55265 3325
rect 55235 3295 55240 3315
rect 55260 3295 55265 3315
rect 55235 3265 55265 3295
rect 55235 3245 55240 3265
rect 55260 3245 55265 3265
rect 55235 3215 55265 3245
rect 55235 3195 55240 3215
rect 55260 3195 55265 3215
rect 55235 3165 55265 3195
rect 55235 3145 55240 3165
rect 55260 3145 55265 3165
rect 55235 3115 55265 3145
rect 55235 3095 55240 3115
rect 55260 3095 55265 3115
rect 55235 3065 55265 3095
rect 55235 3045 55240 3065
rect 55260 3045 55265 3065
rect 55235 3015 55265 3045
rect 55235 2995 55240 3015
rect 55260 2995 55265 3015
rect 55235 2965 55265 2995
rect 55235 2945 55240 2965
rect 55260 2945 55265 2965
rect 55235 2915 55265 2945
rect 55235 2895 55240 2915
rect 55260 2895 55265 2915
rect 55235 2865 55265 2895
rect 55235 2845 55240 2865
rect 55260 2845 55265 2865
rect 55235 2815 55265 2845
rect 55235 2795 55240 2815
rect 55260 2795 55265 2815
rect 55235 2765 55265 2795
rect 55235 2745 55240 2765
rect 55260 2745 55265 2765
rect 55235 2735 55265 2745
rect 55290 3315 55320 3325
rect 55290 3295 55295 3315
rect 55315 3295 55320 3315
rect 55290 3265 55320 3295
rect 55290 3245 55295 3265
rect 55315 3245 55320 3265
rect 55290 3215 55320 3245
rect 55290 3195 55295 3215
rect 55315 3195 55320 3215
rect 55290 3165 55320 3195
rect 55290 3145 55295 3165
rect 55315 3145 55320 3165
rect 55290 3115 55320 3145
rect 55290 3095 55295 3115
rect 55315 3095 55320 3115
rect 55290 3065 55320 3095
rect 55290 3045 55295 3065
rect 55315 3045 55320 3065
rect 55290 3015 55320 3045
rect 55290 2995 55295 3015
rect 55315 2995 55320 3015
rect 55290 2965 55320 2995
rect 55290 2945 55295 2965
rect 55315 2945 55320 2965
rect 55290 2915 55320 2945
rect 55290 2895 55295 2915
rect 55315 2895 55320 2915
rect 55290 2865 55320 2895
rect 55290 2845 55295 2865
rect 55315 2845 55320 2865
rect 55290 2815 55320 2845
rect 55290 2795 55295 2815
rect 55315 2795 55320 2815
rect 55290 2765 55320 2795
rect 55290 2745 55295 2765
rect 55315 2745 55320 2765
rect 55290 2735 55320 2745
rect 55345 3315 55375 3325
rect 55345 3295 55350 3315
rect 55370 3295 55375 3315
rect 55345 3265 55375 3295
rect 55345 3245 55350 3265
rect 55370 3245 55375 3265
rect 55345 3215 55375 3245
rect 55345 3195 55350 3215
rect 55370 3195 55375 3215
rect 55345 3165 55375 3195
rect 55345 3145 55350 3165
rect 55370 3145 55375 3165
rect 55345 3115 55375 3145
rect 55345 3095 55350 3115
rect 55370 3095 55375 3115
rect 55345 3065 55375 3095
rect 55345 3045 55350 3065
rect 55370 3045 55375 3065
rect 55345 3015 55375 3045
rect 55345 2995 55350 3015
rect 55370 2995 55375 3015
rect 55345 2965 55375 2995
rect 55345 2945 55350 2965
rect 55370 2945 55375 2965
rect 55345 2915 55375 2945
rect 55345 2895 55350 2915
rect 55370 2895 55375 2915
rect 55345 2865 55375 2895
rect 55345 2845 55350 2865
rect 55370 2845 55375 2865
rect 55345 2815 55375 2845
rect 55345 2795 55350 2815
rect 55370 2795 55375 2815
rect 55345 2765 55375 2795
rect 55345 2745 55350 2765
rect 55370 2745 55375 2765
rect 55345 2735 55375 2745
rect 55400 3315 55430 3325
rect 55400 3295 55405 3315
rect 55425 3295 55430 3315
rect 55400 3265 55430 3295
rect 55400 3245 55405 3265
rect 55425 3245 55430 3265
rect 55400 3215 55430 3245
rect 55400 3195 55405 3215
rect 55425 3195 55430 3215
rect 55400 3165 55430 3195
rect 55400 3145 55405 3165
rect 55425 3145 55430 3165
rect 55400 3115 55430 3145
rect 55400 3095 55405 3115
rect 55425 3095 55430 3115
rect 55400 3065 55430 3095
rect 55400 3045 55405 3065
rect 55425 3045 55430 3065
rect 55400 3015 55430 3045
rect 55400 2995 55405 3015
rect 55425 2995 55430 3015
rect 55400 2965 55430 2995
rect 55400 2945 55405 2965
rect 55425 2945 55430 2965
rect 55400 2915 55430 2945
rect 55400 2895 55405 2915
rect 55425 2895 55430 2915
rect 55400 2865 55430 2895
rect 55400 2845 55405 2865
rect 55425 2845 55430 2865
rect 55400 2815 55430 2845
rect 55400 2795 55405 2815
rect 55425 2795 55430 2815
rect 55400 2765 55430 2795
rect 55400 2745 55405 2765
rect 55425 2745 55430 2765
rect 55400 2735 55430 2745
rect 55455 3315 55485 3325
rect 55455 3295 55460 3315
rect 55480 3295 55485 3315
rect 55455 3265 55485 3295
rect 55455 3245 55460 3265
rect 55480 3245 55485 3265
rect 55455 3215 55485 3245
rect 55455 3195 55460 3215
rect 55480 3195 55485 3215
rect 55455 3165 55485 3195
rect 55455 3145 55460 3165
rect 55480 3145 55485 3165
rect 55455 3115 55485 3145
rect 55455 3095 55460 3115
rect 55480 3095 55485 3115
rect 55455 3065 55485 3095
rect 55455 3045 55460 3065
rect 55480 3045 55485 3065
rect 55455 3015 55485 3045
rect 55455 2995 55460 3015
rect 55480 2995 55485 3015
rect 55455 2965 55485 2995
rect 55455 2945 55460 2965
rect 55480 2945 55485 2965
rect 55455 2915 55485 2945
rect 55455 2895 55460 2915
rect 55480 2895 55485 2915
rect 55455 2865 55485 2895
rect 55455 2845 55460 2865
rect 55480 2845 55485 2865
rect 55455 2815 55485 2845
rect 55455 2795 55460 2815
rect 55480 2795 55485 2815
rect 55455 2765 55485 2795
rect 55455 2745 55460 2765
rect 55480 2745 55485 2765
rect 55455 2735 55485 2745
rect 55510 3315 55540 3325
rect 55510 3295 55515 3315
rect 55535 3295 55540 3315
rect 55510 3265 55540 3295
rect 55510 3245 55515 3265
rect 55535 3245 55540 3265
rect 55510 3215 55540 3245
rect 55510 3195 55515 3215
rect 55535 3195 55540 3215
rect 55510 3165 55540 3195
rect 55510 3145 55515 3165
rect 55535 3145 55540 3165
rect 55510 3115 55540 3145
rect 55510 3095 55515 3115
rect 55535 3095 55540 3115
rect 55510 3065 55540 3095
rect 55510 3045 55515 3065
rect 55535 3045 55540 3065
rect 55510 3015 55540 3045
rect 55510 2995 55515 3015
rect 55535 2995 55540 3015
rect 55510 2965 55540 2995
rect 55510 2945 55515 2965
rect 55535 2945 55540 2965
rect 55510 2915 55540 2945
rect 55510 2895 55515 2915
rect 55535 2895 55540 2915
rect 55510 2865 55540 2895
rect 55510 2845 55515 2865
rect 55535 2845 55540 2865
rect 55510 2815 55540 2845
rect 55510 2795 55515 2815
rect 55535 2795 55540 2815
rect 55510 2765 55540 2795
rect 55510 2745 55515 2765
rect 55535 2745 55540 2765
rect 55510 2735 55540 2745
rect 55565 3315 55595 3325
rect 55565 3295 55570 3315
rect 55590 3295 55595 3315
rect 55565 3265 55595 3295
rect 55565 3245 55570 3265
rect 55590 3245 55595 3265
rect 55565 3215 55595 3245
rect 55565 3195 55570 3215
rect 55590 3195 55595 3215
rect 55565 3165 55595 3195
rect 55565 3145 55570 3165
rect 55590 3145 55595 3165
rect 55565 3115 55595 3145
rect 55565 3095 55570 3115
rect 55590 3095 55595 3115
rect 55565 3065 55595 3095
rect 55565 3045 55570 3065
rect 55590 3045 55595 3065
rect 55565 3015 55595 3045
rect 55565 2995 55570 3015
rect 55590 2995 55595 3015
rect 55565 2965 55595 2995
rect 55565 2945 55570 2965
rect 55590 2945 55595 2965
rect 55565 2915 55595 2945
rect 55565 2895 55570 2915
rect 55590 2895 55595 2915
rect 55565 2865 55595 2895
rect 55565 2845 55570 2865
rect 55590 2845 55595 2865
rect 55565 2815 55595 2845
rect 55565 2795 55570 2815
rect 55590 2795 55595 2815
rect 55565 2765 55595 2795
rect 55565 2745 55570 2765
rect 55590 2745 55595 2765
rect 55565 2735 55595 2745
rect 55620 3315 55650 3325
rect 55620 3295 55625 3315
rect 55645 3295 55650 3315
rect 55620 3265 55650 3295
rect 55620 3245 55625 3265
rect 55645 3245 55650 3265
rect 55620 3215 55650 3245
rect 55620 3195 55625 3215
rect 55645 3195 55650 3215
rect 55620 3165 55650 3195
rect 55620 3145 55625 3165
rect 55645 3145 55650 3165
rect 55620 3115 55650 3145
rect 55620 3095 55625 3115
rect 55645 3095 55650 3115
rect 55620 3065 55650 3095
rect 55620 3045 55625 3065
rect 55645 3045 55650 3065
rect 55620 3015 55650 3045
rect 55620 2995 55625 3015
rect 55645 2995 55650 3015
rect 55620 2965 55650 2995
rect 55620 2945 55625 2965
rect 55645 2945 55650 2965
rect 55620 2915 55650 2945
rect 55620 2895 55625 2915
rect 55645 2895 55650 2915
rect 55620 2865 55650 2895
rect 55620 2845 55625 2865
rect 55645 2845 55650 2865
rect 55620 2815 55650 2845
rect 55620 2795 55625 2815
rect 55645 2795 55650 2815
rect 55620 2765 55650 2795
rect 55620 2745 55625 2765
rect 55645 2745 55650 2765
rect 55020 2715 55040 2735
rect 55130 2715 55150 2735
rect 55240 2715 55260 2735
rect 55350 2715 55370 2735
rect 55460 2715 55480 2735
rect 55570 2715 55590 2735
rect 54960 2685 54965 2705
rect 54985 2685 54990 2705
rect 54960 2675 54990 2685
rect 55010 2705 55050 2715
rect 55010 2685 55020 2705
rect 55040 2685 55050 2705
rect 55010 2675 55050 2685
rect 55120 2705 55160 2715
rect 55120 2685 55130 2705
rect 55150 2685 55160 2705
rect 55120 2675 55160 2685
rect 55178 2705 55212 2715
rect 55178 2685 55186 2705
rect 55204 2685 55212 2705
rect 55178 2675 55212 2685
rect 55230 2705 55270 2715
rect 55230 2685 55240 2705
rect 55260 2685 55270 2705
rect 55230 2675 55270 2685
rect 55340 2705 55380 2715
rect 55340 2685 55350 2705
rect 55370 2685 55380 2705
rect 55340 2675 55380 2685
rect 55450 2705 55490 2715
rect 55450 2685 55460 2705
rect 55480 2685 55490 2705
rect 55450 2675 55490 2685
rect 55560 2705 55600 2715
rect 55560 2685 55570 2705
rect 55590 2685 55600 2705
rect 55560 2675 55600 2685
rect 55620 2705 55650 2745
rect 55620 2685 55625 2705
rect 55645 2685 55650 2705
rect 55620 2675 55650 2685
rect 55685 3075 55705 3405
rect 56225 3405 56860 3425
rect 56940 3405 57575 3425
rect 56225 3345 56245 3405
rect 56275 3375 56315 3385
rect 56275 3355 56285 3375
rect 56305 3355 56315 3375
rect 56275 3345 56315 3355
rect 56385 3375 56425 3385
rect 56385 3355 56395 3375
rect 56415 3355 56425 3375
rect 56385 3345 56425 3355
rect 56495 3375 56535 3385
rect 56495 3355 56505 3375
rect 56525 3355 56535 3375
rect 56495 3345 56535 3355
rect 56605 3375 56645 3385
rect 56605 3355 56615 3375
rect 56635 3355 56645 3375
rect 56605 3345 56645 3355
rect 56715 3375 56755 3385
rect 56715 3355 56725 3375
rect 56745 3355 56755 3375
rect 56715 3345 56755 3355
rect 56825 3375 56865 3385
rect 56825 3355 56835 3375
rect 56855 3355 56865 3375
rect 56825 3345 56865 3355
rect 56935 3375 56975 3385
rect 56935 3355 56945 3375
rect 56965 3355 56975 3375
rect 56935 3345 56975 3355
rect 57045 3375 57085 3385
rect 57045 3355 57055 3375
rect 57075 3355 57085 3375
rect 57045 3345 57085 3355
rect 57155 3375 57195 3385
rect 57155 3355 57165 3375
rect 57185 3355 57195 3375
rect 57155 3345 57195 3355
rect 57265 3375 57305 3385
rect 57265 3355 57275 3375
rect 57295 3355 57305 3375
rect 57265 3345 57305 3355
rect 57375 3375 57415 3385
rect 57375 3355 57385 3375
rect 57405 3355 57415 3375
rect 57375 3345 57415 3355
rect 57485 3375 57525 3385
rect 57485 3355 57495 3375
rect 57515 3355 57525 3375
rect 57485 3345 57525 3355
rect 57555 3345 57575 3405
rect 56285 3325 56305 3345
rect 56395 3325 56415 3345
rect 56505 3325 56525 3345
rect 56615 3325 56635 3345
rect 56725 3325 56745 3345
rect 56835 3325 56855 3345
rect 56945 3325 56965 3345
rect 57055 3325 57075 3345
rect 57165 3325 57185 3345
rect 57275 3325 57295 3345
rect 57385 3325 57405 3345
rect 57495 3325 57515 3345
rect 56225 3205 56245 3265
rect 56280 3315 56310 3325
rect 56280 3295 56285 3315
rect 56305 3295 56310 3315
rect 56280 3255 56310 3295
rect 56335 3315 56365 3325
rect 56335 3295 56340 3315
rect 56360 3295 56365 3315
rect 56335 3285 56365 3295
rect 56390 3315 56420 3325
rect 56390 3295 56395 3315
rect 56415 3295 56420 3315
rect 56390 3285 56420 3295
rect 56445 3315 56475 3325
rect 56445 3295 56450 3315
rect 56470 3295 56475 3315
rect 56445 3285 56475 3295
rect 56500 3315 56530 3325
rect 56500 3295 56505 3315
rect 56525 3295 56530 3315
rect 56500 3285 56530 3295
rect 56555 3315 56585 3325
rect 56555 3295 56560 3315
rect 56580 3295 56585 3315
rect 56555 3285 56585 3295
rect 56610 3315 56640 3325
rect 56610 3295 56615 3315
rect 56635 3295 56640 3315
rect 56610 3285 56640 3295
rect 56665 3315 56695 3325
rect 56665 3295 56670 3315
rect 56690 3295 56695 3315
rect 56665 3285 56695 3295
rect 56720 3315 56750 3325
rect 56720 3295 56725 3315
rect 56745 3295 56750 3315
rect 56720 3285 56750 3295
rect 56775 3315 56805 3325
rect 56775 3295 56780 3315
rect 56800 3295 56805 3315
rect 56775 3285 56805 3295
rect 56830 3315 56860 3325
rect 56830 3295 56835 3315
rect 56855 3295 56860 3315
rect 56830 3285 56860 3295
rect 56885 3315 56915 3325
rect 56885 3295 56890 3315
rect 56910 3295 56915 3315
rect 56885 3285 56915 3295
rect 56940 3315 56970 3325
rect 56940 3295 56945 3315
rect 56965 3295 56970 3315
rect 56940 3285 56970 3295
rect 56995 3315 57025 3325
rect 56995 3295 57000 3315
rect 57020 3295 57025 3315
rect 56995 3285 57025 3295
rect 57050 3315 57080 3325
rect 57050 3295 57055 3315
rect 57075 3295 57080 3315
rect 57050 3285 57080 3295
rect 57105 3315 57135 3325
rect 57105 3295 57110 3315
rect 57130 3295 57135 3315
rect 57105 3285 57135 3295
rect 57160 3315 57190 3325
rect 57160 3295 57165 3315
rect 57185 3295 57190 3315
rect 57160 3285 57190 3295
rect 57215 3315 57245 3325
rect 57215 3295 57220 3315
rect 57240 3295 57245 3315
rect 57215 3285 57245 3295
rect 57270 3315 57300 3325
rect 57270 3295 57275 3315
rect 57295 3295 57300 3315
rect 57270 3285 57300 3295
rect 57325 3315 57355 3325
rect 57325 3295 57330 3315
rect 57350 3295 57355 3315
rect 57325 3285 57355 3295
rect 57380 3315 57410 3325
rect 57380 3295 57385 3315
rect 57405 3295 57410 3315
rect 57380 3285 57410 3295
rect 57435 3315 57465 3325
rect 57435 3295 57440 3315
rect 57460 3295 57465 3315
rect 57435 3285 57465 3295
rect 57490 3315 57520 3325
rect 57490 3295 57495 3315
rect 57515 3295 57520 3315
rect 56340 3265 56360 3285
rect 56450 3265 56470 3285
rect 56560 3265 56580 3285
rect 56670 3265 56690 3285
rect 56780 3265 56800 3285
rect 56890 3265 56910 3285
rect 57000 3265 57020 3285
rect 57110 3265 57130 3285
rect 57220 3265 57240 3285
rect 57330 3265 57350 3285
rect 57440 3265 57460 3285
rect 56280 3235 56285 3255
rect 56305 3235 56310 3255
rect 56280 3225 56310 3235
rect 56330 3255 56370 3265
rect 56330 3235 56340 3255
rect 56360 3235 56370 3255
rect 56330 3225 56370 3235
rect 56440 3255 56480 3265
rect 56440 3235 56450 3255
rect 56470 3235 56480 3255
rect 56440 3225 56480 3235
rect 56497 3255 56533 3265
rect 56497 3235 56505 3255
rect 56525 3235 56533 3255
rect 56497 3225 56533 3235
rect 56550 3255 56590 3265
rect 56550 3235 56560 3255
rect 56580 3235 56590 3255
rect 56550 3225 56590 3235
rect 56660 3255 56700 3265
rect 56660 3235 56670 3255
rect 56690 3235 56700 3255
rect 56660 3225 56700 3235
rect 56770 3255 56810 3265
rect 56770 3235 56780 3255
rect 56800 3235 56810 3255
rect 56770 3225 56810 3235
rect 56880 3255 56920 3265
rect 56880 3235 56890 3255
rect 56910 3235 56920 3255
rect 56880 3225 56920 3235
rect 56990 3255 57030 3265
rect 56990 3235 57000 3255
rect 57020 3235 57030 3255
rect 56990 3225 57030 3235
rect 57100 3255 57140 3265
rect 57100 3235 57110 3255
rect 57130 3235 57140 3255
rect 57100 3225 57140 3235
rect 57210 3255 57250 3265
rect 57210 3235 57220 3255
rect 57240 3235 57250 3255
rect 57210 3225 57250 3235
rect 57320 3255 57360 3265
rect 57320 3235 57330 3255
rect 57350 3235 57360 3255
rect 57320 3225 57360 3235
rect 57430 3255 57470 3265
rect 57430 3235 57440 3255
rect 57460 3235 57470 3255
rect 57430 3225 57470 3235
rect 57490 3255 57520 3295
rect 57490 3235 57495 3255
rect 57515 3235 57520 3255
rect 57490 3225 57520 3235
rect 56285 3205 56305 3225
rect 57495 3205 57515 3225
rect 57555 3205 57575 3265
rect 56225 3185 56860 3205
rect 56940 3185 57575 3205
rect 58095 3405 58455 3425
rect 58535 3405 58895 3425
rect 54965 2655 54985 2675
rect 55625 2655 55645 2675
rect 55685 2655 55705 2980
rect 58095 3075 58115 3405
rect 58145 3375 58185 3385
rect 58145 3355 58155 3375
rect 58175 3355 58185 3375
rect 58145 3345 58185 3355
rect 58255 3375 58295 3385
rect 58255 3355 58265 3375
rect 58285 3355 58295 3375
rect 58255 3345 58295 3355
rect 58365 3375 58405 3385
rect 58365 3355 58375 3375
rect 58395 3355 58405 3375
rect 58365 3345 58405 3355
rect 58475 3375 58515 3385
rect 58475 3355 58485 3375
rect 58505 3355 58515 3375
rect 58475 3345 58515 3355
rect 58585 3375 58625 3385
rect 58585 3355 58595 3375
rect 58615 3355 58625 3375
rect 58585 3345 58625 3355
rect 58695 3375 58735 3385
rect 58695 3355 58705 3375
rect 58725 3355 58735 3375
rect 58695 3345 58735 3355
rect 58805 3375 58845 3385
rect 58805 3355 58815 3375
rect 58835 3355 58845 3375
rect 58805 3345 58845 3355
rect 58155 3325 58175 3345
rect 58265 3325 58285 3345
rect 58375 3325 58395 3345
rect 58485 3325 58505 3345
rect 58595 3325 58615 3345
rect 58705 3325 58725 3345
rect 58815 3325 58835 3345
rect 56015 2950 56375 2970
rect 56455 2950 56815 2970
rect 56015 2890 56035 2950
rect 56145 2920 56175 2930
rect 56145 2900 56150 2920
rect 56170 2900 56175 2920
rect 56145 2890 56175 2900
rect 56192 2920 56218 2930
rect 56192 2900 56195 2920
rect 56215 2900 56218 2920
rect 56192 2890 56218 2900
rect 56292 2920 56318 2930
rect 56292 2900 56295 2920
rect 56315 2900 56318 2920
rect 56292 2890 56318 2900
rect 56345 2920 56375 2930
rect 56345 2900 56350 2920
rect 56370 2900 56375 2920
rect 56345 2890 56375 2900
rect 56402 2920 56428 2930
rect 56402 2900 56405 2920
rect 56425 2900 56428 2920
rect 56402 2890 56428 2900
rect 56455 2920 56485 2930
rect 56455 2900 56460 2920
rect 56480 2900 56485 2920
rect 56455 2890 56485 2900
rect 56512 2920 56538 2930
rect 56512 2900 56515 2920
rect 56535 2900 56538 2920
rect 56512 2890 56538 2900
rect 56560 2920 56600 2930
rect 56560 2900 56570 2920
rect 56590 2900 56600 2920
rect 56560 2890 56600 2900
rect 56622 2920 56648 2930
rect 56622 2900 56625 2920
rect 56645 2900 56648 2920
rect 56622 2890 56648 2900
rect 56795 2890 56815 2950
rect 56005 2830 56015 2870
rect 56192 2870 56210 2890
rect 56295 2870 56315 2890
rect 56405 2870 56425 2890
rect 56460 2870 56480 2890
rect 56515 2870 56535 2890
rect 56625 2870 56645 2890
rect 56035 2830 56045 2870
rect 56070 2860 56100 2870
rect 56070 2840 56075 2860
rect 56095 2840 56100 2860
rect 56015 2750 56035 2810
rect 56070 2800 56100 2840
rect 56125 2860 56155 2870
rect 56125 2840 56130 2860
rect 56150 2840 56155 2860
rect 56125 2830 56155 2840
rect 56180 2860 56210 2870
rect 56180 2840 56185 2860
rect 56205 2840 56210 2860
rect 56180 2830 56210 2840
rect 56235 2860 56265 2870
rect 56235 2840 56240 2860
rect 56260 2840 56265 2860
rect 56235 2830 56265 2840
rect 56290 2860 56320 2870
rect 56290 2840 56295 2860
rect 56315 2840 56320 2860
rect 56290 2830 56320 2840
rect 56345 2860 56375 2870
rect 56345 2840 56350 2860
rect 56370 2840 56375 2860
rect 56345 2830 56375 2840
rect 56400 2860 56430 2870
rect 56400 2840 56405 2860
rect 56425 2840 56430 2860
rect 56400 2830 56430 2840
rect 56455 2860 56485 2870
rect 56455 2840 56460 2860
rect 56480 2840 56485 2860
rect 56455 2830 56485 2840
rect 56510 2860 56540 2870
rect 56510 2840 56515 2860
rect 56535 2840 56540 2860
rect 56510 2830 56540 2840
rect 56565 2860 56595 2870
rect 56565 2840 56570 2860
rect 56590 2840 56595 2860
rect 56565 2830 56595 2840
rect 56620 2860 56650 2870
rect 56620 2840 56625 2860
rect 56645 2840 56650 2860
rect 56620 2830 56650 2840
rect 56675 2860 56705 2870
rect 56675 2840 56680 2860
rect 56700 2840 56705 2860
rect 56675 2830 56705 2840
rect 56130 2810 56150 2830
rect 56235 2810 56255 2830
rect 56350 2810 56370 2830
rect 56455 2810 56475 2830
rect 56570 2810 56590 2830
rect 56685 2810 56705 2830
rect 56730 2860 56760 2870
rect 56730 2840 56735 2860
rect 56755 2840 56760 2860
rect 56070 2780 56075 2800
rect 56095 2780 56100 2800
rect 56070 2770 56100 2780
rect 56120 2800 56160 2810
rect 56120 2780 56130 2800
rect 56150 2780 56160 2800
rect 56120 2770 56160 2780
rect 56215 2800 56255 2810
rect 56215 2780 56225 2800
rect 56245 2780 56255 2800
rect 56215 2770 56255 2780
rect 56272 2800 56304 2810
rect 56272 2780 56278 2800
rect 56295 2780 56304 2800
rect 56272 2770 56304 2780
rect 56340 2800 56380 2810
rect 56340 2780 56350 2800
rect 56370 2780 56380 2800
rect 56340 2770 56380 2780
rect 56435 2800 56475 2810
rect 56435 2780 56445 2800
rect 56465 2780 56475 2800
rect 56435 2770 56475 2780
rect 56492 2800 56524 2810
rect 56492 2780 56498 2800
rect 56515 2780 56524 2800
rect 56492 2770 56524 2780
rect 56560 2800 56600 2810
rect 56560 2780 56570 2800
rect 56590 2780 56600 2800
rect 56560 2770 56600 2780
rect 56636 2800 56668 2810
rect 56636 2780 56645 2800
rect 56662 2780 56668 2800
rect 56636 2770 56668 2780
rect 56685 2800 56711 2810
rect 56685 2780 56688 2800
rect 56708 2780 56711 2800
rect 56685 2770 56711 2780
rect 56730 2800 56760 2840
rect 56785 2830 56795 2870
rect 56985 2950 57345 2970
rect 57425 2950 57785 2970
rect 56985 2890 57005 2950
rect 57113 2920 57143 2930
rect 57113 2900 57118 2920
rect 57138 2900 57143 2920
rect 57113 2890 57143 2900
rect 57162 2920 57188 2930
rect 57162 2900 57165 2920
rect 57185 2900 57188 2920
rect 57162 2890 57188 2900
rect 57262 2920 57288 2930
rect 57262 2900 57265 2920
rect 57285 2900 57288 2920
rect 57262 2890 57288 2900
rect 57310 2920 57350 2930
rect 57310 2900 57320 2920
rect 57340 2900 57350 2920
rect 57310 2890 57350 2900
rect 57372 2920 57398 2930
rect 57372 2900 57375 2920
rect 57395 2900 57398 2920
rect 57372 2890 57398 2900
rect 57482 2920 57508 2930
rect 57482 2900 57485 2920
rect 57505 2900 57508 2920
rect 57482 2890 57508 2900
rect 57530 2920 57570 2930
rect 57530 2900 57540 2920
rect 57560 2900 57570 2920
rect 57530 2890 57570 2900
rect 57592 2920 57618 2930
rect 57592 2900 57595 2920
rect 57615 2900 57618 2920
rect 57592 2890 57618 2900
rect 57765 2890 57785 2950
rect 56730 2780 56735 2800
rect 56755 2780 56760 2800
rect 56730 2770 56760 2780
rect 56815 2830 56825 2870
rect 56975 2830 56985 2870
rect 57162 2870 57180 2890
rect 57265 2870 57285 2890
rect 57375 2870 57395 2890
rect 57485 2870 57505 2890
rect 57595 2870 57615 2890
rect 56075 2750 56095 2770
rect 56735 2750 56755 2770
rect 56795 2750 56815 2810
rect 56015 2730 56375 2750
rect 56455 2730 56815 2750
rect 57005 2830 57015 2870
rect 57040 2860 57070 2870
rect 57040 2840 57045 2860
rect 57065 2840 57070 2860
rect 56985 2750 57005 2810
rect 57040 2800 57070 2840
rect 57095 2860 57125 2870
rect 57095 2840 57100 2860
rect 57120 2840 57125 2860
rect 57095 2830 57125 2840
rect 57150 2860 57180 2870
rect 57150 2840 57155 2860
rect 57175 2840 57180 2860
rect 57150 2830 57180 2840
rect 57205 2860 57235 2870
rect 57205 2840 57210 2860
rect 57230 2840 57235 2860
rect 57205 2830 57235 2840
rect 57260 2860 57290 2870
rect 57260 2840 57265 2860
rect 57285 2840 57290 2860
rect 57260 2830 57290 2840
rect 57315 2860 57345 2870
rect 57315 2840 57320 2860
rect 57340 2840 57345 2860
rect 57315 2830 57345 2840
rect 57370 2860 57400 2870
rect 57370 2840 57375 2860
rect 57395 2840 57400 2860
rect 57370 2830 57400 2840
rect 57425 2860 57455 2870
rect 57425 2840 57430 2860
rect 57450 2840 57455 2860
rect 57425 2830 57455 2840
rect 57480 2860 57510 2870
rect 57480 2840 57485 2860
rect 57505 2840 57510 2860
rect 57480 2830 57510 2840
rect 57535 2860 57565 2870
rect 57535 2840 57540 2860
rect 57560 2840 57565 2860
rect 57535 2830 57565 2840
rect 57590 2860 57620 2870
rect 57590 2840 57595 2860
rect 57615 2840 57620 2860
rect 57590 2830 57620 2840
rect 57645 2860 57675 2870
rect 57645 2840 57650 2860
rect 57670 2840 57675 2860
rect 57645 2830 57675 2840
rect 57100 2810 57120 2830
rect 57205 2810 57225 2830
rect 57320 2810 57340 2830
rect 57425 2810 57445 2830
rect 57540 2810 57560 2830
rect 57655 2810 57675 2830
rect 57700 2860 57730 2870
rect 57700 2840 57705 2860
rect 57725 2840 57730 2860
rect 57040 2780 57045 2800
rect 57065 2780 57070 2800
rect 57040 2770 57070 2780
rect 57090 2800 57130 2810
rect 57090 2780 57100 2800
rect 57120 2780 57130 2800
rect 57090 2770 57130 2780
rect 57185 2800 57225 2810
rect 57185 2780 57195 2800
rect 57215 2780 57225 2800
rect 57185 2770 57225 2780
rect 57242 2800 57274 2810
rect 57242 2780 57248 2800
rect 57265 2780 57274 2800
rect 57242 2770 57274 2780
rect 57310 2800 57350 2810
rect 57310 2780 57320 2800
rect 57340 2780 57350 2800
rect 57310 2770 57350 2780
rect 57405 2800 57445 2810
rect 57405 2780 57415 2800
rect 57435 2780 57445 2800
rect 57405 2770 57445 2780
rect 57462 2800 57494 2810
rect 57462 2780 57468 2800
rect 57485 2780 57494 2800
rect 57462 2770 57494 2780
rect 57530 2800 57570 2810
rect 57530 2780 57540 2800
rect 57560 2780 57570 2800
rect 57530 2770 57570 2780
rect 57606 2800 57638 2810
rect 57606 2780 57615 2800
rect 57632 2780 57638 2800
rect 57606 2770 57638 2780
rect 57655 2800 57681 2810
rect 57655 2780 57658 2800
rect 57678 2780 57681 2800
rect 57655 2770 57681 2780
rect 57700 2800 57730 2840
rect 57700 2780 57705 2800
rect 57725 2780 57730 2800
rect 57700 2770 57730 2780
rect 57045 2750 57065 2770
rect 57705 2750 57725 2770
rect 57765 2750 57785 2810
rect 56985 2730 57345 2750
rect 57425 2730 57785 2750
rect 56680 2715 56710 2730
rect 54555 2630 54565 2640
rect 54905 2635 55265 2655
rect 55345 2635 55705 2655
rect 58095 2655 58115 2980
rect 58150 3315 58180 3325
rect 58150 3295 58155 3315
rect 58175 3295 58180 3315
rect 58150 3265 58180 3295
rect 58150 3245 58155 3265
rect 58175 3245 58180 3265
rect 58150 3215 58180 3245
rect 58150 3195 58155 3215
rect 58175 3195 58180 3215
rect 58150 3165 58180 3195
rect 58150 3145 58155 3165
rect 58175 3145 58180 3165
rect 58150 3115 58180 3145
rect 58150 3095 58155 3115
rect 58175 3095 58180 3115
rect 58150 3065 58180 3095
rect 58150 3045 58155 3065
rect 58175 3045 58180 3065
rect 58150 3015 58180 3045
rect 58150 2995 58155 3015
rect 58175 2995 58180 3015
rect 58150 2965 58180 2995
rect 58150 2945 58155 2965
rect 58175 2945 58180 2965
rect 58150 2915 58180 2945
rect 58150 2895 58155 2915
rect 58175 2895 58180 2915
rect 58150 2865 58180 2895
rect 58150 2845 58155 2865
rect 58175 2845 58180 2865
rect 58150 2815 58180 2845
rect 58150 2795 58155 2815
rect 58175 2795 58180 2815
rect 58150 2765 58180 2795
rect 58150 2745 58155 2765
rect 58175 2745 58180 2765
rect 58150 2705 58180 2745
rect 58205 3315 58235 3325
rect 58205 3295 58210 3315
rect 58230 3295 58235 3315
rect 58205 3265 58235 3295
rect 58205 3245 58210 3265
rect 58230 3245 58235 3265
rect 58205 3215 58235 3245
rect 58205 3195 58210 3215
rect 58230 3195 58235 3215
rect 58205 3165 58235 3195
rect 58205 3145 58210 3165
rect 58230 3145 58235 3165
rect 58205 3115 58235 3145
rect 58205 3095 58210 3115
rect 58230 3095 58235 3115
rect 58205 3065 58235 3095
rect 58205 3045 58210 3065
rect 58230 3045 58235 3065
rect 58205 3015 58235 3045
rect 58205 2995 58210 3015
rect 58230 2995 58235 3015
rect 58205 2965 58235 2995
rect 58205 2945 58210 2965
rect 58230 2945 58235 2965
rect 58205 2915 58235 2945
rect 58205 2895 58210 2915
rect 58230 2895 58235 2915
rect 58205 2865 58235 2895
rect 58205 2845 58210 2865
rect 58230 2845 58235 2865
rect 58205 2815 58235 2845
rect 58205 2795 58210 2815
rect 58230 2795 58235 2815
rect 58205 2765 58235 2795
rect 58205 2745 58210 2765
rect 58230 2745 58235 2765
rect 58205 2735 58235 2745
rect 58260 3315 58290 3325
rect 58260 3295 58265 3315
rect 58285 3295 58290 3315
rect 58260 3265 58290 3295
rect 58260 3245 58265 3265
rect 58285 3245 58290 3265
rect 58260 3215 58290 3245
rect 58260 3195 58265 3215
rect 58285 3195 58290 3215
rect 58260 3165 58290 3195
rect 58260 3145 58265 3165
rect 58285 3145 58290 3165
rect 58260 3115 58290 3145
rect 58260 3095 58265 3115
rect 58285 3095 58290 3115
rect 58260 3065 58290 3095
rect 58260 3045 58265 3065
rect 58285 3045 58290 3065
rect 58260 3015 58290 3045
rect 58260 2995 58265 3015
rect 58285 2995 58290 3015
rect 58260 2965 58290 2995
rect 58260 2945 58265 2965
rect 58285 2945 58290 2965
rect 58260 2915 58290 2945
rect 58260 2895 58265 2915
rect 58285 2895 58290 2915
rect 58260 2865 58290 2895
rect 58260 2845 58265 2865
rect 58285 2845 58290 2865
rect 58260 2815 58290 2845
rect 58260 2795 58265 2815
rect 58285 2795 58290 2815
rect 58260 2765 58290 2795
rect 58260 2745 58265 2765
rect 58285 2745 58290 2765
rect 58260 2735 58290 2745
rect 58315 3315 58345 3325
rect 58315 3295 58320 3315
rect 58340 3295 58345 3315
rect 58315 3265 58345 3295
rect 58315 3245 58320 3265
rect 58340 3245 58345 3265
rect 58315 3215 58345 3245
rect 58315 3195 58320 3215
rect 58340 3195 58345 3215
rect 58315 3165 58345 3195
rect 58315 3145 58320 3165
rect 58340 3145 58345 3165
rect 58315 3115 58345 3145
rect 58315 3095 58320 3115
rect 58340 3095 58345 3115
rect 58315 3065 58345 3095
rect 58315 3045 58320 3065
rect 58340 3045 58345 3065
rect 58315 3015 58345 3045
rect 58315 2995 58320 3015
rect 58340 2995 58345 3015
rect 58315 2965 58345 2995
rect 58315 2945 58320 2965
rect 58340 2945 58345 2965
rect 58315 2915 58345 2945
rect 58315 2895 58320 2915
rect 58340 2895 58345 2915
rect 58315 2865 58345 2895
rect 58315 2845 58320 2865
rect 58340 2845 58345 2865
rect 58315 2815 58345 2845
rect 58315 2795 58320 2815
rect 58340 2795 58345 2815
rect 58315 2765 58345 2795
rect 58315 2745 58320 2765
rect 58340 2745 58345 2765
rect 58315 2735 58345 2745
rect 58370 3315 58400 3325
rect 58370 3295 58375 3315
rect 58395 3295 58400 3315
rect 58370 3265 58400 3295
rect 58370 3245 58375 3265
rect 58395 3245 58400 3265
rect 58370 3215 58400 3245
rect 58370 3195 58375 3215
rect 58395 3195 58400 3215
rect 58370 3165 58400 3195
rect 58370 3145 58375 3165
rect 58395 3145 58400 3165
rect 58370 3115 58400 3145
rect 58370 3095 58375 3115
rect 58395 3095 58400 3115
rect 58370 3065 58400 3095
rect 58370 3045 58375 3065
rect 58395 3045 58400 3065
rect 58370 3015 58400 3045
rect 58370 2995 58375 3015
rect 58395 2995 58400 3015
rect 58370 2965 58400 2995
rect 58370 2945 58375 2965
rect 58395 2945 58400 2965
rect 58370 2915 58400 2945
rect 58370 2895 58375 2915
rect 58395 2895 58400 2915
rect 58370 2865 58400 2895
rect 58370 2845 58375 2865
rect 58395 2845 58400 2865
rect 58370 2815 58400 2845
rect 58370 2795 58375 2815
rect 58395 2795 58400 2815
rect 58370 2765 58400 2795
rect 58370 2745 58375 2765
rect 58395 2745 58400 2765
rect 58370 2735 58400 2745
rect 58425 3315 58455 3325
rect 58425 3295 58430 3315
rect 58450 3295 58455 3315
rect 58425 3265 58455 3295
rect 58425 3245 58430 3265
rect 58450 3245 58455 3265
rect 58425 3215 58455 3245
rect 58425 3195 58430 3215
rect 58450 3195 58455 3215
rect 58425 3165 58455 3195
rect 58425 3145 58430 3165
rect 58450 3145 58455 3165
rect 58425 3115 58455 3145
rect 58425 3095 58430 3115
rect 58450 3095 58455 3115
rect 58425 3065 58455 3095
rect 58425 3045 58430 3065
rect 58450 3045 58455 3065
rect 58425 3015 58455 3045
rect 58425 2995 58430 3015
rect 58450 2995 58455 3015
rect 58425 2965 58455 2995
rect 58425 2945 58430 2965
rect 58450 2945 58455 2965
rect 58425 2915 58455 2945
rect 58425 2895 58430 2915
rect 58450 2895 58455 2915
rect 58425 2865 58455 2895
rect 58425 2845 58430 2865
rect 58450 2845 58455 2865
rect 58425 2815 58455 2845
rect 58425 2795 58430 2815
rect 58450 2795 58455 2815
rect 58425 2765 58455 2795
rect 58425 2745 58430 2765
rect 58450 2745 58455 2765
rect 58425 2735 58455 2745
rect 58480 3315 58510 3325
rect 58480 3295 58485 3315
rect 58505 3295 58510 3315
rect 58480 3265 58510 3295
rect 58480 3245 58485 3265
rect 58505 3245 58510 3265
rect 58480 3215 58510 3245
rect 58480 3195 58485 3215
rect 58505 3195 58510 3215
rect 58480 3165 58510 3195
rect 58480 3145 58485 3165
rect 58505 3145 58510 3165
rect 58480 3115 58510 3145
rect 58480 3095 58485 3115
rect 58505 3095 58510 3115
rect 58480 3065 58510 3095
rect 58480 3045 58485 3065
rect 58505 3045 58510 3065
rect 58480 3015 58510 3045
rect 58480 2995 58485 3015
rect 58505 2995 58510 3015
rect 58480 2965 58510 2995
rect 58480 2945 58485 2965
rect 58505 2945 58510 2965
rect 58480 2915 58510 2945
rect 58480 2895 58485 2915
rect 58505 2895 58510 2915
rect 58480 2865 58510 2895
rect 58480 2845 58485 2865
rect 58505 2845 58510 2865
rect 58480 2815 58510 2845
rect 58480 2795 58485 2815
rect 58505 2795 58510 2815
rect 58480 2765 58510 2795
rect 58480 2745 58485 2765
rect 58505 2745 58510 2765
rect 58480 2735 58510 2745
rect 58535 3315 58565 3325
rect 58535 3295 58540 3315
rect 58560 3295 58565 3315
rect 58535 3265 58565 3295
rect 58535 3245 58540 3265
rect 58560 3245 58565 3265
rect 58535 3215 58565 3245
rect 58535 3195 58540 3215
rect 58560 3195 58565 3215
rect 58535 3165 58565 3195
rect 58535 3145 58540 3165
rect 58560 3145 58565 3165
rect 58535 3115 58565 3145
rect 58535 3095 58540 3115
rect 58560 3095 58565 3115
rect 58535 3065 58565 3095
rect 58535 3045 58540 3065
rect 58560 3045 58565 3065
rect 58535 3015 58565 3045
rect 58535 2995 58540 3015
rect 58560 2995 58565 3015
rect 58535 2965 58565 2995
rect 58535 2945 58540 2965
rect 58560 2945 58565 2965
rect 58535 2915 58565 2945
rect 58535 2895 58540 2915
rect 58560 2895 58565 2915
rect 58535 2865 58565 2895
rect 58535 2845 58540 2865
rect 58560 2845 58565 2865
rect 58535 2815 58565 2845
rect 58535 2795 58540 2815
rect 58560 2795 58565 2815
rect 58535 2765 58565 2795
rect 58535 2745 58540 2765
rect 58560 2745 58565 2765
rect 58535 2735 58565 2745
rect 58590 3315 58620 3325
rect 58590 3295 58595 3315
rect 58615 3295 58620 3315
rect 58590 3265 58620 3295
rect 58590 3245 58595 3265
rect 58615 3245 58620 3265
rect 58590 3215 58620 3245
rect 58590 3195 58595 3215
rect 58615 3195 58620 3215
rect 58590 3165 58620 3195
rect 58590 3145 58595 3165
rect 58615 3145 58620 3165
rect 58590 3115 58620 3145
rect 58590 3095 58595 3115
rect 58615 3095 58620 3115
rect 58590 3065 58620 3095
rect 58590 3045 58595 3065
rect 58615 3045 58620 3065
rect 58590 3015 58620 3045
rect 58590 2995 58595 3015
rect 58615 2995 58620 3015
rect 58590 2965 58620 2995
rect 58590 2945 58595 2965
rect 58615 2945 58620 2965
rect 58590 2915 58620 2945
rect 58590 2895 58595 2915
rect 58615 2895 58620 2915
rect 58590 2865 58620 2895
rect 58590 2845 58595 2865
rect 58615 2845 58620 2865
rect 58590 2815 58620 2845
rect 58590 2795 58595 2815
rect 58615 2795 58620 2815
rect 58590 2765 58620 2795
rect 58590 2745 58595 2765
rect 58615 2745 58620 2765
rect 58590 2735 58620 2745
rect 58645 3315 58675 3325
rect 58645 3295 58650 3315
rect 58670 3295 58675 3315
rect 58645 3265 58675 3295
rect 58645 3245 58650 3265
rect 58670 3245 58675 3265
rect 58645 3215 58675 3245
rect 58645 3195 58650 3215
rect 58670 3195 58675 3215
rect 58645 3165 58675 3195
rect 58645 3145 58650 3165
rect 58670 3145 58675 3165
rect 58645 3115 58675 3145
rect 58645 3095 58650 3115
rect 58670 3095 58675 3115
rect 58645 3065 58675 3095
rect 58645 3045 58650 3065
rect 58670 3045 58675 3065
rect 58645 3015 58675 3045
rect 58645 2995 58650 3015
rect 58670 2995 58675 3015
rect 58645 2965 58675 2995
rect 58645 2945 58650 2965
rect 58670 2945 58675 2965
rect 58645 2915 58675 2945
rect 58645 2895 58650 2915
rect 58670 2895 58675 2915
rect 58645 2865 58675 2895
rect 58645 2845 58650 2865
rect 58670 2845 58675 2865
rect 58645 2815 58675 2845
rect 58645 2795 58650 2815
rect 58670 2795 58675 2815
rect 58645 2765 58675 2795
rect 58645 2745 58650 2765
rect 58670 2745 58675 2765
rect 58645 2735 58675 2745
rect 58700 3315 58730 3325
rect 58700 3295 58705 3315
rect 58725 3295 58730 3315
rect 58700 3265 58730 3295
rect 58700 3245 58705 3265
rect 58725 3245 58730 3265
rect 58700 3215 58730 3245
rect 58700 3195 58705 3215
rect 58725 3195 58730 3215
rect 58700 3165 58730 3195
rect 58700 3145 58705 3165
rect 58725 3145 58730 3165
rect 58700 3115 58730 3145
rect 58700 3095 58705 3115
rect 58725 3095 58730 3115
rect 58700 3065 58730 3095
rect 58700 3045 58705 3065
rect 58725 3045 58730 3065
rect 58700 3015 58730 3045
rect 58700 2995 58705 3015
rect 58725 2995 58730 3015
rect 58700 2965 58730 2995
rect 58700 2945 58705 2965
rect 58725 2945 58730 2965
rect 58700 2915 58730 2945
rect 58700 2895 58705 2915
rect 58725 2895 58730 2915
rect 58700 2865 58730 2895
rect 58700 2845 58705 2865
rect 58725 2845 58730 2865
rect 58700 2815 58730 2845
rect 58700 2795 58705 2815
rect 58725 2795 58730 2815
rect 58700 2765 58730 2795
rect 58700 2745 58705 2765
rect 58725 2745 58730 2765
rect 58700 2735 58730 2745
rect 58755 3315 58785 3325
rect 58755 3295 58760 3315
rect 58780 3295 58785 3315
rect 58755 3265 58785 3295
rect 58755 3245 58760 3265
rect 58780 3245 58785 3265
rect 58755 3215 58785 3245
rect 58755 3195 58760 3215
rect 58780 3195 58785 3215
rect 58755 3165 58785 3195
rect 58755 3145 58760 3165
rect 58780 3145 58785 3165
rect 58755 3115 58785 3145
rect 58755 3095 58760 3115
rect 58780 3095 58785 3115
rect 58755 3065 58785 3095
rect 58755 3045 58760 3065
rect 58780 3045 58785 3065
rect 58755 3015 58785 3045
rect 58755 2995 58760 3015
rect 58780 2995 58785 3015
rect 58755 2965 58785 2995
rect 58755 2945 58760 2965
rect 58780 2945 58785 2965
rect 58755 2915 58785 2945
rect 58755 2895 58760 2915
rect 58780 2895 58785 2915
rect 58755 2865 58785 2895
rect 58755 2845 58760 2865
rect 58780 2845 58785 2865
rect 58755 2815 58785 2845
rect 58755 2795 58760 2815
rect 58780 2795 58785 2815
rect 58755 2765 58785 2795
rect 58755 2745 58760 2765
rect 58780 2745 58785 2765
rect 58755 2735 58785 2745
rect 58810 3315 58840 3325
rect 58810 3295 58815 3315
rect 58835 3295 58840 3315
rect 58810 3265 58840 3295
rect 58810 3245 58815 3265
rect 58835 3245 58840 3265
rect 58810 3215 58840 3245
rect 58810 3195 58815 3215
rect 58835 3195 58840 3215
rect 58810 3165 58840 3195
rect 58810 3145 58815 3165
rect 58835 3145 58840 3165
rect 58810 3115 58840 3145
rect 58810 3095 58815 3115
rect 58835 3095 58840 3115
rect 58810 3065 58840 3095
rect 58810 3045 58815 3065
rect 58835 3045 58840 3065
rect 58810 3015 58840 3045
rect 58810 2995 58815 3015
rect 58835 2995 58840 3015
rect 58810 2965 58840 2995
rect 58810 2945 58815 2965
rect 58835 2945 58840 2965
rect 58810 2915 58840 2945
rect 58810 2895 58815 2915
rect 58835 2895 58840 2915
rect 58810 2865 58840 2895
rect 58810 2845 58815 2865
rect 58835 2845 58840 2865
rect 58810 2815 58840 2845
rect 58810 2795 58815 2815
rect 58835 2795 58840 2815
rect 58810 2765 58840 2795
rect 58810 2745 58815 2765
rect 58835 2745 58840 2765
rect 58210 2715 58230 2735
rect 58320 2715 58340 2735
rect 58430 2715 58450 2735
rect 58540 2715 58560 2735
rect 58650 2715 58670 2735
rect 58760 2715 58780 2735
rect 58150 2685 58155 2705
rect 58175 2685 58180 2705
rect 58150 2675 58180 2685
rect 58200 2705 58240 2715
rect 58200 2685 58210 2705
rect 58230 2685 58240 2705
rect 58200 2675 58240 2685
rect 58310 2705 58350 2715
rect 58310 2685 58320 2705
rect 58340 2685 58350 2705
rect 58310 2675 58350 2685
rect 58420 2705 58460 2715
rect 58420 2685 58430 2705
rect 58450 2685 58460 2705
rect 58420 2675 58460 2685
rect 58530 2705 58570 2715
rect 58530 2685 58540 2705
rect 58560 2685 58570 2705
rect 58530 2675 58570 2685
rect 58588 2705 58622 2715
rect 58588 2685 58596 2705
rect 58614 2685 58622 2705
rect 58588 2675 58622 2685
rect 58640 2705 58680 2715
rect 58640 2685 58650 2705
rect 58670 2685 58680 2705
rect 58640 2675 58680 2685
rect 58750 2705 58790 2715
rect 58750 2685 58760 2705
rect 58780 2685 58790 2705
rect 58750 2675 58790 2685
rect 58810 2705 58840 2745
rect 58810 2685 58815 2705
rect 58835 2685 58840 2705
rect 58810 2675 58840 2685
rect 58875 3075 58895 3405
rect 58155 2655 58175 2675
rect 58815 2655 58835 2675
rect 58875 2655 58895 2980
rect 58095 2635 58455 2655
rect 58535 2635 58895 2655
rect 59035 3345 59315 3365
rect 59035 3040 59055 3345
rect 59105 3320 59246 3325
rect 59105 3290 59111 3320
rect 59141 3290 59160 3320
rect 59190 3290 59210 3320
rect 59240 3290 59246 3320
rect 59105 3285 59246 3290
rect 59035 2660 59055 2945
rect 59295 3040 59315 3345
rect 59105 2715 59246 2720
rect 59105 2685 59111 2715
rect 59141 2685 59160 2715
rect 59190 2685 59210 2715
rect 59240 2685 59246 2715
rect 59105 2680 59246 2685
rect 59295 2660 59315 2945
rect 59035 2640 59135 2660
rect 59215 2650 59315 2660
rect 59215 2640 59245 2650
rect 54525 2620 54565 2630
rect 55285 2625 55295 2635
rect 55315 2625 55325 2635
rect 55285 2615 55325 2625
rect 58475 2625 58485 2635
rect 58505 2625 58515 2635
rect 58475 2615 58515 2625
rect 59235 2630 59245 2640
rect 59265 2640 59315 2650
rect 59265 2630 59275 2640
rect 59235 2620 59275 2630
rect 56500 2535 56860 2555
rect 56940 2535 57300 2555
rect 55285 2475 55325 2485
rect 55285 2465 55295 2475
rect 55315 2465 55325 2475
rect 56500 2465 56520 2535
rect 56560 2515 56580 2535
rect 57220 2515 57240 2535
rect 54905 2445 55265 2465
rect 55345 2445 55705 2465
rect 54525 2310 54565 2320
rect 54525 2300 54535 2310
rect 54555 2300 54565 2310
rect 54905 2310 54925 2445
rect 55010 2415 55050 2425
rect 55010 2395 55020 2415
rect 55040 2395 55050 2415
rect 55010 2385 55050 2395
rect 55120 2415 55160 2425
rect 55120 2395 55130 2415
rect 55150 2395 55160 2415
rect 55120 2385 55160 2395
rect 55230 2415 55270 2425
rect 55230 2395 55240 2415
rect 55260 2395 55270 2415
rect 55230 2385 55270 2395
rect 55340 2415 55380 2425
rect 55340 2395 55350 2415
rect 55370 2395 55380 2415
rect 55340 2385 55380 2395
rect 55450 2415 55490 2425
rect 55450 2395 55460 2415
rect 55480 2395 55490 2415
rect 55450 2385 55490 2395
rect 55560 2415 55600 2425
rect 55560 2395 55570 2415
rect 55590 2395 55600 2415
rect 55560 2385 55600 2395
rect 55020 2365 55040 2385
rect 55130 2365 55150 2385
rect 55240 2365 55260 2385
rect 55350 2365 55370 2385
rect 55460 2365 55480 2385
rect 55570 2365 55590 2385
rect 54400 2280 54535 2300
rect 54615 2280 54755 2300
rect 54400 1945 54420 2280
rect 54470 2226 54685 2246
rect 54470 2209 54505 2226
rect 54650 2209 54685 2226
rect 54565 2159 54590 2209
rect 54400 1535 54420 1865
rect 54735 1945 54755 2280
rect 54905 2095 54925 2230
rect 54960 2355 54990 2365
rect 54960 2335 54965 2355
rect 54985 2335 54990 2355
rect 54960 2305 54990 2335
rect 54960 2285 54965 2305
rect 54985 2285 54990 2305
rect 54960 2255 54990 2285
rect 54960 2235 54965 2255
rect 54985 2235 54990 2255
rect 54960 2205 54990 2235
rect 54960 2185 54965 2205
rect 54985 2185 54990 2205
rect 54960 2145 54990 2185
rect 55015 2355 55045 2365
rect 55015 2335 55020 2355
rect 55040 2335 55045 2355
rect 55015 2305 55045 2335
rect 55015 2285 55020 2305
rect 55040 2285 55045 2305
rect 55015 2255 55045 2285
rect 55015 2235 55020 2255
rect 55040 2235 55045 2255
rect 55015 2205 55045 2235
rect 55015 2185 55020 2205
rect 55040 2185 55045 2205
rect 55015 2175 55045 2185
rect 55070 2355 55100 2365
rect 55070 2335 55075 2355
rect 55095 2335 55100 2355
rect 55070 2305 55100 2335
rect 55070 2285 55075 2305
rect 55095 2285 55100 2305
rect 55070 2255 55100 2285
rect 55070 2235 55075 2255
rect 55095 2235 55100 2255
rect 55070 2205 55100 2235
rect 55070 2185 55075 2205
rect 55095 2185 55100 2205
rect 55070 2175 55100 2185
rect 55125 2355 55155 2365
rect 55125 2335 55130 2355
rect 55150 2335 55155 2355
rect 55125 2305 55155 2335
rect 55125 2285 55130 2305
rect 55150 2285 55155 2305
rect 55125 2255 55155 2285
rect 55125 2235 55130 2255
rect 55150 2235 55155 2255
rect 55125 2205 55155 2235
rect 55125 2185 55130 2205
rect 55150 2185 55155 2205
rect 55125 2175 55155 2185
rect 55180 2355 55210 2365
rect 55180 2335 55185 2355
rect 55205 2335 55210 2355
rect 55180 2305 55210 2335
rect 55180 2285 55185 2305
rect 55205 2285 55210 2305
rect 55180 2255 55210 2285
rect 55180 2235 55185 2255
rect 55205 2235 55210 2255
rect 55180 2205 55210 2235
rect 55180 2185 55185 2205
rect 55205 2185 55210 2205
rect 55180 2175 55210 2185
rect 55235 2355 55265 2365
rect 55235 2335 55240 2355
rect 55260 2335 55265 2355
rect 55235 2305 55265 2335
rect 55235 2285 55240 2305
rect 55260 2285 55265 2305
rect 55235 2255 55265 2285
rect 55235 2235 55240 2255
rect 55260 2235 55265 2255
rect 55235 2205 55265 2235
rect 55235 2185 55240 2205
rect 55260 2185 55265 2205
rect 55235 2175 55265 2185
rect 55290 2355 55320 2365
rect 55290 2335 55295 2355
rect 55315 2335 55320 2355
rect 55290 2305 55320 2335
rect 55290 2285 55295 2305
rect 55315 2285 55320 2305
rect 55290 2255 55320 2285
rect 55290 2235 55295 2255
rect 55315 2235 55320 2255
rect 55290 2205 55320 2235
rect 55290 2185 55295 2205
rect 55315 2185 55320 2205
rect 55290 2175 55320 2185
rect 55345 2355 55375 2365
rect 55345 2335 55350 2355
rect 55370 2335 55375 2355
rect 55345 2305 55375 2335
rect 55345 2285 55350 2305
rect 55370 2285 55375 2305
rect 55345 2255 55375 2285
rect 55345 2235 55350 2255
rect 55370 2235 55375 2255
rect 55345 2205 55375 2235
rect 55345 2185 55350 2205
rect 55370 2185 55375 2205
rect 55345 2175 55375 2185
rect 55400 2355 55430 2365
rect 55400 2335 55405 2355
rect 55425 2335 55430 2355
rect 55400 2305 55430 2335
rect 55400 2285 55405 2305
rect 55425 2285 55430 2305
rect 55400 2255 55430 2285
rect 55400 2235 55405 2255
rect 55425 2235 55430 2255
rect 55400 2205 55430 2235
rect 55400 2185 55405 2205
rect 55425 2185 55430 2205
rect 55400 2175 55430 2185
rect 55455 2355 55485 2365
rect 55455 2335 55460 2355
rect 55480 2335 55485 2355
rect 55455 2305 55485 2335
rect 55455 2285 55460 2305
rect 55480 2285 55485 2305
rect 55455 2255 55485 2285
rect 55455 2235 55460 2255
rect 55480 2235 55485 2255
rect 55455 2205 55485 2235
rect 55455 2185 55460 2205
rect 55480 2185 55485 2205
rect 55455 2175 55485 2185
rect 55510 2355 55540 2365
rect 55510 2335 55515 2355
rect 55535 2335 55540 2355
rect 55510 2305 55540 2335
rect 55510 2285 55515 2305
rect 55535 2285 55540 2305
rect 55510 2255 55540 2285
rect 55510 2235 55515 2255
rect 55535 2235 55540 2255
rect 55510 2205 55540 2235
rect 55510 2185 55515 2205
rect 55535 2185 55540 2205
rect 55510 2175 55540 2185
rect 55565 2355 55595 2365
rect 55565 2335 55570 2355
rect 55590 2335 55595 2355
rect 55565 2305 55595 2335
rect 55565 2285 55570 2305
rect 55590 2285 55595 2305
rect 55565 2255 55595 2285
rect 55565 2235 55570 2255
rect 55590 2235 55595 2255
rect 55565 2205 55595 2235
rect 55565 2185 55570 2205
rect 55590 2185 55595 2205
rect 55565 2175 55595 2185
rect 55620 2355 55650 2365
rect 55620 2335 55625 2355
rect 55645 2335 55650 2355
rect 55620 2305 55650 2335
rect 55620 2285 55625 2305
rect 55645 2285 55650 2305
rect 55620 2255 55650 2285
rect 55620 2235 55625 2255
rect 55645 2235 55650 2255
rect 55620 2205 55650 2235
rect 55620 2185 55625 2205
rect 55645 2185 55650 2205
rect 55075 2155 55095 2175
rect 55185 2155 55205 2175
rect 55295 2155 55315 2175
rect 55405 2155 55425 2175
rect 55515 2155 55535 2175
rect 54960 2125 54965 2145
rect 54985 2125 54990 2145
rect 54960 2115 54990 2125
rect 55065 2145 55105 2155
rect 55065 2125 55075 2145
rect 55095 2125 55105 2145
rect 55065 2115 55105 2125
rect 55175 2145 55215 2155
rect 55175 2125 55185 2145
rect 55205 2125 55215 2145
rect 55175 2115 55215 2125
rect 55285 2145 55325 2155
rect 55285 2125 55295 2145
rect 55315 2125 55325 2145
rect 55285 2115 55325 2125
rect 55395 2145 55435 2155
rect 55395 2125 55405 2145
rect 55425 2125 55435 2145
rect 55395 2115 55435 2125
rect 55453 2145 55487 2155
rect 55453 2125 55461 2145
rect 55479 2125 55487 2145
rect 55453 2115 55487 2125
rect 55505 2145 55545 2155
rect 55505 2125 55515 2145
rect 55535 2125 55545 2145
rect 55505 2115 55545 2125
rect 55620 2145 55650 2185
rect 55620 2125 55625 2145
rect 55645 2125 55650 2145
rect 55620 2115 55650 2125
rect 55685 2310 55705 2445
rect 56555 2505 56585 2515
rect 56555 2485 56560 2505
rect 56580 2485 56585 2505
rect 56555 2445 56585 2485
rect 56605 2505 56645 2515
rect 56605 2485 56615 2505
rect 56635 2485 56645 2505
rect 56605 2475 56645 2485
rect 56715 2505 56755 2515
rect 56715 2485 56725 2505
rect 56745 2485 56755 2505
rect 56715 2475 56755 2485
rect 56825 2505 56865 2515
rect 56825 2485 56835 2505
rect 56855 2485 56865 2505
rect 56825 2475 56865 2485
rect 56935 2505 56975 2515
rect 56935 2485 56945 2505
rect 56965 2485 56975 2505
rect 56935 2475 56975 2485
rect 57045 2505 57085 2515
rect 57045 2485 57055 2505
rect 57075 2485 57085 2505
rect 57045 2475 57085 2485
rect 57155 2505 57195 2515
rect 57155 2485 57165 2505
rect 57185 2485 57195 2505
rect 57155 2475 57195 2485
rect 57215 2505 57245 2515
rect 57215 2485 57220 2505
rect 57240 2485 57245 2505
rect 56615 2455 56635 2475
rect 56725 2455 56745 2475
rect 56835 2455 56855 2475
rect 56945 2455 56965 2475
rect 57055 2455 57075 2475
rect 57165 2455 57185 2475
rect 56555 2425 56560 2445
rect 56580 2425 56585 2445
rect 56555 2415 56585 2425
rect 56610 2445 56640 2455
rect 56610 2425 56615 2445
rect 56635 2425 56640 2445
rect 56610 2415 56640 2425
rect 56665 2445 56695 2455
rect 56665 2425 56670 2445
rect 56690 2425 56695 2445
rect 56665 2415 56695 2425
rect 56720 2445 56750 2455
rect 56720 2425 56725 2445
rect 56745 2425 56750 2445
rect 56720 2415 56750 2425
rect 56775 2445 56805 2455
rect 56775 2425 56780 2445
rect 56800 2425 56805 2445
rect 56775 2415 56805 2425
rect 56830 2445 56860 2455
rect 56830 2425 56835 2445
rect 56855 2425 56860 2445
rect 56830 2415 56860 2425
rect 56885 2445 56915 2455
rect 56885 2425 56890 2445
rect 56910 2425 56915 2445
rect 56885 2415 56915 2425
rect 56940 2445 56970 2455
rect 56940 2425 56945 2445
rect 56965 2425 56970 2445
rect 56940 2415 56970 2425
rect 56995 2445 57025 2455
rect 56995 2425 57000 2445
rect 57020 2425 57025 2445
rect 56995 2415 57025 2425
rect 57050 2445 57080 2455
rect 57050 2425 57055 2445
rect 57075 2425 57080 2445
rect 57050 2415 57080 2425
rect 57105 2445 57135 2455
rect 57105 2425 57110 2445
rect 57130 2425 57135 2445
rect 57105 2415 57135 2425
rect 57160 2445 57190 2455
rect 57160 2425 57165 2445
rect 57185 2425 57190 2445
rect 57160 2415 57190 2425
rect 57215 2445 57245 2485
rect 57215 2425 57220 2445
rect 57240 2425 57245 2445
rect 57215 2415 57245 2425
rect 57280 2465 57300 2535
rect 58475 2475 58515 2485
rect 58475 2465 58485 2475
rect 58505 2465 58515 2475
rect 56670 2395 56690 2415
rect 56780 2395 56800 2415
rect 56890 2395 56910 2415
rect 57000 2395 57020 2415
rect 57110 2395 57130 2415
rect 56500 2335 56520 2385
rect 56660 2385 56700 2395
rect 56660 2365 56670 2385
rect 56690 2365 56700 2385
rect 56660 2355 56700 2365
rect 56770 2385 56810 2395
rect 56770 2365 56780 2385
rect 56800 2365 56810 2385
rect 56770 2355 56810 2365
rect 56880 2385 56920 2395
rect 56880 2365 56890 2385
rect 56910 2365 56920 2385
rect 56880 2355 56920 2365
rect 56990 2385 57030 2395
rect 56990 2365 57000 2385
rect 57020 2365 57030 2385
rect 56990 2355 57030 2365
rect 57100 2385 57140 2395
rect 57100 2365 57110 2385
rect 57130 2365 57140 2385
rect 57100 2355 57140 2365
rect 57280 2335 57300 2385
rect 56500 2315 56860 2335
rect 56940 2315 57300 2335
rect 58095 2445 58455 2465
rect 58535 2445 58895 2465
rect 56880 2305 56890 2315
rect 56910 2305 56920 2315
rect 56880 2295 56920 2305
rect 58095 2310 58115 2445
rect 58200 2415 58240 2425
rect 58200 2395 58210 2415
rect 58230 2395 58240 2415
rect 58200 2385 58240 2395
rect 58310 2415 58350 2425
rect 58310 2395 58320 2415
rect 58340 2395 58350 2415
rect 58310 2385 58350 2395
rect 58420 2415 58460 2425
rect 58420 2395 58430 2415
rect 58450 2395 58460 2415
rect 58420 2385 58460 2395
rect 58530 2415 58570 2425
rect 58530 2395 58540 2415
rect 58560 2395 58570 2415
rect 58530 2385 58570 2395
rect 58640 2415 58680 2425
rect 58640 2395 58650 2415
rect 58670 2395 58680 2415
rect 58640 2385 58680 2395
rect 58750 2415 58790 2425
rect 58750 2395 58760 2415
rect 58780 2395 58790 2415
rect 58750 2385 58790 2395
rect 58210 2365 58230 2385
rect 58320 2365 58340 2385
rect 58430 2365 58450 2385
rect 58540 2365 58560 2385
rect 58650 2365 58670 2385
rect 58760 2365 58780 2385
rect 54965 2095 54985 2115
rect 55625 2095 55645 2115
rect 55685 2095 55705 2230
rect 54905 2075 55265 2095
rect 55345 2075 55705 2095
rect 56025 2255 56825 2275
rect 56025 2145 56045 2255
rect 56085 2235 56105 2255
rect 56745 2235 56765 2255
rect 54470 1590 54505 1600
rect 54470 1565 54475 1590
rect 54500 1565 54505 1590
rect 54470 1555 54505 1565
rect 54530 1590 54565 1600
rect 54530 1565 54535 1590
rect 54560 1565 54565 1590
rect 54530 1555 54565 1565
rect 54590 1590 54625 1600
rect 54590 1565 54595 1590
rect 54620 1565 54625 1590
rect 54590 1555 54625 1565
rect 54650 1590 54685 1600
rect 54650 1565 54655 1590
rect 54680 1565 54685 1590
rect 54650 1555 54685 1565
rect 54735 1780 54755 1865
rect 54905 1985 55265 2005
rect 55345 1985 55705 2005
rect 54905 1800 54925 1985
rect 54965 1965 54985 1985
rect 55625 1965 55645 1985
rect 54735 1770 54775 1780
rect 54735 1750 54745 1770
rect 54765 1750 54775 1770
rect 54735 1740 54775 1750
rect 54885 1770 54905 1780
rect 54885 1750 54895 1770
rect 54885 1740 54905 1750
rect 54735 1535 54755 1740
rect 54400 1515 54535 1535
rect 54615 1515 54755 1535
rect 54905 1535 54925 1720
rect 54960 1955 54990 1965
rect 54960 1935 54965 1955
rect 54985 1935 54990 1955
rect 54960 1895 54990 1935
rect 55065 1955 55105 1965
rect 55065 1935 55075 1955
rect 55095 1935 55105 1955
rect 55065 1925 55105 1935
rect 55175 1955 55215 1965
rect 55175 1935 55185 1955
rect 55205 1935 55215 1955
rect 55175 1925 55215 1935
rect 55285 1955 55325 1965
rect 55285 1935 55295 1955
rect 55315 1935 55325 1955
rect 55285 1925 55325 1935
rect 55395 1955 55435 1965
rect 55395 1935 55405 1955
rect 55425 1935 55435 1955
rect 55395 1925 55435 1935
rect 55453 1955 55487 1965
rect 55453 1935 55461 1955
rect 55479 1935 55487 1955
rect 55453 1925 55487 1935
rect 55505 1955 55545 1965
rect 55505 1935 55515 1955
rect 55535 1935 55545 1955
rect 55505 1925 55545 1935
rect 55620 1955 55650 1965
rect 55620 1935 55625 1955
rect 55645 1935 55650 1955
rect 55075 1905 55095 1925
rect 55185 1905 55205 1925
rect 55295 1905 55315 1925
rect 55405 1905 55425 1925
rect 55515 1905 55535 1925
rect 54960 1875 54965 1895
rect 54985 1875 54990 1895
rect 54960 1845 54990 1875
rect 54960 1825 54965 1845
rect 54985 1825 54990 1845
rect 54960 1795 54990 1825
rect 54960 1775 54965 1795
rect 54985 1775 54990 1795
rect 54960 1745 54990 1775
rect 54960 1725 54965 1745
rect 54985 1725 54990 1745
rect 54960 1695 54990 1725
rect 54960 1675 54965 1695
rect 54985 1675 54990 1695
rect 54960 1645 54990 1675
rect 54960 1625 54965 1645
rect 54985 1625 54990 1645
rect 54960 1615 54990 1625
rect 55015 1895 55045 1905
rect 55015 1875 55020 1895
rect 55040 1875 55045 1895
rect 55015 1845 55045 1875
rect 55015 1825 55020 1845
rect 55040 1825 55045 1845
rect 55015 1795 55045 1825
rect 55015 1775 55020 1795
rect 55040 1775 55045 1795
rect 55015 1745 55045 1775
rect 55015 1725 55020 1745
rect 55040 1725 55045 1745
rect 55015 1695 55045 1725
rect 55015 1675 55020 1695
rect 55040 1675 55045 1695
rect 55015 1645 55045 1675
rect 55015 1625 55020 1645
rect 55040 1625 55045 1645
rect 55015 1615 55045 1625
rect 55070 1895 55100 1905
rect 55070 1875 55075 1895
rect 55095 1875 55100 1895
rect 55070 1845 55100 1875
rect 55070 1825 55075 1845
rect 55095 1825 55100 1845
rect 55070 1795 55100 1825
rect 55070 1775 55075 1795
rect 55095 1775 55100 1795
rect 55070 1745 55100 1775
rect 55070 1725 55075 1745
rect 55095 1725 55100 1745
rect 55070 1695 55100 1725
rect 55070 1675 55075 1695
rect 55095 1675 55100 1695
rect 55070 1645 55100 1675
rect 55070 1625 55075 1645
rect 55095 1625 55100 1645
rect 55070 1615 55100 1625
rect 55125 1895 55155 1905
rect 55125 1875 55130 1895
rect 55150 1875 55155 1895
rect 55125 1845 55155 1875
rect 55125 1825 55130 1845
rect 55150 1825 55155 1845
rect 55125 1795 55155 1825
rect 55125 1775 55130 1795
rect 55150 1775 55155 1795
rect 55125 1745 55155 1775
rect 55125 1725 55130 1745
rect 55150 1725 55155 1745
rect 55125 1695 55155 1725
rect 55125 1675 55130 1695
rect 55150 1675 55155 1695
rect 55125 1645 55155 1675
rect 55125 1625 55130 1645
rect 55150 1625 55155 1645
rect 55125 1615 55155 1625
rect 55180 1895 55210 1905
rect 55180 1875 55185 1895
rect 55205 1875 55210 1895
rect 55180 1845 55210 1875
rect 55180 1825 55185 1845
rect 55205 1825 55210 1845
rect 55180 1795 55210 1825
rect 55180 1775 55185 1795
rect 55205 1775 55210 1795
rect 55180 1745 55210 1775
rect 55180 1725 55185 1745
rect 55205 1725 55210 1745
rect 55180 1695 55210 1725
rect 55180 1675 55185 1695
rect 55205 1675 55210 1695
rect 55180 1645 55210 1675
rect 55180 1625 55185 1645
rect 55205 1625 55210 1645
rect 55180 1615 55210 1625
rect 55235 1895 55265 1905
rect 55235 1875 55240 1895
rect 55260 1875 55265 1895
rect 55235 1845 55265 1875
rect 55235 1825 55240 1845
rect 55260 1825 55265 1845
rect 55235 1795 55265 1825
rect 55235 1775 55240 1795
rect 55260 1775 55265 1795
rect 55235 1745 55265 1775
rect 55235 1725 55240 1745
rect 55260 1725 55265 1745
rect 55235 1695 55265 1725
rect 55235 1675 55240 1695
rect 55260 1675 55265 1695
rect 55235 1645 55265 1675
rect 55235 1625 55240 1645
rect 55260 1625 55265 1645
rect 55235 1615 55265 1625
rect 55290 1895 55320 1905
rect 55290 1875 55295 1895
rect 55315 1875 55320 1895
rect 55290 1845 55320 1875
rect 55290 1825 55295 1845
rect 55315 1825 55320 1845
rect 55290 1795 55320 1825
rect 55290 1775 55295 1795
rect 55315 1775 55320 1795
rect 55290 1745 55320 1775
rect 55290 1725 55295 1745
rect 55315 1725 55320 1745
rect 55290 1695 55320 1725
rect 55290 1675 55295 1695
rect 55315 1675 55320 1695
rect 55290 1645 55320 1675
rect 55290 1625 55295 1645
rect 55315 1625 55320 1645
rect 55290 1615 55320 1625
rect 55345 1895 55375 1905
rect 55345 1875 55350 1895
rect 55370 1875 55375 1895
rect 55345 1845 55375 1875
rect 55345 1825 55350 1845
rect 55370 1825 55375 1845
rect 55345 1795 55375 1825
rect 55345 1775 55350 1795
rect 55370 1775 55375 1795
rect 55345 1745 55375 1775
rect 55345 1725 55350 1745
rect 55370 1725 55375 1745
rect 55345 1695 55375 1725
rect 55345 1675 55350 1695
rect 55370 1675 55375 1695
rect 55345 1645 55375 1675
rect 55345 1625 55350 1645
rect 55370 1625 55375 1645
rect 55345 1615 55375 1625
rect 55400 1895 55430 1905
rect 55400 1875 55405 1895
rect 55425 1875 55430 1895
rect 55400 1845 55430 1875
rect 55400 1825 55405 1845
rect 55425 1825 55430 1845
rect 55400 1795 55430 1825
rect 55400 1775 55405 1795
rect 55425 1775 55430 1795
rect 55400 1745 55430 1775
rect 55400 1725 55405 1745
rect 55425 1725 55430 1745
rect 55400 1695 55430 1725
rect 55400 1675 55405 1695
rect 55425 1675 55430 1695
rect 55400 1645 55430 1675
rect 55400 1625 55405 1645
rect 55425 1625 55430 1645
rect 55400 1615 55430 1625
rect 55455 1895 55485 1905
rect 55455 1875 55460 1895
rect 55480 1875 55485 1895
rect 55455 1845 55485 1875
rect 55455 1825 55460 1845
rect 55480 1825 55485 1845
rect 55455 1795 55485 1825
rect 55455 1775 55460 1795
rect 55480 1775 55485 1795
rect 55455 1745 55485 1775
rect 55455 1725 55460 1745
rect 55480 1725 55485 1745
rect 55455 1695 55485 1725
rect 55455 1675 55460 1695
rect 55480 1675 55485 1695
rect 55455 1645 55485 1675
rect 55455 1625 55460 1645
rect 55480 1625 55485 1645
rect 55455 1615 55485 1625
rect 55510 1895 55540 1905
rect 55510 1875 55515 1895
rect 55535 1875 55540 1895
rect 55510 1845 55540 1875
rect 55510 1825 55515 1845
rect 55535 1825 55540 1845
rect 55510 1795 55540 1825
rect 55510 1775 55515 1795
rect 55535 1775 55540 1795
rect 55510 1745 55540 1775
rect 55510 1725 55515 1745
rect 55535 1725 55540 1745
rect 55510 1695 55540 1725
rect 55510 1675 55515 1695
rect 55535 1675 55540 1695
rect 55510 1645 55540 1675
rect 55510 1625 55515 1645
rect 55535 1625 55540 1645
rect 55510 1615 55540 1625
rect 55565 1895 55595 1905
rect 55565 1875 55570 1895
rect 55590 1875 55595 1895
rect 55565 1845 55595 1875
rect 55565 1825 55570 1845
rect 55590 1825 55595 1845
rect 55565 1795 55595 1825
rect 55565 1775 55570 1795
rect 55590 1775 55595 1795
rect 55565 1745 55595 1775
rect 55565 1725 55570 1745
rect 55590 1725 55595 1745
rect 55565 1695 55595 1725
rect 55565 1675 55570 1695
rect 55590 1675 55595 1695
rect 55565 1645 55595 1675
rect 55565 1625 55570 1645
rect 55590 1625 55595 1645
rect 55565 1615 55595 1625
rect 55620 1895 55650 1935
rect 55620 1875 55625 1895
rect 55645 1875 55650 1895
rect 55620 1845 55650 1875
rect 55620 1825 55625 1845
rect 55645 1825 55650 1845
rect 55620 1795 55650 1825
rect 55620 1775 55625 1795
rect 55645 1775 55650 1795
rect 55620 1745 55650 1775
rect 55620 1725 55625 1745
rect 55645 1725 55650 1745
rect 55620 1695 55650 1725
rect 55620 1675 55625 1695
rect 55645 1675 55650 1695
rect 55620 1645 55650 1675
rect 55620 1625 55625 1645
rect 55645 1625 55650 1645
rect 55620 1615 55650 1625
rect 55685 1800 55705 1985
rect 56025 1955 56045 2065
rect 56080 2225 56110 2235
rect 56080 2205 56085 2225
rect 56105 2205 56110 2225
rect 56080 2165 56110 2205
rect 56130 2225 56170 2235
rect 56130 2205 56140 2225
rect 56160 2205 56170 2225
rect 56130 2195 56170 2205
rect 56240 2225 56280 2235
rect 56240 2205 56250 2225
rect 56270 2205 56280 2225
rect 56240 2195 56280 2205
rect 56350 2225 56390 2235
rect 56350 2205 56360 2225
rect 56380 2205 56390 2225
rect 56350 2195 56390 2205
rect 56410 2225 56440 2235
rect 56410 2205 56415 2225
rect 56435 2205 56440 2225
rect 56410 2195 56440 2205
rect 56460 2225 56500 2235
rect 56460 2205 56470 2225
rect 56490 2205 56500 2225
rect 56460 2195 56500 2205
rect 56570 2225 56610 2235
rect 56570 2205 56580 2225
rect 56600 2205 56610 2225
rect 56570 2195 56610 2205
rect 56680 2225 56720 2235
rect 56680 2205 56690 2225
rect 56710 2205 56720 2225
rect 56680 2195 56720 2205
rect 56740 2225 56770 2235
rect 56740 2205 56745 2225
rect 56765 2205 56770 2225
rect 56140 2175 56160 2195
rect 56250 2175 56270 2195
rect 56360 2175 56380 2195
rect 56470 2175 56490 2195
rect 56580 2175 56600 2195
rect 56690 2175 56710 2195
rect 56080 2145 56085 2165
rect 56105 2145 56110 2165
rect 56080 2115 56110 2145
rect 56080 2095 56085 2115
rect 56105 2095 56110 2115
rect 56080 2065 56110 2095
rect 56080 2045 56085 2065
rect 56105 2045 56110 2065
rect 56080 2035 56110 2045
rect 56135 2165 56165 2175
rect 56135 2145 56140 2165
rect 56160 2145 56165 2165
rect 56135 2115 56165 2145
rect 56135 2095 56140 2115
rect 56160 2095 56165 2115
rect 56135 2065 56165 2095
rect 56135 2045 56140 2065
rect 56160 2045 56165 2065
rect 56135 2035 56165 2045
rect 56190 2165 56220 2175
rect 56190 2145 56195 2165
rect 56215 2145 56220 2165
rect 56190 2115 56220 2145
rect 56190 2095 56195 2115
rect 56215 2095 56220 2115
rect 56190 2065 56220 2095
rect 56190 2045 56195 2065
rect 56215 2045 56220 2065
rect 56190 2035 56220 2045
rect 56245 2165 56275 2175
rect 56245 2145 56250 2165
rect 56270 2145 56275 2165
rect 56245 2115 56275 2145
rect 56245 2095 56250 2115
rect 56270 2095 56275 2115
rect 56245 2065 56275 2095
rect 56245 2045 56250 2065
rect 56270 2045 56275 2065
rect 56245 2035 56275 2045
rect 56300 2165 56330 2175
rect 56300 2145 56305 2165
rect 56325 2145 56330 2165
rect 56300 2115 56330 2145
rect 56300 2095 56305 2115
rect 56325 2095 56330 2115
rect 56300 2065 56330 2095
rect 56300 2045 56305 2065
rect 56325 2045 56330 2065
rect 56300 2035 56330 2045
rect 56355 2165 56385 2175
rect 56355 2145 56360 2165
rect 56380 2145 56385 2165
rect 56355 2115 56385 2145
rect 56355 2095 56360 2115
rect 56380 2095 56385 2115
rect 56355 2065 56385 2095
rect 56355 2045 56360 2065
rect 56380 2045 56385 2065
rect 56355 2035 56385 2045
rect 56410 2165 56440 2175
rect 56410 2145 56415 2165
rect 56435 2145 56440 2165
rect 56410 2115 56440 2145
rect 56410 2095 56415 2115
rect 56435 2095 56440 2115
rect 56410 2065 56440 2095
rect 56410 2045 56415 2065
rect 56435 2045 56440 2065
rect 56410 2035 56440 2045
rect 56465 2165 56495 2175
rect 56465 2145 56470 2165
rect 56490 2145 56495 2165
rect 56465 2115 56495 2145
rect 56465 2095 56470 2115
rect 56490 2095 56495 2115
rect 56465 2065 56495 2095
rect 56465 2045 56470 2065
rect 56490 2045 56495 2065
rect 56465 2035 56495 2045
rect 56520 2165 56550 2175
rect 56520 2145 56525 2165
rect 56545 2145 56550 2165
rect 56520 2115 56550 2145
rect 56520 2095 56525 2115
rect 56545 2095 56550 2115
rect 56520 2065 56550 2095
rect 56520 2045 56525 2065
rect 56545 2045 56550 2065
rect 56520 2035 56550 2045
rect 56575 2165 56605 2175
rect 56575 2145 56580 2165
rect 56600 2145 56605 2165
rect 56575 2115 56605 2145
rect 56575 2095 56580 2115
rect 56600 2095 56605 2115
rect 56575 2065 56605 2095
rect 56575 2045 56580 2065
rect 56600 2045 56605 2065
rect 56575 2035 56605 2045
rect 56630 2165 56660 2175
rect 56630 2145 56635 2165
rect 56655 2145 56660 2165
rect 56630 2115 56660 2145
rect 56630 2095 56635 2115
rect 56655 2095 56660 2115
rect 56630 2065 56660 2095
rect 56630 2045 56635 2065
rect 56655 2045 56660 2065
rect 56630 2035 56660 2045
rect 56685 2165 56715 2175
rect 56685 2145 56690 2165
rect 56710 2145 56715 2165
rect 56685 2115 56715 2145
rect 56685 2095 56690 2115
rect 56710 2095 56715 2115
rect 56685 2065 56715 2095
rect 56685 2045 56690 2065
rect 56710 2045 56715 2065
rect 56685 2035 56715 2045
rect 56740 2165 56770 2205
rect 56740 2145 56745 2165
rect 56765 2145 56770 2165
rect 56740 2115 56770 2145
rect 56740 2095 56745 2115
rect 56765 2095 56770 2115
rect 56740 2065 56770 2095
rect 56740 2045 56745 2065
rect 56765 2045 56770 2065
rect 56740 2035 56770 2045
rect 56805 2145 56825 2255
rect 56195 2015 56215 2035
rect 56305 2015 56325 2035
rect 56415 2015 56435 2035
rect 56525 2015 56545 2035
rect 56635 2015 56655 2035
rect 56185 2005 56225 2015
rect 56185 1985 56195 2005
rect 56215 1985 56225 2005
rect 56185 1975 56225 1985
rect 56295 2005 56335 2015
rect 56295 1985 56305 2005
rect 56325 1985 56335 2005
rect 56295 1975 56335 1985
rect 56405 2005 56445 2015
rect 56405 1985 56415 2005
rect 56435 1985 56445 2005
rect 56405 1975 56445 1985
rect 56515 2005 56555 2015
rect 56515 1985 56525 2005
rect 56545 1985 56555 2005
rect 56515 1975 56555 1985
rect 56625 2005 56665 2015
rect 56625 1985 56635 2005
rect 56655 1985 56665 2005
rect 56625 1975 56665 1985
rect 56805 1955 56825 2065
rect 56025 1935 56825 1955
rect 56975 2255 57775 2275
rect 56975 2145 56995 2255
rect 57035 2235 57055 2255
rect 57695 2235 57715 2255
rect 56975 1955 56995 2065
rect 57030 2225 57060 2235
rect 57030 2205 57035 2225
rect 57055 2205 57060 2225
rect 57030 2165 57060 2205
rect 57080 2225 57120 2235
rect 57080 2205 57090 2225
rect 57110 2205 57120 2225
rect 57080 2195 57120 2205
rect 57190 2225 57230 2235
rect 57190 2205 57200 2225
rect 57220 2205 57230 2225
rect 57190 2195 57230 2205
rect 57300 2225 57340 2235
rect 57300 2205 57310 2225
rect 57330 2205 57340 2225
rect 57300 2195 57340 2205
rect 57360 2225 57390 2235
rect 57360 2205 57365 2225
rect 57385 2205 57390 2225
rect 57360 2195 57390 2205
rect 57410 2225 57450 2235
rect 57410 2205 57420 2225
rect 57440 2205 57450 2225
rect 57410 2195 57450 2205
rect 57520 2225 57560 2235
rect 57520 2205 57530 2225
rect 57550 2205 57560 2225
rect 57520 2195 57560 2205
rect 57630 2225 57670 2235
rect 57630 2205 57640 2225
rect 57660 2205 57670 2225
rect 57630 2195 57670 2205
rect 57690 2225 57720 2235
rect 57690 2205 57695 2225
rect 57715 2205 57720 2225
rect 57090 2175 57110 2195
rect 57200 2175 57220 2195
rect 57310 2175 57330 2195
rect 57420 2175 57440 2195
rect 57530 2175 57550 2195
rect 57640 2175 57660 2195
rect 57030 2145 57035 2165
rect 57055 2145 57060 2165
rect 57030 2115 57060 2145
rect 57030 2095 57035 2115
rect 57055 2095 57060 2115
rect 57030 2065 57060 2095
rect 57030 2045 57035 2065
rect 57055 2045 57060 2065
rect 57030 2035 57060 2045
rect 57085 2165 57115 2175
rect 57085 2145 57090 2165
rect 57110 2145 57115 2165
rect 57085 2115 57115 2145
rect 57085 2095 57090 2115
rect 57110 2095 57115 2115
rect 57085 2065 57115 2095
rect 57085 2045 57090 2065
rect 57110 2045 57115 2065
rect 57085 2035 57115 2045
rect 57140 2165 57170 2175
rect 57140 2145 57145 2165
rect 57165 2145 57170 2165
rect 57140 2115 57170 2145
rect 57140 2095 57145 2115
rect 57165 2095 57170 2115
rect 57140 2065 57170 2095
rect 57140 2045 57145 2065
rect 57165 2045 57170 2065
rect 57140 2035 57170 2045
rect 57195 2165 57225 2175
rect 57195 2145 57200 2165
rect 57220 2145 57225 2165
rect 57195 2115 57225 2145
rect 57195 2095 57200 2115
rect 57220 2095 57225 2115
rect 57195 2065 57225 2095
rect 57195 2045 57200 2065
rect 57220 2045 57225 2065
rect 57195 2035 57225 2045
rect 57250 2165 57280 2175
rect 57250 2145 57255 2165
rect 57275 2145 57280 2165
rect 57250 2115 57280 2145
rect 57250 2095 57255 2115
rect 57275 2095 57280 2115
rect 57250 2065 57280 2095
rect 57250 2045 57255 2065
rect 57275 2045 57280 2065
rect 57250 2035 57280 2045
rect 57305 2165 57335 2175
rect 57305 2145 57310 2165
rect 57330 2145 57335 2165
rect 57305 2115 57335 2145
rect 57305 2095 57310 2115
rect 57330 2095 57335 2115
rect 57305 2065 57335 2095
rect 57305 2045 57310 2065
rect 57330 2045 57335 2065
rect 57305 2035 57335 2045
rect 57360 2165 57390 2175
rect 57360 2145 57365 2165
rect 57385 2145 57390 2165
rect 57360 2115 57390 2145
rect 57360 2095 57365 2115
rect 57385 2095 57390 2115
rect 57360 2065 57390 2095
rect 57360 2045 57365 2065
rect 57385 2045 57390 2065
rect 57360 2035 57390 2045
rect 57415 2165 57445 2175
rect 57415 2145 57420 2165
rect 57440 2145 57445 2165
rect 57415 2115 57445 2145
rect 57415 2095 57420 2115
rect 57440 2095 57445 2115
rect 57415 2065 57445 2095
rect 57415 2045 57420 2065
rect 57440 2045 57445 2065
rect 57415 2035 57445 2045
rect 57470 2165 57500 2175
rect 57470 2145 57475 2165
rect 57495 2145 57500 2165
rect 57470 2115 57500 2145
rect 57470 2095 57475 2115
rect 57495 2095 57500 2115
rect 57470 2065 57500 2095
rect 57470 2045 57475 2065
rect 57495 2045 57500 2065
rect 57470 2035 57500 2045
rect 57525 2165 57555 2175
rect 57525 2145 57530 2165
rect 57550 2145 57555 2165
rect 57525 2115 57555 2145
rect 57525 2095 57530 2115
rect 57550 2095 57555 2115
rect 57525 2065 57555 2095
rect 57525 2045 57530 2065
rect 57550 2045 57555 2065
rect 57525 2035 57555 2045
rect 57580 2165 57610 2175
rect 57580 2145 57585 2165
rect 57605 2145 57610 2165
rect 57580 2115 57610 2145
rect 57580 2095 57585 2115
rect 57605 2095 57610 2115
rect 57580 2065 57610 2095
rect 57580 2045 57585 2065
rect 57605 2045 57610 2065
rect 57580 2035 57610 2045
rect 57635 2165 57665 2175
rect 57635 2145 57640 2165
rect 57660 2145 57665 2165
rect 57635 2115 57665 2145
rect 57635 2095 57640 2115
rect 57660 2095 57665 2115
rect 57635 2065 57665 2095
rect 57635 2045 57640 2065
rect 57660 2045 57665 2065
rect 57635 2035 57665 2045
rect 57690 2165 57720 2205
rect 57690 2145 57695 2165
rect 57715 2145 57720 2165
rect 57690 2115 57720 2145
rect 57690 2095 57695 2115
rect 57715 2095 57720 2115
rect 57690 2065 57720 2095
rect 57690 2045 57695 2065
rect 57715 2045 57720 2065
rect 57690 2035 57720 2045
rect 57755 2145 57775 2255
rect 58095 2095 58115 2230
rect 58150 2355 58180 2365
rect 58150 2335 58155 2355
rect 58175 2335 58180 2355
rect 58150 2305 58180 2335
rect 58150 2285 58155 2305
rect 58175 2285 58180 2305
rect 58150 2255 58180 2285
rect 58150 2235 58155 2255
rect 58175 2235 58180 2255
rect 58150 2205 58180 2235
rect 58150 2185 58155 2205
rect 58175 2185 58180 2205
rect 58150 2145 58180 2185
rect 58205 2355 58235 2365
rect 58205 2335 58210 2355
rect 58230 2335 58235 2355
rect 58205 2305 58235 2335
rect 58205 2285 58210 2305
rect 58230 2285 58235 2305
rect 58205 2255 58235 2285
rect 58205 2235 58210 2255
rect 58230 2235 58235 2255
rect 58205 2205 58235 2235
rect 58205 2185 58210 2205
rect 58230 2185 58235 2205
rect 58205 2175 58235 2185
rect 58260 2355 58290 2365
rect 58260 2335 58265 2355
rect 58285 2335 58290 2355
rect 58260 2305 58290 2335
rect 58260 2285 58265 2305
rect 58285 2285 58290 2305
rect 58260 2255 58290 2285
rect 58260 2235 58265 2255
rect 58285 2235 58290 2255
rect 58260 2205 58290 2235
rect 58260 2185 58265 2205
rect 58285 2185 58290 2205
rect 58260 2175 58290 2185
rect 58315 2355 58345 2365
rect 58315 2335 58320 2355
rect 58340 2335 58345 2355
rect 58315 2305 58345 2335
rect 58315 2285 58320 2305
rect 58340 2285 58345 2305
rect 58315 2255 58345 2285
rect 58315 2235 58320 2255
rect 58340 2235 58345 2255
rect 58315 2205 58345 2235
rect 58315 2185 58320 2205
rect 58340 2185 58345 2205
rect 58315 2175 58345 2185
rect 58370 2355 58400 2365
rect 58370 2335 58375 2355
rect 58395 2335 58400 2355
rect 58370 2305 58400 2335
rect 58370 2285 58375 2305
rect 58395 2285 58400 2305
rect 58370 2255 58400 2285
rect 58370 2235 58375 2255
rect 58395 2235 58400 2255
rect 58370 2205 58400 2235
rect 58370 2185 58375 2205
rect 58395 2185 58400 2205
rect 58370 2175 58400 2185
rect 58425 2355 58455 2365
rect 58425 2335 58430 2355
rect 58450 2335 58455 2355
rect 58425 2305 58455 2335
rect 58425 2285 58430 2305
rect 58450 2285 58455 2305
rect 58425 2255 58455 2285
rect 58425 2235 58430 2255
rect 58450 2235 58455 2255
rect 58425 2205 58455 2235
rect 58425 2185 58430 2205
rect 58450 2185 58455 2205
rect 58425 2175 58455 2185
rect 58480 2355 58510 2365
rect 58480 2335 58485 2355
rect 58505 2335 58510 2355
rect 58480 2305 58510 2335
rect 58480 2285 58485 2305
rect 58505 2285 58510 2305
rect 58480 2255 58510 2285
rect 58480 2235 58485 2255
rect 58505 2235 58510 2255
rect 58480 2205 58510 2235
rect 58480 2185 58485 2205
rect 58505 2185 58510 2205
rect 58480 2175 58510 2185
rect 58535 2355 58565 2365
rect 58535 2335 58540 2355
rect 58560 2335 58565 2355
rect 58535 2305 58565 2335
rect 58535 2285 58540 2305
rect 58560 2285 58565 2305
rect 58535 2255 58565 2285
rect 58535 2235 58540 2255
rect 58560 2235 58565 2255
rect 58535 2205 58565 2235
rect 58535 2185 58540 2205
rect 58560 2185 58565 2205
rect 58535 2175 58565 2185
rect 58590 2355 58620 2365
rect 58590 2335 58595 2355
rect 58615 2335 58620 2355
rect 58590 2305 58620 2335
rect 58590 2285 58595 2305
rect 58615 2285 58620 2305
rect 58590 2255 58620 2285
rect 58590 2235 58595 2255
rect 58615 2235 58620 2255
rect 58590 2205 58620 2235
rect 58590 2185 58595 2205
rect 58615 2185 58620 2205
rect 58590 2175 58620 2185
rect 58645 2355 58675 2365
rect 58645 2335 58650 2355
rect 58670 2335 58675 2355
rect 58645 2305 58675 2335
rect 58645 2285 58650 2305
rect 58670 2285 58675 2305
rect 58645 2255 58675 2285
rect 58645 2235 58650 2255
rect 58670 2235 58675 2255
rect 58645 2205 58675 2235
rect 58645 2185 58650 2205
rect 58670 2185 58675 2205
rect 58645 2175 58675 2185
rect 58700 2355 58730 2365
rect 58700 2335 58705 2355
rect 58725 2335 58730 2355
rect 58700 2305 58730 2335
rect 58700 2285 58705 2305
rect 58725 2285 58730 2305
rect 58700 2255 58730 2285
rect 58700 2235 58705 2255
rect 58725 2235 58730 2255
rect 58700 2205 58730 2235
rect 58700 2185 58705 2205
rect 58725 2185 58730 2205
rect 58700 2175 58730 2185
rect 58755 2355 58785 2365
rect 58755 2335 58760 2355
rect 58780 2335 58785 2355
rect 58755 2305 58785 2335
rect 58755 2285 58760 2305
rect 58780 2285 58785 2305
rect 58755 2255 58785 2285
rect 58755 2235 58760 2255
rect 58780 2235 58785 2255
rect 58755 2205 58785 2235
rect 58755 2185 58760 2205
rect 58780 2185 58785 2205
rect 58755 2175 58785 2185
rect 58810 2355 58840 2365
rect 58810 2335 58815 2355
rect 58835 2335 58840 2355
rect 58810 2305 58840 2335
rect 58810 2285 58815 2305
rect 58835 2285 58840 2305
rect 58810 2255 58840 2285
rect 58810 2235 58815 2255
rect 58835 2235 58840 2255
rect 58810 2205 58840 2235
rect 58810 2185 58815 2205
rect 58835 2185 58840 2205
rect 58265 2155 58285 2175
rect 58375 2155 58395 2175
rect 58485 2155 58505 2175
rect 58595 2155 58615 2175
rect 58705 2155 58725 2175
rect 58150 2125 58155 2145
rect 58175 2125 58180 2145
rect 58150 2115 58180 2125
rect 58255 2145 58295 2155
rect 58255 2125 58265 2145
rect 58285 2125 58295 2145
rect 58255 2115 58295 2125
rect 58313 2145 58347 2155
rect 58313 2125 58321 2145
rect 58339 2125 58347 2145
rect 58313 2115 58347 2125
rect 58365 2145 58405 2155
rect 58365 2125 58375 2145
rect 58395 2125 58405 2145
rect 58365 2115 58405 2125
rect 58475 2145 58515 2155
rect 58475 2125 58485 2145
rect 58505 2125 58515 2145
rect 58475 2115 58515 2125
rect 58585 2145 58625 2155
rect 58585 2125 58595 2145
rect 58615 2125 58625 2145
rect 58585 2115 58625 2125
rect 58695 2145 58735 2155
rect 58695 2125 58705 2145
rect 58725 2125 58735 2145
rect 58695 2115 58735 2125
rect 58810 2145 58840 2185
rect 58810 2125 58815 2145
rect 58835 2125 58840 2145
rect 58810 2115 58840 2125
rect 58875 2310 58895 2445
rect 59235 2310 59275 2320
rect 59235 2300 59245 2310
rect 59265 2300 59275 2310
rect 58155 2095 58175 2115
rect 58815 2095 58835 2115
rect 58875 2095 58895 2230
rect 58095 2075 58455 2095
rect 58535 2075 58895 2095
rect 59045 2280 59185 2300
rect 59265 2280 59400 2300
rect 57145 2015 57165 2035
rect 57255 2015 57275 2035
rect 57365 2015 57385 2035
rect 57475 2015 57495 2035
rect 57585 2015 57605 2035
rect 57135 2005 57175 2015
rect 57135 1985 57145 2005
rect 57165 1985 57175 2005
rect 57135 1975 57175 1985
rect 57245 2005 57285 2015
rect 57245 1985 57255 2005
rect 57275 1985 57285 2005
rect 57245 1975 57285 1985
rect 57355 2005 57395 2015
rect 57355 1985 57365 2005
rect 57385 1985 57395 2005
rect 57355 1975 57395 1985
rect 57465 2005 57505 2015
rect 57465 1985 57475 2005
rect 57495 1985 57505 2005
rect 57465 1975 57505 1985
rect 57575 2005 57615 2015
rect 57575 1985 57585 2005
rect 57605 1985 57615 2005
rect 57575 1975 57615 1985
rect 57755 1955 57775 2065
rect 56975 1935 57775 1955
rect 58095 1985 58455 2005
rect 58535 1985 58895 2005
rect 56880 1815 56920 1825
rect 56880 1805 56890 1815
rect 56910 1805 56920 1815
rect 55020 1595 55040 1615
rect 55130 1595 55150 1615
rect 55240 1595 55260 1615
rect 55350 1595 55370 1615
rect 55460 1595 55480 1615
rect 55570 1595 55590 1615
rect 55010 1585 55050 1595
rect 55010 1565 55020 1585
rect 55038 1565 55050 1585
rect 55010 1555 55050 1565
rect 55120 1585 55160 1595
rect 55120 1565 55130 1585
rect 55148 1565 55160 1585
rect 55120 1555 55160 1565
rect 55230 1585 55270 1595
rect 55230 1565 55240 1585
rect 55258 1565 55270 1585
rect 55230 1555 55270 1565
rect 55340 1585 55380 1595
rect 55340 1565 55350 1585
rect 55368 1565 55380 1585
rect 55340 1555 55380 1565
rect 55450 1585 55490 1595
rect 55450 1565 55460 1585
rect 55478 1565 55490 1585
rect 55450 1555 55490 1565
rect 55560 1585 55600 1595
rect 55560 1565 55570 1585
rect 55588 1565 55600 1585
rect 55560 1555 55600 1565
rect 55685 1535 55705 1720
rect 54905 1515 55265 1535
rect 55345 1515 55705 1535
rect 55980 1785 56860 1805
rect 56940 1785 57820 1805
rect 55980 1675 56000 1785
rect 56040 1765 56060 1785
rect 56700 1765 56720 1785
rect 56780 1765 56800 1785
rect 57000 1765 57020 1785
rect 57080 1765 57100 1785
rect 57740 1765 57760 1785
rect 55285 1505 55295 1515
rect 55315 1505 55325 1515
rect 55285 1495 55325 1505
rect 55980 1485 56000 1595
rect 56035 1755 56065 1765
rect 56237 1755 56269 1765
rect 56457 1755 56489 1765
rect 56601 1755 56633 1765
rect 56695 1755 56725 1765
rect 56035 1735 56040 1755
rect 56060 1735 56065 1755
rect 56035 1695 56065 1735
rect 56100 1745 56126 1755
rect 56100 1725 56103 1745
rect 56123 1725 56126 1745
rect 56100 1715 56126 1725
rect 56194 1745 56220 1755
rect 56194 1725 56197 1745
rect 56217 1725 56220 1745
rect 56237 1735 56243 1755
rect 56260 1735 56269 1755
rect 56237 1725 56269 1735
rect 56320 1745 56346 1755
rect 56320 1725 56323 1745
rect 56343 1725 56346 1745
rect 56194 1715 56220 1725
rect 56100 1705 56120 1715
rect 56200 1705 56220 1715
rect 56320 1715 56346 1725
rect 56414 1745 56440 1755
rect 56414 1725 56417 1745
rect 56437 1725 56440 1745
rect 56457 1735 56463 1755
rect 56480 1735 56489 1755
rect 56457 1725 56489 1735
rect 56540 1745 56566 1755
rect 56540 1725 56543 1745
rect 56563 1725 56566 1745
rect 56601 1735 56610 1755
rect 56627 1735 56633 1755
rect 56601 1725 56633 1735
rect 56650 1745 56676 1755
rect 56650 1725 56653 1745
rect 56673 1725 56676 1745
rect 56414 1715 56440 1725
rect 56320 1705 56340 1715
rect 56420 1705 56440 1715
rect 56540 1715 56566 1725
rect 56650 1715 56676 1725
rect 56695 1735 56700 1755
rect 56720 1735 56725 1755
rect 56540 1705 56560 1715
rect 56650 1705 56670 1715
rect 56035 1675 56040 1695
rect 56060 1675 56065 1695
rect 56035 1645 56065 1675
rect 56035 1625 56040 1645
rect 56060 1625 56065 1645
rect 56035 1595 56065 1625
rect 56035 1575 56040 1595
rect 56060 1575 56065 1595
rect 56035 1565 56065 1575
rect 56090 1695 56120 1705
rect 56090 1675 56095 1695
rect 56115 1675 56120 1695
rect 56090 1645 56120 1675
rect 56090 1625 56095 1645
rect 56115 1625 56120 1645
rect 56090 1595 56120 1625
rect 56090 1575 56095 1595
rect 56115 1575 56120 1595
rect 56090 1565 56120 1575
rect 56145 1695 56175 1705
rect 56145 1675 56150 1695
rect 56170 1675 56175 1695
rect 56145 1645 56175 1675
rect 56145 1625 56150 1645
rect 56170 1625 56175 1645
rect 56145 1595 56175 1625
rect 56145 1575 56150 1595
rect 56170 1575 56175 1595
rect 56145 1565 56175 1575
rect 56200 1695 56230 1705
rect 56200 1675 56205 1695
rect 56225 1675 56230 1695
rect 56200 1645 56230 1675
rect 56200 1625 56205 1645
rect 56225 1625 56230 1645
rect 56200 1595 56230 1625
rect 56200 1575 56205 1595
rect 56225 1575 56230 1595
rect 56200 1565 56230 1575
rect 56255 1695 56285 1705
rect 56255 1675 56260 1695
rect 56280 1675 56285 1695
rect 56255 1645 56285 1675
rect 56255 1625 56260 1645
rect 56280 1625 56285 1645
rect 56255 1595 56285 1625
rect 56255 1575 56260 1595
rect 56280 1575 56285 1595
rect 56255 1565 56285 1575
rect 56310 1695 56340 1705
rect 56310 1675 56315 1695
rect 56335 1675 56340 1695
rect 56310 1645 56340 1675
rect 56310 1625 56315 1645
rect 56335 1625 56340 1645
rect 56310 1595 56340 1625
rect 56310 1575 56315 1595
rect 56335 1575 56340 1595
rect 56310 1565 56340 1575
rect 56365 1695 56395 1705
rect 56365 1675 56370 1695
rect 56390 1675 56395 1695
rect 56365 1645 56395 1675
rect 56365 1625 56370 1645
rect 56390 1625 56395 1645
rect 56365 1595 56395 1625
rect 56365 1575 56370 1595
rect 56390 1575 56395 1595
rect 56365 1565 56395 1575
rect 56420 1695 56450 1705
rect 56420 1675 56425 1695
rect 56445 1675 56450 1695
rect 56420 1645 56450 1675
rect 56420 1625 56425 1645
rect 56445 1625 56450 1645
rect 56420 1595 56450 1625
rect 56420 1575 56425 1595
rect 56445 1575 56450 1595
rect 56420 1565 56450 1575
rect 56475 1695 56505 1705
rect 56475 1675 56480 1695
rect 56500 1675 56505 1695
rect 56475 1645 56505 1675
rect 56475 1625 56480 1645
rect 56500 1625 56505 1645
rect 56475 1595 56505 1625
rect 56475 1575 56480 1595
rect 56500 1575 56505 1595
rect 56475 1565 56505 1575
rect 56530 1695 56560 1705
rect 56530 1675 56535 1695
rect 56555 1675 56560 1695
rect 56530 1645 56560 1675
rect 56530 1625 56535 1645
rect 56555 1625 56560 1645
rect 56530 1595 56560 1625
rect 56530 1575 56535 1595
rect 56555 1575 56560 1595
rect 56530 1565 56560 1575
rect 56585 1695 56615 1705
rect 56585 1675 56590 1695
rect 56610 1675 56615 1695
rect 56585 1645 56615 1675
rect 56585 1625 56590 1645
rect 56610 1625 56615 1645
rect 56585 1595 56615 1625
rect 56585 1575 56590 1595
rect 56610 1575 56615 1595
rect 56585 1565 56615 1575
rect 56640 1695 56670 1705
rect 56640 1675 56645 1695
rect 56665 1675 56670 1695
rect 56640 1645 56670 1675
rect 56640 1625 56645 1645
rect 56665 1625 56670 1645
rect 56640 1595 56670 1625
rect 56640 1575 56645 1595
rect 56665 1575 56670 1595
rect 56640 1565 56670 1575
rect 56695 1695 56725 1735
rect 56695 1675 56700 1695
rect 56720 1675 56725 1695
rect 56695 1645 56725 1675
rect 56695 1625 56700 1645
rect 56720 1625 56725 1645
rect 56695 1595 56725 1625
rect 56695 1575 56700 1595
rect 56720 1575 56725 1595
rect 56695 1565 56725 1575
rect 56775 1755 56805 1765
rect 56775 1735 56780 1755
rect 56800 1735 56805 1755
rect 56775 1695 56805 1735
rect 56824 1755 56850 1765
rect 56824 1735 56827 1755
rect 56847 1735 56850 1755
rect 56824 1725 56850 1735
rect 56867 1755 56899 1765
rect 56867 1735 56873 1755
rect 56890 1735 56899 1755
rect 56867 1725 56899 1735
rect 56947 1755 56973 1765
rect 56947 1735 56950 1755
rect 56970 1735 56973 1755
rect 56947 1725 56973 1735
rect 56995 1755 57025 1765
rect 56995 1735 57000 1755
rect 57020 1735 57025 1755
rect 56775 1675 56780 1695
rect 56800 1675 56805 1695
rect 56775 1645 56805 1675
rect 56775 1625 56780 1645
rect 56800 1625 56805 1645
rect 56775 1595 56805 1625
rect 56775 1575 56780 1595
rect 56800 1575 56805 1595
rect 56775 1565 56805 1575
rect 56830 1705 56850 1725
rect 56950 1705 56970 1725
rect 56830 1695 56860 1705
rect 56830 1675 56835 1695
rect 56855 1675 56860 1695
rect 56830 1645 56860 1675
rect 56830 1625 56835 1645
rect 56855 1625 56860 1645
rect 56830 1595 56860 1625
rect 56830 1575 56835 1595
rect 56855 1575 56860 1595
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1675 56890 1695
rect 56910 1675 56915 1695
rect 56885 1645 56915 1675
rect 56885 1625 56890 1645
rect 56910 1625 56915 1645
rect 56885 1595 56915 1625
rect 56885 1575 56890 1595
rect 56910 1575 56915 1595
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1675 56945 1695
rect 56965 1675 56970 1695
rect 56940 1645 56970 1675
rect 56940 1625 56945 1645
rect 56965 1625 56970 1645
rect 56940 1595 56970 1625
rect 56940 1575 56945 1595
rect 56965 1575 56970 1595
rect 56940 1565 56970 1575
rect 56995 1695 57025 1735
rect 56995 1675 57000 1695
rect 57020 1675 57025 1695
rect 56995 1645 57025 1675
rect 56995 1625 57000 1645
rect 57020 1625 57025 1645
rect 56995 1595 57025 1625
rect 56995 1575 57000 1595
rect 57020 1575 57025 1595
rect 56995 1565 57025 1575
rect 57075 1755 57105 1765
rect 57277 1755 57309 1765
rect 57497 1755 57529 1765
rect 57641 1755 57673 1765
rect 57735 1755 57765 1765
rect 57075 1735 57080 1755
rect 57100 1735 57105 1755
rect 57075 1695 57105 1735
rect 57140 1745 57166 1755
rect 57140 1725 57143 1745
rect 57163 1725 57166 1745
rect 57140 1715 57166 1725
rect 57234 1745 57260 1755
rect 57234 1725 57237 1745
rect 57257 1725 57260 1745
rect 57277 1735 57283 1755
rect 57300 1735 57309 1755
rect 57277 1725 57309 1735
rect 57360 1745 57386 1755
rect 57360 1725 57363 1745
rect 57383 1725 57386 1745
rect 57234 1715 57260 1725
rect 57140 1705 57160 1715
rect 57240 1705 57260 1715
rect 57360 1715 57386 1725
rect 57454 1745 57480 1755
rect 57454 1725 57457 1745
rect 57477 1725 57480 1745
rect 57497 1735 57503 1755
rect 57520 1735 57529 1755
rect 57497 1725 57529 1735
rect 57580 1745 57606 1755
rect 57580 1725 57583 1745
rect 57603 1725 57606 1745
rect 57641 1735 57650 1755
rect 57667 1735 57673 1755
rect 57641 1725 57673 1735
rect 57690 1745 57716 1755
rect 57690 1725 57693 1745
rect 57713 1725 57716 1745
rect 57454 1715 57480 1725
rect 57360 1705 57380 1715
rect 57460 1705 57480 1715
rect 57580 1715 57606 1725
rect 57690 1715 57716 1725
rect 57735 1735 57740 1755
rect 57760 1735 57765 1755
rect 57580 1705 57600 1715
rect 57690 1705 57710 1715
rect 57075 1675 57080 1695
rect 57100 1675 57105 1695
rect 57075 1645 57105 1675
rect 57075 1625 57080 1645
rect 57100 1625 57105 1645
rect 57075 1595 57105 1625
rect 57075 1575 57080 1595
rect 57100 1575 57105 1595
rect 57075 1565 57105 1575
rect 57130 1695 57160 1705
rect 57130 1675 57135 1695
rect 57155 1675 57160 1695
rect 57130 1645 57160 1675
rect 57130 1625 57135 1645
rect 57155 1625 57160 1645
rect 57130 1595 57160 1625
rect 57130 1575 57135 1595
rect 57155 1575 57160 1595
rect 57130 1565 57160 1575
rect 57185 1695 57215 1705
rect 57185 1675 57190 1695
rect 57210 1675 57215 1695
rect 57185 1645 57215 1675
rect 57185 1625 57190 1645
rect 57210 1625 57215 1645
rect 57185 1595 57215 1625
rect 57185 1575 57190 1595
rect 57210 1575 57215 1595
rect 57185 1565 57215 1575
rect 57240 1695 57270 1705
rect 57240 1675 57245 1695
rect 57265 1675 57270 1695
rect 57240 1645 57270 1675
rect 57240 1625 57245 1645
rect 57265 1625 57270 1645
rect 57240 1595 57270 1625
rect 57240 1575 57245 1595
rect 57265 1575 57270 1595
rect 57240 1565 57270 1575
rect 57295 1695 57325 1705
rect 57295 1675 57300 1695
rect 57320 1675 57325 1695
rect 57295 1645 57325 1675
rect 57295 1625 57300 1645
rect 57320 1625 57325 1645
rect 57295 1595 57325 1625
rect 57295 1575 57300 1595
rect 57320 1575 57325 1595
rect 57295 1565 57325 1575
rect 57350 1695 57380 1705
rect 57350 1675 57355 1695
rect 57375 1675 57380 1695
rect 57350 1645 57380 1675
rect 57350 1625 57355 1645
rect 57375 1625 57380 1645
rect 57350 1595 57380 1625
rect 57350 1575 57355 1595
rect 57375 1575 57380 1595
rect 57350 1565 57380 1575
rect 57405 1695 57435 1705
rect 57405 1675 57410 1695
rect 57430 1675 57435 1695
rect 57405 1645 57435 1675
rect 57405 1625 57410 1645
rect 57430 1625 57435 1645
rect 57405 1595 57435 1625
rect 57405 1575 57410 1595
rect 57430 1575 57435 1595
rect 57405 1565 57435 1575
rect 57460 1695 57490 1705
rect 57460 1675 57465 1695
rect 57485 1675 57490 1695
rect 57460 1645 57490 1675
rect 57460 1625 57465 1645
rect 57485 1625 57490 1645
rect 57460 1595 57490 1625
rect 57460 1575 57465 1595
rect 57485 1575 57490 1595
rect 57460 1565 57490 1575
rect 57515 1695 57545 1705
rect 57515 1675 57520 1695
rect 57540 1675 57545 1695
rect 57515 1645 57545 1675
rect 57515 1625 57520 1645
rect 57540 1625 57545 1645
rect 57515 1595 57545 1625
rect 57515 1575 57520 1595
rect 57540 1575 57545 1595
rect 57515 1565 57545 1575
rect 57570 1695 57600 1705
rect 57570 1675 57575 1695
rect 57595 1675 57600 1695
rect 57570 1645 57600 1675
rect 57570 1625 57575 1645
rect 57595 1625 57600 1645
rect 57570 1595 57600 1625
rect 57570 1575 57575 1595
rect 57595 1575 57600 1595
rect 57570 1565 57600 1575
rect 57625 1695 57655 1705
rect 57625 1675 57630 1695
rect 57650 1675 57655 1695
rect 57625 1645 57655 1675
rect 57625 1625 57630 1645
rect 57650 1625 57655 1645
rect 57625 1595 57655 1625
rect 57625 1575 57630 1595
rect 57650 1575 57655 1595
rect 57625 1565 57655 1575
rect 57680 1695 57710 1705
rect 57680 1675 57685 1695
rect 57705 1675 57710 1695
rect 57680 1645 57710 1675
rect 57680 1625 57685 1645
rect 57705 1625 57710 1645
rect 57680 1595 57710 1625
rect 57680 1575 57685 1595
rect 57705 1575 57710 1595
rect 57680 1565 57710 1575
rect 57735 1695 57765 1735
rect 57735 1675 57740 1695
rect 57760 1675 57765 1695
rect 57735 1645 57765 1675
rect 57800 1675 57820 1785
rect 57735 1625 57740 1645
rect 57760 1625 57765 1645
rect 57735 1595 57765 1625
rect 57790 1615 57800 1655
rect 58095 1800 58115 1985
rect 58155 1965 58175 1985
rect 58815 1965 58835 1985
rect 57735 1575 57740 1595
rect 57760 1575 57765 1595
rect 57735 1565 57765 1575
rect 57820 1615 57830 1655
rect 58095 1645 58115 1720
rect 56155 1545 56175 1565
rect 56260 1545 56280 1565
rect 56370 1545 56390 1565
rect 56480 1545 56500 1565
rect 56590 1545 56610 1565
rect 56830 1545 56850 1565
rect 56885 1545 56905 1565
rect 57195 1545 57215 1565
rect 57300 1545 57320 1565
rect 57410 1545 57430 1565
rect 57520 1545 57540 1565
rect 57630 1545 57650 1565
rect 56106 1535 56138 1545
rect 56106 1515 56112 1535
rect 56129 1515 56138 1535
rect 56106 1505 56138 1515
rect 56155 1535 56181 1545
rect 56155 1515 56158 1535
rect 56178 1515 56181 1535
rect 56155 1505 56181 1515
rect 56256 1535 56283 1545
rect 56256 1515 56260 1535
rect 56280 1515 56283 1535
rect 56256 1505 56283 1515
rect 56305 1535 56345 1545
rect 56305 1515 56315 1535
rect 56335 1515 56345 1535
rect 56305 1505 56345 1515
rect 56366 1535 56393 1545
rect 56366 1515 56370 1535
rect 56390 1515 56393 1535
rect 56366 1505 56393 1515
rect 56476 1535 56503 1545
rect 56476 1515 56480 1535
rect 56500 1515 56503 1535
rect 56476 1505 56503 1515
rect 56525 1535 56565 1545
rect 56525 1515 56535 1535
rect 56555 1515 56565 1535
rect 56525 1505 56565 1515
rect 56586 1535 56613 1545
rect 56586 1515 56590 1535
rect 56610 1515 56613 1535
rect 56586 1505 56613 1515
rect 56825 1535 56855 1545
rect 56825 1515 56830 1535
rect 56850 1515 56855 1535
rect 56825 1505 56855 1515
rect 56875 1535 56905 1545
rect 56875 1515 56880 1535
rect 56900 1515 56905 1535
rect 56875 1505 56905 1515
rect 56922 1535 56954 1545
rect 56922 1515 56928 1535
rect 56945 1515 56954 1535
rect 56922 1505 56954 1515
rect 57146 1535 57178 1545
rect 57146 1515 57152 1535
rect 57169 1515 57178 1535
rect 57146 1505 57178 1515
rect 57195 1535 57221 1545
rect 57195 1515 57198 1535
rect 57218 1515 57221 1535
rect 57195 1505 57221 1515
rect 57296 1535 57323 1545
rect 57296 1515 57300 1535
rect 57320 1515 57323 1535
rect 57296 1505 57323 1515
rect 57345 1535 57385 1545
rect 57345 1515 57355 1535
rect 57375 1515 57385 1535
rect 57345 1505 57385 1515
rect 57406 1535 57433 1545
rect 57406 1515 57410 1535
rect 57430 1515 57433 1535
rect 57406 1505 57433 1515
rect 57516 1535 57543 1545
rect 57516 1515 57520 1535
rect 57540 1515 57543 1535
rect 57516 1505 57543 1515
rect 57565 1535 57605 1545
rect 57565 1515 57575 1535
rect 57595 1515 57605 1535
rect 57565 1505 57605 1515
rect 57626 1535 57653 1545
rect 57626 1515 57630 1535
rect 57650 1515 57653 1535
rect 57626 1505 57653 1515
rect 57800 1485 57820 1595
rect 58095 1535 58115 1625
rect 58150 1955 58180 1965
rect 58150 1935 58155 1955
rect 58175 1935 58180 1955
rect 58150 1895 58180 1935
rect 58255 1955 58295 1965
rect 58255 1935 58265 1955
rect 58285 1935 58295 1955
rect 58255 1925 58295 1935
rect 58313 1955 58347 1965
rect 58313 1935 58321 1955
rect 58339 1935 58347 1955
rect 58313 1925 58347 1935
rect 58365 1955 58405 1965
rect 58365 1935 58375 1955
rect 58395 1935 58405 1955
rect 58365 1925 58405 1935
rect 58475 1955 58515 1965
rect 58475 1935 58485 1955
rect 58505 1935 58515 1955
rect 58475 1925 58515 1935
rect 58585 1955 58625 1965
rect 58585 1935 58595 1955
rect 58615 1935 58625 1955
rect 58585 1925 58625 1935
rect 58695 1955 58735 1965
rect 58695 1935 58705 1955
rect 58725 1935 58735 1955
rect 58695 1925 58735 1935
rect 58810 1955 58840 1965
rect 58810 1935 58815 1955
rect 58835 1935 58840 1955
rect 58265 1905 58285 1925
rect 58375 1905 58395 1925
rect 58485 1905 58505 1925
rect 58595 1905 58615 1925
rect 58705 1905 58725 1925
rect 58150 1875 58155 1895
rect 58175 1875 58180 1895
rect 58150 1845 58180 1875
rect 58150 1825 58155 1845
rect 58175 1825 58180 1845
rect 58150 1795 58180 1825
rect 58150 1775 58155 1795
rect 58175 1775 58180 1795
rect 58150 1745 58180 1775
rect 58150 1725 58155 1745
rect 58175 1725 58180 1745
rect 58150 1695 58180 1725
rect 58150 1675 58155 1695
rect 58175 1675 58180 1695
rect 58150 1645 58180 1675
rect 58150 1625 58155 1645
rect 58175 1625 58180 1645
rect 58150 1615 58180 1625
rect 58205 1895 58235 1905
rect 58205 1875 58210 1895
rect 58230 1875 58235 1895
rect 58205 1845 58235 1875
rect 58205 1825 58210 1845
rect 58230 1825 58235 1845
rect 58205 1795 58235 1825
rect 58205 1775 58210 1795
rect 58230 1775 58235 1795
rect 58205 1745 58235 1775
rect 58205 1725 58210 1745
rect 58230 1725 58235 1745
rect 58205 1695 58235 1725
rect 58205 1675 58210 1695
rect 58230 1675 58235 1695
rect 58205 1645 58235 1675
rect 58205 1625 58210 1645
rect 58230 1625 58235 1645
rect 58205 1615 58235 1625
rect 58260 1895 58290 1905
rect 58260 1875 58265 1895
rect 58285 1875 58290 1895
rect 58260 1845 58290 1875
rect 58260 1825 58265 1845
rect 58285 1825 58290 1845
rect 58260 1795 58290 1825
rect 58260 1775 58265 1795
rect 58285 1775 58290 1795
rect 58260 1745 58290 1775
rect 58260 1725 58265 1745
rect 58285 1725 58290 1745
rect 58260 1695 58290 1725
rect 58260 1675 58265 1695
rect 58285 1675 58290 1695
rect 58260 1645 58290 1675
rect 58260 1625 58265 1645
rect 58285 1625 58290 1645
rect 58260 1615 58290 1625
rect 58315 1895 58345 1905
rect 58315 1875 58320 1895
rect 58340 1875 58345 1895
rect 58315 1845 58345 1875
rect 58315 1825 58320 1845
rect 58340 1825 58345 1845
rect 58315 1795 58345 1825
rect 58315 1775 58320 1795
rect 58340 1775 58345 1795
rect 58315 1745 58345 1775
rect 58315 1725 58320 1745
rect 58340 1725 58345 1745
rect 58315 1695 58345 1725
rect 58315 1675 58320 1695
rect 58340 1675 58345 1695
rect 58315 1645 58345 1675
rect 58315 1625 58320 1645
rect 58340 1625 58345 1645
rect 58315 1615 58345 1625
rect 58370 1895 58400 1905
rect 58370 1875 58375 1895
rect 58395 1875 58400 1895
rect 58370 1845 58400 1875
rect 58370 1825 58375 1845
rect 58395 1825 58400 1845
rect 58370 1795 58400 1825
rect 58370 1775 58375 1795
rect 58395 1775 58400 1795
rect 58370 1745 58400 1775
rect 58370 1725 58375 1745
rect 58395 1725 58400 1745
rect 58370 1695 58400 1725
rect 58370 1675 58375 1695
rect 58395 1675 58400 1695
rect 58370 1645 58400 1675
rect 58370 1625 58375 1645
rect 58395 1625 58400 1645
rect 58370 1615 58400 1625
rect 58425 1895 58455 1905
rect 58425 1875 58430 1895
rect 58450 1875 58455 1895
rect 58425 1845 58455 1875
rect 58425 1825 58430 1845
rect 58450 1825 58455 1845
rect 58425 1795 58455 1825
rect 58425 1775 58430 1795
rect 58450 1775 58455 1795
rect 58425 1745 58455 1775
rect 58425 1725 58430 1745
rect 58450 1725 58455 1745
rect 58425 1695 58455 1725
rect 58425 1675 58430 1695
rect 58450 1675 58455 1695
rect 58425 1645 58455 1675
rect 58425 1625 58430 1645
rect 58450 1625 58455 1645
rect 58425 1615 58455 1625
rect 58480 1895 58510 1905
rect 58480 1875 58485 1895
rect 58505 1875 58510 1895
rect 58480 1845 58510 1875
rect 58480 1825 58485 1845
rect 58505 1825 58510 1845
rect 58480 1795 58510 1825
rect 58480 1775 58485 1795
rect 58505 1775 58510 1795
rect 58480 1745 58510 1775
rect 58480 1725 58485 1745
rect 58505 1725 58510 1745
rect 58480 1695 58510 1725
rect 58480 1675 58485 1695
rect 58505 1675 58510 1695
rect 58480 1645 58510 1675
rect 58480 1625 58485 1645
rect 58505 1625 58510 1645
rect 58480 1615 58510 1625
rect 58535 1895 58565 1905
rect 58535 1875 58540 1895
rect 58560 1875 58565 1895
rect 58535 1845 58565 1875
rect 58535 1825 58540 1845
rect 58560 1825 58565 1845
rect 58535 1795 58565 1825
rect 58535 1775 58540 1795
rect 58560 1775 58565 1795
rect 58535 1745 58565 1775
rect 58535 1725 58540 1745
rect 58560 1725 58565 1745
rect 58535 1695 58565 1725
rect 58535 1675 58540 1695
rect 58560 1675 58565 1695
rect 58535 1645 58565 1675
rect 58535 1625 58540 1645
rect 58560 1625 58565 1645
rect 58535 1615 58565 1625
rect 58590 1895 58620 1905
rect 58590 1875 58595 1895
rect 58615 1875 58620 1895
rect 58590 1845 58620 1875
rect 58590 1825 58595 1845
rect 58615 1825 58620 1845
rect 58590 1795 58620 1825
rect 58590 1775 58595 1795
rect 58615 1775 58620 1795
rect 58590 1745 58620 1775
rect 58590 1725 58595 1745
rect 58615 1725 58620 1745
rect 58590 1695 58620 1725
rect 58590 1675 58595 1695
rect 58615 1675 58620 1695
rect 58590 1645 58620 1675
rect 58590 1625 58595 1645
rect 58615 1625 58620 1645
rect 58590 1615 58620 1625
rect 58645 1895 58675 1905
rect 58645 1875 58650 1895
rect 58670 1875 58675 1895
rect 58645 1845 58675 1875
rect 58645 1825 58650 1845
rect 58670 1825 58675 1845
rect 58645 1795 58675 1825
rect 58645 1775 58650 1795
rect 58670 1775 58675 1795
rect 58645 1745 58675 1775
rect 58645 1725 58650 1745
rect 58670 1725 58675 1745
rect 58645 1695 58675 1725
rect 58645 1675 58650 1695
rect 58670 1675 58675 1695
rect 58645 1645 58675 1675
rect 58645 1625 58650 1645
rect 58670 1625 58675 1645
rect 58645 1615 58675 1625
rect 58700 1895 58730 1905
rect 58700 1875 58705 1895
rect 58725 1875 58730 1895
rect 58700 1845 58730 1875
rect 58700 1825 58705 1845
rect 58725 1825 58730 1845
rect 58700 1795 58730 1825
rect 58700 1775 58705 1795
rect 58725 1775 58730 1795
rect 58700 1745 58730 1775
rect 58700 1725 58705 1745
rect 58725 1725 58730 1745
rect 58700 1695 58730 1725
rect 58700 1675 58705 1695
rect 58725 1675 58730 1695
rect 58700 1645 58730 1675
rect 58700 1625 58705 1645
rect 58725 1625 58730 1645
rect 58700 1615 58730 1625
rect 58755 1895 58785 1905
rect 58755 1875 58760 1895
rect 58780 1875 58785 1895
rect 58755 1845 58785 1875
rect 58755 1825 58760 1845
rect 58780 1825 58785 1845
rect 58755 1795 58785 1825
rect 58755 1775 58760 1795
rect 58780 1775 58785 1795
rect 58755 1745 58785 1775
rect 58755 1725 58760 1745
rect 58780 1725 58785 1745
rect 58755 1695 58785 1725
rect 58755 1675 58760 1695
rect 58780 1675 58785 1695
rect 58755 1645 58785 1675
rect 58755 1625 58760 1645
rect 58780 1625 58785 1645
rect 58755 1615 58785 1625
rect 58810 1895 58840 1935
rect 58810 1875 58815 1895
rect 58835 1875 58840 1895
rect 58810 1845 58840 1875
rect 58810 1825 58815 1845
rect 58835 1825 58840 1845
rect 58810 1795 58840 1825
rect 58810 1775 58815 1795
rect 58835 1775 58840 1795
rect 58810 1745 58840 1775
rect 58810 1725 58815 1745
rect 58835 1725 58840 1745
rect 58810 1695 58840 1725
rect 58810 1675 58815 1695
rect 58835 1675 58840 1695
rect 58810 1645 58840 1675
rect 58810 1625 58815 1645
rect 58835 1625 58840 1645
rect 58810 1615 58840 1625
rect 58875 1800 58895 1985
rect 59045 1945 59065 2280
rect 59115 2216 59330 2236
rect 59115 2199 59150 2216
rect 59295 2199 59330 2216
rect 59210 2149 59235 2199
rect 59045 1780 59065 1865
rect 59380 1945 59400 2280
rect 58895 1770 58915 1780
rect 58905 1750 58915 1770
rect 58895 1740 58915 1750
rect 59025 1770 59065 1780
rect 59025 1750 59035 1770
rect 59055 1750 59065 1770
rect 59025 1740 59065 1750
rect 58210 1595 58230 1615
rect 58320 1595 58340 1615
rect 58430 1595 58450 1615
rect 58540 1595 58560 1615
rect 58650 1595 58670 1615
rect 58760 1595 58780 1615
rect 58200 1585 58240 1595
rect 58200 1565 58212 1585
rect 58230 1565 58240 1585
rect 58200 1555 58240 1565
rect 58310 1585 58350 1595
rect 58310 1565 58322 1585
rect 58340 1565 58350 1585
rect 58310 1555 58350 1565
rect 58420 1585 58460 1595
rect 58420 1565 58432 1585
rect 58450 1565 58460 1585
rect 58420 1555 58460 1565
rect 58530 1585 58570 1595
rect 58530 1565 58542 1585
rect 58560 1565 58570 1585
rect 58530 1555 58570 1565
rect 58640 1585 58680 1595
rect 58640 1565 58652 1585
rect 58670 1565 58680 1585
rect 58640 1555 58680 1565
rect 58750 1585 58790 1595
rect 58750 1565 58762 1585
rect 58780 1565 58790 1585
rect 58750 1555 58790 1565
rect 58875 1535 58895 1720
rect 58095 1515 58455 1535
rect 58535 1515 58895 1535
rect 59045 1535 59065 1740
rect 59115 1590 59150 1600
rect 59115 1565 59120 1590
rect 59145 1565 59150 1590
rect 59115 1555 59150 1565
rect 59175 1590 59210 1600
rect 59175 1565 59180 1590
rect 59205 1565 59210 1590
rect 59175 1555 59210 1565
rect 59235 1590 59270 1600
rect 59235 1565 59240 1590
rect 59265 1565 59270 1590
rect 59235 1555 59270 1565
rect 59295 1590 59330 1600
rect 59295 1565 59300 1590
rect 59325 1565 59330 1590
rect 59295 1555 59330 1565
rect 59380 1535 59400 1865
rect 59045 1515 59185 1535
rect 59265 1515 59400 1535
rect 58475 1505 58485 1515
rect 58505 1505 58515 1515
rect 58475 1495 58515 1505
rect 55980 1465 56860 1485
rect 56940 1465 57820 1485
rect 55285 1425 55325 1435
rect 55285 1415 55295 1425
rect 54985 1405 55295 1415
rect 55315 1415 55325 1425
rect 58475 1425 58515 1435
rect 58475 1415 58485 1425
rect 54985 1395 55315 1405
rect 55395 1395 55725 1415
rect 54660 1340 54735 1360
rect 54815 1340 54895 1360
rect 54660 965 54680 1340
rect 54730 1305 54765 1315
rect 54730 1280 54735 1305
rect 54760 1280 54765 1305
rect 54730 1270 54765 1280
rect 54790 1305 54825 1315
rect 54790 1280 54795 1305
rect 54820 1280 54825 1305
rect 54790 1270 54825 1280
rect 54660 533 54680 885
rect 54875 990 54895 1340
rect 54985 1010 55005 1395
rect 55045 1375 55065 1395
rect 55645 1375 55665 1395
rect 54875 980 54915 990
rect 54875 965 54885 980
rect 54905 960 54915 980
rect 54895 950 54915 960
rect 54965 980 54985 990
rect 54965 960 54975 980
rect 54965 950 54985 960
rect 54765 583 54790 633
rect 54875 533 54895 885
rect 54660 513 54735 533
rect 54815 513 54895 533
rect 54985 545 55005 930
rect 55040 1365 55070 1375
rect 55040 1345 55045 1365
rect 55065 1345 55070 1365
rect 55040 1305 55070 1345
rect 55135 1365 55175 1375
rect 55135 1345 55145 1365
rect 55165 1345 55175 1365
rect 55135 1335 55175 1345
rect 55335 1365 55375 1375
rect 55335 1345 55345 1365
rect 55365 1345 55375 1365
rect 55335 1335 55375 1345
rect 55438 1365 55472 1375
rect 55438 1345 55446 1365
rect 55464 1345 55472 1365
rect 55438 1335 55472 1345
rect 55535 1365 55575 1375
rect 55535 1345 55545 1365
rect 55565 1345 55575 1365
rect 55535 1335 55575 1345
rect 55640 1365 55670 1375
rect 55640 1345 55645 1365
rect 55665 1345 55670 1365
rect 55145 1315 55165 1335
rect 55345 1315 55365 1335
rect 55545 1315 55565 1335
rect 55040 1285 55045 1305
rect 55065 1285 55070 1305
rect 55040 1255 55070 1285
rect 55040 1235 55045 1255
rect 55065 1235 55070 1255
rect 55040 1205 55070 1235
rect 55040 1185 55045 1205
rect 55065 1185 55070 1205
rect 55040 1155 55070 1185
rect 55040 1135 55045 1155
rect 55065 1135 55070 1155
rect 55040 1105 55070 1135
rect 55040 1085 55045 1105
rect 55065 1085 55070 1105
rect 55040 1055 55070 1085
rect 55040 1035 55045 1055
rect 55065 1035 55070 1055
rect 55040 1005 55070 1035
rect 55040 985 55045 1005
rect 55065 985 55070 1005
rect 55040 955 55070 985
rect 55040 935 55045 955
rect 55065 935 55070 955
rect 55040 905 55070 935
rect 55040 885 55045 905
rect 55065 885 55070 905
rect 55040 855 55070 885
rect 55040 835 55045 855
rect 55065 835 55070 855
rect 55040 805 55070 835
rect 55040 785 55045 805
rect 55065 785 55070 805
rect 55040 755 55070 785
rect 55040 735 55045 755
rect 55065 735 55070 755
rect 55040 705 55070 735
rect 55040 685 55045 705
rect 55065 685 55070 705
rect 55040 655 55070 685
rect 55040 635 55045 655
rect 55065 635 55070 655
rect 55040 625 55070 635
rect 55140 1305 55170 1315
rect 55140 1285 55145 1305
rect 55165 1285 55170 1305
rect 55140 1255 55170 1285
rect 55140 1235 55145 1255
rect 55165 1235 55170 1255
rect 55140 1205 55170 1235
rect 55140 1185 55145 1205
rect 55165 1185 55170 1205
rect 55140 1155 55170 1185
rect 55140 1135 55145 1155
rect 55165 1135 55170 1155
rect 55140 1105 55170 1135
rect 55140 1085 55145 1105
rect 55165 1085 55170 1105
rect 55140 1055 55170 1085
rect 55140 1035 55145 1055
rect 55165 1035 55170 1055
rect 55140 1005 55170 1035
rect 55140 985 55145 1005
rect 55165 985 55170 1005
rect 55140 955 55170 985
rect 55140 935 55145 955
rect 55165 935 55170 955
rect 55140 905 55170 935
rect 55140 885 55145 905
rect 55165 885 55170 905
rect 55140 855 55170 885
rect 55140 835 55145 855
rect 55165 835 55170 855
rect 55140 805 55170 835
rect 55140 785 55145 805
rect 55165 785 55170 805
rect 55140 755 55170 785
rect 55140 735 55145 755
rect 55165 735 55170 755
rect 55140 705 55170 735
rect 55140 685 55145 705
rect 55165 685 55170 705
rect 55140 655 55170 685
rect 55140 635 55145 655
rect 55165 635 55170 655
rect 55140 625 55170 635
rect 55240 1305 55270 1315
rect 55240 1285 55245 1305
rect 55265 1285 55270 1305
rect 55240 1255 55270 1285
rect 55240 1235 55245 1255
rect 55265 1235 55270 1255
rect 55240 1205 55270 1235
rect 55240 1185 55245 1205
rect 55265 1185 55270 1205
rect 55240 1155 55270 1185
rect 55240 1135 55245 1155
rect 55265 1135 55270 1155
rect 55240 1105 55270 1135
rect 55240 1085 55245 1105
rect 55265 1085 55270 1105
rect 55240 1055 55270 1085
rect 55240 1035 55245 1055
rect 55265 1035 55270 1055
rect 55240 1005 55270 1035
rect 55240 985 55245 1005
rect 55265 985 55270 1005
rect 55240 955 55270 985
rect 55240 935 55245 955
rect 55265 935 55270 955
rect 55240 905 55270 935
rect 55240 885 55245 905
rect 55265 885 55270 905
rect 55240 855 55270 885
rect 55240 835 55245 855
rect 55265 835 55270 855
rect 55240 805 55270 835
rect 55240 785 55245 805
rect 55265 785 55270 805
rect 55240 755 55270 785
rect 55240 735 55245 755
rect 55265 735 55270 755
rect 55240 705 55270 735
rect 55240 685 55245 705
rect 55265 685 55270 705
rect 55240 655 55270 685
rect 55240 635 55245 655
rect 55265 635 55270 655
rect 55240 625 55270 635
rect 55340 1305 55370 1315
rect 55340 1285 55345 1305
rect 55365 1285 55370 1305
rect 55340 1255 55370 1285
rect 55340 1235 55345 1255
rect 55365 1235 55370 1255
rect 55340 1205 55370 1235
rect 55340 1185 55345 1205
rect 55365 1185 55370 1205
rect 55340 1155 55370 1185
rect 55340 1135 55345 1155
rect 55365 1135 55370 1155
rect 55340 1105 55370 1135
rect 55340 1085 55345 1105
rect 55365 1085 55370 1105
rect 55340 1055 55370 1085
rect 55340 1035 55345 1055
rect 55365 1035 55370 1055
rect 55340 1005 55370 1035
rect 55340 985 55345 1005
rect 55365 985 55370 1005
rect 55340 955 55370 985
rect 55340 935 55345 955
rect 55365 935 55370 955
rect 55340 905 55370 935
rect 55340 885 55345 905
rect 55365 885 55370 905
rect 55340 855 55370 885
rect 55340 835 55345 855
rect 55365 835 55370 855
rect 55340 805 55370 835
rect 55340 785 55345 805
rect 55365 785 55370 805
rect 55340 755 55370 785
rect 55340 735 55345 755
rect 55365 735 55370 755
rect 55340 705 55370 735
rect 55340 685 55345 705
rect 55365 685 55370 705
rect 55340 655 55370 685
rect 55340 635 55345 655
rect 55365 635 55370 655
rect 55340 625 55370 635
rect 55440 1305 55470 1315
rect 55440 1285 55445 1305
rect 55465 1285 55470 1305
rect 55440 1255 55470 1285
rect 55440 1235 55445 1255
rect 55465 1235 55470 1255
rect 55440 1205 55470 1235
rect 55440 1185 55445 1205
rect 55465 1185 55470 1205
rect 55440 1155 55470 1185
rect 55440 1135 55445 1155
rect 55465 1135 55470 1155
rect 55440 1105 55470 1135
rect 55440 1085 55445 1105
rect 55465 1085 55470 1105
rect 55440 1055 55470 1085
rect 55440 1035 55445 1055
rect 55465 1035 55470 1055
rect 55440 1005 55470 1035
rect 55440 985 55445 1005
rect 55465 985 55470 1005
rect 55440 955 55470 985
rect 55440 935 55445 955
rect 55465 935 55470 955
rect 55440 905 55470 935
rect 55440 885 55445 905
rect 55465 885 55470 905
rect 55440 855 55470 885
rect 55440 835 55445 855
rect 55465 835 55470 855
rect 55440 805 55470 835
rect 55440 785 55445 805
rect 55465 785 55470 805
rect 55440 755 55470 785
rect 55440 735 55445 755
rect 55465 735 55470 755
rect 55440 705 55470 735
rect 55440 685 55445 705
rect 55465 685 55470 705
rect 55440 655 55470 685
rect 55440 635 55445 655
rect 55465 635 55470 655
rect 55440 625 55470 635
rect 55540 1305 55570 1315
rect 55540 1285 55545 1305
rect 55565 1285 55570 1305
rect 55540 1255 55570 1285
rect 55540 1235 55545 1255
rect 55565 1235 55570 1255
rect 55540 1205 55570 1235
rect 55540 1185 55545 1205
rect 55565 1185 55570 1205
rect 55540 1155 55570 1185
rect 55540 1135 55545 1155
rect 55565 1135 55570 1155
rect 55540 1105 55570 1135
rect 55540 1085 55545 1105
rect 55565 1085 55570 1105
rect 55540 1055 55570 1085
rect 55540 1035 55545 1055
rect 55565 1035 55570 1055
rect 55540 1005 55570 1035
rect 55540 985 55545 1005
rect 55565 985 55570 1005
rect 55540 955 55570 985
rect 55540 935 55545 955
rect 55565 935 55570 955
rect 55540 905 55570 935
rect 55540 885 55545 905
rect 55565 885 55570 905
rect 55540 855 55570 885
rect 55540 835 55545 855
rect 55565 835 55570 855
rect 55540 805 55570 835
rect 55540 785 55545 805
rect 55565 785 55570 805
rect 55540 755 55570 785
rect 55540 735 55545 755
rect 55565 735 55570 755
rect 55540 705 55570 735
rect 55540 685 55545 705
rect 55565 685 55570 705
rect 55540 655 55570 685
rect 55540 635 55545 655
rect 55565 635 55570 655
rect 55540 625 55570 635
rect 55640 1305 55670 1345
rect 55640 1285 55645 1305
rect 55665 1285 55670 1305
rect 55640 1255 55670 1285
rect 55640 1235 55645 1255
rect 55665 1235 55670 1255
rect 55640 1205 55670 1235
rect 55640 1185 55645 1205
rect 55665 1185 55670 1205
rect 55640 1155 55670 1185
rect 55640 1135 55645 1155
rect 55665 1135 55670 1155
rect 55640 1105 55670 1135
rect 55640 1085 55645 1105
rect 55665 1085 55670 1105
rect 55640 1055 55670 1085
rect 55640 1035 55645 1055
rect 55665 1035 55670 1055
rect 55640 1005 55670 1035
rect 55640 985 55645 1005
rect 55665 985 55670 1005
rect 55640 955 55670 985
rect 55640 935 55645 955
rect 55665 935 55670 955
rect 55640 905 55670 935
rect 55640 885 55645 905
rect 55665 885 55670 905
rect 55640 855 55670 885
rect 55640 835 55645 855
rect 55665 835 55670 855
rect 55640 805 55670 835
rect 55640 785 55645 805
rect 55665 785 55670 805
rect 55640 755 55670 785
rect 55640 735 55645 755
rect 55665 735 55670 755
rect 55640 705 55670 735
rect 55640 685 55645 705
rect 55665 685 55670 705
rect 55640 655 55670 685
rect 55640 635 55645 655
rect 55665 635 55670 655
rect 55640 625 55670 635
rect 55705 1010 55725 1395
rect 58075 1395 58405 1415
rect 58505 1415 58515 1425
rect 58505 1405 58815 1415
rect 58485 1395 58815 1405
rect 55245 605 55265 625
rect 55445 605 55465 625
rect 55235 595 55275 605
rect 55235 575 55245 595
rect 55265 575 55275 595
rect 55235 565 55275 575
rect 55435 595 55475 605
rect 55435 575 55445 595
rect 55465 575 55475 595
rect 55435 565 55475 575
rect 55705 545 55725 930
rect 56170 1280 56860 1300
rect 56940 1280 57440 1300
rect 57520 1280 57635 1300
rect 56170 1100 56190 1280
rect 56330 1250 56370 1260
rect 56330 1230 56340 1250
rect 56360 1230 56370 1250
rect 56330 1220 56370 1230
rect 56440 1250 56480 1260
rect 56440 1230 56450 1250
rect 56470 1230 56480 1250
rect 56440 1220 56480 1230
rect 56550 1250 56590 1260
rect 56550 1230 56560 1250
rect 56580 1230 56590 1250
rect 56550 1220 56590 1230
rect 56660 1250 56700 1260
rect 56660 1230 56670 1250
rect 56690 1230 56700 1250
rect 56660 1220 56700 1230
rect 56770 1250 56810 1260
rect 56770 1230 56780 1250
rect 56800 1230 56810 1250
rect 56770 1220 56810 1230
rect 56830 1250 56860 1260
rect 56830 1230 56835 1250
rect 56855 1230 56860 1250
rect 56830 1220 56860 1230
rect 56880 1250 56920 1260
rect 56880 1230 56890 1250
rect 56910 1230 56920 1250
rect 56880 1220 56920 1230
rect 56990 1250 57030 1260
rect 56990 1230 57000 1250
rect 57020 1230 57030 1250
rect 56990 1220 57030 1230
rect 57100 1250 57140 1260
rect 57100 1230 57110 1250
rect 57130 1230 57140 1250
rect 57100 1220 57140 1230
rect 57210 1250 57250 1260
rect 57210 1230 57220 1250
rect 57240 1230 57250 1250
rect 57210 1220 57250 1230
rect 57320 1250 57360 1260
rect 57320 1230 57330 1250
rect 57350 1230 57360 1250
rect 57320 1220 57360 1230
rect 57415 1250 57455 1260
rect 57415 1230 57425 1250
rect 57445 1230 57455 1250
rect 57415 1220 57455 1230
rect 57474 1250 57504 1260
rect 57474 1230 57479 1250
rect 57499 1230 57504 1250
rect 57474 1220 57504 1230
rect 56340 1200 56360 1220
rect 56450 1200 56470 1220
rect 56560 1200 56580 1220
rect 56670 1200 56690 1220
rect 56780 1200 56800 1220
rect 56890 1200 56910 1220
rect 57000 1200 57020 1220
rect 57110 1200 57130 1220
rect 57220 1200 57240 1220
rect 57330 1200 57350 1220
rect 57435 1200 57455 1220
rect 56170 875 56190 1020
rect 56225 1190 56255 1200
rect 56225 1170 56230 1190
rect 56250 1170 56255 1190
rect 56225 1140 56255 1170
rect 56225 1120 56230 1140
rect 56250 1120 56255 1140
rect 56225 1090 56255 1120
rect 56225 1070 56230 1090
rect 56250 1070 56255 1090
rect 56225 1040 56255 1070
rect 56225 1020 56230 1040
rect 56250 1020 56255 1040
rect 56225 990 56255 1020
rect 56225 970 56230 990
rect 56250 970 56255 990
rect 56225 960 56255 970
rect 56280 1190 56310 1200
rect 56280 1170 56285 1190
rect 56305 1170 56310 1190
rect 56280 1140 56310 1170
rect 56280 1120 56285 1140
rect 56305 1120 56310 1140
rect 56280 1090 56310 1120
rect 56280 1070 56285 1090
rect 56305 1070 56310 1090
rect 56280 1040 56310 1070
rect 56280 1020 56285 1040
rect 56305 1020 56310 1040
rect 56280 990 56310 1020
rect 56280 970 56285 990
rect 56305 970 56310 990
rect 56280 960 56310 970
rect 56335 1190 56365 1200
rect 56335 1170 56340 1190
rect 56360 1170 56365 1190
rect 56335 1140 56365 1170
rect 56335 1120 56340 1140
rect 56360 1120 56365 1140
rect 56335 1090 56365 1120
rect 56335 1070 56340 1090
rect 56360 1070 56365 1090
rect 56335 1040 56365 1070
rect 56335 1020 56340 1040
rect 56360 1020 56365 1040
rect 56335 990 56365 1020
rect 56335 970 56340 990
rect 56360 970 56365 990
rect 56335 960 56365 970
rect 56390 1190 56420 1200
rect 56390 1170 56395 1190
rect 56415 1170 56420 1190
rect 56390 1140 56420 1170
rect 56390 1120 56395 1140
rect 56415 1120 56420 1140
rect 56390 1090 56420 1120
rect 56390 1070 56395 1090
rect 56415 1070 56420 1090
rect 56390 1040 56420 1070
rect 56390 1020 56395 1040
rect 56415 1020 56420 1040
rect 56390 990 56420 1020
rect 56390 970 56395 990
rect 56415 970 56420 990
rect 56390 960 56420 970
rect 56445 1190 56475 1200
rect 56445 1170 56450 1190
rect 56470 1170 56475 1190
rect 56445 1140 56475 1170
rect 56445 1120 56450 1140
rect 56470 1120 56475 1140
rect 56445 1090 56475 1120
rect 56445 1070 56450 1090
rect 56470 1070 56475 1090
rect 56445 1040 56475 1070
rect 56445 1020 56450 1040
rect 56470 1020 56475 1040
rect 56445 990 56475 1020
rect 56445 970 56450 990
rect 56470 970 56475 990
rect 56445 960 56475 970
rect 56500 1190 56530 1200
rect 56500 1170 56505 1190
rect 56525 1170 56530 1190
rect 56500 1140 56530 1170
rect 56500 1120 56505 1140
rect 56525 1120 56530 1140
rect 56500 1090 56530 1120
rect 56500 1070 56505 1090
rect 56525 1070 56530 1090
rect 56500 1040 56530 1070
rect 56500 1020 56505 1040
rect 56525 1020 56530 1040
rect 56500 990 56530 1020
rect 56500 970 56505 990
rect 56525 970 56530 990
rect 56500 960 56530 970
rect 56555 1190 56585 1200
rect 56555 1170 56560 1190
rect 56580 1170 56585 1190
rect 56555 1140 56585 1170
rect 56555 1120 56560 1140
rect 56580 1120 56585 1140
rect 56555 1090 56585 1120
rect 56555 1070 56560 1090
rect 56580 1070 56585 1090
rect 56555 1040 56585 1070
rect 56555 1020 56560 1040
rect 56580 1020 56585 1040
rect 56555 990 56585 1020
rect 56555 970 56560 990
rect 56580 970 56585 990
rect 56555 960 56585 970
rect 56610 1190 56640 1200
rect 56610 1170 56615 1190
rect 56635 1170 56640 1190
rect 56610 1140 56640 1170
rect 56610 1120 56615 1140
rect 56635 1120 56640 1140
rect 56610 1090 56640 1120
rect 56610 1070 56615 1090
rect 56635 1070 56640 1090
rect 56610 1040 56640 1070
rect 56610 1020 56615 1040
rect 56635 1020 56640 1040
rect 56610 990 56640 1020
rect 56610 970 56615 990
rect 56635 970 56640 990
rect 56610 960 56640 970
rect 56665 1190 56695 1200
rect 56665 1170 56670 1190
rect 56690 1170 56695 1190
rect 56665 1140 56695 1170
rect 56665 1120 56670 1140
rect 56690 1120 56695 1140
rect 56665 1090 56695 1120
rect 56665 1070 56670 1090
rect 56690 1070 56695 1090
rect 56665 1040 56695 1070
rect 56665 1020 56670 1040
rect 56690 1020 56695 1040
rect 56665 990 56695 1020
rect 56665 970 56670 990
rect 56690 970 56695 990
rect 56665 960 56695 970
rect 56720 1190 56750 1200
rect 56720 1170 56725 1190
rect 56745 1170 56750 1190
rect 56720 1140 56750 1170
rect 56720 1120 56725 1140
rect 56745 1120 56750 1140
rect 56720 1090 56750 1120
rect 56720 1070 56725 1090
rect 56745 1070 56750 1090
rect 56720 1040 56750 1070
rect 56720 1020 56725 1040
rect 56745 1020 56750 1040
rect 56720 990 56750 1020
rect 56720 970 56725 990
rect 56745 970 56750 990
rect 56720 960 56750 970
rect 56775 1190 56805 1200
rect 56775 1170 56780 1190
rect 56800 1170 56805 1190
rect 56775 1140 56805 1170
rect 56775 1120 56780 1140
rect 56800 1120 56805 1140
rect 56775 1090 56805 1120
rect 56775 1070 56780 1090
rect 56800 1070 56805 1090
rect 56775 1040 56805 1070
rect 56775 1020 56780 1040
rect 56800 1020 56805 1040
rect 56775 990 56805 1020
rect 56775 970 56780 990
rect 56800 970 56805 990
rect 56775 960 56805 970
rect 56830 1190 56860 1200
rect 56830 1170 56835 1190
rect 56855 1170 56860 1190
rect 56830 1140 56860 1170
rect 56830 1120 56835 1140
rect 56855 1120 56860 1140
rect 56830 1090 56860 1120
rect 56830 1070 56835 1090
rect 56855 1070 56860 1090
rect 56830 1040 56860 1070
rect 56830 1020 56835 1040
rect 56855 1020 56860 1040
rect 56830 990 56860 1020
rect 56830 970 56835 990
rect 56855 970 56860 990
rect 56830 960 56860 970
rect 56885 1190 56915 1200
rect 56885 1170 56890 1190
rect 56910 1170 56915 1190
rect 56885 1140 56915 1170
rect 56885 1120 56890 1140
rect 56910 1120 56915 1140
rect 56885 1090 56915 1120
rect 56885 1070 56890 1090
rect 56910 1070 56915 1090
rect 56885 1040 56915 1070
rect 56885 1020 56890 1040
rect 56910 1020 56915 1040
rect 56885 990 56915 1020
rect 56885 970 56890 990
rect 56910 970 56915 990
rect 56885 960 56915 970
rect 56940 1190 56970 1200
rect 56940 1170 56945 1190
rect 56965 1170 56970 1190
rect 56940 1140 56970 1170
rect 56940 1120 56945 1140
rect 56965 1120 56970 1140
rect 56940 1090 56970 1120
rect 56940 1070 56945 1090
rect 56965 1070 56970 1090
rect 56940 1040 56970 1070
rect 56940 1020 56945 1040
rect 56965 1020 56970 1040
rect 56940 990 56970 1020
rect 56940 970 56945 990
rect 56965 970 56970 990
rect 56940 960 56970 970
rect 56995 1190 57025 1200
rect 56995 1170 57000 1190
rect 57020 1170 57025 1190
rect 56995 1140 57025 1170
rect 56995 1120 57000 1140
rect 57020 1120 57025 1140
rect 56995 1090 57025 1120
rect 56995 1070 57000 1090
rect 57020 1070 57025 1090
rect 56995 1040 57025 1070
rect 56995 1020 57000 1040
rect 57020 1020 57025 1040
rect 56995 990 57025 1020
rect 56995 970 57000 990
rect 57020 970 57025 990
rect 56995 960 57025 970
rect 57050 1190 57080 1200
rect 57050 1170 57055 1190
rect 57075 1170 57080 1190
rect 57050 1140 57080 1170
rect 57050 1120 57055 1140
rect 57075 1120 57080 1140
rect 57050 1090 57080 1120
rect 57050 1070 57055 1090
rect 57075 1070 57080 1090
rect 57050 1040 57080 1070
rect 57050 1020 57055 1040
rect 57075 1020 57080 1040
rect 57050 990 57080 1020
rect 57050 970 57055 990
rect 57075 970 57080 990
rect 57050 960 57080 970
rect 57105 1190 57135 1200
rect 57105 1170 57110 1190
rect 57130 1170 57135 1190
rect 57105 1140 57135 1170
rect 57105 1120 57110 1140
rect 57130 1120 57135 1140
rect 57105 1090 57135 1120
rect 57105 1070 57110 1090
rect 57130 1070 57135 1090
rect 57105 1040 57135 1070
rect 57105 1020 57110 1040
rect 57130 1020 57135 1040
rect 57105 990 57135 1020
rect 57105 970 57110 990
rect 57130 970 57135 990
rect 57105 960 57135 970
rect 57160 1190 57190 1200
rect 57160 1170 57165 1190
rect 57185 1170 57190 1190
rect 57160 1140 57190 1170
rect 57160 1120 57165 1140
rect 57185 1120 57190 1140
rect 57160 1090 57190 1120
rect 57160 1070 57165 1090
rect 57185 1070 57190 1090
rect 57160 1040 57190 1070
rect 57160 1020 57165 1040
rect 57185 1020 57190 1040
rect 57160 990 57190 1020
rect 57160 970 57165 990
rect 57185 970 57190 990
rect 57160 960 57190 970
rect 57215 1190 57245 1200
rect 57215 1170 57220 1190
rect 57240 1170 57245 1190
rect 57215 1140 57245 1170
rect 57215 1120 57220 1140
rect 57240 1120 57245 1140
rect 57215 1090 57245 1120
rect 57215 1070 57220 1090
rect 57240 1070 57245 1090
rect 57215 1040 57245 1070
rect 57215 1020 57220 1040
rect 57240 1020 57245 1040
rect 57215 990 57245 1020
rect 57215 970 57220 990
rect 57240 970 57245 990
rect 57215 960 57245 970
rect 57270 1190 57300 1200
rect 57270 1170 57275 1190
rect 57295 1170 57300 1190
rect 57270 1140 57300 1170
rect 57270 1120 57275 1140
rect 57295 1120 57300 1140
rect 57270 1090 57300 1120
rect 57270 1070 57275 1090
rect 57295 1070 57300 1090
rect 57270 1040 57300 1070
rect 57270 1020 57275 1040
rect 57295 1020 57300 1040
rect 57270 990 57300 1020
rect 57270 970 57275 990
rect 57295 970 57300 990
rect 57270 960 57300 970
rect 57325 1190 57355 1200
rect 57325 1170 57330 1190
rect 57350 1170 57355 1190
rect 57325 1140 57355 1170
rect 57325 1120 57330 1140
rect 57350 1120 57355 1140
rect 57325 1090 57355 1120
rect 57325 1070 57330 1090
rect 57350 1070 57355 1090
rect 57325 1040 57355 1070
rect 57325 1020 57330 1040
rect 57350 1020 57355 1040
rect 57325 990 57355 1020
rect 57325 970 57330 990
rect 57350 970 57355 990
rect 57325 960 57355 970
rect 57380 1190 57410 1200
rect 57380 1170 57385 1190
rect 57405 1170 57410 1190
rect 57380 1140 57410 1170
rect 57380 1120 57385 1140
rect 57405 1120 57410 1140
rect 57380 1090 57410 1120
rect 57380 1070 57385 1090
rect 57405 1070 57410 1090
rect 57380 1040 57410 1070
rect 57380 1020 57385 1040
rect 57405 1020 57410 1040
rect 57380 990 57410 1020
rect 57380 970 57385 990
rect 57405 970 57410 990
rect 57380 960 57410 970
rect 57435 1190 57465 1200
rect 57435 1170 57440 1190
rect 57460 1170 57465 1190
rect 57435 1140 57465 1170
rect 57435 1120 57440 1140
rect 57460 1120 57465 1140
rect 57435 1090 57465 1120
rect 57435 1070 57440 1090
rect 57460 1070 57465 1090
rect 57435 1040 57465 1070
rect 57435 1020 57440 1040
rect 57460 1020 57465 1040
rect 57435 990 57465 1020
rect 57435 970 57440 990
rect 57460 970 57465 990
rect 57435 960 57465 970
rect 57490 1190 57520 1200
rect 57490 1170 57495 1190
rect 57515 1170 57520 1190
rect 57490 1140 57520 1170
rect 57490 1120 57495 1140
rect 57515 1120 57520 1140
rect 57490 1090 57520 1120
rect 57490 1070 57495 1090
rect 57515 1070 57520 1090
rect 57490 1040 57520 1070
rect 57490 1020 57495 1040
rect 57515 1020 57520 1040
rect 57490 990 57520 1020
rect 57490 970 57495 990
rect 57515 970 57520 990
rect 57490 960 57520 970
rect 57545 1190 57575 1200
rect 57545 1170 57550 1190
rect 57570 1170 57575 1190
rect 57545 1140 57575 1170
rect 57545 1120 57550 1140
rect 57570 1120 57575 1140
rect 57545 1090 57575 1120
rect 57545 1070 57550 1090
rect 57570 1070 57575 1090
rect 57545 1040 57575 1070
rect 57545 1020 57550 1040
rect 57570 1020 57575 1040
rect 57545 990 57575 1020
rect 57545 970 57550 990
rect 57570 970 57575 990
rect 57545 960 57575 970
rect 57615 1100 57635 1280
rect 56230 940 56250 960
rect 56285 940 56305 960
rect 56395 940 56415 960
rect 56505 940 56525 960
rect 56615 940 56635 960
rect 56725 940 56745 960
rect 56835 940 56855 960
rect 56945 940 56965 960
rect 57055 940 57075 960
rect 57165 940 57185 960
rect 57275 940 57295 960
rect 57385 940 57405 960
rect 57495 940 57515 960
rect 57550 940 57570 960
rect 56210 930 56250 940
rect 56210 910 56220 930
rect 56240 910 56250 930
rect 56210 900 56250 910
rect 56275 930 56315 940
rect 56275 910 56285 930
rect 56305 910 56315 930
rect 56275 900 56315 910
rect 56385 930 56425 940
rect 56385 910 56395 930
rect 56415 910 56425 930
rect 56385 900 56425 910
rect 56495 930 56535 940
rect 56495 910 56505 930
rect 56525 910 56535 930
rect 56495 900 56535 910
rect 56605 930 56645 940
rect 56605 910 56615 930
rect 56635 910 56645 930
rect 56605 900 56645 910
rect 56715 930 56755 940
rect 56715 910 56725 930
rect 56745 910 56755 930
rect 56715 900 56755 910
rect 56825 930 56865 940
rect 56825 910 56835 930
rect 56855 910 56865 930
rect 56825 900 56865 910
rect 56935 930 56975 940
rect 56935 910 56945 930
rect 56965 910 56975 930
rect 56935 900 56975 910
rect 57045 930 57085 940
rect 57045 910 57055 930
rect 57075 910 57085 930
rect 57045 900 57085 910
rect 57155 930 57195 940
rect 57155 910 57165 930
rect 57185 910 57195 930
rect 57155 900 57195 910
rect 57265 930 57305 940
rect 57265 910 57275 930
rect 57295 910 57305 930
rect 57265 900 57305 910
rect 57375 930 57415 940
rect 57375 910 57385 930
rect 57405 910 57415 930
rect 57375 900 57415 910
rect 57485 930 57525 940
rect 57485 910 57495 930
rect 57515 910 57525 930
rect 57485 900 57525 910
rect 57545 930 57585 940
rect 57545 910 57555 930
rect 57575 910 57585 930
rect 57545 900 57585 910
rect 56220 875 56240 900
rect 57555 875 57575 900
rect 57615 875 57635 1020
rect 56170 855 56860 875
rect 56940 855 57440 875
rect 57520 855 57635 875
rect 58075 1010 58095 1395
rect 58135 1375 58155 1395
rect 58735 1375 58755 1395
rect 54985 525 55315 545
rect 55395 525 55725 545
rect 56660 765 56865 785
rect 56935 765 57135 785
rect 56660 695 56680 765
rect 56755 735 56795 745
rect 56755 725 56765 735
rect 56725 715 56765 725
rect 56785 715 56795 735
rect 56725 705 56795 715
rect 56875 735 56915 745
rect 56875 715 56885 735
rect 56905 715 56915 735
rect 56875 705 56915 715
rect 56995 735 57035 745
rect 56995 715 57005 735
rect 57025 715 57035 735
rect 56995 705 57035 715
rect 57055 735 57095 745
rect 57055 715 57065 735
rect 57085 715 57095 735
rect 57055 705 57095 715
rect 56725 685 56745 705
rect 57055 685 57075 705
rect 56660 555 56680 615
rect 56715 675 56745 685
rect 56715 655 56720 675
rect 56740 655 56745 675
rect 56715 625 56745 655
rect 56715 605 56720 625
rect 56740 605 56745 625
rect 56715 595 56745 605
rect 57045 675 57075 685
rect 57045 655 57050 675
rect 57070 655 57075 675
rect 57045 625 57075 655
rect 57045 605 57050 625
rect 57070 605 57075 625
rect 57045 595 57075 605
rect 57115 695 57135 765
rect 57115 555 57135 615
rect 56660 535 56865 555
rect 56935 535 57135 555
rect 58075 545 58095 930
rect 58130 1365 58160 1375
rect 58130 1345 58135 1365
rect 58155 1345 58160 1365
rect 58130 1305 58160 1345
rect 58225 1365 58265 1375
rect 58225 1345 58235 1365
rect 58255 1345 58265 1365
rect 58225 1335 58265 1345
rect 58328 1365 58362 1375
rect 58328 1345 58336 1365
rect 58354 1345 58362 1365
rect 58328 1335 58362 1345
rect 58425 1365 58465 1375
rect 58425 1345 58435 1365
rect 58455 1345 58465 1365
rect 58425 1335 58465 1345
rect 58625 1365 58665 1375
rect 58625 1345 58635 1365
rect 58655 1345 58665 1365
rect 58625 1335 58665 1345
rect 58730 1365 58760 1375
rect 58730 1345 58735 1365
rect 58755 1345 58760 1365
rect 58235 1315 58255 1335
rect 58435 1315 58455 1335
rect 58635 1315 58655 1335
rect 58130 1285 58135 1305
rect 58155 1285 58160 1305
rect 58130 1255 58160 1285
rect 58130 1235 58135 1255
rect 58155 1235 58160 1255
rect 58130 1205 58160 1235
rect 58130 1185 58135 1205
rect 58155 1185 58160 1205
rect 58130 1155 58160 1185
rect 58130 1135 58135 1155
rect 58155 1135 58160 1155
rect 58130 1105 58160 1135
rect 58130 1085 58135 1105
rect 58155 1085 58160 1105
rect 58130 1055 58160 1085
rect 58130 1035 58135 1055
rect 58155 1035 58160 1055
rect 58130 1005 58160 1035
rect 58130 985 58135 1005
rect 58155 985 58160 1005
rect 58130 955 58160 985
rect 58130 935 58135 955
rect 58155 935 58160 955
rect 58130 905 58160 935
rect 58130 885 58135 905
rect 58155 885 58160 905
rect 58130 855 58160 885
rect 58130 835 58135 855
rect 58155 835 58160 855
rect 58130 805 58160 835
rect 58130 785 58135 805
rect 58155 785 58160 805
rect 58130 755 58160 785
rect 58130 735 58135 755
rect 58155 735 58160 755
rect 58130 705 58160 735
rect 58130 685 58135 705
rect 58155 685 58160 705
rect 58130 655 58160 685
rect 58130 635 58135 655
rect 58155 635 58160 655
rect 58130 625 58160 635
rect 58230 1305 58260 1315
rect 58230 1285 58235 1305
rect 58255 1285 58260 1305
rect 58230 1255 58260 1285
rect 58230 1235 58235 1255
rect 58255 1235 58260 1255
rect 58230 1205 58260 1235
rect 58230 1185 58235 1205
rect 58255 1185 58260 1205
rect 58230 1155 58260 1185
rect 58230 1135 58235 1155
rect 58255 1135 58260 1155
rect 58230 1105 58260 1135
rect 58230 1085 58235 1105
rect 58255 1085 58260 1105
rect 58230 1055 58260 1085
rect 58230 1035 58235 1055
rect 58255 1035 58260 1055
rect 58230 1005 58260 1035
rect 58230 985 58235 1005
rect 58255 985 58260 1005
rect 58230 955 58260 985
rect 58230 935 58235 955
rect 58255 935 58260 955
rect 58230 905 58260 935
rect 58230 885 58235 905
rect 58255 885 58260 905
rect 58230 855 58260 885
rect 58230 835 58235 855
rect 58255 835 58260 855
rect 58230 805 58260 835
rect 58230 785 58235 805
rect 58255 785 58260 805
rect 58230 755 58260 785
rect 58230 735 58235 755
rect 58255 735 58260 755
rect 58230 705 58260 735
rect 58230 685 58235 705
rect 58255 685 58260 705
rect 58230 655 58260 685
rect 58230 635 58235 655
rect 58255 635 58260 655
rect 58230 625 58260 635
rect 58330 1305 58360 1315
rect 58330 1285 58335 1305
rect 58355 1285 58360 1305
rect 58330 1255 58360 1285
rect 58330 1235 58335 1255
rect 58355 1235 58360 1255
rect 58330 1205 58360 1235
rect 58330 1185 58335 1205
rect 58355 1185 58360 1205
rect 58330 1155 58360 1185
rect 58330 1135 58335 1155
rect 58355 1135 58360 1155
rect 58330 1105 58360 1135
rect 58330 1085 58335 1105
rect 58355 1085 58360 1105
rect 58330 1055 58360 1085
rect 58330 1035 58335 1055
rect 58355 1035 58360 1055
rect 58330 1005 58360 1035
rect 58330 985 58335 1005
rect 58355 985 58360 1005
rect 58330 955 58360 985
rect 58330 935 58335 955
rect 58355 935 58360 955
rect 58330 905 58360 935
rect 58330 885 58335 905
rect 58355 885 58360 905
rect 58330 855 58360 885
rect 58330 835 58335 855
rect 58355 835 58360 855
rect 58330 805 58360 835
rect 58330 785 58335 805
rect 58355 785 58360 805
rect 58330 755 58360 785
rect 58330 735 58335 755
rect 58355 735 58360 755
rect 58330 705 58360 735
rect 58330 685 58335 705
rect 58355 685 58360 705
rect 58330 655 58360 685
rect 58330 635 58335 655
rect 58355 635 58360 655
rect 58330 625 58360 635
rect 58430 1305 58460 1315
rect 58430 1285 58435 1305
rect 58455 1285 58460 1305
rect 58430 1255 58460 1285
rect 58430 1235 58435 1255
rect 58455 1235 58460 1255
rect 58430 1205 58460 1235
rect 58430 1185 58435 1205
rect 58455 1185 58460 1205
rect 58430 1155 58460 1185
rect 58430 1135 58435 1155
rect 58455 1135 58460 1155
rect 58430 1105 58460 1135
rect 58430 1085 58435 1105
rect 58455 1085 58460 1105
rect 58430 1055 58460 1085
rect 58430 1035 58435 1055
rect 58455 1035 58460 1055
rect 58430 1005 58460 1035
rect 58430 985 58435 1005
rect 58455 985 58460 1005
rect 58430 955 58460 985
rect 58430 935 58435 955
rect 58455 935 58460 955
rect 58430 905 58460 935
rect 58430 885 58435 905
rect 58455 885 58460 905
rect 58430 855 58460 885
rect 58430 835 58435 855
rect 58455 835 58460 855
rect 58430 805 58460 835
rect 58430 785 58435 805
rect 58455 785 58460 805
rect 58430 755 58460 785
rect 58430 735 58435 755
rect 58455 735 58460 755
rect 58430 705 58460 735
rect 58430 685 58435 705
rect 58455 685 58460 705
rect 58430 655 58460 685
rect 58430 635 58435 655
rect 58455 635 58460 655
rect 58430 625 58460 635
rect 58530 1305 58560 1315
rect 58530 1285 58535 1305
rect 58555 1285 58560 1305
rect 58530 1255 58560 1285
rect 58530 1235 58535 1255
rect 58555 1235 58560 1255
rect 58530 1205 58560 1235
rect 58530 1185 58535 1205
rect 58555 1185 58560 1205
rect 58530 1155 58560 1185
rect 58530 1135 58535 1155
rect 58555 1135 58560 1155
rect 58530 1105 58560 1135
rect 58530 1085 58535 1105
rect 58555 1085 58560 1105
rect 58530 1055 58560 1085
rect 58530 1035 58535 1055
rect 58555 1035 58560 1055
rect 58530 1005 58560 1035
rect 58530 985 58535 1005
rect 58555 985 58560 1005
rect 58530 955 58560 985
rect 58530 935 58535 955
rect 58555 935 58560 955
rect 58530 905 58560 935
rect 58530 885 58535 905
rect 58555 885 58560 905
rect 58530 855 58560 885
rect 58530 835 58535 855
rect 58555 835 58560 855
rect 58530 805 58560 835
rect 58530 785 58535 805
rect 58555 785 58560 805
rect 58530 755 58560 785
rect 58530 735 58535 755
rect 58555 735 58560 755
rect 58530 705 58560 735
rect 58530 685 58535 705
rect 58555 685 58560 705
rect 58530 655 58560 685
rect 58530 635 58535 655
rect 58555 635 58560 655
rect 58530 625 58560 635
rect 58630 1305 58660 1315
rect 58630 1285 58635 1305
rect 58655 1285 58660 1305
rect 58630 1255 58660 1285
rect 58630 1235 58635 1255
rect 58655 1235 58660 1255
rect 58630 1205 58660 1235
rect 58630 1185 58635 1205
rect 58655 1185 58660 1205
rect 58630 1155 58660 1185
rect 58630 1135 58635 1155
rect 58655 1135 58660 1155
rect 58630 1105 58660 1135
rect 58630 1085 58635 1105
rect 58655 1085 58660 1105
rect 58630 1055 58660 1085
rect 58630 1035 58635 1055
rect 58655 1035 58660 1055
rect 58630 1005 58660 1035
rect 58630 985 58635 1005
rect 58655 985 58660 1005
rect 58630 955 58660 985
rect 58630 935 58635 955
rect 58655 935 58660 955
rect 58630 905 58660 935
rect 58630 885 58635 905
rect 58655 885 58660 905
rect 58630 855 58660 885
rect 58630 835 58635 855
rect 58655 835 58660 855
rect 58630 805 58660 835
rect 58630 785 58635 805
rect 58655 785 58660 805
rect 58630 755 58660 785
rect 58630 735 58635 755
rect 58655 735 58660 755
rect 58630 705 58660 735
rect 58630 685 58635 705
rect 58655 685 58660 705
rect 58630 655 58660 685
rect 58630 635 58635 655
rect 58655 635 58660 655
rect 58630 625 58660 635
rect 58730 1305 58760 1345
rect 58730 1285 58735 1305
rect 58755 1285 58760 1305
rect 58730 1255 58760 1285
rect 58730 1235 58735 1255
rect 58755 1235 58760 1255
rect 58730 1205 58760 1235
rect 58730 1185 58735 1205
rect 58755 1185 58760 1205
rect 58730 1155 58760 1185
rect 58730 1135 58735 1155
rect 58755 1135 58760 1155
rect 58730 1105 58760 1135
rect 58730 1085 58735 1105
rect 58755 1085 58760 1105
rect 58730 1055 58760 1085
rect 58730 1035 58735 1055
rect 58755 1035 58760 1055
rect 58730 1005 58760 1035
rect 58730 985 58735 1005
rect 58755 985 58760 1005
rect 58730 955 58760 985
rect 58730 935 58735 955
rect 58755 935 58760 955
rect 58730 905 58760 935
rect 58730 885 58735 905
rect 58755 885 58760 905
rect 58730 855 58760 885
rect 58730 835 58735 855
rect 58755 835 58760 855
rect 58730 805 58760 835
rect 58730 785 58735 805
rect 58755 785 58760 805
rect 58730 755 58760 785
rect 58730 735 58735 755
rect 58755 735 58760 755
rect 58730 705 58760 735
rect 58730 685 58735 705
rect 58755 685 58760 705
rect 58730 655 58760 685
rect 58730 635 58735 655
rect 58755 635 58760 655
rect 58730 625 58760 635
rect 58795 1010 58815 1395
rect 58905 1340 58985 1360
rect 59065 1340 59140 1360
rect 58905 990 58925 1340
rect 58975 1305 59010 1315
rect 58975 1280 58980 1305
rect 59005 1280 59010 1305
rect 58975 1270 59010 1280
rect 59035 1305 59070 1315
rect 59035 1280 59040 1305
rect 59065 1280 59070 1305
rect 59035 1270 59070 1280
rect 58815 980 58835 990
rect 58825 960 58835 980
rect 58815 950 58835 960
rect 58885 980 58925 990
rect 58885 960 58895 980
rect 58915 965 58925 980
rect 58885 950 58905 960
rect 58335 605 58355 625
rect 58535 605 58555 625
rect 58325 595 58365 605
rect 58325 575 58335 595
rect 58355 575 58365 595
rect 58325 565 58365 575
rect 58525 595 58565 605
rect 58525 575 58535 595
rect 58555 575 58565 595
rect 58525 565 58565 575
rect 58795 545 58815 930
rect 56875 525 56885 535
rect 56905 525 56915 535
rect 58075 525 58405 545
rect 58485 525 58815 545
rect 58905 533 58925 885
rect 59120 965 59140 1340
rect 59010 583 59035 633
rect 59120 533 59140 885
rect 55335 515 55345 525
rect 55365 515 55375 525
rect 56875 515 56915 525
rect 58425 515 58435 525
rect 58455 515 58465 525
rect 55335 505 55375 515
rect 58425 505 58465 515
rect 58905 513 58985 533
rect 59065 513 59140 533
<< viali >>
rect 56830 4760 56850 4780
rect 56890 4760 56910 4780
rect 56950 4760 56970 4780
rect 57010 4760 57030 4780
rect 56155 4505 56175 4525
rect 56215 4505 56235 4525
rect 56335 4505 56355 4525
rect 56245 4370 56265 4390
rect 56920 4365 56940 4385
rect 57500 4800 57520 4820
rect 57560 4800 57580 4820
rect 57680 4800 57700 4820
rect 57577 4365 57595 4385
rect 57625 4370 57645 4390
rect 55085 4065 55105 4085
rect 55205 4065 55225 4085
rect 55325 4065 55345 4085
rect 55445 4065 55465 4085
rect 55565 4065 55585 4085
rect 55025 3645 55045 3665
rect 55145 3645 55165 3665
rect 55265 3645 55285 3665
rect 55326 3645 55344 3665
rect 55385 3645 55405 3665
rect 55505 3645 55525 3665
rect 55625 3645 55645 3665
rect 56135 4065 56155 4085
rect 56255 4065 56275 4085
rect 56375 4065 56395 4085
rect 56495 4065 56515 4085
rect 56615 4065 56635 4085
rect 56075 3645 56095 3665
rect 56195 3645 56215 3665
rect 56315 3645 56335 3665
rect 56376 3645 56394 3665
rect 56435 3645 56455 3665
rect 56555 3645 56575 3665
rect 56675 3645 56695 3665
rect 57165 4065 57185 4085
rect 57285 4065 57305 4085
rect 57405 4065 57425 4085
rect 57525 4065 57545 4085
rect 57645 4065 57665 4085
rect 57105 3645 57125 3665
rect 57225 3645 57245 3665
rect 57345 3645 57365 3665
rect 57406 3645 57424 3665
rect 57465 3645 57485 3665
rect 57585 3645 57605 3665
rect 57705 3645 57725 3665
rect 58215 4065 58235 4085
rect 58335 4065 58355 4085
rect 58455 4065 58475 4085
rect 58575 4065 58595 4085
rect 58695 4065 58715 4085
rect 58155 3645 58175 3665
rect 58275 3645 58295 3665
rect 58395 3645 58415 3665
rect 58456 3645 58474 3665
rect 58515 3645 58535 3665
rect 58635 3645 58655 3665
rect 58755 3645 58775 3665
rect 54560 3290 54590 3320
rect 54610 3290 54640 3320
rect 54659 3290 54689 3320
rect 54560 2685 54590 2715
rect 54610 2685 54640 2715
rect 54659 2685 54689 2715
rect 54535 2630 54555 2650
rect 54965 3355 54985 3375
rect 55075 3355 55095 3375
rect 55185 3355 55205 3375
rect 55295 3355 55315 3375
rect 55405 3355 55425 3375
rect 55515 3355 55535 3375
rect 55625 3355 55645 3375
rect 55020 2685 55040 2705
rect 55130 2685 55150 2705
rect 55186 2685 55204 2705
rect 55240 2685 55260 2705
rect 55350 2685 55370 2705
rect 55460 2685 55480 2705
rect 55570 2685 55590 2705
rect 56285 3355 56305 3375
rect 56395 3355 56415 3375
rect 56505 3355 56525 3375
rect 56615 3355 56635 3375
rect 56725 3355 56745 3375
rect 56835 3355 56855 3375
rect 56945 3355 56965 3375
rect 57055 3355 57075 3375
rect 57165 3355 57185 3375
rect 57275 3355 57295 3375
rect 57385 3355 57405 3375
rect 57495 3355 57515 3375
rect 56340 3235 56360 3255
rect 56450 3235 56470 3255
rect 56505 3235 56525 3255
rect 56560 3235 56580 3255
rect 56670 3235 56690 3255
rect 56780 3235 56800 3255
rect 56890 3235 56910 3255
rect 57000 3235 57020 3255
rect 57110 3235 57130 3255
rect 57220 3235 57240 3255
rect 57330 3235 57350 3255
rect 57440 3235 57460 3255
rect 58155 3355 58175 3375
rect 58265 3355 58285 3375
rect 58375 3355 58395 3375
rect 58485 3355 58505 3375
rect 58595 3355 58615 3375
rect 58705 3355 58725 3375
rect 58815 3355 58835 3375
rect 56150 2900 56170 2920
rect 56195 2900 56215 2920
rect 56295 2900 56315 2920
rect 56350 2900 56370 2920
rect 56405 2900 56425 2920
rect 56460 2900 56480 2920
rect 56515 2900 56535 2920
rect 56570 2900 56590 2920
rect 56625 2900 56645 2920
rect 56015 2840 56035 2860
rect 56130 2780 56150 2800
rect 56225 2780 56245 2800
rect 56278 2780 56295 2800
rect 56350 2780 56370 2800
rect 56445 2780 56465 2800
rect 56498 2780 56515 2800
rect 56570 2780 56590 2800
rect 56645 2780 56662 2800
rect 56688 2780 56708 2800
rect 57118 2900 57138 2920
rect 57165 2900 57185 2920
rect 57265 2900 57285 2920
rect 57320 2900 57340 2920
rect 57375 2900 57395 2920
rect 57485 2900 57505 2920
rect 57540 2900 57560 2920
rect 57595 2900 57615 2920
rect 56795 2840 56815 2860
rect 56985 2840 57005 2860
rect 57100 2780 57120 2800
rect 57195 2780 57215 2800
rect 57248 2780 57265 2800
rect 57320 2780 57340 2800
rect 57415 2780 57435 2800
rect 57468 2780 57485 2800
rect 57540 2780 57560 2800
rect 57615 2780 57632 2800
rect 57658 2780 57678 2800
rect 55295 2635 55315 2645
rect 58210 2685 58230 2705
rect 58320 2685 58340 2705
rect 58430 2685 58450 2705
rect 58540 2685 58560 2705
rect 58596 2685 58614 2705
rect 58650 2685 58670 2705
rect 58760 2685 58780 2705
rect 58485 2635 58505 2645
rect 59111 3290 59141 3320
rect 59160 3290 59190 3320
rect 59210 3290 59240 3320
rect 59111 2685 59141 2715
rect 59160 2685 59190 2715
rect 59210 2685 59240 2715
rect 55295 2625 55315 2635
rect 58485 2625 58505 2635
rect 59245 2630 59265 2650
rect 55295 2465 55315 2475
rect 55295 2455 55315 2465
rect 54535 2300 54555 2310
rect 55020 2395 55040 2415
rect 55130 2395 55150 2415
rect 55240 2395 55260 2415
rect 55350 2395 55370 2415
rect 55460 2395 55480 2415
rect 55570 2395 55590 2415
rect 54535 2290 54555 2300
rect 55075 2125 55095 2145
rect 55185 2125 55205 2145
rect 55295 2125 55315 2145
rect 55405 2125 55425 2145
rect 55461 2125 55479 2145
rect 55515 2125 55535 2145
rect 56615 2485 56635 2505
rect 56725 2485 56745 2505
rect 56835 2485 56855 2505
rect 56945 2485 56965 2505
rect 57055 2485 57075 2505
rect 57165 2485 57185 2505
rect 58485 2465 58505 2475
rect 56670 2365 56690 2385
rect 56780 2365 56800 2385
rect 56890 2365 56910 2385
rect 57000 2365 57020 2385
rect 57110 2365 57130 2385
rect 56890 2315 56910 2325
rect 58485 2455 58505 2465
rect 56890 2305 56910 2315
rect 58210 2395 58230 2415
rect 58320 2395 58340 2415
rect 58430 2395 58450 2415
rect 58540 2395 58560 2415
rect 58650 2395 58670 2415
rect 58760 2395 58780 2415
rect 54475 1565 54500 1590
rect 54535 1565 54560 1590
rect 54595 1565 54620 1590
rect 54655 1565 54680 1590
rect 54745 1750 54765 1770
rect 54895 1750 54905 1770
rect 54905 1750 54915 1770
rect 55075 1935 55095 1955
rect 55185 1935 55205 1955
rect 55295 1935 55315 1955
rect 55405 1935 55425 1955
rect 55461 1935 55479 1955
rect 55515 1935 55535 1955
rect 56140 2205 56160 2225
rect 56250 2205 56270 2225
rect 56360 2205 56380 2225
rect 56415 2205 56435 2225
rect 56470 2205 56490 2225
rect 56580 2205 56600 2225
rect 56690 2205 56710 2225
rect 56805 2095 56825 2115
rect 56195 1985 56215 2005
rect 56305 1985 56325 2005
rect 56415 1985 56435 2005
rect 56525 1985 56545 2005
rect 56635 1985 56655 2005
rect 56975 2095 56995 2115
rect 57090 2205 57110 2225
rect 57200 2205 57220 2225
rect 57310 2205 57330 2225
rect 57365 2205 57385 2225
rect 57420 2205 57440 2225
rect 57530 2205 57550 2225
rect 57640 2205 57660 2225
rect 58265 2125 58285 2145
rect 58321 2125 58339 2145
rect 58375 2125 58395 2145
rect 58485 2125 58505 2145
rect 58595 2125 58615 2145
rect 58705 2125 58725 2145
rect 59245 2300 59265 2310
rect 59245 2290 59265 2300
rect 57145 1985 57165 2005
rect 57255 1985 57275 2005
rect 57365 1985 57385 2005
rect 57475 1985 57495 2005
rect 57585 1985 57605 2005
rect 56890 1805 56910 1815
rect 55020 1565 55038 1585
rect 55130 1565 55148 1585
rect 55240 1565 55258 1585
rect 55350 1565 55368 1585
rect 55460 1565 55478 1585
rect 55570 1565 55588 1585
rect 55295 1515 55315 1525
rect 56890 1795 56910 1805
rect 55295 1505 55315 1515
rect 56103 1725 56123 1745
rect 56197 1725 56217 1745
rect 56243 1735 56260 1755
rect 56323 1725 56343 1745
rect 56417 1725 56437 1745
rect 56463 1735 56480 1755
rect 56543 1725 56563 1745
rect 56610 1735 56627 1755
rect 56653 1725 56673 1745
rect 56827 1735 56847 1755
rect 56873 1735 56890 1755
rect 56950 1735 56970 1755
rect 57143 1725 57163 1745
rect 57237 1725 57257 1745
rect 57283 1735 57300 1755
rect 57363 1725 57383 1745
rect 57457 1725 57477 1745
rect 57503 1735 57520 1755
rect 57583 1725 57603 1745
rect 57650 1735 57667 1755
rect 57693 1725 57713 1745
rect 57800 1625 57820 1645
rect 58095 1625 58115 1645
rect 56112 1515 56129 1535
rect 56158 1515 56178 1535
rect 56260 1515 56280 1535
rect 56315 1515 56335 1535
rect 56370 1515 56390 1535
rect 56480 1515 56500 1535
rect 56535 1515 56555 1535
rect 56590 1515 56610 1535
rect 56830 1515 56850 1535
rect 56880 1515 56900 1535
rect 56928 1515 56945 1535
rect 57152 1515 57169 1535
rect 57198 1515 57218 1535
rect 57300 1515 57320 1535
rect 57355 1515 57375 1535
rect 57410 1515 57430 1535
rect 57520 1515 57540 1535
rect 57575 1515 57595 1535
rect 57630 1515 57650 1535
rect 58265 1935 58285 1955
rect 58321 1935 58339 1955
rect 58375 1935 58395 1955
rect 58485 1935 58505 1955
rect 58595 1935 58615 1955
rect 58705 1935 58725 1955
rect 58885 1750 58895 1770
rect 58895 1750 58905 1770
rect 59035 1750 59055 1770
rect 58212 1565 58230 1585
rect 58322 1565 58340 1585
rect 58432 1565 58450 1585
rect 58542 1565 58560 1585
rect 58652 1565 58670 1585
rect 58762 1565 58780 1585
rect 58485 1515 58505 1525
rect 59120 1565 59145 1590
rect 59180 1565 59205 1590
rect 59240 1565 59265 1590
rect 59300 1565 59325 1590
rect 58485 1505 58505 1515
rect 55295 1405 55315 1425
rect 54735 1280 54760 1305
rect 54795 1280 54820 1305
rect 54885 965 54905 980
rect 54885 960 54895 965
rect 54895 960 54905 965
rect 54975 960 54985 980
rect 54985 960 54995 980
rect 55145 1345 55165 1365
rect 55345 1345 55365 1365
rect 55446 1345 55464 1365
rect 55545 1345 55565 1365
rect 58485 1405 58505 1425
rect 55245 575 55265 595
rect 55445 575 55465 595
rect 56340 1230 56360 1250
rect 56450 1230 56470 1250
rect 56560 1230 56580 1250
rect 56670 1230 56690 1250
rect 56780 1230 56800 1250
rect 56835 1230 56855 1250
rect 56890 1230 56910 1250
rect 57000 1230 57020 1250
rect 57110 1230 57130 1250
rect 57220 1230 57240 1250
rect 57330 1230 57350 1250
rect 57425 1230 57445 1250
rect 57479 1230 57499 1250
rect 56220 910 56240 930
rect 56285 910 56305 930
rect 56395 910 56415 930
rect 56505 910 56525 930
rect 56615 910 56635 930
rect 56725 910 56745 930
rect 56835 910 56855 930
rect 56945 910 56965 930
rect 57055 910 57075 930
rect 57165 910 57185 930
rect 57275 910 57295 930
rect 57385 910 57405 930
rect 57495 910 57515 930
rect 57555 910 57575 930
rect 55345 525 55365 535
rect 56765 715 56785 735
rect 56885 715 56905 735
rect 57005 715 57025 735
rect 57065 715 57085 735
rect 56885 535 56905 545
rect 58235 1345 58255 1365
rect 58336 1345 58354 1365
rect 58435 1345 58455 1365
rect 58635 1345 58655 1365
rect 58980 1280 59005 1305
rect 59040 1280 59065 1305
rect 58805 960 58815 980
rect 58815 960 58825 980
rect 58895 965 58915 980
rect 58895 960 58905 965
rect 58905 960 58915 965
rect 58335 575 58355 595
rect 58535 575 58555 595
rect 56885 525 56905 535
rect 58435 525 58455 535
rect 55345 515 55365 525
rect 58435 515 58455 525
<< metal1 >>
rect 55785 6185 55825 6190
rect 55785 6155 55790 6185
rect 55820 6155 55825 6185
rect 55785 6150 55825 6155
rect 55795 4535 55815 6150
rect 56880 4880 56920 4885
rect 56880 4850 56885 4880
rect 56915 4850 56920 4880
rect 56880 4845 56920 4850
rect 57550 4880 57590 4885
rect 57550 4850 57555 4880
rect 57585 4850 57590 4880
rect 57550 4845 57590 4850
rect 56890 4790 56910 4845
rect 57560 4830 57580 4845
rect 57490 4825 57530 4830
rect 57490 4795 57495 4825
rect 57525 4795 57530 4825
rect 57490 4790 57530 4795
rect 57550 4825 57590 4830
rect 57550 4795 57555 4825
rect 57585 4795 57590 4825
rect 57550 4790 57590 4795
rect 57670 4825 57710 4830
rect 57670 4795 57675 4825
rect 57705 4795 57710 4825
rect 57670 4790 57710 4795
rect 56325 4785 56365 4790
rect 56325 4755 56330 4785
rect 56360 4755 56365 4785
rect 56325 4750 56365 4755
rect 56820 4785 56860 4790
rect 56820 4755 56825 4785
rect 56855 4755 56860 4785
rect 56820 4750 56860 4755
rect 56887 4780 56913 4790
rect 56887 4760 56890 4780
rect 56910 4760 56913 4780
rect 56887 4750 56913 4760
rect 56940 4785 56980 4790
rect 56940 4755 56945 4785
rect 56975 4755 56980 4785
rect 56940 4750 56980 4755
rect 57000 4785 57040 4790
rect 57000 4755 57005 4785
rect 57035 4755 57040 4785
rect 57000 4750 57040 4755
rect 56335 4535 56355 4750
rect 55785 4530 55825 4535
rect 55785 4500 55790 4530
rect 55820 4500 55825 4530
rect 55785 4495 55825 4500
rect 56145 4530 56185 4535
rect 56145 4500 56150 4530
rect 56180 4500 56185 4530
rect 56145 4495 56185 4500
rect 56205 4530 56245 4535
rect 56205 4500 56210 4530
rect 56240 4500 56245 4530
rect 56205 4495 56245 4500
rect 56325 4530 56365 4535
rect 56325 4500 56330 4530
rect 56360 4500 56365 4530
rect 56325 4495 56365 4500
rect 55795 4205 55815 4495
rect 56235 4390 56275 4400
rect 57620 4395 57650 4400
rect 56235 4370 56245 4390
rect 56265 4370 56275 4390
rect 56235 4360 56275 4370
rect 56910 4390 56950 4395
rect 56910 4360 56915 4390
rect 56945 4360 56950 4390
rect 56245 4295 56265 4360
rect 56910 4355 56950 4360
rect 57571 4385 57603 4395
rect 57571 4365 57577 4385
rect 57595 4365 57603 4385
rect 57571 4355 57603 4365
rect 57620 4360 57650 4365
rect 56235 4290 56275 4295
rect 56235 4260 56240 4290
rect 56270 4260 56275 4290
rect 56235 4255 56275 4260
rect 56850 4290 56890 4295
rect 56850 4260 56855 4290
rect 56885 4260 56890 4290
rect 56850 4255 56890 4260
rect 55315 4200 55355 4205
rect 55315 4170 55320 4200
rect 55350 4170 55355 4200
rect 55315 4165 55355 4170
rect 55785 4200 55825 4205
rect 55785 4170 55790 4200
rect 55820 4170 55825 4200
rect 55785 4165 55825 4170
rect 55325 4095 55345 4165
rect 55075 4090 55115 4095
rect 55075 4060 55080 4090
rect 55110 4060 55115 4090
rect 55075 4055 55115 4060
rect 55195 4090 55235 4095
rect 55195 4060 55200 4090
rect 55230 4060 55235 4090
rect 55195 4055 55235 4060
rect 55315 4090 55355 4095
rect 55315 4060 55320 4090
rect 55350 4060 55355 4090
rect 55315 4055 55355 4060
rect 55435 4090 55475 4095
rect 55435 4060 55440 4090
rect 55470 4060 55475 4090
rect 55435 4055 55475 4060
rect 55555 4090 55595 4095
rect 55555 4060 55560 4090
rect 55590 4060 55595 4090
rect 55555 4055 55595 4060
rect 55015 3670 55055 3675
rect 55015 3640 55020 3670
rect 55050 3640 55055 3670
rect 55015 3635 55055 3640
rect 55135 3670 55175 3675
rect 55135 3640 55140 3670
rect 55170 3640 55175 3670
rect 55135 3635 55175 3640
rect 55255 3670 55295 3675
rect 55255 3640 55260 3670
rect 55290 3640 55295 3670
rect 55255 3635 55295 3640
rect 55318 3665 55352 3675
rect 55318 3645 55326 3665
rect 55344 3645 55352 3665
rect 55318 3635 55352 3645
rect 55375 3670 55415 3675
rect 55375 3640 55380 3670
rect 55410 3640 55415 3670
rect 55375 3635 55415 3640
rect 55495 3670 55535 3675
rect 55495 3640 55500 3670
rect 55530 3640 55535 3670
rect 55495 3635 55535 3640
rect 55615 3670 55655 3675
rect 55615 3640 55620 3670
rect 55650 3640 55655 3670
rect 55615 3635 55655 3640
rect 55325 3575 55345 3635
rect 55315 3570 55355 3575
rect 55315 3540 55320 3570
rect 55350 3540 55355 3570
rect 55315 3535 55355 3540
rect 54605 3400 54645 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 55795 3385 55815 4165
rect 55890 4090 55930 4095
rect 55890 4060 55895 4090
rect 55925 4060 55930 4090
rect 55890 4055 55930 4060
rect 56125 4090 56165 4095
rect 56125 4060 56130 4090
rect 56160 4060 56165 4090
rect 56125 4055 56165 4060
rect 56185 4090 56225 4095
rect 56185 4060 56190 4090
rect 56220 4060 56225 4090
rect 56185 4055 56225 4060
rect 56245 4090 56285 4095
rect 56245 4060 56250 4090
rect 56280 4060 56285 4090
rect 56245 4055 56285 4060
rect 56365 4090 56405 4095
rect 56365 4060 56370 4090
rect 56400 4060 56405 4090
rect 56365 4055 56405 4060
rect 56485 4090 56525 4095
rect 56485 4060 56490 4090
rect 56520 4060 56525 4090
rect 56485 4055 56525 4060
rect 56605 4090 56645 4095
rect 56605 4060 56610 4090
rect 56640 4060 56645 4090
rect 56605 4055 56645 4060
rect 55900 3675 55920 4055
rect 55890 3670 55930 3675
rect 55890 3640 55895 3670
rect 55925 3640 55930 3670
rect 55890 3635 55930 3640
rect 56065 3670 56105 3675
rect 56065 3640 56070 3670
rect 56100 3640 56105 3670
rect 56065 3635 56105 3640
rect 56185 3670 56225 3675
rect 56185 3640 56190 3670
rect 56220 3640 56225 3670
rect 56185 3635 56225 3640
rect 56305 3670 56345 3675
rect 56305 3640 56310 3670
rect 56340 3640 56345 3670
rect 56305 3635 56345 3640
rect 56368 3665 56402 3675
rect 56368 3645 56376 3665
rect 56394 3645 56402 3665
rect 56368 3635 56402 3645
rect 56425 3670 56465 3675
rect 56425 3640 56430 3670
rect 56460 3640 56465 3670
rect 56425 3635 56465 3640
rect 56545 3670 56585 3675
rect 56545 3640 56550 3670
rect 56580 3640 56585 3670
rect 56545 3635 56585 3640
rect 56665 3670 56705 3675
rect 56665 3640 56670 3670
rect 56700 3640 56705 3670
rect 56665 3635 56705 3640
rect 54605 3365 54645 3370
rect 54955 3380 54995 3385
rect 54615 3325 54635 3365
rect 54955 3350 54960 3380
rect 54990 3350 54995 3380
rect 54955 3345 54995 3350
rect 55065 3380 55105 3385
rect 55065 3350 55070 3380
rect 55100 3350 55105 3380
rect 55065 3345 55105 3350
rect 55175 3380 55215 3385
rect 55175 3350 55180 3380
rect 55210 3350 55215 3380
rect 55175 3345 55215 3350
rect 55285 3380 55325 3385
rect 55285 3350 55290 3380
rect 55320 3350 55325 3380
rect 55285 3345 55325 3350
rect 55395 3380 55435 3385
rect 55395 3350 55400 3380
rect 55430 3350 55435 3380
rect 55395 3345 55435 3350
rect 55505 3380 55545 3385
rect 55505 3350 55510 3380
rect 55540 3350 55545 3380
rect 55505 3345 55545 3350
rect 55615 3380 55655 3385
rect 55615 3350 55620 3380
rect 55650 3350 55655 3380
rect 55615 3345 55655 3350
rect 55785 3380 55825 3385
rect 55785 3350 55790 3380
rect 55820 3350 55825 3380
rect 55785 3345 55825 3350
rect 55740 3325 55780 3330
rect 54554 3320 54695 3325
rect 54554 3290 54560 3320
rect 54590 3290 54610 3320
rect 54640 3290 54659 3320
rect 54689 3290 54695 3320
rect 55740 3295 55745 3325
rect 55775 3295 55780 3325
rect 55740 3290 55780 3295
rect 54554 3285 54695 3290
rect 54554 2715 54695 2720
rect 54554 2685 54560 2715
rect 54590 2685 54610 2715
rect 54640 2685 54659 2715
rect 54689 2685 54695 2715
rect 54554 2680 54695 2685
rect 55010 2710 55050 2715
rect 55010 2680 55015 2710
rect 55045 2680 55050 2710
rect 54525 2650 54565 2660
rect 54525 2630 54535 2650
rect 54555 2630 54565 2650
rect 54525 2620 54565 2630
rect 54315 2545 54355 2550
rect 54315 2515 54320 2545
rect 54350 2515 54355 2545
rect 54315 2510 54355 2515
rect 54265 2420 54305 2425
rect 54265 2390 54270 2420
rect 54300 2390 54305 2420
rect 54265 2385 54305 2390
rect 54275 500 54295 2385
rect 54325 1920 54345 2510
rect 54535 2320 54555 2620
rect 54615 2595 54635 2680
rect 55010 2675 55050 2680
rect 55120 2710 55160 2715
rect 55120 2680 55125 2710
rect 55155 2680 55160 2710
rect 55120 2675 55160 2680
rect 55178 2705 55212 2715
rect 55178 2685 55186 2705
rect 55204 2685 55212 2705
rect 55178 2675 55212 2685
rect 55230 2710 55270 2715
rect 55230 2680 55235 2710
rect 55265 2680 55270 2710
rect 55230 2675 55270 2680
rect 55340 2710 55380 2715
rect 55340 2680 55345 2710
rect 55375 2680 55380 2710
rect 55340 2675 55380 2680
rect 55450 2710 55490 2715
rect 55450 2680 55455 2710
rect 55485 2680 55490 2710
rect 55450 2675 55490 2680
rect 55560 2710 55600 2715
rect 55560 2680 55565 2710
rect 55595 2680 55600 2710
rect 55560 2675 55600 2680
rect 55185 2595 55205 2675
rect 55285 2645 55325 2655
rect 55285 2625 55295 2645
rect 55315 2625 55325 2645
rect 55285 2615 55325 2625
rect 54605 2590 54645 2595
rect 54605 2560 54610 2590
rect 54640 2560 54645 2590
rect 54605 2555 54645 2560
rect 55175 2590 55215 2595
rect 55175 2560 55180 2590
rect 55210 2560 55215 2590
rect 55175 2555 55215 2560
rect 55295 2485 55315 2615
rect 55460 2550 55480 2675
rect 55750 2595 55770 3290
rect 55795 2870 55815 3345
rect 56075 3330 56095 3635
rect 56375 3620 56395 3635
rect 56860 3620 56880 4255
rect 56365 3615 56405 3620
rect 56365 3585 56370 3615
rect 56400 3585 56405 3615
rect 56365 3580 56405 3585
rect 56850 3615 56890 3620
rect 56850 3585 56855 3615
rect 56885 3585 56890 3615
rect 56850 3580 56890 3585
rect 56920 3575 56940 4355
rect 57575 4295 57595 4355
rect 57565 4290 57605 4295
rect 57565 4260 57570 4290
rect 57600 4260 57605 4290
rect 57565 4255 57605 4260
rect 57975 4200 58015 4205
rect 57975 4170 57980 4200
rect 58010 4170 58015 4200
rect 57975 4165 58015 4170
rect 58445 4200 58485 4205
rect 58445 4170 58450 4200
rect 58480 4170 58485 4200
rect 58445 4165 58485 4170
rect 57155 4090 57195 4095
rect 57155 4060 57160 4090
rect 57190 4060 57195 4090
rect 57155 4055 57195 4060
rect 57275 4090 57315 4095
rect 57275 4060 57280 4090
rect 57310 4060 57315 4090
rect 57275 4055 57315 4060
rect 57395 4090 57435 4095
rect 57395 4060 57400 4090
rect 57430 4060 57435 4090
rect 57395 4055 57435 4060
rect 57515 4090 57555 4095
rect 57515 4060 57520 4090
rect 57550 4060 57555 4090
rect 57515 4055 57555 4060
rect 57575 4090 57615 4095
rect 57575 4060 57580 4090
rect 57610 4060 57615 4090
rect 57575 4055 57615 4060
rect 57635 4090 57675 4095
rect 57635 4060 57640 4090
rect 57670 4060 57675 4090
rect 57635 4055 57675 4060
rect 57870 4090 57910 4095
rect 57870 4060 57875 4090
rect 57905 4060 57910 4090
rect 57870 4055 57910 4060
rect 57880 3675 57900 4055
rect 57095 3670 57135 3675
rect 57095 3640 57100 3670
rect 57130 3640 57135 3670
rect 57095 3635 57135 3640
rect 57215 3670 57255 3675
rect 57215 3640 57220 3670
rect 57250 3640 57255 3670
rect 57215 3635 57255 3640
rect 57335 3670 57375 3675
rect 57335 3640 57340 3670
rect 57370 3640 57375 3670
rect 57335 3635 57375 3640
rect 57398 3665 57432 3675
rect 57398 3645 57406 3665
rect 57424 3645 57432 3665
rect 57398 3635 57432 3645
rect 57455 3670 57495 3675
rect 57455 3640 57460 3670
rect 57490 3640 57495 3670
rect 57455 3635 57495 3640
rect 57575 3670 57615 3675
rect 57575 3640 57580 3670
rect 57610 3640 57615 3670
rect 57575 3635 57615 3640
rect 57695 3670 57735 3675
rect 57695 3640 57700 3670
rect 57730 3640 57735 3670
rect 57695 3635 57735 3640
rect 57870 3670 57910 3675
rect 57870 3640 57875 3670
rect 57905 3640 57910 3670
rect 57870 3635 57910 3640
rect 57405 3620 57425 3635
rect 57395 3615 57435 3620
rect 57395 3585 57400 3615
rect 57430 3585 57435 3615
rect 57395 3580 57435 3585
rect 56910 3570 56950 3575
rect 56910 3540 56915 3570
rect 56945 3540 56950 3570
rect 56910 3535 56950 3540
rect 57985 3385 58005 4165
rect 58455 4095 58475 4165
rect 58205 4090 58245 4095
rect 58205 4060 58210 4090
rect 58240 4060 58245 4090
rect 58205 4055 58245 4060
rect 58325 4090 58365 4095
rect 58325 4060 58330 4090
rect 58360 4060 58365 4090
rect 58325 4055 58365 4060
rect 58445 4090 58485 4095
rect 58445 4060 58450 4090
rect 58480 4060 58485 4090
rect 58445 4055 58485 4060
rect 58565 4090 58605 4095
rect 58565 4060 58570 4090
rect 58600 4060 58605 4090
rect 58565 4055 58605 4060
rect 58685 4090 58725 4095
rect 58685 4060 58690 4090
rect 58720 4060 58725 4090
rect 58685 4055 58725 4060
rect 58145 3670 58185 3675
rect 58145 3640 58150 3670
rect 58180 3640 58185 3670
rect 58145 3635 58185 3640
rect 58265 3670 58305 3675
rect 58265 3640 58270 3670
rect 58300 3640 58305 3670
rect 58265 3635 58305 3640
rect 58385 3670 58425 3675
rect 58385 3640 58390 3670
rect 58420 3640 58425 3670
rect 58385 3635 58425 3640
rect 58448 3665 58482 3675
rect 58448 3645 58456 3665
rect 58474 3645 58482 3665
rect 58448 3635 58482 3645
rect 58505 3670 58545 3675
rect 58505 3640 58510 3670
rect 58540 3640 58545 3670
rect 58505 3635 58545 3640
rect 58625 3670 58665 3675
rect 58625 3640 58630 3670
rect 58660 3640 58665 3670
rect 58625 3635 58665 3640
rect 58745 3670 58785 3675
rect 58745 3640 58750 3670
rect 58780 3640 58785 3670
rect 58745 3635 58785 3640
rect 58455 3575 58475 3635
rect 58445 3570 58485 3575
rect 58445 3540 58450 3570
rect 58480 3540 58485 3570
rect 59155 3400 59195 3405
rect 56275 3380 56315 3385
rect 56275 3350 56280 3380
rect 56310 3350 56315 3380
rect 56275 3345 56315 3350
rect 56385 3380 56425 3385
rect 56385 3350 56390 3380
rect 56420 3350 56425 3380
rect 56385 3345 56425 3350
rect 56495 3380 56535 3385
rect 56495 3350 56500 3380
rect 56530 3350 56535 3380
rect 56495 3345 56535 3350
rect 56605 3380 56645 3385
rect 56605 3350 56610 3380
rect 56640 3350 56645 3380
rect 56605 3345 56645 3350
rect 56715 3380 56755 3385
rect 56715 3350 56720 3380
rect 56750 3350 56755 3380
rect 56715 3345 56755 3350
rect 56825 3380 56865 3385
rect 56825 3350 56830 3380
rect 56860 3350 56865 3380
rect 56825 3345 56865 3350
rect 56935 3380 56975 3385
rect 56935 3350 56940 3380
rect 56970 3350 56975 3380
rect 56935 3345 56975 3350
rect 57045 3380 57085 3385
rect 57045 3350 57050 3380
rect 57080 3350 57085 3380
rect 57045 3345 57085 3350
rect 57155 3380 57195 3385
rect 57155 3350 57160 3380
rect 57190 3350 57195 3380
rect 57155 3345 57195 3350
rect 57265 3380 57305 3385
rect 57265 3350 57270 3380
rect 57300 3350 57305 3380
rect 57265 3345 57305 3350
rect 57375 3380 57415 3385
rect 57375 3350 57380 3380
rect 57410 3350 57415 3380
rect 57375 3345 57415 3350
rect 57485 3380 57525 3385
rect 57485 3350 57490 3380
rect 57520 3350 57525 3380
rect 57485 3345 57525 3350
rect 57975 3380 58015 3385
rect 57975 3350 57980 3380
rect 58010 3350 58015 3380
rect 57975 3345 58015 3350
rect 58145 3380 58185 3385
rect 58145 3350 58150 3380
rect 58180 3350 58185 3380
rect 58145 3345 58185 3350
rect 58255 3380 58295 3385
rect 58255 3350 58260 3380
rect 58290 3350 58295 3380
rect 58255 3345 58295 3350
rect 58365 3380 58405 3385
rect 58365 3350 58370 3380
rect 58400 3350 58405 3380
rect 58365 3345 58405 3350
rect 58475 3380 58515 3385
rect 58475 3350 58480 3380
rect 58510 3350 58515 3380
rect 58475 3345 58515 3350
rect 58585 3380 58625 3385
rect 58585 3350 58590 3380
rect 58620 3350 58625 3380
rect 58585 3345 58625 3350
rect 58695 3380 58735 3385
rect 58695 3350 58700 3380
rect 58730 3350 58735 3380
rect 58695 3345 58735 3350
rect 58805 3380 58845 3385
rect 58805 3350 58810 3380
rect 58840 3350 58845 3380
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58805 3345 58845 3350
rect 56065 3325 56105 3330
rect 56065 3295 56070 3325
rect 56100 3295 56105 3325
rect 56065 3290 56105 3295
rect 56330 3260 56370 3265
rect 56330 3230 56335 3260
rect 56365 3230 56370 3260
rect 56330 3225 56370 3230
rect 56440 3255 56480 3265
rect 56440 3235 56450 3255
rect 56470 3235 56480 3255
rect 56440 3225 56480 3235
rect 56497 3255 56533 3265
rect 56497 3235 56505 3255
rect 56525 3235 56533 3255
rect 56497 3225 56533 3235
rect 56550 3260 56590 3265
rect 56550 3230 56555 3260
rect 56585 3230 56590 3260
rect 56550 3225 56590 3230
rect 56660 3255 56700 3265
rect 56660 3235 56670 3255
rect 56690 3235 56700 3255
rect 56660 3225 56700 3235
rect 56770 3260 56810 3265
rect 56770 3230 56775 3260
rect 56805 3230 56810 3260
rect 56770 3225 56810 3230
rect 56880 3255 56920 3265
rect 56880 3235 56890 3255
rect 56910 3235 56920 3255
rect 56880 3225 56920 3235
rect 56990 3260 57030 3265
rect 56990 3230 56995 3260
rect 57025 3230 57030 3260
rect 56990 3225 57030 3230
rect 57100 3255 57140 3265
rect 57100 3235 57110 3255
rect 57130 3235 57140 3255
rect 57100 3225 57140 3235
rect 57190 3260 57250 3265
rect 57190 3230 57215 3260
rect 57245 3230 57250 3260
rect 57190 3225 57250 3230
rect 57320 3255 57360 3265
rect 57320 3235 57330 3255
rect 57350 3235 57360 3255
rect 57320 3225 57360 3235
rect 57430 3260 57470 3265
rect 57430 3230 57435 3260
rect 57465 3230 57470 3260
rect 57430 3225 57470 3230
rect 56450 3210 56470 3225
rect 56440 3205 56480 3210
rect 56440 3175 56445 3205
rect 56475 3175 56480 3205
rect 56440 3170 56480 3175
rect 56505 3050 56525 3225
rect 56670 3210 56690 3225
rect 56890 3210 56910 3225
rect 57110 3210 57130 3225
rect 56465 3045 56525 3050
rect 56465 3015 56480 3045
rect 56510 3015 56525 3045
rect 56465 3010 56525 3015
rect 56640 3205 56700 3210
rect 56640 3175 56665 3205
rect 56695 3175 56700 3205
rect 56640 3170 56700 3175
rect 56880 3205 56920 3210
rect 56880 3175 56885 3205
rect 56915 3175 56920 3205
rect 56880 3170 56920 3175
rect 57100 3205 57140 3210
rect 57100 3175 57105 3205
rect 57135 3175 57140 3205
rect 57100 3170 57140 3175
rect 56185 2985 56225 2990
rect 56185 2955 56190 2985
rect 56220 2955 56225 2985
rect 56185 2950 56225 2955
rect 56285 2985 56325 2990
rect 56285 2955 56290 2985
rect 56320 2955 56325 2985
rect 56285 2950 56325 2955
rect 56395 2985 56435 2990
rect 56395 2955 56400 2985
rect 56430 2955 56435 2985
rect 56395 2950 56435 2955
rect 56195 2930 56215 2950
rect 56295 2930 56315 2950
rect 56405 2930 56425 2950
rect 56465 2930 56485 3010
rect 56640 2990 56660 3170
rect 57190 2990 57210 3225
rect 57330 3210 57350 3225
rect 57320 3205 57360 3210
rect 57320 3175 57325 3205
rect 57355 3175 57360 3205
rect 57320 3170 57360 3175
rect 56505 2985 56545 2990
rect 56505 2955 56510 2985
rect 56540 2955 56545 2985
rect 56505 2950 56545 2955
rect 56615 2985 56660 2990
rect 56615 2955 56620 2985
rect 56650 2955 56660 2985
rect 56615 2950 56660 2955
rect 57155 2985 57210 2990
rect 57155 2955 57160 2985
rect 57190 2955 57210 2985
rect 57155 2950 57210 2955
rect 57255 2985 57295 2990
rect 57255 2955 57260 2985
rect 57290 2955 57295 2985
rect 57255 2950 57295 2955
rect 57365 2985 57405 2990
rect 57365 2955 57370 2985
rect 57400 2955 57405 2985
rect 57365 2950 57405 2955
rect 57475 2985 57515 2990
rect 57475 2955 57480 2985
rect 57510 2955 57515 2985
rect 57475 2950 57515 2955
rect 57585 2985 57625 2990
rect 57585 2955 57590 2985
rect 57620 2955 57625 2985
rect 57585 2950 57625 2955
rect 56515 2930 56535 2950
rect 56625 2930 56645 2950
rect 57165 2930 57185 2950
rect 57265 2930 57285 2950
rect 57375 2930 57395 2950
rect 57485 2930 57505 2950
rect 57595 2930 57615 2950
rect 56145 2924 56175 2930
rect 56145 2896 56147 2924
rect 56173 2896 56175 2924
rect 56145 2890 56175 2896
rect 56192 2920 56218 2930
rect 56192 2900 56195 2920
rect 56215 2900 56218 2920
rect 56192 2890 56218 2900
rect 56292 2920 56318 2930
rect 56292 2900 56295 2920
rect 56315 2900 56318 2920
rect 56292 2890 56318 2900
rect 56345 2924 56375 2930
rect 56345 2896 56347 2924
rect 56373 2896 56375 2924
rect 56345 2890 56375 2896
rect 56402 2920 56428 2930
rect 56402 2900 56405 2920
rect 56425 2900 56428 2920
rect 56402 2890 56428 2900
rect 56455 2920 56485 2930
rect 56455 2900 56460 2920
rect 56480 2900 56485 2920
rect 56455 2890 56485 2900
rect 56512 2920 56538 2930
rect 56512 2900 56515 2920
rect 56535 2900 56538 2920
rect 56512 2890 56538 2900
rect 56560 2925 56600 2930
rect 56560 2895 56565 2925
rect 56595 2895 56600 2925
rect 56560 2890 56600 2895
rect 56622 2920 56648 2930
rect 56622 2900 56625 2920
rect 56645 2900 56648 2920
rect 56622 2890 56648 2900
rect 56880 2925 56920 2930
rect 56880 2895 56885 2925
rect 56915 2895 56920 2925
rect 56880 2890 56920 2895
rect 57113 2924 57143 2930
rect 57113 2896 57115 2924
rect 57141 2896 57143 2924
rect 57113 2890 57143 2896
rect 57162 2920 57188 2930
rect 57162 2900 57165 2920
rect 57185 2900 57188 2920
rect 57162 2890 57188 2900
rect 57262 2920 57288 2930
rect 57262 2900 57265 2920
rect 57285 2900 57288 2920
rect 57262 2890 57288 2900
rect 57310 2925 57350 2930
rect 57310 2895 57315 2925
rect 57345 2895 57350 2925
rect 57310 2890 57350 2895
rect 57372 2920 57398 2930
rect 57372 2900 57375 2920
rect 57395 2900 57398 2920
rect 57372 2890 57398 2900
rect 57482 2920 57508 2930
rect 57482 2900 57485 2920
rect 57505 2900 57508 2920
rect 57482 2890 57508 2900
rect 57530 2925 57570 2930
rect 57530 2895 57535 2925
rect 57565 2895 57570 2925
rect 57530 2890 57570 2895
rect 57592 2920 57618 2930
rect 57592 2900 57595 2920
rect 57615 2900 57618 2920
rect 57592 2890 57618 2900
rect 55785 2865 55825 2870
rect 55785 2835 55790 2865
rect 55820 2835 55825 2865
rect 55785 2830 55825 2835
rect 56005 2865 56045 2870
rect 56005 2835 56010 2865
rect 56040 2835 56045 2865
rect 56005 2830 56045 2835
rect 56785 2865 56825 2870
rect 56785 2835 56790 2865
rect 56820 2835 56825 2865
rect 56785 2830 56825 2835
rect 55740 2590 55780 2595
rect 55740 2560 55745 2590
rect 55775 2560 55780 2590
rect 55740 2555 55780 2560
rect 55450 2545 55490 2550
rect 55450 2515 55455 2545
rect 55485 2515 55490 2545
rect 55450 2510 55490 2515
rect 55285 2475 55325 2485
rect 55285 2455 55295 2475
rect 55315 2455 55325 2475
rect 55285 2445 55325 2455
rect 55010 2420 55050 2425
rect 55010 2390 55015 2420
rect 55045 2390 55050 2420
rect 55010 2385 55050 2390
rect 55120 2420 55160 2425
rect 55120 2390 55125 2420
rect 55155 2390 55160 2420
rect 55120 2385 55160 2390
rect 55230 2420 55270 2425
rect 55230 2390 55235 2420
rect 55265 2390 55270 2420
rect 55230 2385 55270 2390
rect 55340 2420 55380 2425
rect 55340 2390 55345 2420
rect 55375 2390 55380 2420
rect 55340 2385 55380 2390
rect 55450 2420 55490 2425
rect 55450 2390 55455 2420
rect 55485 2390 55490 2420
rect 55450 2385 55490 2390
rect 55560 2420 55600 2425
rect 55560 2390 55565 2420
rect 55595 2390 55600 2420
rect 55560 2385 55600 2390
rect 54525 2310 54565 2320
rect 54525 2290 54535 2310
rect 54555 2290 54565 2310
rect 54525 2280 54565 2290
rect 54790 2150 54830 2155
rect 54790 2120 54795 2150
rect 54825 2120 54830 2150
rect 54790 2115 54830 2120
rect 55065 2150 55105 2155
rect 55065 2120 55070 2150
rect 55100 2120 55105 2150
rect 55065 2115 55105 2120
rect 55175 2150 55215 2155
rect 55175 2120 55180 2150
rect 55210 2120 55215 2150
rect 55175 2115 55215 2120
rect 55285 2150 55325 2155
rect 55285 2120 55290 2150
rect 55320 2120 55325 2150
rect 55285 2115 55325 2120
rect 55395 2150 55435 2155
rect 55395 2120 55400 2150
rect 55430 2120 55435 2150
rect 55395 2115 55435 2120
rect 55453 2145 55487 2155
rect 55453 2125 55461 2145
rect 55479 2125 55487 2145
rect 55453 2115 55487 2125
rect 55505 2150 55545 2155
rect 55505 2120 55510 2150
rect 55540 2120 55545 2150
rect 55505 2115 55545 2120
rect 54310 1910 54360 1920
rect 54310 1880 54320 1910
rect 54350 1880 54360 1910
rect 54310 1870 54360 1880
rect 54325 1375 54345 1870
rect 54735 1775 54775 1780
rect 54735 1745 54740 1775
rect 54770 1745 54775 1775
rect 54735 1740 54775 1745
rect 54470 1595 54505 1600
rect 54470 1555 54505 1560
rect 54530 1595 54565 1600
rect 54530 1555 54565 1560
rect 54590 1595 54625 1601
rect 54590 1555 54625 1560
rect 54650 1595 54685 1600
rect 54650 1555 54685 1560
rect 54480 1490 54500 1555
rect 54600 1540 54620 1555
rect 54800 1540 54820 2115
rect 55460 2050 55480 2115
rect 55750 2050 55770 2555
rect 55450 2045 55490 2050
rect 55450 2015 55455 2045
rect 55485 2015 55490 2045
rect 55450 2010 55490 2015
rect 55740 2045 55780 2050
rect 55740 2015 55745 2045
rect 55775 2015 55780 2045
rect 55740 2010 55780 2015
rect 55460 1965 55480 2010
rect 54835 1960 54875 1965
rect 54835 1930 54840 1960
rect 54870 1930 54875 1960
rect 54835 1925 54875 1930
rect 55065 1960 55105 1965
rect 55065 1930 55070 1960
rect 55100 1930 55105 1960
rect 55065 1925 55105 1930
rect 55175 1960 55215 1965
rect 55175 1930 55180 1960
rect 55210 1930 55215 1960
rect 55175 1925 55215 1930
rect 55285 1960 55325 1965
rect 55285 1930 55290 1960
rect 55320 1930 55325 1960
rect 55285 1925 55325 1930
rect 55395 1960 55435 1965
rect 55395 1930 55400 1960
rect 55430 1930 55435 1960
rect 55395 1925 55435 1930
rect 55453 1955 55487 1965
rect 55453 1935 55461 1955
rect 55479 1935 55487 1955
rect 55453 1925 55487 1935
rect 55505 1960 55545 1965
rect 55505 1930 55510 1960
rect 55540 1930 55545 1960
rect 55505 1925 55545 1930
rect 54845 1595 54865 1925
rect 54885 1775 54925 1780
rect 54885 1745 54890 1775
rect 54920 1745 54925 1775
rect 54885 1740 54925 1745
rect 55795 1595 55815 2830
rect 56120 2800 56160 2810
rect 56120 2780 56130 2800
rect 56150 2780 56160 2800
rect 56120 2770 56160 2780
rect 56215 2800 56255 2810
rect 56215 2780 56225 2800
rect 56245 2780 56255 2800
rect 56215 2770 56255 2780
rect 56272 2805 56304 2810
rect 56272 2775 56275 2805
rect 56301 2775 56304 2805
rect 56272 2770 56304 2775
rect 56340 2800 56380 2810
rect 56340 2780 56350 2800
rect 56370 2780 56380 2800
rect 56340 2770 56380 2780
rect 56435 2800 56475 2810
rect 56435 2780 56445 2800
rect 56465 2780 56475 2800
rect 56435 2770 56475 2780
rect 56492 2805 56524 2810
rect 56492 2775 56495 2805
rect 56521 2775 56524 2805
rect 56492 2770 56524 2775
rect 56560 2800 56600 2810
rect 56560 2780 56570 2800
rect 56590 2780 56600 2800
rect 56560 2770 56600 2780
rect 56636 2805 56668 2810
rect 56636 2775 56639 2805
rect 56665 2775 56668 2805
rect 56636 2770 56668 2775
rect 56685 2800 56711 2810
rect 56685 2780 56688 2800
rect 56708 2780 56711 2800
rect 56685 2770 56711 2780
rect 56130 2750 56150 2770
rect 56235 2750 56255 2770
rect 56350 2750 56370 2770
rect 56455 2750 56475 2770
rect 56570 2750 56590 2770
rect 56685 2750 56705 2770
rect 56120 2745 56160 2750
rect 56120 2715 56125 2745
rect 56155 2715 56160 2745
rect 56120 2710 56160 2715
rect 56225 2745 56265 2750
rect 56225 2715 56230 2745
rect 56260 2715 56265 2745
rect 56225 2710 56265 2715
rect 56340 2745 56380 2750
rect 56340 2715 56345 2745
rect 56375 2715 56380 2745
rect 56340 2710 56380 2715
rect 56445 2745 56485 2750
rect 56445 2715 56450 2745
rect 56480 2715 56485 2745
rect 56445 2710 56485 2715
rect 56560 2745 56600 2750
rect 56560 2715 56565 2745
rect 56595 2715 56600 2745
rect 56560 2710 56600 2715
rect 56675 2745 56715 2750
rect 56675 2715 56680 2745
rect 56710 2715 56715 2745
rect 56675 2710 56715 2715
rect 56605 2690 56645 2695
rect 56605 2660 56610 2690
rect 56640 2660 56645 2690
rect 56605 2655 56645 2660
rect 55875 2645 55915 2650
rect 55875 2615 55880 2645
rect 55910 2615 55915 2645
rect 55875 2610 55915 2615
rect 55830 2230 55870 2235
rect 55830 2200 55835 2230
rect 55865 2200 55870 2230
rect 55830 2195 55870 2200
rect 54835 1590 54875 1595
rect 54835 1560 54840 1590
rect 54870 1560 54875 1590
rect 54835 1555 54875 1560
rect 55010 1590 55050 1595
rect 55010 1560 55015 1590
rect 55045 1560 55050 1590
rect 55010 1555 55050 1560
rect 55120 1590 55160 1595
rect 55120 1560 55125 1590
rect 55155 1560 55160 1590
rect 55120 1555 55160 1560
rect 55230 1590 55270 1595
rect 55230 1560 55235 1590
rect 55265 1560 55270 1590
rect 55230 1555 55270 1560
rect 55340 1590 55380 1595
rect 55340 1560 55345 1590
rect 55375 1560 55380 1590
rect 55340 1555 55380 1560
rect 55450 1590 55490 1595
rect 55450 1560 55455 1590
rect 55485 1560 55490 1590
rect 55450 1555 55490 1560
rect 55560 1590 55600 1595
rect 55560 1560 55565 1590
rect 55595 1560 55600 1590
rect 55560 1555 55600 1560
rect 55785 1590 55825 1595
rect 55785 1560 55790 1590
rect 55820 1560 55825 1590
rect 55785 1555 55825 1560
rect 54590 1535 54630 1540
rect 54590 1505 54595 1535
rect 54625 1505 54630 1535
rect 54590 1500 54630 1505
rect 54790 1535 54830 1540
rect 54790 1505 54795 1535
rect 54825 1505 54830 1535
rect 54790 1500 54830 1505
rect 55285 1525 55325 1535
rect 55285 1505 55295 1525
rect 55315 1505 55325 1525
rect 55285 1495 55325 1505
rect 54470 1485 54510 1490
rect 54470 1455 54475 1485
rect 54505 1455 54510 1485
rect 54470 1450 54510 1455
rect 55295 1435 55315 1495
rect 54725 1425 54765 1430
rect 54725 1395 54730 1425
rect 54760 1395 54765 1425
rect 55285 1425 55325 1435
rect 55285 1405 55295 1425
rect 55315 1405 55325 1425
rect 55285 1395 55325 1405
rect 55435 1425 55475 1430
rect 55435 1395 55440 1425
rect 55470 1395 55475 1425
rect 54725 1390 54765 1395
rect 55435 1390 55475 1395
rect 55740 1425 55780 1430
rect 55740 1395 55745 1425
rect 55775 1395 55780 1425
rect 55740 1390 55780 1395
rect 54315 1370 54355 1375
rect 54315 1340 54320 1370
rect 54350 1340 54355 1370
rect 54315 1335 54355 1340
rect 54735 1315 54755 1390
rect 55445 1375 55465 1390
rect 54790 1370 54830 1375
rect 54790 1340 54795 1370
rect 54825 1340 54830 1370
rect 54790 1335 54830 1340
rect 55135 1370 55175 1375
rect 55135 1340 55140 1370
rect 55170 1340 55175 1370
rect 55135 1335 55175 1340
rect 55335 1370 55375 1375
rect 55335 1340 55340 1370
rect 55370 1340 55375 1370
rect 55335 1335 55375 1340
rect 55438 1365 55472 1375
rect 55438 1345 55446 1365
rect 55464 1345 55472 1365
rect 55438 1335 55472 1345
rect 55535 1370 55575 1375
rect 55535 1340 55540 1370
rect 55570 1340 55575 1370
rect 55535 1335 55575 1340
rect 54800 1315 54820 1335
rect 54730 1310 54765 1315
rect 54730 1270 54765 1275
rect 54790 1310 54825 1315
rect 54790 1270 54825 1275
rect 54875 985 54915 990
rect 54875 955 54880 985
rect 54910 955 54915 985
rect 54875 950 54915 955
rect 54965 985 55005 990
rect 54965 955 54970 985
rect 55000 955 55005 985
rect 54965 950 55005 955
rect 55785 935 55825 940
rect 55785 905 55790 935
rect 55820 905 55825 935
rect 55785 900 55825 905
rect 55795 605 55815 900
rect 55840 745 55860 2195
rect 55885 1490 55905 2610
rect 56240 2590 56280 2595
rect 56240 2560 56245 2590
rect 56275 2560 56280 2590
rect 56240 2555 56280 2560
rect 56250 2290 56270 2555
rect 56615 2515 56635 2655
rect 56890 2650 56910 2890
rect 56975 2865 57015 2870
rect 56975 2835 56980 2865
rect 57010 2835 57015 2865
rect 56975 2830 57015 2835
rect 57090 2800 57130 2810
rect 57090 2780 57100 2800
rect 57120 2780 57130 2800
rect 57090 2770 57130 2780
rect 57185 2800 57225 2810
rect 57185 2780 57195 2800
rect 57215 2780 57225 2800
rect 57185 2770 57225 2780
rect 57242 2805 57274 2810
rect 57242 2775 57245 2805
rect 57271 2775 57274 2805
rect 57242 2770 57274 2775
rect 57310 2800 57350 2810
rect 57310 2780 57320 2800
rect 57340 2780 57350 2800
rect 57310 2770 57350 2780
rect 57405 2800 57445 2810
rect 57405 2780 57415 2800
rect 57435 2780 57445 2800
rect 57405 2770 57445 2780
rect 57462 2805 57494 2810
rect 57462 2775 57465 2805
rect 57491 2775 57494 2805
rect 57462 2770 57494 2775
rect 57530 2800 57570 2810
rect 57530 2780 57540 2800
rect 57560 2780 57570 2800
rect 57530 2770 57570 2780
rect 57606 2805 57638 2810
rect 57606 2775 57609 2805
rect 57635 2775 57638 2805
rect 57606 2770 57638 2775
rect 57655 2800 57681 2810
rect 57655 2780 57658 2800
rect 57678 2780 57681 2800
rect 57655 2770 57681 2780
rect 57100 2750 57120 2770
rect 57090 2745 57130 2750
rect 57090 2715 57095 2745
rect 57125 2715 57130 2745
rect 57090 2710 57130 2715
rect 56880 2645 56920 2650
rect 56880 2615 56885 2645
rect 56915 2615 56920 2645
rect 56880 2610 56920 2615
rect 57100 2605 57120 2710
rect 57195 2695 57215 2770
rect 57320 2750 57340 2770
rect 57310 2745 57350 2750
rect 57310 2715 57315 2745
rect 57345 2715 57350 2745
rect 57310 2710 57350 2715
rect 57415 2695 57435 2770
rect 57540 2750 57560 2770
rect 57530 2745 57570 2750
rect 57530 2715 57535 2745
rect 57565 2715 57570 2745
rect 57530 2710 57570 2715
rect 57655 2695 57675 2770
rect 57185 2690 57225 2695
rect 57185 2660 57190 2690
rect 57220 2660 57225 2690
rect 57185 2655 57225 2660
rect 57405 2690 57445 2695
rect 57405 2660 57410 2690
rect 57440 2660 57445 2690
rect 57405 2655 57445 2660
rect 57645 2690 57685 2695
rect 57645 2660 57650 2690
rect 57680 2660 57685 2690
rect 57645 2655 57685 2660
rect 57870 2645 57910 2650
rect 57870 2615 57875 2645
rect 57905 2615 57910 2645
rect 57870 2610 57910 2615
rect 56715 2600 56755 2605
rect 56715 2570 56720 2600
rect 56750 2570 56755 2600
rect 56715 2565 56755 2570
rect 56935 2600 56975 2605
rect 56935 2570 56940 2600
rect 56970 2570 56975 2600
rect 56935 2565 56975 2570
rect 57090 2600 57130 2605
rect 57090 2570 57095 2600
rect 57125 2570 57130 2600
rect 57090 2565 57130 2570
rect 57155 2600 57195 2605
rect 57155 2570 57160 2600
rect 57190 2570 57195 2600
rect 57155 2565 57195 2570
rect 57520 2590 57560 2595
rect 56725 2515 56745 2565
rect 56945 2515 56965 2565
rect 57165 2515 57185 2565
rect 57520 2560 57525 2590
rect 57555 2560 57560 2590
rect 57520 2555 57560 2560
rect 56605 2510 56645 2515
rect 56605 2480 56610 2510
rect 56640 2480 56645 2510
rect 56605 2475 56645 2480
rect 56715 2505 56755 2515
rect 56715 2485 56725 2505
rect 56745 2485 56755 2505
rect 56715 2475 56755 2485
rect 56825 2510 56865 2515
rect 56825 2480 56830 2510
rect 56860 2480 56865 2510
rect 56825 2475 56865 2480
rect 56935 2505 56975 2515
rect 56935 2485 56945 2505
rect 56965 2485 56975 2505
rect 56935 2475 56975 2485
rect 57045 2510 57085 2515
rect 57045 2480 57050 2510
rect 57080 2480 57085 2510
rect 57045 2475 57085 2480
rect 57155 2505 57195 2515
rect 57155 2485 57165 2505
rect 57185 2485 57195 2505
rect 57155 2475 57195 2485
rect 56660 2390 56700 2395
rect 56660 2360 56665 2390
rect 56695 2360 56700 2390
rect 56660 2355 56700 2360
rect 56770 2390 56810 2395
rect 56770 2360 56775 2390
rect 56805 2360 56810 2390
rect 56770 2355 56810 2360
rect 56880 2390 56920 2395
rect 56880 2360 56885 2390
rect 56915 2360 56920 2390
rect 56880 2355 56920 2360
rect 56990 2390 57030 2395
rect 56990 2360 56995 2390
rect 57025 2360 57030 2390
rect 56990 2355 57030 2360
rect 57100 2390 57140 2395
rect 57100 2360 57105 2390
rect 57135 2360 57140 2390
rect 57100 2355 57140 2360
rect 56880 2330 56920 2335
rect 56880 2300 56885 2330
rect 56915 2300 56920 2330
rect 56880 2295 56920 2300
rect 56130 2285 56170 2290
rect 56130 2255 56135 2285
rect 56165 2255 56170 2285
rect 56130 2250 56170 2255
rect 56240 2285 56280 2290
rect 56240 2255 56245 2285
rect 56275 2255 56280 2285
rect 56240 2250 56280 2255
rect 56350 2285 56390 2290
rect 56350 2255 56355 2285
rect 56385 2255 56390 2285
rect 56350 2250 56390 2255
rect 56460 2285 56500 2290
rect 56460 2255 56465 2285
rect 56495 2255 56500 2285
rect 56460 2250 56500 2255
rect 56570 2285 56610 2290
rect 56570 2255 56575 2285
rect 56605 2255 56610 2285
rect 56570 2250 56610 2255
rect 56680 2285 56720 2290
rect 56680 2255 56685 2285
rect 56715 2255 56720 2285
rect 56680 2250 56720 2255
rect 56140 2235 56160 2250
rect 56250 2235 56270 2250
rect 56360 2235 56380 2250
rect 56470 2235 56490 2250
rect 56580 2235 56600 2250
rect 56690 2235 56710 2250
rect 56130 2225 56170 2235
rect 56130 2205 56140 2225
rect 56160 2205 56170 2225
rect 56130 2195 56170 2205
rect 56240 2225 56280 2235
rect 56240 2205 56250 2225
rect 56270 2205 56280 2225
rect 56240 2195 56280 2205
rect 56350 2225 56390 2235
rect 56350 2205 56360 2225
rect 56380 2205 56390 2225
rect 56350 2195 56390 2205
rect 56410 2230 56440 2235
rect 56410 2195 56440 2200
rect 56460 2225 56500 2235
rect 56460 2205 56470 2225
rect 56490 2205 56500 2225
rect 56460 2195 56500 2205
rect 56570 2225 56610 2235
rect 56570 2205 56580 2225
rect 56600 2205 56610 2225
rect 56570 2195 56610 2205
rect 56680 2225 56720 2235
rect 56680 2205 56690 2225
rect 56710 2205 56720 2225
rect 56680 2195 56720 2205
rect 56890 2125 56910 2295
rect 57530 2290 57550 2555
rect 57080 2285 57120 2290
rect 57080 2255 57085 2285
rect 57115 2255 57120 2285
rect 57080 2250 57120 2255
rect 57190 2285 57230 2290
rect 57190 2255 57195 2285
rect 57225 2255 57230 2285
rect 57190 2250 57230 2255
rect 57300 2285 57340 2290
rect 57300 2255 57305 2285
rect 57335 2255 57340 2285
rect 57300 2250 57340 2255
rect 57410 2285 57450 2290
rect 57410 2255 57415 2285
rect 57445 2255 57450 2285
rect 57410 2250 57450 2255
rect 57520 2285 57560 2290
rect 57520 2255 57525 2285
rect 57555 2255 57560 2285
rect 57520 2250 57560 2255
rect 57630 2285 57670 2290
rect 57630 2255 57635 2285
rect 57665 2255 57670 2285
rect 57630 2250 57670 2255
rect 57090 2235 57110 2250
rect 57200 2235 57220 2250
rect 57310 2235 57330 2250
rect 57420 2235 57440 2250
rect 57530 2235 57550 2250
rect 57640 2235 57660 2250
rect 57080 2225 57120 2235
rect 57080 2205 57090 2225
rect 57110 2205 57120 2225
rect 57080 2195 57120 2205
rect 57190 2225 57230 2235
rect 57190 2205 57200 2225
rect 57220 2205 57230 2225
rect 57190 2195 57230 2205
rect 57300 2225 57340 2235
rect 57300 2205 57310 2225
rect 57330 2205 57340 2225
rect 57300 2195 57340 2205
rect 57360 2230 57390 2235
rect 57360 2195 57390 2200
rect 57410 2225 57450 2235
rect 57410 2205 57420 2225
rect 57440 2205 57450 2225
rect 57410 2195 57450 2205
rect 57520 2225 57560 2235
rect 57520 2205 57530 2225
rect 57550 2205 57560 2225
rect 57520 2195 57560 2205
rect 57630 2225 57670 2235
rect 57630 2205 57640 2225
rect 57660 2205 57670 2225
rect 57630 2195 57670 2205
rect 56795 2120 56835 2125
rect 56795 2090 56800 2120
rect 56830 2090 56835 2120
rect 56795 2085 56835 2090
rect 56880 2120 56920 2125
rect 56880 2090 56885 2120
rect 56915 2090 56920 2120
rect 56880 2085 56920 2090
rect 56965 2120 57005 2125
rect 56965 2090 56970 2120
rect 57000 2090 57005 2120
rect 56965 2085 57005 2090
rect 56185 2005 56225 2015
rect 56185 1985 56195 2005
rect 56215 1985 56225 2005
rect 56185 1975 56225 1985
rect 56295 2005 56335 2015
rect 56295 1985 56305 2005
rect 56325 1985 56335 2005
rect 56295 1975 56335 1985
rect 56405 2005 56445 2015
rect 56405 1985 56415 2005
rect 56435 1985 56445 2005
rect 56405 1975 56445 1985
rect 56515 2005 56555 2015
rect 56515 1985 56525 2005
rect 56545 1985 56555 2005
rect 56515 1975 56555 1985
rect 56625 2005 56665 2015
rect 56625 1985 56635 2005
rect 56655 1985 56665 2005
rect 56625 1975 56665 1985
rect 56195 1955 56215 1975
rect 56305 1955 56325 1975
rect 56415 1955 56435 1975
rect 56525 1955 56545 1975
rect 56635 1955 56655 1975
rect 56185 1950 56225 1955
rect 56185 1920 56190 1950
rect 56220 1920 56225 1950
rect 56185 1915 56225 1920
rect 56295 1950 56335 1955
rect 56295 1920 56300 1950
rect 56330 1920 56335 1950
rect 56295 1915 56335 1920
rect 56405 1950 56445 1955
rect 56405 1920 56410 1950
rect 56440 1920 56445 1950
rect 56405 1915 56445 1920
rect 56515 1950 56555 1955
rect 56515 1920 56520 1950
rect 56550 1920 56555 1950
rect 56515 1915 56555 1920
rect 56625 1950 56665 1955
rect 56625 1920 56630 1950
rect 56660 1920 56665 1950
rect 56625 1915 56665 1920
rect 56190 1895 56230 1900
rect 56190 1865 56195 1895
rect 56225 1865 56230 1895
rect 56190 1860 56230 1865
rect 56410 1895 56450 1900
rect 56410 1865 56415 1895
rect 56445 1865 56450 1895
rect 56410 1860 56450 1865
rect 56085 1805 56125 1810
rect 56085 1775 56090 1805
rect 56120 1775 56125 1805
rect 56085 1770 56125 1775
rect 56100 1755 56120 1770
rect 56200 1755 56220 1860
rect 56305 1805 56345 1810
rect 56305 1775 56310 1805
rect 56340 1775 56345 1805
rect 56305 1770 56345 1775
rect 56100 1745 56126 1755
rect 56100 1725 56103 1745
rect 56123 1725 56126 1745
rect 56100 1715 56126 1725
rect 56194 1745 56220 1755
rect 56194 1725 56197 1745
rect 56217 1725 56220 1745
rect 56237 1760 56269 1765
rect 56237 1730 56240 1760
rect 56266 1730 56269 1760
rect 56237 1725 56269 1730
rect 56320 1755 56340 1770
rect 56420 1755 56440 1860
rect 56535 1810 56555 1915
rect 56640 1895 56680 1900
rect 56640 1865 56645 1895
rect 56675 1865 56680 1895
rect 56640 1860 56680 1865
rect 56525 1805 56565 1810
rect 56525 1775 56530 1805
rect 56560 1775 56565 1805
rect 56525 1770 56565 1775
rect 56320 1745 56346 1755
rect 56320 1725 56323 1745
rect 56343 1725 56346 1745
rect 56194 1715 56220 1725
rect 56320 1715 56346 1725
rect 56414 1745 56440 1755
rect 56414 1725 56417 1745
rect 56437 1725 56440 1745
rect 56457 1760 56489 1765
rect 56457 1730 56460 1760
rect 56486 1730 56489 1760
rect 56457 1725 56489 1730
rect 56540 1755 56560 1770
rect 56601 1760 56633 1765
rect 56540 1745 56566 1755
rect 56540 1725 56543 1745
rect 56563 1725 56566 1745
rect 56601 1730 56604 1760
rect 56630 1730 56633 1760
rect 56601 1725 56633 1730
rect 56650 1755 56670 1860
rect 56820 1850 56860 1855
rect 56820 1820 56825 1850
rect 56855 1820 56860 1850
rect 56890 1825 56910 2085
rect 57135 2005 57175 2015
rect 57135 1985 57145 2005
rect 57165 1985 57175 2005
rect 57135 1975 57175 1985
rect 57245 2005 57285 2015
rect 57245 1985 57255 2005
rect 57275 1985 57285 2005
rect 57245 1975 57285 1985
rect 57355 2005 57395 2015
rect 57355 1985 57365 2005
rect 57385 1985 57395 2005
rect 57355 1975 57395 1985
rect 57465 2005 57505 2015
rect 57465 1985 57475 2005
rect 57495 1985 57505 2005
rect 57465 1975 57505 1985
rect 57575 2005 57615 2015
rect 57575 1985 57585 2005
rect 57605 1985 57615 2005
rect 57575 1975 57615 1985
rect 57145 1955 57165 1975
rect 57255 1955 57275 1975
rect 57365 1955 57385 1975
rect 57475 1955 57495 1975
rect 57585 1955 57605 1975
rect 57135 1950 57175 1955
rect 57135 1920 57140 1950
rect 57170 1920 57175 1950
rect 57135 1915 57175 1920
rect 57245 1950 57285 1955
rect 57245 1920 57250 1950
rect 57280 1920 57285 1950
rect 57245 1915 57285 1920
rect 57355 1950 57395 1955
rect 57355 1920 57360 1950
rect 57390 1920 57395 1950
rect 57355 1915 57395 1920
rect 57465 1950 57505 1955
rect 57465 1920 57470 1950
rect 57500 1920 57505 1950
rect 57465 1915 57505 1920
rect 57575 1950 57615 1955
rect 57575 1920 57580 1950
rect 57610 1920 57615 1950
rect 57575 1915 57615 1920
rect 57245 1900 57265 1915
rect 57230 1895 57270 1900
rect 57230 1865 57235 1895
rect 57265 1865 57270 1895
rect 57230 1860 57270 1865
rect 57450 1895 57490 1900
rect 57450 1865 57455 1895
rect 57485 1865 57490 1895
rect 57450 1860 57490 1865
rect 57680 1895 57720 1900
rect 57680 1865 57685 1895
rect 57715 1865 57720 1895
rect 57680 1860 57720 1865
rect 56940 1850 56980 1855
rect 56820 1815 56860 1820
rect 56880 1815 56920 1825
rect 56940 1820 56945 1850
rect 56975 1820 56980 1850
rect 56940 1815 56980 1820
rect 56830 1765 56850 1815
rect 56880 1795 56890 1815
rect 56910 1795 56920 1815
rect 56880 1785 56920 1795
rect 56950 1765 56970 1815
rect 57125 1805 57165 1810
rect 57125 1775 57130 1805
rect 57160 1775 57165 1805
rect 57125 1770 57165 1775
rect 56824 1755 56850 1765
rect 56650 1745 56676 1755
rect 56650 1725 56653 1745
rect 56673 1725 56676 1745
rect 56824 1735 56827 1755
rect 56847 1735 56850 1755
rect 56824 1725 56850 1735
rect 56867 1760 56899 1765
rect 56867 1730 56870 1760
rect 56896 1730 56899 1760
rect 56867 1725 56899 1730
rect 56947 1755 56973 1765
rect 56947 1735 56950 1755
rect 56970 1735 56973 1755
rect 56947 1725 56973 1735
rect 57140 1755 57160 1770
rect 57240 1755 57260 1860
rect 57345 1805 57385 1810
rect 57345 1775 57350 1805
rect 57380 1775 57385 1805
rect 57345 1770 57385 1775
rect 57140 1745 57166 1755
rect 57140 1725 57143 1745
rect 57163 1725 57166 1745
rect 56414 1715 56440 1725
rect 56540 1715 56566 1725
rect 56650 1715 56676 1725
rect 57140 1715 57166 1725
rect 57234 1745 57260 1755
rect 57234 1725 57237 1745
rect 57257 1725 57260 1745
rect 57277 1760 57309 1765
rect 57277 1730 57280 1760
rect 57306 1730 57309 1760
rect 57277 1725 57309 1730
rect 57360 1755 57380 1770
rect 57460 1755 57480 1860
rect 57565 1805 57605 1810
rect 57565 1775 57570 1805
rect 57600 1775 57605 1805
rect 57565 1770 57605 1775
rect 57360 1745 57386 1755
rect 57360 1725 57363 1745
rect 57383 1725 57386 1745
rect 57234 1715 57260 1725
rect 57360 1715 57386 1725
rect 57454 1745 57480 1755
rect 57454 1725 57457 1745
rect 57477 1725 57480 1745
rect 57497 1760 57529 1765
rect 57497 1730 57500 1760
rect 57526 1730 57529 1760
rect 57497 1725 57529 1730
rect 57580 1755 57600 1770
rect 57641 1760 57673 1765
rect 57580 1745 57606 1755
rect 57580 1725 57583 1745
rect 57603 1725 57606 1745
rect 57641 1730 57644 1760
rect 57670 1730 57673 1760
rect 57641 1725 57673 1730
rect 57690 1755 57710 1860
rect 57690 1745 57716 1755
rect 57690 1725 57693 1745
rect 57713 1725 57716 1745
rect 57454 1715 57480 1725
rect 57580 1715 57606 1725
rect 57690 1715 57716 1725
rect 57790 1650 57830 1655
rect 57790 1620 57795 1650
rect 57825 1620 57830 1650
rect 57790 1615 57830 1620
rect 56106 1540 56138 1545
rect 56106 1510 56109 1540
rect 56135 1510 56138 1540
rect 56106 1505 56138 1510
rect 56155 1535 56181 1545
rect 56155 1515 56158 1535
rect 56178 1515 56181 1535
rect 56155 1505 56181 1515
rect 56256 1535 56283 1545
rect 56256 1515 56260 1535
rect 56280 1515 56283 1535
rect 56256 1505 56283 1515
rect 56305 1540 56345 1545
rect 56305 1510 56310 1540
rect 56340 1510 56345 1540
rect 56305 1505 56345 1510
rect 56366 1535 56393 1545
rect 56366 1515 56370 1535
rect 56390 1515 56393 1535
rect 56366 1505 56393 1515
rect 56476 1535 56503 1545
rect 56476 1515 56480 1535
rect 56500 1515 56503 1535
rect 56476 1505 56503 1515
rect 56525 1540 56565 1545
rect 56525 1510 56530 1540
rect 56560 1510 56565 1540
rect 56525 1505 56565 1510
rect 56586 1535 56613 1545
rect 56586 1515 56590 1535
rect 56610 1515 56613 1535
rect 56586 1505 56613 1515
rect 56825 1535 56855 1545
rect 56825 1515 56830 1535
rect 56850 1515 56855 1535
rect 56825 1505 56855 1515
rect 56875 1535 56905 1545
rect 56875 1515 56880 1535
rect 56900 1515 56905 1535
rect 56875 1505 56905 1515
rect 56922 1540 56954 1545
rect 56922 1510 56925 1540
rect 56951 1510 56954 1540
rect 56922 1505 56954 1510
rect 57146 1540 57178 1545
rect 57146 1510 57149 1540
rect 57175 1510 57178 1540
rect 57146 1505 57178 1510
rect 57195 1535 57221 1545
rect 57195 1515 57198 1535
rect 57218 1515 57221 1535
rect 57195 1505 57221 1515
rect 57296 1535 57323 1545
rect 57296 1515 57300 1535
rect 57320 1515 57323 1535
rect 57296 1505 57323 1515
rect 57345 1540 57385 1545
rect 57345 1510 57350 1540
rect 57380 1510 57385 1540
rect 57345 1505 57385 1510
rect 57406 1535 57433 1545
rect 57406 1515 57410 1535
rect 57430 1515 57433 1535
rect 57406 1505 57433 1515
rect 57516 1535 57543 1545
rect 57516 1515 57520 1535
rect 57540 1515 57543 1535
rect 57516 1505 57543 1515
rect 57565 1540 57605 1545
rect 57565 1510 57570 1540
rect 57600 1510 57605 1540
rect 57565 1505 57605 1510
rect 57626 1535 57653 1545
rect 57626 1515 57630 1535
rect 57650 1515 57653 1535
rect 57626 1505 57653 1515
rect 55875 1485 55915 1490
rect 56155 1485 56175 1505
rect 56260 1485 56280 1505
rect 56370 1485 56390 1505
rect 56480 1485 56500 1505
rect 56590 1485 56610 1505
rect 55875 1455 55880 1485
rect 55910 1455 55915 1485
rect 55875 1450 55915 1455
rect 56145 1480 56185 1485
rect 56145 1450 56150 1480
rect 56180 1450 56185 1480
rect 56145 1445 56185 1450
rect 56250 1480 56290 1485
rect 56250 1450 56255 1480
rect 56285 1450 56290 1480
rect 56250 1445 56290 1450
rect 56360 1480 56400 1485
rect 56360 1450 56365 1480
rect 56395 1450 56400 1480
rect 56360 1445 56400 1450
rect 56470 1480 56510 1485
rect 56470 1450 56475 1480
rect 56505 1450 56510 1480
rect 56470 1445 56510 1450
rect 56580 1480 56620 1485
rect 56580 1450 56585 1480
rect 56615 1450 56620 1480
rect 56580 1445 56620 1450
rect 55955 1390 55995 1395
rect 55955 1360 55960 1390
rect 55990 1360 55995 1390
rect 55955 1355 55995 1360
rect 56770 1390 56810 1395
rect 56770 1360 56775 1390
rect 56805 1360 56810 1390
rect 56770 1355 56810 1360
rect 55965 835 55985 1355
rect 56330 1345 56370 1350
rect 56330 1315 56335 1345
rect 56365 1315 56370 1345
rect 56330 1310 56370 1315
rect 56340 1260 56360 1310
rect 56780 1260 56800 1355
rect 56835 1260 56855 1505
rect 56880 1350 56900 1505
rect 57195 1485 57215 1505
rect 57300 1485 57320 1505
rect 57410 1485 57430 1505
rect 57520 1485 57540 1505
rect 57630 1485 57650 1505
rect 57880 1495 57900 2610
rect 57915 2510 57955 2515
rect 57915 2480 57920 2510
rect 57950 2480 57955 2510
rect 57915 2475 57955 2480
rect 57870 1490 57910 1495
rect 57185 1480 57225 1485
rect 57185 1450 57190 1480
rect 57220 1450 57225 1480
rect 57185 1445 57225 1450
rect 57290 1480 57330 1485
rect 57290 1450 57295 1480
rect 57325 1450 57330 1480
rect 57290 1445 57330 1450
rect 57400 1480 57440 1485
rect 57400 1450 57405 1480
rect 57435 1450 57440 1480
rect 57400 1445 57440 1450
rect 57510 1480 57550 1485
rect 57510 1450 57515 1480
rect 57545 1450 57550 1480
rect 57510 1445 57550 1450
rect 57620 1480 57660 1485
rect 57620 1450 57625 1480
rect 57655 1450 57660 1480
rect 57870 1460 57875 1490
rect 57905 1460 57910 1490
rect 57870 1455 57910 1460
rect 57620 1445 57660 1450
rect 56870 1345 56910 1350
rect 56870 1315 56875 1345
rect 56905 1315 56910 1345
rect 56870 1310 56910 1315
rect 57200 1260 57220 1445
rect 57925 1370 57945 2475
rect 57985 1595 58005 3345
rect 59165 3325 59185 3365
rect 59105 3320 59246 3325
rect 59105 3290 59111 3320
rect 59141 3290 59160 3320
rect 59190 3290 59210 3320
rect 59240 3290 59246 3320
rect 59105 3285 59246 3290
rect 59105 2715 59246 2720
rect 58200 2710 58240 2715
rect 58200 2680 58205 2710
rect 58235 2680 58240 2710
rect 58200 2675 58240 2680
rect 58310 2710 58350 2715
rect 58310 2680 58315 2710
rect 58345 2680 58350 2710
rect 58310 2675 58350 2680
rect 58420 2710 58460 2715
rect 58420 2680 58425 2710
rect 58455 2680 58460 2710
rect 58420 2675 58460 2680
rect 58530 2710 58570 2715
rect 58530 2680 58535 2710
rect 58565 2680 58570 2710
rect 58530 2675 58570 2680
rect 58588 2705 58622 2715
rect 58588 2685 58596 2705
rect 58614 2685 58622 2705
rect 58588 2675 58622 2685
rect 58640 2710 58680 2715
rect 58640 2680 58645 2710
rect 58675 2680 58680 2710
rect 58640 2675 58680 2680
rect 58750 2710 58790 2715
rect 58750 2680 58755 2710
rect 58785 2680 58790 2710
rect 59105 2685 59111 2715
rect 59141 2685 59160 2715
rect 59190 2685 59210 2715
rect 59240 2685 59246 2715
rect 59105 2680 59246 2685
rect 58750 2675 58790 2680
rect 58040 2590 58080 2595
rect 58040 2560 58045 2590
rect 58075 2560 58080 2590
rect 58040 2555 58080 2560
rect 58050 2050 58070 2555
rect 58320 2550 58340 2675
rect 58475 2645 58515 2655
rect 58475 2625 58485 2645
rect 58505 2625 58515 2645
rect 58475 2615 58515 2625
rect 58310 2545 58350 2550
rect 58310 2515 58315 2545
rect 58345 2515 58350 2545
rect 58310 2510 58350 2515
rect 58485 2485 58505 2615
rect 58595 2595 58615 2675
rect 59165 2595 59185 2680
rect 59235 2650 59275 2660
rect 59235 2630 59245 2650
rect 59265 2630 59275 2650
rect 59235 2620 59275 2630
rect 58585 2590 58625 2595
rect 58585 2560 58590 2590
rect 58620 2560 58625 2590
rect 58585 2555 58625 2560
rect 59155 2590 59195 2595
rect 59155 2560 59160 2590
rect 59190 2560 59195 2590
rect 59155 2555 59195 2560
rect 58475 2475 58515 2485
rect 58475 2455 58485 2475
rect 58505 2455 58515 2475
rect 58475 2445 58515 2455
rect 58200 2420 58240 2425
rect 58200 2390 58205 2420
rect 58235 2390 58240 2420
rect 58200 2385 58240 2390
rect 58310 2420 58350 2425
rect 58310 2390 58315 2420
rect 58345 2390 58350 2420
rect 58310 2385 58350 2390
rect 58420 2420 58460 2425
rect 58420 2390 58425 2420
rect 58455 2390 58460 2420
rect 58420 2385 58460 2390
rect 58530 2420 58570 2425
rect 58530 2390 58535 2420
rect 58565 2390 58570 2420
rect 58530 2385 58570 2390
rect 58640 2420 58680 2425
rect 58640 2390 58645 2420
rect 58675 2390 58680 2420
rect 58640 2385 58680 2390
rect 58750 2420 58790 2425
rect 58750 2390 58755 2420
rect 58785 2390 58790 2420
rect 58750 2385 58790 2390
rect 59245 2320 59265 2620
rect 59445 2545 59485 2550
rect 59445 2515 59450 2545
rect 59480 2515 59485 2545
rect 59445 2510 59485 2515
rect 59235 2310 59275 2320
rect 59235 2290 59245 2310
rect 59265 2290 59275 2310
rect 59235 2280 59275 2290
rect 58255 2150 58295 2155
rect 58255 2120 58260 2150
rect 58290 2120 58295 2150
rect 58255 2115 58295 2120
rect 58313 2145 58347 2155
rect 58313 2125 58321 2145
rect 58339 2125 58347 2145
rect 58313 2115 58347 2125
rect 58365 2150 58405 2155
rect 58365 2120 58370 2150
rect 58400 2120 58405 2150
rect 58365 2115 58405 2120
rect 58475 2150 58515 2155
rect 58475 2120 58480 2150
rect 58510 2120 58515 2150
rect 58475 2115 58515 2120
rect 58585 2150 58625 2155
rect 58585 2120 58590 2150
rect 58620 2120 58625 2150
rect 58585 2115 58625 2120
rect 58695 2150 58735 2155
rect 58695 2120 58700 2150
rect 58730 2120 58735 2150
rect 58695 2115 58735 2120
rect 58975 2150 59015 2155
rect 58975 2120 58980 2150
rect 59010 2120 59015 2150
rect 58975 2115 59015 2120
rect 58320 2050 58340 2115
rect 58040 2045 58080 2050
rect 58040 2015 58045 2045
rect 58075 2015 58080 2045
rect 58040 2010 58080 2015
rect 58310 2045 58350 2050
rect 58310 2015 58315 2045
rect 58345 2015 58350 2045
rect 58310 2010 58350 2015
rect 58320 1965 58340 2010
rect 58255 1960 58295 1965
rect 58255 1930 58260 1960
rect 58290 1930 58295 1960
rect 58255 1925 58295 1930
rect 58313 1955 58347 1965
rect 58313 1935 58321 1955
rect 58339 1935 58347 1955
rect 58313 1925 58347 1935
rect 58365 1960 58405 1965
rect 58365 1930 58370 1960
rect 58400 1930 58405 1960
rect 58365 1925 58405 1930
rect 58475 1960 58515 1965
rect 58475 1930 58480 1960
rect 58510 1930 58515 1960
rect 58475 1925 58515 1930
rect 58585 1960 58625 1965
rect 58585 1930 58590 1960
rect 58620 1930 58625 1960
rect 58585 1925 58625 1930
rect 58695 1960 58735 1965
rect 58695 1930 58700 1960
rect 58730 1930 58735 1960
rect 58695 1925 58735 1930
rect 58930 1960 58970 1965
rect 58930 1930 58935 1960
rect 58965 1930 58970 1960
rect 58930 1925 58970 1930
rect 58875 1775 58915 1780
rect 58875 1745 58880 1775
rect 58910 1745 58915 1775
rect 58875 1740 58915 1745
rect 58085 1650 58125 1655
rect 58085 1620 58090 1650
rect 58120 1620 58125 1650
rect 58085 1615 58125 1620
rect 58940 1595 58960 1925
rect 57975 1590 58015 1595
rect 57975 1560 57980 1590
rect 58010 1560 58015 1590
rect 57975 1555 58015 1560
rect 58200 1590 58240 1595
rect 58200 1560 58205 1590
rect 58235 1560 58240 1590
rect 58200 1555 58240 1560
rect 58310 1590 58350 1595
rect 58310 1560 58315 1590
rect 58345 1560 58350 1590
rect 58310 1555 58350 1560
rect 58420 1590 58460 1595
rect 58420 1560 58425 1590
rect 58455 1560 58460 1590
rect 58420 1555 58460 1560
rect 58530 1590 58570 1595
rect 58530 1560 58535 1590
rect 58565 1560 58570 1590
rect 58530 1555 58570 1560
rect 58640 1590 58680 1595
rect 58640 1560 58645 1590
rect 58675 1560 58680 1590
rect 58640 1555 58680 1560
rect 58750 1590 58790 1595
rect 58750 1560 58755 1590
rect 58785 1560 58790 1590
rect 58750 1555 58790 1560
rect 58930 1590 58970 1595
rect 58930 1560 58935 1590
rect 58965 1560 58970 1590
rect 58930 1555 58970 1560
rect 58985 1540 59005 2115
rect 59455 1920 59475 2510
rect 59495 2420 59535 2425
rect 59495 2390 59500 2420
rect 59530 2390 59535 2420
rect 59495 2385 59535 2390
rect 59440 1910 59490 1920
rect 59440 1880 59450 1910
rect 59480 1880 59490 1910
rect 59440 1870 59490 1880
rect 59025 1775 59065 1780
rect 59025 1745 59030 1775
rect 59060 1745 59065 1775
rect 59025 1740 59065 1745
rect 59115 1595 59150 1600
rect 59115 1555 59150 1560
rect 59175 1595 59210 1601
rect 59175 1555 59210 1560
rect 59235 1595 59270 1600
rect 59235 1555 59270 1560
rect 59295 1595 59330 1601
rect 59295 1555 59330 1560
rect 59180 1540 59200 1555
rect 58975 1535 59015 1540
rect 58475 1525 58515 1535
rect 58475 1505 58485 1525
rect 58505 1505 58515 1525
rect 58475 1495 58515 1505
rect 58975 1505 58980 1535
rect 59010 1505 59015 1535
rect 58975 1500 59015 1505
rect 59170 1535 59210 1540
rect 59170 1505 59175 1535
rect 59205 1505 59210 1535
rect 59170 1500 59210 1505
rect 59300 1495 59320 1555
rect 58485 1435 58505 1495
rect 59290 1490 59330 1495
rect 59290 1460 59295 1490
rect 59325 1460 59330 1490
rect 59290 1455 59330 1460
rect 58015 1425 58055 1430
rect 58015 1395 58020 1425
rect 58050 1395 58055 1425
rect 58015 1390 58055 1395
rect 58325 1425 58365 1430
rect 58325 1395 58330 1425
rect 58360 1395 58365 1425
rect 58475 1425 58515 1435
rect 58475 1405 58485 1425
rect 58505 1405 58515 1425
rect 58475 1395 58515 1405
rect 59035 1425 59075 1430
rect 59035 1395 59040 1425
rect 59070 1395 59075 1425
rect 58325 1390 58365 1395
rect 59035 1390 59075 1395
rect 58335 1375 58355 1390
rect 58225 1370 58265 1375
rect 57470 1365 57510 1370
rect 57470 1335 57475 1365
rect 57505 1335 57510 1365
rect 57470 1330 57510 1335
rect 57915 1365 57955 1370
rect 57915 1335 57920 1365
rect 57950 1335 57955 1365
rect 58225 1340 58230 1370
rect 58260 1340 58265 1370
rect 58225 1335 58265 1340
rect 58328 1365 58362 1375
rect 58328 1345 58336 1365
rect 58354 1345 58362 1365
rect 58328 1335 58362 1345
rect 58425 1370 58465 1375
rect 58425 1340 58430 1370
rect 58460 1340 58465 1370
rect 58425 1335 58465 1340
rect 58625 1370 58665 1375
rect 58625 1340 58630 1370
rect 58660 1340 58665 1370
rect 58625 1335 58665 1340
rect 58970 1370 59010 1375
rect 58970 1340 58975 1370
rect 59005 1340 59010 1370
rect 58970 1335 59010 1340
rect 57915 1330 57955 1335
rect 57480 1260 57500 1330
rect 58980 1315 59000 1335
rect 59045 1315 59065 1390
rect 59455 1375 59475 1870
rect 59445 1370 59485 1375
rect 59445 1340 59450 1370
rect 59480 1340 59485 1370
rect 59445 1335 59485 1340
rect 58975 1310 59010 1315
rect 58975 1270 59010 1275
rect 59035 1310 59070 1315
rect 59035 1270 59070 1275
rect 56330 1250 56370 1260
rect 56330 1230 56340 1250
rect 56360 1230 56370 1250
rect 56330 1220 56370 1230
rect 56440 1255 56480 1260
rect 56440 1225 56445 1255
rect 56475 1225 56480 1255
rect 56440 1220 56480 1225
rect 56550 1255 56590 1260
rect 56550 1225 56555 1255
rect 56585 1225 56590 1255
rect 56550 1220 56590 1225
rect 56660 1255 56700 1260
rect 56660 1225 56665 1255
rect 56695 1225 56700 1255
rect 56660 1220 56700 1225
rect 56770 1255 56810 1260
rect 56770 1225 56775 1255
rect 56805 1225 56810 1255
rect 56770 1220 56810 1225
rect 56830 1250 56860 1260
rect 56830 1230 56835 1250
rect 56855 1230 56860 1250
rect 56830 1220 56860 1230
rect 56880 1255 56920 1260
rect 56880 1225 56885 1255
rect 56915 1225 56920 1255
rect 56880 1220 56920 1225
rect 56990 1255 57030 1260
rect 56990 1225 56995 1255
rect 57025 1225 57030 1255
rect 56990 1220 57030 1225
rect 57100 1255 57140 1260
rect 57100 1225 57105 1255
rect 57135 1225 57140 1255
rect 57100 1220 57140 1225
rect 57200 1255 57250 1260
rect 57200 1225 57215 1255
rect 57245 1225 57250 1255
rect 57200 1220 57250 1225
rect 57320 1255 57360 1260
rect 57320 1225 57325 1255
rect 57355 1225 57360 1255
rect 57320 1220 57360 1225
rect 57415 1255 57455 1260
rect 57415 1225 57420 1255
rect 57450 1225 57455 1255
rect 57415 1220 57455 1225
rect 57474 1250 57504 1260
rect 57474 1230 57479 1250
rect 57499 1230 57504 1250
rect 57474 1220 57504 1230
rect 58795 985 58835 990
rect 58795 955 58800 985
rect 58830 955 58835 985
rect 58795 950 58835 955
rect 58885 985 58925 990
rect 58885 955 58890 985
rect 58920 955 58925 985
rect 58885 950 58925 955
rect 56210 935 56250 940
rect 56210 905 56215 935
rect 56245 905 56250 935
rect 56210 900 56250 905
rect 56275 935 56315 940
rect 56275 905 56280 935
rect 56310 905 56315 935
rect 56275 900 56315 905
rect 56385 935 56425 940
rect 56385 905 56390 935
rect 56420 905 56425 935
rect 56385 900 56425 905
rect 56495 935 56535 940
rect 56495 905 56500 935
rect 56530 905 56535 935
rect 56495 900 56535 905
rect 56605 935 56645 940
rect 56605 905 56610 935
rect 56640 905 56645 935
rect 56605 900 56645 905
rect 56715 935 56755 940
rect 56715 905 56720 935
rect 56750 905 56755 935
rect 56715 900 56755 905
rect 56825 935 56865 940
rect 56825 905 56830 935
rect 56860 905 56865 935
rect 56825 900 56865 905
rect 56935 935 56975 940
rect 56935 905 56940 935
rect 56970 905 56975 935
rect 56935 900 56975 905
rect 57045 935 57085 940
rect 57045 905 57050 935
rect 57080 905 57085 935
rect 57045 900 57085 905
rect 57155 935 57195 940
rect 57155 905 57160 935
rect 57190 905 57195 935
rect 57155 900 57195 905
rect 57265 935 57305 940
rect 57265 905 57270 935
rect 57300 905 57305 935
rect 57265 900 57305 905
rect 57375 935 57415 940
rect 57375 905 57380 935
rect 57410 905 57415 935
rect 57375 900 57415 905
rect 57485 935 57525 940
rect 57485 905 57490 935
rect 57520 905 57525 935
rect 57485 900 57525 905
rect 57545 935 57585 940
rect 57545 905 57550 935
rect 57580 905 57585 935
rect 57545 900 57585 905
rect 57975 925 58015 930
rect 57975 895 57980 925
rect 58010 895 58015 925
rect 57975 890 58015 895
rect 55955 830 55995 835
rect 55955 800 55960 830
rect 55990 800 55995 830
rect 55955 795 55995 800
rect 57055 830 57095 835
rect 57055 800 57060 830
rect 57090 800 57095 830
rect 57055 795 57095 800
rect 57065 745 57085 795
rect 55830 740 55870 745
rect 55830 710 55835 740
rect 55865 710 55870 740
rect 55830 705 55870 710
rect 56755 740 56795 745
rect 56755 710 56760 740
rect 56790 710 56795 740
rect 56755 705 56795 710
rect 56875 740 56915 745
rect 56875 710 56880 740
rect 56910 710 56915 740
rect 56875 705 56915 710
rect 56995 740 57035 745
rect 56995 710 57000 740
rect 57030 710 57035 740
rect 56995 705 57035 710
rect 57055 735 57095 745
rect 57055 715 57065 735
rect 57085 715 57095 735
rect 57055 705 57095 715
rect 57985 605 58005 890
rect 55235 600 55275 605
rect 55235 570 55240 600
rect 55270 570 55275 600
rect 55235 565 55275 570
rect 55335 600 55375 605
rect 55335 570 55340 600
rect 55370 570 55375 600
rect 55335 565 55375 570
rect 55435 600 55475 605
rect 55435 570 55440 600
rect 55470 570 55475 600
rect 55435 565 55475 570
rect 55785 600 55825 605
rect 55785 570 55790 600
rect 55820 570 55825 600
rect 55785 565 55825 570
rect 57975 600 58015 605
rect 57975 570 57980 600
rect 58010 570 58015 600
rect 57975 565 58015 570
rect 58325 600 58365 605
rect 58325 570 58330 600
rect 58360 570 58365 600
rect 58325 565 58365 570
rect 58425 600 58465 605
rect 58425 570 58430 600
rect 58460 570 58465 600
rect 58425 565 58465 570
rect 58525 600 58565 605
rect 58525 570 58530 600
rect 58560 570 58565 600
rect 58525 565 58565 570
rect 55345 545 55365 565
rect 55335 540 55375 545
rect 55335 510 55340 540
rect 55370 510 55375 540
rect 55335 505 55375 510
rect 55795 500 55815 565
rect 56875 545 56915 555
rect 56875 525 56885 545
rect 56905 525 56915 545
rect 56875 515 56915 525
rect 56885 500 56905 515
rect 57985 500 58005 565
rect 58435 545 58455 565
rect 58425 540 58465 545
rect 58425 510 58430 540
rect 58460 510 58465 540
rect 58425 505 58465 510
rect 59505 500 59525 2385
rect 54265 495 54305 500
rect 54265 465 54270 495
rect 54300 465 54305 495
rect 54265 460 54305 465
rect 55785 495 55825 500
rect 55785 465 55790 495
rect 55820 465 55825 495
rect 55785 460 55825 465
rect 56875 495 56915 500
rect 56875 465 56880 495
rect 56910 465 56915 495
rect 56875 460 56915 465
rect 57975 495 58015 500
rect 57975 465 57980 495
rect 58010 465 58015 495
rect 57975 460 58015 465
rect 59495 495 59535 500
rect 59495 465 59500 495
rect 59530 465 59535 495
rect 59495 460 59535 465
rect 57985 -510 58005 460
rect 57975 -515 58015 -510
rect 57975 -545 57980 -515
rect 58010 -545 58015 -515
rect 57975 -550 58015 -545
<< via1 >>
rect 55790 6155 55820 6185
rect 56885 4850 56915 4880
rect 57555 4850 57585 4880
rect 57495 4820 57525 4825
rect 57495 4800 57500 4820
rect 57500 4800 57520 4820
rect 57520 4800 57525 4820
rect 57495 4795 57525 4800
rect 57555 4820 57585 4825
rect 57555 4800 57560 4820
rect 57560 4800 57580 4820
rect 57580 4800 57585 4820
rect 57555 4795 57585 4800
rect 57675 4820 57705 4825
rect 57675 4800 57680 4820
rect 57680 4800 57700 4820
rect 57700 4800 57705 4820
rect 57675 4795 57705 4800
rect 56330 4755 56360 4785
rect 56825 4780 56855 4785
rect 56825 4760 56830 4780
rect 56830 4760 56850 4780
rect 56850 4760 56855 4780
rect 56825 4755 56855 4760
rect 56945 4780 56975 4785
rect 56945 4760 56950 4780
rect 56950 4760 56970 4780
rect 56970 4760 56975 4780
rect 56945 4755 56975 4760
rect 57005 4780 57035 4785
rect 57005 4760 57010 4780
rect 57010 4760 57030 4780
rect 57030 4760 57035 4780
rect 57005 4755 57035 4760
rect 55790 4500 55820 4530
rect 56150 4525 56180 4530
rect 56150 4505 56155 4525
rect 56155 4505 56175 4525
rect 56175 4505 56180 4525
rect 56150 4500 56180 4505
rect 56210 4525 56240 4530
rect 56210 4505 56215 4525
rect 56215 4505 56235 4525
rect 56235 4505 56240 4525
rect 56210 4500 56240 4505
rect 56330 4525 56360 4530
rect 56330 4505 56335 4525
rect 56335 4505 56355 4525
rect 56355 4505 56360 4525
rect 56330 4500 56360 4505
rect 56915 4385 56945 4390
rect 56915 4365 56920 4385
rect 56920 4365 56940 4385
rect 56940 4365 56945 4385
rect 56915 4360 56945 4365
rect 57620 4390 57650 4395
rect 57620 4370 57625 4390
rect 57625 4370 57645 4390
rect 57645 4370 57650 4390
rect 57620 4365 57650 4370
rect 56240 4260 56270 4290
rect 56855 4260 56885 4290
rect 55320 4170 55350 4200
rect 55790 4170 55820 4200
rect 55080 4085 55110 4090
rect 55080 4065 55085 4085
rect 55085 4065 55105 4085
rect 55105 4065 55110 4085
rect 55080 4060 55110 4065
rect 55200 4085 55230 4090
rect 55200 4065 55205 4085
rect 55205 4065 55225 4085
rect 55225 4065 55230 4085
rect 55200 4060 55230 4065
rect 55320 4085 55350 4090
rect 55320 4065 55325 4085
rect 55325 4065 55345 4085
rect 55345 4065 55350 4085
rect 55320 4060 55350 4065
rect 55440 4085 55470 4090
rect 55440 4065 55445 4085
rect 55445 4065 55465 4085
rect 55465 4065 55470 4085
rect 55440 4060 55470 4065
rect 55560 4085 55590 4090
rect 55560 4065 55565 4085
rect 55565 4065 55585 4085
rect 55585 4065 55590 4085
rect 55560 4060 55590 4065
rect 55020 3665 55050 3670
rect 55020 3645 55025 3665
rect 55025 3645 55045 3665
rect 55045 3645 55050 3665
rect 55020 3640 55050 3645
rect 55140 3665 55170 3670
rect 55140 3645 55145 3665
rect 55145 3645 55165 3665
rect 55165 3645 55170 3665
rect 55140 3640 55170 3645
rect 55260 3665 55290 3670
rect 55260 3645 55265 3665
rect 55265 3645 55285 3665
rect 55285 3645 55290 3665
rect 55260 3640 55290 3645
rect 55380 3665 55410 3670
rect 55380 3645 55385 3665
rect 55385 3645 55405 3665
rect 55405 3645 55410 3665
rect 55380 3640 55410 3645
rect 55500 3665 55530 3670
rect 55500 3645 55505 3665
rect 55505 3645 55525 3665
rect 55525 3645 55530 3665
rect 55500 3640 55530 3645
rect 55620 3665 55650 3670
rect 55620 3645 55625 3665
rect 55625 3645 55645 3665
rect 55645 3645 55650 3665
rect 55620 3640 55650 3645
rect 55320 3540 55350 3570
rect 54610 3370 54640 3400
rect 55895 4060 55925 4090
rect 56130 4085 56160 4090
rect 56130 4065 56135 4085
rect 56135 4065 56155 4085
rect 56155 4065 56160 4085
rect 56130 4060 56160 4065
rect 56190 4060 56220 4090
rect 56250 4085 56280 4090
rect 56250 4065 56255 4085
rect 56255 4065 56275 4085
rect 56275 4065 56280 4085
rect 56250 4060 56280 4065
rect 56370 4085 56400 4090
rect 56370 4065 56375 4085
rect 56375 4065 56395 4085
rect 56395 4065 56400 4085
rect 56370 4060 56400 4065
rect 56490 4085 56520 4090
rect 56490 4065 56495 4085
rect 56495 4065 56515 4085
rect 56515 4065 56520 4085
rect 56490 4060 56520 4065
rect 56610 4085 56640 4090
rect 56610 4065 56615 4085
rect 56615 4065 56635 4085
rect 56635 4065 56640 4085
rect 56610 4060 56640 4065
rect 55895 3640 55925 3670
rect 56070 3665 56100 3670
rect 56070 3645 56075 3665
rect 56075 3645 56095 3665
rect 56095 3645 56100 3665
rect 56070 3640 56100 3645
rect 56190 3665 56220 3670
rect 56190 3645 56195 3665
rect 56195 3645 56215 3665
rect 56215 3645 56220 3665
rect 56190 3640 56220 3645
rect 56310 3665 56340 3670
rect 56310 3645 56315 3665
rect 56315 3645 56335 3665
rect 56335 3645 56340 3665
rect 56310 3640 56340 3645
rect 56430 3665 56460 3670
rect 56430 3645 56435 3665
rect 56435 3645 56455 3665
rect 56455 3645 56460 3665
rect 56430 3640 56460 3645
rect 56550 3665 56580 3670
rect 56550 3645 56555 3665
rect 56555 3645 56575 3665
rect 56575 3645 56580 3665
rect 56550 3640 56580 3645
rect 56670 3665 56700 3670
rect 56670 3645 56675 3665
rect 56675 3645 56695 3665
rect 56695 3645 56700 3665
rect 56670 3640 56700 3645
rect 54960 3375 54990 3380
rect 54960 3355 54965 3375
rect 54965 3355 54985 3375
rect 54985 3355 54990 3375
rect 54960 3350 54990 3355
rect 55070 3375 55100 3380
rect 55070 3355 55075 3375
rect 55075 3355 55095 3375
rect 55095 3355 55100 3375
rect 55070 3350 55100 3355
rect 55180 3375 55210 3380
rect 55180 3355 55185 3375
rect 55185 3355 55205 3375
rect 55205 3355 55210 3375
rect 55180 3350 55210 3355
rect 55290 3375 55320 3380
rect 55290 3355 55295 3375
rect 55295 3355 55315 3375
rect 55315 3355 55320 3375
rect 55290 3350 55320 3355
rect 55400 3375 55430 3380
rect 55400 3355 55405 3375
rect 55405 3355 55425 3375
rect 55425 3355 55430 3375
rect 55400 3350 55430 3355
rect 55510 3375 55540 3380
rect 55510 3355 55515 3375
rect 55515 3355 55535 3375
rect 55535 3355 55540 3375
rect 55510 3350 55540 3355
rect 55620 3375 55650 3380
rect 55620 3355 55625 3375
rect 55625 3355 55645 3375
rect 55645 3355 55650 3375
rect 55620 3350 55650 3355
rect 55790 3350 55820 3380
rect 54560 3290 54590 3320
rect 54610 3290 54640 3320
rect 54659 3290 54689 3320
rect 55745 3295 55775 3325
rect 54560 2685 54590 2715
rect 54610 2685 54640 2715
rect 54659 2685 54689 2715
rect 55015 2705 55045 2710
rect 55015 2685 55020 2705
rect 55020 2685 55040 2705
rect 55040 2685 55045 2705
rect 55015 2680 55045 2685
rect 54320 2515 54350 2545
rect 54270 2390 54300 2420
rect 55125 2705 55155 2710
rect 55125 2685 55130 2705
rect 55130 2685 55150 2705
rect 55150 2685 55155 2705
rect 55125 2680 55155 2685
rect 55235 2705 55265 2710
rect 55235 2685 55240 2705
rect 55240 2685 55260 2705
rect 55260 2685 55265 2705
rect 55235 2680 55265 2685
rect 55345 2705 55375 2710
rect 55345 2685 55350 2705
rect 55350 2685 55370 2705
rect 55370 2685 55375 2705
rect 55345 2680 55375 2685
rect 55455 2705 55485 2710
rect 55455 2685 55460 2705
rect 55460 2685 55480 2705
rect 55480 2685 55485 2705
rect 55455 2680 55485 2685
rect 55565 2705 55595 2710
rect 55565 2685 55570 2705
rect 55570 2685 55590 2705
rect 55590 2685 55595 2705
rect 55565 2680 55595 2685
rect 54610 2560 54640 2590
rect 55180 2560 55210 2590
rect 56370 3585 56400 3615
rect 56855 3585 56885 3615
rect 57570 4260 57600 4290
rect 57980 4170 58010 4200
rect 58450 4170 58480 4200
rect 57160 4085 57190 4090
rect 57160 4065 57165 4085
rect 57165 4065 57185 4085
rect 57185 4065 57190 4085
rect 57160 4060 57190 4065
rect 57280 4085 57310 4090
rect 57280 4065 57285 4085
rect 57285 4065 57305 4085
rect 57305 4065 57310 4085
rect 57280 4060 57310 4065
rect 57400 4085 57430 4090
rect 57400 4065 57405 4085
rect 57405 4065 57425 4085
rect 57425 4065 57430 4085
rect 57400 4060 57430 4065
rect 57520 4085 57550 4090
rect 57520 4065 57525 4085
rect 57525 4065 57545 4085
rect 57545 4065 57550 4085
rect 57520 4060 57550 4065
rect 57580 4060 57610 4090
rect 57640 4085 57670 4090
rect 57640 4065 57645 4085
rect 57645 4065 57665 4085
rect 57665 4065 57670 4085
rect 57640 4060 57670 4065
rect 57875 4060 57905 4090
rect 57100 3665 57130 3670
rect 57100 3645 57105 3665
rect 57105 3645 57125 3665
rect 57125 3645 57130 3665
rect 57100 3640 57130 3645
rect 57220 3665 57250 3670
rect 57220 3645 57225 3665
rect 57225 3645 57245 3665
rect 57245 3645 57250 3665
rect 57220 3640 57250 3645
rect 57340 3665 57370 3670
rect 57340 3645 57345 3665
rect 57345 3645 57365 3665
rect 57365 3645 57370 3665
rect 57340 3640 57370 3645
rect 57460 3665 57490 3670
rect 57460 3645 57465 3665
rect 57465 3645 57485 3665
rect 57485 3645 57490 3665
rect 57460 3640 57490 3645
rect 57580 3665 57610 3670
rect 57580 3645 57585 3665
rect 57585 3645 57605 3665
rect 57605 3645 57610 3665
rect 57580 3640 57610 3645
rect 57700 3665 57730 3670
rect 57700 3645 57705 3665
rect 57705 3645 57725 3665
rect 57725 3645 57730 3665
rect 57700 3640 57730 3645
rect 57875 3640 57905 3670
rect 57400 3585 57430 3615
rect 56915 3540 56945 3570
rect 58210 4085 58240 4090
rect 58210 4065 58215 4085
rect 58215 4065 58235 4085
rect 58235 4065 58240 4085
rect 58210 4060 58240 4065
rect 58330 4085 58360 4090
rect 58330 4065 58335 4085
rect 58335 4065 58355 4085
rect 58355 4065 58360 4085
rect 58330 4060 58360 4065
rect 58450 4085 58480 4090
rect 58450 4065 58455 4085
rect 58455 4065 58475 4085
rect 58475 4065 58480 4085
rect 58450 4060 58480 4065
rect 58570 4085 58600 4090
rect 58570 4065 58575 4085
rect 58575 4065 58595 4085
rect 58595 4065 58600 4085
rect 58570 4060 58600 4065
rect 58690 4085 58720 4090
rect 58690 4065 58695 4085
rect 58695 4065 58715 4085
rect 58715 4065 58720 4085
rect 58690 4060 58720 4065
rect 58150 3665 58180 3670
rect 58150 3645 58155 3665
rect 58155 3645 58175 3665
rect 58175 3645 58180 3665
rect 58150 3640 58180 3645
rect 58270 3665 58300 3670
rect 58270 3645 58275 3665
rect 58275 3645 58295 3665
rect 58295 3645 58300 3665
rect 58270 3640 58300 3645
rect 58390 3665 58420 3670
rect 58390 3645 58395 3665
rect 58395 3645 58415 3665
rect 58415 3645 58420 3665
rect 58390 3640 58420 3645
rect 58510 3665 58540 3670
rect 58510 3645 58515 3665
rect 58515 3645 58535 3665
rect 58535 3645 58540 3665
rect 58510 3640 58540 3645
rect 58630 3665 58660 3670
rect 58630 3645 58635 3665
rect 58635 3645 58655 3665
rect 58655 3645 58660 3665
rect 58630 3640 58660 3645
rect 58750 3665 58780 3670
rect 58750 3645 58755 3665
rect 58755 3645 58775 3665
rect 58775 3645 58780 3665
rect 58750 3640 58780 3645
rect 58450 3540 58480 3570
rect 56280 3375 56310 3380
rect 56280 3355 56285 3375
rect 56285 3355 56305 3375
rect 56305 3355 56310 3375
rect 56280 3350 56310 3355
rect 56390 3375 56420 3380
rect 56390 3355 56395 3375
rect 56395 3355 56415 3375
rect 56415 3355 56420 3375
rect 56390 3350 56420 3355
rect 56500 3375 56530 3380
rect 56500 3355 56505 3375
rect 56505 3355 56525 3375
rect 56525 3355 56530 3375
rect 56500 3350 56530 3355
rect 56610 3375 56640 3380
rect 56610 3355 56615 3375
rect 56615 3355 56635 3375
rect 56635 3355 56640 3375
rect 56610 3350 56640 3355
rect 56720 3375 56750 3380
rect 56720 3355 56725 3375
rect 56725 3355 56745 3375
rect 56745 3355 56750 3375
rect 56720 3350 56750 3355
rect 56830 3375 56860 3380
rect 56830 3355 56835 3375
rect 56835 3355 56855 3375
rect 56855 3355 56860 3375
rect 56830 3350 56860 3355
rect 56940 3375 56970 3380
rect 56940 3355 56945 3375
rect 56945 3355 56965 3375
rect 56965 3355 56970 3375
rect 56940 3350 56970 3355
rect 57050 3375 57080 3380
rect 57050 3355 57055 3375
rect 57055 3355 57075 3375
rect 57075 3355 57080 3375
rect 57050 3350 57080 3355
rect 57160 3375 57190 3380
rect 57160 3355 57165 3375
rect 57165 3355 57185 3375
rect 57185 3355 57190 3375
rect 57160 3350 57190 3355
rect 57270 3375 57300 3380
rect 57270 3355 57275 3375
rect 57275 3355 57295 3375
rect 57295 3355 57300 3375
rect 57270 3350 57300 3355
rect 57380 3375 57410 3380
rect 57380 3355 57385 3375
rect 57385 3355 57405 3375
rect 57405 3355 57410 3375
rect 57380 3350 57410 3355
rect 57490 3375 57520 3380
rect 57490 3355 57495 3375
rect 57495 3355 57515 3375
rect 57515 3355 57520 3375
rect 57490 3350 57520 3355
rect 57980 3350 58010 3380
rect 58150 3375 58180 3380
rect 58150 3355 58155 3375
rect 58155 3355 58175 3375
rect 58175 3355 58180 3375
rect 58150 3350 58180 3355
rect 58260 3375 58290 3380
rect 58260 3355 58265 3375
rect 58265 3355 58285 3375
rect 58285 3355 58290 3375
rect 58260 3350 58290 3355
rect 58370 3375 58400 3380
rect 58370 3355 58375 3375
rect 58375 3355 58395 3375
rect 58395 3355 58400 3375
rect 58370 3350 58400 3355
rect 58480 3375 58510 3380
rect 58480 3355 58485 3375
rect 58485 3355 58505 3375
rect 58505 3355 58510 3375
rect 58480 3350 58510 3355
rect 58590 3375 58620 3380
rect 58590 3355 58595 3375
rect 58595 3355 58615 3375
rect 58615 3355 58620 3375
rect 58590 3350 58620 3355
rect 58700 3375 58730 3380
rect 58700 3355 58705 3375
rect 58705 3355 58725 3375
rect 58725 3355 58730 3375
rect 58700 3350 58730 3355
rect 58810 3375 58840 3380
rect 58810 3355 58815 3375
rect 58815 3355 58835 3375
rect 58835 3355 58840 3375
rect 58810 3350 58840 3355
rect 59160 3370 59190 3400
rect 56070 3295 56100 3325
rect 56335 3255 56365 3260
rect 56335 3235 56340 3255
rect 56340 3235 56360 3255
rect 56360 3235 56365 3255
rect 56335 3230 56365 3235
rect 56555 3255 56585 3260
rect 56555 3235 56560 3255
rect 56560 3235 56580 3255
rect 56580 3235 56585 3255
rect 56555 3230 56585 3235
rect 56775 3255 56805 3260
rect 56775 3235 56780 3255
rect 56780 3235 56800 3255
rect 56800 3235 56805 3255
rect 56775 3230 56805 3235
rect 56995 3255 57025 3260
rect 56995 3235 57000 3255
rect 57000 3235 57020 3255
rect 57020 3235 57025 3255
rect 56995 3230 57025 3235
rect 57215 3255 57245 3260
rect 57215 3235 57220 3255
rect 57220 3235 57240 3255
rect 57240 3235 57245 3255
rect 57215 3230 57245 3235
rect 57435 3255 57465 3260
rect 57435 3235 57440 3255
rect 57440 3235 57460 3255
rect 57460 3235 57465 3255
rect 57435 3230 57465 3235
rect 56445 3175 56475 3205
rect 56480 3015 56510 3045
rect 56665 3175 56695 3205
rect 56885 3175 56915 3205
rect 57105 3175 57135 3205
rect 56190 2955 56220 2985
rect 56290 2955 56320 2985
rect 56400 2955 56430 2985
rect 57325 3175 57355 3205
rect 56510 2955 56540 2985
rect 56620 2955 56650 2985
rect 57160 2955 57190 2985
rect 57260 2955 57290 2985
rect 57370 2955 57400 2985
rect 57480 2955 57510 2985
rect 57590 2955 57620 2985
rect 56147 2920 56173 2924
rect 56147 2900 56150 2920
rect 56150 2900 56170 2920
rect 56170 2900 56173 2920
rect 56147 2896 56173 2900
rect 56347 2920 56373 2924
rect 56347 2900 56350 2920
rect 56350 2900 56370 2920
rect 56370 2900 56373 2920
rect 56347 2896 56373 2900
rect 56565 2920 56595 2925
rect 56565 2900 56570 2920
rect 56570 2900 56590 2920
rect 56590 2900 56595 2920
rect 56565 2895 56595 2900
rect 56885 2895 56915 2925
rect 57115 2920 57141 2924
rect 57115 2900 57118 2920
rect 57118 2900 57138 2920
rect 57138 2900 57141 2920
rect 57115 2896 57141 2900
rect 57315 2920 57345 2925
rect 57315 2900 57320 2920
rect 57320 2900 57340 2920
rect 57340 2900 57345 2920
rect 57315 2895 57345 2900
rect 57535 2920 57565 2925
rect 57535 2900 57540 2920
rect 57540 2900 57560 2920
rect 57560 2900 57565 2920
rect 57535 2895 57565 2900
rect 55790 2835 55820 2865
rect 56010 2860 56040 2865
rect 56010 2840 56015 2860
rect 56015 2840 56035 2860
rect 56035 2840 56040 2860
rect 56010 2835 56040 2840
rect 56790 2860 56820 2865
rect 56790 2840 56795 2860
rect 56795 2840 56815 2860
rect 56815 2840 56820 2860
rect 56790 2835 56820 2840
rect 55745 2560 55775 2590
rect 55455 2515 55485 2545
rect 55015 2415 55045 2420
rect 55015 2395 55020 2415
rect 55020 2395 55040 2415
rect 55040 2395 55045 2415
rect 55015 2390 55045 2395
rect 55125 2415 55155 2420
rect 55125 2395 55130 2415
rect 55130 2395 55150 2415
rect 55150 2395 55155 2415
rect 55125 2390 55155 2395
rect 55235 2415 55265 2420
rect 55235 2395 55240 2415
rect 55240 2395 55260 2415
rect 55260 2395 55265 2415
rect 55235 2390 55265 2395
rect 55345 2415 55375 2420
rect 55345 2395 55350 2415
rect 55350 2395 55370 2415
rect 55370 2395 55375 2415
rect 55345 2390 55375 2395
rect 55455 2415 55485 2420
rect 55455 2395 55460 2415
rect 55460 2395 55480 2415
rect 55480 2395 55485 2415
rect 55455 2390 55485 2395
rect 55565 2415 55595 2420
rect 55565 2395 55570 2415
rect 55570 2395 55590 2415
rect 55590 2395 55595 2415
rect 55565 2390 55595 2395
rect 54795 2120 54825 2150
rect 55070 2145 55100 2150
rect 55070 2125 55075 2145
rect 55075 2125 55095 2145
rect 55095 2125 55100 2145
rect 55070 2120 55100 2125
rect 55180 2145 55210 2150
rect 55180 2125 55185 2145
rect 55185 2125 55205 2145
rect 55205 2125 55210 2145
rect 55180 2120 55210 2125
rect 55290 2145 55320 2150
rect 55290 2125 55295 2145
rect 55295 2125 55315 2145
rect 55315 2125 55320 2145
rect 55290 2120 55320 2125
rect 55400 2145 55430 2150
rect 55400 2125 55405 2145
rect 55405 2125 55425 2145
rect 55425 2125 55430 2145
rect 55400 2120 55430 2125
rect 55510 2145 55540 2150
rect 55510 2125 55515 2145
rect 55515 2125 55535 2145
rect 55535 2125 55540 2145
rect 55510 2120 55540 2125
rect 54320 1880 54350 1910
rect 54740 1770 54770 1775
rect 54740 1750 54745 1770
rect 54745 1750 54765 1770
rect 54765 1750 54770 1770
rect 54740 1745 54770 1750
rect 54470 1590 54505 1595
rect 54470 1565 54475 1590
rect 54475 1565 54500 1590
rect 54500 1565 54505 1590
rect 54470 1560 54505 1565
rect 54530 1590 54565 1595
rect 54530 1565 54535 1590
rect 54535 1565 54560 1590
rect 54560 1565 54565 1590
rect 54530 1560 54565 1565
rect 54590 1590 54625 1595
rect 54590 1565 54595 1590
rect 54595 1565 54620 1590
rect 54620 1565 54625 1590
rect 54590 1560 54625 1565
rect 54650 1590 54685 1595
rect 54650 1565 54655 1590
rect 54655 1565 54680 1590
rect 54680 1565 54685 1590
rect 54650 1560 54685 1565
rect 55455 2015 55485 2045
rect 55745 2015 55775 2045
rect 54840 1930 54870 1960
rect 55070 1955 55100 1960
rect 55070 1935 55075 1955
rect 55075 1935 55095 1955
rect 55095 1935 55100 1955
rect 55070 1930 55100 1935
rect 55180 1955 55210 1960
rect 55180 1935 55185 1955
rect 55185 1935 55205 1955
rect 55205 1935 55210 1955
rect 55180 1930 55210 1935
rect 55290 1955 55320 1960
rect 55290 1935 55295 1955
rect 55295 1935 55315 1955
rect 55315 1935 55320 1955
rect 55290 1930 55320 1935
rect 55400 1955 55430 1960
rect 55400 1935 55405 1955
rect 55405 1935 55425 1955
rect 55425 1935 55430 1955
rect 55400 1930 55430 1935
rect 55510 1955 55540 1960
rect 55510 1935 55515 1955
rect 55515 1935 55535 1955
rect 55535 1935 55540 1955
rect 55510 1930 55540 1935
rect 54890 1770 54920 1775
rect 54890 1750 54895 1770
rect 54895 1750 54915 1770
rect 54915 1750 54920 1770
rect 54890 1745 54920 1750
rect 56275 2800 56301 2805
rect 56275 2780 56278 2800
rect 56278 2780 56295 2800
rect 56295 2780 56301 2800
rect 56275 2775 56301 2780
rect 56495 2800 56521 2805
rect 56495 2780 56498 2800
rect 56498 2780 56515 2800
rect 56515 2780 56521 2800
rect 56495 2775 56521 2780
rect 56639 2800 56665 2805
rect 56639 2780 56645 2800
rect 56645 2780 56662 2800
rect 56662 2780 56665 2800
rect 56639 2775 56665 2780
rect 56125 2715 56155 2745
rect 56230 2715 56260 2745
rect 56345 2715 56375 2745
rect 56450 2715 56480 2745
rect 56565 2715 56595 2745
rect 56680 2715 56710 2745
rect 56610 2660 56640 2690
rect 55880 2615 55910 2645
rect 55835 2200 55865 2230
rect 54840 1560 54870 1590
rect 55015 1585 55045 1590
rect 55015 1565 55020 1585
rect 55020 1565 55038 1585
rect 55038 1565 55045 1585
rect 55015 1560 55045 1565
rect 55125 1585 55155 1590
rect 55125 1565 55130 1585
rect 55130 1565 55148 1585
rect 55148 1565 55155 1585
rect 55125 1560 55155 1565
rect 55235 1585 55265 1590
rect 55235 1565 55240 1585
rect 55240 1565 55258 1585
rect 55258 1565 55265 1585
rect 55235 1560 55265 1565
rect 55345 1585 55375 1590
rect 55345 1565 55350 1585
rect 55350 1565 55368 1585
rect 55368 1565 55375 1585
rect 55345 1560 55375 1565
rect 55455 1585 55485 1590
rect 55455 1565 55460 1585
rect 55460 1565 55478 1585
rect 55478 1565 55485 1585
rect 55455 1560 55485 1565
rect 55565 1585 55595 1590
rect 55565 1565 55570 1585
rect 55570 1565 55588 1585
rect 55588 1565 55595 1585
rect 55565 1560 55595 1565
rect 55790 1560 55820 1590
rect 54595 1505 54625 1535
rect 54795 1505 54825 1535
rect 54475 1455 54505 1485
rect 54730 1395 54760 1425
rect 55440 1395 55470 1425
rect 55745 1395 55775 1425
rect 54320 1340 54350 1370
rect 54795 1340 54825 1370
rect 55140 1365 55170 1370
rect 55140 1345 55145 1365
rect 55145 1345 55165 1365
rect 55165 1345 55170 1365
rect 55140 1340 55170 1345
rect 55340 1365 55370 1370
rect 55340 1345 55345 1365
rect 55345 1345 55365 1365
rect 55365 1345 55370 1365
rect 55340 1340 55370 1345
rect 55540 1365 55570 1370
rect 55540 1345 55545 1365
rect 55545 1345 55565 1365
rect 55565 1345 55570 1365
rect 55540 1340 55570 1345
rect 54730 1305 54765 1310
rect 54730 1280 54735 1305
rect 54735 1280 54760 1305
rect 54760 1280 54765 1305
rect 54730 1275 54765 1280
rect 54790 1305 54825 1310
rect 54790 1280 54795 1305
rect 54795 1280 54820 1305
rect 54820 1280 54825 1305
rect 54790 1275 54825 1280
rect 54880 980 54910 985
rect 54880 960 54885 980
rect 54885 960 54905 980
rect 54905 960 54910 980
rect 54880 955 54910 960
rect 54970 980 55000 985
rect 54970 960 54975 980
rect 54975 960 54995 980
rect 54995 960 55000 980
rect 54970 955 55000 960
rect 55790 905 55820 935
rect 56245 2560 56275 2590
rect 56980 2860 57010 2865
rect 56980 2840 56985 2860
rect 56985 2840 57005 2860
rect 57005 2840 57010 2860
rect 56980 2835 57010 2840
rect 57245 2800 57271 2805
rect 57245 2780 57248 2800
rect 57248 2780 57265 2800
rect 57265 2780 57271 2800
rect 57245 2775 57271 2780
rect 57465 2800 57491 2805
rect 57465 2780 57468 2800
rect 57468 2780 57485 2800
rect 57485 2780 57491 2800
rect 57465 2775 57491 2780
rect 57609 2800 57635 2805
rect 57609 2780 57615 2800
rect 57615 2780 57632 2800
rect 57632 2780 57635 2800
rect 57609 2775 57635 2780
rect 57095 2715 57125 2745
rect 56885 2615 56915 2645
rect 57315 2715 57345 2745
rect 57535 2715 57565 2745
rect 57190 2660 57220 2690
rect 57410 2660 57440 2690
rect 57650 2660 57680 2690
rect 57875 2615 57905 2645
rect 56720 2570 56750 2600
rect 56940 2570 56970 2600
rect 57095 2570 57125 2600
rect 57160 2570 57190 2600
rect 57525 2560 57555 2590
rect 56610 2505 56640 2510
rect 56610 2485 56615 2505
rect 56615 2485 56635 2505
rect 56635 2485 56640 2505
rect 56610 2480 56640 2485
rect 56830 2505 56860 2510
rect 56830 2485 56835 2505
rect 56835 2485 56855 2505
rect 56855 2485 56860 2505
rect 56830 2480 56860 2485
rect 57050 2505 57080 2510
rect 57050 2485 57055 2505
rect 57055 2485 57075 2505
rect 57075 2485 57080 2505
rect 57050 2480 57080 2485
rect 56665 2385 56695 2390
rect 56665 2365 56670 2385
rect 56670 2365 56690 2385
rect 56690 2365 56695 2385
rect 56665 2360 56695 2365
rect 56775 2385 56805 2390
rect 56775 2365 56780 2385
rect 56780 2365 56800 2385
rect 56800 2365 56805 2385
rect 56775 2360 56805 2365
rect 56885 2385 56915 2390
rect 56885 2365 56890 2385
rect 56890 2365 56910 2385
rect 56910 2365 56915 2385
rect 56885 2360 56915 2365
rect 56995 2385 57025 2390
rect 56995 2365 57000 2385
rect 57000 2365 57020 2385
rect 57020 2365 57025 2385
rect 56995 2360 57025 2365
rect 57105 2385 57135 2390
rect 57105 2365 57110 2385
rect 57110 2365 57130 2385
rect 57130 2365 57135 2385
rect 57105 2360 57135 2365
rect 56885 2325 56915 2330
rect 56885 2305 56890 2325
rect 56890 2305 56910 2325
rect 56910 2305 56915 2325
rect 56885 2300 56915 2305
rect 56135 2255 56165 2285
rect 56245 2255 56275 2285
rect 56355 2255 56385 2285
rect 56465 2255 56495 2285
rect 56575 2255 56605 2285
rect 56685 2255 56715 2285
rect 56410 2225 56440 2230
rect 56410 2205 56415 2225
rect 56415 2205 56435 2225
rect 56435 2205 56440 2225
rect 56410 2200 56440 2205
rect 57085 2255 57115 2285
rect 57195 2255 57225 2285
rect 57305 2255 57335 2285
rect 57415 2255 57445 2285
rect 57525 2255 57555 2285
rect 57635 2255 57665 2285
rect 57360 2225 57390 2230
rect 57360 2205 57365 2225
rect 57365 2205 57385 2225
rect 57385 2205 57390 2225
rect 57360 2200 57390 2205
rect 56800 2115 56830 2120
rect 56800 2095 56805 2115
rect 56805 2095 56825 2115
rect 56825 2095 56830 2115
rect 56800 2090 56830 2095
rect 56885 2090 56915 2120
rect 56970 2115 57000 2120
rect 56970 2095 56975 2115
rect 56975 2095 56995 2115
rect 56995 2095 57000 2115
rect 56970 2090 57000 2095
rect 56190 1920 56220 1950
rect 56300 1920 56330 1950
rect 56410 1920 56440 1950
rect 56520 1920 56550 1950
rect 56630 1920 56660 1950
rect 56195 1865 56225 1895
rect 56415 1865 56445 1895
rect 56090 1775 56120 1805
rect 56310 1775 56340 1805
rect 56240 1755 56266 1760
rect 56240 1735 56243 1755
rect 56243 1735 56260 1755
rect 56260 1735 56266 1755
rect 56240 1730 56266 1735
rect 56645 1865 56675 1895
rect 56530 1775 56560 1805
rect 56460 1755 56486 1760
rect 56460 1735 56463 1755
rect 56463 1735 56480 1755
rect 56480 1735 56486 1755
rect 56460 1730 56486 1735
rect 56604 1755 56630 1760
rect 56604 1735 56610 1755
rect 56610 1735 56627 1755
rect 56627 1735 56630 1755
rect 56604 1730 56630 1735
rect 56825 1820 56855 1850
rect 57140 1920 57170 1950
rect 57250 1920 57280 1950
rect 57360 1920 57390 1950
rect 57470 1920 57500 1950
rect 57580 1920 57610 1950
rect 57235 1865 57265 1895
rect 57455 1865 57485 1895
rect 57685 1865 57715 1895
rect 56945 1820 56975 1850
rect 57130 1775 57160 1805
rect 56870 1755 56896 1760
rect 56870 1735 56873 1755
rect 56873 1735 56890 1755
rect 56890 1735 56896 1755
rect 56870 1730 56896 1735
rect 57350 1775 57380 1805
rect 57280 1755 57306 1760
rect 57280 1735 57283 1755
rect 57283 1735 57300 1755
rect 57300 1735 57306 1755
rect 57280 1730 57306 1735
rect 57570 1775 57600 1805
rect 57500 1755 57526 1760
rect 57500 1735 57503 1755
rect 57503 1735 57520 1755
rect 57520 1735 57526 1755
rect 57500 1730 57526 1735
rect 57644 1755 57670 1760
rect 57644 1735 57650 1755
rect 57650 1735 57667 1755
rect 57667 1735 57670 1755
rect 57644 1730 57670 1735
rect 57795 1645 57825 1650
rect 57795 1625 57800 1645
rect 57800 1625 57820 1645
rect 57820 1625 57825 1645
rect 57795 1620 57825 1625
rect 56109 1535 56135 1540
rect 56109 1515 56112 1535
rect 56112 1515 56129 1535
rect 56129 1515 56135 1535
rect 56109 1510 56135 1515
rect 56310 1535 56340 1540
rect 56310 1515 56315 1535
rect 56315 1515 56335 1535
rect 56335 1515 56340 1535
rect 56310 1510 56340 1515
rect 56530 1535 56560 1540
rect 56530 1515 56535 1535
rect 56535 1515 56555 1535
rect 56555 1515 56560 1535
rect 56530 1510 56560 1515
rect 56925 1535 56951 1540
rect 56925 1515 56928 1535
rect 56928 1515 56945 1535
rect 56945 1515 56951 1535
rect 56925 1510 56951 1515
rect 57149 1535 57175 1540
rect 57149 1515 57152 1535
rect 57152 1515 57169 1535
rect 57169 1515 57175 1535
rect 57149 1510 57175 1515
rect 57350 1535 57380 1540
rect 57350 1515 57355 1535
rect 57355 1515 57375 1535
rect 57375 1515 57380 1535
rect 57350 1510 57380 1515
rect 57570 1535 57600 1540
rect 57570 1515 57575 1535
rect 57575 1515 57595 1535
rect 57595 1515 57600 1535
rect 57570 1510 57600 1515
rect 55880 1455 55910 1485
rect 56150 1450 56180 1480
rect 56255 1450 56285 1480
rect 56365 1450 56395 1480
rect 56475 1450 56505 1480
rect 56585 1450 56615 1480
rect 55960 1360 55990 1390
rect 56775 1360 56805 1390
rect 56335 1315 56365 1345
rect 57920 2480 57950 2510
rect 57190 1450 57220 1480
rect 57295 1450 57325 1480
rect 57405 1450 57435 1480
rect 57515 1450 57545 1480
rect 57625 1450 57655 1480
rect 57875 1460 57905 1490
rect 56875 1315 56905 1345
rect 59111 3290 59141 3320
rect 59160 3290 59190 3320
rect 59210 3290 59240 3320
rect 58205 2705 58235 2710
rect 58205 2685 58210 2705
rect 58210 2685 58230 2705
rect 58230 2685 58235 2705
rect 58205 2680 58235 2685
rect 58315 2705 58345 2710
rect 58315 2685 58320 2705
rect 58320 2685 58340 2705
rect 58340 2685 58345 2705
rect 58315 2680 58345 2685
rect 58425 2705 58455 2710
rect 58425 2685 58430 2705
rect 58430 2685 58450 2705
rect 58450 2685 58455 2705
rect 58425 2680 58455 2685
rect 58535 2705 58565 2710
rect 58535 2685 58540 2705
rect 58540 2685 58560 2705
rect 58560 2685 58565 2705
rect 58535 2680 58565 2685
rect 58645 2705 58675 2710
rect 58645 2685 58650 2705
rect 58650 2685 58670 2705
rect 58670 2685 58675 2705
rect 58645 2680 58675 2685
rect 58755 2705 58785 2710
rect 58755 2685 58760 2705
rect 58760 2685 58780 2705
rect 58780 2685 58785 2705
rect 58755 2680 58785 2685
rect 59111 2685 59141 2715
rect 59160 2685 59190 2715
rect 59210 2685 59240 2715
rect 58045 2560 58075 2590
rect 58315 2515 58345 2545
rect 58590 2560 58620 2590
rect 59160 2560 59190 2590
rect 58205 2415 58235 2420
rect 58205 2395 58210 2415
rect 58210 2395 58230 2415
rect 58230 2395 58235 2415
rect 58205 2390 58235 2395
rect 58315 2415 58345 2420
rect 58315 2395 58320 2415
rect 58320 2395 58340 2415
rect 58340 2395 58345 2415
rect 58315 2390 58345 2395
rect 58425 2415 58455 2420
rect 58425 2395 58430 2415
rect 58430 2395 58450 2415
rect 58450 2395 58455 2415
rect 58425 2390 58455 2395
rect 58535 2415 58565 2420
rect 58535 2395 58540 2415
rect 58540 2395 58560 2415
rect 58560 2395 58565 2415
rect 58535 2390 58565 2395
rect 58645 2415 58675 2420
rect 58645 2395 58650 2415
rect 58650 2395 58670 2415
rect 58670 2395 58675 2415
rect 58645 2390 58675 2395
rect 58755 2415 58785 2420
rect 58755 2395 58760 2415
rect 58760 2395 58780 2415
rect 58780 2395 58785 2415
rect 58755 2390 58785 2395
rect 59450 2515 59480 2545
rect 58260 2145 58290 2150
rect 58260 2125 58265 2145
rect 58265 2125 58285 2145
rect 58285 2125 58290 2145
rect 58260 2120 58290 2125
rect 58370 2145 58400 2150
rect 58370 2125 58375 2145
rect 58375 2125 58395 2145
rect 58395 2125 58400 2145
rect 58370 2120 58400 2125
rect 58480 2145 58510 2150
rect 58480 2125 58485 2145
rect 58485 2125 58505 2145
rect 58505 2125 58510 2145
rect 58480 2120 58510 2125
rect 58590 2145 58620 2150
rect 58590 2125 58595 2145
rect 58595 2125 58615 2145
rect 58615 2125 58620 2145
rect 58590 2120 58620 2125
rect 58700 2145 58730 2150
rect 58700 2125 58705 2145
rect 58705 2125 58725 2145
rect 58725 2125 58730 2145
rect 58700 2120 58730 2125
rect 58980 2120 59010 2150
rect 58045 2015 58075 2045
rect 58315 2015 58345 2045
rect 58260 1955 58290 1960
rect 58260 1935 58265 1955
rect 58265 1935 58285 1955
rect 58285 1935 58290 1955
rect 58260 1930 58290 1935
rect 58370 1955 58400 1960
rect 58370 1935 58375 1955
rect 58375 1935 58395 1955
rect 58395 1935 58400 1955
rect 58370 1930 58400 1935
rect 58480 1955 58510 1960
rect 58480 1935 58485 1955
rect 58485 1935 58505 1955
rect 58505 1935 58510 1955
rect 58480 1930 58510 1935
rect 58590 1955 58620 1960
rect 58590 1935 58595 1955
rect 58595 1935 58615 1955
rect 58615 1935 58620 1955
rect 58590 1930 58620 1935
rect 58700 1955 58730 1960
rect 58700 1935 58705 1955
rect 58705 1935 58725 1955
rect 58725 1935 58730 1955
rect 58700 1930 58730 1935
rect 58935 1930 58965 1960
rect 58880 1770 58910 1775
rect 58880 1750 58885 1770
rect 58885 1750 58905 1770
rect 58905 1750 58910 1770
rect 58880 1745 58910 1750
rect 58090 1645 58120 1650
rect 58090 1625 58095 1645
rect 58095 1625 58115 1645
rect 58115 1625 58120 1645
rect 58090 1620 58120 1625
rect 57980 1560 58010 1590
rect 58205 1585 58235 1590
rect 58205 1565 58212 1585
rect 58212 1565 58230 1585
rect 58230 1565 58235 1585
rect 58205 1560 58235 1565
rect 58315 1585 58345 1590
rect 58315 1565 58322 1585
rect 58322 1565 58340 1585
rect 58340 1565 58345 1585
rect 58315 1560 58345 1565
rect 58425 1585 58455 1590
rect 58425 1565 58432 1585
rect 58432 1565 58450 1585
rect 58450 1565 58455 1585
rect 58425 1560 58455 1565
rect 58535 1585 58565 1590
rect 58535 1565 58542 1585
rect 58542 1565 58560 1585
rect 58560 1565 58565 1585
rect 58535 1560 58565 1565
rect 58645 1585 58675 1590
rect 58645 1565 58652 1585
rect 58652 1565 58670 1585
rect 58670 1565 58675 1585
rect 58645 1560 58675 1565
rect 58755 1585 58785 1590
rect 58755 1565 58762 1585
rect 58762 1565 58780 1585
rect 58780 1565 58785 1585
rect 58755 1560 58785 1565
rect 58935 1560 58965 1590
rect 59500 2390 59530 2420
rect 59450 1880 59480 1910
rect 59030 1770 59060 1775
rect 59030 1750 59035 1770
rect 59035 1750 59055 1770
rect 59055 1750 59060 1770
rect 59030 1745 59060 1750
rect 59115 1590 59150 1595
rect 59115 1565 59120 1590
rect 59120 1565 59145 1590
rect 59145 1565 59150 1590
rect 59115 1560 59150 1565
rect 59175 1590 59210 1595
rect 59175 1565 59180 1590
rect 59180 1565 59205 1590
rect 59205 1565 59210 1590
rect 59175 1560 59210 1565
rect 59235 1590 59270 1595
rect 59235 1565 59240 1590
rect 59240 1565 59265 1590
rect 59265 1565 59270 1590
rect 59235 1560 59270 1565
rect 59295 1590 59330 1595
rect 59295 1565 59300 1590
rect 59300 1565 59325 1590
rect 59325 1565 59330 1590
rect 59295 1560 59330 1565
rect 58980 1505 59010 1535
rect 59175 1505 59205 1535
rect 59295 1460 59325 1490
rect 58020 1395 58050 1425
rect 58330 1395 58360 1425
rect 59040 1395 59070 1425
rect 57475 1335 57505 1365
rect 57920 1335 57950 1365
rect 58230 1365 58260 1370
rect 58230 1345 58235 1365
rect 58235 1345 58255 1365
rect 58255 1345 58260 1365
rect 58230 1340 58260 1345
rect 58430 1365 58460 1370
rect 58430 1345 58435 1365
rect 58435 1345 58455 1365
rect 58455 1345 58460 1365
rect 58430 1340 58460 1345
rect 58630 1365 58660 1370
rect 58630 1345 58635 1365
rect 58635 1345 58655 1365
rect 58655 1345 58660 1365
rect 58630 1340 58660 1345
rect 58975 1340 59005 1370
rect 59450 1340 59480 1370
rect 58975 1305 59010 1310
rect 58975 1280 58980 1305
rect 58980 1280 59005 1305
rect 59005 1280 59010 1305
rect 58975 1275 59010 1280
rect 59035 1305 59070 1310
rect 59035 1280 59040 1305
rect 59040 1280 59065 1305
rect 59065 1280 59070 1305
rect 59035 1275 59070 1280
rect 56445 1250 56475 1255
rect 56445 1230 56450 1250
rect 56450 1230 56470 1250
rect 56470 1230 56475 1250
rect 56445 1225 56475 1230
rect 56555 1250 56585 1255
rect 56555 1230 56560 1250
rect 56560 1230 56580 1250
rect 56580 1230 56585 1250
rect 56555 1225 56585 1230
rect 56665 1250 56695 1255
rect 56665 1230 56670 1250
rect 56670 1230 56690 1250
rect 56690 1230 56695 1250
rect 56665 1225 56695 1230
rect 56775 1250 56805 1255
rect 56775 1230 56780 1250
rect 56780 1230 56800 1250
rect 56800 1230 56805 1250
rect 56775 1225 56805 1230
rect 56885 1250 56915 1255
rect 56885 1230 56890 1250
rect 56890 1230 56910 1250
rect 56910 1230 56915 1250
rect 56885 1225 56915 1230
rect 56995 1250 57025 1255
rect 56995 1230 57000 1250
rect 57000 1230 57020 1250
rect 57020 1230 57025 1250
rect 56995 1225 57025 1230
rect 57105 1250 57135 1255
rect 57105 1230 57110 1250
rect 57110 1230 57130 1250
rect 57130 1230 57135 1250
rect 57105 1225 57135 1230
rect 57215 1250 57245 1255
rect 57215 1230 57220 1250
rect 57220 1230 57240 1250
rect 57240 1230 57245 1250
rect 57215 1225 57245 1230
rect 57325 1250 57355 1255
rect 57325 1230 57330 1250
rect 57330 1230 57350 1250
rect 57350 1230 57355 1250
rect 57325 1225 57355 1230
rect 57420 1250 57450 1255
rect 57420 1230 57425 1250
rect 57425 1230 57445 1250
rect 57445 1230 57450 1250
rect 57420 1225 57450 1230
rect 58800 980 58830 985
rect 58800 960 58805 980
rect 58805 960 58825 980
rect 58825 960 58830 980
rect 58800 955 58830 960
rect 58890 980 58920 985
rect 58890 960 58895 980
rect 58895 960 58915 980
rect 58915 960 58920 980
rect 58890 955 58920 960
rect 56215 930 56245 935
rect 56215 910 56220 930
rect 56220 910 56240 930
rect 56240 910 56245 930
rect 56215 905 56245 910
rect 56280 930 56310 935
rect 56280 910 56285 930
rect 56285 910 56305 930
rect 56305 910 56310 930
rect 56280 905 56310 910
rect 56390 930 56420 935
rect 56390 910 56395 930
rect 56395 910 56415 930
rect 56415 910 56420 930
rect 56390 905 56420 910
rect 56500 930 56530 935
rect 56500 910 56505 930
rect 56505 910 56525 930
rect 56525 910 56530 930
rect 56500 905 56530 910
rect 56610 930 56640 935
rect 56610 910 56615 930
rect 56615 910 56635 930
rect 56635 910 56640 930
rect 56610 905 56640 910
rect 56720 930 56750 935
rect 56720 910 56725 930
rect 56725 910 56745 930
rect 56745 910 56750 930
rect 56720 905 56750 910
rect 56830 930 56860 935
rect 56830 910 56835 930
rect 56835 910 56855 930
rect 56855 910 56860 930
rect 56830 905 56860 910
rect 56940 930 56970 935
rect 56940 910 56945 930
rect 56945 910 56965 930
rect 56965 910 56970 930
rect 56940 905 56970 910
rect 57050 930 57080 935
rect 57050 910 57055 930
rect 57055 910 57075 930
rect 57075 910 57080 930
rect 57050 905 57080 910
rect 57160 930 57190 935
rect 57160 910 57165 930
rect 57165 910 57185 930
rect 57185 910 57190 930
rect 57160 905 57190 910
rect 57270 930 57300 935
rect 57270 910 57275 930
rect 57275 910 57295 930
rect 57295 910 57300 930
rect 57270 905 57300 910
rect 57380 930 57410 935
rect 57380 910 57385 930
rect 57385 910 57405 930
rect 57405 910 57410 930
rect 57380 905 57410 910
rect 57490 930 57520 935
rect 57490 910 57495 930
rect 57495 910 57515 930
rect 57515 910 57520 930
rect 57490 905 57520 910
rect 57550 930 57580 935
rect 57550 910 57555 930
rect 57555 910 57575 930
rect 57575 910 57580 930
rect 57550 905 57580 910
rect 57980 895 58010 925
rect 55960 800 55990 830
rect 57060 800 57090 830
rect 55835 710 55865 740
rect 56760 735 56790 740
rect 56760 715 56765 735
rect 56765 715 56785 735
rect 56785 715 56790 735
rect 56760 710 56790 715
rect 56880 735 56910 740
rect 56880 715 56885 735
rect 56885 715 56905 735
rect 56905 715 56910 735
rect 56880 710 56910 715
rect 57000 735 57030 740
rect 57000 715 57005 735
rect 57005 715 57025 735
rect 57025 715 57030 735
rect 57000 710 57030 715
rect 55240 595 55270 600
rect 55240 575 55245 595
rect 55245 575 55265 595
rect 55265 575 55270 595
rect 55240 570 55270 575
rect 55340 570 55370 600
rect 55440 595 55470 600
rect 55440 575 55445 595
rect 55445 575 55465 595
rect 55465 575 55470 595
rect 55440 570 55470 575
rect 55790 570 55820 600
rect 57980 570 58010 600
rect 58330 595 58360 600
rect 58330 575 58335 595
rect 58335 575 58355 595
rect 58355 575 58360 595
rect 58330 570 58360 575
rect 58430 570 58460 600
rect 58530 595 58560 600
rect 58530 575 58535 595
rect 58535 575 58555 595
rect 58555 575 58560 595
rect 58530 570 58560 575
rect 55340 535 55370 540
rect 55340 515 55345 535
rect 55345 515 55365 535
rect 55365 515 55370 535
rect 55340 510 55370 515
rect 58430 535 58460 540
rect 58430 515 58435 535
rect 58435 515 58455 535
rect 58455 515 58460 535
rect 58430 510 58460 515
rect 54270 465 54300 495
rect 55790 465 55820 495
rect 56880 465 56910 495
rect 57980 465 58010 495
rect 59500 465 59530 495
rect 57980 -545 58010 -515
<< metal2 >>
rect 55785 6185 55825 6190
rect 55785 6155 55790 6185
rect 55820 6155 55825 6185
rect 55785 6150 55825 6155
rect 56880 4880 56920 4885
rect 56880 4850 56885 4880
rect 56915 4875 56920 4880
rect 57550 4880 57590 4885
rect 57550 4875 57555 4880
rect 56915 4855 57555 4875
rect 56915 4850 56920 4855
rect 56880 4845 56920 4850
rect 57550 4850 57555 4855
rect 57585 4850 57590 4880
rect 57550 4845 57590 4850
rect 57490 4825 57530 4830
rect 57490 4795 57495 4825
rect 57525 4820 57530 4825
rect 57550 4825 57590 4830
rect 57550 4820 57555 4825
rect 57525 4800 57555 4820
rect 57525 4795 57530 4800
rect 57490 4790 57530 4795
rect 57550 4795 57555 4800
rect 57585 4820 57590 4825
rect 57670 4825 57710 4830
rect 57670 4820 57675 4825
rect 57585 4800 57675 4820
rect 57585 4795 57590 4800
rect 57550 4790 57590 4795
rect 57670 4795 57675 4800
rect 57705 4795 57710 4825
rect 57670 4790 57710 4795
rect 56325 4785 56365 4790
rect 56325 4755 56330 4785
rect 56360 4780 56365 4785
rect 56820 4785 56860 4790
rect 56820 4780 56825 4785
rect 56360 4760 56825 4780
rect 56360 4755 56365 4760
rect 56325 4750 56365 4755
rect 56820 4755 56825 4760
rect 56855 4780 56860 4785
rect 56940 4785 56980 4790
rect 56940 4780 56945 4785
rect 56855 4760 56945 4780
rect 56855 4755 56860 4760
rect 56820 4750 56860 4755
rect 56940 4755 56945 4760
rect 56975 4780 56980 4785
rect 57000 4785 57040 4790
rect 57000 4780 57005 4785
rect 56975 4760 57005 4780
rect 56975 4755 56980 4760
rect 56940 4750 56980 4755
rect 57000 4755 57005 4760
rect 57035 4755 57040 4785
rect 57000 4750 57040 4755
rect 55785 4530 55825 4535
rect 55785 4500 55790 4530
rect 55820 4525 55825 4530
rect 56145 4530 56185 4535
rect 56145 4525 56150 4530
rect 55820 4505 56150 4525
rect 55820 4500 55825 4505
rect 55785 4495 55825 4500
rect 56145 4500 56150 4505
rect 56180 4525 56185 4530
rect 56205 4530 56245 4535
rect 56205 4525 56210 4530
rect 56180 4505 56210 4525
rect 56180 4500 56185 4505
rect 56145 4495 56185 4500
rect 56205 4500 56210 4505
rect 56240 4525 56245 4530
rect 56325 4530 56365 4535
rect 56325 4525 56330 4530
rect 56240 4505 56330 4525
rect 56240 4500 56245 4505
rect 56205 4495 56245 4500
rect 56325 4500 56330 4505
rect 56360 4500 56365 4530
rect 56325 4495 56365 4500
rect 57620 4395 57650 4400
rect 56910 4390 56950 4395
rect 56910 4360 56915 4390
rect 56945 4385 56950 4390
rect 56945 4365 57620 4385
rect 56945 4360 56950 4365
rect 57620 4360 57650 4365
rect 56910 4355 56950 4360
rect 56235 4290 56275 4295
rect 56235 4260 56240 4290
rect 56270 4285 56275 4290
rect 56850 4290 56890 4295
rect 56850 4285 56855 4290
rect 56270 4265 56855 4285
rect 56270 4260 56275 4265
rect 56235 4255 56275 4260
rect 56850 4260 56855 4265
rect 56885 4285 56890 4290
rect 57565 4290 57605 4295
rect 57565 4285 57570 4290
rect 56885 4265 57570 4285
rect 56885 4260 56890 4265
rect 56850 4255 56890 4260
rect 57565 4260 57570 4265
rect 57600 4260 57605 4290
rect 57565 4255 57605 4260
rect 55315 4200 55355 4205
rect 55315 4170 55320 4200
rect 55350 4195 55355 4200
rect 55785 4200 55825 4205
rect 55785 4195 55790 4200
rect 55350 4175 55790 4195
rect 55350 4170 55355 4175
rect 55315 4165 55355 4170
rect 55785 4170 55790 4175
rect 55820 4195 55825 4200
rect 57975 4200 58015 4205
rect 57975 4195 57980 4200
rect 55820 4175 57980 4195
rect 55820 4170 55825 4175
rect 55785 4165 55825 4170
rect 57975 4170 57980 4175
rect 58010 4195 58015 4200
rect 58445 4200 58485 4205
rect 58445 4195 58450 4200
rect 58010 4175 58450 4195
rect 58010 4170 58015 4175
rect 57975 4165 58015 4170
rect 58445 4170 58450 4175
rect 58480 4170 58485 4200
rect 58445 4165 58485 4170
rect 55075 4090 55115 4095
rect 55075 4060 55080 4090
rect 55110 4085 55115 4090
rect 55195 4090 55235 4095
rect 55195 4085 55200 4090
rect 55110 4065 55200 4085
rect 55110 4060 55115 4065
rect 55075 4055 55115 4060
rect 55195 4060 55200 4065
rect 55230 4085 55235 4090
rect 55315 4090 55355 4095
rect 55315 4085 55320 4090
rect 55230 4065 55320 4085
rect 55230 4060 55235 4065
rect 55195 4055 55235 4060
rect 55315 4060 55320 4065
rect 55350 4085 55355 4090
rect 55435 4090 55475 4095
rect 55435 4085 55440 4090
rect 55350 4065 55440 4085
rect 55350 4060 55355 4065
rect 55315 4055 55355 4060
rect 55435 4060 55440 4065
rect 55470 4085 55475 4090
rect 55555 4090 55595 4095
rect 55555 4085 55560 4090
rect 55470 4065 55560 4085
rect 55470 4060 55475 4065
rect 55435 4055 55475 4060
rect 55555 4060 55560 4065
rect 55590 4060 55595 4090
rect 55555 4055 55595 4060
rect 55890 4090 55930 4095
rect 55890 4060 55895 4090
rect 55925 4085 55930 4090
rect 56125 4090 56165 4095
rect 56125 4085 56130 4090
rect 55925 4065 56130 4085
rect 55925 4060 55930 4065
rect 55890 4055 55930 4060
rect 56125 4060 56130 4065
rect 56160 4085 56165 4090
rect 56185 4090 56225 4095
rect 56185 4085 56190 4090
rect 56160 4065 56190 4085
rect 56160 4060 56165 4065
rect 56125 4055 56165 4060
rect 56185 4060 56190 4065
rect 56220 4085 56225 4090
rect 56245 4090 56285 4095
rect 56245 4085 56250 4090
rect 56220 4065 56250 4085
rect 56220 4060 56225 4065
rect 56185 4055 56225 4060
rect 56245 4060 56250 4065
rect 56280 4085 56285 4090
rect 56365 4090 56405 4095
rect 56365 4085 56370 4090
rect 56280 4065 56370 4085
rect 56280 4060 56285 4065
rect 56245 4055 56285 4060
rect 56365 4060 56370 4065
rect 56400 4085 56405 4090
rect 56485 4090 56525 4095
rect 56485 4085 56490 4090
rect 56400 4065 56490 4085
rect 56400 4060 56405 4065
rect 56365 4055 56405 4060
rect 56485 4060 56490 4065
rect 56520 4085 56525 4090
rect 56605 4090 56645 4095
rect 56605 4085 56610 4090
rect 56520 4065 56610 4085
rect 56520 4060 56525 4065
rect 56485 4055 56525 4060
rect 56605 4060 56610 4065
rect 56640 4060 56645 4090
rect 56605 4055 56645 4060
rect 57155 4090 57195 4095
rect 57155 4060 57160 4090
rect 57190 4085 57195 4090
rect 57275 4090 57315 4095
rect 57275 4085 57280 4090
rect 57190 4065 57280 4085
rect 57190 4060 57195 4065
rect 57155 4055 57195 4060
rect 57275 4060 57280 4065
rect 57310 4085 57315 4090
rect 57395 4090 57435 4095
rect 57395 4085 57400 4090
rect 57310 4065 57400 4085
rect 57310 4060 57315 4065
rect 57275 4055 57315 4060
rect 57395 4060 57400 4065
rect 57430 4085 57435 4090
rect 57515 4090 57555 4095
rect 57515 4085 57520 4090
rect 57430 4065 57520 4085
rect 57430 4060 57435 4065
rect 57395 4055 57435 4060
rect 57515 4060 57520 4065
rect 57550 4085 57555 4090
rect 57575 4090 57615 4095
rect 57575 4085 57580 4090
rect 57550 4065 57580 4085
rect 57550 4060 57555 4065
rect 57515 4055 57555 4060
rect 57575 4060 57580 4065
rect 57610 4085 57615 4090
rect 57635 4090 57675 4095
rect 57635 4085 57640 4090
rect 57610 4065 57640 4085
rect 57610 4060 57615 4065
rect 57575 4055 57615 4060
rect 57635 4060 57640 4065
rect 57670 4085 57675 4090
rect 57870 4090 57910 4095
rect 57870 4085 57875 4090
rect 57670 4065 57875 4085
rect 57670 4060 57675 4065
rect 57635 4055 57675 4060
rect 57870 4060 57875 4065
rect 57905 4060 57910 4090
rect 57870 4055 57910 4060
rect 58205 4090 58245 4095
rect 58205 4060 58210 4090
rect 58240 4085 58245 4090
rect 58325 4090 58365 4095
rect 58325 4085 58330 4090
rect 58240 4065 58330 4085
rect 58240 4060 58245 4065
rect 58205 4055 58245 4060
rect 58325 4060 58330 4065
rect 58360 4085 58365 4090
rect 58445 4090 58485 4095
rect 58445 4085 58450 4090
rect 58360 4065 58450 4085
rect 58360 4060 58365 4065
rect 58325 4055 58365 4060
rect 58445 4060 58450 4065
rect 58480 4085 58485 4090
rect 58565 4090 58605 4095
rect 58565 4085 58570 4090
rect 58480 4065 58570 4085
rect 58480 4060 58485 4065
rect 58445 4055 58485 4060
rect 58565 4060 58570 4065
rect 58600 4085 58605 4090
rect 58685 4090 58725 4095
rect 58685 4085 58690 4090
rect 58600 4065 58690 4085
rect 58600 4060 58605 4065
rect 58565 4055 58605 4060
rect 58685 4060 58690 4065
rect 58720 4060 58725 4090
rect 58685 4055 58725 4060
rect 55015 3670 55055 3675
rect 55015 3640 55020 3670
rect 55050 3665 55055 3670
rect 55135 3670 55175 3675
rect 55135 3665 55140 3670
rect 55050 3645 55140 3665
rect 55050 3640 55055 3645
rect 55015 3635 55055 3640
rect 55135 3640 55140 3645
rect 55170 3665 55175 3670
rect 55255 3670 55295 3675
rect 55255 3665 55260 3670
rect 55170 3645 55260 3665
rect 55170 3640 55175 3645
rect 55135 3635 55175 3640
rect 55255 3640 55260 3645
rect 55290 3665 55295 3670
rect 55375 3670 55415 3675
rect 55375 3665 55380 3670
rect 55290 3645 55380 3665
rect 55290 3640 55295 3645
rect 55255 3635 55295 3640
rect 55375 3640 55380 3645
rect 55410 3665 55415 3670
rect 55495 3670 55535 3675
rect 55495 3665 55500 3670
rect 55410 3645 55500 3665
rect 55410 3640 55415 3645
rect 55375 3635 55415 3640
rect 55495 3640 55500 3645
rect 55530 3665 55535 3670
rect 55615 3670 55655 3675
rect 55615 3665 55620 3670
rect 55530 3645 55620 3665
rect 55530 3640 55535 3645
rect 55495 3635 55535 3640
rect 55615 3640 55620 3645
rect 55650 3665 55655 3670
rect 55890 3670 55930 3675
rect 55890 3665 55895 3670
rect 55650 3645 55895 3665
rect 55650 3640 55655 3645
rect 55615 3635 55655 3640
rect 55890 3640 55895 3645
rect 55925 3640 55930 3670
rect 55890 3635 55930 3640
rect 56065 3670 56105 3675
rect 56065 3640 56070 3670
rect 56100 3665 56105 3670
rect 56185 3670 56225 3675
rect 56185 3665 56190 3670
rect 56100 3645 56190 3665
rect 56100 3640 56105 3645
rect 56065 3635 56105 3640
rect 56185 3640 56190 3645
rect 56220 3665 56225 3670
rect 56305 3670 56345 3675
rect 56305 3665 56310 3670
rect 56220 3645 56310 3665
rect 56220 3640 56225 3645
rect 56185 3635 56225 3640
rect 56305 3640 56310 3645
rect 56340 3665 56345 3670
rect 56425 3670 56465 3675
rect 56425 3665 56430 3670
rect 56340 3645 56430 3665
rect 56340 3640 56345 3645
rect 56305 3635 56345 3640
rect 56425 3640 56430 3645
rect 56460 3665 56465 3670
rect 56545 3670 56585 3675
rect 56545 3665 56550 3670
rect 56460 3645 56550 3665
rect 56460 3640 56465 3645
rect 56425 3635 56465 3640
rect 56545 3640 56550 3645
rect 56580 3665 56585 3670
rect 56665 3670 56705 3675
rect 56665 3665 56670 3670
rect 56580 3645 56670 3665
rect 56580 3640 56585 3645
rect 56545 3635 56585 3640
rect 56665 3640 56670 3645
rect 56700 3640 56705 3670
rect 56665 3635 56705 3640
rect 57095 3670 57135 3675
rect 57095 3640 57100 3670
rect 57130 3665 57135 3670
rect 57215 3670 57255 3675
rect 57215 3665 57220 3670
rect 57130 3645 57220 3665
rect 57130 3640 57135 3645
rect 57095 3635 57135 3640
rect 57215 3640 57220 3645
rect 57250 3665 57255 3670
rect 57335 3670 57375 3675
rect 57335 3665 57340 3670
rect 57250 3645 57340 3665
rect 57250 3640 57255 3645
rect 57215 3635 57255 3640
rect 57335 3640 57340 3645
rect 57370 3665 57375 3670
rect 57455 3670 57495 3675
rect 57455 3665 57460 3670
rect 57370 3645 57460 3665
rect 57370 3640 57375 3645
rect 57335 3635 57375 3640
rect 57455 3640 57460 3645
rect 57490 3665 57495 3670
rect 57575 3670 57615 3675
rect 57575 3665 57580 3670
rect 57490 3645 57580 3665
rect 57490 3640 57495 3645
rect 57455 3635 57495 3640
rect 57575 3640 57580 3645
rect 57610 3665 57615 3670
rect 57695 3670 57735 3675
rect 57695 3665 57700 3670
rect 57610 3645 57700 3665
rect 57610 3640 57615 3645
rect 57575 3635 57615 3640
rect 57695 3640 57700 3645
rect 57730 3640 57735 3670
rect 57695 3635 57735 3640
rect 57870 3670 57910 3675
rect 57870 3640 57875 3670
rect 57905 3665 57910 3670
rect 58145 3670 58185 3675
rect 58145 3665 58150 3670
rect 57905 3645 58150 3665
rect 57905 3640 57910 3645
rect 57870 3635 57910 3640
rect 58145 3640 58150 3645
rect 58180 3665 58185 3670
rect 58265 3670 58305 3675
rect 58265 3665 58270 3670
rect 58180 3645 58270 3665
rect 58180 3640 58185 3645
rect 58145 3635 58185 3640
rect 58265 3640 58270 3645
rect 58300 3665 58305 3670
rect 58385 3670 58425 3675
rect 58385 3665 58390 3670
rect 58300 3645 58390 3665
rect 58300 3640 58305 3645
rect 58265 3635 58305 3640
rect 58385 3640 58390 3645
rect 58420 3665 58425 3670
rect 58505 3670 58545 3675
rect 58505 3665 58510 3670
rect 58420 3645 58510 3665
rect 58420 3640 58425 3645
rect 58385 3635 58425 3640
rect 58505 3640 58510 3645
rect 58540 3665 58545 3670
rect 58625 3670 58665 3675
rect 58625 3665 58630 3670
rect 58540 3645 58630 3665
rect 58540 3640 58545 3645
rect 58505 3635 58545 3640
rect 58625 3640 58630 3645
rect 58660 3665 58665 3670
rect 58745 3670 58785 3675
rect 58745 3665 58750 3670
rect 58660 3645 58750 3665
rect 58660 3640 58665 3645
rect 58625 3635 58665 3640
rect 58745 3640 58750 3645
rect 58780 3640 58785 3670
rect 58745 3635 58785 3640
rect 56365 3615 56405 3620
rect 56365 3585 56370 3615
rect 56400 3610 56405 3615
rect 56850 3615 56890 3620
rect 56850 3610 56855 3615
rect 56400 3590 56855 3610
rect 56400 3585 56405 3590
rect 56365 3580 56405 3585
rect 56850 3585 56855 3590
rect 56885 3610 56890 3615
rect 57395 3615 57435 3620
rect 57395 3610 57400 3615
rect 56885 3590 57400 3610
rect 56885 3585 56890 3590
rect 56850 3580 56890 3585
rect 57395 3585 57400 3590
rect 57430 3585 57435 3615
rect 57395 3580 57435 3585
rect 55315 3570 55355 3575
rect 55315 3540 55320 3570
rect 55350 3565 55355 3570
rect 56910 3570 56950 3575
rect 56910 3565 56915 3570
rect 55350 3545 56915 3565
rect 55350 3540 55355 3545
rect 55315 3535 55355 3540
rect 56910 3540 56915 3545
rect 56945 3565 56950 3570
rect 58445 3570 58485 3575
rect 58445 3565 58450 3570
rect 56945 3545 58450 3565
rect 56945 3540 56950 3545
rect 58445 3540 58450 3545
rect 58480 3540 58485 3570
rect 56910 3535 56950 3540
rect 54605 3400 54645 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 59155 3400 59195 3405
rect 54605 3365 54645 3370
rect 54955 3380 54995 3385
rect 54955 3350 54960 3380
rect 54990 3375 54995 3380
rect 55065 3380 55105 3385
rect 55065 3375 55070 3380
rect 54990 3355 55070 3375
rect 54990 3350 54995 3355
rect 54955 3345 54995 3350
rect 55065 3350 55070 3355
rect 55100 3375 55105 3380
rect 55175 3380 55215 3385
rect 55175 3375 55180 3380
rect 55100 3355 55180 3375
rect 55100 3350 55105 3355
rect 55065 3345 55105 3350
rect 55175 3350 55180 3355
rect 55210 3375 55215 3380
rect 55285 3380 55325 3385
rect 55285 3375 55290 3380
rect 55210 3355 55290 3375
rect 55210 3350 55215 3355
rect 55175 3345 55215 3350
rect 55285 3350 55290 3355
rect 55320 3375 55325 3380
rect 55395 3380 55435 3385
rect 55395 3375 55400 3380
rect 55320 3355 55400 3375
rect 55320 3350 55325 3355
rect 55285 3345 55325 3350
rect 55395 3350 55400 3355
rect 55430 3375 55435 3380
rect 55505 3380 55545 3385
rect 55505 3375 55510 3380
rect 55430 3355 55510 3375
rect 55430 3350 55435 3355
rect 55395 3345 55435 3350
rect 55505 3350 55510 3355
rect 55540 3375 55545 3380
rect 55615 3380 55655 3385
rect 55615 3375 55620 3380
rect 55540 3355 55620 3375
rect 55540 3350 55545 3355
rect 55505 3345 55545 3350
rect 55615 3350 55620 3355
rect 55650 3375 55655 3380
rect 55785 3380 55825 3385
rect 55785 3375 55790 3380
rect 55650 3355 55790 3375
rect 55650 3350 55655 3355
rect 55615 3345 55655 3350
rect 55785 3350 55790 3355
rect 55820 3350 55825 3380
rect 55785 3345 55825 3350
rect 56275 3380 56315 3385
rect 56275 3350 56280 3380
rect 56310 3375 56315 3380
rect 56385 3380 56425 3385
rect 56385 3375 56390 3380
rect 56310 3355 56390 3375
rect 56310 3350 56315 3355
rect 56275 3345 56315 3350
rect 56385 3350 56390 3355
rect 56420 3375 56425 3380
rect 56495 3380 56535 3385
rect 56495 3375 56500 3380
rect 56420 3355 56500 3375
rect 56420 3350 56425 3355
rect 56385 3345 56425 3350
rect 56495 3350 56500 3355
rect 56530 3375 56535 3380
rect 56605 3380 56645 3385
rect 56605 3375 56610 3380
rect 56530 3355 56610 3375
rect 56530 3350 56535 3355
rect 56495 3345 56535 3350
rect 56605 3350 56610 3355
rect 56640 3375 56645 3380
rect 56715 3380 56755 3385
rect 56715 3375 56720 3380
rect 56640 3355 56720 3375
rect 56640 3350 56645 3355
rect 56605 3345 56645 3350
rect 56715 3350 56720 3355
rect 56750 3375 56755 3380
rect 56825 3380 56865 3385
rect 56825 3375 56830 3380
rect 56750 3355 56830 3375
rect 56750 3350 56755 3355
rect 56715 3345 56755 3350
rect 56825 3350 56830 3355
rect 56860 3375 56865 3380
rect 56935 3380 56975 3385
rect 56935 3375 56940 3380
rect 56860 3355 56940 3375
rect 56860 3350 56865 3355
rect 56825 3345 56865 3350
rect 56935 3350 56940 3355
rect 56970 3375 56975 3380
rect 57045 3380 57085 3385
rect 57045 3375 57050 3380
rect 56970 3355 57050 3375
rect 56970 3350 56975 3355
rect 56935 3345 56975 3350
rect 57045 3350 57050 3355
rect 57080 3375 57085 3380
rect 57155 3380 57195 3385
rect 57155 3375 57160 3380
rect 57080 3355 57160 3375
rect 57080 3350 57085 3355
rect 57045 3345 57085 3350
rect 57155 3350 57160 3355
rect 57190 3375 57195 3380
rect 57265 3380 57305 3385
rect 57265 3375 57270 3380
rect 57190 3355 57270 3375
rect 57190 3350 57195 3355
rect 57155 3345 57195 3350
rect 57265 3350 57270 3355
rect 57300 3375 57305 3380
rect 57375 3380 57415 3385
rect 57375 3375 57380 3380
rect 57300 3355 57380 3375
rect 57300 3350 57305 3355
rect 57265 3345 57305 3350
rect 57375 3350 57380 3355
rect 57410 3375 57415 3380
rect 57485 3380 57525 3385
rect 57485 3375 57490 3380
rect 57410 3355 57490 3375
rect 57410 3350 57415 3355
rect 57375 3345 57415 3350
rect 57485 3350 57490 3355
rect 57520 3375 57525 3380
rect 57975 3380 58015 3385
rect 57975 3375 57980 3380
rect 57520 3355 57980 3375
rect 57520 3350 57525 3355
rect 57485 3345 57525 3350
rect 57975 3350 57980 3355
rect 58010 3375 58015 3380
rect 58145 3380 58185 3385
rect 58145 3375 58150 3380
rect 58010 3355 58150 3375
rect 58010 3350 58015 3355
rect 57975 3345 58015 3350
rect 58145 3350 58150 3355
rect 58180 3375 58185 3380
rect 58255 3380 58295 3385
rect 58255 3375 58260 3380
rect 58180 3355 58260 3375
rect 58180 3350 58185 3355
rect 58145 3345 58185 3350
rect 58255 3350 58260 3355
rect 58290 3375 58295 3380
rect 58365 3380 58405 3385
rect 58365 3375 58370 3380
rect 58290 3355 58370 3375
rect 58290 3350 58295 3355
rect 58255 3345 58295 3350
rect 58365 3350 58370 3355
rect 58400 3375 58405 3380
rect 58475 3380 58515 3385
rect 58475 3375 58480 3380
rect 58400 3355 58480 3375
rect 58400 3350 58405 3355
rect 58365 3345 58405 3350
rect 58475 3350 58480 3355
rect 58510 3375 58515 3380
rect 58585 3380 58625 3385
rect 58585 3375 58590 3380
rect 58510 3355 58590 3375
rect 58510 3350 58515 3355
rect 58475 3345 58515 3350
rect 58585 3350 58590 3355
rect 58620 3375 58625 3380
rect 58695 3380 58735 3385
rect 58695 3375 58700 3380
rect 58620 3355 58700 3375
rect 58620 3350 58625 3355
rect 58585 3345 58625 3350
rect 58695 3350 58700 3355
rect 58730 3375 58735 3380
rect 58805 3380 58845 3385
rect 58805 3375 58810 3380
rect 58730 3355 58810 3375
rect 58730 3350 58735 3355
rect 58695 3345 58735 3350
rect 58805 3350 58810 3355
rect 58840 3350 58845 3380
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58805 3345 58845 3350
rect 55740 3325 55780 3330
rect 54554 3320 54695 3325
rect 54554 3290 54560 3320
rect 54590 3290 54610 3320
rect 54640 3290 54659 3320
rect 54689 3290 54695 3320
rect 55740 3295 55745 3325
rect 55775 3320 55780 3325
rect 56065 3325 56105 3330
rect 56065 3320 56070 3325
rect 55775 3300 56070 3320
rect 55775 3295 55780 3300
rect 55740 3290 55780 3295
rect 56065 3295 56070 3300
rect 56100 3295 56105 3325
rect 56065 3290 56105 3295
rect 59105 3320 59246 3325
rect 59105 3290 59111 3320
rect 59141 3290 59160 3320
rect 59190 3290 59210 3320
rect 59240 3290 59246 3320
rect 54554 3285 54695 3290
rect 59105 3285 59246 3290
rect 56330 3260 56370 3265
rect 56330 3230 56335 3260
rect 56365 3255 56370 3260
rect 56550 3260 56590 3265
rect 56550 3255 56555 3260
rect 56365 3235 56555 3255
rect 56365 3230 56370 3235
rect 56330 3225 56370 3230
rect 56550 3230 56555 3235
rect 56585 3255 56590 3260
rect 56770 3260 56810 3265
rect 56770 3255 56775 3260
rect 56585 3235 56775 3255
rect 56585 3230 56590 3235
rect 56550 3225 56590 3230
rect 56770 3230 56775 3235
rect 56805 3255 56810 3260
rect 56990 3260 57030 3265
rect 56990 3255 56995 3260
rect 56805 3235 56995 3255
rect 56805 3230 56810 3235
rect 56770 3225 56810 3230
rect 56990 3230 56995 3235
rect 57025 3255 57030 3260
rect 57210 3260 57250 3265
rect 57210 3255 57215 3260
rect 57025 3235 57215 3255
rect 57025 3230 57030 3235
rect 56990 3225 57030 3230
rect 57210 3230 57215 3235
rect 57245 3255 57250 3260
rect 57430 3260 57470 3265
rect 57430 3255 57435 3260
rect 57245 3235 57435 3255
rect 57245 3230 57250 3235
rect 57210 3225 57250 3230
rect 57430 3230 57435 3235
rect 57465 3230 57470 3260
rect 57430 3225 57470 3230
rect 56440 3205 56480 3210
rect 56440 3175 56445 3205
rect 56475 3200 56480 3205
rect 56660 3205 56700 3210
rect 56660 3200 56665 3205
rect 56475 3180 56665 3200
rect 56475 3175 56480 3180
rect 56440 3170 56480 3175
rect 56660 3175 56665 3180
rect 56695 3200 56700 3205
rect 56880 3205 56920 3210
rect 56880 3200 56885 3205
rect 56695 3180 56885 3200
rect 56695 3175 56700 3180
rect 56660 3170 56700 3175
rect 56880 3175 56885 3180
rect 56915 3200 56920 3205
rect 57100 3205 57140 3210
rect 57100 3200 57105 3205
rect 56915 3180 57105 3200
rect 56915 3175 56920 3180
rect 56880 3170 56920 3175
rect 57100 3175 57105 3180
rect 57135 3200 57140 3205
rect 57320 3205 57360 3210
rect 57320 3200 57325 3205
rect 57135 3180 57325 3200
rect 57135 3175 57140 3180
rect 57100 3170 57140 3175
rect 57320 3175 57325 3180
rect 57355 3175 57360 3205
rect 57320 3170 57360 3175
rect 56475 3045 56515 3050
rect 56475 3015 56480 3045
rect 56510 3015 56515 3045
rect 56475 3010 56515 3015
rect 56185 2985 56225 2990
rect 56185 2955 56190 2985
rect 56220 2980 56225 2985
rect 56285 2985 56325 2990
rect 56285 2980 56290 2985
rect 56220 2960 56290 2980
rect 56220 2955 56225 2960
rect 56185 2950 56225 2955
rect 56285 2955 56290 2960
rect 56320 2980 56325 2985
rect 56395 2985 56435 2990
rect 56395 2980 56400 2985
rect 56320 2960 56400 2980
rect 56320 2955 56325 2960
rect 56285 2950 56325 2955
rect 56395 2955 56400 2960
rect 56430 2980 56435 2985
rect 56505 2985 56545 2990
rect 56505 2980 56510 2985
rect 56430 2960 56510 2980
rect 56430 2955 56435 2960
rect 56395 2950 56435 2955
rect 56505 2955 56510 2960
rect 56540 2980 56545 2985
rect 56615 2985 56655 2990
rect 56615 2980 56620 2985
rect 56540 2960 56620 2980
rect 56540 2955 56545 2960
rect 56505 2950 56545 2955
rect 56615 2955 56620 2960
rect 56650 2955 56655 2985
rect 56615 2950 56655 2955
rect 57155 2985 57195 2990
rect 57155 2955 57160 2985
rect 57190 2980 57195 2985
rect 57255 2985 57295 2990
rect 57255 2980 57260 2985
rect 57190 2960 57260 2980
rect 57190 2955 57195 2960
rect 57155 2950 57195 2955
rect 57255 2955 57260 2960
rect 57290 2980 57295 2985
rect 57365 2985 57405 2990
rect 57365 2980 57370 2985
rect 57290 2960 57370 2980
rect 57290 2955 57295 2960
rect 57255 2950 57295 2955
rect 57365 2955 57370 2960
rect 57400 2980 57405 2985
rect 57475 2985 57515 2990
rect 57475 2980 57480 2985
rect 57400 2960 57480 2980
rect 57400 2955 57405 2960
rect 57365 2950 57405 2955
rect 57475 2955 57480 2960
rect 57510 2980 57515 2985
rect 57585 2985 57625 2990
rect 57585 2980 57590 2985
rect 57510 2960 57590 2980
rect 57510 2955 57515 2960
rect 57475 2950 57515 2955
rect 57585 2955 57590 2960
rect 57620 2955 57625 2985
rect 57585 2950 57625 2955
rect 56145 2924 56175 2930
rect 56145 2896 56147 2924
rect 56173 2920 56175 2924
rect 56345 2924 56375 2930
rect 56345 2920 56347 2924
rect 56173 2900 56347 2920
rect 56173 2896 56175 2900
rect 56145 2890 56175 2896
rect 56345 2896 56347 2900
rect 56373 2920 56375 2924
rect 56560 2925 56600 2930
rect 56560 2920 56565 2925
rect 56373 2900 56565 2920
rect 56373 2896 56375 2900
rect 56345 2890 56375 2896
rect 56560 2895 56565 2900
rect 56595 2920 56600 2925
rect 56880 2925 56920 2930
rect 56880 2920 56885 2925
rect 56595 2900 56885 2920
rect 56595 2895 56600 2900
rect 56560 2890 56600 2895
rect 56880 2895 56885 2900
rect 56915 2920 56920 2925
rect 57113 2924 57143 2930
rect 57113 2920 57115 2924
rect 56915 2900 57115 2920
rect 56915 2895 56920 2900
rect 56880 2890 56920 2895
rect 57113 2896 57115 2900
rect 57141 2920 57143 2924
rect 57310 2925 57350 2930
rect 57310 2920 57315 2925
rect 57141 2900 57315 2920
rect 57141 2896 57143 2900
rect 57113 2890 57143 2896
rect 57310 2895 57315 2900
rect 57345 2920 57350 2925
rect 57530 2925 57570 2930
rect 57530 2920 57535 2925
rect 57345 2900 57535 2920
rect 57345 2895 57350 2900
rect 57310 2890 57350 2895
rect 57530 2895 57535 2900
rect 57565 2895 57570 2925
rect 57530 2890 57570 2895
rect 55785 2865 55825 2870
rect 55785 2835 55790 2865
rect 55820 2860 55825 2865
rect 56005 2865 56045 2870
rect 56005 2860 56010 2865
rect 55820 2840 56010 2860
rect 55820 2835 55825 2840
rect 55785 2830 55825 2835
rect 56005 2835 56010 2840
rect 56040 2835 56045 2865
rect 56005 2830 56045 2835
rect 56785 2865 56825 2870
rect 56785 2835 56790 2865
rect 56820 2860 56825 2865
rect 56975 2865 57015 2870
rect 56975 2860 56980 2865
rect 56820 2840 56980 2860
rect 56820 2835 56825 2840
rect 56785 2830 56825 2835
rect 56975 2835 56980 2840
rect 57010 2835 57015 2865
rect 56975 2830 57015 2835
rect 56272 2805 56304 2810
rect 56272 2800 56275 2805
rect 55955 2780 56275 2800
rect 56272 2775 56275 2780
rect 56301 2800 56304 2805
rect 56492 2805 56524 2810
rect 56492 2800 56495 2805
rect 56301 2780 56495 2800
rect 56301 2775 56304 2780
rect 56272 2770 56304 2775
rect 56492 2775 56495 2780
rect 56521 2800 56524 2805
rect 56636 2805 56668 2810
rect 56636 2800 56639 2805
rect 56521 2780 56639 2800
rect 56521 2775 56524 2780
rect 56492 2770 56524 2775
rect 56636 2775 56639 2780
rect 56665 2800 56668 2805
rect 57242 2805 57274 2810
rect 57242 2800 57245 2805
rect 56665 2780 57245 2800
rect 56665 2775 56668 2780
rect 56636 2770 56668 2775
rect 57242 2775 57245 2780
rect 57271 2800 57274 2805
rect 57462 2805 57494 2810
rect 57462 2800 57465 2805
rect 57271 2780 57465 2800
rect 57271 2775 57274 2780
rect 57242 2770 57274 2775
rect 57462 2775 57465 2780
rect 57491 2800 57494 2805
rect 57606 2805 57638 2810
rect 57606 2800 57609 2805
rect 57491 2780 57609 2800
rect 57491 2775 57494 2780
rect 57462 2770 57494 2775
rect 57606 2775 57609 2780
rect 57635 2800 57638 2805
rect 57635 2780 57640 2800
rect 57635 2775 57638 2780
rect 57606 2770 57638 2775
rect 56120 2745 56160 2750
rect 54554 2715 54695 2720
rect 56120 2715 56125 2745
rect 56155 2740 56160 2745
rect 56225 2745 56265 2750
rect 56225 2740 56230 2745
rect 56155 2720 56230 2740
rect 56155 2715 56160 2720
rect 54554 2685 54560 2715
rect 54590 2685 54610 2715
rect 54640 2685 54659 2715
rect 54689 2685 54695 2715
rect 54554 2680 54695 2685
rect 55010 2710 55050 2715
rect 55010 2680 55015 2710
rect 55045 2705 55050 2710
rect 55120 2710 55160 2715
rect 55120 2705 55125 2710
rect 55045 2685 55125 2705
rect 55045 2680 55050 2685
rect 55010 2675 55050 2680
rect 55120 2680 55125 2685
rect 55155 2705 55160 2710
rect 55230 2710 55270 2715
rect 55230 2705 55235 2710
rect 55155 2685 55235 2705
rect 55155 2680 55160 2685
rect 55120 2675 55160 2680
rect 55230 2680 55235 2685
rect 55265 2705 55270 2710
rect 55340 2710 55380 2715
rect 55340 2705 55345 2710
rect 55265 2685 55345 2705
rect 55265 2680 55270 2685
rect 55230 2675 55270 2680
rect 55340 2680 55345 2685
rect 55375 2705 55380 2710
rect 55450 2710 55490 2715
rect 55450 2705 55455 2710
rect 55375 2685 55455 2705
rect 55375 2680 55380 2685
rect 55340 2675 55380 2680
rect 55450 2680 55455 2685
rect 55485 2705 55490 2710
rect 55560 2710 55600 2715
rect 56120 2710 56160 2715
rect 56225 2715 56230 2720
rect 56260 2740 56265 2745
rect 56340 2745 56380 2750
rect 56340 2740 56345 2745
rect 56260 2720 56345 2740
rect 56260 2715 56265 2720
rect 56225 2710 56265 2715
rect 56340 2715 56345 2720
rect 56375 2740 56380 2745
rect 56445 2745 56485 2750
rect 56445 2740 56450 2745
rect 56375 2720 56450 2740
rect 56375 2715 56380 2720
rect 56340 2710 56380 2715
rect 56445 2715 56450 2720
rect 56480 2740 56485 2745
rect 56560 2745 56600 2750
rect 56560 2740 56565 2745
rect 56480 2720 56565 2740
rect 56480 2715 56485 2720
rect 56445 2710 56485 2715
rect 56560 2715 56565 2720
rect 56595 2740 56600 2745
rect 56675 2745 56715 2750
rect 56675 2740 56680 2745
rect 56595 2720 56680 2740
rect 56595 2715 56600 2720
rect 56560 2710 56600 2715
rect 56675 2715 56680 2720
rect 56710 2715 56715 2745
rect 56675 2710 56715 2715
rect 57090 2745 57130 2750
rect 57090 2715 57095 2745
rect 57125 2740 57130 2745
rect 57310 2745 57350 2750
rect 57310 2740 57315 2745
rect 57125 2720 57315 2740
rect 57125 2715 57130 2720
rect 57090 2710 57130 2715
rect 57310 2715 57315 2720
rect 57345 2740 57350 2745
rect 57530 2745 57570 2750
rect 57530 2740 57535 2745
rect 57345 2720 57535 2740
rect 57345 2715 57350 2720
rect 57310 2710 57350 2715
rect 57530 2715 57535 2720
rect 57565 2715 57570 2745
rect 59105 2715 59246 2720
rect 57530 2710 57570 2715
rect 58200 2710 58240 2715
rect 55560 2705 55565 2710
rect 55485 2685 55565 2705
rect 55485 2680 55490 2685
rect 55450 2675 55490 2680
rect 55560 2680 55565 2685
rect 55595 2680 55600 2710
rect 55560 2675 55600 2680
rect 56605 2690 56645 2695
rect 56605 2660 56610 2690
rect 56640 2685 56645 2690
rect 57185 2690 57225 2695
rect 57185 2685 57190 2690
rect 56640 2665 57190 2685
rect 56640 2660 56645 2665
rect 56605 2655 56645 2660
rect 57185 2660 57190 2665
rect 57220 2685 57225 2690
rect 57405 2690 57445 2695
rect 57405 2685 57410 2690
rect 57220 2665 57410 2685
rect 57220 2660 57225 2665
rect 57185 2655 57225 2660
rect 57405 2660 57410 2665
rect 57440 2685 57445 2690
rect 57645 2690 57685 2695
rect 57645 2685 57650 2690
rect 57440 2665 57650 2685
rect 57440 2660 57445 2665
rect 57405 2655 57445 2660
rect 57645 2660 57650 2665
rect 57680 2660 57685 2690
rect 58200 2680 58205 2710
rect 58235 2705 58240 2710
rect 58310 2710 58350 2715
rect 58310 2705 58315 2710
rect 58235 2685 58315 2705
rect 58235 2680 58240 2685
rect 58200 2675 58240 2680
rect 58310 2680 58315 2685
rect 58345 2705 58350 2710
rect 58420 2710 58460 2715
rect 58420 2705 58425 2710
rect 58345 2685 58425 2705
rect 58345 2680 58350 2685
rect 58310 2675 58350 2680
rect 58420 2680 58425 2685
rect 58455 2705 58460 2710
rect 58530 2710 58570 2715
rect 58530 2705 58535 2710
rect 58455 2685 58535 2705
rect 58455 2680 58460 2685
rect 58420 2675 58460 2680
rect 58530 2680 58535 2685
rect 58565 2705 58570 2710
rect 58640 2710 58680 2715
rect 58640 2705 58645 2710
rect 58565 2685 58645 2705
rect 58565 2680 58570 2685
rect 58530 2675 58570 2680
rect 58640 2680 58645 2685
rect 58675 2705 58680 2710
rect 58750 2710 58790 2715
rect 58750 2705 58755 2710
rect 58675 2685 58755 2705
rect 58675 2680 58680 2685
rect 58640 2675 58680 2680
rect 58750 2680 58755 2685
rect 58785 2680 58790 2710
rect 59105 2685 59111 2715
rect 59141 2685 59160 2715
rect 59190 2685 59210 2715
rect 59240 2685 59246 2715
rect 59105 2680 59246 2685
rect 58750 2675 58790 2680
rect 57645 2655 57685 2660
rect 55875 2645 55915 2650
rect 55875 2615 55880 2645
rect 55910 2640 55915 2645
rect 56880 2645 56920 2650
rect 56880 2640 56885 2645
rect 55910 2620 56885 2640
rect 55910 2615 55915 2620
rect 55875 2610 55915 2615
rect 56880 2615 56885 2620
rect 56915 2640 56920 2645
rect 57870 2645 57910 2650
rect 57870 2640 57875 2645
rect 56915 2620 57875 2640
rect 56915 2615 56920 2620
rect 56880 2610 56920 2615
rect 57870 2615 57875 2620
rect 57905 2615 57910 2645
rect 57870 2610 57910 2615
rect 56715 2600 56755 2605
rect 54605 2590 54645 2595
rect 54605 2560 54610 2590
rect 54640 2585 54645 2590
rect 55175 2590 55215 2595
rect 55175 2585 55180 2590
rect 54640 2565 55180 2585
rect 54640 2560 54645 2565
rect 54605 2555 54645 2560
rect 55175 2560 55180 2565
rect 55210 2585 55215 2590
rect 55740 2590 55780 2595
rect 55740 2585 55745 2590
rect 55210 2565 55745 2585
rect 55210 2560 55215 2565
rect 55175 2555 55215 2560
rect 55740 2560 55745 2565
rect 55775 2585 55780 2590
rect 56240 2590 56280 2595
rect 56240 2585 56245 2590
rect 55775 2565 56245 2585
rect 55775 2560 55780 2565
rect 55740 2555 55780 2560
rect 56240 2560 56245 2565
rect 56275 2560 56280 2590
rect 56715 2570 56720 2600
rect 56750 2595 56755 2600
rect 56935 2600 56975 2605
rect 56935 2595 56940 2600
rect 56750 2575 56940 2595
rect 56750 2570 56755 2575
rect 56715 2565 56755 2570
rect 56935 2570 56940 2575
rect 56970 2595 56975 2600
rect 57090 2600 57130 2605
rect 57090 2595 57095 2600
rect 56970 2575 57095 2595
rect 56970 2570 56975 2575
rect 56935 2565 56975 2570
rect 57090 2570 57095 2575
rect 57125 2595 57130 2600
rect 57155 2600 57195 2605
rect 57155 2595 57160 2600
rect 57125 2575 57160 2595
rect 57125 2570 57130 2575
rect 57090 2565 57130 2570
rect 57155 2570 57160 2575
rect 57190 2570 57195 2600
rect 57155 2565 57195 2570
rect 57520 2590 57560 2595
rect 56240 2555 56280 2560
rect 57520 2560 57525 2590
rect 57555 2585 57560 2590
rect 58040 2590 58080 2595
rect 58040 2585 58045 2590
rect 57555 2565 58045 2585
rect 57555 2560 57560 2565
rect 57520 2555 57560 2560
rect 58040 2560 58045 2565
rect 58075 2585 58080 2590
rect 58585 2590 58625 2595
rect 58585 2585 58590 2590
rect 58075 2565 58590 2585
rect 58075 2560 58080 2565
rect 58040 2555 58080 2560
rect 58585 2560 58590 2565
rect 58620 2585 58625 2590
rect 59155 2590 59195 2595
rect 59155 2585 59160 2590
rect 58620 2565 59160 2585
rect 58620 2560 58625 2565
rect 58585 2555 58625 2560
rect 59155 2560 59160 2565
rect 59190 2560 59195 2590
rect 59155 2555 59195 2560
rect 54315 2545 54355 2550
rect 54315 2515 54320 2545
rect 54350 2540 54355 2545
rect 55450 2545 55490 2550
rect 55450 2540 55455 2545
rect 54350 2520 55455 2540
rect 54350 2515 54355 2520
rect 54315 2510 54355 2515
rect 55450 2515 55455 2520
rect 55485 2515 55490 2545
rect 58310 2545 58350 2550
rect 58310 2515 58315 2545
rect 58345 2540 58350 2545
rect 59445 2545 59485 2550
rect 59445 2540 59450 2545
rect 58345 2520 59450 2540
rect 58345 2515 58350 2520
rect 55450 2510 55490 2515
rect 56605 2510 56645 2515
rect 56605 2480 56610 2510
rect 56640 2505 56645 2510
rect 56825 2510 56865 2515
rect 56825 2505 56830 2510
rect 56640 2485 56830 2505
rect 56640 2480 56645 2485
rect 56605 2475 56645 2480
rect 56825 2480 56830 2485
rect 56860 2505 56865 2510
rect 57045 2510 57085 2515
rect 57045 2505 57050 2510
rect 56860 2485 57050 2505
rect 56860 2480 56865 2485
rect 56825 2475 56865 2480
rect 57045 2480 57050 2485
rect 57080 2505 57085 2510
rect 57915 2510 57955 2515
rect 58310 2510 58350 2515
rect 59445 2515 59450 2520
rect 59480 2515 59485 2545
rect 59445 2510 59485 2515
rect 57915 2505 57920 2510
rect 57080 2485 57920 2505
rect 57080 2480 57085 2485
rect 57045 2475 57085 2480
rect 57915 2480 57920 2485
rect 57950 2480 57955 2510
rect 57915 2475 57955 2480
rect 54265 2420 54305 2425
rect 54265 2390 54270 2420
rect 54300 2415 54305 2420
rect 55010 2420 55050 2425
rect 55010 2415 55015 2420
rect 54300 2395 55015 2415
rect 54300 2390 54305 2395
rect 54265 2385 54305 2390
rect 55010 2390 55015 2395
rect 55045 2415 55050 2420
rect 55120 2420 55160 2425
rect 55120 2415 55125 2420
rect 55045 2395 55125 2415
rect 55045 2390 55050 2395
rect 55010 2385 55050 2390
rect 55120 2390 55125 2395
rect 55155 2415 55160 2420
rect 55230 2420 55270 2425
rect 55230 2415 55235 2420
rect 55155 2395 55235 2415
rect 55155 2390 55160 2395
rect 55120 2385 55160 2390
rect 55230 2390 55235 2395
rect 55265 2415 55270 2420
rect 55340 2420 55380 2425
rect 55340 2415 55345 2420
rect 55265 2395 55345 2415
rect 55265 2390 55270 2395
rect 55230 2385 55270 2390
rect 55340 2390 55345 2395
rect 55375 2415 55380 2420
rect 55450 2420 55490 2425
rect 55450 2415 55455 2420
rect 55375 2395 55455 2415
rect 55375 2390 55380 2395
rect 55340 2385 55380 2390
rect 55450 2390 55455 2395
rect 55485 2415 55490 2420
rect 55560 2420 55600 2425
rect 55560 2415 55565 2420
rect 55485 2395 55565 2415
rect 55485 2390 55490 2395
rect 55450 2385 55490 2390
rect 55560 2390 55565 2395
rect 55595 2390 55600 2420
rect 58200 2420 58240 2425
rect 55560 2385 55600 2390
rect 56660 2390 56700 2395
rect 56660 2360 56665 2390
rect 56695 2385 56700 2390
rect 56770 2390 56810 2395
rect 56770 2385 56775 2390
rect 56695 2365 56775 2385
rect 56695 2360 56700 2365
rect 56660 2355 56700 2360
rect 56770 2360 56775 2365
rect 56805 2385 56810 2390
rect 56880 2390 56920 2395
rect 56880 2385 56885 2390
rect 56805 2365 56885 2385
rect 56805 2360 56810 2365
rect 56770 2355 56810 2360
rect 56880 2360 56885 2365
rect 56915 2385 56920 2390
rect 56990 2390 57030 2395
rect 56990 2385 56995 2390
rect 56915 2365 56995 2385
rect 56915 2360 56920 2365
rect 56880 2355 56920 2360
rect 56990 2360 56995 2365
rect 57025 2385 57030 2390
rect 57100 2390 57140 2395
rect 57100 2385 57105 2390
rect 57025 2365 57105 2385
rect 57025 2360 57030 2365
rect 56990 2355 57030 2360
rect 57100 2360 57105 2365
rect 57135 2360 57140 2390
rect 58200 2390 58205 2420
rect 58235 2415 58240 2420
rect 58310 2420 58350 2425
rect 58310 2415 58315 2420
rect 58235 2395 58315 2415
rect 58235 2390 58240 2395
rect 58200 2385 58240 2390
rect 58310 2390 58315 2395
rect 58345 2415 58350 2420
rect 58420 2420 58460 2425
rect 58420 2415 58425 2420
rect 58345 2395 58425 2415
rect 58345 2390 58350 2395
rect 58310 2385 58350 2390
rect 58420 2390 58425 2395
rect 58455 2415 58460 2420
rect 58530 2420 58570 2425
rect 58530 2415 58535 2420
rect 58455 2395 58535 2415
rect 58455 2390 58460 2395
rect 58420 2385 58460 2390
rect 58530 2390 58535 2395
rect 58565 2415 58570 2420
rect 58640 2420 58680 2425
rect 58640 2415 58645 2420
rect 58565 2395 58645 2415
rect 58565 2390 58570 2395
rect 58530 2385 58570 2390
rect 58640 2390 58645 2395
rect 58675 2415 58680 2420
rect 58750 2420 58790 2425
rect 58750 2415 58755 2420
rect 58675 2395 58755 2415
rect 58675 2390 58680 2395
rect 58640 2385 58680 2390
rect 58750 2390 58755 2395
rect 58785 2415 58790 2420
rect 59495 2420 59535 2425
rect 59495 2415 59500 2420
rect 58785 2395 59500 2415
rect 58785 2390 58790 2395
rect 58750 2385 58790 2390
rect 59495 2390 59500 2395
rect 59530 2390 59535 2420
rect 59495 2385 59535 2390
rect 57100 2355 57140 2360
rect 56880 2330 56920 2335
rect 56880 2300 56885 2330
rect 56915 2300 56920 2330
rect 56880 2295 56920 2300
rect 56130 2285 56170 2290
rect 56130 2255 56135 2285
rect 56165 2280 56170 2285
rect 56240 2285 56280 2290
rect 56240 2280 56245 2285
rect 56165 2260 56245 2280
rect 56165 2255 56170 2260
rect 56130 2250 56170 2255
rect 56240 2255 56245 2260
rect 56275 2280 56280 2285
rect 56350 2285 56390 2290
rect 56350 2280 56355 2285
rect 56275 2260 56355 2280
rect 56275 2255 56280 2260
rect 56240 2250 56280 2255
rect 56350 2255 56355 2260
rect 56385 2280 56390 2285
rect 56460 2285 56500 2290
rect 56460 2280 56465 2285
rect 56385 2260 56465 2280
rect 56385 2255 56390 2260
rect 56350 2250 56390 2255
rect 56460 2255 56465 2260
rect 56495 2280 56500 2285
rect 56570 2285 56610 2290
rect 56570 2280 56575 2285
rect 56495 2260 56575 2280
rect 56495 2255 56500 2260
rect 56460 2250 56500 2255
rect 56570 2255 56575 2260
rect 56605 2280 56610 2285
rect 56680 2285 56720 2290
rect 56680 2280 56685 2285
rect 56605 2260 56685 2280
rect 56605 2255 56610 2260
rect 56570 2250 56610 2255
rect 56680 2255 56685 2260
rect 56715 2255 56720 2285
rect 56680 2250 56720 2255
rect 57080 2285 57120 2290
rect 57080 2255 57085 2285
rect 57115 2280 57120 2285
rect 57190 2285 57230 2290
rect 57190 2280 57195 2285
rect 57115 2260 57195 2280
rect 57115 2255 57120 2260
rect 57080 2250 57120 2255
rect 57190 2255 57195 2260
rect 57225 2280 57230 2285
rect 57300 2285 57340 2290
rect 57300 2280 57305 2285
rect 57225 2260 57305 2280
rect 57225 2255 57230 2260
rect 57190 2250 57230 2255
rect 57300 2255 57305 2260
rect 57335 2280 57340 2285
rect 57410 2285 57450 2290
rect 57410 2280 57415 2285
rect 57335 2260 57415 2280
rect 57335 2255 57340 2260
rect 57300 2250 57340 2255
rect 57410 2255 57415 2260
rect 57445 2280 57450 2285
rect 57520 2285 57560 2290
rect 57520 2280 57525 2285
rect 57445 2260 57525 2280
rect 57445 2255 57450 2260
rect 57410 2250 57450 2255
rect 57520 2255 57525 2260
rect 57555 2280 57560 2285
rect 57630 2285 57670 2290
rect 57630 2280 57635 2285
rect 57555 2260 57635 2280
rect 57555 2255 57560 2260
rect 57520 2250 57560 2255
rect 57630 2255 57635 2260
rect 57665 2255 57670 2285
rect 57630 2250 57670 2255
rect 55830 2230 55870 2235
rect 55830 2200 55835 2230
rect 55865 2225 55870 2230
rect 56410 2230 56440 2235
rect 55865 2205 56410 2225
rect 55865 2200 55870 2205
rect 55830 2195 55870 2200
rect 57360 2230 57390 2235
rect 56440 2205 56775 2225
rect 57025 2205 57360 2225
rect 56410 2195 56440 2200
rect 57360 2195 57390 2200
rect 54790 2150 54830 2155
rect 54790 2120 54795 2150
rect 54825 2145 54830 2150
rect 55065 2150 55105 2155
rect 55065 2145 55070 2150
rect 54825 2125 55070 2145
rect 54825 2120 54830 2125
rect 54790 2115 54830 2120
rect 55065 2120 55070 2125
rect 55100 2145 55105 2150
rect 55175 2150 55215 2155
rect 55175 2145 55180 2150
rect 55100 2125 55180 2145
rect 55100 2120 55105 2125
rect 55065 2115 55105 2120
rect 55175 2120 55180 2125
rect 55210 2145 55215 2150
rect 55285 2150 55325 2155
rect 55285 2145 55290 2150
rect 55210 2125 55290 2145
rect 55210 2120 55215 2125
rect 55175 2115 55215 2120
rect 55285 2120 55290 2125
rect 55320 2145 55325 2150
rect 55395 2150 55435 2155
rect 55395 2145 55400 2150
rect 55320 2125 55400 2145
rect 55320 2120 55325 2125
rect 55285 2115 55325 2120
rect 55395 2120 55400 2125
rect 55430 2145 55435 2150
rect 55505 2150 55545 2155
rect 55505 2145 55510 2150
rect 55430 2125 55510 2145
rect 55430 2120 55435 2125
rect 55395 2115 55435 2120
rect 55505 2120 55510 2125
rect 55540 2120 55545 2150
rect 58255 2150 58295 2155
rect 55505 2115 55545 2120
rect 56795 2120 56835 2125
rect 56795 2090 56800 2120
rect 56830 2115 56835 2120
rect 56880 2120 56920 2125
rect 56880 2115 56885 2120
rect 56830 2095 56885 2115
rect 56830 2090 56835 2095
rect 56795 2085 56835 2090
rect 56880 2090 56885 2095
rect 56915 2115 56920 2120
rect 56965 2120 57005 2125
rect 56965 2115 56970 2120
rect 56915 2095 56970 2115
rect 56915 2090 56920 2095
rect 56880 2085 56920 2090
rect 56965 2090 56970 2095
rect 57000 2090 57005 2120
rect 58255 2120 58260 2150
rect 58290 2145 58295 2150
rect 58365 2150 58405 2155
rect 58365 2145 58370 2150
rect 58290 2125 58370 2145
rect 58290 2120 58295 2125
rect 58255 2115 58295 2120
rect 58365 2120 58370 2125
rect 58400 2145 58405 2150
rect 58475 2150 58515 2155
rect 58475 2145 58480 2150
rect 58400 2125 58480 2145
rect 58400 2120 58405 2125
rect 58365 2115 58405 2120
rect 58475 2120 58480 2125
rect 58510 2145 58515 2150
rect 58585 2150 58625 2155
rect 58585 2145 58590 2150
rect 58510 2125 58590 2145
rect 58510 2120 58515 2125
rect 58475 2115 58515 2120
rect 58585 2120 58590 2125
rect 58620 2145 58625 2150
rect 58695 2150 58735 2155
rect 58695 2145 58700 2150
rect 58620 2125 58700 2145
rect 58620 2120 58625 2125
rect 58585 2115 58625 2120
rect 58695 2120 58700 2125
rect 58730 2145 58735 2150
rect 58975 2150 59015 2155
rect 58975 2145 58980 2150
rect 58730 2125 58980 2145
rect 58730 2120 58735 2125
rect 58695 2115 58735 2120
rect 58975 2120 58980 2125
rect 59010 2120 59015 2150
rect 58975 2115 59015 2120
rect 56965 2085 57005 2090
rect 55450 2045 55490 2050
rect 55450 2015 55455 2045
rect 55485 2040 55490 2045
rect 55740 2045 55780 2050
rect 55740 2040 55745 2045
rect 55485 2020 55745 2040
rect 55485 2015 55490 2020
rect 55450 2010 55490 2015
rect 55740 2015 55745 2020
rect 55775 2015 55780 2045
rect 55740 2010 55780 2015
rect 58040 2045 58080 2050
rect 58040 2015 58045 2045
rect 58075 2040 58080 2045
rect 58310 2045 58350 2050
rect 58310 2040 58315 2045
rect 58075 2020 58315 2040
rect 58075 2015 58080 2020
rect 58040 2010 58080 2015
rect 58310 2015 58315 2020
rect 58345 2015 58350 2045
rect 58310 2010 58350 2015
rect 54835 1960 54875 1965
rect 54835 1930 54840 1960
rect 54870 1955 54875 1960
rect 55065 1960 55105 1965
rect 55065 1955 55070 1960
rect 54870 1935 55070 1955
rect 54870 1930 54875 1935
rect 54835 1925 54875 1930
rect 55065 1930 55070 1935
rect 55100 1955 55105 1960
rect 55175 1960 55215 1965
rect 55175 1955 55180 1960
rect 55100 1935 55180 1955
rect 55100 1930 55105 1935
rect 55065 1925 55105 1930
rect 55175 1930 55180 1935
rect 55210 1955 55215 1960
rect 55285 1960 55325 1965
rect 55285 1955 55290 1960
rect 55210 1935 55290 1955
rect 55210 1930 55215 1935
rect 55175 1925 55215 1930
rect 55285 1930 55290 1935
rect 55320 1955 55325 1960
rect 55395 1960 55435 1965
rect 55395 1955 55400 1960
rect 55320 1935 55400 1955
rect 55320 1930 55325 1935
rect 55285 1925 55325 1930
rect 55395 1930 55400 1935
rect 55430 1955 55435 1960
rect 55505 1960 55545 1965
rect 55505 1955 55510 1960
rect 55430 1935 55510 1955
rect 55430 1930 55435 1935
rect 55395 1925 55435 1930
rect 55505 1930 55510 1935
rect 55540 1930 55545 1960
rect 58255 1960 58295 1965
rect 55505 1925 55545 1930
rect 56185 1950 56225 1955
rect 56185 1920 56190 1950
rect 56220 1945 56225 1950
rect 56295 1950 56335 1955
rect 56295 1945 56300 1950
rect 56220 1925 56300 1945
rect 56220 1920 56225 1925
rect 54310 1910 54360 1920
rect 56185 1915 56225 1920
rect 56295 1920 56300 1925
rect 56330 1945 56335 1950
rect 56405 1950 56445 1955
rect 56405 1945 56410 1950
rect 56330 1925 56410 1945
rect 56330 1920 56335 1925
rect 56295 1915 56335 1920
rect 56405 1920 56410 1925
rect 56440 1945 56445 1950
rect 56515 1950 56555 1955
rect 56515 1945 56520 1950
rect 56440 1925 56520 1945
rect 56440 1920 56445 1925
rect 56405 1915 56445 1920
rect 56515 1920 56520 1925
rect 56550 1945 56555 1950
rect 56625 1950 56665 1955
rect 56625 1945 56630 1950
rect 56550 1925 56630 1945
rect 56550 1920 56555 1925
rect 56515 1915 56555 1920
rect 56625 1920 56630 1925
rect 56660 1920 56665 1950
rect 56625 1915 56665 1920
rect 57135 1950 57175 1955
rect 57135 1920 57140 1950
rect 57170 1945 57175 1950
rect 57245 1950 57285 1955
rect 57245 1945 57250 1950
rect 57170 1925 57250 1945
rect 57170 1920 57175 1925
rect 57135 1915 57175 1920
rect 57245 1920 57250 1925
rect 57280 1945 57285 1950
rect 57355 1950 57395 1955
rect 57355 1945 57360 1950
rect 57280 1925 57360 1945
rect 57280 1920 57285 1925
rect 57245 1915 57285 1920
rect 57355 1920 57360 1925
rect 57390 1945 57395 1950
rect 57465 1950 57505 1955
rect 57465 1945 57470 1950
rect 57390 1925 57470 1945
rect 57390 1920 57395 1925
rect 57355 1915 57395 1920
rect 57465 1920 57470 1925
rect 57500 1945 57505 1950
rect 57575 1950 57615 1955
rect 57575 1945 57580 1950
rect 57500 1925 57580 1945
rect 57500 1920 57505 1925
rect 57465 1915 57505 1920
rect 57575 1920 57580 1925
rect 57610 1920 57615 1950
rect 58255 1930 58260 1960
rect 58290 1955 58295 1960
rect 58365 1960 58405 1965
rect 58365 1955 58370 1960
rect 58290 1935 58370 1955
rect 58290 1930 58295 1935
rect 58255 1925 58295 1930
rect 58365 1930 58370 1935
rect 58400 1955 58405 1960
rect 58475 1960 58515 1965
rect 58475 1955 58480 1960
rect 58400 1935 58480 1955
rect 58400 1930 58405 1935
rect 58365 1925 58405 1930
rect 58475 1930 58480 1935
rect 58510 1955 58515 1960
rect 58585 1960 58625 1965
rect 58585 1955 58590 1960
rect 58510 1935 58590 1955
rect 58510 1930 58515 1935
rect 58475 1925 58515 1930
rect 58585 1930 58590 1935
rect 58620 1955 58625 1960
rect 58695 1960 58735 1965
rect 58695 1955 58700 1960
rect 58620 1935 58700 1955
rect 58620 1930 58625 1935
rect 58585 1925 58625 1930
rect 58695 1930 58700 1935
rect 58730 1955 58735 1960
rect 58930 1960 58970 1965
rect 58930 1955 58935 1960
rect 58730 1935 58935 1955
rect 58730 1930 58735 1935
rect 58695 1925 58735 1930
rect 58930 1930 58935 1935
rect 58965 1930 58970 1960
rect 58930 1925 58970 1930
rect 57575 1915 57615 1920
rect 54310 1880 54320 1910
rect 54350 1880 54360 1910
rect 59440 1910 59490 1920
rect 54310 1870 54360 1880
rect 56190 1895 56230 1900
rect 56190 1865 56195 1895
rect 56225 1890 56230 1895
rect 56410 1895 56450 1900
rect 56410 1890 56415 1895
rect 56225 1870 56415 1890
rect 56225 1865 56230 1870
rect 56190 1860 56230 1865
rect 56410 1865 56415 1870
rect 56445 1890 56450 1895
rect 56640 1895 56680 1900
rect 56640 1890 56645 1895
rect 56445 1870 56645 1890
rect 56445 1865 56450 1870
rect 56410 1860 56450 1865
rect 56640 1865 56645 1870
rect 56675 1890 56680 1895
rect 57230 1895 57270 1900
rect 57230 1890 57235 1895
rect 56675 1870 57235 1890
rect 56675 1865 56680 1870
rect 56640 1860 56680 1865
rect 57230 1865 57235 1870
rect 57265 1890 57270 1895
rect 57450 1895 57490 1900
rect 57450 1890 57455 1895
rect 57265 1870 57455 1890
rect 57265 1865 57270 1870
rect 57230 1860 57270 1865
rect 57450 1865 57455 1870
rect 57485 1890 57490 1895
rect 57680 1895 57720 1900
rect 57680 1890 57685 1895
rect 57485 1870 57685 1890
rect 57485 1865 57490 1870
rect 57450 1860 57490 1865
rect 57680 1865 57685 1870
rect 57715 1865 57720 1895
rect 59440 1880 59450 1910
rect 59480 1880 59490 1910
rect 59440 1870 59490 1880
rect 57680 1860 57720 1865
rect 56820 1850 56860 1855
rect 56820 1820 56825 1850
rect 56855 1845 56860 1850
rect 56940 1850 56980 1855
rect 56940 1845 56945 1850
rect 56855 1825 56945 1845
rect 56855 1820 56860 1825
rect 56820 1815 56860 1820
rect 56940 1820 56945 1825
rect 56975 1820 56980 1850
rect 56940 1815 56980 1820
rect 56085 1805 56125 1810
rect 54735 1775 54775 1780
rect 54735 1745 54740 1775
rect 54770 1770 54775 1775
rect 54885 1775 54925 1780
rect 54885 1770 54890 1775
rect 54770 1750 54890 1770
rect 54770 1745 54775 1750
rect 54735 1740 54775 1745
rect 54885 1745 54890 1750
rect 54920 1745 54925 1775
rect 56085 1775 56090 1805
rect 56120 1800 56125 1805
rect 56305 1805 56345 1810
rect 56305 1800 56310 1805
rect 56120 1780 56310 1800
rect 56120 1775 56125 1780
rect 56085 1770 56125 1775
rect 56305 1775 56310 1780
rect 56340 1800 56345 1805
rect 56525 1805 56565 1810
rect 56525 1800 56530 1805
rect 56340 1780 56530 1800
rect 56340 1775 56345 1780
rect 56305 1770 56345 1775
rect 56525 1775 56530 1780
rect 56560 1800 56565 1805
rect 57125 1805 57165 1810
rect 57125 1800 57130 1805
rect 56560 1780 57130 1800
rect 56560 1775 56565 1780
rect 56525 1770 56565 1775
rect 57125 1775 57130 1780
rect 57160 1800 57165 1805
rect 57345 1805 57385 1810
rect 57345 1800 57350 1805
rect 57160 1780 57350 1800
rect 57160 1775 57165 1780
rect 57125 1770 57165 1775
rect 57345 1775 57350 1780
rect 57380 1800 57385 1805
rect 57565 1805 57605 1810
rect 57565 1800 57570 1805
rect 57380 1780 57570 1800
rect 57380 1775 57385 1780
rect 57345 1770 57385 1775
rect 57565 1775 57570 1780
rect 57600 1775 57605 1805
rect 57565 1770 57605 1775
rect 58875 1775 58915 1780
rect 56237 1760 56269 1765
rect 56237 1755 56240 1760
rect 54885 1740 54925 1745
rect 55960 1735 56240 1755
rect 56237 1730 56240 1735
rect 56266 1755 56269 1760
rect 56457 1760 56489 1765
rect 56457 1755 56460 1760
rect 56266 1735 56460 1755
rect 56266 1730 56269 1735
rect 56237 1725 56269 1730
rect 56457 1730 56460 1735
rect 56486 1755 56489 1760
rect 56601 1760 56633 1765
rect 56601 1755 56604 1760
rect 56486 1735 56604 1755
rect 56486 1730 56489 1735
rect 56457 1725 56489 1730
rect 56601 1730 56604 1735
rect 56630 1755 56633 1760
rect 56867 1760 56899 1765
rect 56867 1755 56870 1760
rect 56630 1735 56870 1755
rect 56630 1730 56633 1735
rect 56601 1725 56633 1730
rect 56867 1730 56870 1735
rect 56896 1755 56899 1760
rect 57277 1760 57309 1765
rect 57277 1755 57280 1760
rect 56896 1735 57280 1755
rect 56896 1730 56899 1735
rect 56867 1725 56899 1730
rect 57277 1730 57280 1735
rect 57306 1755 57309 1760
rect 57497 1760 57529 1765
rect 57497 1755 57500 1760
rect 57306 1735 57500 1755
rect 57306 1730 57309 1735
rect 57277 1725 57309 1730
rect 57497 1730 57500 1735
rect 57526 1755 57529 1760
rect 57641 1760 57673 1765
rect 57641 1755 57644 1760
rect 57526 1735 57644 1755
rect 57526 1730 57529 1735
rect 57497 1725 57529 1730
rect 57641 1730 57644 1735
rect 57670 1730 57673 1760
rect 58875 1745 58880 1775
rect 58910 1770 58915 1775
rect 59025 1775 59065 1780
rect 59025 1770 59030 1775
rect 58910 1750 59030 1770
rect 58910 1745 58915 1750
rect 58875 1740 58915 1745
rect 59025 1745 59030 1750
rect 59060 1745 59065 1775
rect 59025 1740 59065 1745
rect 57641 1725 57673 1730
rect 57790 1650 57830 1655
rect 57790 1620 57795 1650
rect 57825 1645 57830 1650
rect 58085 1650 58125 1655
rect 58085 1645 58090 1650
rect 57825 1625 58090 1645
rect 57825 1620 57830 1625
rect 57790 1615 57830 1620
rect 58085 1620 58090 1625
rect 58120 1620 58125 1650
rect 58085 1615 58125 1620
rect 54470 1595 54565 1600
rect 54505 1560 54530 1595
rect 54470 1555 54565 1560
rect 54590 1595 54625 1601
rect 54590 1555 54625 1560
rect 54650 1595 54685 1600
rect 59115 1595 59150 1600
rect 54835 1590 54875 1595
rect 54835 1585 54840 1590
rect 54685 1565 54840 1585
rect 54650 1555 54685 1560
rect 54835 1560 54840 1565
rect 54870 1560 54875 1590
rect 54835 1555 54875 1560
rect 55010 1590 55050 1595
rect 55010 1560 55015 1590
rect 55045 1585 55050 1590
rect 55120 1590 55160 1595
rect 55120 1585 55125 1590
rect 55045 1565 55125 1585
rect 55045 1560 55050 1565
rect 55010 1555 55050 1560
rect 55120 1560 55125 1565
rect 55155 1585 55160 1590
rect 55230 1590 55270 1595
rect 55230 1585 55235 1590
rect 55155 1565 55235 1585
rect 55155 1560 55160 1565
rect 55120 1555 55160 1560
rect 55230 1560 55235 1565
rect 55265 1585 55270 1590
rect 55340 1590 55380 1595
rect 55340 1585 55345 1590
rect 55265 1565 55345 1585
rect 55265 1560 55270 1565
rect 55230 1555 55270 1560
rect 55340 1560 55345 1565
rect 55375 1585 55380 1590
rect 55450 1590 55490 1595
rect 55450 1585 55455 1590
rect 55375 1565 55455 1585
rect 55375 1560 55380 1565
rect 55340 1555 55380 1560
rect 55450 1560 55455 1565
rect 55485 1585 55490 1590
rect 55560 1590 55600 1595
rect 55560 1585 55565 1590
rect 55485 1565 55565 1585
rect 55485 1560 55490 1565
rect 55450 1555 55490 1560
rect 55560 1560 55565 1565
rect 55595 1585 55600 1590
rect 55785 1590 55825 1595
rect 55785 1585 55790 1590
rect 55595 1565 55790 1585
rect 55595 1560 55600 1565
rect 55560 1555 55600 1560
rect 55785 1560 55790 1565
rect 55820 1560 55825 1590
rect 55785 1555 55825 1560
rect 57975 1590 58015 1595
rect 57975 1560 57980 1590
rect 58010 1585 58015 1590
rect 58200 1590 58240 1595
rect 58200 1585 58205 1590
rect 58010 1565 58205 1585
rect 58010 1560 58015 1565
rect 57975 1555 58015 1560
rect 58200 1560 58205 1565
rect 58235 1585 58240 1590
rect 58310 1590 58350 1595
rect 58310 1585 58315 1590
rect 58235 1565 58315 1585
rect 58235 1560 58240 1565
rect 58200 1555 58240 1560
rect 58310 1560 58315 1565
rect 58345 1585 58350 1590
rect 58420 1590 58460 1595
rect 58420 1585 58425 1590
rect 58345 1565 58425 1585
rect 58345 1560 58350 1565
rect 58310 1555 58350 1560
rect 58420 1560 58425 1565
rect 58455 1585 58460 1590
rect 58530 1590 58570 1595
rect 58530 1585 58535 1590
rect 58455 1565 58535 1585
rect 58455 1560 58460 1565
rect 58420 1555 58460 1560
rect 58530 1560 58535 1565
rect 58565 1585 58570 1590
rect 58640 1590 58680 1595
rect 58640 1585 58645 1590
rect 58565 1565 58645 1585
rect 58565 1560 58570 1565
rect 58530 1555 58570 1560
rect 58640 1560 58645 1565
rect 58675 1585 58680 1590
rect 58750 1590 58790 1595
rect 58750 1585 58755 1590
rect 58675 1565 58755 1585
rect 58675 1560 58680 1565
rect 58640 1555 58680 1560
rect 58750 1560 58755 1565
rect 58785 1560 58790 1590
rect 58750 1555 58790 1560
rect 58930 1590 58970 1595
rect 58930 1560 58935 1590
rect 58965 1585 58970 1590
rect 58965 1565 59115 1585
rect 58965 1560 58970 1565
rect 58930 1555 58970 1560
rect 59115 1555 59150 1560
rect 59175 1595 59210 1601
rect 59295 1600 59330 1601
rect 59175 1555 59210 1560
rect 59235 1595 59330 1600
rect 59270 1560 59295 1595
rect 59235 1555 59330 1560
rect 56106 1540 56138 1545
rect 54590 1535 54630 1540
rect 54590 1505 54595 1535
rect 54625 1530 54630 1535
rect 54790 1535 54830 1540
rect 56106 1535 56109 1540
rect 54790 1530 54795 1535
rect 54625 1510 54795 1530
rect 54625 1505 54630 1510
rect 54590 1500 54630 1505
rect 54790 1505 54795 1510
rect 54825 1505 54830 1535
rect 55960 1515 56109 1535
rect 56106 1510 56109 1515
rect 56135 1535 56138 1540
rect 56305 1540 56345 1545
rect 56305 1535 56310 1540
rect 56135 1515 56310 1535
rect 56135 1510 56138 1515
rect 56106 1505 56138 1510
rect 56305 1510 56310 1515
rect 56340 1535 56345 1540
rect 56525 1540 56565 1545
rect 56525 1535 56530 1540
rect 56340 1515 56530 1535
rect 56340 1510 56345 1515
rect 56305 1505 56345 1510
rect 56525 1510 56530 1515
rect 56560 1535 56565 1540
rect 56922 1540 56954 1545
rect 56922 1535 56925 1540
rect 56560 1515 56925 1535
rect 56560 1510 56565 1515
rect 56525 1505 56565 1510
rect 56922 1510 56925 1515
rect 56951 1535 56954 1540
rect 57146 1540 57178 1545
rect 57146 1535 57149 1540
rect 56951 1515 57149 1535
rect 56951 1510 56954 1515
rect 56922 1505 56954 1510
rect 57146 1510 57149 1515
rect 57175 1535 57178 1540
rect 57345 1540 57385 1545
rect 57345 1535 57350 1540
rect 57175 1515 57350 1535
rect 57175 1510 57178 1515
rect 57146 1505 57178 1510
rect 57345 1510 57350 1515
rect 57380 1535 57385 1540
rect 57565 1540 57605 1545
rect 57565 1535 57570 1540
rect 57380 1515 57570 1535
rect 57380 1510 57385 1515
rect 57345 1505 57385 1510
rect 57565 1510 57570 1515
rect 57600 1510 57605 1540
rect 57565 1505 57605 1510
rect 58975 1535 59015 1540
rect 58975 1505 58980 1535
rect 59010 1530 59015 1535
rect 59170 1535 59210 1540
rect 59170 1530 59175 1535
rect 59010 1510 59175 1530
rect 59010 1505 59015 1510
rect 54790 1500 54830 1505
rect 58975 1500 59015 1505
rect 59170 1505 59175 1510
rect 59205 1505 59210 1535
rect 59170 1500 59210 1505
rect 57870 1490 57910 1495
rect 54470 1485 54510 1490
rect 54470 1455 54475 1485
rect 54505 1480 54510 1485
rect 55875 1485 55915 1490
rect 55875 1480 55880 1485
rect 54505 1460 55880 1480
rect 54505 1455 54510 1460
rect 54470 1450 54510 1455
rect 55875 1455 55880 1460
rect 55910 1455 55915 1485
rect 55875 1450 55915 1455
rect 56145 1480 56185 1485
rect 56145 1450 56150 1480
rect 56180 1475 56185 1480
rect 56250 1480 56290 1485
rect 56250 1475 56255 1480
rect 56180 1455 56255 1475
rect 56180 1450 56185 1455
rect 56145 1445 56185 1450
rect 56250 1450 56255 1455
rect 56285 1475 56290 1480
rect 56360 1480 56400 1485
rect 56360 1475 56365 1480
rect 56285 1455 56365 1475
rect 56285 1450 56290 1455
rect 56250 1445 56290 1450
rect 56360 1450 56365 1455
rect 56395 1475 56400 1480
rect 56470 1480 56510 1485
rect 56470 1475 56475 1480
rect 56395 1455 56475 1475
rect 56395 1450 56400 1455
rect 56360 1445 56400 1450
rect 56470 1450 56475 1455
rect 56505 1475 56510 1480
rect 56580 1480 56620 1485
rect 56580 1475 56585 1480
rect 56505 1455 56585 1475
rect 56505 1450 56510 1455
rect 56470 1445 56510 1450
rect 56580 1450 56585 1455
rect 56615 1475 56620 1480
rect 57185 1480 57225 1485
rect 57185 1475 57190 1480
rect 56615 1455 57190 1475
rect 56615 1450 56620 1455
rect 56580 1445 56620 1450
rect 57185 1450 57190 1455
rect 57220 1475 57225 1480
rect 57290 1480 57330 1485
rect 57290 1475 57295 1480
rect 57220 1455 57295 1475
rect 57220 1450 57225 1455
rect 57185 1445 57225 1450
rect 57290 1450 57295 1455
rect 57325 1475 57330 1480
rect 57400 1480 57440 1485
rect 57400 1475 57405 1480
rect 57325 1455 57405 1475
rect 57325 1450 57330 1455
rect 57290 1445 57330 1450
rect 57400 1450 57405 1455
rect 57435 1475 57440 1480
rect 57510 1480 57550 1485
rect 57510 1475 57515 1480
rect 57435 1455 57515 1475
rect 57435 1450 57440 1455
rect 57400 1445 57440 1450
rect 57510 1450 57515 1455
rect 57545 1475 57550 1480
rect 57620 1480 57660 1485
rect 57620 1475 57625 1480
rect 57545 1455 57625 1475
rect 57545 1450 57550 1455
rect 57510 1445 57550 1450
rect 57620 1450 57625 1455
rect 57655 1450 57660 1480
rect 57870 1460 57875 1490
rect 57905 1485 57910 1490
rect 59290 1490 59330 1495
rect 59290 1485 59295 1490
rect 57905 1465 59295 1485
rect 57905 1460 57910 1465
rect 57870 1455 57910 1460
rect 59290 1460 59295 1465
rect 59325 1460 59330 1490
rect 59290 1455 59330 1460
rect 57620 1445 57660 1450
rect 54725 1425 54765 1430
rect 54725 1395 54730 1425
rect 54760 1420 54765 1425
rect 55435 1425 55475 1430
rect 55435 1420 55440 1425
rect 54760 1400 55440 1420
rect 54760 1395 54765 1400
rect 54725 1390 54765 1395
rect 55435 1395 55440 1400
rect 55470 1420 55475 1425
rect 55740 1425 58055 1430
rect 55740 1420 55745 1425
rect 55470 1400 55745 1420
rect 55470 1395 55475 1400
rect 55435 1390 55475 1395
rect 55740 1395 55745 1400
rect 55775 1410 58020 1425
rect 55775 1395 55780 1410
rect 58015 1395 58020 1410
rect 58050 1420 58055 1425
rect 58325 1425 58365 1430
rect 58325 1420 58330 1425
rect 58050 1400 58330 1420
rect 58050 1395 58055 1400
rect 55740 1390 55780 1395
rect 55955 1390 55995 1395
rect 54315 1370 54355 1375
rect 54315 1340 54320 1370
rect 54350 1365 54355 1370
rect 54790 1370 54830 1375
rect 54790 1365 54795 1370
rect 54350 1345 54795 1365
rect 54350 1340 54355 1345
rect 54315 1335 54355 1340
rect 54790 1340 54795 1345
rect 54825 1365 54830 1370
rect 55135 1370 55175 1375
rect 55135 1365 55140 1370
rect 54825 1345 55140 1365
rect 54825 1340 54830 1345
rect 54790 1335 54830 1340
rect 55135 1340 55140 1345
rect 55170 1365 55175 1370
rect 55335 1370 55375 1375
rect 55335 1365 55340 1370
rect 55170 1345 55340 1365
rect 55170 1340 55175 1345
rect 55135 1335 55175 1340
rect 55335 1340 55340 1345
rect 55370 1365 55375 1370
rect 55535 1370 55575 1375
rect 55535 1365 55540 1370
rect 55370 1345 55540 1365
rect 55370 1340 55375 1345
rect 55335 1335 55375 1340
rect 55535 1340 55540 1345
rect 55570 1340 55575 1370
rect 55955 1360 55960 1390
rect 55990 1385 55995 1390
rect 56770 1390 56810 1395
rect 58015 1390 58055 1395
rect 58325 1395 58330 1400
rect 58360 1420 58365 1425
rect 59035 1425 59075 1430
rect 59035 1420 59040 1425
rect 58360 1400 59040 1420
rect 58360 1395 58365 1400
rect 58325 1390 58365 1395
rect 59035 1395 59040 1400
rect 59070 1395 59075 1425
rect 59035 1390 59075 1395
rect 56770 1385 56775 1390
rect 55990 1365 56775 1385
rect 55990 1360 55995 1365
rect 55955 1355 55995 1360
rect 56770 1360 56775 1365
rect 56805 1360 56810 1390
rect 58225 1370 58265 1375
rect 56770 1355 56810 1360
rect 57470 1365 57510 1370
rect 55535 1335 55575 1340
rect 56330 1345 56370 1350
rect 56330 1315 56335 1345
rect 56365 1340 56370 1345
rect 56870 1345 56910 1350
rect 56870 1340 56875 1345
rect 56365 1320 56875 1340
rect 56365 1315 56370 1320
rect 54730 1310 54765 1315
rect 54730 1270 54765 1275
rect 54790 1310 54825 1315
rect 56330 1310 56370 1315
rect 56870 1315 56875 1320
rect 56905 1315 56910 1345
rect 57470 1335 57475 1365
rect 57505 1360 57510 1365
rect 57915 1365 57955 1370
rect 57915 1360 57920 1365
rect 57505 1340 57920 1360
rect 57505 1335 57510 1340
rect 57470 1330 57510 1335
rect 57915 1335 57920 1340
rect 57950 1335 57955 1365
rect 58225 1340 58230 1370
rect 58260 1365 58265 1370
rect 58425 1370 58465 1375
rect 58425 1365 58430 1370
rect 58260 1345 58430 1365
rect 58260 1340 58265 1345
rect 58225 1335 58265 1340
rect 58425 1340 58430 1345
rect 58460 1365 58465 1370
rect 58625 1370 58665 1375
rect 58625 1365 58630 1370
rect 58460 1345 58630 1365
rect 58460 1340 58465 1345
rect 58425 1335 58465 1340
rect 58625 1340 58630 1345
rect 58660 1365 58665 1370
rect 58970 1370 59010 1375
rect 58970 1365 58975 1370
rect 58660 1345 58975 1365
rect 58660 1340 58665 1345
rect 58625 1335 58665 1340
rect 58970 1340 58975 1345
rect 59005 1365 59010 1370
rect 59445 1370 59485 1375
rect 59445 1365 59450 1370
rect 59005 1345 59450 1365
rect 59005 1340 59010 1345
rect 58970 1335 59010 1340
rect 59445 1340 59450 1345
rect 59480 1340 59485 1370
rect 59445 1335 59485 1340
rect 57915 1330 57955 1335
rect 56870 1310 56910 1315
rect 58975 1310 59010 1315
rect 54790 1270 54825 1275
rect 58975 1270 59010 1275
rect 59035 1310 59070 1315
rect 59035 1270 59070 1275
rect 56440 1255 56480 1260
rect 56440 1225 56445 1255
rect 56475 1250 56480 1255
rect 56550 1255 56590 1260
rect 56550 1250 56555 1255
rect 56475 1230 56555 1250
rect 56475 1225 56480 1230
rect 56440 1220 56480 1225
rect 56550 1225 56555 1230
rect 56585 1250 56590 1255
rect 56660 1255 56700 1260
rect 56660 1250 56665 1255
rect 56585 1230 56665 1250
rect 56585 1225 56590 1230
rect 56550 1220 56590 1225
rect 56660 1225 56665 1230
rect 56695 1250 56700 1255
rect 56770 1255 56810 1260
rect 56770 1250 56775 1255
rect 56695 1230 56775 1250
rect 56695 1225 56700 1230
rect 56660 1220 56700 1225
rect 56770 1225 56775 1230
rect 56805 1250 56810 1255
rect 56880 1255 56920 1260
rect 56880 1250 56885 1255
rect 56805 1230 56885 1250
rect 56805 1225 56810 1230
rect 56770 1220 56810 1225
rect 56880 1225 56885 1230
rect 56915 1250 56920 1255
rect 56990 1255 57030 1260
rect 56990 1250 56995 1255
rect 56915 1230 56995 1250
rect 56915 1225 56920 1230
rect 56880 1220 56920 1225
rect 56990 1225 56995 1230
rect 57025 1250 57030 1255
rect 57100 1255 57140 1260
rect 57100 1250 57105 1255
rect 57025 1230 57105 1250
rect 57025 1225 57030 1230
rect 56990 1220 57030 1225
rect 57100 1225 57105 1230
rect 57135 1250 57140 1255
rect 57210 1255 57250 1260
rect 57210 1250 57215 1255
rect 57135 1230 57215 1250
rect 57135 1225 57140 1230
rect 57100 1220 57140 1225
rect 57210 1225 57215 1230
rect 57245 1250 57250 1255
rect 57320 1255 57360 1260
rect 57320 1250 57325 1255
rect 57245 1230 57325 1250
rect 57245 1225 57250 1230
rect 57210 1220 57250 1225
rect 57320 1225 57325 1230
rect 57355 1250 57360 1255
rect 57415 1255 57455 1260
rect 57415 1250 57420 1255
rect 57355 1230 57420 1250
rect 57355 1225 57360 1230
rect 57320 1220 57360 1225
rect 57415 1225 57420 1230
rect 57450 1225 57455 1255
rect 57415 1220 57455 1225
rect 54875 985 54915 990
rect 54875 955 54880 985
rect 54910 980 54915 985
rect 54965 985 55005 990
rect 54965 980 54970 985
rect 54910 960 54970 980
rect 54910 955 54915 960
rect 54875 950 54915 955
rect 54965 955 54970 960
rect 55000 955 55005 985
rect 54965 950 55005 955
rect 58795 985 58835 990
rect 58795 955 58800 985
rect 58830 980 58835 985
rect 58885 985 58925 990
rect 58885 980 58890 985
rect 58830 960 58890 980
rect 58830 955 58835 960
rect 58795 950 58835 955
rect 58885 955 58890 960
rect 58920 955 58925 985
rect 58885 950 58925 955
rect 55785 935 55825 940
rect 55785 905 55790 935
rect 55820 930 55825 935
rect 56210 935 56250 940
rect 56210 930 56215 935
rect 55820 910 56215 930
rect 55820 905 55825 910
rect 55785 900 55825 905
rect 56210 905 56215 910
rect 56245 930 56250 935
rect 56275 935 56315 940
rect 56275 930 56280 935
rect 56245 910 56280 930
rect 56245 905 56250 910
rect 56210 900 56250 905
rect 56275 905 56280 910
rect 56310 930 56315 935
rect 56385 935 56425 940
rect 56385 930 56390 935
rect 56310 910 56390 930
rect 56310 905 56315 910
rect 56275 900 56315 905
rect 56385 905 56390 910
rect 56420 930 56425 935
rect 56495 935 56535 940
rect 56495 930 56500 935
rect 56420 910 56500 930
rect 56420 905 56425 910
rect 56385 900 56425 905
rect 56495 905 56500 910
rect 56530 930 56535 935
rect 56605 935 56645 940
rect 56605 930 56610 935
rect 56530 910 56610 930
rect 56530 905 56535 910
rect 56495 900 56535 905
rect 56605 905 56610 910
rect 56640 930 56645 935
rect 56715 935 56755 940
rect 56715 930 56720 935
rect 56640 910 56720 930
rect 56640 905 56645 910
rect 56605 900 56645 905
rect 56715 905 56720 910
rect 56750 930 56755 935
rect 56825 935 56865 940
rect 56825 930 56830 935
rect 56750 910 56830 930
rect 56750 905 56755 910
rect 56715 900 56755 905
rect 56825 905 56830 910
rect 56860 930 56865 935
rect 56935 935 56975 940
rect 56935 930 56940 935
rect 56860 910 56940 930
rect 56860 905 56865 910
rect 56825 900 56865 905
rect 56935 905 56940 910
rect 56970 930 56975 935
rect 57045 935 57085 940
rect 57045 930 57050 935
rect 56970 910 57050 930
rect 56970 905 56975 910
rect 56935 900 56975 905
rect 57045 905 57050 910
rect 57080 930 57085 935
rect 57155 935 57195 940
rect 57155 930 57160 935
rect 57080 910 57160 930
rect 57080 905 57085 910
rect 57045 900 57085 905
rect 57155 905 57160 910
rect 57190 930 57195 935
rect 57265 935 57305 940
rect 57265 930 57270 935
rect 57190 910 57270 930
rect 57190 905 57195 910
rect 57155 900 57195 905
rect 57265 905 57270 910
rect 57300 930 57305 935
rect 57375 935 57415 940
rect 57375 930 57380 935
rect 57300 910 57380 930
rect 57300 905 57305 910
rect 57265 900 57305 905
rect 57375 905 57380 910
rect 57410 930 57415 935
rect 57485 935 57525 940
rect 57485 930 57490 935
rect 57410 910 57490 930
rect 57410 905 57415 910
rect 57375 900 57415 905
rect 57485 905 57490 910
rect 57520 930 57525 935
rect 57545 935 57585 940
rect 57545 930 57550 935
rect 57520 910 57550 930
rect 57520 905 57525 910
rect 57485 900 57525 905
rect 57545 905 57550 910
rect 57580 930 57585 935
rect 57580 925 58015 930
rect 57580 910 57980 925
rect 57580 905 57585 910
rect 57545 900 57585 905
rect 57975 895 57980 910
rect 58010 895 58015 925
rect 57975 890 58015 895
rect 55955 830 55995 835
rect 55955 800 55960 830
rect 55990 825 55995 830
rect 57055 830 57095 835
rect 57055 825 57060 830
rect 55990 805 57060 825
rect 55990 800 55995 805
rect 55955 795 55995 800
rect 57055 800 57060 805
rect 57090 800 57095 830
rect 57055 795 57095 800
rect 55830 740 55870 745
rect 55830 710 55835 740
rect 55865 735 55870 740
rect 56755 740 56795 745
rect 56755 735 56760 740
rect 55865 715 56760 735
rect 55865 710 55870 715
rect 55830 705 55870 710
rect 56755 710 56760 715
rect 56790 735 56795 740
rect 56875 740 56915 745
rect 56875 735 56880 740
rect 56790 715 56880 735
rect 56790 710 56795 715
rect 56755 705 56795 710
rect 56875 710 56880 715
rect 56910 735 56915 740
rect 56995 740 57035 745
rect 56995 735 57000 740
rect 56910 715 57000 735
rect 56910 710 56915 715
rect 56875 705 56915 710
rect 56995 710 57000 715
rect 57030 710 57035 740
rect 56995 705 57035 710
rect 55235 600 55275 605
rect 55235 570 55240 600
rect 55270 595 55275 600
rect 55335 600 55375 605
rect 55335 595 55340 600
rect 55270 575 55340 595
rect 55270 570 55275 575
rect 55235 565 55275 570
rect 55335 570 55340 575
rect 55370 595 55375 600
rect 55435 600 55475 605
rect 55435 595 55440 600
rect 55370 575 55440 595
rect 55370 570 55375 575
rect 55335 565 55375 570
rect 55435 570 55440 575
rect 55470 595 55475 600
rect 55785 600 55825 605
rect 55785 595 55790 600
rect 55470 575 55790 595
rect 55470 570 55475 575
rect 55435 565 55475 570
rect 55785 570 55790 575
rect 55820 570 55825 600
rect 55785 565 55825 570
rect 57975 600 58015 605
rect 57975 570 57980 600
rect 58010 595 58015 600
rect 58325 600 58365 605
rect 58325 595 58330 600
rect 58010 575 58330 595
rect 58010 570 58015 575
rect 57975 565 58015 570
rect 58325 570 58330 575
rect 58360 595 58365 600
rect 58425 600 58465 605
rect 58425 595 58430 600
rect 58360 575 58430 595
rect 58360 570 58365 575
rect 58325 565 58365 570
rect 58425 570 58430 575
rect 58460 595 58465 600
rect 58525 600 58565 605
rect 58525 595 58530 600
rect 58460 575 58530 595
rect 58460 570 58465 575
rect 58425 565 58465 570
rect 58525 570 58530 575
rect 58560 570 58565 600
rect 58525 565 58565 570
rect 55335 540 55375 545
rect 55335 510 55340 540
rect 55370 510 55375 540
rect 55335 505 55375 510
rect 58425 540 58465 545
rect 58425 510 58430 540
rect 58460 510 58465 540
rect 58425 505 58465 510
rect 54265 495 54305 500
rect 54265 465 54270 495
rect 54300 490 54305 495
rect 55785 495 55825 500
rect 55785 490 55790 495
rect 54300 470 55790 490
rect 54300 465 54305 470
rect 54265 460 54305 465
rect 55785 465 55790 470
rect 55820 490 55825 495
rect 56875 495 56915 500
rect 56875 490 56880 495
rect 55820 470 56880 490
rect 55820 465 55825 470
rect 55785 460 55825 465
rect 56875 465 56880 470
rect 56910 490 56915 495
rect 57975 495 58015 500
rect 57975 490 57980 495
rect 56910 470 57980 490
rect 56910 465 56915 470
rect 56875 460 56915 465
rect 57975 465 57980 470
rect 58010 490 58015 495
rect 59495 495 59535 500
rect 59495 490 59500 495
rect 58010 470 59500 490
rect 58010 465 58015 470
rect 57975 460 58015 465
rect 59495 465 59500 470
rect 59530 465 59535 495
rect 59495 460 59535 465
rect 57975 -515 58015 -510
rect 57975 -545 57980 -515
rect 58010 -545 58015 -515
rect 57975 -550 58015 -545
<< via2 >>
rect 55790 6155 55820 6185
rect 54610 3370 54640 3400
rect 59160 3370 59190 3400
rect 54320 1880 54350 1910
rect 59450 1880 59480 1910
rect 57980 -545 58010 -515
<< metal3 >>
rect 55780 6190 55830 6195
rect 55780 6150 55785 6190
rect 55825 6150 55830 6190
rect 55780 6145 55830 6150
rect 52410 5770 52640 5855
rect 52760 5770 52990 5855
rect 53110 5770 53340 5855
rect 52410 5720 53340 5770
rect 52410 5625 52640 5720
rect 52760 5625 52990 5720
rect 53110 5625 53340 5720
rect 53460 5625 53690 5855
rect 53810 5625 54040 5855
rect 54160 5625 54390 5855
rect 54510 5625 54740 5855
rect 54860 5625 55090 5855
rect 55210 5625 55440 5855
rect 55560 5625 55790 5855
rect 55910 5625 56140 5855
rect 56260 5625 56490 5855
rect 56610 5625 56840 5855
rect 56960 5625 57190 5855
rect 57310 5625 57540 5855
rect 57660 5625 57890 5855
rect 58010 5625 58240 5855
rect 58360 5625 58590 5855
rect 58710 5625 58940 5855
rect 59060 5625 59290 5855
rect 59410 5625 59640 5855
rect 59760 5625 59990 5855
rect 60110 5625 60340 5855
rect 60460 5770 60690 5855
rect 60810 5770 61040 5855
rect 61160 5770 61390 5855
rect 60460 5720 61390 5770
rect 60460 5625 60690 5720
rect 60810 5625 61040 5720
rect 61160 5625 61390 5720
rect 53200 5505 53250 5625
rect 53550 5505 53600 5625
rect 53900 5505 53950 5625
rect 54250 5505 54300 5625
rect 54600 5505 54650 5625
rect 54950 5505 55000 5625
rect 55300 5505 55350 5625
rect 55650 5505 55700 5625
rect 56000 5505 56050 5625
rect 56350 5505 56400 5625
rect 56700 5505 56750 5625
rect 57050 5505 57100 5625
rect 57400 5505 57450 5625
rect 57750 5505 57800 5625
rect 58100 5505 58150 5625
rect 58450 5505 58500 5625
rect 58800 5505 58850 5625
rect 59150 5505 59200 5625
rect 59500 5505 59550 5625
rect 59850 5505 59900 5625
rect 60200 5505 60250 5625
rect 60550 5505 60600 5625
rect 52410 5420 52640 5505
rect 52760 5420 52990 5505
rect 53110 5420 53340 5505
rect 53460 5420 53690 5505
rect 53810 5420 54040 5505
rect 54160 5420 54390 5505
rect 54510 5420 54740 5505
rect 54860 5420 55090 5505
rect 55210 5420 55440 5505
rect 55560 5420 55790 5505
rect 55910 5420 56140 5505
rect 56260 5420 56490 5505
rect 56610 5420 56840 5505
rect 52410 5370 56840 5420
rect 52410 5275 52640 5370
rect 52760 5275 52990 5370
rect 53110 5275 53340 5370
rect 53460 5275 53690 5370
rect 53810 5275 54040 5370
rect 54160 5275 54390 5370
rect 54510 5275 54740 5370
rect 54860 5275 55090 5370
rect 55210 5275 55440 5370
rect 55560 5275 55790 5370
rect 55910 5275 56140 5370
rect 56260 5275 56490 5370
rect 56610 5275 56840 5370
rect 56960 5420 57190 5505
rect 57310 5420 57540 5505
rect 57660 5420 57890 5505
rect 58010 5420 58240 5505
rect 58360 5420 58590 5505
rect 58710 5420 58940 5505
rect 59060 5420 59290 5505
rect 59410 5420 59640 5505
rect 59760 5420 59990 5505
rect 60110 5420 60340 5505
rect 60460 5420 60690 5505
rect 60810 5420 61040 5505
rect 61160 5420 61390 5505
rect 56960 5370 61390 5420
rect 56960 5275 57190 5370
rect 57310 5275 57540 5370
rect 57660 5275 57890 5370
rect 58010 5275 58240 5370
rect 58360 5275 58590 5370
rect 58710 5275 58940 5370
rect 59060 5275 59290 5370
rect 59410 5275 59640 5370
rect 59760 5275 59990 5370
rect 60110 5275 60340 5370
rect 60460 5275 60690 5370
rect 60810 5275 61040 5370
rect 61160 5275 61390 5370
rect 53200 5155 53250 5275
rect 54250 5155 54300 5275
rect 54600 5155 54650 5275
rect 54950 5155 55000 5275
rect 55300 5155 55350 5275
rect 55650 5155 55700 5275
rect 56000 5155 56050 5275
rect 56350 5155 56400 5275
rect 56700 5155 56750 5275
rect 57050 5155 57100 5275
rect 57400 5155 57450 5275
rect 57750 5155 57800 5275
rect 58100 5155 58150 5275
rect 58450 5155 58500 5275
rect 58800 5155 58850 5275
rect 59150 5155 59200 5275
rect 59500 5155 59550 5275
rect 60550 5155 60600 5275
rect 52410 5070 52640 5155
rect 52760 5070 52990 5155
rect 53110 5070 53340 5155
rect 53460 5070 53690 5155
rect 53810 5070 54040 5155
rect 52410 5020 54040 5070
rect 52410 4925 52640 5020
rect 52760 4925 52990 5020
rect 53110 4925 53340 5020
rect 53460 4925 53690 5020
rect 53810 4925 54040 5020
rect 54160 4925 54390 5155
rect 54510 4925 54740 5155
rect 54860 4925 55090 5155
rect 55210 4925 55440 5155
rect 55560 4925 55790 5155
rect 55910 4925 56140 5155
rect 56260 4925 56490 5155
rect 56610 4925 56840 5155
rect 56960 4925 57190 5155
rect 57310 4925 57540 5155
rect 57660 4925 57890 5155
rect 58010 4925 58240 5155
rect 58360 4925 58590 5155
rect 58710 4925 58940 5155
rect 59060 4925 59290 5155
rect 59410 4925 59640 5155
rect 59760 5070 59990 5155
rect 60110 5070 60340 5155
rect 60460 5070 60690 5155
rect 60810 5070 61040 5155
rect 61160 5070 61390 5155
rect 59760 5020 61390 5070
rect 59760 4925 59990 5020
rect 60110 4925 60340 5020
rect 60460 4925 60690 5020
rect 60810 4925 61040 5020
rect 61160 4925 61390 5020
rect 53200 4805 53250 4925
rect 54250 4805 54300 4925
rect 54600 4805 54650 4925
rect 54950 4805 55000 4925
rect 55300 4805 55350 4925
rect 58450 4805 58500 4925
rect 58800 4805 58850 4925
rect 59150 4805 59200 4925
rect 59500 4805 59550 4925
rect 60550 4805 60600 4925
rect 52410 4720 52640 4805
rect 52760 4720 52990 4805
rect 53110 4720 53340 4805
rect 53460 4720 53690 4805
rect 53810 4720 54040 4805
rect 52410 4670 54040 4720
rect 52410 4575 52640 4670
rect 52760 4575 52990 4670
rect 53110 4575 53340 4670
rect 53460 4575 53690 4670
rect 53810 4575 54040 4670
rect 54160 4575 54390 4805
rect 54510 4575 54740 4805
rect 54860 4575 55090 4805
rect 55210 4575 55440 4805
rect 58360 4575 58590 4805
rect 58710 4575 58940 4805
rect 59060 4575 59290 4805
rect 59410 4575 59640 4805
rect 59760 4720 59990 4805
rect 60110 4720 60340 4805
rect 60460 4720 60690 4805
rect 60810 4720 61040 4805
rect 61160 4720 61390 4805
rect 59760 4670 61390 4720
rect 59760 4575 59990 4670
rect 60110 4575 60340 4670
rect 60460 4575 60690 4670
rect 60810 4575 61040 4670
rect 61160 4575 61390 4670
rect 53200 4455 53250 4575
rect 54250 4455 54300 4575
rect 54600 4455 54650 4575
rect 54950 4455 55000 4575
rect 55300 4455 55350 4575
rect 58450 4455 58500 4575
rect 58800 4455 58850 4575
rect 59150 4455 59200 4575
rect 59500 4455 59550 4575
rect 60550 4455 60600 4575
rect 52410 4370 52640 4455
rect 52760 4370 52990 4455
rect 53110 4370 53340 4455
rect 53460 4370 53690 4455
rect 53810 4370 54040 4455
rect 52410 4320 54040 4370
rect 52410 4225 52640 4320
rect 52760 4225 52990 4320
rect 53110 4225 53340 4320
rect 53460 4225 53690 4320
rect 53810 4225 54040 4320
rect 54160 4225 54390 4455
rect 54510 4225 54740 4455
rect 54860 4225 55090 4455
rect 55210 4225 55440 4455
rect 58360 4225 58590 4455
rect 58710 4225 58940 4455
rect 59060 4225 59290 4455
rect 59410 4225 59640 4455
rect 59760 4370 59990 4455
rect 60110 4370 60340 4455
rect 60460 4370 60690 4455
rect 60810 4370 61040 4455
rect 61160 4370 61390 4455
rect 59760 4320 61390 4370
rect 59760 4225 59990 4320
rect 60110 4225 60340 4320
rect 60460 4225 60690 4320
rect 60810 4225 61040 4320
rect 61160 4225 61390 4320
rect 53200 4105 53250 4225
rect 52410 4020 52640 4105
rect 52760 4020 52990 4105
rect 53110 4020 53340 4105
rect 53460 4020 53690 4105
rect 53810 4020 54040 4105
rect 52410 3970 54040 4020
rect 52410 3875 52640 3970
rect 52760 3875 52990 3970
rect 53110 3875 53340 3970
rect 53460 3875 53690 3970
rect 53810 3875 54040 3970
rect 53200 3755 53250 3875
rect 52410 3670 52640 3755
rect 52760 3670 52990 3755
rect 53110 3670 53340 3755
rect 53460 3670 53690 3755
rect 53810 3670 54040 3755
rect 52410 3620 54040 3670
rect 52410 3525 52640 3620
rect 52760 3525 52990 3620
rect 53110 3525 53340 3620
rect 53460 3525 53690 3620
rect 53810 3525 54040 3620
rect 53200 3405 53250 3525
rect 52410 3320 52640 3405
rect 52760 3320 52990 3405
rect 53110 3320 53340 3405
rect 53460 3320 53690 3405
rect 53810 3320 54040 3405
rect 54605 3400 54645 4225
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 59155 3400 59195 4225
rect 60550 4105 60600 4225
rect 59760 4020 59990 4105
rect 60110 4020 60340 4105
rect 60460 4020 60690 4105
rect 60810 4020 61040 4105
rect 61160 4020 61390 4105
rect 59760 3970 61390 4020
rect 59760 3875 59990 3970
rect 60110 3875 60340 3970
rect 60460 3875 60690 3970
rect 60810 3875 61040 3970
rect 61160 3875 61390 3970
rect 60550 3755 60600 3875
rect 59760 3670 59990 3755
rect 60110 3670 60340 3755
rect 60460 3670 60690 3755
rect 60810 3670 61040 3755
rect 61160 3670 61390 3755
rect 59760 3620 61390 3670
rect 59760 3525 59990 3620
rect 60110 3525 60340 3620
rect 60460 3525 60690 3620
rect 60810 3525 61040 3620
rect 61160 3525 61390 3620
rect 60550 3405 60600 3525
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 52410 3270 54040 3320
rect 52410 3175 52640 3270
rect 52760 3175 52990 3270
rect 53110 3175 53340 3270
rect 53460 3175 53690 3270
rect 53810 3175 54040 3270
rect 59760 3320 59990 3405
rect 60110 3320 60340 3405
rect 60460 3320 60690 3405
rect 60810 3320 61040 3405
rect 61160 3320 61390 3405
rect 59760 3270 61390 3320
rect 59760 3175 59990 3270
rect 60110 3175 60340 3270
rect 60460 3175 60690 3270
rect 60810 3175 61040 3270
rect 61160 3175 61390 3270
rect 53200 3055 53250 3175
rect 60550 3055 60600 3175
rect 52410 2970 52640 3055
rect 52760 2970 52990 3055
rect 53110 2970 53340 3055
rect 53460 2970 53690 3055
rect 53810 2970 54040 3055
rect 52410 2920 54040 2970
rect 52410 2825 52640 2920
rect 52760 2825 52990 2920
rect 53110 2825 53340 2920
rect 53460 2825 53690 2920
rect 53810 2825 54040 2920
rect 59760 2970 59990 3055
rect 60110 2970 60340 3055
rect 60460 2970 60690 3055
rect 60810 2970 61040 3055
rect 61160 2970 61390 3055
rect 59760 2920 61390 2970
rect 59760 2825 59990 2920
rect 60110 2825 60340 2920
rect 60460 2825 60690 2920
rect 60810 2825 61040 2920
rect 61160 2825 61390 2920
rect 53200 2705 53250 2825
rect 60550 2705 60600 2825
rect 52410 2620 52640 2705
rect 52760 2620 52990 2705
rect 53110 2620 53340 2705
rect 53460 2620 53690 2705
rect 53810 2620 54040 2705
rect 52410 2570 54040 2620
rect 52410 2475 52640 2570
rect 52760 2475 52990 2570
rect 53110 2475 53340 2570
rect 53460 2475 53690 2570
rect 53810 2475 54040 2570
rect 59760 2620 59990 2705
rect 60110 2620 60340 2705
rect 60460 2620 60690 2705
rect 60810 2620 61040 2705
rect 61160 2620 61390 2705
rect 59760 2570 61390 2620
rect 59760 2475 59990 2570
rect 60110 2475 60340 2570
rect 60460 2475 60690 2570
rect 60810 2475 61040 2570
rect 61160 2475 61390 2570
rect 53200 2355 53250 2475
rect 60550 2355 60600 2475
rect 52410 2270 52640 2355
rect 52760 2270 52990 2355
rect 53110 2270 53340 2355
rect 53460 2270 53690 2355
rect 53810 2270 54040 2355
rect 52410 2220 54040 2270
rect 52410 2125 52640 2220
rect 52760 2125 52990 2220
rect 53110 2125 53340 2220
rect 53460 2125 53690 2220
rect 53810 2125 54040 2220
rect 59760 2270 59990 2355
rect 60110 2270 60340 2355
rect 60460 2270 60690 2355
rect 60810 2270 61040 2355
rect 61160 2270 61390 2355
rect 59760 2220 61390 2270
rect 59760 2125 59990 2220
rect 60110 2125 60340 2220
rect 60460 2125 60690 2220
rect 60810 2125 61040 2220
rect 61160 2125 61390 2220
rect 53200 2005 53250 2125
rect 60550 2005 60600 2125
rect 52410 1920 52640 2005
rect 52760 1920 52990 2005
rect 53110 1920 53340 2005
rect 53460 1920 53690 2005
rect 53810 1920 54040 2005
rect 59760 1920 59990 2005
rect 60110 1920 60340 2005
rect 60460 1920 60690 2005
rect 60810 1920 61040 2005
rect 61160 1920 61390 2005
rect 52410 1870 54040 1920
rect 54310 1915 54360 1920
rect 54310 1875 54315 1915
rect 54355 1875 54360 1915
rect 54310 1870 54360 1875
rect 59440 1915 59490 1920
rect 59440 1875 59445 1915
rect 59485 1875 59490 1915
rect 59440 1870 59490 1875
rect 59760 1870 61390 1920
rect 52410 1775 52640 1870
rect 52760 1775 52990 1870
rect 53110 1775 53340 1870
rect 53460 1775 53690 1870
rect 53810 1775 54040 1870
rect 59760 1775 59990 1870
rect 60110 1775 60340 1870
rect 60460 1775 60690 1870
rect 60810 1775 61040 1870
rect 61160 1775 61390 1870
rect 53200 1655 53250 1775
rect 60550 1655 60600 1775
rect 52410 1570 52640 1655
rect 52760 1570 52990 1655
rect 53110 1570 53340 1655
rect 53460 1570 53690 1655
rect 53810 1570 54040 1655
rect 52410 1520 54040 1570
rect 52410 1425 52640 1520
rect 52760 1425 52990 1520
rect 53110 1425 53340 1520
rect 53460 1425 53690 1520
rect 53810 1425 54040 1520
rect 59760 1570 59990 1655
rect 60110 1570 60340 1655
rect 60460 1570 60690 1655
rect 60810 1570 61040 1655
rect 61160 1570 61390 1655
rect 59760 1520 61390 1570
rect 59760 1425 59990 1520
rect 60110 1425 60340 1520
rect 60460 1425 60690 1520
rect 60810 1425 61040 1520
rect 61160 1425 61390 1520
rect 53200 1305 53250 1425
rect 60550 1305 60600 1425
rect 52410 1220 52640 1305
rect 52760 1220 52990 1305
rect 53110 1220 53340 1305
rect 53460 1220 53690 1305
rect 53810 1220 54040 1305
rect 52410 1170 54040 1220
rect 52410 1075 52640 1170
rect 52760 1075 52990 1170
rect 53110 1075 53340 1170
rect 53460 1075 53690 1170
rect 53810 1075 54040 1170
rect 59760 1220 59990 1305
rect 60110 1220 60340 1305
rect 60460 1220 60690 1305
rect 60810 1220 61040 1305
rect 61160 1220 61390 1305
rect 59760 1170 61390 1220
rect 59760 1075 59990 1170
rect 60110 1075 60340 1170
rect 60460 1075 60690 1170
rect 60810 1075 61040 1170
rect 61160 1075 61390 1170
rect 53200 955 53250 1075
rect 60550 955 60600 1075
rect 52410 870 52640 955
rect 52760 870 52990 955
rect 53110 870 53340 955
rect 53460 870 53690 955
rect 53810 870 54040 955
rect 52410 820 54040 870
rect 52410 725 52640 820
rect 52760 725 52990 820
rect 53110 725 53340 820
rect 53460 725 53690 820
rect 53810 725 54040 820
rect 59760 870 59990 955
rect 60110 870 60340 955
rect 60460 870 60690 955
rect 60810 870 61040 955
rect 61160 870 61390 955
rect 59760 820 61390 870
rect 59760 725 59990 820
rect 60110 725 60340 820
rect 60460 725 60690 820
rect 60810 725 61040 820
rect 61160 725 61390 820
rect 53200 605 53250 725
rect 60550 605 60600 725
rect 52410 520 52640 605
rect 52760 520 52990 605
rect 53110 520 53340 605
rect 53460 520 53690 605
rect 53810 520 54040 605
rect 52410 470 54040 520
rect 52410 375 52640 470
rect 52760 375 52990 470
rect 53110 375 53340 470
rect 53460 375 53690 470
rect 53810 375 54040 470
rect 59760 520 59990 605
rect 60110 520 60340 605
rect 60460 520 60690 605
rect 60810 520 61040 605
rect 61160 520 61390 605
rect 59760 470 61390 520
rect 59760 375 59990 470
rect 60110 375 60340 470
rect 60460 375 60690 470
rect 60810 375 61040 470
rect 61160 375 61390 470
rect 53200 255 53250 375
rect 60550 255 60600 375
rect 52410 170 52640 255
rect 52760 170 52990 255
rect 53110 170 53340 255
rect 53460 170 53690 255
rect 53810 170 54040 255
rect 54160 170 54390 255
rect 54510 170 54740 255
rect 54860 170 55090 255
rect 55210 170 55440 255
rect 55560 170 55790 255
rect 55910 170 56140 255
rect 56260 170 56490 255
rect 56610 170 56840 255
rect 52410 120 56840 170
rect 52410 25 52640 120
rect 52760 25 52990 120
rect 53110 25 53340 120
rect 53460 25 53690 120
rect 53810 25 54040 120
rect 54160 25 54390 120
rect 54510 25 54740 120
rect 54860 25 55090 120
rect 55210 25 55440 120
rect 55560 25 55790 120
rect 55910 25 56140 120
rect 56260 25 56490 120
rect 56610 25 56840 120
rect 56960 170 57190 255
rect 57310 170 57540 255
rect 57660 170 57890 255
rect 58010 170 58240 255
rect 58360 170 58590 255
rect 58710 170 58940 255
rect 59060 170 59290 255
rect 59410 170 59640 255
rect 59760 170 59990 255
rect 60110 170 60340 255
rect 60460 170 60690 255
rect 60810 170 61040 255
rect 61160 170 61390 255
rect 56960 120 61390 170
rect 56960 25 57190 120
rect 57310 25 57540 120
rect 57660 25 57890 120
rect 58010 25 58240 120
rect 58360 25 58590 120
rect 58710 25 58940 120
rect 59060 25 59290 120
rect 59410 25 59640 120
rect 59760 25 59990 120
rect 60110 25 60340 120
rect 60460 25 60690 120
rect 60810 25 61040 120
rect 61160 25 61390 120
rect 53200 -95 53250 25
rect 53550 -95 53600 25
rect 53900 -95 53950 25
rect 54250 -95 54300 25
rect 54600 -95 54650 25
rect 54950 -95 55000 25
rect 55300 -95 55350 25
rect 55650 -95 55700 25
rect 56000 -95 56050 25
rect 56350 -95 56400 25
rect 56700 -95 56750 25
rect 57050 -95 57100 25
rect 57400 -95 57450 25
rect 57750 -95 57800 25
rect 58100 -95 58150 25
rect 58450 -95 58500 25
rect 58800 -95 58850 25
rect 59150 -95 59200 25
rect 59500 -95 59550 25
rect 59850 -95 59900 25
rect 60200 -95 60250 25
rect 60550 -95 60600 25
rect 52410 -180 52640 -95
rect 52760 -180 52990 -95
rect 53110 -180 53340 -95
rect 52410 -230 53340 -180
rect 52410 -325 52640 -230
rect 52760 -325 52990 -230
rect 53110 -325 53340 -230
rect 53460 -325 53690 -95
rect 53810 -325 54040 -95
rect 54160 -325 54390 -95
rect 54510 -325 54740 -95
rect 54860 -325 55090 -95
rect 55210 -325 55440 -95
rect 55560 -325 55790 -95
rect 55910 -325 56140 -95
rect 56260 -325 56490 -95
rect 56610 -325 56840 -95
rect 56960 -325 57190 -95
rect 57310 -325 57540 -95
rect 57660 -325 57890 -95
rect 58010 -325 58240 -95
rect 58360 -325 58590 -95
rect 58710 -325 58940 -95
rect 59060 -325 59290 -95
rect 59410 -325 59640 -95
rect 59760 -325 59990 -95
rect 60110 -325 60340 -95
rect 60460 -180 60690 -95
rect 60810 -180 61040 -95
rect 61160 -180 61390 -95
rect 60460 -230 61390 -180
rect 60460 -325 60690 -230
rect 60810 -325 61040 -230
rect 61160 -325 61390 -230
rect 57970 -510 58020 -505
rect 57970 -550 57975 -510
rect 58015 -550 58020 -510
rect 57970 -555 58020 -550
<< via3 >>
rect 55785 6185 55825 6190
rect 55785 6155 55790 6185
rect 55790 6155 55820 6185
rect 55820 6155 55825 6185
rect 55785 6150 55825 6155
rect 54315 1910 54355 1915
rect 54315 1880 54320 1910
rect 54320 1880 54350 1910
rect 54350 1880 54355 1910
rect 54315 1875 54355 1880
rect 59445 1910 59485 1915
rect 59445 1880 59450 1910
rect 59450 1880 59480 1910
rect 59480 1880 59485 1910
rect 59445 1875 59485 1880
rect 57975 -515 58015 -510
rect 57975 -545 57980 -515
rect 57980 -545 58010 -515
rect 58010 -545 58015 -515
rect 57975 -550 58015 -545
<< mimcap >>
rect 52425 5765 52625 5840
rect 52425 5725 52505 5765
rect 52545 5725 52625 5765
rect 52425 5640 52625 5725
rect 52775 5765 52975 5840
rect 52775 5725 52855 5765
rect 52895 5725 52975 5765
rect 52775 5640 52975 5725
rect 53125 5765 53325 5840
rect 53125 5725 53205 5765
rect 53245 5725 53325 5765
rect 53125 5640 53325 5725
rect 53475 5765 53675 5840
rect 53475 5725 53555 5765
rect 53595 5725 53675 5765
rect 53475 5640 53675 5725
rect 53825 5765 54025 5840
rect 53825 5725 53905 5765
rect 53945 5725 54025 5765
rect 53825 5640 54025 5725
rect 54175 5765 54375 5840
rect 54175 5725 54255 5765
rect 54295 5725 54375 5765
rect 54175 5640 54375 5725
rect 54525 5765 54725 5840
rect 54525 5725 54605 5765
rect 54645 5725 54725 5765
rect 54525 5640 54725 5725
rect 54875 5765 55075 5840
rect 54875 5725 54955 5765
rect 54995 5725 55075 5765
rect 54875 5640 55075 5725
rect 55225 5765 55425 5840
rect 55225 5725 55305 5765
rect 55345 5725 55425 5765
rect 55225 5640 55425 5725
rect 55575 5765 55775 5840
rect 55575 5725 55655 5765
rect 55695 5725 55775 5765
rect 55575 5640 55775 5725
rect 55925 5765 56125 5840
rect 55925 5725 56005 5765
rect 56045 5725 56125 5765
rect 55925 5640 56125 5725
rect 56275 5765 56475 5840
rect 56275 5725 56355 5765
rect 56395 5725 56475 5765
rect 56275 5640 56475 5725
rect 56625 5765 56825 5840
rect 56625 5725 56705 5765
rect 56745 5725 56825 5765
rect 56625 5640 56825 5725
rect 56975 5765 57175 5840
rect 56975 5725 57055 5765
rect 57095 5725 57175 5765
rect 56975 5640 57175 5725
rect 57325 5765 57525 5840
rect 57325 5725 57405 5765
rect 57445 5725 57525 5765
rect 57325 5640 57525 5725
rect 57675 5765 57875 5840
rect 57675 5725 57755 5765
rect 57795 5725 57875 5765
rect 57675 5640 57875 5725
rect 58025 5765 58225 5840
rect 58025 5725 58105 5765
rect 58145 5725 58225 5765
rect 58025 5640 58225 5725
rect 58375 5765 58575 5840
rect 58375 5725 58455 5765
rect 58495 5725 58575 5765
rect 58375 5640 58575 5725
rect 58725 5765 58925 5840
rect 58725 5725 58805 5765
rect 58845 5725 58925 5765
rect 58725 5640 58925 5725
rect 59075 5765 59275 5840
rect 59075 5725 59155 5765
rect 59195 5725 59275 5765
rect 59075 5640 59275 5725
rect 59425 5765 59625 5840
rect 59425 5725 59505 5765
rect 59545 5725 59625 5765
rect 59425 5640 59625 5725
rect 59775 5765 59975 5840
rect 59775 5725 59855 5765
rect 59895 5725 59975 5765
rect 59775 5640 59975 5725
rect 60125 5765 60325 5840
rect 60125 5725 60205 5765
rect 60245 5725 60325 5765
rect 60125 5640 60325 5725
rect 60475 5765 60675 5840
rect 60475 5725 60555 5765
rect 60595 5725 60675 5765
rect 60475 5640 60675 5725
rect 60825 5765 61025 5840
rect 60825 5725 60905 5765
rect 60945 5725 61025 5765
rect 60825 5640 61025 5725
rect 61175 5765 61375 5840
rect 61175 5725 61255 5765
rect 61295 5725 61375 5765
rect 61175 5640 61375 5725
rect 52425 5415 52625 5490
rect 52425 5375 52505 5415
rect 52545 5375 52625 5415
rect 52425 5290 52625 5375
rect 52775 5415 52975 5490
rect 52775 5375 52855 5415
rect 52895 5375 52975 5415
rect 52775 5290 52975 5375
rect 53125 5415 53325 5490
rect 53125 5375 53205 5415
rect 53245 5375 53325 5415
rect 53125 5290 53325 5375
rect 53475 5415 53675 5490
rect 53475 5375 53555 5415
rect 53595 5375 53675 5415
rect 53475 5290 53675 5375
rect 53825 5415 54025 5490
rect 53825 5375 53905 5415
rect 53945 5375 54025 5415
rect 53825 5290 54025 5375
rect 54175 5415 54375 5490
rect 54175 5375 54255 5415
rect 54295 5375 54375 5415
rect 54175 5290 54375 5375
rect 54525 5415 54725 5490
rect 54525 5375 54605 5415
rect 54645 5375 54725 5415
rect 54525 5290 54725 5375
rect 54875 5415 55075 5490
rect 54875 5375 54955 5415
rect 54995 5375 55075 5415
rect 54875 5290 55075 5375
rect 55225 5415 55425 5490
rect 55225 5375 55305 5415
rect 55345 5375 55425 5415
rect 55225 5290 55425 5375
rect 55575 5415 55775 5490
rect 55575 5375 55655 5415
rect 55695 5375 55775 5415
rect 55575 5290 55775 5375
rect 55925 5415 56125 5490
rect 55925 5375 56005 5415
rect 56045 5375 56125 5415
rect 55925 5290 56125 5375
rect 56275 5415 56475 5490
rect 56275 5375 56355 5415
rect 56395 5375 56475 5415
rect 56275 5290 56475 5375
rect 56625 5415 56825 5490
rect 56625 5375 56705 5415
rect 56745 5375 56825 5415
rect 56625 5290 56825 5375
rect 56975 5415 57175 5490
rect 56975 5375 57055 5415
rect 57095 5375 57175 5415
rect 56975 5290 57175 5375
rect 57325 5415 57525 5490
rect 57325 5375 57405 5415
rect 57445 5375 57525 5415
rect 57325 5290 57525 5375
rect 57675 5415 57875 5490
rect 57675 5375 57755 5415
rect 57795 5375 57875 5415
rect 57675 5290 57875 5375
rect 58025 5415 58225 5490
rect 58025 5375 58105 5415
rect 58145 5375 58225 5415
rect 58025 5290 58225 5375
rect 58375 5415 58575 5490
rect 58375 5375 58455 5415
rect 58495 5375 58575 5415
rect 58375 5290 58575 5375
rect 58725 5415 58925 5490
rect 58725 5375 58805 5415
rect 58845 5375 58925 5415
rect 58725 5290 58925 5375
rect 59075 5415 59275 5490
rect 59075 5375 59155 5415
rect 59195 5375 59275 5415
rect 59075 5290 59275 5375
rect 59425 5415 59625 5490
rect 59425 5375 59505 5415
rect 59545 5375 59625 5415
rect 59425 5290 59625 5375
rect 59775 5415 59975 5490
rect 59775 5375 59855 5415
rect 59895 5375 59975 5415
rect 59775 5290 59975 5375
rect 60125 5415 60325 5490
rect 60125 5375 60205 5415
rect 60245 5375 60325 5415
rect 60125 5290 60325 5375
rect 60475 5415 60675 5490
rect 60475 5375 60555 5415
rect 60595 5375 60675 5415
rect 60475 5290 60675 5375
rect 60825 5415 61025 5490
rect 60825 5375 60905 5415
rect 60945 5375 61025 5415
rect 60825 5290 61025 5375
rect 61175 5415 61375 5490
rect 61175 5375 61255 5415
rect 61295 5375 61375 5415
rect 61175 5290 61375 5375
rect 52425 5065 52625 5140
rect 52425 5025 52505 5065
rect 52545 5025 52625 5065
rect 52425 4940 52625 5025
rect 52775 5065 52975 5140
rect 52775 5025 52855 5065
rect 52895 5025 52975 5065
rect 52775 4940 52975 5025
rect 53125 5065 53325 5140
rect 53125 5025 53205 5065
rect 53245 5025 53325 5065
rect 53125 4940 53325 5025
rect 53475 5065 53675 5140
rect 53475 5025 53555 5065
rect 53595 5025 53675 5065
rect 53475 4940 53675 5025
rect 53825 5065 54025 5140
rect 53825 5025 53905 5065
rect 53945 5025 54025 5065
rect 53825 4940 54025 5025
rect 54175 5065 54375 5140
rect 54175 5025 54255 5065
rect 54295 5025 54375 5065
rect 54175 4940 54375 5025
rect 54525 5065 54725 5140
rect 54525 5025 54605 5065
rect 54645 5025 54725 5065
rect 54525 4940 54725 5025
rect 54875 5065 55075 5140
rect 54875 5025 54955 5065
rect 54995 5025 55075 5065
rect 54875 4940 55075 5025
rect 55225 5065 55425 5140
rect 55225 5025 55305 5065
rect 55345 5025 55425 5065
rect 55225 4940 55425 5025
rect 55575 5055 55775 5140
rect 55575 5015 55655 5055
rect 55695 5015 55775 5055
rect 55575 4940 55775 5015
rect 55925 5055 56125 5140
rect 55925 5015 56005 5055
rect 56045 5015 56125 5055
rect 55925 4940 56125 5015
rect 56275 5055 56475 5140
rect 56275 5015 56355 5055
rect 56395 5015 56475 5055
rect 56275 4940 56475 5015
rect 56625 5055 56825 5140
rect 56625 5015 56705 5055
rect 56745 5015 56825 5055
rect 56625 4940 56825 5015
rect 56975 5055 57175 5140
rect 56975 5015 57055 5055
rect 57095 5015 57175 5055
rect 56975 4940 57175 5015
rect 57325 5055 57525 5140
rect 57325 5015 57405 5055
rect 57445 5015 57525 5055
rect 57325 4940 57525 5015
rect 57675 5055 57875 5140
rect 57675 5015 57755 5055
rect 57795 5015 57875 5055
rect 57675 4940 57875 5015
rect 58025 5055 58225 5140
rect 58025 5015 58105 5055
rect 58145 5015 58225 5055
rect 58025 4940 58225 5015
rect 58375 5065 58575 5140
rect 58375 5025 58455 5065
rect 58495 5025 58575 5065
rect 58375 4940 58575 5025
rect 58725 5065 58925 5140
rect 58725 5025 58805 5065
rect 58845 5025 58925 5065
rect 58725 4940 58925 5025
rect 59075 5065 59275 5140
rect 59075 5025 59155 5065
rect 59195 5025 59275 5065
rect 59075 4940 59275 5025
rect 59425 5065 59625 5140
rect 59425 5025 59505 5065
rect 59545 5025 59625 5065
rect 59425 4940 59625 5025
rect 59775 5065 59975 5140
rect 59775 5025 59855 5065
rect 59895 5025 59975 5065
rect 59775 4940 59975 5025
rect 60125 5065 60325 5140
rect 60125 5025 60205 5065
rect 60245 5025 60325 5065
rect 60125 4940 60325 5025
rect 60475 5065 60675 5140
rect 60475 5025 60555 5065
rect 60595 5025 60675 5065
rect 60475 4940 60675 5025
rect 60825 5065 61025 5140
rect 60825 5025 60905 5065
rect 60945 5025 61025 5065
rect 60825 4940 61025 5025
rect 61175 5065 61375 5140
rect 61175 5025 61255 5065
rect 61295 5025 61375 5065
rect 61175 4940 61375 5025
rect 52425 4715 52625 4790
rect 52425 4675 52505 4715
rect 52545 4675 52625 4715
rect 52425 4590 52625 4675
rect 52775 4715 52975 4790
rect 52775 4675 52855 4715
rect 52895 4675 52975 4715
rect 52775 4590 52975 4675
rect 53125 4715 53325 4790
rect 53125 4675 53205 4715
rect 53245 4675 53325 4715
rect 53125 4590 53325 4675
rect 53475 4715 53675 4790
rect 53475 4675 53555 4715
rect 53595 4675 53675 4715
rect 53475 4590 53675 4675
rect 53825 4715 54025 4790
rect 53825 4675 53905 4715
rect 53945 4675 54025 4715
rect 53825 4590 54025 4675
rect 54175 4715 54375 4790
rect 54175 4675 54255 4715
rect 54295 4675 54375 4715
rect 54175 4590 54375 4675
rect 54525 4715 54725 4790
rect 54525 4675 54605 4715
rect 54645 4675 54725 4715
rect 54525 4590 54725 4675
rect 54875 4715 55075 4790
rect 54875 4675 54955 4715
rect 54995 4675 55075 4715
rect 54875 4590 55075 4675
rect 55225 4715 55425 4790
rect 55225 4675 55305 4715
rect 55345 4675 55425 4715
rect 55225 4590 55425 4675
rect 58375 4715 58575 4790
rect 58375 4675 58455 4715
rect 58495 4675 58575 4715
rect 58375 4590 58575 4675
rect 58725 4715 58925 4790
rect 58725 4675 58805 4715
rect 58845 4675 58925 4715
rect 58725 4590 58925 4675
rect 59075 4715 59275 4790
rect 59075 4675 59155 4715
rect 59195 4675 59275 4715
rect 59075 4590 59275 4675
rect 59425 4715 59625 4790
rect 59425 4675 59505 4715
rect 59545 4675 59625 4715
rect 59425 4590 59625 4675
rect 59775 4715 59975 4790
rect 59775 4675 59855 4715
rect 59895 4675 59975 4715
rect 59775 4590 59975 4675
rect 60125 4715 60325 4790
rect 60125 4675 60205 4715
rect 60245 4675 60325 4715
rect 60125 4590 60325 4675
rect 60475 4715 60675 4790
rect 60475 4675 60555 4715
rect 60595 4675 60675 4715
rect 60475 4590 60675 4675
rect 60825 4715 61025 4790
rect 60825 4675 60905 4715
rect 60945 4675 61025 4715
rect 60825 4590 61025 4675
rect 61175 4715 61375 4790
rect 61175 4675 61255 4715
rect 61295 4675 61375 4715
rect 61175 4590 61375 4675
rect 52425 4365 52625 4440
rect 52425 4325 52505 4365
rect 52545 4325 52625 4365
rect 52425 4240 52625 4325
rect 52775 4365 52975 4440
rect 52775 4325 52855 4365
rect 52895 4325 52975 4365
rect 52775 4240 52975 4325
rect 53125 4365 53325 4440
rect 53125 4325 53205 4365
rect 53245 4325 53325 4365
rect 53125 4240 53325 4325
rect 53475 4365 53675 4440
rect 53475 4325 53555 4365
rect 53595 4325 53675 4365
rect 53475 4240 53675 4325
rect 53825 4365 54025 4440
rect 53825 4325 53905 4365
rect 53945 4325 54025 4365
rect 53825 4240 54025 4325
rect 54175 4365 54375 4440
rect 54175 4325 54255 4365
rect 54295 4325 54375 4365
rect 54175 4240 54375 4325
rect 54525 4365 54725 4440
rect 54525 4325 54605 4365
rect 54645 4325 54725 4365
rect 54525 4240 54725 4325
rect 54875 4365 55075 4440
rect 54875 4325 54955 4365
rect 54995 4325 55075 4365
rect 54875 4240 55075 4325
rect 55225 4365 55425 4440
rect 55225 4325 55305 4365
rect 55345 4325 55425 4365
rect 55225 4240 55425 4325
rect 58375 4365 58575 4440
rect 58375 4325 58455 4365
rect 58495 4325 58575 4365
rect 58375 4240 58575 4325
rect 58725 4365 58925 4440
rect 58725 4325 58805 4365
rect 58845 4325 58925 4365
rect 58725 4240 58925 4325
rect 59075 4365 59275 4440
rect 59075 4325 59155 4365
rect 59195 4325 59275 4365
rect 59075 4240 59275 4325
rect 59425 4365 59625 4440
rect 59425 4325 59505 4365
rect 59545 4325 59625 4365
rect 59425 4240 59625 4325
rect 59775 4365 59975 4440
rect 59775 4325 59855 4365
rect 59895 4325 59975 4365
rect 59775 4240 59975 4325
rect 60125 4365 60325 4440
rect 60125 4325 60205 4365
rect 60245 4325 60325 4365
rect 60125 4240 60325 4325
rect 60475 4365 60675 4440
rect 60475 4325 60555 4365
rect 60595 4325 60675 4365
rect 60475 4240 60675 4325
rect 60825 4365 61025 4440
rect 60825 4325 60905 4365
rect 60945 4325 61025 4365
rect 60825 4240 61025 4325
rect 61175 4365 61375 4440
rect 61175 4325 61255 4365
rect 61295 4325 61375 4365
rect 61175 4240 61375 4325
rect 52425 4015 52625 4090
rect 52425 3975 52505 4015
rect 52545 3975 52625 4015
rect 52425 3890 52625 3975
rect 52775 4015 52975 4090
rect 52775 3975 52855 4015
rect 52895 3975 52975 4015
rect 52775 3890 52975 3975
rect 53125 4015 53325 4090
rect 53125 3975 53205 4015
rect 53245 3975 53325 4015
rect 53125 3890 53325 3975
rect 53475 4015 53675 4090
rect 53475 3975 53555 4015
rect 53595 3975 53675 4015
rect 53475 3890 53675 3975
rect 53825 4015 54025 4090
rect 53825 3975 53905 4015
rect 53945 3975 54025 4015
rect 53825 3890 54025 3975
rect 59775 4015 59975 4090
rect 59775 3975 59855 4015
rect 59895 3975 59975 4015
rect 59775 3890 59975 3975
rect 60125 4015 60325 4090
rect 60125 3975 60205 4015
rect 60245 3975 60325 4015
rect 60125 3890 60325 3975
rect 60475 4015 60675 4090
rect 60475 3975 60555 4015
rect 60595 3975 60675 4015
rect 60475 3890 60675 3975
rect 60825 4015 61025 4090
rect 60825 3975 60905 4015
rect 60945 3975 61025 4015
rect 60825 3890 61025 3975
rect 61175 4015 61375 4090
rect 61175 3975 61255 4015
rect 61295 3975 61375 4015
rect 61175 3890 61375 3975
rect 52425 3665 52625 3740
rect 52425 3625 52505 3665
rect 52545 3625 52625 3665
rect 52425 3540 52625 3625
rect 52775 3665 52975 3740
rect 52775 3625 52855 3665
rect 52895 3625 52975 3665
rect 52775 3540 52975 3625
rect 53125 3665 53325 3740
rect 53125 3625 53205 3665
rect 53245 3625 53325 3665
rect 53125 3540 53325 3625
rect 53475 3665 53675 3740
rect 53475 3625 53555 3665
rect 53595 3625 53675 3665
rect 53475 3540 53675 3625
rect 53825 3665 54025 3740
rect 53825 3625 53905 3665
rect 53945 3625 54025 3665
rect 53825 3540 54025 3625
rect 59775 3665 59975 3740
rect 59775 3625 59855 3665
rect 59895 3625 59975 3665
rect 59775 3540 59975 3625
rect 60125 3665 60325 3740
rect 60125 3625 60205 3665
rect 60245 3625 60325 3665
rect 60125 3540 60325 3625
rect 60475 3665 60675 3740
rect 60475 3625 60555 3665
rect 60595 3625 60675 3665
rect 60475 3540 60675 3625
rect 60825 3665 61025 3740
rect 60825 3625 60905 3665
rect 60945 3625 61025 3665
rect 60825 3540 61025 3625
rect 61175 3665 61375 3740
rect 61175 3625 61255 3665
rect 61295 3625 61375 3665
rect 61175 3540 61375 3625
rect 52425 3315 52625 3390
rect 52425 3275 52505 3315
rect 52545 3275 52625 3315
rect 52425 3190 52625 3275
rect 52775 3315 52975 3390
rect 52775 3275 52855 3315
rect 52895 3275 52975 3315
rect 52775 3190 52975 3275
rect 53125 3315 53325 3390
rect 53125 3275 53205 3315
rect 53245 3275 53325 3315
rect 53125 3190 53325 3275
rect 53475 3315 53675 3390
rect 53475 3275 53555 3315
rect 53595 3275 53675 3315
rect 53475 3190 53675 3275
rect 53825 3315 54025 3390
rect 53825 3275 53905 3315
rect 53945 3275 54025 3315
rect 53825 3190 54025 3275
rect 59775 3315 59975 3390
rect 59775 3275 59855 3315
rect 59895 3275 59975 3315
rect 59775 3190 59975 3275
rect 60125 3315 60325 3390
rect 60125 3275 60205 3315
rect 60245 3275 60325 3315
rect 60125 3190 60325 3275
rect 60475 3315 60675 3390
rect 60475 3275 60555 3315
rect 60595 3275 60675 3315
rect 60475 3190 60675 3275
rect 60825 3315 61025 3390
rect 60825 3275 60905 3315
rect 60945 3275 61025 3315
rect 60825 3190 61025 3275
rect 61175 3315 61375 3390
rect 61175 3275 61255 3315
rect 61295 3275 61375 3315
rect 61175 3190 61375 3275
rect 52425 2965 52625 3040
rect 52425 2925 52505 2965
rect 52545 2925 52625 2965
rect 52425 2840 52625 2925
rect 52775 2965 52975 3040
rect 52775 2925 52855 2965
rect 52895 2925 52975 2965
rect 52775 2840 52975 2925
rect 53125 2965 53325 3040
rect 53125 2925 53205 2965
rect 53245 2925 53325 2965
rect 53125 2840 53325 2925
rect 53475 2965 53675 3040
rect 53475 2925 53555 2965
rect 53595 2925 53675 2965
rect 53475 2840 53675 2925
rect 53825 2965 54025 3040
rect 53825 2925 53905 2965
rect 53945 2925 54025 2965
rect 53825 2840 54025 2925
rect 59775 2965 59975 3040
rect 59775 2925 59855 2965
rect 59895 2925 59975 2965
rect 59775 2840 59975 2925
rect 60125 2965 60325 3040
rect 60125 2925 60205 2965
rect 60245 2925 60325 2965
rect 60125 2840 60325 2925
rect 60475 2965 60675 3040
rect 60475 2925 60555 2965
rect 60595 2925 60675 2965
rect 60475 2840 60675 2925
rect 60825 2965 61025 3040
rect 60825 2925 60905 2965
rect 60945 2925 61025 2965
rect 60825 2840 61025 2925
rect 61175 2965 61375 3040
rect 61175 2925 61255 2965
rect 61295 2925 61375 2965
rect 61175 2840 61375 2925
rect 52425 2615 52625 2690
rect 52425 2575 52505 2615
rect 52545 2575 52625 2615
rect 52425 2490 52625 2575
rect 52775 2615 52975 2690
rect 52775 2575 52855 2615
rect 52895 2575 52975 2615
rect 52775 2490 52975 2575
rect 53125 2615 53325 2690
rect 53125 2575 53205 2615
rect 53245 2575 53325 2615
rect 53125 2490 53325 2575
rect 53475 2615 53675 2690
rect 53475 2575 53555 2615
rect 53595 2575 53675 2615
rect 53475 2490 53675 2575
rect 53825 2615 54025 2690
rect 53825 2575 53905 2615
rect 53945 2575 54025 2615
rect 53825 2490 54025 2575
rect 59775 2615 59975 2690
rect 59775 2575 59855 2615
rect 59895 2575 59975 2615
rect 59775 2490 59975 2575
rect 60125 2615 60325 2690
rect 60125 2575 60205 2615
rect 60245 2575 60325 2615
rect 60125 2490 60325 2575
rect 60475 2615 60675 2690
rect 60475 2575 60555 2615
rect 60595 2575 60675 2615
rect 60475 2490 60675 2575
rect 60825 2615 61025 2690
rect 60825 2575 60905 2615
rect 60945 2575 61025 2615
rect 60825 2490 61025 2575
rect 61175 2615 61375 2690
rect 61175 2575 61255 2615
rect 61295 2575 61375 2615
rect 61175 2490 61375 2575
rect 52425 2265 52625 2340
rect 52425 2225 52505 2265
rect 52545 2225 52625 2265
rect 52425 2140 52625 2225
rect 52775 2265 52975 2340
rect 52775 2225 52855 2265
rect 52895 2225 52975 2265
rect 52775 2140 52975 2225
rect 53125 2265 53325 2340
rect 53125 2225 53205 2265
rect 53245 2225 53325 2265
rect 53125 2140 53325 2225
rect 53475 2265 53675 2340
rect 53475 2225 53555 2265
rect 53595 2225 53675 2265
rect 53475 2140 53675 2225
rect 53825 2265 54025 2340
rect 53825 2225 53905 2265
rect 53945 2225 54025 2265
rect 53825 2140 54025 2225
rect 59775 2265 59975 2340
rect 59775 2225 59855 2265
rect 59895 2225 59975 2265
rect 59775 2140 59975 2225
rect 60125 2265 60325 2340
rect 60125 2225 60205 2265
rect 60245 2225 60325 2265
rect 60125 2140 60325 2225
rect 60475 2265 60675 2340
rect 60475 2225 60555 2265
rect 60595 2225 60675 2265
rect 60475 2140 60675 2225
rect 60825 2265 61025 2340
rect 60825 2225 60905 2265
rect 60945 2225 61025 2265
rect 60825 2140 61025 2225
rect 61175 2265 61375 2340
rect 61175 2225 61255 2265
rect 61295 2225 61375 2265
rect 61175 2140 61375 2225
rect 52425 1915 52625 1990
rect 52425 1875 52505 1915
rect 52545 1875 52625 1915
rect 52425 1790 52625 1875
rect 52775 1915 52975 1990
rect 52775 1875 52855 1915
rect 52895 1875 52975 1915
rect 52775 1790 52975 1875
rect 53125 1915 53325 1990
rect 53125 1875 53205 1915
rect 53245 1875 53325 1915
rect 53125 1790 53325 1875
rect 53475 1915 53675 1990
rect 53475 1875 53555 1915
rect 53595 1875 53675 1915
rect 53475 1790 53675 1875
rect 53825 1915 54025 1990
rect 53825 1875 53905 1915
rect 53945 1875 54025 1915
rect 53825 1790 54025 1875
rect 59775 1915 59975 1990
rect 59775 1875 59855 1915
rect 59895 1875 59975 1915
rect 59775 1790 59975 1875
rect 60125 1915 60325 1990
rect 60125 1875 60205 1915
rect 60245 1875 60325 1915
rect 60125 1790 60325 1875
rect 60475 1915 60675 1990
rect 60475 1875 60555 1915
rect 60595 1875 60675 1915
rect 60475 1790 60675 1875
rect 60825 1915 61025 1990
rect 60825 1875 60905 1915
rect 60945 1875 61025 1915
rect 60825 1790 61025 1875
rect 61175 1915 61375 1990
rect 61175 1875 61255 1915
rect 61295 1875 61375 1915
rect 61175 1790 61375 1875
rect 52425 1565 52625 1640
rect 52425 1525 52505 1565
rect 52545 1525 52625 1565
rect 52425 1440 52625 1525
rect 52775 1565 52975 1640
rect 52775 1525 52855 1565
rect 52895 1525 52975 1565
rect 52775 1440 52975 1525
rect 53125 1565 53325 1640
rect 53125 1525 53205 1565
rect 53245 1525 53325 1565
rect 53125 1440 53325 1525
rect 53475 1565 53675 1640
rect 53475 1525 53555 1565
rect 53595 1525 53675 1565
rect 53475 1440 53675 1525
rect 53825 1565 54025 1640
rect 53825 1525 53905 1565
rect 53945 1525 54025 1565
rect 53825 1440 54025 1525
rect 59775 1565 59975 1640
rect 59775 1525 59855 1565
rect 59895 1525 59975 1565
rect 59775 1440 59975 1525
rect 60125 1565 60325 1640
rect 60125 1525 60205 1565
rect 60245 1525 60325 1565
rect 60125 1440 60325 1525
rect 60475 1565 60675 1640
rect 60475 1525 60555 1565
rect 60595 1525 60675 1565
rect 60475 1440 60675 1525
rect 60825 1565 61025 1640
rect 60825 1525 60905 1565
rect 60945 1525 61025 1565
rect 60825 1440 61025 1525
rect 61175 1565 61375 1640
rect 61175 1525 61255 1565
rect 61295 1525 61375 1565
rect 61175 1440 61375 1525
rect 52425 1215 52625 1290
rect 52425 1175 52505 1215
rect 52545 1175 52625 1215
rect 52425 1090 52625 1175
rect 52775 1215 52975 1290
rect 52775 1175 52855 1215
rect 52895 1175 52975 1215
rect 52775 1090 52975 1175
rect 53125 1215 53325 1290
rect 53125 1175 53205 1215
rect 53245 1175 53325 1215
rect 53125 1090 53325 1175
rect 53475 1215 53675 1290
rect 53475 1175 53555 1215
rect 53595 1175 53675 1215
rect 53475 1090 53675 1175
rect 53825 1215 54025 1290
rect 53825 1175 53905 1215
rect 53945 1175 54025 1215
rect 53825 1090 54025 1175
rect 59775 1215 59975 1290
rect 59775 1175 59855 1215
rect 59895 1175 59975 1215
rect 59775 1090 59975 1175
rect 60125 1215 60325 1290
rect 60125 1175 60205 1215
rect 60245 1175 60325 1215
rect 60125 1090 60325 1175
rect 60475 1215 60675 1290
rect 60475 1175 60555 1215
rect 60595 1175 60675 1215
rect 60475 1090 60675 1175
rect 60825 1215 61025 1290
rect 60825 1175 60905 1215
rect 60945 1175 61025 1215
rect 60825 1090 61025 1175
rect 61175 1215 61375 1290
rect 61175 1175 61255 1215
rect 61295 1175 61375 1215
rect 61175 1090 61375 1175
rect 52425 865 52625 940
rect 52425 825 52505 865
rect 52545 825 52625 865
rect 52425 740 52625 825
rect 52775 865 52975 940
rect 52775 825 52855 865
rect 52895 825 52975 865
rect 52775 740 52975 825
rect 53125 865 53325 940
rect 53125 825 53205 865
rect 53245 825 53325 865
rect 53125 740 53325 825
rect 53475 865 53675 940
rect 53475 825 53555 865
rect 53595 825 53675 865
rect 53475 740 53675 825
rect 53825 865 54025 940
rect 53825 825 53905 865
rect 53945 825 54025 865
rect 53825 740 54025 825
rect 59775 865 59975 940
rect 59775 825 59855 865
rect 59895 825 59975 865
rect 59775 740 59975 825
rect 60125 865 60325 940
rect 60125 825 60205 865
rect 60245 825 60325 865
rect 60125 740 60325 825
rect 60475 865 60675 940
rect 60475 825 60555 865
rect 60595 825 60675 865
rect 60475 740 60675 825
rect 60825 865 61025 940
rect 60825 825 60905 865
rect 60945 825 61025 865
rect 60825 740 61025 825
rect 61175 865 61375 940
rect 61175 825 61255 865
rect 61295 825 61375 865
rect 61175 740 61375 825
rect 52425 515 52625 590
rect 52425 475 52505 515
rect 52545 475 52625 515
rect 52425 390 52625 475
rect 52775 515 52975 590
rect 52775 475 52855 515
rect 52895 475 52975 515
rect 52775 390 52975 475
rect 53125 515 53325 590
rect 53125 475 53205 515
rect 53245 475 53325 515
rect 53125 390 53325 475
rect 53475 515 53675 590
rect 53475 475 53555 515
rect 53595 475 53675 515
rect 53475 390 53675 475
rect 53825 515 54025 590
rect 53825 475 53905 515
rect 53945 475 54025 515
rect 53825 390 54025 475
rect 59775 515 59975 590
rect 59775 475 59855 515
rect 59895 475 59975 515
rect 59775 390 59975 475
rect 60125 515 60325 590
rect 60125 475 60205 515
rect 60245 475 60325 515
rect 60125 390 60325 475
rect 60475 515 60675 590
rect 60475 475 60555 515
rect 60595 475 60675 515
rect 60475 390 60675 475
rect 60825 515 61025 590
rect 60825 475 60905 515
rect 60945 475 61025 515
rect 60825 390 61025 475
rect 61175 515 61375 590
rect 61175 475 61255 515
rect 61295 475 61375 515
rect 61175 390 61375 475
rect 52425 165 52625 240
rect 52425 125 52505 165
rect 52545 125 52625 165
rect 52425 40 52625 125
rect 52775 165 52975 240
rect 52775 125 52855 165
rect 52895 125 52975 165
rect 52775 40 52975 125
rect 53125 165 53325 240
rect 53125 125 53205 165
rect 53245 125 53325 165
rect 53125 40 53325 125
rect 53475 165 53675 240
rect 53475 125 53555 165
rect 53595 125 53675 165
rect 53475 40 53675 125
rect 53825 165 54025 240
rect 53825 125 53905 165
rect 53945 125 54025 165
rect 53825 40 54025 125
rect 54175 165 54375 240
rect 54175 125 54255 165
rect 54295 125 54375 165
rect 54175 40 54375 125
rect 54525 165 54725 240
rect 54525 125 54605 165
rect 54645 125 54725 165
rect 54525 40 54725 125
rect 54875 165 55075 240
rect 54875 125 54955 165
rect 54995 125 55075 165
rect 54875 40 55075 125
rect 55225 165 55425 240
rect 55225 125 55305 165
rect 55345 125 55425 165
rect 55225 40 55425 125
rect 55575 165 55775 240
rect 55575 125 55655 165
rect 55695 125 55775 165
rect 55575 40 55775 125
rect 55925 165 56125 240
rect 55925 125 56005 165
rect 56045 125 56125 165
rect 55925 40 56125 125
rect 56275 165 56475 240
rect 56275 125 56355 165
rect 56395 125 56475 165
rect 56275 40 56475 125
rect 56625 165 56825 240
rect 56625 125 56705 165
rect 56745 125 56825 165
rect 56625 40 56825 125
rect 56975 165 57175 240
rect 56975 125 57055 165
rect 57095 125 57175 165
rect 56975 40 57175 125
rect 57325 165 57525 240
rect 57325 125 57405 165
rect 57445 125 57525 165
rect 57325 40 57525 125
rect 57675 165 57875 240
rect 57675 125 57755 165
rect 57795 125 57875 165
rect 57675 40 57875 125
rect 58025 165 58225 240
rect 58025 125 58105 165
rect 58145 125 58225 165
rect 58025 40 58225 125
rect 58375 165 58575 240
rect 58375 125 58455 165
rect 58495 125 58575 165
rect 58375 40 58575 125
rect 58725 165 58925 240
rect 58725 125 58805 165
rect 58845 125 58925 165
rect 58725 40 58925 125
rect 59075 165 59275 240
rect 59075 125 59155 165
rect 59195 125 59275 165
rect 59075 40 59275 125
rect 59425 165 59625 240
rect 59425 125 59505 165
rect 59545 125 59625 165
rect 59425 40 59625 125
rect 59775 165 59975 240
rect 59775 125 59855 165
rect 59895 125 59975 165
rect 59775 40 59975 125
rect 60125 165 60325 240
rect 60125 125 60205 165
rect 60245 125 60325 165
rect 60125 40 60325 125
rect 60475 165 60675 240
rect 60475 125 60555 165
rect 60595 125 60675 165
rect 60475 40 60675 125
rect 60825 165 61025 240
rect 60825 125 60905 165
rect 60945 125 61025 165
rect 60825 40 61025 125
rect 61175 165 61375 240
rect 61175 125 61255 165
rect 61295 125 61375 165
rect 61175 40 61375 125
rect 52425 -185 52625 -110
rect 52425 -225 52505 -185
rect 52545 -225 52625 -185
rect 52425 -310 52625 -225
rect 52775 -185 52975 -110
rect 52775 -225 52855 -185
rect 52895 -225 52975 -185
rect 52775 -310 52975 -225
rect 53125 -185 53325 -110
rect 53125 -225 53205 -185
rect 53245 -225 53325 -185
rect 53125 -310 53325 -225
rect 53475 -185 53675 -110
rect 53475 -225 53555 -185
rect 53595 -225 53675 -185
rect 53475 -310 53675 -225
rect 53825 -185 54025 -110
rect 53825 -225 53905 -185
rect 53945 -225 54025 -185
rect 53825 -310 54025 -225
rect 54175 -185 54375 -110
rect 54175 -225 54255 -185
rect 54295 -225 54375 -185
rect 54175 -310 54375 -225
rect 54525 -185 54725 -110
rect 54525 -225 54605 -185
rect 54645 -225 54725 -185
rect 54525 -310 54725 -225
rect 54875 -185 55075 -110
rect 54875 -225 54955 -185
rect 54995 -225 55075 -185
rect 54875 -310 55075 -225
rect 55225 -185 55425 -110
rect 55225 -225 55305 -185
rect 55345 -225 55425 -185
rect 55225 -310 55425 -225
rect 55575 -185 55775 -110
rect 55575 -225 55655 -185
rect 55695 -225 55775 -185
rect 55575 -310 55775 -225
rect 55925 -185 56125 -110
rect 55925 -225 56005 -185
rect 56045 -225 56125 -185
rect 55925 -310 56125 -225
rect 56275 -185 56475 -110
rect 56275 -225 56355 -185
rect 56395 -225 56475 -185
rect 56275 -310 56475 -225
rect 56625 -185 56825 -110
rect 56625 -225 56705 -185
rect 56745 -225 56825 -185
rect 56625 -310 56825 -225
rect 56975 -185 57175 -110
rect 56975 -225 57055 -185
rect 57095 -225 57175 -185
rect 56975 -310 57175 -225
rect 57325 -185 57525 -110
rect 57325 -225 57405 -185
rect 57445 -225 57525 -185
rect 57325 -310 57525 -225
rect 57675 -185 57875 -110
rect 57675 -225 57755 -185
rect 57795 -225 57875 -185
rect 57675 -310 57875 -225
rect 58025 -185 58225 -110
rect 58025 -225 58105 -185
rect 58145 -225 58225 -185
rect 58025 -310 58225 -225
rect 58375 -185 58575 -110
rect 58375 -225 58455 -185
rect 58495 -225 58575 -185
rect 58375 -310 58575 -225
rect 58725 -185 58925 -110
rect 58725 -225 58805 -185
rect 58845 -225 58925 -185
rect 58725 -310 58925 -225
rect 59075 -185 59275 -110
rect 59075 -225 59155 -185
rect 59195 -225 59275 -185
rect 59075 -310 59275 -225
rect 59425 -185 59625 -110
rect 59425 -225 59505 -185
rect 59545 -225 59625 -185
rect 59425 -310 59625 -225
rect 59775 -185 59975 -110
rect 59775 -225 59855 -185
rect 59895 -225 59975 -185
rect 59775 -310 59975 -225
rect 60125 -185 60325 -110
rect 60125 -225 60205 -185
rect 60245 -225 60325 -185
rect 60125 -310 60325 -225
rect 60475 -185 60675 -110
rect 60475 -225 60555 -185
rect 60595 -225 60675 -185
rect 60475 -310 60675 -225
rect 60825 -185 61025 -110
rect 60825 -225 60905 -185
rect 60945 -225 61025 -185
rect 60825 -310 61025 -225
rect 61175 -185 61375 -110
rect 61175 -225 61255 -185
rect 61295 -225 61375 -185
rect 61175 -310 61375 -225
<< mimcapcontact >>
rect 52505 5725 52545 5765
rect 52855 5725 52895 5765
rect 53205 5725 53245 5765
rect 53555 5725 53595 5765
rect 53905 5725 53945 5765
rect 54255 5725 54295 5765
rect 54605 5725 54645 5765
rect 54955 5725 54995 5765
rect 55305 5725 55345 5765
rect 55655 5725 55695 5765
rect 56005 5725 56045 5765
rect 56355 5725 56395 5765
rect 56705 5725 56745 5765
rect 57055 5725 57095 5765
rect 57405 5725 57445 5765
rect 57755 5725 57795 5765
rect 58105 5725 58145 5765
rect 58455 5725 58495 5765
rect 58805 5725 58845 5765
rect 59155 5725 59195 5765
rect 59505 5725 59545 5765
rect 59855 5725 59895 5765
rect 60205 5725 60245 5765
rect 60555 5725 60595 5765
rect 60905 5725 60945 5765
rect 61255 5725 61295 5765
rect 52505 5375 52545 5415
rect 52855 5375 52895 5415
rect 53205 5375 53245 5415
rect 53555 5375 53595 5415
rect 53905 5375 53945 5415
rect 54255 5375 54295 5415
rect 54605 5375 54645 5415
rect 54955 5375 54995 5415
rect 55305 5375 55345 5415
rect 55655 5375 55695 5415
rect 56005 5375 56045 5415
rect 56355 5375 56395 5415
rect 56705 5375 56745 5415
rect 57055 5375 57095 5415
rect 57405 5375 57445 5415
rect 57755 5375 57795 5415
rect 58105 5375 58145 5415
rect 58455 5375 58495 5415
rect 58805 5375 58845 5415
rect 59155 5375 59195 5415
rect 59505 5375 59545 5415
rect 59855 5375 59895 5415
rect 60205 5375 60245 5415
rect 60555 5375 60595 5415
rect 60905 5375 60945 5415
rect 61255 5375 61295 5415
rect 52505 5025 52545 5065
rect 52855 5025 52895 5065
rect 53205 5025 53245 5065
rect 53555 5025 53595 5065
rect 53905 5025 53945 5065
rect 54255 5025 54295 5065
rect 54605 5025 54645 5065
rect 54955 5025 54995 5065
rect 55305 5025 55345 5065
rect 55655 5015 55695 5055
rect 56005 5015 56045 5055
rect 56355 5015 56395 5055
rect 56705 5015 56745 5055
rect 57055 5015 57095 5055
rect 57405 5015 57445 5055
rect 57755 5015 57795 5055
rect 58105 5015 58145 5055
rect 58455 5025 58495 5065
rect 58805 5025 58845 5065
rect 59155 5025 59195 5065
rect 59505 5025 59545 5065
rect 59855 5025 59895 5065
rect 60205 5025 60245 5065
rect 60555 5025 60595 5065
rect 60905 5025 60945 5065
rect 61255 5025 61295 5065
rect 52505 4675 52545 4715
rect 52855 4675 52895 4715
rect 53205 4675 53245 4715
rect 53555 4675 53595 4715
rect 53905 4675 53945 4715
rect 54255 4675 54295 4715
rect 54605 4675 54645 4715
rect 54955 4675 54995 4715
rect 55305 4675 55345 4715
rect 58455 4675 58495 4715
rect 58805 4675 58845 4715
rect 59155 4675 59195 4715
rect 59505 4675 59545 4715
rect 59855 4675 59895 4715
rect 60205 4675 60245 4715
rect 60555 4675 60595 4715
rect 60905 4675 60945 4715
rect 61255 4675 61295 4715
rect 52505 4325 52545 4365
rect 52855 4325 52895 4365
rect 53205 4325 53245 4365
rect 53555 4325 53595 4365
rect 53905 4325 53945 4365
rect 54255 4325 54295 4365
rect 54605 4325 54645 4365
rect 54955 4325 54995 4365
rect 55305 4325 55345 4365
rect 58455 4325 58495 4365
rect 58805 4325 58845 4365
rect 59155 4325 59195 4365
rect 59505 4325 59545 4365
rect 59855 4325 59895 4365
rect 60205 4325 60245 4365
rect 60555 4325 60595 4365
rect 60905 4325 60945 4365
rect 61255 4325 61295 4365
rect 52505 3975 52545 4015
rect 52855 3975 52895 4015
rect 53205 3975 53245 4015
rect 53555 3975 53595 4015
rect 53905 3975 53945 4015
rect 59855 3975 59895 4015
rect 60205 3975 60245 4015
rect 60555 3975 60595 4015
rect 60905 3975 60945 4015
rect 61255 3975 61295 4015
rect 52505 3625 52545 3665
rect 52855 3625 52895 3665
rect 53205 3625 53245 3665
rect 53555 3625 53595 3665
rect 53905 3625 53945 3665
rect 59855 3625 59895 3665
rect 60205 3625 60245 3665
rect 60555 3625 60595 3665
rect 60905 3625 60945 3665
rect 61255 3625 61295 3665
rect 52505 3275 52545 3315
rect 52855 3275 52895 3315
rect 53205 3275 53245 3315
rect 53555 3275 53595 3315
rect 53905 3275 53945 3315
rect 59855 3275 59895 3315
rect 60205 3275 60245 3315
rect 60555 3275 60595 3315
rect 60905 3275 60945 3315
rect 61255 3275 61295 3315
rect 52505 2925 52545 2965
rect 52855 2925 52895 2965
rect 53205 2925 53245 2965
rect 53555 2925 53595 2965
rect 53905 2925 53945 2965
rect 59855 2925 59895 2965
rect 60205 2925 60245 2965
rect 60555 2925 60595 2965
rect 60905 2925 60945 2965
rect 61255 2925 61295 2965
rect 52505 2575 52545 2615
rect 52855 2575 52895 2615
rect 53205 2575 53245 2615
rect 53555 2575 53595 2615
rect 53905 2575 53945 2615
rect 59855 2575 59895 2615
rect 60205 2575 60245 2615
rect 60555 2575 60595 2615
rect 60905 2575 60945 2615
rect 61255 2575 61295 2615
rect 52505 2225 52545 2265
rect 52855 2225 52895 2265
rect 53205 2225 53245 2265
rect 53555 2225 53595 2265
rect 53905 2225 53945 2265
rect 59855 2225 59895 2265
rect 60205 2225 60245 2265
rect 60555 2225 60595 2265
rect 60905 2225 60945 2265
rect 61255 2225 61295 2265
rect 52505 1875 52545 1915
rect 52855 1875 52895 1915
rect 53205 1875 53245 1915
rect 53555 1875 53595 1915
rect 53905 1875 53945 1915
rect 59855 1875 59895 1915
rect 60205 1875 60245 1915
rect 60555 1875 60595 1915
rect 60905 1875 60945 1915
rect 61255 1875 61295 1915
rect 52505 1525 52545 1565
rect 52855 1525 52895 1565
rect 53205 1525 53245 1565
rect 53555 1525 53595 1565
rect 53905 1525 53945 1565
rect 59855 1525 59895 1565
rect 60205 1525 60245 1565
rect 60555 1525 60595 1565
rect 60905 1525 60945 1565
rect 61255 1525 61295 1565
rect 52505 1175 52545 1215
rect 52855 1175 52895 1215
rect 53205 1175 53245 1215
rect 53555 1175 53595 1215
rect 53905 1175 53945 1215
rect 59855 1175 59895 1215
rect 60205 1175 60245 1215
rect 60555 1175 60595 1215
rect 60905 1175 60945 1215
rect 61255 1175 61295 1215
rect 52505 825 52545 865
rect 52855 825 52895 865
rect 53205 825 53245 865
rect 53555 825 53595 865
rect 53905 825 53945 865
rect 59855 825 59895 865
rect 60205 825 60245 865
rect 60555 825 60595 865
rect 60905 825 60945 865
rect 61255 825 61295 865
rect 52505 475 52545 515
rect 52855 475 52895 515
rect 53205 475 53245 515
rect 53555 475 53595 515
rect 53905 475 53945 515
rect 59855 475 59895 515
rect 60205 475 60245 515
rect 60555 475 60595 515
rect 60905 475 60945 515
rect 61255 475 61295 515
rect 52505 125 52545 165
rect 52855 125 52895 165
rect 53205 125 53245 165
rect 53555 125 53595 165
rect 53905 125 53945 165
rect 54255 125 54295 165
rect 54605 125 54645 165
rect 54955 125 54995 165
rect 55305 125 55345 165
rect 55655 125 55695 165
rect 56005 125 56045 165
rect 56355 125 56395 165
rect 56705 125 56745 165
rect 57055 125 57095 165
rect 57405 125 57445 165
rect 57755 125 57795 165
rect 58105 125 58145 165
rect 58455 125 58495 165
rect 58805 125 58845 165
rect 59155 125 59195 165
rect 59505 125 59545 165
rect 59855 125 59895 165
rect 60205 125 60245 165
rect 60555 125 60595 165
rect 60905 125 60945 165
rect 61255 125 61295 165
rect 52505 -225 52545 -185
rect 52855 -225 52895 -185
rect 53205 -225 53245 -185
rect 53555 -225 53595 -185
rect 53905 -225 53945 -185
rect 54255 -225 54295 -185
rect 54605 -225 54645 -185
rect 54955 -225 54995 -185
rect 55305 -225 55345 -185
rect 55655 -225 55695 -185
rect 56005 -225 56045 -185
rect 56355 -225 56395 -185
rect 56705 -225 56745 -185
rect 57055 -225 57095 -185
rect 57405 -225 57445 -185
rect 57755 -225 57795 -185
rect 58105 -225 58145 -185
rect 58455 -225 58495 -185
rect 58805 -225 58845 -185
rect 59155 -225 59195 -185
rect 59505 -225 59545 -185
rect 59855 -225 59895 -185
rect 60205 -225 60245 -185
rect 60555 -225 60595 -185
rect 60905 -225 60945 -185
rect 61255 -225 61295 -185
<< metal4 >>
rect 51855 6190 61545 6195
rect 51855 6150 55785 6190
rect 55825 6150 61545 6190
rect 51855 6145 61545 6150
rect 52500 5765 53250 5770
rect 52500 5725 52505 5765
rect 52545 5725 52855 5765
rect 52895 5725 53205 5765
rect 53245 5725 53250 5765
rect 52500 5720 53250 5725
rect 53200 5420 53250 5720
rect 53550 5765 53600 5770
rect 53550 5725 53555 5765
rect 53595 5725 53600 5765
rect 53550 5420 53600 5725
rect 53900 5765 53950 5770
rect 53900 5725 53905 5765
rect 53945 5725 53950 5765
rect 53900 5420 53950 5725
rect 54250 5765 54300 5770
rect 54250 5725 54255 5765
rect 54295 5725 54300 5765
rect 54250 5420 54300 5725
rect 54600 5765 54650 5770
rect 54600 5725 54605 5765
rect 54645 5725 54650 5765
rect 54600 5420 54650 5725
rect 54950 5765 55000 5770
rect 54950 5725 54955 5765
rect 54995 5725 55000 5765
rect 54950 5420 55000 5725
rect 55300 5765 55350 5770
rect 55300 5725 55305 5765
rect 55345 5725 55350 5765
rect 55300 5420 55350 5725
rect 55650 5765 55700 5770
rect 55650 5725 55655 5765
rect 55695 5725 55700 5765
rect 55650 5420 55700 5725
rect 56000 5765 56050 5770
rect 56000 5725 56005 5765
rect 56045 5725 56050 5765
rect 56000 5420 56050 5725
rect 56350 5765 56400 5770
rect 56350 5725 56355 5765
rect 56395 5725 56400 5765
rect 56350 5420 56400 5725
rect 56700 5765 56750 5770
rect 56700 5725 56705 5765
rect 56745 5725 56750 5765
rect 56700 5420 56750 5725
rect 52500 5415 56750 5420
rect 52500 5375 52505 5415
rect 52545 5375 52855 5415
rect 52895 5375 53205 5415
rect 53245 5375 53555 5415
rect 53595 5375 53905 5415
rect 53945 5375 54255 5415
rect 54295 5375 54605 5415
rect 54645 5375 54955 5415
rect 54995 5375 55305 5415
rect 55345 5375 55655 5415
rect 55695 5375 56005 5415
rect 56045 5375 56355 5415
rect 56395 5375 56705 5415
rect 56745 5375 56750 5415
rect 52500 5370 56750 5375
rect 53200 5070 53250 5370
rect 52500 5065 53950 5070
rect 52500 5025 52505 5065
rect 52545 5025 52855 5065
rect 52895 5025 53205 5065
rect 53245 5025 53555 5065
rect 53595 5025 53905 5065
rect 53945 5025 53950 5065
rect 52500 5020 53950 5025
rect 54250 5065 54300 5370
rect 54250 5025 54255 5065
rect 54295 5025 54300 5065
rect 53200 4720 53250 5020
rect 52500 4715 53950 4720
rect 52500 4675 52505 4715
rect 52545 4675 52855 4715
rect 52895 4675 53205 4715
rect 53245 4675 53555 4715
rect 53595 4675 53905 4715
rect 53945 4675 53950 4715
rect 52500 4670 53950 4675
rect 54250 4715 54300 5025
rect 54250 4675 54255 4715
rect 54295 4675 54300 4715
rect 53200 4370 53250 4670
rect 52500 4365 53950 4370
rect 52500 4325 52505 4365
rect 52545 4325 52855 4365
rect 52895 4325 53205 4365
rect 53245 4325 53555 4365
rect 53595 4325 53905 4365
rect 53945 4325 53950 4365
rect 52500 4320 53950 4325
rect 54250 4365 54300 4675
rect 54250 4325 54255 4365
rect 54295 4325 54300 4365
rect 54250 4320 54300 4325
rect 54600 5065 54650 5370
rect 54600 5025 54605 5065
rect 54645 5025 54650 5065
rect 54600 4715 54650 5025
rect 54600 4675 54605 4715
rect 54645 4675 54650 4715
rect 54600 4365 54650 4675
rect 54600 4325 54605 4365
rect 54645 4325 54650 4365
rect 54600 4320 54650 4325
rect 54950 5065 55000 5370
rect 54950 5025 54955 5065
rect 54995 5025 55000 5065
rect 54950 4715 55000 5025
rect 54950 4675 54955 4715
rect 54995 4675 55000 4715
rect 54950 4365 55000 4675
rect 54950 4325 54955 4365
rect 54995 4325 55000 4365
rect 54950 4320 55000 4325
rect 55300 5065 55350 5370
rect 55300 5025 55305 5065
rect 55345 5025 55350 5065
rect 55300 4715 55350 5025
rect 55650 5055 55700 5370
rect 55650 5015 55655 5055
rect 55695 5015 55700 5055
rect 55650 5010 55700 5015
rect 56000 5055 56050 5370
rect 56000 5015 56005 5055
rect 56045 5015 56050 5055
rect 56000 5010 56050 5015
rect 56350 5055 56400 5370
rect 56350 5015 56355 5055
rect 56395 5015 56400 5055
rect 56350 5010 56400 5015
rect 56700 5055 56750 5370
rect 56700 5015 56705 5055
rect 56745 5015 56750 5055
rect 56700 5010 56750 5015
rect 57050 5765 57100 5770
rect 57050 5725 57055 5765
rect 57095 5725 57100 5765
rect 57050 5420 57100 5725
rect 57400 5765 57450 5770
rect 57400 5725 57405 5765
rect 57445 5725 57450 5765
rect 57400 5420 57450 5725
rect 57750 5765 57800 5770
rect 57750 5725 57755 5765
rect 57795 5725 57800 5765
rect 57750 5420 57800 5725
rect 58100 5765 58150 5770
rect 58100 5725 58105 5765
rect 58145 5725 58150 5765
rect 58100 5420 58150 5725
rect 58450 5765 58500 5770
rect 58450 5725 58455 5765
rect 58495 5725 58500 5765
rect 58450 5420 58500 5725
rect 58800 5765 58850 5770
rect 58800 5725 58805 5765
rect 58845 5725 58850 5765
rect 58800 5420 58850 5725
rect 59150 5765 59200 5770
rect 59150 5725 59155 5765
rect 59195 5725 59200 5765
rect 59150 5420 59200 5725
rect 59500 5765 59550 5770
rect 59500 5725 59505 5765
rect 59545 5725 59550 5765
rect 59500 5420 59550 5725
rect 59850 5765 59900 5770
rect 59850 5725 59855 5765
rect 59895 5725 59900 5765
rect 59850 5420 59900 5725
rect 60200 5765 60250 5770
rect 60200 5725 60205 5765
rect 60245 5725 60250 5765
rect 60200 5420 60250 5725
rect 60550 5765 61300 5770
rect 60550 5725 60555 5765
rect 60595 5725 60905 5765
rect 60945 5725 61255 5765
rect 61295 5725 61300 5765
rect 60550 5720 61300 5725
rect 60550 5420 60600 5720
rect 57050 5415 61300 5420
rect 57050 5375 57055 5415
rect 57095 5375 57405 5415
rect 57445 5375 57755 5415
rect 57795 5375 58105 5415
rect 58145 5375 58455 5415
rect 58495 5375 58805 5415
rect 58845 5375 59155 5415
rect 59195 5375 59505 5415
rect 59545 5375 59855 5415
rect 59895 5375 60205 5415
rect 60245 5375 60555 5415
rect 60595 5375 60905 5415
rect 60945 5375 61255 5415
rect 61295 5375 61300 5415
rect 57050 5370 61300 5375
rect 57050 5055 57100 5370
rect 57050 5015 57055 5055
rect 57095 5015 57100 5055
rect 57050 5010 57100 5015
rect 57400 5055 57450 5370
rect 57400 5015 57405 5055
rect 57445 5015 57450 5055
rect 57400 5010 57450 5015
rect 57750 5055 57800 5370
rect 57750 5015 57755 5055
rect 57795 5015 57800 5055
rect 57750 5010 57800 5015
rect 58100 5055 58150 5370
rect 58100 5015 58105 5055
rect 58145 5015 58150 5055
rect 58100 5010 58150 5015
rect 58450 5065 58500 5370
rect 58450 5025 58455 5065
rect 58495 5025 58500 5065
rect 55300 4675 55305 4715
rect 55345 4675 55350 4715
rect 55300 4365 55350 4675
rect 55300 4325 55305 4365
rect 55345 4325 55350 4365
rect 55300 4320 55350 4325
rect 58450 4715 58500 5025
rect 58450 4675 58455 4715
rect 58495 4675 58500 4715
rect 58450 4365 58500 4675
rect 58450 4325 58455 4365
rect 58495 4325 58500 4365
rect 58450 4320 58500 4325
rect 58800 5065 58850 5370
rect 58800 5025 58805 5065
rect 58845 5025 58850 5065
rect 58800 4715 58850 5025
rect 58800 4675 58805 4715
rect 58845 4675 58850 4715
rect 58800 4365 58850 4675
rect 58800 4325 58805 4365
rect 58845 4325 58850 4365
rect 58800 4320 58850 4325
rect 59150 5065 59200 5370
rect 59150 5025 59155 5065
rect 59195 5025 59200 5065
rect 59150 4715 59200 5025
rect 59150 4675 59155 4715
rect 59195 4675 59200 4715
rect 59150 4365 59200 4675
rect 59150 4325 59155 4365
rect 59195 4325 59200 4365
rect 59150 4320 59200 4325
rect 59500 5065 59550 5370
rect 60550 5070 60600 5370
rect 59500 5025 59505 5065
rect 59545 5025 59550 5065
rect 59500 4715 59550 5025
rect 59850 5065 61300 5070
rect 59850 5025 59855 5065
rect 59895 5025 60205 5065
rect 60245 5025 60555 5065
rect 60595 5025 60905 5065
rect 60945 5025 61255 5065
rect 61295 5025 61300 5065
rect 59850 5020 61300 5025
rect 60550 4720 60600 5020
rect 59500 4675 59505 4715
rect 59545 4675 59550 4715
rect 59500 4365 59550 4675
rect 59850 4715 61300 4720
rect 59850 4675 59855 4715
rect 59895 4675 60205 4715
rect 60245 4675 60555 4715
rect 60595 4675 60905 4715
rect 60945 4675 61255 4715
rect 61295 4675 61300 4715
rect 59850 4670 61300 4675
rect 60550 4370 60600 4670
rect 59500 4325 59505 4365
rect 59545 4325 59550 4365
rect 59500 4320 59550 4325
rect 59850 4365 61300 4370
rect 59850 4325 59855 4365
rect 59895 4325 60205 4365
rect 60245 4325 60555 4365
rect 60595 4325 60905 4365
rect 60945 4325 61255 4365
rect 61295 4325 61300 4365
rect 59850 4320 61300 4325
rect 53200 4020 53250 4320
rect 60550 4020 60600 4320
rect 52500 4015 53950 4020
rect 52500 3975 52505 4015
rect 52545 3975 52855 4015
rect 52895 3975 53205 4015
rect 53245 3975 53555 4015
rect 53595 3975 53905 4015
rect 53945 3975 53950 4015
rect 52500 3970 53950 3975
rect 59850 4015 61300 4020
rect 59850 3975 59855 4015
rect 59895 3975 60205 4015
rect 60245 3975 60555 4015
rect 60595 3975 60905 4015
rect 60945 3975 61255 4015
rect 61295 3975 61300 4015
rect 59850 3970 61300 3975
rect 53200 3670 53250 3970
rect 60550 3670 60600 3970
rect 52500 3665 53950 3670
rect 52500 3625 52505 3665
rect 52545 3625 52855 3665
rect 52895 3625 53205 3665
rect 53245 3625 53555 3665
rect 53595 3625 53905 3665
rect 53945 3625 53950 3665
rect 52500 3620 53950 3625
rect 59850 3665 61300 3670
rect 59850 3625 59855 3665
rect 59895 3625 60205 3665
rect 60245 3625 60555 3665
rect 60595 3625 60905 3665
rect 60945 3625 61255 3665
rect 61295 3625 61300 3665
rect 59850 3620 61300 3625
rect 53200 3320 53250 3620
rect 60550 3320 60600 3620
rect 52500 3315 53950 3320
rect 52500 3275 52505 3315
rect 52545 3275 52855 3315
rect 52895 3275 53205 3315
rect 53245 3275 53555 3315
rect 53595 3275 53905 3315
rect 53945 3275 53950 3315
rect 52500 3270 53950 3275
rect 59850 3315 61300 3320
rect 59850 3275 59855 3315
rect 59895 3275 60205 3315
rect 60245 3275 60555 3315
rect 60595 3275 60905 3315
rect 60945 3275 61255 3315
rect 61295 3275 61300 3315
rect 59850 3270 61300 3275
rect 53200 2970 53250 3270
rect 60550 2970 60600 3270
rect 52500 2965 53950 2970
rect 52500 2925 52505 2965
rect 52545 2925 52855 2965
rect 52895 2925 53205 2965
rect 53245 2925 53555 2965
rect 53595 2925 53905 2965
rect 53945 2925 53950 2965
rect 52500 2920 53950 2925
rect 59850 2965 61300 2970
rect 59850 2925 59855 2965
rect 59895 2925 60205 2965
rect 60245 2925 60555 2965
rect 60595 2925 60905 2965
rect 60945 2925 61255 2965
rect 61295 2925 61300 2965
rect 59850 2920 61300 2925
rect 53200 2620 53250 2920
rect 60550 2620 60600 2920
rect 52500 2615 53950 2620
rect 52500 2575 52505 2615
rect 52545 2575 52855 2615
rect 52895 2575 53205 2615
rect 53245 2575 53555 2615
rect 53595 2575 53905 2615
rect 53945 2575 53950 2615
rect 52500 2570 53950 2575
rect 59850 2615 61300 2620
rect 59850 2575 59855 2615
rect 59895 2575 60205 2615
rect 60245 2575 60555 2615
rect 60595 2575 60905 2615
rect 60945 2575 61255 2615
rect 61295 2575 61300 2615
rect 59850 2570 61300 2575
rect 53200 2270 53250 2570
rect 60550 2270 60600 2570
rect 52500 2265 53950 2270
rect 52500 2225 52505 2265
rect 52545 2225 52855 2265
rect 52895 2225 53205 2265
rect 53245 2225 53555 2265
rect 53595 2225 53905 2265
rect 53945 2225 53950 2265
rect 52500 2220 53950 2225
rect 59850 2265 61300 2270
rect 59850 2225 59855 2265
rect 59895 2225 60205 2265
rect 60245 2225 60555 2265
rect 60595 2225 60905 2265
rect 60945 2225 61255 2265
rect 61295 2225 61300 2265
rect 59850 2220 61300 2225
rect 53200 1920 53250 2220
rect 60550 1920 60600 2220
rect 52500 1915 54360 1920
rect 52500 1875 52505 1915
rect 52545 1875 52855 1915
rect 52895 1875 53205 1915
rect 53245 1875 53555 1915
rect 53595 1875 53905 1915
rect 53945 1875 54315 1915
rect 54355 1875 54360 1915
rect 52500 1870 54360 1875
rect 59440 1915 61300 1920
rect 59440 1875 59445 1915
rect 59485 1875 59855 1915
rect 59895 1875 60205 1915
rect 60245 1875 60555 1915
rect 60595 1875 60905 1915
rect 60945 1875 61255 1915
rect 61295 1875 61300 1915
rect 59440 1870 61300 1875
rect 53200 1570 53250 1870
rect 60550 1570 60600 1870
rect 52500 1565 53950 1570
rect 52500 1525 52505 1565
rect 52545 1525 52855 1565
rect 52895 1525 53205 1565
rect 53245 1525 53555 1565
rect 53595 1525 53905 1565
rect 53945 1525 53950 1565
rect 52500 1520 53950 1525
rect 59850 1565 61300 1570
rect 59850 1525 59855 1565
rect 59895 1525 60205 1565
rect 60245 1525 60555 1565
rect 60595 1525 60905 1565
rect 60945 1525 61255 1565
rect 61295 1525 61300 1565
rect 59850 1520 61300 1525
rect 53200 1220 53250 1520
rect 60550 1220 60600 1520
rect 52500 1215 53950 1220
rect 52500 1175 52505 1215
rect 52545 1175 52855 1215
rect 52895 1175 53205 1215
rect 53245 1175 53555 1215
rect 53595 1175 53905 1215
rect 53945 1175 53950 1215
rect 52500 1170 53950 1175
rect 59850 1215 61300 1220
rect 59850 1175 59855 1215
rect 59895 1175 60205 1215
rect 60245 1175 60555 1215
rect 60595 1175 60905 1215
rect 60945 1175 61255 1215
rect 61295 1175 61300 1215
rect 59850 1170 61300 1175
rect 53200 870 53250 1170
rect 60550 870 60600 1170
rect 52500 865 53950 870
rect 52500 825 52505 865
rect 52545 825 52855 865
rect 52895 825 53205 865
rect 53245 825 53555 865
rect 53595 825 53905 865
rect 53945 825 53950 865
rect 52500 820 53950 825
rect 59850 865 61300 870
rect 59850 825 59855 865
rect 59895 825 60205 865
rect 60245 825 60555 865
rect 60595 825 60905 865
rect 60945 825 61255 865
rect 61295 825 61300 865
rect 59850 820 61300 825
rect 53200 520 53250 820
rect 60550 520 60600 820
rect 52500 515 53950 520
rect 52500 475 52505 515
rect 52545 475 52855 515
rect 52895 475 53205 515
rect 53245 475 53555 515
rect 53595 475 53905 515
rect 53945 475 53950 515
rect 52500 470 53950 475
rect 59850 515 61300 520
rect 59850 475 59855 515
rect 59895 475 60205 515
rect 60245 475 60555 515
rect 60595 475 60905 515
rect 60945 475 61255 515
rect 61295 475 61300 515
rect 59850 470 61300 475
rect 53200 170 53250 470
rect 60550 170 60600 470
rect 52500 165 56750 170
rect 52500 125 52505 165
rect 52545 125 52855 165
rect 52895 125 53205 165
rect 53245 125 53555 165
rect 53595 125 53905 165
rect 53945 125 54255 165
rect 54295 125 54605 165
rect 54645 125 54955 165
rect 54995 125 55305 165
rect 55345 125 55655 165
rect 55695 125 56005 165
rect 56045 125 56355 165
rect 56395 125 56705 165
rect 56745 125 56750 165
rect 52500 120 56750 125
rect 53200 -180 53250 120
rect 52500 -185 53250 -180
rect 52500 -225 52505 -185
rect 52545 -225 52855 -185
rect 52895 -225 53205 -185
rect 53245 -225 53250 -185
rect 52500 -230 53250 -225
rect 53550 -185 53600 120
rect 53550 -225 53555 -185
rect 53595 -225 53600 -185
rect 53550 -230 53600 -225
rect 53900 -185 53950 120
rect 53900 -225 53905 -185
rect 53945 -225 53950 -185
rect 53900 -230 53950 -225
rect 54250 -185 54300 120
rect 54250 -225 54255 -185
rect 54295 -225 54300 -185
rect 54250 -230 54300 -225
rect 54600 -185 54650 120
rect 54600 -225 54605 -185
rect 54645 -225 54650 -185
rect 54600 -230 54650 -225
rect 54950 -185 55000 120
rect 54950 -225 54955 -185
rect 54995 -225 55000 -185
rect 54950 -230 55000 -225
rect 55300 -185 55350 120
rect 55300 -225 55305 -185
rect 55345 -225 55350 -185
rect 55300 -230 55350 -225
rect 55650 -185 55700 120
rect 55650 -225 55655 -185
rect 55695 -225 55700 -185
rect 55650 -230 55700 -225
rect 56000 -185 56050 120
rect 56000 -225 56005 -185
rect 56045 -225 56050 -185
rect 56000 -230 56050 -225
rect 56350 -185 56400 120
rect 56350 -225 56355 -185
rect 56395 -225 56400 -185
rect 56350 -230 56400 -225
rect 56700 -185 56750 120
rect 56700 -225 56705 -185
rect 56745 -225 56750 -185
rect 56700 -230 56750 -225
rect 57050 165 61300 170
rect 57050 125 57055 165
rect 57095 125 57405 165
rect 57445 125 57755 165
rect 57795 125 58105 165
rect 58145 125 58455 165
rect 58495 125 58805 165
rect 58845 125 59155 165
rect 59195 125 59505 165
rect 59545 125 59855 165
rect 59895 125 60205 165
rect 60245 125 60555 165
rect 60595 125 60905 165
rect 60945 125 61255 165
rect 61295 125 61300 165
rect 57050 120 61300 125
rect 57050 -185 57100 120
rect 57050 -225 57055 -185
rect 57095 -225 57100 -185
rect 57050 -230 57100 -225
rect 57400 -185 57450 120
rect 57400 -225 57405 -185
rect 57445 -225 57450 -185
rect 57400 -230 57450 -225
rect 57750 -185 57800 120
rect 57750 -225 57755 -185
rect 57795 -225 57800 -185
rect 57750 -230 57800 -225
rect 58100 -185 58150 120
rect 58100 -225 58105 -185
rect 58145 -225 58150 -185
rect 58100 -230 58150 -225
rect 58450 -185 58500 120
rect 58450 -225 58455 -185
rect 58495 -225 58500 -185
rect 58450 -230 58500 -225
rect 58800 -185 58850 120
rect 58800 -225 58805 -185
rect 58845 -225 58850 -185
rect 58800 -230 58850 -225
rect 59150 -185 59200 120
rect 59150 -225 59155 -185
rect 59195 -225 59200 -185
rect 59150 -230 59200 -225
rect 59500 -185 59550 120
rect 59500 -225 59505 -185
rect 59545 -225 59550 -185
rect 59500 -230 59550 -225
rect 59850 -185 59900 120
rect 59850 -225 59855 -185
rect 59895 -225 59900 -185
rect 59850 -230 59900 -225
rect 60200 -185 60250 120
rect 60200 -225 60205 -185
rect 60245 -225 60250 -185
rect 60200 -230 60250 -225
rect 60550 -180 60600 120
rect 60550 -185 61300 -180
rect 60550 -225 60555 -185
rect 60595 -225 60905 -185
rect 60945 -225 61255 -185
rect 61295 -225 61300 -185
rect 60550 -230 61300 -225
rect 51855 -510 61545 -505
rect 51855 -550 57975 -510
rect 58015 -550 61545 -510
rect 51855 -555 61545 -550
<< labels >>
flabel metal4 51855 -530 51855 -530 7 FreeSans 800 0 -400 0 GNDA
port 16 w
flabel metal1 55850 2235 55850 2235 1 FreeSans 200 0 0 80 Vb1
port 6 n
flabel metal2 56190 1880 56190 1880 7 FreeSans 200 0 -80 0 VD1
flabel metal1 56555 1840 56555 1840 3 FreeSans 200 0 80 0 VD2
flabel metal2 57720 1410 57720 1410 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal1 56900 1375 56900 1375 3 FreeSans 200 0 80 0 V_p_mir
flabel metal1 57220 1360 57220 1360 3 FreeSans 200 0 80 0 V_p
flabel metal1 56920 2910 56920 2910 3 FreeSans 200 0 80 0 V_tot
flabel metal2 57570 2730 57570 2730 3 FreeSans 200 0 80 0 err_amp_mir
flabel metal2 55960 2790 55960 2790 7 FreeSans 200 0 -80 0 V_err_amp_ref
port 12 w
flabel metal2 57185 2675 57185 2675 7 FreeSans 200 0 -80 0 err_amp_out
flabel metal1 57210 3065 57210 3065 3 FreeSans 200 0 80 0 V_err_p
flabel metal1 56660 3030 56660 3030 3 FreeSans 200 0 80 0 V_err_mir_p
flabel metal1 56505 3045 56505 3045 7 FreeSans 200 0 -80 0 V_err_gate
port 13 w
flabel metal2 54810 2155 54810 2155 1 FreeSans 200 0 0 80 V_CMFB_S1
port 2 n
flabel metal2 54855 1965 54855 1965 1 FreeSans 200 0 0 80 V_CMFB_S2
port 7 n
flabel metal3 54605 3460 54605 3460 7 FreeSans 200 0 -80 0 cap_res_X
flabel metal2 54335 1335 54335 1335 5 FreeSans 200 0 0 -80 VOUT-
port 9 s
flabel metal2 59465 1335 59465 1335 5 FreeSans 200 0 0 -80 VOUT+
port 10 s
flabel metal3 59195 3460 59195 3460 3 FreeSans 200 0 80 0 cap_res_Y
flabel metal2 58950 1965 58950 1965 1 FreeSans 200 0 0 80 V_CMFB_S4
port 8 n
flabel metal2 58995 2155 58995 2155 1 FreeSans 200 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 56280 2575 56280 2575 3 FreeSans 200 0 80 0 X
flabel metal1 57520 2575 57520 2575 7 FreeSans 200 0 -80 0 Y
flabel metal1 57900 4040 57900 4040 3 FreeSans 200 0 80 0 VD4
flabel metal1 55900 4030 55900 4030 7 FreeSans 200 0 -80 0 VD3
flabel metal2 57000 3545 57000 3545 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56870 3580 56870 3580 5 FreeSans 200 0 0 -80 Vb2
port 5 s
flabel metal2 57320 4870 57320 4870 1 FreeSans 200 0 0 80 Vb2_Vb3
flabel metal4 51855 6170 51855 6170 7 FreeSans 800 0 -400 0 VDDA
port 1 w
flabel metal2 55960 1745 55960 1745 7 FreeSans 200 0 -80 0 VIN-
port 15 w
flabel metal2 55960 1525 55960 1525 7 FreeSans 200 0 -80 0 VIN+
port 14 w
<< end >>
