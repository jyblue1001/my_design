** sch_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/phase_frequency_detector.sch
**.subckt phase_frequency_detector F_REF F_VCO QA QB VPWR VPB VGND
*.ipin F_REF
*.opin QA
*.ipin F_VCO
*.opin QB
*.ipin VDDA
*.ipin GNDA
x1 F_REF QA VGND VNB VPB VPWR QA_b sky130_fd_sc_hd__nor2_1
x2 E QA_b VGND VNB VPB VPWR QA sky130_fd_sc_hd__nor2_1
x3 QA_b E_b VGND VNB VPB VPWR E sky130_fd_sc_hd__nor2_1
x4 Reset E VGND VNB VPB VPWR E_b sky130_fd_sc_hd__nor2_1
x5 F_VCO QB VGND VNB VPB VPWR QB_b sky130_fd_sc_hd__nor2_1
x6 F QB_b VGND VNB VPB VPWR QB sky130_fd_sc_hd__nor2_1
x7 QB_b F_b VGND VNB VPB VPWR F sky130_fd_sc_hd__nor2_1
x8 Reset F VGND VNB VPB VPWR F_b sky130_fd_sc_hd__nor2_1
x9 QB QA VGND VNB VPB VPWR before_Reset sky130_fd_sc_hd__nand2_1
x10 before_Reset VGND VNB VPB VPWR net1 sky130_fd_sc_hd__inv_1
x11 net1 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__inv_1
x12 net2 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_1
x13 net3 VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_1
x14 net4 VGND VNB VPB VPWR Reset sky130_fd_sc_hd__inv_1
**.ends
.end
