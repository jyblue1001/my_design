magic
tech sky130A
timestamp 1751775419
<< error_s >>
rect 4011 4080 4079 4084
rect 4025 4066 4065 4070
rect 3961 3686 3970 3754
rect 3975 3700 3984 3740
rect 5286 3595 5354 3604
rect 5386 3595 5454 3604
rect 5496 3595 5564 3604
rect 5606 3595 5674 3604
rect 5716 3595 5784 3604
rect 5300 3581 5340 3590
rect 5400 3581 5440 3590
rect 5510 3581 5550 3590
rect 5620 3581 5660 3590
rect 5730 3581 5770 3590
rect 6101 3585 6110 3625
rect 6115 3571 6124 3639
rect 5011 3265 5020 3305
rect 4071 2410 4080 3240
rect 4085 2410 4094 3254
rect 5025 3251 5034 3319
rect 5025 2875 5065 2887
rect 5035 2858 5055 2870
<< locali >>
rect 5035 2830 5055 2870
<< metal1 >>
rect 2055 11725 2095 11730
rect 2055 11695 2060 11725
rect 2090 11695 2095 11725
rect 2055 11690 2095 11695
rect 3315 11725 3355 11730
rect 3315 11695 3320 11725
rect 3350 11695 3355 11725
rect 3315 11690 3355 11695
rect 2005 11670 2045 11675
rect 2005 11640 2010 11670
rect 2040 11640 2045 11670
rect 2005 11635 2045 11640
rect 1855 10085 1895 10090
rect 1855 10055 1860 10085
rect 1890 10055 1895 10085
rect 1855 10050 1895 10055
rect 475 9335 515 9340
rect 475 9305 480 9335
rect 510 9305 515 9335
rect 475 9300 515 9305
rect 485 890 505 9300
rect 1865 6445 1885 10050
rect 1905 9015 1945 9020
rect 1905 8985 1910 9015
rect 1940 8985 1945 9015
rect 1905 8980 1945 8985
rect 1915 6495 1935 8980
rect 1955 8770 1995 8775
rect 1955 8740 1960 8770
rect 1990 8740 1995 8770
rect 1955 8735 1995 8740
rect 1965 6545 1985 8735
rect 2015 6595 2035 11635
rect 2065 6645 2085 11690
rect 3205 11670 3245 11675
rect 3205 11640 3210 11670
rect 3240 11640 3245 11670
rect 3205 11635 3245 11640
rect 3215 11550 3235 11635
rect 3325 11550 3345 11690
rect 4655 11590 4695 11595
rect 4655 11560 4660 11590
rect 4690 11560 4695 11590
rect 4655 11555 4695 11560
rect 8435 11590 8475 11595
rect 8435 11560 8440 11590
rect 8470 11560 8475 11590
rect 8435 11555 8475 11560
rect 4665 11550 4685 11555
rect 4040 11545 4080 11550
rect 4040 11515 4045 11545
rect 4075 11515 4080 11545
rect 4040 11510 4080 11515
rect 8365 11545 8405 11550
rect 8365 11515 8370 11545
rect 8400 11515 8405 11545
rect 8365 11510 8405 11515
rect 3820 11495 3860 11500
rect 3820 11465 3825 11495
rect 3855 11465 3860 11495
rect 3820 11460 3860 11465
rect 8315 11495 8355 11500
rect 8315 11465 8320 11495
rect 8350 11465 8355 11495
rect 8315 11460 8355 11465
rect 2105 8495 2145 8500
rect 2105 8465 2110 8495
rect 2140 8465 2145 8495
rect 2105 8460 2145 8465
rect 2115 6695 2135 8460
rect 2105 6690 2145 6695
rect 2105 6660 2110 6690
rect 2140 6660 2145 6690
rect 2105 6655 2145 6660
rect 7120 6690 7160 6695
rect 7120 6660 7125 6690
rect 7155 6660 7160 6690
rect 7120 6655 7160 6660
rect 2055 6640 2095 6645
rect 2055 6610 2060 6640
rect 2090 6610 2095 6640
rect 2055 6605 2095 6610
rect 7070 6640 7110 6645
rect 7070 6610 7075 6640
rect 7105 6610 7110 6640
rect 7070 6605 7110 6610
rect 2005 6590 2045 6595
rect 2005 6560 2010 6590
rect 2040 6560 2045 6590
rect 2005 6555 2045 6560
rect 2985 6590 3025 6595
rect 2985 6560 2990 6590
rect 3020 6560 3025 6590
rect 2985 6555 3025 6560
rect 6070 6590 6110 6595
rect 6070 6560 6075 6590
rect 6105 6560 6110 6590
rect 6070 6555 6110 6560
rect 1955 6540 1995 6545
rect 1955 6510 1960 6540
rect 1990 6510 1995 6540
rect 1955 6505 1995 6510
rect 2935 6540 2975 6545
rect 2935 6510 2940 6540
rect 2970 6510 2975 6540
rect 2935 6505 2975 6510
rect 1905 6490 1945 6495
rect 1905 6460 1910 6490
rect 1940 6460 1945 6490
rect 1905 6455 1945 6460
rect 1855 6440 1895 6445
rect 1855 6410 1860 6440
rect 1890 6410 1895 6440
rect 1855 6405 1895 6410
rect 2890 6440 2930 6445
rect 2890 6410 2895 6440
rect 2925 6410 2930 6440
rect 2890 6405 2930 6410
rect 2900 4070 2920 6405
rect 2890 4065 2930 4070
rect 2890 4035 2895 4065
rect 2925 4035 2930 4065
rect 2890 4030 2930 4035
rect 2945 2710 2965 6505
rect 2990 2520 3010 6555
rect 3975 6490 4015 6495
rect 3975 6460 3980 6490
rect 4010 6460 4015 6490
rect 3975 6455 4015 6460
rect 3985 3740 4005 6455
rect 4025 4065 4065 4070
rect 4025 4035 4030 4065
rect 4060 4035 4065 4065
rect 4025 4030 4065 4035
rect 3975 3735 4015 3740
rect 3975 3705 3980 3735
rect 4010 3705 4015 3735
rect 3975 3700 4015 3705
rect 4035 3365 4055 4030
rect 4075 3735 4115 3740
rect 4075 3705 4080 3735
rect 4110 3705 4115 3735
rect 4075 3700 4115 3705
rect 4025 3360 4065 3365
rect 4025 3330 4030 3360
rect 4060 3330 4065 3360
rect 4025 3325 4065 3330
rect 4085 2410 4105 3700
rect 6080 3625 6100 6555
rect 6120 6540 6160 6545
rect 6120 6510 6125 6540
rect 6155 6510 6160 6540
rect 6120 6505 6160 6510
rect 6130 4950 6150 6505
rect 6425 6495 6465 6500
rect 6425 6465 6430 6495
rect 6460 6465 6465 6495
rect 6425 6460 6465 6465
rect 6120 4945 6160 4950
rect 6120 4915 6125 4945
rect 6155 4915 6160 4945
rect 6120 4910 6160 4915
rect 6435 4850 6455 6460
rect 6425 4845 6465 4850
rect 6425 4815 6430 4845
rect 6460 4815 6465 4845
rect 6425 4810 6465 4815
rect 4980 3620 5020 3625
rect 4980 3590 4985 3620
rect 5015 3590 5020 3620
rect 4980 3585 5020 3590
rect 6070 3620 6110 3625
rect 6070 3590 6075 3620
rect 6105 3590 6110 3620
rect 6070 3585 6110 3590
rect 4990 3305 5010 3585
rect 4980 3300 5020 3305
rect 4980 3270 4985 3300
rect 5015 3270 5020 3300
rect 4980 3265 5020 3270
rect 7085 2520 7105 6605
rect 7130 2710 7150 6655
rect 8325 6545 8345 11460
rect 8375 6595 8395 11510
rect 8365 6590 8405 6595
rect 8365 6560 8370 6590
rect 8400 6560 8405 6590
rect 8365 6555 8405 6560
rect 8315 6540 8355 6545
rect 8315 6510 8320 6540
rect 8350 6510 8355 6540
rect 8315 6505 8355 6510
rect 8445 6500 8465 11555
rect 8435 6495 8475 6500
rect 8435 6465 8440 6495
rect 8470 6465 8475 6495
rect 8435 6460 8475 6465
rect 4075 2405 4115 2410
rect 4075 2375 4080 2405
rect 4110 2375 4115 2405
rect 4075 2370 4115 2375
rect 2460 2225 2500 2265
rect 7590 2225 7630 2265
rect 3985 890 4005 1260
rect 475 885 515 890
rect 475 855 480 885
rect 510 855 515 885
rect 475 850 515 855
rect 3975 885 4015 890
rect 3975 855 3980 885
rect 4010 855 4015 885
rect 3975 850 4015 855
<< via1 >>
rect 2060 11695 2090 11725
rect 3320 11695 3350 11725
rect 2010 11640 2040 11670
rect 1860 10055 1890 10085
rect 480 9305 510 9335
rect 1910 8985 1940 9015
rect 1960 8740 1990 8770
rect 3210 11640 3240 11670
rect 4660 11560 4690 11590
rect 8440 11560 8470 11590
rect 4045 11515 4075 11545
rect 8370 11515 8400 11545
rect 3825 11465 3855 11495
rect 8320 11465 8350 11495
rect 2110 8465 2140 8495
rect 2110 6660 2140 6690
rect 7125 6660 7155 6690
rect 2060 6610 2090 6640
rect 7075 6610 7105 6640
rect 2010 6560 2040 6590
rect 2990 6560 3020 6590
rect 6075 6560 6105 6590
rect 1960 6510 1990 6540
rect 2940 6510 2970 6540
rect 1910 6460 1940 6490
rect 1860 6410 1890 6440
rect 2895 6410 2925 6440
rect 2895 4035 2925 4065
rect 3980 6460 4010 6490
rect 4030 4035 4060 4065
rect 3980 3705 4010 3735
rect 4080 3705 4110 3735
rect 4030 3330 4060 3360
rect 6125 6510 6155 6540
rect 6430 6465 6460 6495
rect 6125 4915 6155 4945
rect 6430 4815 6460 4845
rect 4985 3590 5015 3620
rect 6075 3590 6105 3620
rect 4985 3270 5015 3300
rect 8370 6560 8400 6590
rect 8320 6510 8350 6540
rect 8440 6465 8470 6495
rect 4080 2375 4110 2405
rect 480 855 510 885
rect 3980 855 4010 885
<< metal2 >>
rect 2055 11725 2095 11730
rect 2055 11695 2060 11725
rect 2090 11720 2095 11725
rect 3315 11725 3355 11730
rect 3315 11720 3320 11725
rect 2090 11700 3320 11720
rect 2090 11695 2095 11700
rect 2055 11690 2095 11695
rect 3315 11695 3320 11700
rect 3350 11695 3355 11725
rect 3315 11690 3355 11695
rect 2005 11670 2045 11675
rect 2005 11640 2010 11670
rect 2040 11665 2045 11670
rect 3205 11670 3245 11675
rect 3205 11665 3210 11670
rect 2040 11645 3210 11665
rect 2040 11640 2045 11645
rect 2005 11635 2045 11640
rect 3205 11640 3210 11645
rect 3240 11640 3245 11670
rect 3205 11635 3245 11640
rect 4655 11590 4695 11595
rect 4655 11560 4660 11590
rect 4690 11585 4695 11590
rect 8435 11590 8475 11595
rect 8435 11585 8440 11590
rect 4690 11565 8440 11585
rect 4690 11560 4695 11565
rect 4655 11555 4695 11560
rect 8435 11560 8440 11565
rect 8470 11560 8475 11590
rect 8435 11555 8475 11560
rect 4040 11545 4080 11550
rect 4040 11515 4045 11545
rect 4075 11540 4080 11545
rect 8365 11545 8405 11550
rect 8365 11540 8370 11545
rect 4075 11520 8370 11540
rect 4075 11515 4080 11520
rect 4040 11510 4080 11515
rect 8365 11515 8370 11520
rect 8400 11515 8405 11545
rect 8365 11510 8405 11515
rect 3820 11495 3860 11500
rect 3820 11465 3825 11495
rect 3855 11490 3860 11495
rect 8315 11495 8355 11500
rect 8315 11490 8320 11495
rect 3855 11470 8320 11490
rect 3855 11465 3860 11470
rect 3820 11460 3860 11465
rect 8315 11465 8320 11470
rect 8350 11465 8355 11495
rect 8315 11460 8355 11465
rect 1855 10085 1895 10090
rect 1855 10055 1860 10085
rect 1890 10080 1895 10085
rect 1890 10060 1930 10080
rect 1890 10055 1895 10060
rect 1855 10050 1895 10055
rect 475 9335 515 9340
rect 475 9305 480 9335
rect 510 9330 515 9335
rect 510 9310 1930 9330
rect 510 9305 515 9310
rect 475 9300 515 9305
rect 1905 9015 1945 9020
rect 1905 8985 1910 9015
rect 1940 8985 1945 9015
rect 1905 8980 1945 8985
rect 1955 8770 1995 8775
rect 1955 8740 1960 8770
rect 1990 8740 1995 8770
rect 1955 8735 1995 8740
rect 2105 8495 2145 8500
rect 2105 8465 2110 8495
rect 2140 8465 2145 8495
rect 2105 8460 2145 8465
rect 2105 6690 2145 6695
rect 2105 6660 2110 6690
rect 2140 6685 2145 6690
rect 7120 6690 7160 6695
rect 7120 6685 7125 6690
rect 2140 6665 7125 6685
rect 2140 6660 2145 6665
rect 2105 6655 2145 6660
rect 7120 6660 7125 6665
rect 7155 6660 7160 6690
rect 7120 6655 7160 6660
rect 2055 6640 2095 6645
rect 2055 6610 2060 6640
rect 2090 6635 2095 6640
rect 7070 6640 7110 6645
rect 7070 6635 7075 6640
rect 2090 6615 7075 6635
rect 2090 6610 2095 6615
rect 2055 6605 2095 6610
rect 7070 6610 7075 6615
rect 7105 6610 7110 6640
rect 7070 6605 7110 6610
rect 2005 6590 2045 6595
rect 2005 6560 2010 6590
rect 2040 6585 2045 6590
rect 2985 6590 3025 6595
rect 2985 6585 2990 6590
rect 2040 6565 2990 6585
rect 2040 6560 2045 6565
rect 2005 6555 2045 6560
rect 2985 6560 2990 6565
rect 3020 6560 3025 6590
rect 2985 6555 3025 6560
rect 6070 6590 6110 6595
rect 6070 6560 6075 6590
rect 6105 6585 6110 6590
rect 8365 6590 8405 6595
rect 8365 6585 8370 6590
rect 6105 6565 8370 6585
rect 6105 6560 6110 6565
rect 6070 6555 6110 6560
rect 8365 6560 8370 6565
rect 8400 6560 8405 6590
rect 8365 6555 8405 6560
rect 1955 6540 1995 6545
rect 1955 6510 1960 6540
rect 1990 6535 1995 6540
rect 2935 6540 2975 6545
rect 2935 6535 2940 6540
rect 1990 6515 2940 6535
rect 1990 6510 1995 6515
rect 1955 6505 1995 6510
rect 2935 6510 2940 6515
rect 2970 6510 2975 6540
rect 2935 6505 2975 6510
rect 6120 6540 6160 6545
rect 6120 6510 6125 6540
rect 6155 6535 6160 6540
rect 8315 6540 8355 6545
rect 8315 6535 8320 6540
rect 6155 6515 8320 6535
rect 6155 6510 6160 6515
rect 6120 6505 6160 6510
rect 8315 6510 8320 6515
rect 8350 6510 8355 6540
rect 8315 6505 8355 6510
rect 6425 6495 6465 6500
rect 1905 6490 1945 6495
rect 1905 6460 1910 6490
rect 1940 6485 1945 6490
rect 3975 6490 4015 6495
rect 3975 6485 3980 6490
rect 1940 6465 3980 6485
rect 1940 6460 1945 6465
rect 1905 6455 1945 6460
rect 3975 6460 3980 6465
rect 4010 6460 4015 6490
rect 6425 6465 6430 6495
rect 6460 6490 6465 6495
rect 8435 6495 8475 6500
rect 8435 6490 8440 6495
rect 6460 6470 8440 6490
rect 6460 6465 6465 6470
rect 6425 6460 6465 6465
rect 8435 6465 8440 6470
rect 8470 6465 8475 6495
rect 8435 6460 8475 6465
rect 3975 6455 4015 6460
rect 1855 6440 1895 6445
rect 1855 6410 1860 6440
rect 1890 6435 1895 6440
rect 2890 6440 2930 6445
rect 2890 6435 2895 6440
rect 1890 6415 2895 6435
rect 1890 6410 1895 6415
rect 1855 6405 1895 6410
rect 2890 6410 2895 6415
rect 2925 6410 2930 6440
rect 2890 6405 2930 6410
rect 6120 4945 6160 4950
rect 6120 4940 6125 4945
rect 5795 4920 6125 4940
rect 6120 4915 6125 4920
rect 6155 4915 6160 4945
rect 6120 4910 6160 4915
rect 6425 4845 6465 4850
rect 6425 4840 6430 4845
rect 5745 4820 6430 4840
rect 6425 4815 6430 4820
rect 6460 4815 6465 4845
rect 6425 4810 6465 4815
rect 2890 4065 2930 4070
rect 2890 4035 2895 4065
rect 2925 4060 2930 4065
rect 4025 4065 4065 4070
rect 4025 4060 4030 4065
rect 2925 4040 4030 4060
rect 2925 4035 2930 4040
rect 2890 4030 2930 4035
rect 4025 4035 4030 4040
rect 4060 4035 4065 4065
rect 4025 4030 4065 4035
rect 3975 3735 4015 3740
rect 3975 3705 3980 3735
rect 4010 3730 4015 3735
rect 4075 3735 4115 3740
rect 4075 3730 4080 3735
rect 4010 3710 4080 3730
rect 4010 3705 4015 3710
rect 3975 3700 4015 3705
rect 4075 3705 4080 3710
rect 4110 3705 4115 3735
rect 4075 3700 4115 3705
rect 4980 3620 5020 3625
rect 4980 3590 4985 3620
rect 5015 3615 5020 3620
rect 6070 3620 6110 3625
rect 6070 3615 6075 3620
rect 5015 3595 6075 3615
rect 5015 3590 5020 3595
rect 4980 3585 5020 3590
rect 6070 3590 6075 3595
rect 6105 3590 6110 3620
rect 6070 3585 6110 3590
rect 4025 3360 4065 3365
rect 4025 3330 4030 3360
rect 4060 3355 4065 3360
rect 4060 3335 4110 3355
rect 4060 3330 4065 3335
rect 4025 3325 4065 3330
rect 4980 3300 5020 3305
rect 4980 3295 4985 3300
rect 4860 3275 4985 3295
rect 4980 3270 4985 3275
rect 5015 3270 5020 3300
rect 4980 3265 5020 3270
rect 4075 2405 4115 2410
rect 4075 2375 4080 2405
rect 4110 2400 4115 2405
rect 4110 2380 4965 2400
rect 4110 2375 4115 2380
rect 4075 2370 4115 2375
rect 4090 2290 4105 2310
rect 2460 2225 2500 2265
rect 7590 2225 7630 2265
rect 4090 2070 4105 2090
rect 475 885 515 890
rect 475 855 480 885
rect 510 880 515 885
rect 3975 885 4015 890
rect 3975 880 3980 885
rect 510 860 3980 880
rect 510 855 515 860
rect 475 850 515 855
rect 3975 855 3980 860
rect 4010 855 4015 885
rect 3975 850 4015 855
<< metal3 >>
rect 9840 6880 9890 6885
rect 9840 6840 9845 6880
rect 9885 6840 9890 6880
rect 9840 6835 9890 6840
rect 9845 50 9885 6835
rect 9840 45 9890 50
rect 9840 5 9845 45
rect 9885 5 9890 45
rect 9840 0 9890 5
<< via3 >>
rect 9845 6840 9885 6880
rect 9845 5 9885 45
<< metal4 >>
rect 8145 6880 9890 6885
rect 8145 6840 9845 6880
rect 9885 6840 9890 6880
rect 8145 6835 9890 6840
rect 940 6700 990 6750
rect 975 0 1025 50
rect 9685 45 9890 50
rect 9685 5 9845 45
rect 9885 5 9890 45
rect 9685 0 9890 5
use bgr  bgr_0
timestamp 1751725295
transform -1 0 8030 0 -1 12100
box -200 535 6100 5350
use two_stage_opamp_dummy_magic  two_stage_opamp_dummy_magic_0
timestamp 1751775338
transform 1 0 -51855 0 1 555
box 51855 -555 61545 6195
<< labels >>
flabel metal4 965 6750 965 6750 1 FreeSans 800 0 0 400 VDDA
port 1 n
flabel metal4 1000 0 1000 0 5 FreeSans 800 0 0 -400 GNDA
port 2 s
flabel metal2 2480 2225 2480 2225 5 FreeSans 400 0 0 -200 VOUT-
port 4 s
flabel metal2 7610 2225 7610 2225 5 FreeSans 400 0 0 -200 VOUT+
port 3 s
flabel metal2 4090 2300 4090 2300 7 FreeSans 400 0 -200 0 VIN-
port 6 w
flabel metal2 4090 2080 4090 2080 7 FreeSans 400 0 -200 0 VIN+
port 5 w
<< end >>
