magic
tech sky130A
timestamp 1751783180
<< metal1 >>
rect 3315 11775 3355 11780
rect 3315 11745 3320 11775
rect 3350 11745 3355 11775
rect 2005 11670 2045 11675
rect 2005 11640 2010 11670
rect 2040 11640 2045 11670
rect 1840 10085 1880 10090
rect 1840 10055 1845 10085
rect 1875 10055 1880 10085
rect 475 9335 515 9340
rect 475 9305 480 9335
rect 510 9305 515 9335
rect 475 885 515 9305
rect 1840 6450 1880 10055
rect 1895 9015 1935 9020
rect 1895 8985 1900 9015
rect 1930 8985 1935 9015
rect 1895 6505 1935 8985
rect 1950 8770 1990 8775
rect 1950 8740 1955 8770
rect 1985 8740 1990 8770
rect 1950 6560 1990 8740
rect 2005 6615 2045 11640
rect 3205 11670 3245 11675
rect 3205 11640 3210 11670
rect 3240 11640 3245 11670
rect 3205 11325 3245 11640
rect 3315 11380 3355 11745
rect 8505 11775 8545 11780
rect 8505 11745 8510 11775
rect 8540 11745 8545 11775
rect 4655 11720 4695 11725
rect 4655 11690 4660 11720
rect 4690 11690 4695 11720
rect 4040 11665 4080 11670
rect 4040 11635 4045 11665
rect 4075 11635 4080 11665
rect 3820 11610 3860 11615
rect 3820 11580 3825 11610
rect 3855 11580 3860 11610
rect 3820 11325 3860 11580
rect 4040 11325 4080 11635
rect 4655 11325 4695 11690
rect 8435 11720 8475 11725
rect 8435 11690 8440 11720
rect 8470 11690 8475 11720
rect 8370 11665 8410 11670
rect 8370 11635 8375 11665
rect 8405 11635 8410 11665
rect 8315 11610 8355 11615
rect 8315 11580 8320 11610
rect 8350 11580 8355 11610
rect 2105 8495 2145 8500
rect 2105 8465 2110 8495
rect 2140 8465 2145 8495
rect 2105 6680 2145 8465
rect 2105 6650 2110 6680
rect 2140 6650 2145 6680
rect 2105 6645 2145 6650
rect 7150 6680 7190 6685
rect 7150 6650 7155 6680
rect 7185 6650 7190 6680
rect 2005 6585 2010 6615
rect 2040 6585 2045 6615
rect 2005 6580 2045 6585
rect 2955 6615 2995 6620
rect 2955 6585 2960 6615
rect 2990 6585 2995 6615
rect 1950 6530 1955 6560
rect 1985 6530 1990 6560
rect 1950 6525 1990 6530
rect 2900 6560 2940 6565
rect 2900 6530 2905 6560
rect 2935 6530 2940 6560
rect 1895 6475 1900 6505
rect 1930 6475 1935 6505
rect 1895 6470 1935 6475
rect 2550 6505 2590 6510
rect 2550 6475 2555 6505
rect 2585 6475 2590 6505
rect 1840 6420 1845 6450
rect 1875 6420 1880 6450
rect 1840 6415 1880 6420
rect 2550 4065 2590 6475
rect 2550 4035 2555 4065
rect 2585 4035 2590 4065
rect 2550 4030 2590 4035
rect 2605 6450 2645 6455
rect 2605 6420 2610 6450
rect 2640 6420 2645 6450
rect 2605 4010 2645 6420
rect 2605 3980 2610 4010
rect 2640 3980 2645 4010
rect 2605 3975 2645 3980
rect 2900 2710 2940 6530
rect 2955 2520 2995 6585
rect 7095 6615 7135 6620
rect 7095 6585 7100 6615
rect 7130 6585 7135 6615
rect 6060 6560 6100 6565
rect 6060 6530 6065 6560
rect 6095 6530 6100 6560
rect 4095 4065 4135 4070
rect 4095 4035 4100 4065
rect 4130 4035 4135 4065
rect 4025 4010 4065 4015
rect 4025 3980 4030 4010
rect 4060 3980 4065 4010
rect 4025 3405 4065 3980
rect 4025 3375 4030 3405
rect 4060 3375 4065 3405
rect 4025 3370 4065 3375
rect 4095 2415 4135 4035
rect 4995 3640 5035 3645
rect 4995 3610 5000 3640
rect 5030 3610 5035 3640
rect 4995 3345 5035 3610
rect 6060 3640 6100 6530
rect 6120 6505 6160 6510
rect 6120 6475 6125 6505
rect 6155 6475 6160 6505
rect 6120 4945 6160 6475
rect 6120 4915 6125 4945
rect 6155 4915 6160 4945
rect 6120 4910 6160 4915
rect 6425 6450 6465 6455
rect 6425 6420 6430 6450
rect 6460 6420 6465 6450
rect 6425 4845 6465 6420
rect 6425 4815 6430 4845
rect 6460 4815 6465 4845
rect 6425 4810 6465 4815
rect 6060 3610 6065 3640
rect 6095 3610 6100 3640
rect 6060 3605 6100 3610
rect 4995 3315 5000 3345
rect 5030 3315 5035 3345
rect 4995 3310 5035 3315
rect 7095 2520 7135 6585
rect 7150 2710 7190 6650
rect 8315 6505 8355 11580
rect 8370 6560 8410 11635
rect 8370 6530 8375 6560
rect 8405 6530 8410 6560
rect 8370 6525 8410 6530
rect 8315 6475 8320 6505
rect 8350 6475 8355 6505
rect 8315 6470 8355 6475
rect 8435 6450 8475 11690
rect 8505 6615 8545 11745
rect 8505 6585 8510 6615
rect 8540 6585 8545 6615
rect 8505 6580 8545 6585
rect 8435 6420 8440 6450
rect 8470 6420 8475 6450
rect 8435 6415 8475 6420
rect 4095 2385 4100 2415
rect 4130 2385 4135 2415
rect 4095 2380 4135 2385
rect 2440 1790 2480 1830
rect 7610 1790 7650 1830
rect 475 855 480 885
rect 510 855 515 885
rect 475 850 515 855
rect 3985 885 4025 1235
rect 3985 855 3990 885
rect 4020 855 4025 885
rect 3985 850 4025 855
<< via1 >>
rect 3320 11745 3350 11775
rect 2010 11640 2040 11670
rect 1845 10055 1875 10085
rect 480 9305 510 9335
rect 1900 8985 1930 9015
rect 1955 8740 1985 8770
rect 3210 11640 3240 11670
rect 8510 11745 8540 11775
rect 4660 11690 4690 11720
rect 4045 11635 4075 11665
rect 3825 11580 3855 11610
rect 8440 11690 8470 11720
rect 8375 11635 8405 11665
rect 8320 11580 8350 11610
rect 2110 8465 2140 8495
rect 2110 6650 2140 6680
rect 7155 6650 7185 6680
rect 2010 6585 2040 6615
rect 2960 6585 2990 6615
rect 1955 6530 1985 6560
rect 2905 6530 2935 6560
rect 1900 6475 1930 6505
rect 2555 6475 2585 6505
rect 1845 6420 1875 6450
rect 2555 4035 2585 4065
rect 2610 6420 2640 6450
rect 2610 3980 2640 4010
rect 7100 6585 7130 6615
rect 6065 6530 6095 6560
rect 4100 4035 4130 4065
rect 4030 3980 4060 4010
rect 4030 3375 4060 3405
rect 5000 3610 5030 3640
rect 6125 6475 6155 6505
rect 6125 4915 6155 4945
rect 6430 6420 6460 6450
rect 6430 4815 6460 4845
rect 6065 3610 6095 3640
rect 5000 3315 5030 3345
rect 8375 6530 8405 6560
rect 8320 6475 8350 6505
rect 8510 6585 8540 6615
rect 8440 6420 8470 6450
rect 4100 2385 4130 2415
rect 480 855 510 885
rect 3990 855 4020 885
<< metal2 >>
rect 3315 11775 8545 11780
rect 3315 11745 3320 11775
rect 3350 11745 8510 11775
rect 8540 11745 8545 11775
rect 3315 11740 8545 11745
rect 4655 11720 8475 11725
rect 4655 11690 4660 11720
rect 4690 11690 8440 11720
rect 8470 11690 8475 11720
rect 4655 11685 8475 11690
rect 2005 11670 3245 11675
rect 2005 11640 2010 11670
rect 2040 11640 3210 11670
rect 3240 11640 3245 11670
rect 2005 11635 3245 11640
rect 4040 11665 8410 11670
rect 4040 11635 4045 11665
rect 4075 11635 8375 11665
rect 8405 11635 8410 11665
rect 4040 11630 8410 11635
rect 3820 11610 8355 11615
rect 3820 11580 3825 11610
rect 3855 11580 8320 11610
rect 8350 11580 8355 11610
rect 3820 11575 8355 11580
rect 1840 10085 2430 10090
rect 1840 10055 1845 10085
rect 1875 10055 2430 10085
rect 1840 10050 2430 10055
rect 475 9335 2640 9340
rect 475 9305 480 9335
rect 510 9305 2640 9335
rect 475 9300 2640 9305
rect 1895 9015 1935 9020
rect 1895 8985 1900 9015
rect 1930 8985 1935 9015
rect 1895 8980 1935 8985
rect 1950 8770 3220 8775
rect 1950 8740 1955 8770
rect 1985 8740 3220 8770
rect 1950 8735 3220 8740
rect 2105 8495 2145 8500
rect 2105 8465 2110 8495
rect 2140 8465 2145 8495
rect 2105 8460 2145 8465
rect 2105 6680 7190 6685
rect 2105 6650 2110 6680
rect 2140 6650 7155 6680
rect 7185 6650 7190 6680
rect 2105 6645 7190 6650
rect 2005 6615 2995 6620
rect 2005 6585 2010 6615
rect 2040 6585 2960 6615
rect 2990 6585 2995 6615
rect 2005 6580 2995 6585
rect 7095 6615 8545 6620
rect 7095 6585 7100 6615
rect 7130 6585 8510 6615
rect 8540 6585 8545 6615
rect 7095 6580 8545 6585
rect 1950 6560 2940 6565
rect 1950 6530 1955 6560
rect 1985 6530 2905 6560
rect 2935 6530 2940 6560
rect 1950 6525 2940 6530
rect 6060 6560 8410 6565
rect 6060 6530 6065 6560
rect 6095 6530 8375 6560
rect 8405 6530 8410 6560
rect 6060 6525 8410 6530
rect 1895 6505 2590 6510
rect 1895 6475 1900 6505
rect 1930 6475 2555 6505
rect 2585 6475 2590 6505
rect 1895 6470 2590 6475
rect 6120 6505 8355 6510
rect 6120 6475 6125 6505
rect 6155 6475 8320 6505
rect 8350 6475 8355 6505
rect 6120 6470 8355 6475
rect 1840 6450 2645 6455
rect 1840 6420 1845 6450
rect 1875 6420 2610 6450
rect 2640 6420 2645 6450
rect 1840 6415 2645 6420
rect 6425 6450 8475 6455
rect 6425 6420 6430 6450
rect 6460 6420 8440 6450
rect 8470 6420 8475 6450
rect 6425 6415 8475 6420
rect 5795 4945 6160 4950
rect 5795 4915 6125 4945
rect 6155 4915 6160 4945
rect 5795 4910 6160 4915
rect 5750 4845 6465 4850
rect 5750 4840 6430 4845
rect 5745 4820 6430 4840
rect 5750 4815 6430 4820
rect 6460 4815 6465 4845
rect 5750 4810 6465 4815
rect 2550 4065 4135 4070
rect 2550 4035 2555 4065
rect 2585 4035 4100 4065
rect 4130 4035 4135 4065
rect 2550 4030 4135 4035
rect 2605 4010 4065 4015
rect 2605 3980 2610 4010
rect 2640 3980 4030 4010
rect 4060 3980 4065 4010
rect 2605 3975 4065 3980
rect 4995 3640 6100 3645
rect 4995 3610 5000 3640
rect 5030 3610 6065 3640
rect 6095 3610 6100 3640
rect 4995 3605 6100 3610
rect 4025 3405 4105 3410
rect 4025 3375 4030 3405
rect 4060 3375 4105 3405
rect 4025 3370 4105 3375
rect 4860 3345 5035 3350
rect 4860 3315 5000 3345
rect 5030 3315 5035 3345
rect 4860 3310 5035 3315
rect 4095 2415 4965 2420
rect 4095 2385 4100 2415
rect 4130 2385 4965 2415
rect 4095 2380 4965 2385
rect 4090 2280 4105 2310
rect 4090 2060 4105 2100
rect 2440 1790 2480 1830
rect 7610 1790 7650 1830
rect 475 885 4025 890
rect 475 855 480 885
rect 510 855 3990 885
rect 4020 855 4025 885
rect 475 850 4025 855
<< metal3 >>
rect 9840 6880 9890 6885
rect 9840 6840 9845 6880
rect 9885 6840 9890 6880
rect 9840 6835 9890 6840
rect 9845 50 9885 6835
rect 9840 45 9890 50
rect 9840 5 9845 45
rect 9885 5 9890 45
rect 9840 0 9890 5
<< via3 >>
rect 9845 6840 9885 6880
rect 9845 5 9885 45
<< metal4 >>
rect 8145 6880 9890 6885
rect 8145 6840 9845 6880
rect 9885 6840 9890 6880
rect 8145 6835 9890 6840
rect 940 6700 990 6750
rect 975 0 1025 50
rect 9685 45 9890 50
rect 9685 5 9845 45
rect 9885 5 9890 45
rect 9685 0 9890 5
use bgr  bgr_0
timestamp 1751725295
transform -1 0 8030 0 -1 12100
box -200 535 6100 5350
use two_stage_opamp_dummy_magic  two_stage_opamp_dummy_magic_0
timestamp 1751779601
transform 1 0 -51855 0 1 555
box 51855 -555 61545 6195
<< labels >>
flabel metal4 965 6750 965 6750 1 FreeSans 800 0 0 400 VDDA
port 1 n
flabel metal4 1000 0 1000 0 5 FreeSans 800 0 0 -400 GNDA
port 2 s
flabel metal2 4090 2300 4090 2300 7 FreeSans 400 0 -200 0 VIN-
port 6 w
flabel metal2 4090 2080 4090 2080 7 FreeSans 400 0 -200 0 VIN+
port 5 w
flabel metal2 2460 1790 2460 1790 5 FreeSans 400 0 0 -200 VOUT-
port 4 s
flabel metal2 7630 1790 7630 1790 5 FreeSans 400 0 0 -200 VOUT+
port 3 s
<< end >>
