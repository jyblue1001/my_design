magic
tech sky130A
timestamp 1738052034
<< nwell >>
rect 885 150 2005 2565
<< nmos >>
rect 1185 -225 1200 -125
rect 1350 -225 1365 -125
rect 1515 -225 1530 -125
rect 1680 -225 1695 -125
rect 1845 -225 1860 -125
rect 1615 -1420 1665 -420
rect 1815 -1420 1865 -420
<< pmos >>
rect 1115 510 1165 2510
rect 1315 510 1365 2510
rect 1185 175 1200 375
rect 1350 175 1365 375
rect 1515 175 1530 375
rect 1680 175 1695 375
rect 1845 175 1860 375
<< ndiff >>
rect 1135 -140 1185 -125
rect 1135 -210 1150 -140
rect 1170 -210 1185 -140
rect 1135 -225 1185 -210
rect 1200 -140 1250 -125
rect 1200 -210 1215 -140
rect 1235 -210 1250 -140
rect 1200 -225 1250 -210
rect 1300 -140 1350 -125
rect 1300 -210 1315 -140
rect 1335 -210 1350 -140
rect 1300 -225 1350 -210
rect 1365 -140 1415 -125
rect 1365 -210 1380 -140
rect 1400 -210 1415 -140
rect 1365 -225 1415 -210
rect 1465 -140 1515 -125
rect 1465 -210 1480 -140
rect 1500 -210 1515 -140
rect 1465 -225 1515 -210
rect 1530 -140 1580 -125
rect 1530 -210 1545 -140
rect 1565 -210 1580 -140
rect 1530 -225 1580 -210
rect 1630 -140 1680 -125
rect 1630 -210 1645 -140
rect 1665 -210 1680 -140
rect 1630 -225 1680 -210
rect 1695 -140 1745 -125
rect 1695 -210 1710 -140
rect 1730 -210 1745 -140
rect 1695 -225 1745 -210
rect 1795 -140 1845 -125
rect 1795 -210 1810 -140
rect 1830 -210 1845 -140
rect 1795 -225 1845 -210
rect 1860 -140 1910 -125
rect 1860 -210 1875 -140
rect 1895 -210 1910 -140
rect 1860 -225 1910 -210
rect 1565 -435 1615 -420
rect 1565 -1405 1580 -435
rect 1600 -1405 1615 -435
rect 1565 -1420 1615 -1405
rect 1665 -435 1715 -420
rect 1665 -1405 1680 -435
rect 1700 -1405 1715 -435
rect 1665 -1420 1715 -1405
rect 1765 -435 1815 -420
rect 1765 -1405 1780 -435
rect 1800 -1405 1815 -435
rect 1765 -1420 1815 -1405
rect 1865 -435 1915 -420
rect 1865 -1405 1880 -435
rect 1900 -1405 1915 -435
rect 1865 -1420 1915 -1405
<< pdiff >>
rect 1065 2495 1115 2510
rect 1065 525 1080 2495
rect 1100 525 1115 2495
rect 1065 510 1115 525
rect 1165 2495 1215 2510
rect 1165 525 1180 2495
rect 1200 525 1215 2495
rect 1165 510 1215 525
rect 1265 2495 1315 2510
rect 1265 525 1280 2495
rect 1300 525 1315 2495
rect 1265 510 1315 525
rect 1365 2495 1415 2510
rect 1365 525 1380 2495
rect 1400 525 1415 2495
rect 1365 510 1415 525
rect 1135 360 1185 375
rect 1135 190 1150 360
rect 1170 190 1185 360
rect 1135 175 1185 190
rect 1200 360 1250 375
rect 1200 190 1215 360
rect 1235 190 1250 360
rect 1200 175 1250 190
rect 1300 360 1350 375
rect 1300 190 1315 360
rect 1335 190 1350 360
rect 1300 175 1350 190
rect 1365 360 1415 375
rect 1365 190 1380 360
rect 1400 190 1415 360
rect 1365 175 1415 190
rect 1465 360 1515 375
rect 1465 190 1480 360
rect 1500 190 1515 360
rect 1465 175 1515 190
rect 1530 360 1580 375
rect 1530 190 1545 360
rect 1565 190 1580 360
rect 1530 175 1580 190
rect 1630 360 1680 375
rect 1630 190 1645 360
rect 1665 190 1680 360
rect 1630 175 1680 190
rect 1695 360 1745 375
rect 1695 190 1710 360
rect 1730 190 1745 360
rect 1695 175 1745 190
rect 1795 360 1845 375
rect 1795 190 1810 360
rect 1830 190 1845 360
rect 1795 175 1845 190
rect 1860 360 1910 375
rect 1860 190 1875 360
rect 1895 190 1910 360
rect 1860 175 1910 190
<< ndiffc >>
rect 1150 -210 1170 -140
rect 1215 -210 1235 -140
rect 1315 -210 1335 -140
rect 1380 -210 1400 -140
rect 1480 -210 1500 -140
rect 1545 -210 1565 -140
rect 1645 -210 1665 -140
rect 1710 -210 1730 -140
rect 1810 -210 1830 -140
rect 1875 -210 1895 -140
rect 1580 -1405 1600 -435
rect 1680 -1405 1700 -435
rect 1780 -1405 1800 -435
rect 1880 -1405 1900 -435
<< pdiffc >>
rect 1080 525 1100 2495
rect 1180 525 1200 2495
rect 1280 525 1300 2495
rect 1380 525 1400 2495
rect 1150 190 1170 360
rect 1215 190 1235 360
rect 1315 190 1335 360
rect 1380 190 1400 360
rect 1480 190 1500 360
rect 1545 190 1565 360
rect 1645 190 1665 360
rect 1710 190 1730 360
rect 1810 190 1830 360
rect 1875 190 1895 360
<< psubdiff >>
rect 1225 -270 1325 -255
rect 1225 -290 1240 -270
rect 1310 -290 1325 -270
rect 1225 -305 1325 -290
rect 1725 -270 1825 -255
rect 1725 -290 1740 -270
rect 1810 -290 1825 -270
rect 1725 -305 1825 -290
rect 1970 -460 2020 -445
rect 1970 -480 1985 -460
rect 2005 -480 2020 -460
rect 1970 -495 2020 -480
<< nsubdiff >>
rect 1595 485 1795 500
rect 1595 465 1610 485
rect 1780 465 1795 485
rect 1595 450 1795 465
<< psubdiffcont >>
rect 1240 -290 1310 -270
rect 1740 -290 1810 -270
rect 1985 -480 2005 -460
<< nsubdiffcont >>
rect 1610 465 1780 485
<< poly >>
rect 1320 2555 1360 2560
rect 1320 2535 1330 2555
rect 1350 2535 1360 2555
rect 1320 2525 1360 2535
rect 1115 2510 1165 2525
rect 1315 2510 1365 2525
rect 1115 500 1165 510
rect 1315 500 1365 510
rect 1115 475 1365 500
rect 720 435 910 450
rect 895 405 910 435
rect 895 390 1200 405
rect 895 345 910 390
rect 1185 375 1200 390
rect 1350 375 1365 390
rect 1515 375 1530 390
rect 1680 375 1695 390
rect 1845 375 1860 390
rect 615 330 910 345
rect 615 -330 630 330
rect 1185 160 1200 175
rect 1350 85 1365 175
rect 1515 165 1530 175
rect 1680 165 1695 175
rect 1515 160 1695 165
rect 1845 160 1860 175
rect 1480 145 1695 160
rect 1805 150 2105 160
rect 1805 145 2075 150
rect 1480 125 1495 145
rect 1515 125 1530 145
rect 1480 110 1530 125
rect 1805 125 1820 145
rect 1840 125 1860 145
rect 1805 110 1860 125
rect 2065 130 2075 145
rect 2095 130 2105 150
rect 2065 120 2105 130
rect 945 70 1590 85
rect 945 -85 960 70
rect 1540 50 1555 70
rect 1575 50 1590 70
rect 1540 35 1590 50
rect 1350 10 1400 25
rect 1350 -10 1365 10
rect 1385 5 1400 10
rect 1385 -10 1860 5
rect 1350 -25 1400 -10
rect 800 -100 960 -85
rect 1150 -75 1200 -60
rect 1150 -95 1165 -75
rect 1185 -95 1200 -75
rect 1525 -75 1575 -60
rect 1525 -95 1540 -75
rect 1560 -95 1575 -75
rect 1150 -100 1200 -95
rect 1150 -110 1365 -100
rect 1185 -115 1365 -110
rect 1185 -125 1200 -115
rect 1350 -125 1365 -115
rect 1515 -110 1575 -95
rect 1515 -125 1530 -110
rect 1680 -125 1695 -110
rect 1845 -125 1860 -10
rect 2065 -220 2105 -210
rect 1185 -240 1200 -225
rect 1350 -240 1365 -225
rect 1515 -240 1530 -225
rect 1680 -330 1695 -225
rect 1845 -235 1860 -225
rect 2065 -235 2075 -220
rect 1845 -240 2075 -235
rect 2095 -240 2105 -220
rect 1845 -250 2105 -240
rect 615 -345 1695 -330
rect 1615 -420 1665 -405
rect 1815 -420 1865 -405
rect 1615 -1430 1665 -1420
rect 1815 -1430 1865 -1420
rect 1615 -1440 1865 -1430
rect 1615 -1445 1830 -1440
rect 1820 -1460 1830 -1445
rect 1850 -1445 1865 -1440
rect 1850 -1460 1860 -1445
rect 1820 -1470 1860 -1460
<< polycont >>
rect 1330 2535 1350 2555
rect 1495 125 1515 145
rect 1820 125 1840 145
rect 2075 130 2095 150
rect 1555 50 1575 70
rect 1365 -10 1385 10
rect 1165 -95 1185 -75
rect 1540 -95 1560 -75
rect 2075 -240 2095 -220
rect 1830 -1460 1850 -1440
<< xpolycontact >>
rect 2070 545 2105 765
rect 2070 210 2105 430
rect 960 -705 1180 -420
rect 1230 -705 1450 -420
rect 2070 -525 2105 -305
rect 2070 -830 2105 -610
<< xpolyres >>
rect 2070 430 2105 545
rect 1180 -705 1230 -420
rect 2070 -610 2105 -525
<< locali >>
rect 1320 2555 1360 2560
rect 1320 2550 1330 2555
rect 905 2535 1330 2550
rect 1350 2545 1360 2555
rect 1350 2535 1400 2545
rect 905 2530 1400 2535
rect 905 -420 925 2530
rect 1320 2525 1400 2530
rect 1320 2520 1360 2525
rect 1380 2505 1400 2525
rect 1065 2495 1110 2505
rect 1065 525 1080 2495
rect 1100 525 1110 2495
rect 1065 515 1110 525
rect 1170 2495 1215 2505
rect 1170 525 1180 2495
rect 1200 525 1215 2495
rect 1170 515 1215 525
rect 1265 2495 1310 2505
rect 1265 525 1280 2495
rect 1300 525 1310 2495
rect 1265 515 1310 525
rect 1370 2495 1415 2505
rect 1370 525 1380 2495
rect 1400 525 1415 2495
rect 2125 880 2175 890
rect 2125 870 2135 880
rect 2085 850 2135 870
rect 2165 850 2175 880
rect 2085 765 2105 850
rect 2125 840 2175 850
rect 1370 515 1415 525
rect 1080 410 1100 515
rect 1180 485 1200 515
rect 1280 485 1300 515
rect 1600 485 1790 495
rect 1180 465 1610 485
rect 1780 465 1830 485
rect 1080 390 1335 410
rect 1215 370 1235 390
rect 1315 370 1335 390
rect 1545 370 1565 465
rect 1600 455 1790 465
rect 1645 370 1665 455
rect 1810 370 1830 465
rect 1135 360 1180 370
rect 1135 190 1150 360
rect 1170 190 1180 360
rect 1135 180 1180 190
rect 1205 360 1250 370
rect 1205 190 1215 360
rect 1235 190 1250 360
rect 1205 180 1250 190
rect 1300 360 1345 370
rect 1300 190 1315 360
rect 1335 190 1345 360
rect 1300 180 1345 190
rect 1370 360 1415 370
rect 1370 190 1380 360
rect 1400 190 1415 360
rect 1370 180 1415 190
rect 1465 360 1510 370
rect 1465 190 1480 360
rect 1500 190 1510 360
rect 1465 180 1510 190
rect 1535 360 1580 370
rect 1535 190 1545 360
rect 1565 190 1580 360
rect 1535 180 1580 190
rect 1630 360 1675 370
rect 1630 190 1645 360
rect 1665 190 1675 360
rect 1630 180 1675 190
rect 1700 360 1745 370
rect 1700 190 1710 360
rect 1730 190 1745 360
rect 1700 180 1745 190
rect 1795 360 1840 370
rect 1795 190 1810 360
rect 1830 190 1840 360
rect 1795 180 1840 190
rect 1865 360 1910 370
rect 1865 190 1875 360
rect 1895 190 1910 360
rect 1865 180 1910 190
rect 1150 -60 1170 180
rect 1380 25 1400 180
rect 1350 10 1400 25
rect 1350 -10 1365 10
rect 1385 -10 1400 10
rect 1350 -25 1400 -10
rect 1150 -75 1200 -60
rect 1150 -95 1165 -75
rect 1185 -95 1200 -75
rect 1150 -110 1200 -95
rect 1150 -130 1170 -110
rect 1380 -130 1400 -25
rect 1480 160 1500 180
rect 1710 160 1730 180
rect 1480 145 1530 160
rect 1480 125 1495 145
rect 1515 125 1530 145
rect 1480 110 1530 125
rect 1710 145 1855 160
rect 1710 140 1820 145
rect 1480 -130 1500 110
rect 1540 70 1590 85
rect 1540 50 1555 70
rect 1575 50 1590 70
rect 1540 35 1590 50
rect 1540 -60 1560 35
rect 1525 -75 1575 -60
rect 1525 -95 1540 -75
rect 1560 -95 1575 -75
rect 1525 -110 1575 -95
rect 1710 -130 1730 140
rect 1805 125 1820 140
rect 1840 125 1855 145
rect 1805 110 1855 125
rect 1875 30 1895 180
rect 2070 160 2090 210
rect 2065 150 2105 160
rect 2065 130 2075 150
rect 2095 130 2105 150
rect 2065 120 2105 130
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2125 30 2145 70
rect 1875 10 2285 30
rect 2265 -50 2285 10
rect 1875 -70 2285 -50
rect 1875 -130 1895 -70
rect 2125 -125 2145 -70
rect 1135 -140 1180 -130
rect 1135 -210 1150 -140
rect 1170 -210 1180 -140
rect 1135 -220 1180 -210
rect 1205 -140 1250 -130
rect 1205 -210 1215 -140
rect 1235 -210 1250 -140
rect 1205 -220 1250 -210
rect 1230 -260 1250 -220
rect 1300 -140 1345 -130
rect 1300 -210 1315 -140
rect 1335 -210 1345 -140
rect 1300 -220 1345 -210
rect 1370 -140 1415 -130
rect 1370 -210 1380 -140
rect 1400 -210 1415 -140
rect 1370 -220 1415 -210
rect 1465 -140 1510 -130
rect 1465 -210 1480 -140
rect 1500 -210 1510 -140
rect 1465 -220 1510 -210
rect 1535 -140 1580 -130
rect 1535 -210 1545 -140
rect 1565 -210 1580 -140
rect 1535 -220 1580 -210
rect 1630 -140 1675 -130
rect 1630 -210 1645 -140
rect 1665 -210 1675 -140
rect 1630 -220 1675 -210
rect 1700 -140 1745 -130
rect 1700 -210 1710 -140
rect 1730 -210 1745 -140
rect 1700 -220 1745 -210
rect 1795 -140 1840 -130
rect 1795 -210 1810 -140
rect 1830 -210 1840 -140
rect 1795 -220 1840 -210
rect 1865 -140 1910 -130
rect 1865 -210 1875 -140
rect 1895 -210 1910 -140
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 1865 -220 1910 -210
rect 2065 -220 2105 -210
rect 1300 -260 1320 -220
rect 1230 -270 1320 -260
rect 1230 -290 1240 -270
rect 1310 -290 1320 -270
rect 1230 -300 1320 -290
rect 1545 -315 1565 -220
rect 1645 -315 1665 -220
rect 1800 -260 1820 -220
rect 2065 -240 2075 -220
rect 2095 -240 2105 -220
rect 2065 -250 2105 -240
rect 1730 -270 1820 -260
rect 1730 -280 1740 -270
rect 1545 -335 1665 -315
rect 1695 -290 1740 -280
rect 1810 -290 1820 -270
rect 1695 -300 1820 -290
rect 905 -440 960 -420
rect 1580 -425 1600 -335
rect 1695 -425 1715 -300
rect 1780 -425 1800 -300
rect 2085 -305 2105 -250
rect 1430 -1435 1450 -705
rect 1565 -435 1610 -425
rect 1565 -1405 1580 -435
rect 1600 -1405 1610 -435
rect 1565 -1415 1610 -1405
rect 1670 -435 1715 -425
rect 1670 -1405 1680 -435
rect 1700 -1405 1715 -435
rect 1670 -1415 1715 -1405
rect 1765 -435 1810 -425
rect 1765 -1405 1780 -435
rect 1800 -1405 1810 -435
rect 1765 -1415 1810 -1405
rect 1870 -435 1915 -425
rect 1870 -1405 1880 -435
rect 1900 -1405 1915 -435
rect 1975 -460 2015 -450
rect 1975 -480 1985 -460
rect 2005 -480 2015 -460
rect 1975 -490 2015 -480
rect 2085 -905 2105 -830
rect 2125 -905 2175 -895
rect 2085 -925 2135 -905
rect 2125 -935 2135 -925
rect 2165 -935 2175 -905
rect 2125 -945 2175 -935
rect 1870 -1415 1915 -1405
rect 1820 -1435 1860 -1430
rect 1880 -1435 1900 -1415
rect 1430 -1440 1900 -1435
rect 1430 -1455 1830 -1440
rect 1820 -1460 1830 -1455
rect 1850 -1455 1900 -1440
rect 1850 -1460 1860 -1455
rect 1820 -1470 1860 -1460
<< viali >>
rect 1180 525 1200 2495
rect 1280 525 1300 2495
rect 2135 850 2165 880
rect 1610 465 1780 485
rect 1545 190 1565 360
rect 1645 190 1665 360
rect 1810 190 1830 360
rect 2135 80 2170 115
rect 1215 -210 1235 -140
rect 1315 -210 1335 -140
rect 1810 -210 1830 -140
rect 2135 -170 2170 -135
rect 1240 -290 1310 -270
rect 1740 -290 1810 -270
rect 1680 -1405 1700 -435
rect 1780 -1405 1800 -435
rect 2135 -935 2165 -905
<< metal1 >>
rect 855 2495 2025 2565
rect 855 525 1180 2495
rect 1200 525 1280 2495
rect 1300 525 2025 2495
rect 2125 880 2175 890
rect 2125 850 2135 880
rect 2165 850 2175 880
rect 2125 840 2175 850
rect 855 485 2025 525
rect 855 465 1610 485
rect 1780 465 2025 485
rect 855 360 2025 465
rect 855 190 1545 360
rect 1565 190 1645 360
rect 1665 190 1810 360
rect 1830 190 2025 360
rect 855 150 2025 190
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 955 -140 1955 -85
rect 955 -210 1215 -140
rect 1235 -210 1315 -140
rect 1335 -210 1810 -140
rect 1830 -210 1955 -140
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 955 -270 1955 -210
rect 955 -290 1240 -270
rect 1310 -290 1740 -270
rect 1810 -290 1955 -270
rect 955 -435 1955 -290
rect 955 -745 1680 -435
rect 1515 -1405 1680 -745
rect 1700 -1405 1780 -435
rect 1800 -1405 1955 -435
rect 2125 -905 2175 -895
rect 2125 -935 2135 -905
rect 2165 -935 2175 -905
rect 2125 -945 2175 -935
rect 1515 -1420 1955 -1405
rect 1560 -1475 1920 -1420
<< via1 >>
rect 2135 850 2165 880
rect 2135 80 2170 115
rect 2135 -170 2170 -135
rect 2135 -935 2165 -905
<< metal2 >>
rect 2125 880 2175 890
rect 2125 850 2135 880
rect 2165 850 2175 880
rect 2125 840 2175 850
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 2125 -905 2175 -895
rect 2125 -935 2135 -905
rect 2165 -935 2175 -905
rect 2125 -945 2175 -935
<< via2 >>
rect 2135 850 2165 880
rect 2135 80 2170 115
rect 2135 -170 2170 -135
rect 2135 -935 2165 -905
<< metal3 >>
rect 2125 885 2175 890
rect 2125 880 3130 885
rect 2125 850 2135 880
rect 2165 850 3130 880
rect 2125 840 3130 850
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2300 55 3130 840
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 2300 -895 3130 -110
rect 2125 -905 3130 -895
rect 2125 -935 2135 -905
rect 2165 -935 3130 -905
rect 2125 -940 3130 -935
rect 2125 -945 2175 -940
<< via3 >>
rect 2135 80 2170 115
rect 2135 -170 2170 -135
<< mimcap >>
rect 2315 115 3115 870
rect 2315 80 2325 115
rect 2360 80 3115 115
rect 2315 70 3115 80
rect 2315 -135 3115 -125
rect 2315 -170 2325 -135
rect 2360 -170 3115 -135
rect 2315 -925 3115 -170
<< mimcapcontact >>
rect 2325 80 2360 115
rect 2325 -170 2360 -135
<< metal4 >>
rect 2125 115 2365 125
rect 2125 80 2135 115
rect 2170 80 2325 115
rect 2360 80 2365 115
rect 2125 70 2365 80
rect 2125 -135 2365 -125
rect 2125 -170 2135 -135
rect 2170 -170 2325 -135
rect 2360 -170 2365 -135
rect 2125 -180 2365 -170
<< labels >>
flabel metal1 855 795 855 795 7 FreeSans 400 0 0 0 VDDA
flabel metal1 955 -360 955 -360 7 FreeSans 400 0 0 0 GNDA
flabel locali 2285 -20 2285 -20 3 FreeSans 400 0 0 0 VOUT
flabel poly 720 445 720 445 7 FreeSans 400 0 0 0 VIN-
flabel poly 800 -90 800 -90 7 FreeSans 400 0 0 0 VIN+
<< end >>
