* PEX produced on Wed Jul  2 09:26:20 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 a_n8798_9160.t1 a_n7190_9280.t1 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X1 a_14640_5738.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA.t176 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X2 VDDA.t259 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t4 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 bgr_0.NFET_GATE_10uA.t5 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X4 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA.t308 GNDA.t310 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X5 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_0.V_err_gate.t12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDDA.t169 bgr_0.V_mir1.t12 bgr_0.V_mir1.t13 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X13 GNDA.t63 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X14 GNDA.t41 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X15 two_stage_opamp_dummy_magic_0.X.t19 GNDA.t311 GNDA.t313 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X16 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VDDA.t206 two_stage_opamp_dummy_magic_0.X.t26 VOUT-.t2 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X20 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_0.Y.t25 VDDA.t381 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X21 bgr_0.V_p_2.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 bgr_0.V_mir2.t2 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X22 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 GNDA.t227 GNDA.t315 bgr_0.Vbe2.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X24 VDDA.t454 bgr_0.V_TOP.t14 bgr_0.START_UP.t3 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X25 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5750_2946.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X26 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VDDA.t139 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X30 bgr_0.V_p_1.t7 bgr_0.Vin+.t6 bgr_0.1st_Vout_1.t2 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X31 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.VD3.t23 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X32 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VDDA.t456 bgr_0.V_TOP.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X36 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 GNDA.t175 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X38 GNDA.t225 GNDA.t314 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X39 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VDDA.t217 two_stage_opamp_dummy_magic_0.Vb3.t8 two_stage_opamp_dummy_magic_0.VD3.t19 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X42 VDDA.t121 VDDA.t119 two_stage_opamp_dummy_magic_0.V_err_gate.t1 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X43 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 two_stage_opamp_dummy_magic_0.Y.t20 GNDA.t319 GNDA.t321 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X46 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD1.t9 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X47 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X50 VOUT-.t3 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t208 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X51 bgr_0.V_TOP.t16 VDDA.t458 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 two_stage_opamp_dummy_magic_0.V_err_p.t4 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 VDDA.t428 bgr_0.1st_Vout_2.t13 bgr_0.PFET_GATE_10uA.t9 VDDA.t427 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X54 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 two_stage_opamp_dummy_magic_0.VD1.t17 VIN-.t0 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X56 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X60 VDDA.t460 bgr_0.V_TOP.t17 bgr_0.Vin+.t3 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X61 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 GNDA.t151 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X64 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 two_stage_opamp_dummy_magic_0.Vb2.t8 bgr_0.NFET_GATE_10uA.t7 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X67 GNDA.t46 bgr_0.START_UP_NFET1.t1 bgr_0.START_UP_NFET1.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X68 two_stage_opamp_dummy_magic_0.VD1.t21 VIN-.t1 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA.t332 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X69 VDDA.t145 two_stage_opamp_dummy_magic_0.Vb3.t9 two_stage_opamp_dummy_magic_0.VD3.t7 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X70 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.VD3.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X72 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 VDDA.t116 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X73 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 GNDA.t342 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 VOUT+.t18 GNDA.t341 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X75 GNDA.t14 two_stage_opamp_dummy_magic_0.X.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X76 GNDA.t89 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X77 VDDA.t426 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t8 VDDA.t425 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X78 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 GNDA.t318 GNDA.t316 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X81 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 two_stage_opamp_dummy_magic_0.Vb2.t7 bgr_0.NFET_GATE_10uA.t8 GNDA.t100 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X85 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT+.t15 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t294 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X87 GNDA.t307 GNDA.t305 GNDA.t307 GNDA.t306 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X88 GNDA.t304 GNDA.t302 two_stage_opamp_dummy_magic_0.VD1.t19 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X89 VDDA.t359 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t358 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X90 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 bgr_0.PFET_GATE_10uA.t10 VDDA.t284 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X92 GNDA.t301 GNDA.t299 VOUT+.t17 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X93 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_0.X.t29 VDDA.t151 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X94 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X96 GNDA.t298 GNDA.t296 two_stage_opamp_dummy_magic_0.X.t18 GNDA.t297 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X97 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t147 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X98 VOUT-.t7 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X99 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 bgr_0.1st_Vout_2.t10 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t10 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X106 a_14640_5738.t0 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X107 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 bgr_0.1st_Vout_2.t5 bgr_0.V_mir2.t18 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X111 VDDA.t115 VDDA.t113 two_stage_opamp_dummy_magic_0.VD3.t1 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X112 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 bgr_0.V_TOP.t18 VDDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 GNDA.t18 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X115 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 bgr_0.NFET_GATE_10uA.t9 GNDA.t102 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X118 VDDA.t262 two_stage_opamp_dummy_magic_0.X.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X119 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X120 bgr_0.V_TOP.t19 VDDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 bgr_0.V_mir1.t11 bgr_0.V_mir1.t10 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X122 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 bgr_0.PFET_GATE_10uA.t11 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X124 GNDA.t295 GNDA.t293 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X125 GNDA.t292 GNDA.t290 two_stage_opamp_dummy_magic_0.Y.t19 GNDA.t291 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X126 GNDA.t134 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X127 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 GNDA.t150 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X129 GNDA.t135 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t321 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X130 two_stage_opamp_dummy_magic_0.X.t17 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X131 bgr_0.Vin+.t2 bgr_0.V_TOP.t20 VDDA.t300 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X132 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 two_stage_opamp_dummy_magic_0.V_p.t36 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X135 bgr_0.V_mir2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 bgr_0.V_p_2.t5 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X136 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 VOUT-.t4 a_5750_2946.t1 GNDA.t54 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X138 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 bgr_0.V_TOP.t21 VDDA.t301 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 bgr_0.1st_Vout_1.t0 bgr_0.Vin+.t7 bgr_0.V_p_1.t6 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X142 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t287 GNDA.t289 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X143 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT+.t14 two_stage_opamp_dummy_magic_0.Y.t29 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X145 two_stage_opamp_dummy_magic_0.V_p.t4 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA.t31 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X146 two_stage_opamp_dummy_magic_0.V_p.t27 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X147 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VDDA.t437 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t10 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X150 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X151 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t12 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X153 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 a_n9700_9790.t1 GNDA.t86 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X157 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT+.t16 GNDA.t284 GNDA.t286 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X159 bgr_0.V_TOP.t22 VDDA.t445 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 bgr_0.PFET_GATE_10uA.t7 bgr_0.1st_Vout_2.t16 VDDA.t424 VDDA.t423 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X161 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 two_stage_opamp_dummy_magic_0.VD2.t20 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t23 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X164 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT-.t10 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X167 VOUT-.t11 two_stage_opamp_dummy_magic_0.X.t35 VDDA.t313 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X168 VDDA.t339 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X169 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VOUT-.t8 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X172 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t4 GNDA.t21 sky130_fd_pr__res_high_po_1p41 l=1.41
X174 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 GNDA.t20 two_stage_opamp_dummy_magic_0.Y.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X176 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.Vb3.t11 VDDA.t416 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X178 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 VDDA.t414 bgr_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X180 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X181 two_stage_opamp_dummy_magic_0.err_amp_out.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X182 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA.t281 GNDA.t283 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X183 VDDA.t263 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X184 GNDA.t227 GNDA.t280 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X185 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP.t4 bgr_0.START_UP.t5 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X187 bgr_0.1st_Vout_2.t6 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t1 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X188 two_stage_opamp_dummy_magic_0.VD1.t8 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.Y.t13 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X189 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 bgr_0.PFET_GATE_10uA.t6 bgr_0.1st_Vout_2.t18 VDDA.t422 VDDA.t421 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X193 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 bgr_0.PFET_GATE_10uA.t14 VDDA.t370 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X194 VDDA.t112 VDDA.t110 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X195 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 GNDA.t5 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X199 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X200 GNDA.t84 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X201 a_5230_5758.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t17 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X202 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VDDA.t223 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X204 VDDA.t441 bgr_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X205 two_stage_opamp_dummy_magic_0.Vb2.t6 bgr_0.NFET_GATE_10uA.t10 GNDA.t346 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X206 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 two_stage_opamp_dummy_magic_0.V_p.t7 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X212 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_0.V_p.t40 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA.t353 GNDA.t352 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X214 VDDA.t195 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD4.t11 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X215 VOUT+.t13 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t324 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X216 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 two_stage_opamp_dummy_magic_0.Y.t18 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X218 two_stage_opamp_dummy_magic_0.V_p.t17 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t11 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X219 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t277 GNDA.t279 GNDA.t278 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X220 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 bgr_0.V_CUR_REF_REG.t1 bgr_0.PFET_GATE_10uA.t16 VDDA.t133 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X222 bgr_0.PFET_GATE_10uA.t1 VDDA.t107 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X223 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X224 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 two_stage_opamp_dummy_magic_0.VD2.t18 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t20 GNDA.t331 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X229 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 bgr_0.V_p_2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 bgr_0.V_mir2.t0 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X231 a_14520_5738.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t67 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X232 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 bgr_0.cap_res1.t0 bgr_0.V_TOP.t9 GNDA.t44 sky130_fd_pr__res_high_po_0p35 l=2.05
X234 VOUT-.t12 two_stage_opamp_dummy_magic_0.X.t38 VDDA.t318 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X235 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VDDA.t200 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X237 VDDA.t468 bgr_0.V_mir1.t6 bgr_0.V_mir1.t7 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X238 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 two_stage_opamp_dummy_magic_0.V_err_p.t0 VDDA.t104 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X244 GNDA.t157 two_stage_opamp_dummy_magic_0.Y.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X245 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 two_stage_opamp_dummy_magic_0.Y.t12 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD4.t29 two_stage_opamp_dummy_magic_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X248 GNDA.t351 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 VDDA.t463 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X249 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t131 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X252 VDDA.t153 bgr_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X253 VDDA.t272 bgr_0.1st_Vout_1.t20 bgr_0.V_TOP.t8 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X254 bgr_0.V_TOP.t23 VDDA.t446 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X256 VDDA.t319 two_stage_opamp_dummy_magic_0.X.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X257 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X259 VDDA.t308 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X260 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 VDDA.t164 bgr_0.V_TOP.t24 bgr_0.Vin-.t3 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X262 VDDA.t380 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t379 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X263 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 two_stage_opamp_dummy_magic_0.VD1.t7 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t3 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X265 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VDDA.t149 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t11 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X267 VDDA.t187 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X268 GNDA.t56 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X269 bgr_0.V_p_2.t8 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t8 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X270 GNDA.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X271 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t15 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X272 GNDA.t199 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 VOUT-.t14 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X273 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X274 two_stage_opamp_dummy_magic_0.V_p.t16 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X275 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 GNDA.t349 two_stage_opamp_dummy_magic_0.err_amp_out.t12 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA.t348 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X277 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 VDDA.t103 VDDA.t101 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X281 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 VDDA.t439 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X283 VDDA.t185 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD3.t13 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X284 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 bgr_0.NFET_GATE_10uA.t12 GNDA.t82 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X285 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VDDA.t100 VDDA.t98 two_stage_opamp_dummy_magic_0.Vb1.t3 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X287 bgr_0.1st_Vout_1.t9 bgr_0.V_mir1.t18 VDDA.t286 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X288 VOUT+.t12 two_stage_opamp_dummy_magic_0.Y.t36 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X289 two_stage_opamp_dummy_magic_0.V_p.t15 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X290 two_stage_opamp_dummy_magic_0.V_p.t3 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X291 VOUT+.t11 two_stage_opamp_dummy_magic_0.Y.t37 VDDA.t448 VDDA.t447 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X292 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 GNDA.t87 a_n9700_9790.t0 GNDA.t86 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X296 bgr_0.V_p_2.t0 VDDA.t469 GNDA.t215 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X297 VDDA.t255 bgr_0.V_mir2.t14 bgr_0.V_mir2.t15 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X298 bgr_0.V_TOP.t6 VDDA.t470 GNDA.t216 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X299 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 GNDA.t238 GNDA.t276 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X303 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t7 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X304 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t3 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X305 bgr_0.NFET_GATE_10uA.t4 GNDA.t273 GNDA.t275 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X306 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X307 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VDDA.t302 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X310 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 bgr_0.START_UP.t2 bgr_0.V_TOP.t25 VDDA.t166 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X314 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_0.VD4.t1 VDDA.t95 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X318 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X319 GNDA.t219 VDDA.t92 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X320 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA.t181 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X322 bgr_0.V_p_2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 bgr_0.V_mir2.t1 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X323 VDDA.t253 bgr_0.V_mir2.t8 bgr_0.V_mir2.t9 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X324 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VDDA.t309 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X328 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 two_stage_opamp_dummy_magic_0.VD1.t6 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.Y.t6 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X331 VDDA.t135 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 a_5350_5758.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t115 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X333 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 GNDA.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_p_mir.t2 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X335 bgr_0.V_TOP.t12 bgr_0.START_UP.t6 bgr_0.Vin-.t6 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X336 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X337 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t292 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X338 GNDA.t1 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X339 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 GNDA.t197 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X343 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_0.V_err_p.t18 VDDA.t289 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X344 two_stage_opamp_dummy_magic_0.V_p.t38 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t333 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X345 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 bgr_0.V_p_1.t2 bgr_0.Vin-.t8 bgr_0.V_mir1.t1 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X348 bgr_0.V_TOP.t26 VDDA.t231 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.Vb3.t14 VDDA.t334 VDDA.t333 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X350 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X351 GNDA.t227 GNDA.t226 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X352 VDDA.t88 VDDA.t85 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X353 VOUT+.t1 VDDA.t89 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X354 two_stage_opamp_dummy_magic_0.V_p.t35 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t327 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X355 two_stage_opamp_dummy_magic_0.V_p.t5 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X356 GNDA.t225 GNDA.t224 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X357 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t23 VDDA.t420 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X358 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 bgr_0.cap_res2.t0 bgr_0.PFET_GATE_10uA.t3 GNDA.t44 sky130_fd_pr__res_high_po_0p35 l=2.05
X361 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 bgr_0.V_mir2.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 bgr_0.V_p_2.t2 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X363 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VDDA.t84 VDDA.t82 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X365 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t10 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X366 two_stage_opamp_dummy_magic_0.V_err_gate.t5 bgr_0.NFET_GATE_10uA.t14 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X367 two_stage_opamp_dummy_magic_0.VD2.t1 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t3 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X368 bgr_0.V_mir1.t3 bgr_0.V_mir1.t2 VDDA.t432 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X369 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VDDA.t282 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X372 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VDDA.t279 two_stage_opamp_dummy_magic_0.Y.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X374 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VDDA.t251 bgr_0.V_mir2.t19 bgr_0.1st_Vout_2.t2 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X376 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t2 GNDA.t19 sky130_fd_pr__res_high_po_1p41 l=1.41
X378 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Y.t9 two_stage_opamp_dummy_magic_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X379 bgr_0.V_TOP.t27 VDDA.t232 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 VDDA.t79 VDDA.t81 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X381 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 two_stage_opamp_dummy_magic_0.V_err_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t137 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X383 bgr_0.V_mir1.t14 bgr_0.Vin-.t9 bgr_0.V_p_1.t8 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X384 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X386 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t78 VDDA.t76 bgr_0.V_CUR_REF_REG.t0 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X388 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA.t138 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X389 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VDDA.t191 bgr_0.PFET_GATE_10uA.t20 bgr_0.NFET_GATE_10uA.t1 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X391 bgr_0.V_TOP.t28 VDDA.t347 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 VDDA.t349 bgr_0.V_TOP.t29 bgr_0.Vin-.t2 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X394 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.Vb3.t15 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X395 two_stage_opamp_dummy_magic_0.VD1.t5 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t11 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X396 VDDA.t219 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X397 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X398 two_stage_opamp_dummy_magic_0.VD1.t4 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.Y.t17 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X399 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 GNDA.t272 GNDA.t269 GNDA.t271 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X403 two_stage_opamp_dummy_magic_0.err_amp_out.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X404 GNDA.t37 VDDA.t73 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X405 VDDA.t173 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0.64 ps=3.6 w=3.2 l=0.2
X406 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 two_stage_opamp_dummy_magic_0.V_p.t14 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t10 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X408 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 VDDA.t221 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t8 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X413 VDDA.t72 VDDA.t70 GNDA.t335 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X414 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 GNDA.t65 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X417 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t249 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X418 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 GNDA.t71 bgr_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X420 bgr_0.V_TOP.t30 VDDA.t340 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+.t3 a_14240_2946.t0 GNDA.t61 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X422 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VDDA.t342 bgr_0.V_TOP.t31 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X426 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t181 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X428 VDDA.t69 VDDA.t67 bgr_0.V_TOP.t5 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X429 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X433 VDDA.t66 VDDA.t64 bgr_0.PFET_GATE_10uA.t0 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X434 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X435 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_0.X.t42 GNDA.t62 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X436 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT-.t1 VDDA.t58 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X438 bgr_0.1st_Vout_1.t4 bgr_0.Vin+.t8 bgr_0.V_p_1.t5 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X439 VDDA.t412 GNDA.t266 GNDA.t268 GNDA.t267 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X440 VDDA.t355 two_stage_opamp_dummy_magic_0.Vb3.t17 two_stage_opamp_dummy_magic_0.VD4.t8 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X441 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 GNDA.t188 bgr_0.NFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X443 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 bgr_0.V_mir2.t5 bgr_0.V_mir2.t4 VDDA.t247 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X447 VDDA.t63 VDDA.t61 VOUT+.t0 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X448 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X450 bgr_0.V_TOP.t4 VDDA.t55 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X451 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA.t264 GNDA.t265 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X455 VOUT+.t4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t75 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X456 GNDA.t227 GNDA.t254 bgr_0.Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X457 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 a_5350_5758.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA.t112 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X460 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 GNDA.t225 GNDA.t253 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X462 two_stage_opamp_dummy_magic_0.V_err_gate.t9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X463 VDDA.t4 bgr_0.1st_Vout_1.t24 bgr_0.V_TOP.t0 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X464 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VDDA.t330 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X466 VDDA.t226 two_stage_opamp_dummy_magic_0.X.t43 VOUT-.t5 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X467 bgr_0.V_mir1.t15 bgr_0.Vin-.t10 bgr_0.V_p_1.t9 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X468 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 VDDA.t52 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X469 bgr_0.V_TOP.t32 VDDA.t385 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VDDA.t234 two_stage_opamp_dummy_magic_0.Vb3.t18 two_stage_opamp_dummy_magic_0.VD4.t7 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X471 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 two_stage_opamp_dummy_magic_0.Y.t1 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X475 two_stage_opamp_dummy_magic_0.V_p.t33 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t325 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X476 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t430 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X477 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VOUT+.t5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X479 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X480 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 two_stage_opamp_dummy_magic_0.Y.t41 GNDA.t340 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X483 bgr_0.V_TOP.t33 VDDA.t386 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 bgr_0.Vin-.t1 bgr_0.V_TOP.t34 VDDA.t363 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X486 GNDA.t190 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X487 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VDDA.t6 bgr_0.1st_Vout_1.t25 bgr_0.V_TOP.t1 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X489 VDDA.t143 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.VD4.t6 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X490 VDDA.t51 VDDA.t49 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X491 VDDA.t450 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 VDDA.t449 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X492 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 GNDA.t113 VDDA.t471 bgr_0.PFET_GATE_10uA.t2 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X494 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 two_stage_opamp_dummy_magic_0.V_p.t26 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA.t173 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X496 two_stage_opamp_dummy_magic_0.V_p.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA.t160 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X497 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_0.X.t44 GNDA.t126 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X498 two_stage_opamp_dummy_magic_0.VD2.t0 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.X.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X499 bgr_0.1st_Vout_2.t0 bgr_0.V_mir2.t20 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X500 VDDA.t48 VDDA.t46 GNDA.t11 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X501 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 GNDA.t114 VDDA.t472 bgr_0.V_p_1.t0 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X504 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 two_stage_opamp_dummy_magic_0.VD1.t16 VIN-.t6 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X506 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 bgr_0.V_p_1.t4 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t1 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X512 GNDA.t263 GNDA.t261 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X513 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 bgr_0.V_TOP.t35 VDDA.t364 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t22 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X516 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 GNDA.t203 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X518 VDDA.t462 two_stage_opamp_dummy_magic_0.Y.t42 VOUT+.t10 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X519 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 bgr_0.V_TOP.t36 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X520 two_stage_opamp_dummy_magic_0.VD1.t18 VIN-.t7 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X521 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VDDA.t131 bgr_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X526 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VDDA.t336 two_stage_opamp_dummy_magic_0.Vb3.t21 two_stage_opamp_dummy_magic_0.VD4.t5 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X529 VDDA.t411 GNDA.t258 GNDA.t260 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X530 two_stage_opamp_dummy_magic_0.Y.t0 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X531 VDDA.t243 bgr_0.V_mir2.t6 bgr_0.V_mir2.t7 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X532 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X533 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VDDA.t307 two_stage_opamp_dummy_magic_0.X.t45 VOUT-.t9 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X535 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 VDDA.t45 VDDA.t43 VOUT-.t0 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X537 GNDA.t257 GNDA.t255 VDDA.t410 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X538 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 bgr_0.V_TOP.t3 VDDA.t40 VDDA.t42 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X541 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VDDA.t241 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t1 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X545 VDDA.t288 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t8 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X546 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_2946.t1 GNDA.t350 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X549 bgr_0.Vin-.t0 bgr_0.V_TOP.t37 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X550 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 two_stage_opamp_dummy_magic_0.Y.t43 GNDA.t330 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X551 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 bgr_0.PFET_GATE_10uA.t23 VDDA.t374 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X554 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 GNDA.t252 GNDA.t250 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X556 two_stage_opamp_dummy_magic_0.X.t16 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X557 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 two_stage_opamp_dummy_magic_0.X.t46 VDDA.t397 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X558 bgr_0.V_TOP.t11 bgr_0.1st_Vout_1.t27 VDDA.t304 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X559 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 two_stage_opamp_dummy_magic_0.Y.t4 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X562 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t9 GNDA.t343 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X563 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VDDA.t352 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X566 bgr_0.V_p_1.t10 bgr_0.Vin-.t11 bgr_0.V_mir1.t16 GNDA.t354 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X567 GNDA.t73 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 VOUT-.t6 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X568 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 two_stage_opamp_dummy_magic_0.Y.t16 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.VD1.t3 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X570 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.Vb3.t22 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X572 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 two_stage_opamp_dummy_magic_0.VD2.t3 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.X.t8 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X574 two_stage_opamp_dummy_magic_0.V_p.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA.t170 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X575 VDDA.t39 VDDA.t37 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X576 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_0.X.t47 GNDA.t210 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X577 VDDA.t175 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD3.t12 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X578 GNDA.t50 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 VOUT+.t2 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X579 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t34 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X581 GNDA.t184 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X582 GNDA.t162 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X583 VDDA.t316 two_stage_opamp_dummy_magic_0.Y.t44 VOUT+.t9 VDDA.t315 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X584 a_5230_5758.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA.t124 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X585 GNDA.t249 GNDA.t247 VOUT-.t18 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X586 two_stage_opamp_dummy_magic_0.VD2.t12 VIN+.t7 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X587 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 bgr_0.V_TOP.t7 bgr_0.1st_Vout_1.t28 VDDA.t210 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X589 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 VDDA.t372 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X591 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 two_stage_opamp_dummy_magic_0.V_err_gate.t4 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X594 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 VDDA.t31 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=1.28 ps=7.2 w=3.2 l=0.2
X596 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X597 bgr_0.V_p_1.t3 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t3 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X598 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X601 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VDDA.t395 two_stage_opamp_dummy_magic_0.X.t48 VOUT-.t15 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X604 VDDA.t298 two_stage_opamp_dummy_magic_0.Vb3.t24 two_stage_opamp_dummy_magic_0.VD3.t30 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X605 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 two_stage_opamp_dummy_magic_0.Y.t45 VDDA.t167 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X606 VDDA.t1 bgr_0.V_TOP.t38 bgr_0.Vin+.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X607 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X608 bgr_0.V_TOP.t39 VDDA.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t46 GNDA.t142 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X611 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t132 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X614 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 bgr_0.V_TOP.t10 bgr_0.1st_Vout_1.t30 VDDA.t281 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X616 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t408 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X617 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 bgr_0.V_TOP.t40 VDDA.t360 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 bgr_0.PFET_GATE_10uA.t26 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X620 GNDA.t140 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X621 GNDA.t186 bgr_0.NFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X622 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t396 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X623 GNDA.t246 GNDA.t244 VDDA.t409 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X624 two_stage_opamp_dummy_magic_0.Vb1.t2 VDDA.t28 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X625 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 VDDA.t418 bgr_0.1st_Vout_2.t31 bgr_0.PFET_GATE_10uA.t4 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X628 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X629 VDDA.t27 VDDA.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X630 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t332 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X633 two_stage_opamp_dummy_magic_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t20 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X634 two_stage_opamp_dummy_magic_0.V_p.t24 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA.t165 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X635 two_stage_opamp_dummy_magic_0.V_err_p.t21 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 VDDA.t403 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X636 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_0.X.t50 GNDA.t220 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X637 two_stage_opamp_dummy_magic_0.VD2.t11 VIN+.t8 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X638 bgr_0.V_TOP.t41 VDDA.t361 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 GNDA.t243 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X640 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X641 GNDA.t240 GNDA.t239 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X642 VDDA.t443 bgr_0.V_TOP.t42 bgr_0.START_UP.t1 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X643 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 bgr_0.1st_Vout_1.t7 bgr_0.V_mir1.t20 VDDA.t212 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X645 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 bgr_0.PFET_GATE_10uA.t27 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X648 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 bgr_0.PFET_GATE_10uA.t28 VDDA.t275 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X650 two_stage_opamp_dummy_magic_0.VD3.t0 VDDA.t22 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X651 GNDA.t119 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X652 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 two_stage_opamp_dummy_magic_0.Vb1.t4 bgr_0.PFET_GATE_10uA.t29 VDDA.t156 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X654 VDDA.t199 two_stage_opamp_dummy_magic_0.Y.t48 VOUT+.t8 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X655 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 two_stage_opamp_dummy_magic_0.VD2.t14 VIN+.t9 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X658 a_n8798_9040.t1 a_n7190_9400.t0 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X659 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t402 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X660 VDDA.t278 two_stage_opamp_dummy_magic_0.Y.t49 VOUT+.t7 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X661 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 GNDA.t59 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X664 a_14520_5738.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t136 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X665 a_n8798_9040.t0 bgr_0.Vin+.t4 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X666 GNDA.t238 GNDA.t237 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X667 bgr_0.V_mir2.t13 bgr_0.V_mir2.t12 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X668 GNDA.t96 a_n9760_9260.t0 GNDA.t95 sky130_fd_pr__res_xhigh_po_0p35 l=6
X669 VOUT-.t17 GNDA.t234 GNDA.t236 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X670 two_stage_opamp_dummy_magic_0.V_err_gate.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X671 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA.t355 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X673 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_0.V_p.t0 two_stage_opamp_dummy_magic_0.Vb1.t0 two_stage_opamp_dummy_magic_0.Vb1.t1 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X675 VDDA.t406 two_stage_opamp_dummy_magic_0.X.t51 VOUT-.t16 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X676 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_0.Y.t50 VDDA.t265 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X677 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 bgr_0.1st_Vout_1.t6 bgr_0.V_mir1.t21 VDDA.t214 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X679 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VOUT-.t13 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA.t179 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X684 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VDDA.t177 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X686 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 two_stage_opamp_dummy_magic_0.Y.t51 GNDA.t338 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X687 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.Y.t24 two_stage_opamp_dummy_magic_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X689 GNDA.t213 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X690 two_stage_opamp_dummy_magic_0.Vb2.t2 two_stage_opamp_dummy_magic_0.Vb2.t1 VDDA.t376 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X691 bgr_0.1st_Vout_2.t7 bgr_0.V_CUR_REF_REG.t7 bgr_0.V_p_2.t7 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X692 bgr_0.V_TOP.t43 VDDA.t444 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 bgr_0.V_mir1.t0 bgr_0.Vin-.t12 bgr_0.V_p_1.t1 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X695 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t392 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X696 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t1 GNDA.t347 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X698 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 two_stage_opamp_dummy_magic_0.V_err_p.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t179 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X700 bgr_0.Vin+.t0 bgr_0.V_TOP.t44 VDDA.t229 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X701 bgr_0.V_TOP.t45 VDDA.t230 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.Vb3.t27 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X703 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 bgr_0.Vin-.t5 bgr_0.START_UP.t7 bgr_0.V_TOP.t13 VDDA.t465 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X705 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X706 two_stage_opamp_dummy_magic_0.Vb3.t2 bgr_0.NFET_GATE_10uA.t22 GNDA.t145 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X707 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 two_stage_opamp_dummy_magic_0.V_p.t21 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X709 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t7 VDDA.t267 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X710 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA.t231 GNDA.t233 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X711 two_stage_opamp_dummy_magic_0.V_p_mir.t3 VIN-.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X712 two_stage_opamp_dummy_magic_0.VD1.t12 VIN-.t9 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X713 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 bgr_0.V_TOP.t46 VDDA.t344 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 GNDA.t344 a_n7190_9400.t1 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X719 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VDDA.t435 bgr_0.V_mir1.t22 bgr_0.1st_Vout_1.t5 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X722 VDDA.t366 two_stage_opamp_dummy_magic_0.Y.t52 VOUT+.t6 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X723 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 a_n8798_9160.t0 bgr_0.Vin-.t4 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X725 two_stage_opamp_dummy_magic_0.VD1.t13 VIN-.t10 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X726 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 GNDA.t104 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X728 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X729 bgr_0.V_CUR_REF_REG.t2 a_n9760_9260.t1 GNDA.t95 sky130_fd_pr__res_xhigh_po_0p35 l=6
X730 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 bgr_0.V_TOP.t47 VDDA.t346 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X733 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 bgr_0.V_TOP.t48 VDDA.t382 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 bgr_0.START_UP.t0 bgr_0.V_TOP.t49 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X737 two_stage_opamp_dummy_magic_0.V_err_gate.t0 VDDA.t19 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X738 two_stage_opamp_dummy_magic_0.V_err_gate.t13 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X739 GNDA.t167 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.t3 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X740 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.Vb3.t28 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X742 two_stage_opamp_dummy_magic_0.X.t15 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X743 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.VD3.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X744 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_0.Y.t53 VDDA.t276 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X746 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 two_stage_opamp_dummy_magic_0.Y.t54 VDDA.t452 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X749 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 bgr_0.1st_Vout_2.t3 bgr_0.V_mir2.t22 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X753 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VDDA.t18 VDDA.t16 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0 ps=0 w=3.2 l=0.2
X755 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 VDDA.t326 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t5 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X760 bgr_0.Vbe2.t0 bgr_0.Vin+.t5 GNDA.t123 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X761 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 GNDA.t111 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X763 GNDA.t230 GNDA.t228 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t229 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X764 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 bgr_0.NFET_GATE_10uA.t0 VDDA.t13 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X767 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 two_stage_opamp_dummy_magic_0.X.t53 VDDA.t393 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X769 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD1.t0 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X772 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t328 VDDA.t327 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X773 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.VD3.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X774 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 two_stage_opamp_dummy_magic_0.V_p_mir.t1 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X779 VDDA.t12 VDDA.t10 bgr_0.V_TOP.t2 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X780 two_stage_opamp_dummy_magic_0.V_err_p.t19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t6 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X781 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t205 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X782 two_stage_opamp_dummy_magic_0.Vb3.t1 bgr_0.NFET_GATE_10uA.t23 GNDA.t147 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X783 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA.t221 GNDA.t223 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X785 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 GNDA.t122 a_n7190_9280.t0 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X787 two_stage_opamp_dummy_magic_0.VD2.t17 VIN+.t10 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X788 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X789 VDDA.t9 VDDA.t7 two_stage_opamp_dummy_magic_0.VD4.t0 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X790 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 a_n8798_9160.t0 a_n8798_9160.t1 258.591
R1 a_n7190_9280.t0 a_n7190_9280.t1 376.99
R2 GNDA.n856 GNDA.n779 299369
R3 GNDA.n1012 GNDA.n994 68623.1
R4 GNDA.n856 GNDA.n855 64900
R5 GNDA.n1009 GNDA.n994 56607.7
R6 GNDA.n990 GNDA.n949 41223.8
R7 GNDA.n1013 GNDA.n993 35482.9
R8 GNDA.n1011 GNDA.n995 34650
R9 GNDA.n1014 GNDA.n927 32661.5
R10 GNDA.n992 GNDA.n927 32661.5
R11 GNDA.n853 GNDA.n778 30676.6
R12 GNDA.n1850 GNDA.n1849 29091.6
R13 GNDA.n1175 GNDA.n868 28430.8
R14 GNDA.n1016 GNDA.n990 28430.8
R15 GNDA.n1015 GNDA.n1013 28372.4
R16 GNDA.n1012 GNDA.n1011 27818.3
R17 GNDA.n1849 GNDA.n779 26648.4
R18 GNDA.n1013 GNDA.n927 19630.8
R19 GNDA.n1110 GNDA.n927 19630.8
R20 GNDA.n1850 GNDA.n778 18723.2
R21 GNDA.n994 GNDA.n991 18063.2
R22 GNDA.n855 GNDA.n854 17370.4
R23 GNDA.n1008 GNDA.n991 15462.2
R24 GNDA.n1015 GNDA.n1014 14773.1
R25 GNDA.n993 GNDA.n992 14449.6
R26 GNDA.n784 GNDA.n780 12361.8
R27 GNDA.n783 GNDA.n780 12312.5
R28 GNDA.n1010 GNDA.n1009 12184.6
R29 GNDA.n2468 GNDA.n2467 12175.2
R30 GNDA.n1847 GNDA.n784 11918.5
R31 GNDA.n1847 GNDA.n783 11869.2
R32 GNDA.n778 GNDA.n777 11338.5
R33 GNDA.n854 GNDA.n779 11169.2
R34 GNDA.n1010 GNDA.n1007 10968.3
R35 GNDA.n1098 GNDA.n882 10835
R36 GNDA.n1149 GNDA.n882 10835
R37 GNDA.n1098 GNDA.n883 10835
R38 GNDA.n1149 GNDA.n883 10835
R39 GNDA.n854 GNDA.n853 10831.8
R40 GNDA.n1849 GNDA.n1848 10371.4
R41 GNDA.n1151 GNDA.n868 10371.4
R42 GNDA.n1013 GNDA.n1012 9476.92
R43 GNDA.n929 GNDA.n928 9308.25
R44 GNDA.n934 GNDA.n928 9308.25
R45 GNDA.n1109 GNDA.n929 9308.25
R46 GNDA.n1109 GNDA.n934 9308.25
R47 GNDA.n1137 GNDA.n892 9259
R48 GNDA.n1137 GNDA.n1136 8914.25
R49 GNDA.n1009 GNDA.n1008 8800
R50 GNDA.n1011 GNDA.n1010 8695.24
R51 GNDA.n1853 GNDA.n773 8175.5
R52 GNDA.n893 GNDA.n892 8175.5
R53 GNDA.n1853 GNDA.n774 8126.25
R54 GNDA.n823 GNDA.n816 7880
R55 GNDA.n1838 GNDA.n816 7880
R56 GNDA.n1195 GNDA.n1186 7880
R57 GNDA.n1195 GNDA.n1188 7880
R58 GNDA.n823 GNDA.n818 7830.75
R59 GNDA.n1838 GNDA.n818 7830.75
R60 GNDA.n1186 GNDA.n850 7830.75
R61 GNDA.n1188 GNDA.n850 7830.75
R62 GNDA.n1136 GNDA.n893 7830.75
R63 GNDA.n1857 GNDA.n773 7732.25
R64 GNDA.n880 GNDA.n874 7732.25
R65 GNDA.n1161 GNDA.n874 7732.25
R66 GNDA.n1160 GNDA.n880 7732.25
R67 GNDA.n1161 GNDA.n1160 7732.25
R68 GNDA.n1054 GNDA.n966 7732.25
R69 GNDA.n1054 GNDA.n967 7732.25
R70 GNDA.n1056 GNDA.n966 7732.25
R71 GNDA.n1056 GNDA.n967 7732.25
R72 GNDA.n1857 GNDA.n774 7683
R73 GNDA.n1166 GNDA.n857 7338.25
R74 GNDA.n1033 GNDA.n983 7338.25
R75 GNDA.n1182 GNDA.n857 7289
R76 GNDA.n853 GNDA.n852 7287.5
R77 GNDA.n1028 GNDA.n983 7092
R78 GNDA.n1940 GNDA.n1939 6917.5
R79 GNDA.n1879 GNDA.n1872 6845.75
R80 GNDA.n1879 GNDA.n1873 6845.75
R81 GNDA.n1872 GNDA.n648 6796.5
R82 GNDA.n1873 GNDA.n648 6796.5
R83 GNDA.n1934 GNDA.n466 6698
R84 GNDA.n1938 GNDA.n466 6698
R85 GNDA.n1934 GNDA.n467 6648.75
R86 GNDA.n1938 GNDA.n467 6648.75
R87 GNDA.n1157 GNDA.n865 6057.75
R88 GNDA.n1177 GNDA.n865 6057.75
R89 GNDA.n1157 GNDA.n866 6057.75
R90 GNDA.n1177 GNDA.n866 6057.75
R91 GNDA.n1044 GNDA.n974 6057.75
R92 GNDA.n1047 GNDA.n1044 6057.75
R93 GNDA.n974 GNDA.n971 6057.75
R94 GNDA.n1047 GNDA.n971 6057.75
R95 GNDA.n855 GNDA.n852 5525.52
R96 GNDA.n1771 GNDA.n1656 5502.84
R97 GNDA.n1851 GNDA.n777 5325.97
R98 GNDA.n1166 GNDA.n858 5319
R99 GNDA.n1033 GNDA.n984 5319
R100 GNDA.n1182 GNDA.n858 5269.75
R101 GNDA.n1028 GNDA.n984 5269.75
R102 GNDA.n1174 GNDA.n869 5171.25
R103 GNDA.n1040 GNDA.n978 5171.25
R104 GNDA.n1170 GNDA.n869 5122
R105 GNDA.n1036 GNDA.n978 5122
R106 GNDA.n1896 GNDA.n465 5090.53
R107 GNDA.n1222 GNDA.n820 4974.25
R108 GNDA.n1226 GNDA.n820 4974.25
R109 GNDA.n1174 GNDA.n870 4944.7
R110 GNDA.n1040 GNDA.n979 4944.7
R111 GNDA.n956 GNDA.n926 4925
R112 GNDA.n1112 GNDA.n926 4925
R113 GNDA.n1170 GNDA.n870 4895.45
R114 GNDA.n1036 GNDA.n979 4895.45
R115 GNDA.n956 GNDA.n920 4728
R116 GNDA.n1112 GNDA.n920 4728
R117 GNDA.n1016 GNDA.n1015 4727.03
R118 GNDA.n1779 GNDA.n1615 4678.75
R119 GNDA.n1783 GNDA.n1615 4629.5
R120 GNDA.n1779 GNDA.n1616 4629.5
R121 GNDA.n1923 GNDA.n481 4580.25
R122 GNDA.n1923 GNDA.n482 4580.25
R123 GNDA.n1783 GNDA.n1616 4580.25
R124 GNDA.n1919 GNDA.n479 4580.25
R125 GNDA.n488 GNDA.n479 4580.25
R126 GNDA.n1222 GNDA.n821 4531
R127 GNDA.n1226 GNDA.n821 4531
R128 GNDA.n842 GNDA.n781 4531
R129 GNDA.n1219 GNDA.n781 4531
R130 GNDA.n842 GNDA.n782 4531
R131 GNDA.n1219 GNDA.n782 4531
R132 GNDA.n1894 GNDA.n481 4481.75
R133 GNDA.n1894 GNDA.n482 4481.75
R134 GNDA.n1919 GNDA.n486 4481.75
R135 GNDA.n488 GNDA.n486 4481.75
R136 GNDA.n1851 GNDA.n1850 3770.78
R137 GNDA.n1095 GNDA.n950 3595.25
R138 GNDA.n961 GNDA.n950 3595.25
R139 GNDA.n931 GNDA.n894 3349
R140 GNDA.n1133 GNDA.n894 3299.75
R141 GNDA.n1095 GNDA.n951 3250.5
R142 GNDA.n961 GNDA.n951 3250.5
R143 GNDA.n931 GNDA.n895 3250.5
R144 GNDA.n1133 GNDA.n895 3201.25
R145 GNDA.n1008 GNDA.n1007 3174.4
R146 GNDA.n1006 GNDA.n995 3148.62
R147 GNDA.n1939 GNDA.n465 2978.29
R148 GNDA.n1014 GNDA.n990 2933.33
R149 GNDA.n992 GNDA.n868 2933.33
R150 GNDA.n852 GNDA.n777 2569.8
R151 GNDA.n1205 GNDA.n847 2371.15
R152 GNDA.n1208 GNDA.n847 2371.15
R153 GNDA.n1185 GNDA.n1184 2341.03
R154 GNDA.n1007 GNDA.n1006 2331.19
R155 GNDA.n1004 GNDA.n997 2326.02
R156 GNDA.n998 GNDA.n997 2326.02
R157 GNDA.n1024 GNDA.n988 2326.02
R158 GNDA.n1017 GNDA.n988 2326.02
R159 GNDA.n1027 GNDA.n1025 2324.65
R160 GNDA.n1184 GNDA.n856 2237.35
R161 GNDA.n835 GNDA.n834 2142.38
R162 GNDA.n1202 GNDA.n846 2142.38
R163 GNDA.n834 GNDA.n827 1846.88
R164 GNDA.n1212 GNDA.n846 1846.88
R165 GNDA.n1184 GNDA.n851 1707.72
R166 GNDA.n995 GNDA.n993 1564
R167 GNDA.n1184 GNDA.n1183 1469.8
R168 GNDA.n848 GNDA.n847 1301.55
R169 GNDA.n640 GNDA.n495 1214.72
R170 GNDA.n640 GNDA.n507 1214.72
R171 GNDA.n598 GNDA.n507 1214.72
R172 GNDA.n606 GNDA.n598 1214.72
R173 GNDA.n606 GNDA.n605 1214.72
R174 GNDA.n621 GNDA.n589 1214.72
R175 GNDA.n621 GNDA.n585 1214.72
R176 GNDA.n628 GNDA.n585 1214.72
R177 GNDA.n628 GNDA.n410 1214.72
R178 GNDA.n2132 GNDA.n410 1214.72
R179 GNDA.n1001 GNDA.n997 1114.8
R180 GNDA.n1020 GNDA.n988 1114.8
R181 GNDA.n834 GNDA.n833 991.841
R182 GNDA.n1197 GNDA.n846 991.841
R183 GNDA.n1967 GNDA.n1966 949.682
R184 GNDA.n2498 GNDA.t227 949.682
R185 GNDA.n1771 GNDA.t225 875.452
R186 GNDA.n589 GNDA.t225 823.313
R187 GNDA.n1845 GNDA.n1844 803.201
R188 GNDA.n1844 GNDA.n785 800
R189 GNDA.n1846 GNDA.n1845 774.4
R190 GNDA.n1846 GNDA.n785 771.201
R191 GNDA.n862 GNDA.t258 734.418
R192 GNDA.n1153 GNDA.t244 734.418
R193 GNDA.n972 GNDA.t266 734.418
R194 GNDA.n975 GNDA.t255 734.418
R195 GNDA.n1099 GNDA.n886 704
R196 GNDA.n1148 GNDA.n886 697.601
R197 GNDA.n1090 GNDA.t231 682.201
R198 GNDA.n1140 GNDA.t269 682.201
R199 GNDA.n2515 GNDA.n2514 669.307
R200 GNDA.n953 GNDA.t241 666.134
R201 GNDA.n1087 GNDA.t305 666.134
R202 GNDA.n1837 GNDA.n1836 628.034
R203 GNDA.n1016 GNDA.n991 624.324
R204 GNDA.n1982 GNDA.n1967 623.755
R205 GNDA.n2492 GNDA.t227 623.755
R206 GNDA.n1003 GNDA.n999 617.601
R207 GNDA.n1023 GNDA.n989 617.601
R208 GNDA.n1138 GNDA.n891 601.601
R209 GNDA.n1108 GNDA.n945 598.4
R210 GNDA.n1108 GNDA.n935 598.4
R211 GNDA.n1831 GNDA.n1235 588.271
R212 GNDA.n1564 GNDA.n1343 588.271
R213 GNDA.n2495 GNDA.n15 585
R214 GNDA.n205 GNDA.n14 585
R215 GNDA.n2373 GNDA.n2369 585
R216 GNDA.n2374 GNDA.n204 585
R217 GNDA.n2375 GNDA.n203 585
R218 GNDA.n2364 GNDA.n200 585
R219 GNDA.n2380 GNDA.n199 585
R220 GNDA.n2381 GNDA.n198 585
R221 GNDA.n2382 GNDA.n197 585
R222 GNDA.n2361 GNDA.n195 585
R223 GNDA.n2360 GNDA.n192 585
R224 GNDA.n2390 GNDA.n2389 585
R225 GNDA.n2393 GNDA.n2392 585
R226 GNDA.n2392 GNDA.n46 585
R227 GNDA.n2496 GNDA.n2495 585
R228 GNDA.n2371 GNDA.n14 585
R229 GNDA.n2373 GNDA.n2372 585
R230 GNDA.n2374 GNDA.n202 585
R231 GNDA.n2376 GNDA.n2375 585
R232 GNDA.n2378 GNDA.n200 585
R233 GNDA.n2380 GNDA.n2379 585
R234 GNDA.n2381 GNDA.n196 585
R235 GNDA.n2383 GNDA.n2382 585
R236 GNDA.n2385 GNDA.n195 585
R237 GNDA.n2386 GNDA.n192 585
R238 GNDA.n2389 GNDA.n2388 585
R239 GNDA.n2128 GNDA.n2127 585
R240 GNDA.n2015 GNDA.n2009 585
R241 GNDA.n2123 GNDA.n2122 585
R242 GNDA.n2017 GNDA.n2014 585
R243 GNDA.n2045 GNDA.n2044 585
R244 GNDA.n2049 GNDA.n2048 585
R245 GNDA.n2047 GNDA.n2038 585
R246 GNDA.n2056 GNDA.n2055 585
R247 GNDA.n2058 GNDA.n2057 585
R248 GNDA.n2063 GNDA.n2060 585
R249 GNDA.n2065 GNDA.n2064 585
R250 GNDA.n2061 GNDA.n193 585
R251 GNDA.n2325 GNDA.n69 585
R252 GNDA.n2319 GNDA.n364 585
R253 GNDA.n2321 GNDA.n2320 585
R254 GNDA.n2318 GNDA.n369 585
R255 GNDA.n2317 GNDA.n2316 585
R256 GNDA.n2315 GNDA.n2314 585
R257 GNDA.n2313 GNDA.n2312 585
R258 GNDA.n2311 GNDA.n2310 585
R259 GNDA.n2309 GNDA.n2308 585
R260 GNDA.n2307 GNDA.n2306 585
R261 GNDA.n2305 GNDA.n2304 585
R262 GNDA.n2303 GNDA.n2302 585
R263 GNDA.n2269 GNDA.n2268 585
R264 GNDA.n2266 GNDA.n388 585
R265 GNDA.n2159 GNDA.n2158 585
R266 GNDA.n2187 GNDA.n2186 585
R267 GNDA.n2189 GNDA.n2188 585
R268 GNDA.n2194 GNDA.n2193 585
R269 GNDA.n2196 GNDA.n2195 585
R270 GNDA.n2201 GNDA.n2200 585
R271 GNDA.n2203 GNDA.n2202 585
R272 GNDA.n2257 GNDA.n2205 585
R273 GNDA.n2259 GNDA.n2258 585
R274 GNDA.n2255 GNDA.n346 585
R275 GNDA.n2133 GNDA.n409 585
R276 GNDA.n2133 GNDA.n2132 585
R277 GNDA.n625 GNDA.n408 585
R278 GNDA.n410 GNDA.n408 585
R279 GNDA.n627 GNDA.n626 585
R280 GNDA.n628 GNDA.n627 585
R281 GNDA.n624 GNDA.n586 585
R282 GNDA.n586 GNDA.n585 585
R283 GNDA.n623 GNDA.n622 585
R284 GNDA.n622 GNDA.n621 585
R285 GNDA.n588 GNDA.n587 585
R286 GNDA.n589 GNDA.n588 585
R287 GNDA.n604 GNDA.n603 585
R288 GNDA.n605 GNDA.n604 585
R289 GNDA.n602 GNDA.n599 585
R290 GNDA.n606 GNDA.n599 585
R291 GNDA.n601 GNDA.n600 585
R292 GNDA.n600 GNDA.n598 585
R293 GNDA.n506 GNDA.n505 585
R294 GNDA.n507 GNDA.n506 585
R295 GNDA.n642 GNDA.n641 585
R296 GNDA.n641 GNDA.n640 585
R297 GNDA.n643 GNDA.n498 585
R298 GNDA.n498 GNDA.n495 585
R299 GNDA.n508 GNDA.n493 585
R300 GNDA.n508 GNDA.n495 585
R301 GNDA.n639 GNDA.n638 585
R302 GNDA.n640 GNDA.n639 585
R303 GNDA.n511 GNDA.n509 585
R304 GNDA.n509 GNDA.n507 585
R305 GNDA.n596 GNDA.n595 585
R306 GNDA.n598 GNDA.n596 585
R307 GNDA.n608 GNDA.n607 585
R308 GNDA.n607 GNDA.n606 585
R309 GNDA.n597 GNDA.n591 585
R310 GNDA.n605 GNDA.n597 585
R311 GNDA.n613 GNDA.n590 585
R312 GNDA.n590 GNDA.n589 585
R313 GNDA.n620 GNDA.n619 585
R314 GNDA.n621 GNDA.n620 585
R315 GNDA.n615 GNDA.n584 585
R316 GNDA.n585 GNDA.n584 585
R317 GNDA.n630 GNDA.n629 585
R318 GNDA.n629 GNDA.n628 585
R319 GNDA.n631 GNDA.n411 585
R320 GNDA.n411 GNDA.n410 585
R321 GNDA.n2131 GNDA.n2130 585
R322 GNDA.n2132 GNDA.n2131 585
R323 GNDA.n1527 GNDA.n1342 585
R324 GNDA.n1525 GNDA.n1524 585
R325 GNDA.n1346 GNDA.n1344 585
R326 GNDA.n1427 GNDA.n1425 585
R327 GNDA.n1434 GNDA.n1433 585
R328 GNDA.n1436 GNDA.n1423 585
R329 GNDA.n1439 GNDA.n1438 585
R330 GNDA.n1421 GNDA.n1420 585
R331 GNDA.n1446 GNDA.n1445 585
R332 GNDA.n1448 GNDA.n1368 585
R333 GNDA.n1517 GNDA.n1516 585
R334 GNDA.n1514 GNDA.n1513 585
R335 GNDA.n504 GNDA.n497 585
R336 GNDA.n497 GNDA.n496 585
R337 GNDA.n503 GNDA.n502 585
R338 GNDA.n502 GNDA.n501 585
R339 GNDA.n500 GNDA.n499 585
R340 GNDA.n500 GNDA.n480 585
R341 GNDA.n477 GNDA.n476 585
R342 GNDA.n1925 GNDA.n477 585
R343 GNDA.n1928 GNDA.n1927 585
R344 GNDA.n1927 GNDA.n1926 585
R345 GNDA.n1929 GNDA.n474 585
R346 GNDA.n478 GNDA.n474 585
R347 GNDA.n1931 GNDA.n1930 585
R348 GNDA.n1932 GNDA.n1931 585
R349 GNDA.n475 GNDA.n473 585
R350 GNDA.n473 GNDA.n472 585
R351 GNDA.n1869 GNDA.n1868 585
R352 GNDA.n1870 GNDA.n1869 585
R353 GNDA.n1867 GNDA.n650 585
R354 GNDA.n650 GNDA.n649 585
R355 GNDA.n1860 GNDA.n1859 585
R356 GNDA.n1862 GNDA.n1861 585
R357 GNDA.n1865 GNDA.n1864 585
R358 GNDA.n1864 GNDA.n1863 585
R359 GNDA.n645 GNDA.n644 585
R360 GNDA.n646 GNDA.n645 585
R361 GNDA.n1898 GNDA.n1897 585
R362 GNDA.n1897 GNDA.n1896 585
R363 GNDA.n1900 GNDA.n1899 585
R364 GNDA.n1901 GNDA.n1900 585
R365 GNDA.n1893 GNDA.n1892 585
R366 GNDA.n1902 GNDA.n1893 585
R367 GNDA.n1905 GNDA.n1904 585
R368 GNDA.n1904 GNDA.n1903 585
R369 GNDA.n1906 GNDA.n1891 585
R370 GNDA.n1891 GNDA.n1890 585
R371 GNDA.n1908 GNDA.n1907 585
R372 GNDA.n1909 GNDA.n1908 585
R373 GNDA.n1889 GNDA.n1888 585
R374 GNDA.n1910 GNDA.n1889 585
R375 GNDA.n1913 GNDA.n1912 585
R376 GNDA.n1912 GNDA.n1911 585
R377 GNDA.n1914 GNDA.n491 585
R378 GNDA.n491 GNDA.n489 585
R379 GNDA.n1916 GNDA.n1915 585
R380 GNDA.n1917 GNDA.n1916 585
R381 GNDA.n1881 GNDA.n490 585
R382 GNDA.n1883 GNDA.n1882 585
R383 GNDA.n1886 GNDA.n1885 585
R384 GNDA.n1885 GNDA.n1884 585
R385 GNDA.n2134 GNDA.n371 585
R386 GNDA.n425 GNDA.n406 585
R387 GNDA.n2139 GNDA.n405 585
R388 GNDA.n2140 GNDA.n404 585
R389 GNDA.n2141 GNDA.n403 585
R390 GNDA.n422 GNDA.n400 585
R391 GNDA.n2146 GNDA.n399 585
R392 GNDA.n2147 GNDA.n398 585
R393 GNDA.n2148 GNDA.n397 585
R394 GNDA.n419 GNDA.n395 585
R395 GNDA.n418 GNDA.n392 585
R396 GNDA.n2155 GNDA.n391 585
R397 GNDA.n380 GNDA.n374 585
R398 GNDA.n2300 GNDA.n374 585
R399 GNDA.n2301 GNDA.n372 585
R400 GNDA.n2301 GNDA.n2300 585
R401 GNDA.n1985 GNDA.n451 585
R402 GNDA.n449 GNDA.n446 585
R403 GNDA.n1990 GNDA.n445 585
R404 GNDA.n1991 GNDA.n443 585
R405 GNDA.n1992 GNDA.n442 585
R406 GNDA.n440 GNDA.n437 585
R407 GNDA.n1997 GNDA.n436 585
R408 GNDA.n1998 GNDA.n434 585
R409 GNDA.n1999 GNDA.n433 585
R410 GNDA.n429 GNDA.n428 585
R411 GNDA.n2005 GNDA.n2004 585
R412 GNDA.n2007 GNDA.n415 585
R413 GNDA.n414 GNDA.n373 585
R414 GNDA.n2300 GNDA.n373 585
R415 GNDA.n2135 GNDA.n2134 585
R416 GNDA.n2137 GNDA.n406 585
R417 GNDA.n2139 GNDA.n2138 585
R418 GNDA.n2140 GNDA.n402 585
R419 GNDA.n2142 GNDA.n2141 585
R420 GNDA.n2144 GNDA.n400 585
R421 GNDA.n2146 GNDA.n2145 585
R422 GNDA.n2147 GNDA.n396 585
R423 GNDA.n2149 GNDA.n2148 585
R424 GNDA.n2151 GNDA.n395 585
R425 GNDA.n2152 GNDA.n392 585
R426 GNDA.n2155 GNDA.n2154 585
R427 GNDA.n1986 GNDA.n1985 585
R428 GNDA.n1988 GNDA.n446 585
R429 GNDA.n1990 GNDA.n1989 585
R430 GNDA.n1991 GNDA.n439 585
R431 GNDA.n1993 GNDA.n1992 585
R432 GNDA.n1995 GNDA.n437 585
R433 GNDA.n1997 GNDA.n1996 585
R434 GNDA.n1998 GNDA.n431 585
R435 GNDA.n2000 GNDA.n1999 585
R436 GNDA.n2002 GNDA.n429 585
R437 GNDA.n2004 GNDA.n2003 585
R438 GNDA.n415 GNDA.n412 585
R439 GNDA.n771 GNDA.n652 585
R440 GNDA.n663 GNDA.n653 585
R441 GNDA.n767 GNDA.n766 585
R442 GNDA.n660 GNDA.n658 585
R443 GNDA.n690 GNDA.n689 585
R444 GNDA.n694 GNDA.n693 585
R445 GNDA.n692 GNDA.n683 585
R446 GNDA.n701 GNDA.n700 585
R447 GNDA.n703 GNDA.n702 585
R448 GNDA.n707 GNDA.n705 585
R449 GNDA.n709 GNDA.n708 585
R450 GNDA.n393 GNDA.n390 585
R451 GNDA.n1810 GNDA.n379 585
R452 GNDA.n1804 GNDA.n1606 585
R453 GNDA.n1806 GNDA.n1805 585
R454 GNDA.n1803 GNDA.n1611 585
R455 GNDA.n1802 GNDA.n1801 585
R456 GNDA.n1800 GNDA.n1799 585
R457 GNDA.n1798 GNDA.n1797 585
R458 GNDA.n1796 GNDA.n1795 585
R459 GNDA.n1794 GNDA.n1793 585
R460 GNDA.n1792 GNDA.n1791 585
R461 GNDA.n1790 GNDA.n1789 585
R462 GNDA.n1788 GNDA.n1787 585
R463 GNDA.n1630 GNDA.n1613 585
R464 GNDA.n1614 GNDA.n1613 585
R465 GNDA.n1632 GNDA.n1631 585
R466 GNDA.n1633 GNDA.n1632 585
R467 GNDA.n1636 GNDA.n1635 585
R468 GNDA.n1635 GNDA.n1634 585
R469 GNDA.n1637 GNDA.n1629 585
R470 GNDA.n1629 GNDA.n1628 585
R471 GNDA.n1639 GNDA.n1638 585
R472 GNDA.n1640 GNDA.n1639 585
R473 GNDA.n1625 GNDA.n1624 585
R474 GNDA.n1641 GNDA.n1625 585
R475 GNDA.n1644 GNDA.n1643 585
R476 GNDA.n1643 GNDA.n1642 585
R477 GNDA.n1645 GNDA.n1623 585
R478 GNDA.n1627 GNDA.n1623 585
R479 GNDA.n1647 GNDA.n1646 585
R480 GNDA.n1648 GNDA.n1647 585
R481 GNDA.n1622 GNDA.n1620 585
R482 GNDA.n1649 GNDA.n1622 585
R483 GNDA.n1786 GNDA.n1612 585
R484 GNDA.n1786 GNDA.n1785 585
R485 GNDA.n1651 GNDA.n1650 585
R486 GNDA.n1621 GNDA.n1618 585
R487 GNDA.n1776 GNDA.n1775 585
R488 GNDA.n1777 GNDA.n1776 585
R489 GNDA.n1774 GNDA.n1773 585
R490 GNDA.n1658 GNDA.n1655 585
R491 GNDA.n1769 GNDA.n1768 585
R492 GNDA.n1660 GNDA.n1657 585
R493 GNDA.n1691 GNDA.n1690 585
R494 GNDA.n1692 GNDA.n1691 585
R495 GNDA.n1695 GNDA.n1694 585
R496 GNDA.n1694 GNDA.n1693 585
R497 GNDA.n1696 GNDA.n1683 585
R498 GNDA.n1683 GNDA.n1682 585
R499 GNDA.n1705 GNDA.n1704 585
R500 GNDA.n1706 GNDA.n1705 585
R501 GNDA.n1685 GNDA.n1681 585
R502 GNDA.n1707 GNDA.n1681 585
R503 GNDA.n1710 GNDA.n1709 585
R504 GNDA.n1709 GNDA.n1708 585
R505 GNDA.n1711 GNDA.n1231 585
R506 GNDA.n1231 GNDA.n1230 585
R507 GNDA.n1833 GNDA.n1832 585
R508 GNDA.n1834 GNDA.n1833 585
R509 GNDA.n1579 GNDA.n1234 585
R510 GNDA.n1577 GNDA.n1576 585
R511 GNDA.n1238 GNDA.n1236 585
R512 GNDA.n1319 GNDA.n1317 585
R513 GNDA.n1326 GNDA.n1325 585
R514 GNDA.n1328 GNDA.n1315 585
R515 GNDA.n1331 GNDA.n1330 585
R516 GNDA.n1313 GNDA.n1312 585
R517 GNDA.n1338 GNDA.n1337 585
R518 GNDA.n1340 GNDA.n1260 585
R519 GNDA.n1569 GNDA.n1568 585
R520 GNDA.n1566 GNDA.n1565 585
R521 GNDA.n378 GNDA.n376 585
R522 GNDA.n1604 GNDA.n1603 585
R523 GNDA.n1815 GNDA.n1601 585
R524 GNDA.n1816 GNDA.n1599 585
R525 GNDA.n1817 GNDA.n1598 585
R526 GNDA.n1596 GNDA.n1593 585
R527 GNDA.n1822 GNDA.n1592 585
R528 GNDA.n1823 GNDA.n1590 585
R529 GNDA.n1824 GNDA.n1589 585
R530 GNDA.n1587 GNDA.n1584 585
R531 GNDA.n1829 GNDA.n1583 585
R532 GNDA.n1830 GNDA.n1581 585
R533 GNDA.n1235 GNDA.n1229 585
R534 GNDA.n2299 GNDA.n2298 585
R535 GNDA.n2300 GNDA.n2299 585
R536 GNDA.n1811 GNDA.n378 585
R537 GNDA.n1813 GNDA.n1604 585
R538 GNDA.n1815 GNDA.n1814 585
R539 GNDA.n1816 GNDA.n1595 585
R540 GNDA.n1818 GNDA.n1817 585
R541 GNDA.n1820 GNDA.n1593 585
R542 GNDA.n1822 GNDA.n1821 585
R543 GNDA.n1823 GNDA.n1586 585
R544 GNDA.n1825 GNDA.n1824 585
R545 GNDA.n1827 GNDA.n1584 585
R546 GNDA.n1829 GNDA.n1828 585
R547 GNDA.n1830 GNDA.n1232 585
R548 GNDA.n2355 GNDA.n2354 585
R549 GNDA.n2279 GNDA.n223 585
R550 GNDA.n2281 GNDA.n2280 585
R551 GNDA.n2282 GNDA.n2277 585
R552 GNDA.n2284 GNDA.n2283 585
R553 GNDA.n2286 GNDA.n2275 585
R554 GNDA.n2288 GNDA.n2287 585
R555 GNDA.n2289 GNDA.n2274 585
R556 GNDA.n2291 GNDA.n2290 585
R557 GNDA.n2293 GNDA.n381 585
R558 GNDA.n2295 GNDA.n2294 585
R559 GNDA.n2296 GNDA.n377 585
R560 GNDA.n1489 GNDA.n1461 585
R561 GNDA.n1487 GNDA.n1486 585
R562 GNDA.n1485 GNDA.n1462 585
R563 GNDA.n1484 GNDA.n1483 585
R564 GNDA.n1481 GNDA.n1463 585
R565 GNDA.n1479 GNDA.n1478 585
R566 GNDA.n1477 GNDA.n1464 585
R567 GNDA.n1476 GNDA.n1475 585
R568 GNDA.n1473 GNDA.n1465 585
R569 GNDA.n1471 GNDA.n1470 585
R570 GNDA.n1469 GNDA.n1468 585
R571 GNDA.n1466 GNDA.n224 585
R572 GNDA.n2358 GNDA.n2357 585
R573 GNDA.n219 GNDA.n217 585
R574 GNDA.n1548 GNDA.n1544 585
R575 GNDA.n1549 GNDA.n1543 585
R576 GNDA.n1550 GNDA.n1542 585
R577 GNDA.n1539 GNDA.n1538 585
R578 GNDA.n1555 GNDA.n1537 585
R579 GNDA.n1556 GNDA.n1536 585
R580 GNDA.n1557 GNDA.n1535 585
R581 GNDA.n1532 GNDA.n1531 585
R582 GNDA.n1562 GNDA.n1530 585
R583 GNDA.n1563 GNDA.n1529 585
R584 GNDA.n1343 GNDA.n1229 585
R585 GNDA.n220 GNDA.n218 585
R586 GNDA.n218 GNDA.n46 585
R587 GNDA.n2357 GNDA.n2356 585
R588 GNDA.n1546 GNDA.n219 585
R589 GNDA.n1548 GNDA.n1547 585
R590 GNDA.n1549 GNDA.n1541 585
R591 GNDA.n1551 GNDA.n1550 585
R592 GNDA.n1553 GNDA.n1539 585
R593 GNDA.n1555 GNDA.n1554 585
R594 GNDA.n1556 GNDA.n1534 585
R595 GNDA.n1558 GNDA.n1557 585
R596 GNDA.n1560 GNDA.n1532 585
R597 GNDA.n1562 GNDA.n1561 585
R598 GNDA.n1563 GNDA.n1341 585
R599 GNDA.n2327 GNDA.n2326 585
R600 GNDA.n362 GNDA.n361 585
R601 GNDA.n2332 GNDA.n360 585
R602 GNDA.n2333 GNDA.n359 585
R603 GNDA.n2334 GNDA.n358 585
R604 GNDA.n355 GNDA.n354 585
R605 GNDA.n2339 GNDA.n353 585
R606 GNDA.n2340 GNDA.n352 585
R607 GNDA.n2341 GNDA.n351 585
R608 GNDA.n349 GNDA.n348 585
R609 GNDA.n347 GNDA.n345 585
R610 GNDA.n2349 GNDA.n2348 585
R611 GNDA.n2352 GNDA.n2351 585
R612 GNDA.n2351 GNDA.n46 585
R613 GNDA.n70 GNDA.n68 585
R614 GNDA.n68 GNDA.n46 585
R615 GNDA.n2328 GNDA.n2327 585
R616 GNDA.n2330 GNDA.n362 585
R617 GNDA.n2332 GNDA.n2331 585
R618 GNDA.n2333 GNDA.n357 585
R619 GNDA.n2335 GNDA.n2334 585
R620 GNDA.n2337 GNDA.n355 585
R621 GNDA.n2339 GNDA.n2338 585
R622 GNDA.n2340 GNDA.n350 585
R623 GNDA.n2342 GNDA.n2341 585
R624 GNDA.n2344 GNDA.n349 585
R625 GNDA.n2345 GNDA.n345 585
R626 GNDA.n2348 GNDA.n2347 585
R627 GNDA.n344 GNDA.n343 585
R628 GNDA.n341 GNDA.n340 585
R629 GNDA.n339 GNDA.n338 585
R630 GNDA.n257 GNDA.n230 585
R631 GNDA.n261 GNDA.n260 585
R632 GNDA.n263 GNDA.n256 585
R633 GNDA.n266 GNDA.n265 585
R634 GNDA.n252 GNDA.n251 585
R635 GNDA.n276 GNDA.n275 585
R636 GNDA.n278 GNDA.n249 585
R637 GNDA.n281 GNDA.n280 585
R638 GNDA.n52 GNDA.n50 585
R639 GNDA.n2418 GNDA.n2417 585
R640 GNDA.n2416 GNDA.n2415 585
R641 GNDA.n2414 GNDA.n63 585
R642 GNDA.n2412 GNDA.n2411 585
R643 GNDA.n2410 GNDA.n64 585
R644 GNDA.n2409 GNDA.n2408 585
R645 GNDA.n2406 GNDA.n65 585
R646 GNDA.n2404 GNDA.n2403 585
R647 GNDA.n2402 GNDA.n66 585
R648 GNDA.n2401 GNDA.n2400 585
R649 GNDA.n2398 GNDA.n67 585
R650 GNDA.n2396 GNDA.n2395 585
R651 GNDA.n190 GNDA.n189 585
R652 GNDA.n187 GNDA.n186 585
R653 GNDA.n185 GNDA.n184 585
R654 GNDA.n103 GNDA.n76 585
R655 GNDA.n107 GNDA.n106 585
R656 GNDA.n109 GNDA.n102 585
R657 GNDA.n112 GNDA.n111 585
R658 GNDA.n98 GNDA.n97 585
R659 GNDA.n122 GNDA.n121 585
R660 GNDA.n124 GNDA.n95 585
R661 GNDA.n127 GNDA.n126 585
R662 GNDA.n41 GNDA.n40 585
R663 GNDA.n1490 GNDA.n1460 585
R664 GNDA.n1490 GNDA.n48 585
R665 GNDA.n1493 GNDA.n1492 585
R666 GNDA.n1492 GNDA.n1491 585
R667 GNDA.n1494 GNDA.n1458 585
R668 GNDA.n1458 GNDA.n1457 585
R669 GNDA.n1496 GNDA.n1495 585
R670 GNDA.n1497 GNDA.n1496 585
R671 GNDA.n1459 GNDA.n1456 585
R672 GNDA.n1498 GNDA.n1456 585
R673 GNDA.n1500 GNDA.n1455 585
R674 GNDA.n1500 GNDA.n1499 585
R675 GNDA.n1503 GNDA.n1502 585
R676 GNDA.n1502 GNDA.n1501 585
R677 GNDA.n1504 GNDA.n1454 585
R678 GNDA.n1454 GNDA.n1453 585
R679 GNDA.n1506 GNDA.n1505 585
R680 GNDA.n1507 GNDA.n1506 585
R681 GNDA.n1451 GNDA.n1450 585
R682 GNDA.n1508 GNDA.n1451 585
R683 GNDA.n1510 GNDA.n1509 585
R684 GNDA.n1452 GNDA.n1449 585
R685 GNDA.n2419 GNDA.n61 585
R686 GNDA.n2419 GNDA.n43 585
R687 GNDA.n2422 GNDA.n2421 585
R688 GNDA.n2421 GNDA.n2420 585
R689 GNDA.n2423 GNDA.n60 585
R690 GNDA.n60 GNDA.n59 585
R691 GNDA.n2425 GNDA.n2424 585
R692 GNDA.n2426 GNDA.n2425 585
R693 GNDA.n58 GNDA.n57 585
R694 GNDA.n2427 GNDA.n58 585
R695 GNDA.n2430 GNDA.n2429 585
R696 GNDA.n2429 GNDA.n2428 585
R697 GNDA.n2431 GNDA.n56 585
R698 GNDA.n56 GNDA.n55 585
R699 GNDA.n2433 GNDA.n2432 585
R700 GNDA.n2434 GNDA.n2433 585
R701 GNDA.n54 GNDA.n53 585
R702 GNDA.n2435 GNDA.n54 585
R703 GNDA.n2438 GNDA.n2437 585
R704 GNDA.n2437 GNDA.n2436 585
R705 GNDA.n51 GNDA.n49 585
R706 GNDA.n2442 GNDA.n2441 585
R707 GNDA.n30 GNDA.n29 585
R708 GNDA.n2467 GNDA.n30 585
R709 GNDA.n2465 GNDA.n2464 585
R710 GNDA.n2466 GNDA.n2465 585
R711 GNDA.n2463 GNDA.n32 585
R712 GNDA.n32 GNDA.n31 585
R713 GNDA.n2462 GNDA.n2461 585
R714 GNDA.n2461 GNDA.n2460 585
R715 GNDA.n34 GNDA.n33 585
R716 GNDA.n2459 GNDA.n34 585
R717 GNDA.n2457 GNDA.n2456 585
R718 GNDA.n2458 GNDA.n2457 585
R719 GNDA.n2455 GNDA.n35 585
R720 GNDA.n2451 GNDA.n35 585
R721 GNDA.n2454 GNDA.n2453 585
R722 GNDA.n2453 GNDA.n2452 585
R723 GNDA.n37 GNDA.n36 585
R724 GNDA.n2450 GNDA.n37 585
R725 GNDA.n2448 GNDA.n2447 585
R726 GNDA.n2449 GNDA.n2448 585
R727 GNDA.n39 GNDA.n38 585
R728 GNDA.n2444 GNDA.n2443 585
R729 GNDA.n2494 GNDA.n2493 585
R730 GNDA.n2493 GNDA.n2492 585
R731 GNDA.n2470 GNDA.n2469 585
R732 GNDA.n2469 GNDA.n2468 585
R733 GNDA.n2471 GNDA.n28 585
R734 GNDA.n28 GNDA.n27 585
R735 GNDA.n2473 GNDA.n2472 585
R736 GNDA.n2474 GNDA.n2473 585
R737 GNDA.n25 GNDA.n24 585
R738 GNDA.n2475 GNDA.n25 585
R739 GNDA.n2478 GNDA.n2477 585
R740 GNDA.n2477 GNDA.n2476 585
R741 GNDA.n2479 GNDA.n23 585
R742 GNDA.n26 GNDA.n23 585
R743 GNDA.n2481 GNDA.n2480 585
R744 GNDA.n2482 GNDA.n2481 585
R745 GNDA.n22 GNDA.n21 585
R746 GNDA.n2483 GNDA.n22 585
R747 GNDA.n2486 GNDA.n2485 585
R748 GNDA.n2485 GNDA.n2484 585
R749 GNDA.n2487 GNDA.n19 585
R750 GNDA.n19 GNDA.n18 585
R751 GNDA.n2489 GNDA.n2488 585
R752 GNDA.n2490 GNDA.n2489 585
R753 GNDA.n20 GNDA.n17 585
R754 GNDA.n2491 GNDA.n17 585
R755 GNDA.n4 GNDA.n3 585
R756 GNDA.n2512 GNDA.n2511 585
R757 GNDA.n2513 GNDA.n2512 585
R758 GNDA.n1984 GNDA.n1983 585
R759 GNDA.n1983 GNDA.n1982 585
R760 GNDA.n2497 GNDA.n12 585
R761 GNDA.n2498 GNDA.n2497 585
R762 GNDA.n2501 GNDA.n2500 585
R763 GNDA.n2500 GNDA.n2499 585
R764 GNDA.n2502 GNDA.n11 585
R765 GNDA.n11 GNDA.n10 585
R766 GNDA.n2504 GNDA.n2503 585
R767 GNDA.n2505 GNDA.n2504 585
R768 GNDA.n9 GNDA.n7 585
R769 GNDA.n2506 GNDA.n9 585
R770 GNDA.n2509 GNDA.n2508 585
R771 GNDA.n2508 GNDA.n2507 585
R772 GNDA.n8 GNDA.n6 585
R773 GNDA.n8 GNDA.n5 585
R774 GNDA.n1972 GNDA.n1971 585
R775 GNDA.n1973 GNDA.n1972 585
R776 GNDA.n1976 GNDA.n1975 585
R777 GNDA.n1975 GNDA.n1974 585
R778 GNDA.n1977 GNDA.n1969 585
R779 GNDA.n1969 GNDA.n1968 585
R780 GNDA.n1979 GNDA.n1978 585
R781 GNDA.n1980 GNDA.n1979 585
R782 GNDA.n1970 GNDA.n453 585
R783 GNDA.n1981 GNDA.n453 585
R784 GNDA.n464 GNDA.n463 585
R785 GNDA.n1940 GNDA.n464 585
R786 GNDA.n1962 GNDA.n448 585
R787 GNDA.n1966 GNDA.n448 585
R788 GNDA.n1964 GNDA.n1963 585
R789 GNDA.n1965 GNDA.n1964 585
R790 GNDA.n1961 GNDA.n455 585
R791 GNDA.n455 GNDA.n454 585
R792 GNDA.n1960 GNDA.n1959 585
R793 GNDA.n1959 GNDA.n1958 585
R794 GNDA.n457 GNDA.n456 585
R795 GNDA.n1957 GNDA.n457 585
R796 GNDA.n1955 GNDA.n1954 585
R797 GNDA.n1956 GNDA.n1955 585
R798 GNDA.n1953 GNDA.n458 585
R799 GNDA.n1949 GNDA.n458 585
R800 GNDA.n1952 GNDA.n1951 585
R801 GNDA.n1951 GNDA.n1950 585
R802 GNDA.n460 GNDA.n459 585
R803 GNDA.n1948 GNDA.n460 585
R804 GNDA.n1946 GNDA.n1945 585
R805 GNDA.n1947 GNDA.n1946 585
R806 GNDA.n1944 GNDA.n462 585
R807 GNDA.n462 GNDA.n461 585
R808 GNDA.n1943 GNDA.n1942 585
R809 GNDA.n1942 GNDA.n1941 585
R810 GNDA.n871 GNDA.t234 535.191
R811 GNDA.n875 GNDA.t247 535.191
R812 GNDA.n968 GNDA.t299 535.191
R813 GNDA.n1051 GNDA.t284 535.191
R814 GNDA.n1855 GNDA.n1854 531.201
R815 GNDA.n1085 GNDA.n891 531.201
R816 GNDA.n1854 GNDA.n775 528
R817 GNDA.n647 GNDA.n495 512.884
R818 GNDA.n1840 GNDA.n815 512
R819 GNDA.n1840 GNDA.n1839 512
R820 GNDA.n1194 GNDA.n1189 512
R821 GNDA.n1194 GNDA.n1191 512
R822 GNDA.n817 GNDA.n815 508.8
R823 GNDA.n1839 GNDA.n817 508.8
R824 GNDA.n1190 GNDA.n1189 508.8
R825 GNDA.n1191 GNDA.n1190 508.8
R826 GNDA.n1941 GNDA.n1940 505.748
R827 GNDA.n1941 GNDA.n461 505.748
R828 GNDA.n1947 GNDA.n461 505.748
R829 GNDA.n1948 GNDA.n1947 505.748
R830 GNDA.n1950 GNDA.n1948 505.748
R831 GNDA.n1950 GNDA.n1949 505.748
R832 GNDA.n1957 GNDA.n1956 505.748
R833 GNDA.n1958 GNDA.n1957 505.748
R834 GNDA.n1958 GNDA.n454 505.748
R835 GNDA.n1965 GNDA.n454 505.748
R836 GNDA.n1966 GNDA.n1965 505.748
R837 GNDA.n1982 GNDA.n1981 505.748
R838 GNDA.n1981 GNDA.n1980 505.748
R839 GNDA.n1980 GNDA.n1968 505.748
R840 GNDA.n1974 GNDA.n1968 505.748
R841 GNDA.n1974 GNDA.n1973 505.748
R842 GNDA.n1973 GNDA.n5 505.748
R843 GNDA.n2507 GNDA.n2506 505.748
R844 GNDA.n2506 GNDA.n2505 505.748
R845 GNDA.n2505 GNDA.n10 505.748
R846 GNDA.n2499 GNDA.n10 505.748
R847 GNDA.n2499 GNDA.n2498 505.748
R848 GNDA.n2492 GNDA.n2491 505.748
R849 GNDA.n2491 GNDA.n2490 505.748
R850 GNDA.n2490 GNDA.n18 505.748
R851 GNDA.n2484 GNDA.n18 505.748
R852 GNDA.n2484 GNDA.n2483 505.748
R853 GNDA.n2483 GNDA.n2482 505.748
R854 GNDA.n2476 GNDA.n26 505.748
R855 GNDA.n2476 GNDA.n2475 505.748
R856 GNDA.n2475 GNDA.n2474 505.748
R857 GNDA.n2474 GNDA.n27 505.748
R858 GNDA.n2468 GNDA.n27 505.748
R859 GNDA.n1856 GNDA.n1855 499.2
R860 GNDA.n879 GNDA.n873 496
R861 GNDA.n1057 GNDA.n965 496
R862 GNDA.n936 GNDA.t311 493.418
R863 GNDA.n937 GNDA.t296 493.418
R864 GNDA.n938 GNDA.t319 493.418
R865 GNDA.n939 GNDA.t290 493.418
R866 GNDA.n884 GNDA.t308 493.418
R867 GNDA.n1104 GNDA.t302 493.418
R868 GNDA.n1103 GNDA.t277 493.418
R869 GNDA.n946 GNDA.t239 493.418
R870 GNDA.n947 GNDA.t221 493.418
R871 GNDA.n948 GNDA.t316 493.418
R872 GNDA.n1162 GNDA.n873 489.601
R873 GNDA.n1057 GNDA.n964 489.601
R874 GNDA.n775 GNDA.n471 486.401
R875 GNDA.n861 GNDA.n860 476.8
R876 GNDA.n1032 GNDA.n985 476.8
R877 GNDA.n1181 GNDA.n859 448
R878 GNDA.n1029 GNDA.n986 448
R879 GNDA.n1878 GNDA.n1874 444.8
R880 GNDA.n1878 GNDA.n1877 444.8
R881 GNDA.n1206 GNDA.n1205 444.695
R882 GNDA.n1875 GNDA.n1874 441.601
R883 GNDA.n1877 GNDA.n1876 438.401
R884 GNDA.n1937 GNDA.n468 435.2
R885 GNDA.n1139 GNDA.n890 428.8
R886 GNDA.n1937 GNDA.n1936 425.601
R887 GNDA.n941 GNDA.n940 422.401
R888 GNDA.n944 GNDA.n943 422.401
R889 GNDA.n1105 GNDA.n885 422.401
R890 GNDA.n1101 GNDA.n1100 422.401
R891 GNDA.n1935 GNDA.n470 422.401
R892 GNDA.n1936 GNDA.n1935 419.2
R893 GNDA.n841 GNDA.t293 413.084
R894 GNDA.n840 GNDA.t273 413.084
R895 GNDA.n828 GNDA.t228 413.084
R896 GNDA.n829 GNDA.t281 413.084
R897 GNDA.n1199 GNDA.t261 413.084
R898 GNDA.n844 GNDA.t287 413.084
R899 GNDA.n605 GNDA.t225 391.411
R900 GNDA.n1156 GNDA.n864 387.2
R901 GNDA.n1049 GNDA.n1048 387.2
R902 GNDA.n1178 GNDA.n864 380.8
R903 GNDA.n1049 GNDA.n970 380.8
R904 GNDA.n1206 GNDA.n848 377.149
R905 GNDA.n1086 GNDA.n890 355.2
R906 GNDA.n1693 GNDA.n1692 352.627
R907 GNDA.n1706 GNDA.n1682 352.627
R908 GNDA.n1707 GNDA.n1706 352.627
R909 GNDA.n1708 GNDA.n1707 352.627
R910 GNDA.n1708 GNDA.n1230 352.627
R911 GNDA.n1834 GNDA.n1230 352.627
R912 GNDA.n1956 GNDA.t225 342.784
R913 GNDA.n2507 GNDA.t227 342.784
R914 GNDA.n26 GNDA.t227 342.784
R915 GNDA.n1181 GNDA.n1180 342.401
R916 GNDA.n1030 GNDA.n1029 342.401
R917 GNDA.n1171 GNDA.n1164 332.8
R918 GNDA.n1037 GNDA.n981 332.8
R919 GNDA.n921 GNDA.t264 332.75
R920 GNDA.n923 GNDA.t250 332.75
R921 GNDA.t227 GNDA.n47 172.876
R922 GNDA.n44 GNDA.t227 172.876
R923 GNDA.n42 GNDA.t227 172.615
R924 GNDA.t227 GNDA.n45 172.615
R925 GNDA.n1225 GNDA.n822 323.2
R926 GNDA.n1173 GNDA.n1172 321.281
R927 GNDA.n1039 GNDA.n1038 321.281
R928 GNDA.n1172 GNDA.n1171 318.08
R929 GNDA.n1038 GNDA.n1037 318.08
R930 GNDA.n1223 GNDA.n822 316.8
R931 GNDA.n879 GNDA.n878 310.401
R932 GNDA.n1052 GNDA.n965 310.401
R933 GNDA.n1780 GNDA.n1617 304
R934 GNDA.n1162 GNDA.n872 304
R935 GNDA.n969 GNDA.n964 304
R936 GNDA.n1836 GNDA.n1229 303.363
R937 GNDA.n1782 GNDA.n1617 300.8
R938 GNDA.n1781 GNDA.n1780 300.8
R939 GNDA.n1114 GNDA.n1113 300.8
R940 GNDA.n1114 GNDA.n919 300.8
R941 GNDA.n1164 GNDA.n1163 300.8
R942 GNDA.n981 GNDA.n980 300.8
R943 GNDA.n1853 GNDA.n1852 300.257
R944 GNDA.n1782 GNDA.n1781 297.601
R945 GNDA.n1922 GNDA.n469 297.601
R946 GNDA.n1922 GNDA.n1921 297.601
R947 GNDA.n1920 GNDA.n484 297.601
R948 GNDA.n487 GNDA.n484 297.601
R949 GNDA.n1778 GNDA.n1777 296.411
R950 GNDA.n1003 GNDA.n1002 296
R951 GNDA.n1021 GNDA.n989 296
R952 GNDA.n1225 GNDA.n1224 294.401
R953 GNDA.n1214 GNDA.n825 294.401
R954 GNDA.n1218 GNDA.n825 294.401
R955 GNDA.n1040 GNDA.n1039 292.5
R956 GNDA.n1041 GNDA.n1040 292.5
R957 GNDA.n1038 GNDA.n979 292.5
R958 GNDA.n982 GNDA.n979 292.5
R959 GNDA.n1037 GNDA.n1036 292.5
R960 GNDA.n1036 GNDA.n1035 292.5
R961 GNDA.n981 GNDA.n978 292.5
R962 GNDA.n982 GNDA.n978 292.5
R963 GNDA.n967 GNDA.n965 292.5
R964 GNDA.n1045 GNDA.n967 292.5
R965 GNDA.n1057 GNDA.n1056 292.5
R966 GNDA.n1056 GNDA.n1055 292.5
R967 GNDA.n966 GNDA.n964 292.5
R968 GNDA.n1043 GNDA.n966 292.5
R969 GNDA.n1054 GNDA.n1053 292.5
R970 GNDA.n1055 GNDA.n1054 292.5
R971 GNDA.n1048 GNDA.n1047 292.5
R972 GNDA.n1047 GNDA.n1046 292.5
R973 GNDA.n1049 GNDA.n971 292.5
R974 GNDA.t341 GNDA.n971 292.5
R975 GNDA.n974 GNDA.n970 292.5
R976 GNDA.n1042 GNDA.n974 292.5
R977 GNDA.n1044 GNDA.n977 292.5
R978 GNDA.n1044 GNDA.t341 292.5
R979 GNDA.n1033 GNDA.n1032 292.5
R980 GNDA.n1034 GNDA.n1033 292.5
R981 GNDA.n1030 GNDA.n984 292.5
R982 GNDA.n1026 GNDA.n984 292.5
R983 GNDA.n1029 GNDA.n1028 292.5
R984 GNDA.n1028 GNDA.n1027 292.5
R985 GNDA.n985 GNDA.n983 292.5
R986 GNDA.n987 GNDA.n983 292.5
R987 GNDA.n1021 GNDA.n1020 292.5
R988 GNDA.n1020 GNDA.n1019 292.5
R989 GNDA.n1113 GNDA.n1112 292.5
R990 GNDA.n1112 GNDA.n1111 292.5
R991 GNDA.n1114 GNDA.n920 292.5
R992 GNDA.n958 GNDA.n920 292.5
R993 GNDA.n956 GNDA.n919 292.5
R994 GNDA.n957 GNDA.n956 292.5
R995 GNDA.n926 GNDA.n925 292.5
R996 GNDA.n958 GNDA.n926 292.5
R997 GNDA.n931 GNDA.n897 292.5
R998 GNDA.n932 GNDA.n931 292.5
R999 GNDA.n1131 GNDA.n895 292.5
R1000 GNDA.n930 GNDA.n895 292.5
R1001 GNDA.n1133 GNDA.n1132 292.5
R1002 GNDA.n1134 GNDA.n1133 292.5
R1003 GNDA.n896 GNDA.n894 292.5
R1004 GNDA.n930 GNDA.n894 292.5
R1005 GNDA.n962 GNDA.n961 292.5
R1006 GNDA.n961 GNDA.n960 292.5
R1007 GNDA.n1092 GNDA.n951 292.5
R1008 GNDA.n955 GNDA.n951 292.5
R1009 GNDA.n1095 GNDA.n1094 292.5
R1010 GNDA.n1096 GNDA.n1095 292.5
R1011 GNDA.n952 GNDA.n950 292.5
R1012 GNDA.n955 GNDA.n950 292.5
R1013 GNDA.n1138 GNDA.n1137 292.5
R1014 GNDA.n1137 GNDA.n881 292.5
R1015 GNDA.n1136 GNDA.n890 292.5
R1016 GNDA.n1136 GNDA.n1135 292.5
R1017 GNDA.n1085 GNDA.n893 292.5
R1018 GNDA.n959 GNDA.n893 292.5
R1019 GNDA.n892 GNDA.n891 292.5
R1020 GNDA.n1135 GNDA.n892 292.5
R1021 GNDA.n1149 GNDA.n1148 292.5
R1022 GNDA.n1150 GNDA.n1149 292.5
R1023 GNDA.n886 GNDA.n883 292.5
R1024 GNDA.n1110 GNDA.n883 292.5
R1025 GNDA.n1099 GNDA.n1098 292.5
R1026 GNDA.n1098 GNDA.n1097 292.5
R1027 GNDA.n1107 GNDA.n882 292.5
R1028 GNDA.n1110 GNDA.n882 292.5
R1029 GNDA.n945 GNDA.n934 292.5
R1030 GNDA.n934 GNDA.n933 292.5
R1031 GNDA.n1109 GNDA.n1108 292.5
R1032 GNDA.n1110 GNDA.n1109 292.5
R1033 GNDA.n935 GNDA.n929 292.5
R1034 GNDA.n954 GNDA.n929 292.5
R1035 GNDA.n942 GNDA.n928 292.5
R1036 GNDA.n1110 GNDA.n928 292.5
R1037 GNDA.n1174 GNDA.n1173 292.5
R1038 GNDA.n1175 GNDA.n1174 292.5
R1039 GNDA.n1162 GNDA.n1161 292.5
R1040 GNDA.n1161 GNDA.n867 292.5
R1041 GNDA.n1160 GNDA.n873 292.5
R1042 GNDA.n1160 GNDA.n1159 292.5
R1043 GNDA.n880 GNDA.n879 292.5
R1044 GNDA.n1152 GNDA.n880 292.5
R1045 GNDA.n877 GNDA.n874 292.5
R1046 GNDA.n1159 GNDA.n874 292.5
R1047 GNDA.n1178 GNDA.n1177 292.5
R1048 GNDA.n1177 GNDA.n1176 292.5
R1049 GNDA.n866 GNDA.n864 292.5
R1050 GNDA.t178 GNDA.n866 292.5
R1051 GNDA.n1157 GNDA.n1156 292.5
R1052 GNDA.n1158 GNDA.n1157 292.5
R1053 GNDA.n1154 GNDA.n865 292.5
R1054 GNDA.t178 GNDA.n865 292.5
R1055 GNDA.n1002 GNDA.n1001 292.5
R1056 GNDA.n1001 GNDA.n996 292.5
R1057 GNDA.n1171 GNDA.n1170 292.5
R1058 GNDA.n1170 GNDA.n1169 292.5
R1059 GNDA.n1172 GNDA.n870 292.5
R1060 GNDA.n1165 GNDA.n870 292.5
R1061 GNDA.n1164 GNDA.n869 292.5
R1062 GNDA.n1165 GNDA.n869 292.5
R1063 GNDA.n1213 GNDA.n1212 292.5
R1064 GNDA.n1212 GNDA.n1211 292.5
R1065 GNDA.n1202 GNDA.n1201 292.5
R1066 GNDA.n1203 GNDA.n1202 292.5
R1067 GNDA.n1197 GNDA.n843 292.5
R1068 GNDA.n1198 GNDA.n1197 292.5
R1069 GNDA.n1219 GNDA.n1218 292.5
R1070 GNDA.n1220 GNDA.n1219 292.5
R1071 GNDA.n1216 GNDA.n782 292.5
R1072 GNDA.n1848 GNDA.n782 292.5
R1073 GNDA.n1214 GNDA.n842 292.5
R1074 GNDA.n1210 GNDA.n842 292.5
R1075 GNDA.n825 GNDA.n781 292.5
R1076 GNDA.n1848 GNDA.n781 292.5
R1077 GNDA.n836 GNDA.n835 292.5
R1078 GNDA.n835 GNDA.n819 292.5
R1079 GNDA.n839 GNDA.n827 292.5
R1080 GNDA.n830 GNDA.n827 292.5
R1081 GNDA.n833 GNDA.n826 292.5
R1082 GNDA.n833 GNDA.n832 292.5
R1083 GNDA.n1845 GNDA.n784 292.5
R1084 GNDA.n1228 GNDA.n784 292.5
R1085 GNDA.n1847 GNDA.n1846 292.5
R1086 GNDA.n1848 GNDA.n1847 292.5
R1087 GNDA.n785 GNDA.n783 292.5
R1088 GNDA.n849 GNDA.n783 292.5
R1089 GNDA.n1844 GNDA.n780 292.5
R1090 GNDA.n1848 GNDA.n780 292.5
R1091 GNDA.n1191 GNDA.n1188 292.5
R1092 GNDA.n1188 GNDA.n1187 292.5
R1093 GNDA.n1195 GNDA.n1194 292.5
R1094 GNDA.n1196 GNDA.n1195 292.5
R1095 GNDA.n1189 GNDA.n1186 292.5
R1096 GNDA.n1186 GNDA.n1185 292.5
R1097 GNDA.n1190 GNDA.n850 292.5
R1098 GNDA.n1196 GNDA.n850 292.5
R1099 GNDA.n1839 GNDA.n1838 292.5
R1100 GNDA.n1838 GNDA.n1837 292.5
R1101 GNDA.n1840 GNDA.n816 292.5
R1102 GNDA.n831 GNDA.n816 292.5
R1103 GNDA.n823 GNDA.n815 292.5
R1104 GNDA.n824 GNDA.n823 292.5
R1105 GNDA.n818 GNDA.n817 292.5
R1106 GNDA.n831 GNDA.n818 292.5
R1107 GNDA.n1182 GNDA.n1181 292.5
R1108 GNDA.n1183 GNDA.n1182 292.5
R1109 GNDA.n1180 GNDA.n858 292.5
R1110 GNDA.n1168 GNDA.n858 292.5
R1111 GNDA.n1166 GNDA.n861 292.5
R1112 GNDA.n1167 GNDA.n1166 292.5
R1113 GNDA.n860 GNDA.n857 292.5
R1114 GNDA.n1168 GNDA.n857 292.5
R1115 GNDA.n1208 GNDA.n1207 292.5
R1116 GNDA.n1209 GNDA.n1208 292.5
R1117 GNDA.n1205 GNDA.n1204 292.5
R1118 GNDA.n1196 GNDA.n848 292.5
R1119 GNDA.n1226 GNDA.n1225 292.5
R1120 GNDA.n1227 GNDA.n1226 292.5
R1121 GNDA.n1224 GNDA.n821 292.5
R1122 GNDA.n831 GNDA.n821 292.5
R1123 GNDA.n1223 GNDA.n1222 292.5
R1124 GNDA.n1222 GNDA.n1221 292.5
R1125 GNDA.n822 GNDA.n820 292.5
R1126 GNDA.n831 GNDA.n820 292.5
R1127 GNDA.n486 GNDA.n485 292.5
R1128 GNDA.n1895 GNDA.n486 292.5
R1129 GNDA.n488 GNDA.n487 292.5
R1130 GNDA.n1918 GNDA.n488 292.5
R1131 GNDA.n484 GNDA.n479 292.5
R1132 GNDA.n1924 GNDA.n479 292.5
R1133 GNDA.n1920 GNDA.n1919 292.5
R1134 GNDA.n1919 GNDA.n1918 292.5
R1135 GNDA.n1783 GNDA.n1782 292.5
R1136 GNDA.n1784 GNDA.n1783 292.5
R1137 GNDA.n1781 GNDA.n1616 292.5
R1138 GNDA.n1626 GNDA.n1616 292.5
R1139 GNDA.n1780 GNDA.n1779 292.5
R1140 GNDA.n1779 GNDA.n1778 292.5
R1141 GNDA.n1617 GNDA.n1615 292.5
R1142 GNDA.n1626 GNDA.n1615 292.5
R1143 GNDA.n1894 GNDA.n483 292.5
R1144 GNDA.n1895 GNDA.n1894 292.5
R1145 GNDA.n1921 GNDA.n482 292.5
R1146 GNDA.n1918 GNDA.n482 292.5
R1147 GNDA.n1923 GNDA.n1922 292.5
R1148 GNDA.n1924 GNDA.n1923 292.5
R1149 GNDA.n481 GNDA.n469 292.5
R1150 GNDA.n1918 GNDA.n481 292.5
R1151 GNDA.n1857 GNDA.n1856 292.5
R1152 GNDA.n1858 GNDA.n1857 292.5
R1153 GNDA.n775 GNDA.n774 292.5
R1154 GNDA.n1626 GNDA.n774 292.5
R1155 GNDA.n1854 GNDA.n1853 292.5
R1156 GNDA.n1855 GNDA.n773 292.5
R1157 GNDA.n1626 GNDA.n773 292.5
R1158 GNDA.n1875 GNDA.n648 292.5
R1159 GNDA.n1880 GNDA.n648 292.5
R1160 GNDA.n1874 GNDA.n1872 292.5
R1161 GNDA.n1872 GNDA.n1871 292.5
R1162 GNDA.n1879 GNDA.n1878 292.5
R1163 GNDA.n1880 GNDA.n1879 292.5
R1164 GNDA.n1877 GNDA.n1873 292.5
R1165 GNDA.n1873 GNDA.n465 292.5
R1166 GNDA.n1938 GNDA.n1937 292.5
R1167 GNDA.n1939 GNDA.n1938 292.5
R1168 GNDA.n468 GNDA.n466 292.5
R1169 GNDA.n1918 GNDA.n466 292.5
R1170 GNDA.n1935 GNDA.n1934 292.5
R1171 GNDA.n1934 GNDA.n1933 292.5
R1172 GNDA.n1936 GNDA.n467 292.5
R1173 GNDA.n1918 GNDA.n467 292.5
R1174 GNDA.n483 GNDA.n469 291.2
R1175 GNDA.n1921 GNDA.n483 291.2
R1176 GNDA.n1920 GNDA.n485 291.2
R1177 GNDA.n487 GNDA.n485 291.2
R1178 GNDA.n1224 GNDA.n1223 288
R1179 GNDA.n838 GNDA.n837 281.601
R1180 GNDA.n1200 GNDA.n845 281.601
R1181 GNDA.n836 GNDA.n826 278.401
R1182 GNDA.n1201 GNDA.n843 278.401
R1183 GNDA.n921 GNDA.t265 258.601
R1184 GNDA.n923 GNDA.t252 258.601
R1185 GNDA.n301 GNDA.n242 258.334
R1186 GNDA.n1294 GNDA.n1249 258.334
R1187 GNDA.n1731 GNDA.n1673 258.334
R1188 GNDA.n2085 GNDA.n2030 258.334
R1189 GNDA.n147 GNDA.n88 258.334
R1190 GNDA.n564 GNDA.n522 258.334
R1191 GNDA.n2238 GNDA.n2170 258.334
R1192 GNDA.n729 GNDA.n675 258.334
R1193 GNDA.n1402 GNDA.n1357 258.334
R1194 GNDA.n2441 GNDA.n50 257.466
R1195 GNDA.n1566 GNDA.n1341 257.466
R1196 GNDA.n2131 GNDA.n412 257.466
R1197 GNDA.n2154 GNDA.n393 257.466
R1198 GNDA.n2388 GNDA.n193 257.466
R1199 GNDA.n2444 GNDA.n41 257.466
R1200 GNDA.n2347 GNDA.n346 257.466
R1201 GNDA.n1514 GNDA.n1449 257.466
R1202 GNDA.n1833 GNDA.n1232 257.466
R1203 GNDA.n1512 GNDA.n1511 254.442
R1204 GNDA.n2367 GNDA.n2366 254.34
R1205 GNDA.n2368 GNDA.n2367 254.34
R1206 GNDA.n2367 GNDA.n2365 254.34
R1207 GNDA.n2367 GNDA.n2363 254.34
R1208 GNDA.n2367 GNDA.n2362 254.34
R1209 GNDA.n2367 GNDA.n191 254.34
R1210 GNDA.n194 GNDA.n13 254.34
R1211 GNDA.n2370 GNDA.n194 254.34
R1212 GNDA.n2377 GNDA.n194 254.34
R1213 GNDA.n201 GNDA.n194 254.34
R1214 GNDA.n2384 GNDA.n194 254.34
R1215 GNDA.n2387 GNDA.n194 254.34
R1216 GNDA.n2126 GNDA.n2125 254.34
R1217 GNDA.n2125 GNDA.n2124 254.34
R1218 GNDA.n2125 GNDA.n2013 254.34
R1219 GNDA.n2125 GNDA.n2012 254.34
R1220 GNDA.n2125 GNDA.n2011 254.34
R1221 GNDA.n2125 GNDA.n2010 254.34
R1222 GNDA.n2324 GNDA.n2323 254.34
R1223 GNDA.n2323 GNDA.n2322 254.34
R1224 GNDA.n2323 GNDA.n368 254.34
R1225 GNDA.n2323 GNDA.n367 254.34
R1226 GNDA.n2323 GNDA.n366 254.34
R1227 GNDA.n2323 GNDA.n365 254.34
R1228 GNDA.n2271 GNDA.n2270 254.34
R1229 GNDA.n2271 GNDA.n387 254.34
R1230 GNDA.n2271 GNDA.n386 254.34
R1231 GNDA.n2271 GNDA.n385 254.34
R1232 GNDA.n2271 GNDA.n384 254.34
R1233 GNDA.n2271 GNDA.n383 254.34
R1234 GNDA.n1526 GNDA.n1229 254.34
R1235 GNDA.n1424 GNDA.n1229 254.34
R1236 GNDA.n1435 GNDA.n1229 254.34
R1237 GNDA.n1437 GNDA.n1229 254.34
R1238 GNDA.n1447 GNDA.n1229 254.34
R1239 GNDA.n1515 GNDA.n1229 254.34
R1240 GNDA.n1866 GNDA.n651 254.34
R1241 GNDA.n1887 GNDA.n492 254.34
R1242 GNDA.n427 GNDA.n426 254.34
R1243 GNDA.n427 GNDA.n424 254.34
R1244 GNDA.n427 GNDA.n423 254.34
R1245 GNDA.n427 GNDA.n421 254.34
R1246 GNDA.n427 GNDA.n420 254.34
R1247 GNDA.n427 GNDA.n417 254.34
R1248 GNDA.n450 GNDA.n427 254.34
R1249 GNDA.n444 GNDA.n427 254.34
R1250 GNDA.n441 GNDA.n427 254.34
R1251 GNDA.n435 GNDA.n427 254.34
R1252 GNDA.n432 GNDA.n427 254.34
R1253 GNDA.n2006 GNDA.n427 254.34
R1254 GNDA.n2136 GNDA.n394 254.34
R1255 GNDA.n407 GNDA.n394 254.34
R1256 GNDA.n2143 GNDA.n394 254.34
R1257 GNDA.n401 GNDA.n394 254.34
R1258 GNDA.n2150 GNDA.n394 254.34
R1259 GNDA.n2153 GNDA.n394 254.34
R1260 GNDA.n1987 GNDA.n394 254.34
R1261 GNDA.n447 GNDA.n394 254.34
R1262 GNDA.n1994 GNDA.n394 254.34
R1263 GNDA.n438 GNDA.n394 254.34
R1264 GNDA.n2001 GNDA.n394 254.34
R1265 GNDA.n430 GNDA.n394 254.34
R1266 GNDA.n770 GNDA.n769 254.34
R1267 GNDA.n769 GNDA.n768 254.34
R1268 GNDA.n769 GNDA.n657 254.34
R1269 GNDA.n769 GNDA.n656 254.34
R1270 GNDA.n769 GNDA.n655 254.34
R1271 GNDA.n769 GNDA.n654 254.34
R1272 GNDA.n1809 GNDA.n1808 254.34
R1273 GNDA.n1808 GNDA.n1807 254.34
R1274 GNDA.n1808 GNDA.n1610 254.34
R1275 GNDA.n1808 GNDA.n1609 254.34
R1276 GNDA.n1808 GNDA.n1608 254.34
R1277 GNDA.n1808 GNDA.n1607 254.34
R1278 GNDA.n1653 GNDA.n1652 254.34
R1279 GNDA.n1772 GNDA.n1771 254.34
R1280 GNDA.n1771 GNDA.n1770 254.34
R1281 GNDA.n1578 GNDA.n1229 254.34
R1282 GNDA.n1316 GNDA.n1229 254.34
R1283 GNDA.n1327 GNDA.n1229 254.34
R1284 GNDA.n1329 GNDA.n1229 254.34
R1285 GNDA.n1339 GNDA.n1229 254.34
R1286 GNDA.n1567 GNDA.n1229 254.34
R1287 GNDA.n1602 GNDA.n427 254.34
R1288 GNDA.n1600 GNDA.n427 254.34
R1289 GNDA.n1597 GNDA.n427 254.34
R1290 GNDA.n1591 GNDA.n427 254.34
R1291 GNDA.n1588 GNDA.n427 254.34
R1292 GNDA.n1582 GNDA.n427 254.34
R1293 GNDA.n1812 GNDA.n394 254.34
R1294 GNDA.n1605 GNDA.n394 254.34
R1295 GNDA.n1819 GNDA.n394 254.34
R1296 GNDA.n1594 GNDA.n394 254.34
R1297 GNDA.n1826 GNDA.n394 254.34
R1298 GNDA.n1585 GNDA.n394 254.34
R1299 GNDA.n2273 GNDA.n222 254.34
R1300 GNDA.n2278 GNDA.n2273 254.34
R1301 GNDA.n2285 GNDA.n2273 254.34
R1302 GNDA.n2276 GNDA.n2273 254.34
R1303 GNDA.n2292 GNDA.n2273 254.34
R1304 GNDA.n2273 GNDA.n382 254.34
R1305 GNDA.n1488 GNDA.n42 254.34
R1306 GNDA.n1482 GNDA.n42 254.34
R1307 GNDA.n1480 GNDA.n42 254.34
R1308 GNDA.n1474 GNDA.n42 254.34
R1309 GNDA.n1472 GNDA.n42 254.34
R1310 GNDA.n1467 GNDA.n42 254.34
R1311 GNDA.n2367 GNDA.n2359 254.34
R1312 GNDA.n2367 GNDA.n216 254.34
R1313 GNDA.n2367 GNDA.n215 254.34
R1314 GNDA.n2367 GNDA.n214 254.34
R1315 GNDA.n2367 GNDA.n213 254.34
R1316 GNDA.n2367 GNDA.n212 254.34
R1317 GNDA.n221 GNDA.n194 254.34
R1318 GNDA.n1545 GNDA.n194 254.34
R1319 GNDA.n1552 GNDA.n194 254.34
R1320 GNDA.n1540 GNDA.n194 254.34
R1321 GNDA.n1559 GNDA.n194 254.34
R1322 GNDA.n1533 GNDA.n194 254.34
R1323 GNDA.n2367 GNDA.n211 254.34
R1324 GNDA.n2367 GNDA.n210 254.34
R1325 GNDA.n2367 GNDA.n209 254.34
R1326 GNDA.n2367 GNDA.n208 254.34
R1327 GNDA.n2367 GNDA.n207 254.34
R1328 GNDA.n2367 GNDA.n206 254.34
R1329 GNDA.n2329 GNDA.n194 254.34
R1330 GNDA.n363 GNDA.n194 254.34
R1331 GNDA.n2336 GNDA.n194 254.34
R1332 GNDA.n356 GNDA.n194 254.34
R1333 GNDA.n2343 GNDA.n194 254.34
R1334 GNDA.n2346 GNDA.n194 254.34
R1335 GNDA.n226 GNDA.n47 254.34
R1336 GNDA.n229 GNDA.n47 254.34
R1337 GNDA.n262 GNDA.n47 254.34
R1338 GNDA.n264 GNDA.n47 254.34
R1339 GNDA.n277 GNDA.n47 254.34
R1340 GNDA.n279 GNDA.n47 254.34
R1341 GNDA.n62 GNDA.n45 254.34
R1342 GNDA.n2413 GNDA.n45 254.34
R1343 GNDA.n2407 GNDA.n45 254.34
R1344 GNDA.n2405 GNDA.n45 254.34
R1345 GNDA.n2399 GNDA.n45 254.34
R1346 GNDA.n2397 GNDA.n45 254.34
R1347 GNDA.n72 GNDA.n44 254.34
R1348 GNDA.n75 GNDA.n44 254.34
R1349 GNDA.n108 GNDA.n44 254.34
R1350 GNDA.n110 GNDA.n44 254.34
R1351 GNDA.n123 GNDA.n44 254.34
R1352 GNDA.n125 GNDA.n44 254.34
R1353 GNDA.n2440 GNDA.n2439 254.34
R1354 GNDA.n2446 GNDA.n2445 254.34
R1355 GNDA.n2419 GNDA.n2418 251.614
R1356 GNDA.n2356 GNDA.n2355 251.614
R1357 GNDA.n1986 GNDA.n448 251.614
R1358 GNDA.n2135 GNDA.n2133 251.614
R1359 GNDA.n2497 GNDA.n2496 251.614
R1360 GNDA.n2469 GNDA.n30 251.614
R1361 GNDA.n2328 GNDA.n2325 251.614
R1362 GNDA.n1490 GNDA.n1489 251.614
R1363 GNDA.n1811 GNDA.n1810 251.614
R1364 GNDA.n2514 GNDA.n2513 250.349
R1365 GNDA.n1180 GNDA.n1179 246.4
R1366 GNDA.n1031 GNDA.n1030 246.4
R1367 GNDA.n839 GNDA.n826 240
R1368 GNDA.n1213 GNDA.n843 240
R1369 GNDA.n1682 GNDA.t225 239.004
R1370 GNDA.n1000 GNDA.n999 238.4
R1371 GNDA.n1023 GNDA.n1022 238.4
R1372 GNDA.n1094 GNDA.n952 233.601
R1373 GNDA.n962 GNDA.n952 233.601
R1374 GNDA.n915 GNDA.n913 227.096
R1375 GNDA.n912 GNDA.n910 227.096
R1376 GNDA.n1852 GNDA.n1851 226.805
R1377 GNDA.n915 GNDA.n914 226.534
R1378 GNDA.n912 GNDA.n911 226.534
R1379 GNDA.n871 GNDA.t236 224.525
R1380 GNDA.n875 GNDA.t249 224.525
R1381 GNDA.n968 GNDA.t301 224.525
R1382 GNDA.n1051 GNDA.t286 224.525
R1383 GNDA.n918 GNDA.n917 222.034
R1384 GNDA.n897 GNDA.n896 217.601
R1385 GNDA.n1132 GNDA.n896 214.4
R1386 GNDA.n925 GNDA.n924 211.201
R1387 GNDA.n925 GNDA.n922 211.201
R1388 GNDA.n1155 GNDA.n1154 211.201
R1389 GNDA.n1154 GNDA.n863 211.201
R1390 GNDA.n977 GNDA.n976 211.201
R1391 GNDA.n977 GNDA.n973 211.201
R1392 GNDA.n1852 GNDA.n776 209.417
R1393 GNDA.n1119 GNDA.n1117 206.052
R1394 GNDA.n900 GNDA.n898 206.052
R1395 GNDA.n1127 GNDA.n1126 205.488
R1396 GNDA.n1125 GNDA.n1124 205.488
R1397 GNDA.n1123 GNDA.n1122 205.488
R1398 GNDA.n1121 GNDA.n1120 205.488
R1399 GNDA.n1119 GNDA.n1118 205.488
R1400 GNDA.n908 GNDA.n907 205.488
R1401 GNDA.n906 GNDA.n905 205.488
R1402 GNDA.n904 GNDA.n903 205.488
R1403 GNDA.n902 GNDA.n901 205.488
R1404 GNDA.n900 GNDA.n899 205.488
R1405 GNDA.n1132 GNDA.n1131 203.201
R1406 GNDA.n1130 GNDA.n897 201.601
R1407 GNDA.n2512 GNDA.n4 197
R1408 GNDA.n2350 GNDA.n2349 195.049
R1409 GNDA.n1581 GNDA.n1580 195.049
R1410 GNDA.n1882 GNDA.n494 195.049
R1411 GNDA.n1861 GNDA.n772 195.049
R1412 GNDA.n2008 GNDA.n2007 195.049
R1413 GNDA.n2391 GNDA.n2390 195.049
R1414 GNDA.n391 GNDA.n389 195.049
R1415 GNDA.n1529 GNDA.n1528 195.049
R1416 GNDA.n1621 GNDA.n1619 195.049
R1417 GNDA.n1017 GNDA.n989 195
R1418 GNDA.n1018 GNDA.n1017 195
R1419 GNDA.n1024 GNDA.n1023 195
R1420 GNDA.n1025 GNDA.n1024 195
R1421 GNDA.n999 GNDA.n998 195
R1422 GNDA.n998 GNDA.n851 195
R1423 GNDA.n1004 GNDA.n1003 195
R1424 GNDA.n1005 GNDA.n1004 195
R1425 GNDA.n878 GNDA.n877 192
R1426 GNDA.n1053 GNDA.n1052 192
R1427 GNDA.t227 GNDA.n2442 190.773
R1428 GNDA.n2443 GNDA.t227 190.773
R1429 GNDA.n2326 GNDA.n68 187.249
R1430 GNDA.n2299 GNDA.n376 187.249
R1431 GNDA.n1897 GNDA.n464 187.249
R1432 GNDA.n645 GNDA.n497 187.249
R1433 GNDA.n1983 GNDA.n451 187.249
R1434 GNDA.n2493 GNDA.n15 187.249
R1435 GNDA.n2301 GNDA.n371 187.249
R1436 GNDA.n2358 GNDA.n218 187.249
R1437 GNDA.n1786 GNDA.n1613 187.249
R1438 GNDA.t227 GNDA.n48 186.691
R1439 GNDA.t227 GNDA.n43 186.691
R1440 GNDA.n299 GNDA.n242 185
R1441 GNDA.n242 GNDA.t276 185
R1442 GNDA.n298 GNDA.n297 185
R1443 GNDA.n295 GNDA.n243 185
R1444 GNDA.n294 GNDA.n244 185
R1445 GNDA.n292 GNDA.n291 185
R1446 GNDA.n290 GNDA.n245 185
R1447 GNDA.n289 GNDA.n288 185
R1448 GNDA.n286 GNDA.n246 185
R1449 GNDA.n286 GNDA.t276 185
R1450 GNDA.n285 GNDA.n247 185
R1451 GNDA.n301 GNDA.n300 185
R1452 GNDA.n303 GNDA.n240 185
R1453 GNDA.n305 GNDA.n304 185
R1454 GNDA.n306 GNDA.n239 185
R1455 GNDA.n308 GNDA.n307 185
R1456 GNDA.n310 GNDA.n237 185
R1457 GNDA.n312 GNDA.n311 185
R1458 GNDA.n313 GNDA.n236 185
R1459 GNDA.n315 GNDA.n314 185
R1460 GNDA.n317 GNDA.n235 185
R1461 GNDA.n320 GNDA.n319 185
R1462 GNDA.n321 GNDA.n234 185
R1463 GNDA.n323 GNDA.n322 185
R1464 GNDA.n325 GNDA.n233 185
R1465 GNDA.n328 GNDA.n327 185
R1466 GNDA.n329 GNDA.n232 185
R1467 GNDA.n331 GNDA.n330 185
R1468 GNDA.n333 GNDA.n227 185
R1469 GNDA.n1296 GNDA.n1249 185
R1470 GNDA.t226 GNDA.n1249 185
R1471 GNDA.n1298 GNDA.n1297 185
R1472 GNDA.n1300 GNDA.n1299 185
R1473 GNDA.n1302 GNDA.n1301 185
R1474 GNDA.n1304 GNDA.n1303 185
R1475 GNDA.n1306 GNDA.n1305 185
R1476 GNDA.n1308 GNDA.n1307 185
R1477 GNDA.n1309 GNDA.n1254 185
R1478 GNDA.t226 GNDA.n1254 185
R1479 GNDA.n1310 GNDA.n1258 185
R1480 GNDA.n1295 GNDA.n1294 185
R1481 GNDA.n1293 GNDA.n1292 185
R1482 GNDA.n1291 GNDA.n1290 185
R1483 GNDA.n1289 GNDA.n1288 185
R1484 GNDA.n1287 GNDA.n1286 185
R1485 GNDA.n1285 GNDA.n1284 185
R1486 GNDA.n1283 GNDA.n1282 185
R1487 GNDA.n1281 GNDA.n1280 185
R1488 GNDA.n1279 GNDA.n1278 185
R1489 GNDA.n1277 GNDA.n1276 185
R1490 GNDA.n1275 GNDA.n1274 185
R1491 GNDA.n1273 GNDA.n1272 185
R1492 GNDA.n1271 GNDA.n1270 185
R1493 GNDA.n1269 GNDA.n1268 185
R1494 GNDA.n1267 GNDA.n1266 185
R1495 GNDA.n1265 GNDA.n1264 185
R1496 GNDA.n1263 GNDA.n1262 185
R1497 GNDA.n1261 GNDA.n1239 185
R1498 GNDA.n1729 GNDA.n1673 185
R1499 GNDA.n1673 GNDA.t224 185
R1500 GNDA.n1728 GNDA.n1727 185
R1501 GNDA.n1725 GNDA.n1674 185
R1502 GNDA.n1724 GNDA.n1675 185
R1503 GNDA.n1722 GNDA.n1721 185
R1504 GNDA.n1720 GNDA.n1676 185
R1505 GNDA.n1719 GNDA.n1718 185
R1506 GNDA.n1716 GNDA.n1677 185
R1507 GNDA.n1716 GNDA.t224 185
R1508 GNDA.n1715 GNDA.n1678 185
R1509 GNDA.n1731 GNDA.n1730 185
R1510 GNDA.n1733 GNDA.n1671 185
R1511 GNDA.n1735 GNDA.n1734 185
R1512 GNDA.n1736 GNDA.n1670 185
R1513 GNDA.n1738 GNDA.n1737 185
R1514 GNDA.n1740 GNDA.n1668 185
R1515 GNDA.n1742 GNDA.n1741 185
R1516 GNDA.n1743 GNDA.n1667 185
R1517 GNDA.n1745 GNDA.n1744 185
R1518 GNDA.n1747 GNDA.n1666 185
R1519 GNDA.n1749 GNDA.n1748 185
R1520 GNDA.n1751 GNDA.n1750 185
R1521 GNDA.n1754 GNDA.n1753 185
R1522 GNDA.n1755 GNDA.n1664 185
R1523 GNDA.n1757 GNDA.n1756 185
R1524 GNDA.n1759 GNDA.n1663 185
R1525 GNDA.n1761 GNDA.n1760 185
R1526 GNDA.n1763 GNDA.n1762 185
R1527 GNDA.n2083 GNDA.n2030 185
R1528 GNDA.n2030 GNDA.t315 185
R1529 GNDA.n2082 GNDA.n2081 185
R1530 GNDA.n2079 GNDA.n2031 185
R1531 GNDA.n2078 GNDA.n2032 185
R1532 GNDA.n2076 GNDA.n2075 185
R1533 GNDA.n2074 GNDA.n2033 185
R1534 GNDA.n2073 GNDA.n2072 185
R1535 GNDA.n2070 GNDA.n2034 185
R1536 GNDA.n2070 GNDA.t315 185
R1537 GNDA.n2069 GNDA.n2035 185
R1538 GNDA.n2085 GNDA.n2084 185
R1539 GNDA.n2087 GNDA.n2028 185
R1540 GNDA.n2089 GNDA.n2088 185
R1541 GNDA.n2090 GNDA.n2027 185
R1542 GNDA.n2092 GNDA.n2091 185
R1543 GNDA.n2094 GNDA.n2025 185
R1544 GNDA.n2096 GNDA.n2095 185
R1545 GNDA.n2097 GNDA.n2024 185
R1546 GNDA.n2099 GNDA.n2098 185
R1547 GNDA.n2101 GNDA.n2023 185
R1548 GNDA.n2103 GNDA.n2102 185
R1549 GNDA.n2105 GNDA.n2104 185
R1550 GNDA.n2108 GNDA.n2107 185
R1551 GNDA.n2109 GNDA.n2021 185
R1552 GNDA.n2111 GNDA.n2110 185
R1553 GNDA.n2113 GNDA.n2020 185
R1554 GNDA.n2115 GNDA.n2114 185
R1555 GNDA.n2117 GNDA.n2116 185
R1556 GNDA.n145 GNDA.n88 185
R1557 GNDA.n88 GNDA.t237 185
R1558 GNDA.n144 GNDA.n143 185
R1559 GNDA.n141 GNDA.n89 185
R1560 GNDA.n140 GNDA.n90 185
R1561 GNDA.n138 GNDA.n137 185
R1562 GNDA.n136 GNDA.n91 185
R1563 GNDA.n135 GNDA.n134 185
R1564 GNDA.n132 GNDA.n92 185
R1565 GNDA.n132 GNDA.t237 185
R1566 GNDA.n131 GNDA.n93 185
R1567 GNDA.n147 GNDA.n146 185
R1568 GNDA.n149 GNDA.n86 185
R1569 GNDA.n151 GNDA.n150 185
R1570 GNDA.n152 GNDA.n85 185
R1571 GNDA.n154 GNDA.n153 185
R1572 GNDA.n156 GNDA.n83 185
R1573 GNDA.n158 GNDA.n157 185
R1574 GNDA.n159 GNDA.n82 185
R1575 GNDA.n161 GNDA.n160 185
R1576 GNDA.n163 GNDA.n81 185
R1577 GNDA.n166 GNDA.n165 185
R1578 GNDA.n167 GNDA.n80 185
R1579 GNDA.n169 GNDA.n168 185
R1580 GNDA.n171 GNDA.n79 185
R1581 GNDA.n174 GNDA.n173 185
R1582 GNDA.n175 GNDA.n78 185
R1583 GNDA.n177 GNDA.n176 185
R1584 GNDA.n179 GNDA.n73 185
R1585 GNDA.n180 GNDA.n74 185
R1586 GNDA.n183 GNDA.n182 185
R1587 GNDA.n104 GNDA.n77 185
R1588 GNDA.n105 GNDA.n101 185
R1589 GNDA.n114 GNDA.n113 185
R1590 GNDA.n116 GNDA.n99 185
R1591 GNDA.n119 GNDA.n118 185
R1592 GNDA.n120 GNDA.n94 185
R1593 GNDA.n129 GNDA.n128 185
R1594 GNDA.n566 GNDA.n522 185
R1595 GNDA.t314 GNDA.n522 185
R1596 GNDA.n568 GNDA.n567 185
R1597 GNDA.n570 GNDA.n569 185
R1598 GNDA.n572 GNDA.n571 185
R1599 GNDA.n574 GNDA.n573 185
R1600 GNDA.n576 GNDA.n575 185
R1601 GNDA.n578 GNDA.n577 185
R1602 GNDA.n579 GNDA.n527 185
R1603 GNDA.t314 GNDA.n527 185
R1604 GNDA.n581 GNDA.n580 185
R1605 GNDA.n565 GNDA.n564 185
R1606 GNDA.n563 GNDA.n562 185
R1607 GNDA.n561 GNDA.n560 185
R1608 GNDA.n559 GNDA.n558 185
R1609 GNDA.n557 GNDA.n556 185
R1610 GNDA.n555 GNDA.n554 185
R1611 GNDA.n553 GNDA.n552 185
R1612 GNDA.n551 GNDA.n550 185
R1613 GNDA.n549 GNDA.n548 185
R1614 GNDA.n547 GNDA.n546 185
R1615 GNDA.n545 GNDA.n544 185
R1616 GNDA.n543 GNDA.n542 185
R1617 GNDA.n541 GNDA.n540 185
R1618 GNDA.n539 GNDA.n538 185
R1619 GNDA.n537 GNDA.n536 185
R1620 GNDA.n535 GNDA.n534 185
R1621 GNDA.n533 GNDA.n532 185
R1622 GNDA.n531 GNDA.n512 185
R1623 GNDA.n637 GNDA.n636 185
R1624 GNDA.n594 GNDA.n513 185
R1625 GNDA.n593 GNDA.n592 185
R1626 GNDA.n610 GNDA.n609 185
R1627 GNDA.n612 GNDA.n611 185
R1628 GNDA.n616 GNDA.n614 185
R1629 GNDA.n618 GNDA.n617 185
R1630 GNDA.n583 GNDA.n582 185
R1631 GNDA.n633 GNDA.n632 185
R1632 GNDA.n2118 GNDA.n2016 185
R1633 GNDA.n2121 GNDA.n2120 185
R1634 GNDA.n2043 GNDA.n2018 185
R1635 GNDA.n2046 GNDA.n2042 185
R1636 GNDA.n2051 GNDA.n2050 185
R1637 GNDA.n2054 GNDA.n2053 185
R1638 GNDA.n2040 GNDA.n2037 185
R1639 GNDA.n2059 GNDA.n2036 185
R1640 GNDA.n2067 GNDA.n2066 185
R1641 GNDA.n2240 GNDA.n2170 185
R1642 GNDA.t254 GNDA.n2170 185
R1643 GNDA.n2242 GNDA.n2241 185
R1644 GNDA.n2244 GNDA.n2243 185
R1645 GNDA.n2246 GNDA.n2245 185
R1646 GNDA.n2248 GNDA.n2247 185
R1647 GNDA.n2250 GNDA.n2249 185
R1648 GNDA.n2252 GNDA.n2251 185
R1649 GNDA.n2253 GNDA.n2175 185
R1650 GNDA.t254 GNDA.n2175 185
R1651 GNDA.n2254 GNDA.n2179 185
R1652 GNDA.n2239 GNDA.n2238 185
R1653 GNDA.n2237 GNDA.n2236 185
R1654 GNDA.n2235 GNDA.n2234 185
R1655 GNDA.n2233 GNDA.n2232 185
R1656 GNDA.n2231 GNDA.n2230 185
R1657 GNDA.n2229 GNDA.n2228 185
R1658 GNDA.n2227 GNDA.n2226 185
R1659 GNDA.n2225 GNDA.n2224 185
R1660 GNDA.n2223 GNDA.n2222 185
R1661 GNDA.n2221 GNDA.n2220 185
R1662 GNDA.n2219 GNDA.n2218 185
R1663 GNDA.n2217 GNDA.n2216 185
R1664 GNDA.n2215 GNDA.n2214 185
R1665 GNDA.n2213 GNDA.n2212 185
R1666 GNDA.n2211 GNDA.n2210 185
R1667 GNDA.n2209 GNDA.n2208 185
R1668 GNDA.n2207 GNDA.n2206 185
R1669 GNDA.n2160 GNDA.n2157 185
R1670 GNDA.n727 GNDA.n675 185
R1671 GNDA.n675 GNDA.t253 185
R1672 GNDA.n726 GNDA.n725 185
R1673 GNDA.n723 GNDA.n676 185
R1674 GNDA.n722 GNDA.n677 185
R1675 GNDA.n720 GNDA.n719 185
R1676 GNDA.n718 GNDA.n678 185
R1677 GNDA.n717 GNDA.n716 185
R1678 GNDA.n714 GNDA.n679 185
R1679 GNDA.n714 GNDA.t253 185
R1680 GNDA.n713 GNDA.n680 185
R1681 GNDA.n729 GNDA.n728 185
R1682 GNDA.n731 GNDA.n673 185
R1683 GNDA.n733 GNDA.n732 185
R1684 GNDA.n734 GNDA.n672 185
R1685 GNDA.n736 GNDA.n735 185
R1686 GNDA.n738 GNDA.n670 185
R1687 GNDA.n740 GNDA.n739 185
R1688 GNDA.n741 GNDA.n669 185
R1689 GNDA.n743 GNDA.n742 185
R1690 GNDA.n745 GNDA.n668 185
R1691 GNDA.n747 GNDA.n746 185
R1692 GNDA.n749 GNDA.n748 185
R1693 GNDA.n752 GNDA.n751 185
R1694 GNDA.n753 GNDA.n666 185
R1695 GNDA.n755 GNDA.n754 185
R1696 GNDA.n757 GNDA.n665 185
R1697 GNDA.n759 GNDA.n758 185
R1698 GNDA.n761 GNDA.n760 185
R1699 GNDA.n762 GNDA.n659 185
R1700 GNDA.n765 GNDA.n764 185
R1701 GNDA.n688 GNDA.n661 185
R1702 GNDA.n691 GNDA.n687 185
R1703 GNDA.n696 GNDA.n695 185
R1704 GNDA.n699 GNDA.n698 185
R1705 GNDA.n685 GNDA.n682 185
R1706 GNDA.n704 GNDA.n681 185
R1707 GNDA.n711 GNDA.n710 185
R1708 GNDA.n2265 GNDA.n2264 185
R1709 GNDA.n2185 GNDA.n2161 185
R1710 GNDA.n2184 GNDA.n2183 185
R1711 GNDA.n2192 GNDA.n2191 185
R1712 GNDA.n2190 GNDA.n2182 185
R1713 GNDA.n2199 GNDA.n2198 185
R1714 GNDA.n2197 GNDA.n2181 185
R1715 GNDA.n2204 GNDA.n2180 185
R1716 GNDA.n2261 GNDA.n2260 185
R1717 GNDA.n1404 GNDA.n1357 185
R1718 GNDA.t280 GNDA.n1357 185
R1719 GNDA.n1406 GNDA.n1405 185
R1720 GNDA.n1408 GNDA.n1407 185
R1721 GNDA.n1410 GNDA.n1409 185
R1722 GNDA.n1412 GNDA.n1411 185
R1723 GNDA.n1414 GNDA.n1413 185
R1724 GNDA.n1416 GNDA.n1415 185
R1725 GNDA.n1417 GNDA.n1362 185
R1726 GNDA.t280 GNDA.n1362 185
R1727 GNDA.n1418 GNDA.n1366 185
R1728 GNDA.n1403 GNDA.n1402 185
R1729 GNDA.n1401 GNDA.n1400 185
R1730 GNDA.n1399 GNDA.n1398 185
R1731 GNDA.n1397 GNDA.n1396 185
R1732 GNDA.n1395 GNDA.n1394 185
R1733 GNDA.n1393 GNDA.n1392 185
R1734 GNDA.n1391 GNDA.n1390 185
R1735 GNDA.n1389 GNDA.n1388 185
R1736 GNDA.n1387 GNDA.n1386 185
R1737 GNDA.n1385 GNDA.n1384 185
R1738 GNDA.n1383 GNDA.n1382 185
R1739 GNDA.n1381 GNDA.n1380 185
R1740 GNDA.n1379 GNDA.n1378 185
R1741 GNDA.n1377 GNDA.n1376 185
R1742 GNDA.n1375 GNDA.n1374 185
R1743 GNDA.n1373 GNDA.n1372 185
R1744 GNDA.n1371 GNDA.n1370 185
R1745 GNDA.n1369 GNDA.n1347 185
R1746 GNDA.n1523 GNDA.n1522 185
R1747 GNDA.n1426 GNDA.n1348 185
R1748 GNDA.n1429 GNDA.n1428 185
R1749 GNDA.n1432 GNDA.n1431 185
R1750 GNDA.n1430 GNDA.n1422 185
R1751 GNDA.n1441 GNDA.n1440 185
R1752 GNDA.n1443 GNDA.n1442 185
R1753 GNDA.n1444 GNDA.n1367 185
R1754 GNDA.n1519 GNDA.n1518 185
R1755 GNDA.n1764 GNDA.n1659 185
R1756 GNDA.n1767 GNDA.n1766 185
R1757 GNDA.n1689 GNDA.n1661 185
R1758 GNDA.n1688 GNDA.n1687 185
R1759 GNDA.n1698 GNDA.n1697 185
R1760 GNDA.n1700 GNDA.n1684 185
R1761 GNDA.n1703 GNDA.n1702 185
R1762 GNDA.n1680 GNDA.n1679 185
R1763 GNDA.n1713 GNDA.n1712 185
R1764 GNDA.n1575 GNDA.n1574 185
R1765 GNDA.n1318 GNDA.n1240 185
R1766 GNDA.n1321 GNDA.n1320 185
R1767 GNDA.n1324 GNDA.n1323 185
R1768 GNDA.n1322 GNDA.n1314 185
R1769 GNDA.n1333 GNDA.n1332 185
R1770 GNDA.n1335 GNDA.n1334 185
R1771 GNDA.n1336 GNDA.n1259 185
R1772 GNDA.n1571 GNDA.n1570 185
R1773 GNDA.n334 GNDA.n228 185
R1774 GNDA.n337 GNDA.n336 185
R1775 GNDA.n258 GNDA.n231 185
R1776 GNDA.n259 GNDA.n255 185
R1777 GNDA.n268 GNDA.n267 185
R1778 GNDA.n270 GNDA.n253 185
R1779 GNDA.n273 GNDA.n272 185
R1780 GNDA.n274 GNDA.n248 185
R1781 GNDA.n283 GNDA.n282 185
R1782 GNDA.n1156 GNDA.n1155 182.4
R1783 GNDA.n1048 GNDA.n973 182.4
R1784 GNDA.n1151 GNDA.n1150 179.363
R1785 GNDA.n1006 GNDA.n1005 176.543
R1786 GNDA.n1005 GNDA.n996 176.543
R1787 GNDA.n1216 GNDA.n1215 176
R1788 GNDA.n1217 GNDA.n1216 176
R1789 GNDA.n1178 GNDA.n863 176
R1790 GNDA.n976 GNDA.n970 176
R1791 GNDA.t21 GNDA.n851 175.864
R1792 GNDA.n2400 GNDA.n2398 175.546
R1793 GNDA.n2404 GNDA.n66 175.546
R1794 GNDA.n2408 GNDA.n2406 175.546
R1795 GNDA.n2412 GNDA.n64 175.546
R1796 GNDA.n2415 GNDA.n2414 175.546
R1797 GNDA.n2437 GNDA.n51 175.546
R1798 GNDA.n2437 GNDA.n54 175.546
R1799 GNDA.n2433 GNDA.n54 175.546
R1800 GNDA.n2433 GNDA.n56 175.546
R1801 GNDA.n2429 GNDA.n56 175.546
R1802 GNDA.n2429 GNDA.n58 175.546
R1803 GNDA.n2425 GNDA.n58 175.546
R1804 GNDA.n2425 GNDA.n60 175.546
R1805 GNDA.n2421 GNDA.n60 175.546
R1806 GNDA.n2421 GNDA.n2419 175.546
R1807 GNDA.n340 GNDA.n339 175.546
R1808 GNDA.n261 GNDA.n257 175.546
R1809 GNDA.n265 GNDA.n263 175.546
R1810 GNDA.n276 GNDA.n251 175.546
R1811 GNDA.n280 GNDA.n278 175.546
R1812 GNDA.n348 GNDA.n347 175.546
R1813 GNDA.n352 GNDA.n351 175.546
R1814 GNDA.n354 GNDA.n353 175.546
R1815 GNDA.n359 GNDA.n358 175.546
R1816 GNDA.n361 GNDA.n360 175.546
R1817 GNDA.n1587 GNDA.n1583 175.546
R1818 GNDA.n1590 GNDA.n1589 175.546
R1819 GNDA.n1596 GNDA.n1592 175.546
R1820 GNDA.n1599 GNDA.n1598 175.546
R1821 GNDA.n1603 GNDA.n1601 175.546
R1822 GNDA.n2294 GNDA.n2293 175.546
R1823 GNDA.n2291 GNDA.n2274 175.546
R1824 GNDA.n2287 GNDA.n2286 175.546
R1825 GNDA.n2284 GNDA.n2277 175.546
R1826 GNDA.n2280 GNDA.n2279 175.546
R1827 GNDA.n1561 GNDA.n1560 175.546
R1828 GNDA.n1558 GNDA.n1534 175.546
R1829 GNDA.n1554 GNDA.n1553 175.546
R1830 GNDA.n1551 GNDA.n1541 175.546
R1831 GNDA.n1547 GNDA.n1546 175.546
R1832 GNDA.n1577 GNDA.n1236 175.546
R1833 GNDA.n1326 GNDA.n1317 175.546
R1834 GNDA.n1330 GNDA.n1328 175.546
R1835 GNDA.n1338 GNDA.n1312 175.546
R1836 GNDA.n1568 GNDA.n1340 175.546
R1837 GNDA.n1916 GNDA.n490 175.546
R1838 GNDA.n1916 GNDA.n491 175.546
R1839 GNDA.n1912 GNDA.n491 175.546
R1840 GNDA.n1912 GNDA.n1889 175.546
R1841 GNDA.n1908 GNDA.n1889 175.546
R1842 GNDA.n1908 GNDA.n1891 175.546
R1843 GNDA.n1904 GNDA.n1891 175.546
R1844 GNDA.n1904 GNDA.n1893 175.546
R1845 GNDA.n1900 GNDA.n1893 175.546
R1846 GNDA.n1900 GNDA.n1897 175.546
R1847 GNDA.n1942 GNDA.n462 175.546
R1848 GNDA.n1946 GNDA.n462 175.546
R1849 GNDA.n1946 GNDA.n460 175.546
R1850 GNDA.n1951 GNDA.n460 175.546
R1851 GNDA.n1951 GNDA.n458 175.546
R1852 GNDA.n1955 GNDA.n458 175.546
R1853 GNDA.n1955 GNDA.n457 175.546
R1854 GNDA.n1959 GNDA.n457 175.546
R1855 GNDA.n1959 GNDA.n455 175.546
R1856 GNDA.n1964 GNDA.n455 175.546
R1857 GNDA.n1964 GNDA.n448 175.546
R1858 GNDA.n2003 GNDA.n2002 175.546
R1859 GNDA.n2000 GNDA.n431 175.546
R1860 GNDA.n1996 GNDA.n1995 175.546
R1861 GNDA.n1993 GNDA.n439 175.546
R1862 GNDA.n1989 GNDA.n1988 175.546
R1863 GNDA.n639 GNDA.n508 175.546
R1864 GNDA.n639 GNDA.n509 175.546
R1865 GNDA.n596 GNDA.n509 175.546
R1866 GNDA.n607 GNDA.n596 175.546
R1867 GNDA.n607 GNDA.n597 175.546
R1868 GNDA.n597 GNDA.n590 175.546
R1869 GNDA.n620 GNDA.n590 175.546
R1870 GNDA.n620 GNDA.n584 175.546
R1871 GNDA.n629 GNDA.n584 175.546
R1872 GNDA.n629 GNDA.n411 175.546
R1873 GNDA.n2131 GNDA.n411 175.546
R1874 GNDA.n1859 GNDA.n650 175.546
R1875 GNDA.n1869 GNDA.n650 175.546
R1876 GNDA.n1869 GNDA.n473 175.546
R1877 GNDA.n1931 GNDA.n473 175.546
R1878 GNDA.n1931 GNDA.n474 175.546
R1879 GNDA.n1927 GNDA.n474 175.546
R1880 GNDA.n1927 GNDA.n477 175.546
R1881 GNDA.n500 GNDA.n477 175.546
R1882 GNDA.n502 GNDA.n500 175.546
R1883 GNDA.n502 GNDA.n497 175.546
R1884 GNDA.n767 GNDA.n653 175.546
R1885 GNDA.n689 GNDA.n658 175.546
R1886 GNDA.n693 GNDA.n692 175.546
R1887 GNDA.n702 GNDA.n701 175.546
R1888 GNDA.n708 GNDA.n707 175.546
R1889 GNDA.n2152 GNDA.n2151 175.546
R1890 GNDA.n2149 GNDA.n396 175.546
R1891 GNDA.n2145 GNDA.n2144 175.546
R1892 GNDA.n2142 GNDA.n402 175.546
R1893 GNDA.n2138 GNDA.n2137 175.546
R1894 GNDA.n641 GNDA.n498 175.546
R1895 GNDA.n641 GNDA.n506 175.546
R1896 GNDA.n600 GNDA.n506 175.546
R1897 GNDA.n600 GNDA.n599 175.546
R1898 GNDA.n604 GNDA.n599 175.546
R1899 GNDA.n604 GNDA.n588 175.546
R1900 GNDA.n622 GNDA.n588 175.546
R1901 GNDA.n622 GNDA.n586 175.546
R1902 GNDA.n627 GNDA.n586 175.546
R1903 GNDA.n627 GNDA.n408 175.546
R1904 GNDA.n2133 GNDA.n408 175.546
R1905 GNDA.n2123 GNDA.n2009 175.546
R1906 GNDA.n2044 GNDA.n2014 175.546
R1907 GNDA.n2048 GNDA.n2047 175.546
R1908 GNDA.n2057 GNDA.n2056 175.546
R1909 GNDA.n2064 GNDA.n2063 175.546
R1910 GNDA.n2005 GNDA.n428 175.546
R1911 GNDA.n434 GNDA.n433 175.546
R1912 GNDA.n440 GNDA.n436 175.546
R1913 GNDA.n443 GNDA.n442 175.546
R1914 GNDA.n449 GNDA.n445 175.546
R1915 GNDA.n1979 GNDA.n453 175.546
R1916 GNDA.n1979 GNDA.n1969 175.546
R1917 GNDA.n1975 GNDA.n1969 175.546
R1918 GNDA.n1975 GNDA.n1972 175.546
R1919 GNDA.n1972 GNDA.n8 175.546
R1920 GNDA.n2508 GNDA.n8 175.546
R1921 GNDA.n2508 GNDA.n9 175.546
R1922 GNDA.n2504 GNDA.n9 175.546
R1923 GNDA.n2504 GNDA.n11 175.546
R1924 GNDA.n2500 GNDA.n11 175.546
R1925 GNDA.n2500 GNDA.n2497 175.546
R1926 GNDA.n2386 GNDA.n2385 175.546
R1927 GNDA.n2383 GNDA.n196 175.546
R1928 GNDA.n2379 GNDA.n2378 175.546
R1929 GNDA.n2376 GNDA.n202 175.546
R1930 GNDA.n2372 GNDA.n2371 175.546
R1931 GNDA.n2489 GNDA.n17 175.546
R1932 GNDA.n2489 GNDA.n19 175.546
R1933 GNDA.n2485 GNDA.n19 175.546
R1934 GNDA.n2485 GNDA.n22 175.546
R1935 GNDA.n2481 GNDA.n22 175.546
R1936 GNDA.n2481 GNDA.n23 175.546
R1937 GNDA.n2477 GNDA.n23 175.546
R1938 GNDA.n2477 GNDA.n25 175.546
R1939 GNDA.n2473 GNDA.n25 175.546
R1940 GNDA.n2473 GNDA.n28 175.546
R1941 GNDA.n2469 GNDA.n28 175.546
R1942 GNDA.n2448 GNDA.n39 175.546
R1943 GNDA.n2448 GNDA.n37 175.546
R1944 GNDA.n2453 GNDA.n37 175.546
R1945 GNDA.n2453 GNDA.n35 175.546
R1946 GNDA.n2457 GNDA.n35 175.546
R1947 GNDA.n2457 GNDA.n34 175.546
R1948 GNDA.n2461 GNDA.n34 175.546
R1949 GNDA.n2461 GNDA.n32 175.546
R1950 GNDA.n2465 GNDA.n32 175.546
R1951 GNDA.n2465 GNDA.n30 175.546
R1952 GNDA.n186 GNDA.n185 175.546
R1953 GNDA.n107 GNDA.n103 175.546
R1954 GNDA.n111 GNDA.n109 175.546
R1955 GNDA.n122 GNDA.n97 175.546
R1956 GNDA.n126 GNDA.n124 175.546
R1957 GNDA.n2361 GNDA.n2360 175.546
R1958 GNDA.n198 GNDA.n197 175.546
R1959 GNDA.n2364 GNDA.n199 175.546
R1960 GNDA.n204 GNDA.n203 175.546
R1961 GNDA.n2369 GNDA.n205 175.546
R1962 GNDA.n419 GNDA.n418 175.546
R1963 GNDA.n398 GNDA.n397 175.546
R1964 GNDA.n422 GNDA.n399 175.546
R1965 GNDA.n404 GNDA.n403 175.546
R1966 GNDA.n425 GNDA.n405 175.546
R1967 GNDA.n2306 GNDA.n2305 175.546
R1968 GNDA.n2310 GNDA.n2309 175.546
R1969 GNDA.n2314 GNDA.n2313 175.546
R1970 GNDA.n2316 GNDA.n369 175.546
R1971 GNDA.n2321 GNDA.n364 175.546
R1972 GNDA.n2345 GNDA.n2344 175.546
R1973 GNDA.n2342 GNDA.n350 175.546
R1974 GNDA.n2338 GNDA.n2337 175.546
R1975 GNDA.n2335 GNDA.n357 175.546
R1976 GNDA.n2331 GNDA.n2330 175.546
R1977 GNDA.n2158 GNDA.n388 175.546
R1978 GNDA.n2188 GNDA.n2187 175.546
R1979 GNDA.n2195 GNDA.n2194 175.546
R1980 GNDA.n2202 GNDA.n2201 175.546
R1981 GNDA.n2258 GNDA.n2257 175.546
R1982 GNDA.n1531 GNDA.n1530 175.546
R1983 GNDA.n1536 GNDA.n1535 175.546
R1984 GNDA.n1538 GNDA.n1537 175.546
R1985 GNDA.n1543 GNDA.n1542 175.546
R1986 GNDA.n1544 GNDA.n217 175.546
R1987 GNDA.n1471 GNDA.n1468 175.546
R1988 GNDA.n1475 GNDA.n1473 175.546
R1989 GNDA.n1479 GNDA.n1464 175.546
R1990 GNDA.n1483 GNDA.n1481 175.546
R1991 GNDA.n1487 GNDA.n1462 175.546
R1992 GNDA.n1510 GNDA.n1451 175.546
R1993 GNDA.n1506 GNDA.n1451 175.546
R1994 GNDA.n1506 GNDA.n1454 175.546
R1995 GNDA.n1502 GNDA.n1454 175.546
R1996 GNDA.n1502 GNDA.n1500 175.546
R1997 GNDA.n1500 GNDA.n1456 175.546
R1998 GNDA.n1496 GNDA.n1456 175.546
R1999 GNDA.n1496 GNDA.n1458 175.546
R2000 GNDA.n1492 GNDA.n1458 175.546
R2001 GNDA.n1492 GNDA.n1490 175.546
R2002 GNDA.n1525 GNDA.n1344 175.546
R2003 GNDA.n1434 GNDA.n1425 175.546
R2004 GNDA.n1438 GNDA.n1436 175.546
R2005 GNDA.n1446 GNDA.n1420 175.546
R2006 GNDA.n1516 GNDA.n1448 175.546
R2007 GNDA.n1651 GNDA.n1622 175.546
R2008 GNDA.n1647 GNDA.n1622 175.546
R2009 GNDA.n1647 GNDA.n1623 175.546
R2010 GNDA.n1643 GNDA.n1623 175.546
R2011 GNDA.n1643 GNDA.n1625 175.546
R2012 GNDA.n1639 GNDA.n1625 175.546
R2013 GNDA.n1639 GNDA.n1629 175.546
R2014 GNDA.n1635 GNDA.n1629 175.546
R2015 GNDA.n1635 GNDA.n1632 175.546
R2016 GNDA.n1632 GNDA.n1613 175.546
R2017 GNDA.n1769 GNDA.n1655 175.546
R2018 GNDA.n1691 GNDA.n1657 175.546
R2019 GNDA.n1694 GNDA.n1691 175.546
R2020 GNDA.n1694 GNDA.n1683 175.546
R2021 GNDA.n1705 GNDA.n1683 175.546
R2022 GNDA.n1705 GNDA.n1681 175.546
R2023 GNDA.n1709 GNDA.n1681 175.546
R2024 GNDA.n1709 GNDA.n1231 175.546
R2025 GNDA.n1833 GNDA.n1231 175.546
R2026 GNDA.n1828 GNDA.n1827 175.546
R2027 GNDA.n1825 GNDA.n1586 175.546
R2028 GNDA.n1821 GNDA.n1820 175.546
R2029 GNDA.n1818 GNDA.n1595 175.546
R2030 GNDA.n1814 GNDA.n1813 175.546
R2031 GNDA.n1791 GNDA.n1790 175.546
R2032 GNDA.n1795 GNDA.n1794 175.546
R2033 GNDA.n1799 GNDA.n1798 175.546
R2034 GNDA.n1801 GNDA.n1611 175.546
R2035 GNDA.n1806 GNDA.n1606 175.546
R2036 GNDA.n1228 GNDA.n1227 175.5
R2037 GNDA.n2272 GNDA.n2271 173.881
R2038 GNDA.n2125 GNDA.t227 172.876
R2039 GNDA.n769 GNDA.t225 172.876
R2040 GNDA.n2323 GNDA.t227 172.615
R2041 GNDA.n1808 GNDA.t225 172.615
R2042 GNDA.n1152 GNDA.n1151 171.817
R2043 GNDA.n2273 GNDA.n2272 171.624
R2044 GNDA.n1656 GNDA.n776 170.543
R2045 GNDA.n1204 GNDA.n849 169.232
R2046 GNDA.n1150 GNDA.n881 164.906
R2047 GNDA.n334 GNDA.n333 163.333
R2048 GNDA.n1574 GNDA.n1239 163.333
R2049 GNDA.n1764 GNDA.n1763 163.333
R2050 GNDA.n2118 GNDA.n2117 163.333
R2051 GNDA.n180 GNDA.n179 163.333
R2052 GNDA.n636 GNDA.n512 163.333
R2053 GNDA.n2264 GNDA.n2160 163.333
R2054 GNDA.n762 GNDA.n761 163.333
R2055 GNDA.n1522 GNDA.n1347 163.333
R2056 GNDA.n1949 GNDA.t225 162.964
R2057 GNDA.n2482 GNDA.t227 162.964
R2058 GNDA.n841 GNDA.t295 160.725
R2059 GNDA.n840 GNDA.t275 160.725
R2060 GNDA.n828 GNDA.t230 160.725
R2061 GNDA.n829 GNDA.t283 160.725
R2062 GNDA.n1199 GNDA.t263 160.725
R2063 GNDA.n844 GNDA.t289 160.725
R2064 GNDA.n945 GNDA.n944 160
R2065 GNDA.n940 GNDA.n935 160
R2066 GNDA.n1100 GNDA.n1099 160
R2067 GNDA.n788 GNDA.t87 157.555
R2068 GNDA.n787 GNDA.t96 157.555
R2069 GNDA.n1094 GNDA.n1093 156.8
R2070 GNDA.n1086 GNDA.n1085 153.601
R2071 GNDA.n1148 GNDA.n885 153.601
R2072 GNDA.n876 GNDA.n872 153.601
R2073 GNDA.n1050 GNDA.n969 153.601
R2074 GNDA.n811 GNDA.t46 153.294
R2075 GNDA.n862 GNDA.t260 152.994
R2076 GNDA.n1153 GNDA.t246 152.994
R2077 GNDA.n972 GNDA.t268 152.994
R2078 GNDA.n975 GNDA.t257 152.994
R2079 GNDA.n1091 GNDA.n962 150.4
R2080 GNDA.n1139 GNDA.n1138 150.4
R2081 GNDA.n1019 GNDA.n1018 150.329
R2082 GNDA.n1018 GNDA.n1016 150.329
R2083 GNDA.n336 GNDA.n231 150
R2084 GNDA.n268 GNDA.n255 150
R2085 GNDA.n272 GNDA.n270 150
R2086 GNDA.n283 GNDA.n248 150
R2087 GNDA.n331 GNDA.n232 150
R2088 GNDA.n327 GNDA.n325 150
R2089 GNDA.n323 GNDA.n234 150
R2090 GNDA.n319 GNDA.n317 150
R2091 GNDA.n315 GNDA.n236 150
R2092 GNDA.n311 GNDA.n310 150
R2093 GNDA.n308 GNDA.n239 150
R2094 GNDA.n304 GNDA.n303 150
R2095 GNDA.n286 GNDA.n285 150
R2096 GNDA.n288 GNDA.n286 150
R2097 GNDA.n292 GNDA.n245 150
R2098 GNDA.n295 GNDA.n294 150
R2099 GNDA.n297 GNDA.n242 150
R2100 GNDA.n1320 GNDA.n1240 150
R2101 GNDA.n1323 GNDA.n1322 150
R2102 GNDA.n1334 GNDA.n1333 150
R2103 GNDA.n1571 GNDA.n1259 150
R2104 GNDA.n1264 GNDA.n1263 150
R2105 GNDA.n1268 GNDA.n1267 150
R2106 GNDA.n1272 GNDA.n1271 150
R2107 GNDA.n1276 GNDA.n1275 150
R2108 GNDA.n1280 GNDA.n1279 150
R2109 GNDA.n1284 GNDA.n1283 150
R2110 GNDA.n1288 GNDA.n1287 150
R2111 GNDA.n1292 GNDA.n1291 150
R2112 GNDA.n1258 GNDA.n1254 150
R2113 GNDA.n1307 GNDA.n1254 150
R2114 GNDA.n1305 GNDA.n1304 150
R2115 GNDA.n1301 GNDA.n1300 150
R2116 GNDA.n1297 GNDA.n1249 150
R2117 GNDA.n1766 GNDA.n1661 150
R2118 GNDA.n1698 GNDA.n1687 150
R2119 GNDA.n1702 GNDA.n1700 150
R2120 GNDA.n1713 GNDA.n1679 150
R2121 GNDA.n1760 GNDA.n1759 150
R2122 GNDA.n1757 GNDA.n1664 150
R2123 GNDA.n1753 GNDA.n1751 150
R2124 GNDA.n1748 GNDA.n1747 150
R2125 GNDA.n1745 GNDA.n1667 150
R2126 GNDA.n1741 GNDA.n1740 150
R2127 GNDA.n1738 GNDA.n1670 150
R2128 GNDA.n1734 GNDA.n1733 150
R2129 GNDA.n1716 GNDA.n1715 150
R2130 GNDA.n1718 GNDA.n1716 150
R2131 GNDA.n1722 GNDA.n1676 150
R2132 GNDA.n1725 GNDA.n1724 150
R2133 GNDA.n1727 GNDA.n1673 150
R2134 GNDA.n2120 GNDA.n2018 150
R2135 GNDA.n2051 GNDA.n2042 150
R2136 GNDA.n2053 GNDA.n2040 150
R2137 GNDA.n2067 GNDA.n2036 150
R2138 GNDA.n2114 GNDA.n2113 150
R2139 GNDA.n2111 GNDA.n2021 150
R2140 GNDA.n2107 GNDA.n2105 150
R2141 GNDA.n2102 GNDA.n2101 150
R2142 GNDA.n2099 GNDA.n2024 150
R2143 GNDA.n2095 GNDA.n2094 150
R2144 GNDA.n2092 GNDA.n2027 150
R2145 GNDA.n2088 GNDA.n2087 150
R2146 GNDA.n2070 GNDA.n2069 150
R2147 GNDA.n2072 GNDA.n2070 150
R2148 GNDA.n2076 GNDA.n2033 150
R2149 GNDA.n2079 GNDA.n2078 150
R2150 GNDA.n2081 GNDA.n2030 150
R2151 GNDA.n182 GNDA.n77 150
R2152 GNDA.n114 GNDA.n101 150
R2153 GNDA.n118 GNDA.n116 150
R2154 GNDA.n129 GNDA.n94 150
R2155 GNDA.n177 GNDA.n78 150
R2156 GNDA.n173 GNDA.n171 150
R2157 GNDA.n169 GNDA.n80 150
R2158 GNDA.n165 GNDA.n163 150
R2159 GNDA.n161 GNDA.n82 150
R2160 GNDA.n157 GNDA.n156 150
R2161 GNDA.n154 GNDA.n85 150
R2162 GNDA.n150 GNDA.n149 150
R2163 GNDA.n132 GNDA.n131 150
R2164 GNDA.n134 GNDA.n132 150
R2165 GNDA.n138 GNDA.n91 150
R2166 GNDA.n141 GNDA.n140 150
R2167 GNDA.n143 GNDA.n88 150
R2168 GNDA.n592 GNDA.n513 150
R2169 GNDA.n611 GNDA.n610 150
R2170 GNDA.n617 GNDA.n616 150
R2171 GNDA.n633 GNDA.n582 150
R2172 GNDA.n534 GNDA.n533 150
R2173 GNDA.n538 GNDA.n537 150
R2174 GNDA.n542 GNDA.n541 150
R2175 GNDA.n546 GNDA.n545 150
R2176 GNDA.n550 GNDA.n549 150
R2177 GNDA.n554 GNDA.n553 150
R2178 GNDA.n558 GNDA.n557 150
R2179 GNDA.n562 GNDA.n561 150
R2180 GNDA.n581 GNDA.n527 150
R2181 GNDA.n577 GNDA.n527 150
R2182 GNDA.n575 GNDA.n574 150
R2183 GNDA.n571 GNDA.n570 150
R2184 GNDA.n567 GNDA.n522 150
R2185 GNDA.n2183 GNDA.n2161 150
R2186 GNDA.n2191 GNDA.n2190 150
R2187 GNDA.n2198 GNDA.n2197 150
R2188 GNDA.n2261 GNDA.n2180 150
R2189 GNDA.n2208 GNDA.n2207 150
R2190 GNDA.n2212 GNDA.n2211 150
R2191 GNDA.n2216 GNDA.n2215 150
R2192 GNDA.n2220 GNDA.n2219 150
R2193 GNDA.n2224 GNDA.n2223 150
R2194 GNDA.n2228 GNDA.n2227 150
R2195 GNDA.n2232 GNDA.n2231 150
R2196 GNDA.n2236 GNDA.n2235 150
R2197 GNDA.n2179 GNDA.n2175 150
R2198 GNDA.n2251 GNDA.n2175 150
R2199 GNDA.n2249 GNDA.n2248 150
R2200 GNDA.n2245 GNDA.n2244 150
R2201 GNDA.n2241 GNDA.n2170 150
R2202 GNDA.n764 GNDA.n661 150
R2203 GNDA.n696 GNDA.n687 150
R2204 GNDA.n698 GNDA.n685 150
R2205 GNDA.n711 GNDA.n681 150
R2206 GNDA.n758 GNDA.n757 150
R2207 GNDA.n755 GNDA.n666 150
R2208 GNDA.n751 GNDA.n749 150
R2209 GNDA.n746 GNDA.n745 150
R2210 GNDA.n743 GNDA.n669 150
R2211 GNDA.n739 GNDA.n738 150
R2212 GNDA.n736 GNDA.n672 150
R2213 GNDA.n732 GNDA.n731 150
R2214 GNDA.n714 GNDA.n713 150
R2215 GNDA.n716 GNDA.n714 150
R2216 GNDA.n720 GNDA.n678 150
R2217 GNDA.n723 GNDA.n722 150
R2218 GNDA.n725 GNDA.n675 150
R2219 GNDA.n1428 GNDA.n1348 150
R2220 GNDA.n1431 GNDA.n1430 150
R2221 GNDA.n1442 GNDA.n1441 150
R2222 GNDA.n1519 GNDA.n1367 150
R2223 GNDA.n1372 GNDA.n1371 150
R2224 GNDA.n1376 GNDA.n1375 150
R2225 GNDA.n1380 GNDA.n1379 150
R2226 GNDA.n1384 GNDA.n1383 150
R2227 GNDA.n1388 GNDA.n1387 150
R2228 GNDA.n1392 GNDA.n1391 150
R2229 GNDA.n1396 GNDA.n1395 150
R2230 GNDA.n1400 GNDA.n1399 150
R2231 GNDA.n1366 GNDA.n1362 150
R2232 GNDA.n1415 GNDA.n1362 150
R2233 GNDA.n1413 GNDA.n1412 150
R2234 GNDA.n1409 GNDA.n1408 150
R2235 GNDA.n1405 GNDA.n1357 150
R2236 GNDA.n1207 GNDA.n1206 149.181
R2237 GNDA.n789 GNDA.t344 148.906
R2238 GNDA.n789 GNDA.t122 148.653
R2239 GNDA.n793 GNDA.n791 139.639
R2240 GNDA.n809 GNDA.n808 139.077
R2241 GNDA.n807 GNDA.n806 139.077
R2242 GNDA.n805 GNDA.n804 139.077
R2243 GNDA.n803 GNDA.n802 139.077
R2244 GNDA.n801 GNDA.n800 139.077
R2245 GNDA.n799 GNDA.n798 139.077
R2246 GNDA.n797 GNDA.n796 139.077
R2247 GNDA.n795 GNDA.n794 139.077
R2248 GNDA.n793 GNDA.n792 139.077
R2249 GNDA.n1185 GNDA.n849 131.625
R2250 GNDA.n1046 GNDA.t267 130.731
R2251 GNDA.t245 GNDA.n1158 130.731
R2252 GNDA.n1097 GNDA.n949 127.249
R2253 GNDA.n2396 GNDA.n68 126.782
R2254 GNDA.n2299 GNDA.n377 126.782
R2255 GNDA.n1942 GNDA.n464 126.782
R2256 GNDA.n645 GNDA.n498 126.782
R2257 GNDA.n1983 GNDA.n453 126.782
R2258 GNDA.n2493 GNDA.n17 126.782
R2259 GNDA.n2302 GNDA.n2301 126.782
R2260 GNDA.n1466 GNDA.n218 126.782
R2261 GNDA.n1787 GNDA.n1786 126.782
R2262 GNDA.n1837 GNDA.n1228 125.356
R2263 GNDA.n2350 GNDA.n344 124.832
R2264 GNDA.n1580 GNDA.n1579 124.832
R2265 GNDA.n508 GNDA.n494 124.832
R2266 GNDA.n772 GNDA.n771 124.832
R2267 GNDA.n2127 GNDA.n2008 124.832
R2268 GNDA.n2391 GNDA.n190 124.832
R2269 GNDA.n2269 GNDA.n389 124.832
R2270 GNDA.n1528 GNDA.n1527 124.832
R2271 GNDA.n1773 GNDA.n1619 124.832
R2272 GNDA.n1043 GNDA.n1042 119.525
R2273 GNDA.n1176 GNDA.n867 119.525
R2274 GNDA.n837 GNDA.n836 118.4
R2275 GNDA.n839 GNDA.n838 118.4
R2276 GNDA.n1218 GNDA.n1217 118.4
R2277 GNDA.n1215 GNDA.n1214 118.4
R2278 GNDA.n1201 GNDA.n1200 118.4
R2279 GNDA.n1213 GNDA.n845 118.4
R2280 GNDA.n1027 GNDA.t67 115.79
R2281 GNDA.n1041 GNDA.t61 115.79
R2282 GNDA.n936 GNDA.t313 113.974
R2283 GNDA.n937 GNDA.t298 113.974
R2284 GNDA.n938 GNDA.t321 113.974
R2285 GNDA.n939 GNDA.t292 113.974
R2286 GNDA.n884 GNDA.t310 113.974
R2287 GNDA.n1104 GNDA.t304 113.974
R2288 GNDA.n1103 GNDA.t279 113.974
R2289 GNDA.n946 GNDA.t240 113.974
R2290 GNDA.n947 GNDA.t223 113.974
R2291 GNDA.n948 GNDA.t318 113.974
R2292 GNDA.n1693 GNDA.t225 113.624
R2293 GNDA.n2513 GNDA.t227 112.388
R2294 GNDA.n1035 GNDA.n1034 112.055
R2295 GNDA.n1113 GNDA.n922 108.8
R2296 GNDA.n924 GNDA.n919 108.8
R2297 GNDA.n1778 GNDA.n776 107.713
R2298 GNDA.n2367 GNDA.n0 14.555
R2299 GNDA.n1096 GNDA.t317 101.194
R2300 GNDA.n1967 GNDA.n394 99.6276
R2301 GNDA.n1064 GNDA.n1063 99.0842
R2302 GNDA.n1084 GNDA.n1083 99.0842
R2303 GNDA.n1082 GNDA.n1081 99.0842
R2304 GNDA.n1080 GNDA.n1079 99.0842
R2305 GNDA.n1078 GNDA.n1077 99.0842
R2306 GNDA.n1076 GNDA.n1075 99.0842
R2307 GNDA.n1074 GNDA.n1073 99.0842
R2308 GNDA.n1072 GNDA.n1071 99.0842
R2309 GNDA.n1070 GNDA.n1069 99.0842
R2310 GNDA.n1068 GNDA.n1067 99.0842
R2311 GNDA.n1066 GNDA.n1065 99.0842
R2312 GNDA.n889 GNDA.n888 99.0842
R2313 GNDA.n1175 GNDA.t54 97.1515
R2314 GNDA.n1183 GNDA.t17 97.1515
R2315 GNDA.n1143 GNDA.n1142 95.101
R2316 GNDA.n1058 GNDA.n963 95.101
R2317 GNDA.n1090 GNDA.t233 94.8842
R2318 GNDA.t243 GNDA.n953 94.8842
R2319 GNDA.n1140 GNDA.t272 94.8842
R2320 GNDA.n1087 GNDA.t307 94.8842
R2321 GNDA.n1060 GNDA.n1059 94.601
R2322 GNDA.n1145 GNDA.n1144 94.601
R2323 GNDA.n1169 GNDA.n1167 94.0176
R2324 GNDA.n1025 GNDA.n987 92.5103
R2325 GNDA.n1509 GNDA.n1452 91.8159
R2326 GNDA.n1509 GNDA.n1508 91.8159
R2327 GNDA.n1508 GNDA.n1507 91.8159
R2328 GNDA.n1507 GNDA.n1453 91.8159
R2329 GNDA.n1501 GNDA.n1453 91.8159
R2330 GNDA.n1499 GNDA.n1498 91.8159
R2331 GNDA.n1498 GNDA.n1497 91.8159
R2332 GNDA.n1497 GNDA.n1457 91.8159
R2333 GNDA.n1491 GNDA.n1457 91.8159
R2334 GNDA.n1491 GNDA.n48 91.8159
R2335 GNDA.n2442 GNDA.n49 91.8159
R2336 GNDA.n2436 GNDA.n49 91.8159
R2337 GNDA.n2436 GNDA.n2435 91.8159
R2338 GNDA.n2435 GNDA.n2434 91.8159
R2339 GNDA.n2434 GNDA.n55 91.8159
R2340 GNDA.n2428 GNDA.n2427 91.8159
R2341 GNDA.n2427 GNDA.n2426 91.8159
R2342 GNDA.n2426 GNDA.n59 91.8159
R2343 GNDA.n2420 GNDA.n59 91.8159
R2344 GNDA.n2420 GNDA.n43 91.8159
R2345 GNDA.n2443 GNDA.n38 91.8159
R2346 GNDA.n2449 GNDA.n38 91.8159
R2347 GNDA.n2450 GNDA.n2449 91.8159
R2348 GNDA.n2452 GNDA.n2450 91.8159
R2349 GNDA.n2452 GNDA.n2451 91.8159
R2350 GNDA.n2459 GNDA.n2458 91.8159
R2351 GNDA.n2460 GNDA.n2459 91.8159
R2352 GNDA.n2460 GNDA.n31 91.8159
R2353 GNDA.n2466 GNDA.n31 91.8159
R2354 GNDA.n2467 GNDA.n2466 91.8159
R2355 GNDA.n1097 GNDA.n1096 89.9494
R2356 GNDA.t67 GNDA.t90 89.644
R2357 GNDA.t176 GNDA.t136 89.644
R2358 GNDA.n1179 GNDA.n861 86.4005
R2359 GNDA.n1032 GNDA.n1031 86.4005
R2360 GNDA.n1841 GNDA.n814 85.2842
R2361 GNDA.n1193 GNDA.n1192 85.2842
R2362 GNDA.n2514 GNDA.n4 84.306
R2363 GNDA.n1835 GNDA.n394 83.2184
R2364 GNDA.t141 GNDA.t256 82.1737
R2365 GNDA.t48 GNDA.t22 82.1737
R2366 GNDA.t125 GNDA.t85 82.1737
R2367 GNDA.t105 GNDA.t97 82.1737
R2368 GNDA.t128 GNDA.t206 82.1737
R2369 GNDA.t209 GNDA.t83 82.1737
R2370 GNDA.t208 GNDA.t133 82.1737
R2371 GNDA.t15 GNDA.t259 82.1737
R2372 GNDA.n1777 GNDA.n1618 81.7969
R2373 GNDA.n1863 GNDA.n1862 81.7969
R2374 GNDA.n1884 GNDA.n1883 81.7969
R2375 GNDA.n1210 GNDA.n1209 81.482
R2376 GNDA.n1221 GNDA.n1220 81.482
R2377 GNDA.n2132 GNDA.t225 80.9821
R2378 GNDA.t285 GNDA.t182 78.4385
R2379 GNDA.t127 GNDA.t248 78.4385
R2380 GNDA.n1785 GNDA.n1614 77.7476
R2381 GNDA.n646 GNDA.n496 77.7476
R2382 GNDA.n2272 GNDA.t227 76.3879
R2383 GNDA.n2398 GNDA.n2397 76.3222
R2384 GNDA.n2399 GNDA.n66 76.3222
R2385 GNDA.n2406 GNDA.n2405 76.3222
R2386 GNDA.n2407 GNDA.n64 76.3222
R2387 GNDA.n2414 GNDA.n2413 76.3222
R2388 GNDA.n2418 GNDA.n62 76.3222
R2389 GNDA.n2441 GNDA.n2440 76.3222
R2390 GNDA.n344 GNDA.n226 76.3222
R2391 GNDA.n339 GNDA.n229 76.3222
R2392 GNDA.n262 GNDA.n261 76.3222
R2393 GNDA.n265 GNDA.n264 76.3222
R2394 GNDA.n277 GNDA.n276 76.3222
R2395 GNDA.n280 GNDA.n279 76.3222
R2396 GNDA.n2349 GNDA.n206 76.3222
R2397 GNDA.n348 GNDA.n207 76.3222
R2398 GNDA.n352 GNDA.n208 76.3222
R2399 GNDA.n354 GNDA.n209 76.3222
R2400 GNDA.n359 GNDA.n210 76.3222
R2401 GNDA.n2326 GNDA.n211 76.3222
R2402 GNDA.n1583 GNDA.n1582 76.3222
R2403 GNDA.n1589 GNDA.n1588 76.3222
R2404 GNDA.n1592 GNDA.n1591 76.3222
R2405 GNDA.n1598 GNDA.n1597 76.3222
R2406 GNDA.n1601 GNDA.n1600 76.3222
R2407 GNDA.n1602 GNDA.n376 76.3222
R2408 GNDA.n2294 GNDA.n382 76.3222
R2409 GNDA.n2292 GNDA.n2291 76.3222
R2410 GNDA.n2287 GNDA.n2276 76.3222
R2411 GNDA.n2285 GNDA.n2284 76.3222
R2412 GNDA.n2280 GNDA.n2278 76.3222
R2413 GNDA.n2355 GNDA.n222 76.3222
R2414 GNDA.n1561 GNDA.n1533 76.3222
R2415 GNDA.n1559 GNDA.n1558 76.3222
R2416 GNDA.n1554 GNDA.n1540 76.3222
R2417 GNDA.n1552 GNDA.n1551 76.3222
R2418 GNDA.n1547 GNDA.n1545 76.3222
R2419 GNDA.n2356 GNDA.n221 76.3222
R2420 GNDA.n1579 GNDA.n1578 76.3222
R2421 GNDA.n1316 GNDA.n1236 76.3222
R2422 GNDA.n1327 GNDA.n1326 76.3222
R2423 GNDA.n1330 GNDA.n1329 76.3222
R2424 GNDA.n1339 GNDA.n1338 76.3222
R2425 GNDA.n1568 GNDA.n1567 76.3222
R2426 GNDA.n492 GNDA.n490 76.3222
R2427 GNDA.n2003 GNDA.n430 76.3222
R2428 GNDA.n2001 GNDA.n2000 76.3222
R2429 GNDA.n1996 GNDA.n438 76.3222
R2430 GNDA.n1994 GNDA.n1993 76.3222
R2431 GNDA.n1989 GNDA.n447 76.3222
R2432 GNDA.n1987 GNDA.n1986 76.3222
R2433 GNDA.n1859 GNDA.n651 76.3222
R2434 GNDA.n771 GNDA.n770 76.3222
R2435 GNDA.n768 GNDA.n767 76.3222
R2436 GNDA.n689 GNDA.n657 76.3222
R2437 GNDA.n692 GNDA.n656 76.3222
R2438 GNDA.n702 GNDA.n655 76.3222
R2439 GNDA.n708 GNDA.n654 76.3222
R2440 GNDA.n2153 GNDA.n2152 76.3222
R2441 GNDA.n2150 GNDA.n2149 76.3222
R2442 GNDA.n2145 GNDA.n401 76.3222
R2443 GNDA.n2143 GNDA.n2142 76.3222
R2444 GNDA.n2138 GNDA.n407 76.3222
R2445 GNDA.n2136 GNDA.n2135 76.3222
R2446 GNDA.n2127 GNDA.n2126 76.3222
R2447 GNDA.n2124 GNDA.n2123 76.3222
R2448 GNDA.n2044 GNDA.n2013 76.3222
R2449 GNDA.n2047 GNDA.n2012 76.3222
R2450 GNDA.n2057 GNDA.n2011 76.3222
R2451 GNDA.n2064 GNDA.n2010 76.3222
R2452 GNDA.n2006 GNDA.n2005 76.3222
R2453 GNDA.n433 GNDA.n432 76.3222
R2454 GNDA.n436 GNDA.n435 76.3222
R2455 GNDA.n442 GNDA.n441 76.3222
R2456 GNDA.n445 GNDA.n444 76.3222
R2457 GNDA.n451 GNDA.n450 76.3222
R2458 GNDA.n2387 GNDA.n2386 76.3222
R2459 GNDA.n2384 GNDA.n2383 76.3222
R2460 GNDA.n2379 GNDA.n201 76.3222
R2461 GNDA.n2377 GNDA.n2376 76.3222
R2462 GNDA.n2372 GNDA.n2370 76.3222
R2463 GNDA.n2496 GNDA.n13 76.3222
R2464 GNDA.n2445 GNDA.n39 76.3222
R2465 GNDA.n190 GNDA.n72 76.3222
R2466 GNDA.n185 GNDA.n75 76.3222
R2467 GNDA.n108 GNDA.n107 76.3222
R2468 GNDA.n111 GNDA.n110 76.3222
R2469 GNDA.n123 GNDA.n122 76.3222
R2470 GNDA.n126 GNDA.n125 76.3222
R2471 GNDA.n2390 GNDA.n191 76.3222
R2472 GNDA.n2362 GNDA.n2361 76.3222
R2473 GNDA.n2363 GNDA.n198 76.3222
R2474 GNDA.n2365 GNDA.n2364 76.3222
R2475 GNDA.n2368 GNDA.n204 76.3222
R2476 GNDA.n2366 GNDA.n205 76.3222
R2477 GNDA.n2366 GNDA.n15 76.3222
R2478 GNDA.n2369 GNDA.n2368 76.3222
R2479 GNDA.n2365 GNDA.n203 76.3222
R2480 GNDA.n2363 GNDA.n199 76.3222
R2481 GNDA.n2362 GNDA.n197 76.3222
R2482 GNDA.n2360 GNDA.n191 76.3222
R2483 GNDA.n2371 GNDA.n13 76.3222
R2484 GNDA.n2370 GNDA.n202 76.3222
R2485 GNDA.n2378 GNDA.n2377 76.3222
R2486 GNDA.n201 GNDA.n196 76.3222
R2487 GNDA.n2385 GNDA.n2384 76.3222
R2488 GNDA.n2388 GNDA.n2387 76.3222
R2489 GNDA.n2126 GNDA.n2009 76.3222
R2490 GNDA.n2124 GNDA.n2014 76.3222
R2491 GNDA.n2048 GNDA.n2013 76.3222
R2492 GNDA.n2056 GNDA.n2012 76.3222
R2493 GNDA.n2063 GNDA.n2011 76.3222
R2494 GNDA.n2010 GNDA.n193 76.3222
R2495 GNDA.n418 GNDA.n417 76.3222
R2496 GNDA.n420 GNDA.n397 76.3222
R2497 GNDA.n421 GNDA.n399 76.3222
R2498 GNDA.n423 GNDA.n403 76.3222
R2499 GNDA.n424 GNDA.n405 76.3222
R2500 GNDA.n426 GNDA.n371 76.3222
R2501 GNDA.n2302 GNDA.n365 76.3222
R2502 GNDA.n2306 GNDA.n366 76.3222
R2503 GNDA.n2310 GNDA.n367 76.3222
R2504 GNDA.n2314 GNDA.n368 76.3222
R2505 GNDA.n2322 GNDA.n369 76.3222
R2506 GNDA.n2324 GNDA.n364 76.3222
R2507 GNDA.n2325 GNDA.n2324 76.3222
R2508 GNDA.n2322 GNDA.n2321 76.3222
R2509 GNDA.n2316 GNDA.n368 76.3222
R2510 GNDA.n2313 GNDA.n367 76.3222
R2511 GNDA.n2309 GNDA.n366 76.3222
R2512 GNDA.n2305 GNDA.n365 76.3222
R2513 GNDA.n2346 GNDA.n2345 76.3222
R2514 GNDA.n2343 GNDA.n2342 76.3222
R2515 GNDA.n2338 GNDA.n356 76.3222
R2516 GNDA.n2336 GNDA.n2335 76.3222
R2517 GNDA.n2331 GNDA.n363 76.3222
R2518 GNDA.n2329 GNDA.n2328 76.3222
R2519 GNDA.n2270 GNDA.n388 76.3222
R2520 GNDA.n2187 GNDA.n387 76.3222
R2521 GNDA.n2194 GNDA.n386 76.3222
R2522 GNDA.n2201 GNDA.n385 76.3222
R2523 GNDA.n2257 GNDA.n384 76.3222
R2524 GNDA.n383 GNDA.n346 76.3222
R2525 GNDA.n2270 GNDA.n2269 76.3222
R2526 GNDA.n2158 GNDA.n387 76.3222
R2527 GNDA.n2188 GNDA.n386 76.3222
R2528 GNDA.n2195 GNDA.n385 76.3222
R2529 GNDA.n2202 GNDA.n384 76.3222
R2530 GNDA.n2258 GNDA.n383 76.3222
R2531 GNDA.n1529 GNDA.n212 76.3222
R2532 GNDA.n1531 GNDA.n213 76.3222
R2533 GNDA.n1536 GNDA.n214 76.3222
R2534 GNDA.n1538 GNDA.n215 76.3222
R2535 GNDA.n1543 GNDA.n216 76.3222
R2536 GNDA.n2359 GNDA.n217 76.3222
R2537 GNDA.n1467 GNDA.n1466 76.3222
R2538 GNDA.n1472 GNDA.n1471 76.3222
R2539 GNDA.n1475 GNDA.n1474 76.3222
R2540 GNDA.n1480 GNDA.n1479 76.3222
R2541 GNDA.n1483 GNDA.n1482 76.3222
R2542 GNDA.n1488 GNDA.n1487 76.3222
R2543 GNDA.n1511 GNDA.n1510 76.3222
R2544 GNDA.n1527 GNDA.n1526 76.3222
R2545 GNDA.n1424 GNDA.n1344 76.3222
R2546 GNDA.n1435 GNDA.n1434 76.3222
R2547 GNDA.n1438 GNDA.n1437 76.3222
R2548 GNDA.n1447 GNDA.n1446 76.3222
R2549 GNDA.n1516 GNDA.n1515 76.3222
R2550 GNDA.n1526 GNDA.n1525 76.3222
R2551 GNDA.n1425 GNDA.n1424 76.3222
R2552 GNDA.n1436 GNDA.n1435 76.3222
R2553 GNDA.n1437 GNDA.n1420 76.3222
R2554 GNDA.n1448 GNDA.n1447 76.3222
R2555 GNDA.n1515 GNDA.n1514 76.3222
R2556 GNDA.n1861 GNDA.n651 76.3222
R2557 GNDA.n1882 GNDA.n492 76.3222
R2558 GNDA.n426 GNDA.n425 76.3222
R2559 GNDA.n424 GNDA.n404 76.3222
R2560 GNDA.n423 GNDA.n422 76.3222
R2561 GNDA.n421 GNDA.n398 76.3222
R2562 GNDA.n420 GNDA.n419 76.3222
R2563 GNDA.n417 GNDA.n391 76.3222
R2564 GNDA.n450 GNDA.n449 76.3222
R2565 GNDA.n444 GNDA.n443 76.3222
R2566 GNDA.n441 GNDA.n440 76.3222
R2567 GNDA.n435 GNDA.n434 76.3222
R2568 GNDA.n432 GNDA.n428 76.3222
R2569 GNDA.n2007 GNDA.n2006 76.3222
R2570 GNDA.n2137 GNDA.n2136 76.3222
R2571 GNDA.n407 GNDA.n402 76.3222
R2572 GNDA.n2144 GNDA.n2143 76.3222
R2573 GNDA.n401 GNDA.n396 76.3222
R2574 GNDA.n2151 GNDA.n2150 76.3222
R2575 GNDA.n2154 GNDA.n2153 76.3222
R2576 GNDA.n1988 GNDA.n1987 76.3222
R2577 GNDA.n447 GNDA.n439 76.3222
R2578 GNDA.n1995 GNDA.n1994 76.3222
R2579 GNDA.n438 GNDA.n431 76.3222
R2580 GNDA.n2002 GNDA.n2001 76.3222
R2581 GNDA.n430 GNDA.n412 76.3222
R2582 GNDA.n770 GNDA.n653 76.3222
R2583 GNDA.n768 GNDA.n658 76.3222
R2584 GNDA.n693 GNDA.n657 76.3222
R2585 GNDA.n701 GNDA.n656 76.3222
R2586 GNDA.n707 GNDA.n655 76.3222
R2587 GNDA.n654 GNDA.n393 76.3222
R2588 GNDA.n1652 GNDA.n1651 76.3222
R2589 GNDA.n1773 GNDA.n1772 76.3222
R2590 GNDA.n1770 GNDA.n1769 76.3222
R2591 GNDA.n1828 GNDA.n1585 76.3222
R2592 GNDA.n1826 GNDA.n1825 76.3222
R2593 GNDA.n1821 GNDA.n1594 76.3222
R2594 GNDA.n1819 GNDA.n1818 76.3222
R2595 GNDA.n1814 GNDA.n1605 76.3222
R2596 GNDA.n1812 GNDA.n1811 76.3222
R2597 GNDA.n1787 GNDA.n1607 76.3222
R2598 GNDA.n1791 GNDA.n1608 76.3222
R2599 GNDA.n1795 GNDA.n1609 76.3222
R2600 GNDA.n1799 GNDA.n1610 76.3222
R2601 GNDA.n1807 GNDA.n1611 76.3222
R2602 GNDA.n1809 GNDA.n1606 76.3222
R2603 GNDA.n1810 GNDA.n1809 76.3222
R2604 GNDA.n1807 GNDA.n1806 76.3222
R2605 GNDA.n1801 GNDA.n1610 76.3222
R2606 GNDA.n1798 GNDA.n1609 76.3222
R2607 GNDA.n1794 GNDA.n1608 76.3222
R2608 GNDA.n1790 GNDA.n1607 76.3222
R2609 GNDA.n1652 GNDA.n1621 76.3222
R2610 GNDA.n1772 GNDA.n1655 76.3222
R2611 GNDA.n1770 GNDA.n1657 76.3222
R2612 GNDA.n1578 GNDA.n1577 76.3222
R2613 GNDA.n1317 GNDA.n1316 76.3222
R2614 GNDA.n1328 GNDA.n1327 76.3222
R2615 GNDA.n1329 GNDA.n1312 76.3222
R2616 GNDA.n1340 GNDA.n1339 76.3222
R2617 GNDA.n1567 GNDA.n1566 76.3222
R2618 GNDA.n1603 GNDA.n1602 76.3222
R2619 GNDA.n1600 GNDA.n1599 76.3222
R2620 GNDA.n1597 GNDA.n1596 76.3222
R2621 GNDA.n1591 GNDA.n1590 76.3222
R2622 GNDA.n1588 GNDA.n1587 76.3222
R2623 GNDA.n1582 GNDA.n1581 76.3222
R2624 GNDA.n1813 GNDA.n1812 76.3222
R2625 GNDA.n1605 GNDA.n1595 76.3222
R2626 GNDA.n1820 GNDA.n1819 76.3222
R2627 GNDA.n1594 GNDA.n1586 76.3222
R2628 GNDA.n1827 GNDA.n1826 76.3222
R2629 GNDA.n1585 GNDA.n1232 76.3222
R2630 GNDA.n2279 GNDA.n222 76.3222
R2631 GNDA.n2278 GNDA.n2277 76.3222
R2632 GNDA.n2286 GNDA.n2285 76.3222
R2633 GNDA.n2276 GNDA.n2274 76.3222
R2634 GNDA.n2293 GNDA.n2292 76.3222
R2635 GNDA.n382 GNDA.n377 76.3222
R2636 GNDA.n1489 GNDA.n1488 76.3222
R2637 GNDA.n1482 GNDA.n1462 76.3222
R2638 GNDA.n1481 GNDA.n1480 76.3222
R2639 GNDA.n1474 GNDA.n1464 76.3222
R2640 GNDA.n1473 GNDA.n1472 76.3222
R2641 GNDA.n1468 GNDA.n1467 76.3222
R2642 GNDA.n2359 GNDA.n2358 76.3222
R2643 GNDA.n1544 GNDA.n216 76.3222
R2644 GNDA.n1542 GNDA.n215 76.3222
R2645 GNDA.n1537 GNDA.n214 76.3222
R2646 GNDA.n1535 GNDA.n213 76.3222
R2647 GNDA.n1530 GNDA.n212 76.3222
R2648 GNDA.n1546 GNDA.n221 76.3222
R2649 GNDA.n1545 GNDA.n1541 76.3222
R2650 GNDA.n1553 GNDA.n1552 76.3222
R2651 GNDA.n1540 GNDA.n1534 76.3222
R2652 GNDA.n1560 GNDA.n1559 76.3222
R2653 GNDA.n1533 GNDA.n1341 76.3222
R2654 GNDA.n361 GNDA.n211 76.3222
R2655 GNDA.n360 GNDA.n210 76.3222
R2656 GNDA.n358 GNDA.n209 76.3222
R2657 GNDA.n353 GNDA.n208 76.3222
R2658 GNDA.n351 GNDA.n207 76.3222
R2659 GNDA.n347 GNDA.n206 76.3222
R2660 GNDA.n2330 GNDA.n2329 76.3222
R2661 GNDA.n363 GNDA.n357 76.3222
R2662 GNDA.n2337 GNDA.n2336 76.3222
R2663 GNDA.n356 GNDA.n350 76.3222
R2664 GNDA.n2344 GNDA.n2343 76.3222
R2665 GNDA.n2347 GNDA.n2346 76.3222
R2666 GNDA.n340 GNDA.n226 76.3222
R2667 GNDA.n257 GNDA.n229 76.3222
R2668 GNDA.n263 GNDA.n262 76.3222
R2669 GNDA.n264 GNDA.n251 76.3222
R2670 GNDA.n278 GNDA.n277 76.3222
R2671 GNDA.n279 GNDA.n50 76.3222
R2672 GNDA.n2415 GNDA.n62 76.3222
R2673 GNDA.n2413 GNDA.n2412 76.3222
R2674 GNDA.n2408 GNDA.n2407 76.3222
R2675 GNDA.n2405 GNDA.n2404 76.3222
R2676 GNDA.n2400 GNDA.n2399 76.3222
R2677 GNDA.n2397 GNDA.n2396 76.3222
R2678 GNDA.n186 GNDA.n72 76.3222
R2679 GNDA.n103 GNDA.n75 76.3222
R2680 GNDA.n109 GNDA.n108 76.3222
R2681 GNDA.n110 GNDA.n97 76.3222
R2682 GNDA.n124 GNDA.n123 76.3222
R2683 GNDA.n125 GNDA.n41 76.3222
R2684 GNDA.n1511 GNDA.n1449 76.3222
R2685 GNDA.n2440 GNDA.n51 76.3222
R2686 GNDA.n2445 GNDA.n2444 76.3222
R2687 GNDA.t124 GNDA.t112 75.2142
R2688 GNDA.t115 GNDA.t17 75.2142
R2689 GNDA.n284 GNDA.n283 74.5978
R2690 GNDA.n285 GNDA.n284 74.5978
R2691 GNDA.n1572 GNDA.n1571 74.5978
R2692 GNDA.n1572 GNDA.n1258 74.5978
R2693 GNDA.n1714 GNDA.n1713 74.5978
R2694 GNDA.n1715 GNDA.n1714 74.5978
R2695 GNDA.n2068 GNDA.n2067 74.5978
R2696 GNDA.n2069 GNDA.n2068 74.5978
R2697 GNDA.n130 GNDA.n129 74.5978
R2698 GNDA.n131 GNDA.n130 74.5978
R2699 GNDA.n634 GNDA.n633 74.5978
R2700 GNDA.n634 GNDA.n581 74.5978
R2701 GNDA.n2262 GNDA.n2261 74.5978
R2702 GNDA.n2262 GNDA.n2179 74.5978
R2703 GNDA.n712 GNDA.n711 74.5978
R2704 GNDA.n713 GNDA.n712 74.5978
R2705 GNDA.n1520 GNDA.n1519 74.5978
R2706 GNDA.n1520 GNDA.n1366 74.5978
R2707 GNDA.n1650 GNDA.n1618 72.8884
R2708 GNDA.n1650 GNDA.n1649 72.8884
R2709 GNDA.n1649 GNDA.n1648 72.8884
R2710 GNDA.n1642 GNDA.n1627 72.8884
R2711 GNDA.n1641 GNDA.n1640 72.8884
R2712 GNDA.n1640 GNDA.n1628 72.8884
R2713 GNDA.n1634 GNDA.n1628 72.8884
R2714 GNDA.n1634 GNDA.n1633 72.8884
R2715 GNDA.n1633 GNDA.n1614 72.8884
R2716 GNDA.n1862 GNDA.n1860 72.8884
R2717 GNDA.n1870 GNDA.n649 72.8884
R2718 GNDA.n1926 GNDA.n478 72.8884
R2719 GNDA.n1926 GNDA.n1925 72.8884
R2720 GNDA.n501 GNDA.n480 72.8884
R2721 GNDA.n501 GNDA.n496 72.8884
R2722 GNDA.n1883 GNDA.n1881 72.8884
R2723 GNDA.n1917 GNDA.n489 72.8884
R2724 GNDA.n1911 GNDA.n489 72.8884
R2725 GNDA.n1911 GNDA.n1910 72.8884
R2726 GNDA.n1909 GNDA.n1890 72.8884
R2727 GNDA.n1903 GNDA.n1890 72.8884
R2728 GNDA.n1903 GNDA.n1902 72.8884
R2729 GNDA.n1902 GNDA.n1901 72.8884
R2730 GNDA.t288 GNDA.t152 72.0803
R2731 GNDA.t229 GNDA.t153 72.0803
R2732 GNDA.t300 GNDA.t141 70.9682
R2733 GNDA.t182 GNDA.t49 70.9682
R2734 GNDA.t91 GNDA.t127 70.9682
R2735 GNDA.t235 GNDA.t15 70.9682
R2736 GNDA.n1933 GNDA.n1932 70.4588
R2737 GNDA.n647 GNDA.n646 70.4588
R2738 GNDA.n1863 GNDA.t225 69.6489
R2739 GNDA.n1884 GNDA.n647 69.6489
R2740 GNDA.n317 GNDA.n316 69.3109
R2741 GNDA.n316 GNDA.n315 69.3109
R2742 GNDA.n1276 GNDA.n1248 69.3109
R2743 GNDA.n1279 GNDA.n1248 69.3109
R2744 GNDA.n1747 GNDA.n1746 69.3109
R2745 GNDA.n1746 GNDA.n1745 69.3109
R2746 GNDA.n2101 GNDA.n2100 69.3109
R2747 GNDA.n2100 GNDA.n2099 69.3109
R2748 GNDA.n163 GNDA.n162 69.3109
R2749 GNDA.n162 GNDA.n161 69.3109
R2750 GNDA.n546 GNDA.n521 69.3109
R2751 GNDA.n549 GNDA.n521 69.3109
R2752 GNDA.n2220 GNDA.n2169 69.3109
R2753 GNDA.n2223 GNDA.n2169 69.3109
R2754 GNDA.n745 GNDA.n744 69.3109
R2755 GNDA.n744 GNDA.n743 69.3109
R2756 GNDA.n1384 GNDA.n1356 69.3109
R2757 GNDA.n1387 GNDA.n1356 69.3109
R2758 GNDA.t146 GNDA.t294 68.9464
R2759 GNDA.t0 GNDA.t146 68.9464
R2760 GNDA.t144 GNDA.t0 68.9464
R2761 GNDA.t68 GNDA.t40 68.9464
R2762 GNDA.t166 GNDA.t68 68.9464
R2763 GNDA.t274 GNDA.t166 68.9464
R2764 GNDA.n296 GNDA.t276 65.8183
R2765 GNDA.n293 GNDA.t276 65.8183
R2766 GNDA.n287 GNDA.t276 65.8183
R2767 GNDA.n302 GNDA.t276 65.8183
R2768 GNDA.n241 GNDA.t276 65.8183
R2769 GNDA.n309 GNDA.t276 65.8183
R2770 GNDA.n238 GNDA.t276 65.8183
R2771 GNDA.n318 GNDA.t276 65.8183
R2772 GNDA.n324 GNDA.t276 65.8183
R2773 GNDA.n326 GNDA.t276 65.8183
R2774 GNDA.n332 GNDA.t276 65.8183
R2775 GNDA.t226 GNDA.n1247 65.8183
R2776 GNDA.t226 GNDA.n1245 65.8183
R2777 GNDA.t226 GNDA.n1243 65.8183
R2778 GNDA.t226 GNDA.n1250 65.8183
R2779 GNDA.t226 GNDA.n1251 65.8183
R2780 GNDA.t226 GNDA.n1252 65.8183
R2781 GNDA.t226 GNDA.n1253 65.8183
R2782 GNDA.t226 GNDA.n1246 65.8183
R2783 GNDA.t226 GNDA.n1244 65.8183
R2784 GNDA.t226 GNDA.n1242 65.8183
R2785 GNDA.t226 GNDA.n1241 65.8183
R2786 GNDA.n1726 GNDA.t224 65.8183
R2787 GNDA.n1723 GNDA.t224 65.8183
R2788 GNDA.n1717 GNDA.t224 65.8183
R2789 GNDA.n1732 GNDA.t224 65.8183
R2790 GNDA.n1672 GNDA.t224 65.8183
R2791 GNDA.n1739 GNDA.t224 65.8183
R2792 GNDA.n1669 GNDA.t224 65.8183
R2793 GNDA.n1665 GNDA.t224 65.8183
R2794 GNDA.n1752 GNDA.t224 65.8183
R2795 GNDA.n1758 GNDA.t224 65.8183
R2796 GNDA.n1662 GNDA.t224 65.8183
R2797 GNDA.n2080 GNDA.t315 65.8183
R2798 GNDA.n2077 GNDA.t315 65.8183
R2799 GNDA.n2071 GNDA.t315 65.8183
R2800 GNDA.n2086 GNDA.t315 65.8183
R2801 GNDA.n2029 GNDA.t315 65.8183
R2802 GNDA.n2093 GNDA.t315 65.8183
R2803 GNDA.n2026 GNDA.t315 65.8183
R2804 GNDA.n2022 GNDA.t315 65.8183
R2805 GNDA.n2106 GNDA.t315 65.8183
R2806 GNDA.n2112 GNDA.t315 65.8183
R2807 GNDA.n2019 GNDA.t315 65.8183
R2808 GNDA.n142 GNDA.t237 65.8183
R2809 GNDA.n139 GNDA.t237 65.8183
R2810 GNDA.n133 GNDA.t237 65.8183
R2811 GNDA.n148 GNDA.t237 65.8183
R2812 GNDA.n87 GNDA.t237 65.8183
R2813 GNDA.n155 GNDA.t237 65.8183
R2814 GNDA.n84 GNDA.t237 65.8183
R2815 GNDA.n164 GNDA.t237 65.8183
R2816 GNDA.n170 GNDA.t237 65.8183
R2817 GNDA.n172 GNDA.t237 65.8183
R2818 GNDA.n178 GNDA.t237 65.8183
R2819 GNDA.n181 GNDA.t237 65.8183
R2820 GNDA.n100 GNDA.t237 65.8183
R2821 GNDA.n115 GNDA.t237 65.8183
R2822 GNDA.n117 GNDA.t237 65.8183
R2823 GNDA.t314 GNDA.n520 65.8183
R2824 GNDA.t314 GNDA.n518 65.8183
R2825 GNDA.t314 GNDA.n516 65.8183
R2826 GNDA.t314 GNDA.n523 65.8183
R2827 GNDA.t314 GNDA.n524 65.8183
R2828 GNDA.t314 GNDA.n525 65.8183
R2829 GNDA.t314 GNDA.n526 65.8183
R2830 GNDA.t314 GNDA.n519 65.8183
R2831 GNDA.t314 GNDA.n517 65.8183
R2832 GNDA.t314 GNDA.n515 65.8183
R2833 GNDA.t314 GNDA.n514 65.8183
R2834 GNDA.n635 GNDA.t314 65.8183
R2835 GNDA.t314 GNDA.n528 65.8183
R2836 GNDA.t314 GNDA.n529 65.8183
R2837 GNDA.t314 GNDA.n530 65.8183
R2838 GNDA.n2119 GNDA.t315 65.8183
R2839 GNDA.n2041 GNDA.t315 65.8183
R2840 GNDA.n2052 GNDA.t315 65.8183
R2841 GNDA.n2039 GNDA.t315 65.8183
R2842 GNDA.t254 GNDA.n2168 65.8183
R2843 GNDA.t254 GNDA.n2166 65.8183
R2844 GNDA.t254 GNDA.n2164 65.8183
R2845 GNDA.t254 GNDA.n2171 65.8183
R2846 GNDA.t254 GNDA.n2172 65.8183
R2847 GNDA.t254 GNDA.n2173 65.8183
R2848 GNDA.t254 GNDA.n2174 65.8183
R2849 GNDA.t254 GNDA.n2167 65.8183
R2850 GNDA.t254 GNDA.n2165 65.8183
R2851 GNDA.t254 GNDA.n2163 65.8183
R2852 GNDA.t254 GNDA.n2162 65.8183
R2853 GNDA.n724 GNDA.t253 65.8183
R2854 GNDA.n721 GNDA.t253 65.8183
R2855 GNDA.n715 GNDA.t253 65.8183
R2856 GNDA.n730 GNDA.t253 65.8183
R2857 GNDA.n674 GNDA.t253 65.8183
R2858 GNDA.n737 GNDA.t253 65.8183
R2859 GNDA.n671 GNDA.t253 65.8183
R2860 GNDA.n667 GNDA.t253 65.8183
R2861 GNDA.n750 GNDA.t253 65.8183
R2862 GNDA.n756 GNDA.t253 65.8183
R2863 GNDA.n662 GNDA.t253 65.8183
R2864 GNDA.n763 GNDA.t253 65.8183
R2865 GNDA.n686 GNDA.t253 65.8183
R2866 GNDA.n697 GNDA.t253 65.8183
R2867 GNDA.n684 GNDA.t253 65.8183
R2868 GNDA.n2263 GNDA.t254 65.8183
R2869 GNDA.t254 GNDA.n2176 65.8183
R2870 GNDA.t254 GNDA.n2177 65.8183
R2871 GNDA.t254 GNDA.n2178 65.8183
R2872 GNDA.t280 GNDA.n1355 65.8183
R2873 GNDA.t280 GNDA.n1353 65.8183
R2874 GNDA.t280 GNDA.n1351 65.8183
R2875 GNDA.t280 GNDA.n1358 65.8183
R2876 GNDA.t280 GNDA.n1359 65.8183
R2877 GNDA.t280 GNDA.n1360 65.8183
R2878 GNDA.t280 GNDA.n1361 65.8183
R2879 GNDA.t280 GNDA.n1354 65.8183
R2880 GNDA.t280 GNDA.n1352 65.8183
R2881 GNDA.t280 GNDA.n1350 65.8183
R2882 GNDA.t280 GNDA.n1349 65.8183
R2883 GNDA.n1521 GNDA.t280 65.8183
R2884 GNDA.t280 GNDA.n1363 65.8183
R2885 GNDA.t280 GNDA.n1364 65.8183
R2886 GNDA.t280 GNDA.n1365 65.8183
R2887 GNDA.n1765 GNDA.t224 65.8183
R2888 GNDA.n1686 GNDA.t224 65.8183
R2889 GNDA.n1699 GNDA.t224 65.8183
R2890 GNDA.n1701 GNDA.t224 65.8183
R2891 GNDA.n1573 GNDA.t226 65.8183
R2892 GNDA.t226 GNDA.n1255 65.8183
R2893 GNDA.t226 GNDA.n1256 65.8183
R2894 GNDA.t226 GNDA.n1257 65.8183
R2895 GNDA.n335 GNDA.t276 65.8183
R2896 GNDA.n254 GNDA.t276 65.8183
R2897 GNDA.n269 GNDA.t276 65.8183
R2898 GNDA.n271 GNDA.t276 65.8183
R2899 GNDA.n1187 GNDA.t144 65.8125
R2900 GNDA.t40 GNDA.n824 65.8125
R2901 GNDA.n1107 GNDA.n1106 64.0005
R2902 GNDA.n1107 GNDA.n1102 64.0005
R2903 GNDA.n1203 GNDA.t214 62.6786
R2904 GNDA.t36 GNDA.n819 62.6786
R2905 GNDA.n1924 GNDA.n480 62.3602
R2906 GNDA.t227 GNDA.n0 32.9056
R2907 GNDA.n1092 GNDA.n1091 60.8005
R2908 GNDA.t345 GNDA.t79 59.5447
R2909 GNDA.t189 GNDA.t354 59.5447
R2910 GNDA.n316 GNDA.t276 57.8461
R2911 GNDA.t226 GNDA.n1248 57.8461
R2912 GNDA.n1746 GNDA.t224 57.8461
R2913 GNDA.n2100 GNDA.t315 57.8461
R2914 GNDA.n162 GNDA.t237 57.8461
R2915 GNDA.t314 GNDA.n521 57.8461
R2916 GNDA.t254 GNDA.n2169 57.8461
R2917 GNDA.n744 GNDA.t253 57.8461
R2918 GNDA.t280 GNDA.n1356 57.8461
R2919 GNDA.t19 GNDA.n987 57.241
R2920 GNDA.t106 GNDA.t48 56.0277
R2921 GNDA.t97 GNDA.t74 56.0277
R2922 GNDA.t72 GNDA.t128 56.0277
R2923 GNDA.t198 GNDA.t208 56.0277
R2924 GNDA.n130 GNDA.t237 55.2026
R2925 GNDA.t314 GNDA.n634 55.2026
R2926 GNDA.n2068 GNDA.t315 55.2026
R2927 GNDA.n712 GNDA.t253 55.2026
R2928 GNDA.t254 GNDA.n2262 55.2026
R2929 GNDA.t280 GNDA.n1520 55.2026
R2930 GNDA.n1714 GNDA.t224 55.2026
R2931 GNDA.t226 GNDA.n1572 55.2026
R2932 GNDA.n284 GNDA.t276 55.2026
R2933 GNDA.n1093 GNDA.n1092 54.4005
R2934 GNDA.n1858 GNDA.n649 54.2615
R2935 GNDA.n335 GNDA.n334 53.3664
R2936 GNDA.n254 GNDA.n231 53.3664
R2937 GNDA.n269 GNDA.n268 53.3664
R2938 GNDA.n272 GNDA.n271 53.3664
R2939 GNDA.n333 GNDA.n332 53.3664
R2940 GNDA.n326 GNDA.n232 53.3664
R2941 GNDA.n325 GNDA.n324 53.3664
R2942 GNDA.n318 GNDA.n234 53.3664
R2943 GNDA.n311 GNDA.n238 53.3664
R2944 GNDA.n309 GNDA.n308 53.3664
R2945 GNDA.n304 GNDA.n241 53.3664
R2946 GNDA.n302 GNDA.n301 53.3664
R2947 GNDA.n288 GNDA.n287 53.3664
R2948 GNDA.n293 GNDA.n292 53.3664
R2949 GNDA.n296 GNDA.n295 53.3664
R2950 GNDA.n297 GNDA.n296 53.3664
R2951 GNDA.n294 GNDA.n293 53.3664
R2952 GNDA.n287 GNDA.n245 53.3664
R2953 GNDA.n303 GNDA.n302 53.3664
R2954 GNDA.n241 GNDA.n239 53.3664
R2955 GNDA.n310 GNDA.n309 53.3664
R2956 GNDA.n238 GNDA.n236 53.3664
R2957 GNDA.n319 GNDA.n318 53.3664
R2958 GNDA.n324 GNDA.n323 53.3664
R2959 GNDA.n327 GNDA.n326 53.3664
R2960 GNDA.n332 GNDA.n331 53.3664
R2961 GNDA.n1574 GNDA.n1573 53.3664
R2962 GNDA.n1320 GNDA.n1255 53.3664
R2963 GNDA.n1322 GNDA.n1256 53.3664
R2964 GNDA.n1334 GNDA.n1257 53.3664
R2965 GNDA.n1241 GNDA.n1239 53.3664
R2966 GNDA.n1264 GNDA.n1242 53.3664
R2967 GNDA.n1268 GNDA.n1244 53.3664
R2968 GNDA.n1272 GNDA.n1246 53.3664
R2969 GNDA.n1283 GNDA.n1253 53.3664
R2970 GNDA.n1287 GNDA.n1252 53.3664
R2971 GNDA.n1291 GNDA.n1251 53.3664
R2972 GNDA.n1294 GNDA.n1250 53.3664
R2973 GNDA.n1307 GNDA.n1243 53.3664
R2974 GNDA.n1304 GNDA.n1245 53.3664
R2975 GNDA.n1300 GNDA.n1247 53.3664
R2976 GNDA.n1297 GNDA.n1247 53.3664
R2977 GNDA.n1301 GNDA.n1245 53.3664
R2978 GNDA.n1305 GNDA.n1243 53.3664
R2979 GNDA.n1292 GNDA.n1250 53.3664
R2980 GNDA.n1288 GNDA.n1251 53.3664
R2981 GNDA.n1284 GNDA.n1252 53.3664
R2982 GNDA.n1280 GNDA.n1253 53.3664
R2983 GNDA.n1275 GNDA.n1246 53.3664
R2984 GNDA.n1271 GNDA.n1244 53.3664
R2985 GNDA.n1267 GNDA.n1242 53.3664
R2986 GNDA.n1263 GNDA.n1241 53.3664
R2987 GNDA.n1765 GNDA.n1764 53.3664
R2988 GNDA.n1686 GNDA.n1661 53.3664
R2989 GNDA.n1699 GNDA.n1698 53.3664
R2990 GNDA.n1702 GNDA.n1701 53.3664
R2991 GNDA.n1763 GNDA.n1662 53.3664
R2992 GNDA.n1759 GNDA.n1758 53.3664
R2993 GNDA.n1752 GNDA.n1664 53.3664
R2994 GNDA.n1751 GNDA.n1665 53.3664
R2995 GNDA.n1741 GNDA.n1669 53.3664
R2996 GNDA.n1739 GNDA.n1738 53.3664
R2997 GNDA.n1734 GNDA.n1672 53.3664
R2998 GNDA.n1732 GNDA.n1731 53.3664
R2999 GNDA.n1718 GNDA.n1717 53.3664
R3000 GNDA.n1723 GNDA.n1722 53.3664
R3001 GNDA.n1726 GNDA.n1725 53.3664
R3002 GNDA.n1727 GNDA.n1726 53.3664
R3003 GNDA.n1724 GNDA.n1723 53.3664
R3004 GNDA.n1717 GNDA.n1676 53.3664
R3005 GNDA.n1733 GNDA.n1732 53.3664
R3006 GNDA.n1672 GNDA.n1670 53.3664
R3007 GNDA.n1740 GNDA.n1739 53.3664
R3008 GNDA.n1669 GNDA.n1667 53.3664
R3009 GNDA.n1748 GNDA.n1665 53.3664
R3010 GNDA.n1753 GNDA.n1752 53.3664
R3011 GNDA.n1758 GNDA.n1757 53.3664
R3012 GNDA.n1760 GNDA.n1662 53.3664
R3013 GNDA.n2119 GNDA.n2118 53.3664
R3014 GNDA.n2041 GNDA.n2018 53.3664
R3015 GNDA.n2052 GNDA.n2051 53.3664
R3016 GNDA.n2040 GNDA.n2039 53.3664
R3017 GNDA.n2117 GNDA.n2019 53.3664
R3018 GNDA.n2113 GNDA.n2112 53.3664
R3019 GNDA.n2106 GNDA.n2021 53.3664
R3020 GNDA.n2105 GNDA.n2022 53.3664
R3021 GNDA.n2095 GNDA.n2026 53.3664
R3022 GNDA.n2093 GNDA.n2092 53.3664
R3023 GNDA.n2088 GNDA.n2029 53.3664
R3024 GNDA.n2086 GNDA.n2085 53.3664
R3025 GNDA.n2072 GNDA.n2071 53.3664
R3026 GNDA.n2077 GNDA.n2076 53.3664
R3027 GNDA.n2080 GNDA.n2079 53.3664
R3028 GNDA.n2081 GNDA.n2080 53.3664
R3029 GNDA.n2078 GNDA.n2077 53.3664
R3030 GNDA.n2071 GNDA.n2033 53.3664
R3031 GNDA.n2087 GNDA.n2086 53.3664
R3032 GNDA.n2029 GNDA.n2027 53.3664
R3033 GNDA.n2094 GNDA.n2093 53.3664
R3034 GNDA.n2026 GNDA.n2024 53.3664
R3035 GNDA.n2102 GNDA.n2022 53.3664
R3036 GNDA.n2107 GNDA.n2106 53.3664
R3037 GNDA.n2112 GNDA.n2111 53.3664
R3038 GNDA.n2114 GNDA.n2019 53.3664
R3039 GNDA.n181 GNDA.n180 53.3664
R3040 GNDA.n100 GNDA.n77 53.3664
R3041 GNDA.n115 GNDA.n114 53.3664
R3042 GNDA.n118 GNDA.n117 53.3664
R3043 GNDA.n179 GNDA.n178 53.3664
R3044 GNDA.n172 GNDA.n78 53.3664
R3045 GNDA.n171 GNDA.n170 53.3664
R3046 GNDA.n164 GNDA.n80 53.3664
R3047 GNDA.n157 GNDA.n84 53.3664
R3048 GNDA.n155 GNDA.n154 53.3664
R3049 GNDA.n150 GNDA.n87 53.3664
R3050 GNDA.n148 GNDA.n147 53.3664
R3051 GNDA.n134 GNDA.n133 53.3664
R3052 GNDA.n139 GNDA.n138 53.3664
R3053 GNDA.n142 GNDA.n141 53.3664
R3054 GNDA.n143 GNDA.n142 53.3664
R3055 GNDA.n140 GNDA.n139 53.3664
R3056 GNDA.n133 GNDA.n91 53.3664
R3057 GNDA.n149 GNDA.n148 53.3664
R3058 GNDA.n87 GNDA.n85 53.3664
R3059 GNDA.n156 GNDA.n155 53.3664
R3060 GNDA.n84 GNDA.n82 53.3664
R3061 GNDA.n165 GNDA.n164 53.3664
R3062 GNDA.n170 GNDA.n169 53.3664
R3063 GNDA.n173 GNDA.n172 53.3664
R3064 GNDA.n178 GNDA.n177 53.3664
R3065 GNDA.n182 GNDA.n181 53.3664
R3066 GNDA.n101 GNDA.n100 53.3664
R3067 GNDA.n116 GNDA.n115 53.3664
R3068 GNDA.n117 GNDA.n94 53.3664
R3069 GNDA.n636 GNDA.n635 53.3664
R3070 GNDA.n592 GNDA.n528 53.3664
R3071 GNDA.n611 GNDA.n529 53.3664
R3072 GNDA.n617 GNDA.n530 53.3664
R3073 GNDA.n514 GNDA.n512 53.3664
R3074 GNDA.n534 GNDA.n515 53.3664
R3075 GNDA.n538 GNDA.n517 53.3664
R3076 GNDA.n542 GNDA.n519 53.3664
R3077 GNDA.n553 GNDA.n526 53.3664
R3078 GNDA.n557 GNDA.n525 53.3664
R3079 GNDA.n561 GNDA.n524 53.3664
R3080 GNDA.n564 GNDA.n523 53.3664
R3081 GNDA.n577 GNDA.n516 53.3664
R3082 GNDA.n574 GNDA.n518 53.3664
R3083 GNDA.n570 GNDA.n520 53.3664
R3084 GNDA.n567 GNDA.n520 53.3664
R3085 GNDA.n571 GNDA.n518 53.3664
R3086 GNDA.n575 GNDA.n516 53.3664
R3087 GNDA.n562 GNDA.n523 53.3664
R3088 GNDA.n558 GNDA.n524 53.3664
R3089 GNDA.n554 GNDA.n525 53.3664
R3090 GNDA.n550 GNDA.n526 53.3664
R3091 GNDA.n545 GNDA.n519 53.3664
R3092 GNDA.n541 GNDA.n517 53.3664
R3093 GNDA.n537 GNDA.n515 53.3664
R3094 GNDA.n533 GNDA.n514 53.3664
R3095 GNDA.n635 GNDA.n513 53.3664
R3096 GNDA.n610 GNDA.n528 53.3664
R3097 GNDA.n616 GNDA.n529 53.3664
R3098 GNDA.n582 GNDA.n530 53.3664
R3099 GNDA.n2120 GNDA.n2119 53.3664
R3100 GNDA.n2042 GNDA.n2041 53.3664
R3101 GNDA.n2053 GNDA.n2052 53.3664
R3102 GNDA.n2039 GNDA.n2036 53.3664
R3103 GNDA.n2264 GNDA.n2263 53.3664
R3104 GNDA.n2183 GNDA.n2176 53.3664
R3105 GNDA.n2190 GNDA.n2177 53.3664
R3106 GNDA.n2197 GNDA.n2178 53.3664
R3107 GNDA.n2162 GNDA.n2160 53.3664
R3108 GNDA.n2208 GNDA.n2163 53.3664
R3109 GNDA.n2212 GNDA.n2165 53.3664
R3110 GNDA.n2216 GNDA.n2167 53.3664
R3111 GNDA.n2227 GNDA.n2174 53.3664
R3112 GNDA.n2231 GNDA.n2173 53.3664
R3113 GNDA.n2235 GNDA.n2172 53.3664
R3114 GNDA.n2238 GNDA.n2171 53.3664
R3115 GNDA.n2251 GNDA.n2164 53.3664
R3116 GNDA.n2248 GNDA.n2166 53.3664
R3117 GNDA.n2244 GNDA.n2168 53.3664
R3118 GNDA.n2241 GNDA.n2168 53.3664
R3119 GNDA.n2245 GNDA.n2166 53.3664
R3120 GNDA.n2249 GNDA.n2164 53.3664
R3121 GNDA.n2236 GNDA.n2171 53.3664
R3122 GNDA.n2232 GNDA.n2172 53.3664
R3123 GNDA.n2228 GNDA.n2173 53.3664
R3124 GNDA.n2224 GNDA.n2174 53.3664
R3125 GNDA.n2219 GNDA.n2167 53.3664
R3126 GNDA.n2215 GNDA.n2165 53.3664
R3127 GNDA.n2211 GNDA.n2163 53.3664
R3128 GNDA.n2207 GNDA.n2162 53.3664
R3129 GNDA.n763 GNDA.n762 53.3664
R3130 GNDA.n686 GNDA.n661 53.3664
R3131 GNDA.n697 GNDA.n696 53.3664
R3132 GNDA.n685 GNDA.n684 53.3664
R3133 GNDA.n761 GNDA.n662 53.3664
R3134 GNDA.n757 GNDA.n756 53.3664
R3135 GNDA.n750 GNDA.n666 53.3664
R3136 GNDA.n749 GNDA.n667 53.3664
R3137 GNDA.n739 GNDA.n671 53.3664
R3138 GNDA.n737 GNDA.n736 53.3664
R3139 GNDA.n732 GNDA.n674 53.3664
R3140 GNDA.n730 GNDA.n729 53.3664
R3141 GNDA.n716 GNDA.n715 53.3664
R3142 GNDA.n721 GNDA.n720 53.3664
R3143 GNDA.n724 GNDA.n723 53.3664
R3144 GNDA.n725 GNDA.n724 53.3664
R3145 GNDA.n722 GNDA.n721 53.3664
R3146 GNDA.n715 GNDA.n678 53.3664
R3147 GNDA.n731 GNDA.n730 53.3664
R3148 GNDA.n674 GNDA.n672 53.3664
R3149 GNDA.n738 GNDA.n737 53.3664
R3150 GNDA.n671 GNDA.n669 53.3664
R3151 GNDA.n746 GNDA.n667 53.3664
R3152 GNDA.n751 GNDA.n750 53.3664
R3153 GNDA.n756 GNDA.n755 53.3664
R3154 GNDA.n758 GNDA.n662 53.3664
R3155 GNDA.n764 GNDA.n763 53.3664
R3156 GNDA.n687 GNDA.n686 53.3664
R3157 GNDA.n698 GNDA.n697 53.3664
R3158 GNDA.n684 GNDA.n681 53.3664
R3159 GNDA.n2263 GNDA.n2161 53.3664
R3160 GNDA.n2191 GNDA.n2176 53.3664
R3161 GNDA.n2198 GNDA.n2177 53.3664
R3162 GNDA.n2180 GNDA.n2178 53.3664
R3163 GNDA.n1522 GNDA.n1521 53.3664
R3164 GNDA.n1428 GNDA.n1363 53.3664
R3165 GNDA.n1430 GNDA.n1364 53.3664
R3166 GNDA.n1442 GNDA.n1365 53.3664
R3167 GNDA.n1349 GNDA.n1347 53.3664
R3168 GNDA.n1372 GNDA.n1350 53.3664
R3169 GNDA.n1376 GNDA.n1352 53.3664
R3170 GNDA.n1380 GNDA.n1354 53.3664
R3171 GNDA.n1391 GNDA.n1361 53.3664
R3172 GNDA.n1395 GNDA.n1360 53.3664
R3173 GNDA.n1399 GNDA.n1359 53.3664
R3174 GNDA.n1402 GNDA.n1358 53.3664
R3175 GNDA.n1415 GNDA.n1351 53.3664
R3176 GNDA.n1412 GNDA.n1353 53.3664
R3177 GNDA.n1408 GNDA.n1355 53.3664
R3178 GNDA.n1405 GNDA.n1355 53.3664
R3179 GNDA.n1409 GNDA.n1353 53.3664
R3180 GNDA.n1413 GNDA.n1351 53.3664
R3181 GNDA.n1400 GNDA.n1358 53.3664
R3182 GNDA.n1396 GNDA.n1359 53.3664
R3183 GNDA.n1392 GNDA.n1360 53.3664
R3184 GNDA.n1388 GNDA.n1361 53.3664
R3185 GNDA.n1383 GNDA.n1354 53.3664
R3186 GNDA.n1379 GNDA.n1352 53.3664
R3187 GNDA.n1375 GNDA.n1350 53.3664
R3188 GNDA.n1371 GNDA.n1349 53.3664
R3189 GNDA.n1521 GNDA.n1348 53.3664
R3190 GNDA.n1431 GNDA.n1363 53.3664
R3191 GNDA.n1441 GNDA.n1364 53.3664
R3192 GNDA.n1367 GNDA.n1365 53.3664
R3193 GNDA.n1766 GNDA.n1765 53.3664
R3194 GNDA.n1687 GNDA.n1686 53.3664
R3195 GNDA.n1700 GNDA.n1699 53.3664
R3196 GNDA.n1701 GNDA.n1679 53.3664
R3197 GNDA.n1573 GNDA.n1240 53.3664
R3198 GNDA.n1323 GNDA.n1255 53.3664
R3199 GNDA.n1333 GNDA.n1256 53.3664
R3200 GNDA.n1259 GNDA.n1257 53.3664
R3201 GNDA.n336 GNDA.n335 53.3664
R3202 GNDA.n255 GNDA.n254 53.3664
R3203 GNDA.n270 GNDA.n269 53.3664
R3204 GNDA.n271 GNDA.n248 53.3664
R3205 GNDA.t322 GNDA.t137 52.4707
R3206 GNDA.t158 GNDA.t174 52.4707
R3207 GNDA.t320 GNDA.t163 52.4707
R3208 GNDA.n1106 GNDA.n1105 51.2005
R3209 GNDA.n1102 GNDA.n1101 51.2005
R3210 GNDA.n1835 GNDA.n1834 50.9355
R3211 GNDA.n2513 GNDA.n5 50.5752
R3212 GNDA.n1204 GNDA.n1203 50.1429
R3213 GNDA.t45 GNDA.t337 50.1429
R3214 GNDA.t154 GNDA.t129 50.1429
R3215 GNDA.n1227 GNDA.n819 50.1429
R3216 GNDA.t270 GNDA.n932 48.7228
R3217 GNDA.n1026 GNDA.t176 48.5574
R3218 GNDA.n982 GNDA.t61 48.5574
R3219 GNDA.n1055 GNDA.t98 48.5574
R3220 GNDA.n1159 GNDA.t207 48.5574
R3221 GNDA.n1229 GNDA.t227 48.2626
R3222 GNDA.n917 GNDA.t131 48.0005
R3223 GNDA.n917 GNDA.t213 48.0005
R3224 GNDA.n914 GNDA.t181 48.0005
R3225 GNDA.n914 GNDA.t111 48.0005
R3226 GNDA.n913 GNDA.t138 48.0005
R3227 GNDA.n913 GNDA.t175 48.0005
R3228 GNDA.n911 GNDA.t52 48.0005
R3229 GNDA.n911 GNDA.t65 48.0005
R3230 GNDA.n910 GNDA.t7 48.0005
R3231 GNDA.n910 GNDA.t140 48.0005
R3232 GNDA.n1499 GNDA.t227 47.9486
R3233 GNDA.n2428 GNDA.t227 47.9486
R3234 GNDA.n2458 GNDA.t227 47.9486
R3235 GNDA.n194 GNDA.t227 47.6748
R3236 GNDA.t214 GNDA.t262 47.009
R3237 GNDA.t81 GNDA.t195 47.009
R3238 GNDA.t10 GNDA.t70 47.009
R3239 GNDA.t282 GNDA.t36 47.009
R3240 GNDA.n1785 GNDA.n1784 46.1628
R3241 GNDA.n1871 GNDA.n472 46.1628
R3242 GNDA.n1896 GNDA.n1895 46.1628
R3243 GNDA.t334 GNDA.t149 44.9749
R3244 GNDA.t191 GNDA.t169 44.9749
R3245 GNDA.t4 GNDA.t331 44.9749
R3246 GNDA.t164 GNDA.t355 44.9749
R3247 GNDA.t12 GNDA.t2 44.9749
R3248 GNDA.t155 GNDA.t218 44.9749
R3249 GNDA.t196 GNDA.t38 44.9749
R3250 GNDA.t159 GNDA.t192 44.9749
R3251 GNDA.t24 GNDA.t16 44.9749
R3252 GNDA.t120 GNDA.t312 44.9749
R3253 GNDA.n1042 GNDA.n1041 44.8222
R3254 GNDA.n1176 GNDA.n1175 44.8222
R3255 GNDA.n1002 GNDA.n1000 44.8005
R3256 GNDA.n1022 GNDA.n1021 44.8005
R3257 GNDA.n1501 GNDA.t227 43.8679
R3258 GNDA.t227 GNDA.n55 43.8679
R3259 GNDA.n2451 GNDA.t227 43.8679
R3260 GNDA.n1692 GNDA.n1656 43.0993
R3261 GNDA.t171 GNDA.n954 41.2271
R3262 GNDA.t47 GNDA.n1110 41.2271
R3263 GNDA.n1135 GNDA.t172 41.2271
R3264 GNDA.n933 GNDA.t327 41.2271
R3265 GNDA.n933 GNDA.t309 41.2271
R3266 GNDA.t90 GNDA.n1026 41.0871
R3267 GNDA.t350 GNDA.n982 41.0871
R3268 GNDA.t341 GNDA.t125 41.0871
R3269 GNDA.t341 GNDA.t339 41.0871
R3270 GNDA.t80 GNDA.t178 41.0871
R3271 GNDA.t178 GNDA.t209 41.0871
R3272 GNDA.n1165 GNDA.t54 40.7412
R3273 GNDA.t112 GNDA.n1168 40.7412
R3274 GNDA.t76 GNDA.t99 40.7412
R3275 GNDA.t187 GNDA.t343 40.7412
R3276 GNDA.t53 GNDA.t8 40.7412
R3277 GNDA.t185 GNDA.t336 40.7412
R3278 GNDA.t225 GNDA.n1641 38.0642
R3279 GNDA.n478 GNDA.t225 38.0642
R3280 GNDA.t225 GNDA.n1909 38.0642
R3281 GNDA.n1196 GNDA.t78 37.6073
R3282 GNDA.n1211 GNDA.t152 37.6073
R3283 GNDA.n1211 GNDA.t77 37.6073
R3284 GNDA.n830 GNDA.t194 37.6073
R3285 GNDA.t153 GNDA.n830 37.6073
R3286 GNDA.n831 GNDA.t32 37.6073
R3287 GNDA.t242 GNDA.t317 37.4792
R3288 GNDA.t232 GNDA.t328 37.4792
R3289 GNDA.t251 GNDA.t329 37.4792
R3290 GNDA.t201 GNDA.t139 37.4792
R3291 GNDA.t323 GNDA.t64 37.4792
R3292 GNDA.t168 GNDA.t130 37.4792
R3293 GNDA.t94 GNDA.t212 37.4792
R3294 GNDA.t333 GNDA.t180 37.4792
R3295 GNDA.t222 GNDA.t110 37.4792
R3296 GNDA.t88 GNDA.t35 37.4792
R3297 GNDA.t172 GNDA.t334 37.4792
R3298 GNDA.n1128 GNDA.n1127 36.9067
R3299 GNDA.n909 GNDA.n908 36.6567
R3300 GNDA.n1642 GNDA.t225 34.8247
R3301 GNDA.n1932 GNDA.t225 34.8247
R3302 GNDA.n1910 GNDA.t225 34.8247
R3303 GNDA.t3 GNDA.n1165 34.4734
R3304 GNDA.n1168 GNDA.t115 34.4734
R3305 GNDA.t99 GNDA.t109 34.4734
R3306 GNDA.t109 GNDA.t187 34.4734
R3307 GNDA.n1848 GNDA.t55 34.4734
R3308 GNDA.n1848 GNDA.t116 34.4734
R3309 GNDA.t8 GNDA.t39 34.4734
R3310 GNDA.t39 GNDA.t185 34.4734
R3311 GNDA.n955 GNDA.t171 33.7313
R3312 GNDA.n957 GNDA.t348 33.7313
R3313 GNDA.n960 GNDA.t6 33.7313
R3314 GNDA.n959 GNDA.t51 33.7313
R3315 GNDA.n1111 GNDA.t33 33.7313
R3316 GNDA.n1055 GNDA.t339 33.6168
R3317 GNDA.n1159 GNDA.t80 33.6168
R3318 GNDA.t123 GNDA.t66 32.3951
R3319 GNDA.n375 GNDA.t227 31.6472
R3320 GNDA.t77 GNDA.n1210 31.3395
R3321 GNDA.n1220 GNDA.t194 31.3395
R3322 GNDA.t291 GNDA.t232 29.9835
R3323 GNDA.t211 GNDA.t251 29.9835
R3324 GNDA.t6 GNDA.t217 29.9835
R3325 GNDA.t139 GNDA.t200 29.9835
R3326 GNDA.t51 GNDA.t193 29.9835
R3327 GNDA.t297 GNDA.t278 29.9835
R3328 GNDA.n1046 GNDA.n1045 29.8817
R3329 GNDA.n1158 GNDA.n1152 29.8817
R3330 GNDA.n1179 GNDA.n1178 28.413
R3331 GNDA.n1031 GNDA.n970 28.413
R3332 GNDA.t262 GNDA.t76 28.2056
R3333 GNDA.t343 GNDA.t81 28.2056
R3334 GNDA.n1209 GNDA.t294 28.2056
R3335 GNDA.n1221 GNDA.t274 28.2056
R3336 GNDA.t70 GNDA.t53 28.2056
R3337 GNDA.t336 GNDA.t282 28.2056
R3338 GNDA.n1935 GNDA.n471 28.1318
R3339 GNDA.n1163 GNDA.n1162 28.038
R3340 GNDA.n980 GNDA.n964 28.038
R3341 GNDA.n1218 GNDA.n839 27.8193
R3342 GNDA.n1214 GNDA.n1213 27.8193
R3343 GNDA.n300 GNDA.n299 27.5561
R3344 GNDA.n1296 GNDA.n1295 27.5561
R3345 GNDA.n1730 GNDA.n1729 27.5561
R3346 GNDA.n2084 GNDA.n2083 27.5561
R3347 GNDA.n146 GNDA.n145 27.5561
R3348 GNDA.n566 GNDA.n565 27.5561
R3349 GNDA.n2240 GNDA.n2239 27.5561
R3350 GNDA.n728 GNDA.n727 27.5561
R3351 GNDA.n1404 GNDA.n1403 27.5561
R3352 GNDA.n0 GNDA.n46 8.60107
R3353 GNDA.n1871 GNDA.n1870 26.7261
R3354 GNDA.n1901 GNDA.n1895 26.7261
R3355 GNDA.n1110 GNDA.t103 26.2356
R3356 GNDA.t309 GNDA.n881 26.2356
R3357 GNDA.t85 GNDA.t106 26.1465
R3358 GNDA.t74 GNDA.t98 26.1465
R3359 GNDA.t207 GNDA.t72 26.1465
R3360 GNDA.t83 GNDA.t198 26.1465
R3361 GNDA.n877 GNDA.n876 25.6005
R3362 GNDA.n1053 GNDA.n1050 25.6005
R3363 GNDA.n1452 GNDA.t227 24.4846
R3364 GNDA.n1784 GNDA.t225 24.2965
R3365 GNDA.n808 GNDA.t100 24.0005
R3366 GNDA.n808 GNDA.t188 24.0005
R3367 GNDA.n806 GNDA.t82 24.0005
R3368 GNDA.n806 GNDA.t119 24.0005
R3369 GNDA.n804 GNDA.t346 24.0005
R3370 GNDA.n804 GNDA.t184 24.0005
R3371 GNDA.n802 GNDA.t147 24.0005
R3372 GNDA.n802 GNDA.t1 24.0005
R3373 GNDA.n800 GNDA.t145 24.0005
R3374 GNDA.n800 GNDA.t56 24.0005
R3375 GNDA.n798 GNDA.t117 24.0005
R3376 GNDA.n798 GNDA.t41 24.0005
R3377 GNDA.n796 GNDA.t69 24.0005
R3378 GNDA.n796 GNDA.t167 24.0005
R3379 GNDA.n794 GNDA.t102 24.0005
R3380 GNDA.n794 GNDA.t190 24.0005
R3381 GNDA.n792 GNDA.t43 24.0005
R3382 GNDA.n792 GNDA.t71 24.0005
R3383 GNDA.n791 GNDA.t9 24.0005
R3384 GNDA.n791 GNDA.t186 24.0005
R3385 GNDA.n314 GNDA.n235 23.6449
R3386 GNDA.n1278 GNDA.n1277 23.6449
R3387 GNDA.n1744 GNDA.n1666 23.6449
R3388 GNDA.n2098 GNDA.n2023 23.6449
R3389 GNDA.n160 GNDA.n81 23.6449
R3390 GNDA.n548 GNDA.n547 23.6449
R3391 GNDA.n2222 GNDA.n2221 23.6449
R3392 GNDA.n742 GNDA.n668 23.6449
R3393 GNDA.n1386 GNDA.n1385 23.6449
R3394 GNDA.n1836 GNDA.n1835 23.509
R3395 GNDA.n1148 GNDA.n1147 23.488
R3396 GNDA.t149 GNDA.t303 22.4877
R3397 GNDA.t177 GNDA.t4 22.4877
R3398 GNDA.t324 GNDA.t164 22.4877
R3399 GNDA.t57 GNDA.t12 22.4877
R3400 GNDA.t60 GNDA.t196 22.4877
R3401 GNDA.t326 GNDA.t159 22.4877
R3402 GNDA.t148 GNDA.t24 22.4877
R3403 GNDA.t143 GNDA.t120 22.4877
R3404 GNDA.t327 GNDA.t270 22.4877
R3405 GNDA.n1093 GNDA.n953 22.4005
R3406 GNDA.n1091 GNDA.n1090 22.4005
R3407 GNDA.n1087 GNDA.n1086 22.4005
R3408 GNDA.n1140 GNDA.n1139 22.4005
R3409 GNDA.n942 GNDA.n941 22.4005
R3410 GNDA.n943 GNDA.n942 22.4005
R3411 GNDA.n1173 GNDA.n1163 22.4005
R3412 GNDA.n1039 GNDA.n980 22.4005
R3413 GNDA.t195 GNDA.t118 21.9378
R3414 GNDA.t42 GNDA.t10 21.9378
R3415 GNDA.n1648 GNDA.t66 21.8669
R3416 GNDA.n1881 GNDA.t86 21.8669
R3417 GNDA.n1936 GNDA.n2 21.4917
R3418 GNDA.n1215 GNDA.n841 21.3338
R3419 GNDA.n1217 GNDA.n840 21.3338
R3420 GNDA.n838 GNDA.n828 21.3338
R3421 GNDA.n837 GNDA.n829 21.3338
R3422 GNDA.n1200 GNDA.n1199 21.3338
R3423 GNDA.n845 GNDA.n844 21.3338
R3424 GNDA.n944 GNDA.n936 21.3338
R3425 GNDA.n943 GNDA.n937 21.3338
R3426 GNDA.n941 GNDA.n938 21.3338
R3427 GNDA.n940 GNDA.n939 21.3338
R3428 GNDA.n885 GNDA.n884 21.3338
R3429 GNDA.n1105 GNDA.n1104 21.3338
R3430 GNDA.n1106 GNDA.n1103 21.3338
R3431 GNDA.n1102 GNDA.n946 21.3338
R3432 GNDA.n1101 GNDA.n947 21.3338
R3433 GNDA.n1100 GNDA.n948 21.3338
R3434 GNDA.n922 GNDA.n921 21.3338
R3435 GNDA.n924 GNDA.n923 21.3338
R3436 GNDA.n863 GNDA.n862 21.3338
R3437 GNDA.n1155 GNDA.n1153 21.3338
R3438 GNDA.n872 GNDA.n871 21.3338
R3439 GNDA.n878 GNDA.n875 21.3338
R3440 GNDA.n973 GNDA.n972 21.3338
R3441 GNDA.n976 GNDA.n975 21.3338
R3442 GNDA.n969 GNDA.n968 21.3338
R3443 GNDA.n1052 GNDA.n1051 21.3338
R3444 GNDA.n1201 GNDA.n1 21.1792
R3445 GNDA.n887 GNDA 20.281
R3446 GNDA.n1126 GNDA.t205 19.7005
R3447 GNDA.n1126 GNDA.t37 19.7005
R3448 GNDA.n1124 GNDA.t126 19.7005
R3449 GNDA.n1124 GNDA.t134 19.7005
R3450 GNDA.n1122 GNDA.t62 19.7005
R3451 GNDA.n1122 GNDA.t14 19.7005
R3452 GNDA.n1120 GNDA.t220 19.7005
R3453 GNDA.n1120 GNDA.t63 19.7005
R3454 GNDA.n1118 GNDA.t210 19.7005
R3455 GNDA.n1118 GNDA.t84 19.7005
R3456 GNDA.n1117 GNDA.t11 19.7005
R3457 GNDA.n1117 GNDA.t135 19.7005
R3458 GNDA.n907 GNDA.t335 19.7005
R3459 GNDA.n907 GNDA.t151 19.7005
R3460 GNDA.n905 GNDA.t340 19.7005
R3461 GNDA.n905 GNDA.t18 19.7005
R3462 GNDA.n903 GNDA.t330 19.7005
R3463 GNDA.n903 GNDA.t20 19.7005
R3464 GNDA.n901 GNDA.t132 19.7005
R3465 GNDA.n901 GNDA.t351 19.7005
R3466 GNDA.n899 GNDA.t142 19.7005
R3467 GNDA.n899 GNDA.t157 19.7005
R3468 GNDA.n898 GNDA.t338 19.7005
R3469 GNDA.n898 GNDA.t219 19.7005
R3470 GNDA.n790 GNDA.n789 19.4279
R3471 GNDA.n1000 GNDA.n859 19.3505
R3472 GNDA.n1022 GNDA.n986 19.3505
R3473 GNDA.n1108 GNDA.n1107 19.288
R3474 GNDA.n1876 GNDA.n470 19.2005
R3475 GNDA.n1936 GNDA.n469 19.2005
R3476 GNDA.n1617 GNDA.n775 19.2005
R3477 GNDA.n1921 GNDA.n1920 19.2005
R3478 GNDA.n1841 GNDA.n1840 19.2005
R3479 GNDA.n1194 GNDA.n1193 19.2005
R3480 GNDA.n876 GNDA.n864 19.1005
R3481 GNDA.n1050 GNDA.n1049 19.1005
R3482 GNDA.n930 GNDA.t155 18.7399
R3483 GNDA.n1860 GNDA.n1858 18.6274
R3484 GNDA.n812 GNDA.n790 18.3825
R3485 GNDA.n1842 GNDA.n1841 17.613
R3486 GNDA.n2516 GNDA.n2515 17.4917
R3487 GNDA.n2470 GNDA.n29 17.0672
R3488 GNDA.n1461 GNDA.n1460 17.0672
R3489 GNDA.n2417 GNDA.n61 17.0672
R3490 GNDA.n2511 GNDA.n2510 16.9605
R3491 GNDA.n247 GNDA.n246 16.0005
R3492 GNDA.n289 GNDA.n246 16.0005
R3493 GNDA.n290 GNDA.n289 16.0005
R3494 GNDA.n291 GNDA.n290 16.0005
R3495 GNDA.n291 GNDA.n244 16.0005
R3496 GNDA.n244 GNDA.n243 16.0005
R3497 GNDA.n298 GNDA.n243 16.0005
R3498 GNDA.n299 GNDA.n298 16.0005
R3499 GNDA.n314 GNDA.n313 16.0005
R3500 GNDA.n313 GNDA.n312 16.0005
R3501 GNDA.n312 GNDA.n237 16.0005
R3502 GNDA.n307 GNDA.n237 16.0005
R3503 GNDA.n307 GNDA.n306 16.0005
R3504 GNDA.n306 GNDA.n305 16.0005
R3505 GNDA.n305 GNDA.n240 16.0005
R3506 GNDA.n300 GNDA.n240 16.0005
R3507 GNDA.n330 GNDA.n227 16.0005
R3508 GNDA.n330 GNDA.n329 16.0005
R3509 GNDA.n329 GNDA.n328 16.0005
R3510 GNDA.n328 GNDA.n233 16.0005
R3511 GNDA.n322 GNDA.n233 16.0005
R3512 GNDA.n321 GNDA.n320 16.0005
R3513 GNDA.n320 GNDA.n235 16.0005
R3514 GNDA.n1310 GNDA.n1309 16.0005
R3515 GNDA.n1309 GNDA.n1308 16.0005
R3516 GNDA.n1308 GNDA.n1306 16.0005
R3517 GNDA.n1306 GNDA.n1303 16.0005
R3518 GNDA.n1303 GNDA.n1302 16.0005
R3519 GNDA.n1302 GNDA.n1299 16.0005
R3520 GNDA.n1299 GNDA.n1298 16.0005
R3521 GNDA.n1298 GNDA.n1296 16.0005
R3522 GNDA.n1281 GNDA.n1278 16.0005
R3523 GNDA.n1282 GNDA.n1281 16.0005
R3524 GNDA.n1285 GNDA.n1282 16.0005
R3525 GNDA.n1286 GNDA.n1285 16.0005
R3526 GNDA.n1289 GNDA.n1286 16.0005
R3527 GNDA.n1290 GNDA.n1289 16.0005
R3528 GNDA.n1293 GNDA.n1290 16.0005
R3529 GNDA.n1295 GNDA.n1293 16.0005
R3530 GNDA.n1262 GNDA.n1261 16.0005
R3531 GNDA.n1265 GNDA.n1262 16.0005
R3532 GNDA.n1266 GNDA.n1265 16.0005
R3533 GNDA.n1269 GNDA.n1266 16.0005
R3534 GNDA.n1270 GNDA.n1269 16.0005
R3535 GNDA.n1274 GNDA.n1273 16.0005
R3536 GNDA.n1277 GNDA.n1274 16.0005
R3537 GNDA.n1678 GNDA.n1677 16.0005
R3538 GNDA.n1719 GNDA.n1677 16.0005
R3539 GNDA.n1720 GNDA.n1719 16.0005
R3540 GNDA.n1721 GNDA.n1720 16.0005
R3541 GNDA.n1721 GNDA.n1675 16.0005
R3542 GNDA.n1675 GNDA.n1674 16.0005
R3543 GNDA.n1728 GNDA.n1674 16.0005
R3544 GNDA.n1729 GNDA.n1728 16.0005
R3545 GNDA.n1744 GNDA.n1743 16.0005
R3546 GNDA.n1743 GNDA.n1742 16.0005
R3547 GNDA.n1742 GNDA.n1668 16.0005
R3548 GNDA.n1737 GNDA.n1668 16.0005
R3549 GNDA.n1737 GNDA.n1736 16.0005
R3550 GNDA.n1736 GNDA.n1735 16.0005
R3551 GNDA.n1735 GNDA.n1671 16.0005
R3552 GNDA.n1730 GNDA.n1671 16.0005
R3553 GNDA.n1762 GNDA.n1761 16.0005
R3554 GNDA.n1761 GNDA.n1663 16.0005
R3555 GNDA.n1756 GNDA.n1663 16.0005
R3556 GNDA.n1756 GNDA.n1755 16.0005
R3557 GNDA.n1755 GNDA.n1754 16.0005
R3558 GNDA.n1750 GNDA.n1749 16.0005
R3559 GNDA.n1749 GNDA.n1666 16.0005
R3560 GNDA.n2035 GNDA.n2034 16.0005
R3561 GNDA.n2073 GNDA.n2034 16.0005
R3562 GNDA.n2074 GNDA.n2073 16.0005
R3563 GNDA.n2075 GNDA.n2074 16.0005
R3564 GNDA.n2075 GNDA.n2032 16.0005
R3565 GNDA.n2032 GNDA.n2031 16.0005
R3566 GNDA.n2082 GNDA.n2031 16.0005
R3567 GNDA.n2083 GNDA.n2082 16.0005
R3568 GNDA.n2098 GNDA.n2097 16.0005
R3569 GNDA.n2097 GNDA.n2096 16.0005
R3570 GNDA.n2096 GNDA.n2025 16.0005
R3571 GNDA.n2091 GNDA.n2025 16.0005
R3572 GNDA.n2091 GNDA.n2090 16.0005
R3573 GNDA.n2090 GNDA.n2089 16.0005
R3574 GNDA.n2089 GNDA.n2028 16.0005
R3575 GNDA.n2084 GNDA.n2028 16.0005
R3576 GNDA.n2116 GNDA.n2115 16.0005
R3577 GNDA.n2115 GNDA.n2020 16.0005
R3578 GNDA.n2110 GNDA.n2020 16.0005
R3579 GNDA.n2110 GNDA.n2109 16.0005
R3580 GNDA.n2109 GNDA.n2108 16.0005
R3581 GNDA.n2104 GNDA.n2103 16.0005
R3582 GNDA.n2103 GNDA.n2023 16.0005
R3583 GNDA.n93 GNDA.n92 16.0005
R3584 GNDA.n135 GNDA.n92 16.0005
R3585 GNDA.n136 GNDA.n135 16.0005
R3586 GNDA.n137 GNDA.n136 16.0005
R3587 GNDA.n137 GNDA.n90 16.0005
R3588 GNDA.n90 GNDA.n89 16.0005
R3589 GNDA.n144 GNDA.n89 16.0005
R3590 GNDA.n145 GNDA.n144 16.0005
R3591 GNDA.n160 GNDA.n159 16.0005
R3592 GNDA.n159 GNDA.n158 16.0005
R3593 GNDA.n158 GNDA.n83 16.0005
R3594 GNDA.n153 GNDA.n83 16.0005
R3595 GNDA.n153 GNDA.n152 16.0005
R3596 GNDA.n152 GNDA.n151 16.0005
R3597 GNDA.n151 GNDA.n86 16.0005
R3598 GNDA.n146 GNDA.n86 16.0005
R3599 GNDA.n176 GNDA.n73 16.0005
R3600 GNDA.n176 GNDA.n175 16.0005
R3601 GNDA.n175 GNDA.n174 16.0005
R3602 GNDA.n174 GNDA.n79 16.0005
R3603 GNDA.n168 GNDA.n79 16.0005
R3604 GNDA.n167 GNDA.n166 16.0005
R3605 GNDA.n166 GNDA.n81 16.0005
R3606 GNDA.n2511 GNDA.n3 16.0005
R3607 GNDA.n2515 GNDA.n3 16.0005
R3608 GNDA.n580 GNDA.n579 16.0005
R3609 GNDA.n579 GNDA.n578 16.0005
R3610 GNDA.n578 GNDA.n576 16.0005
R3611 GNDA.n576 GNDA.n573 16.0005
R3612 GNDA.n573 GNDA.n572 16.0005
R3613 GNDA.n572 GNDA.n569 16.0005
R3614 GNDA.n569 GNDA.n568 16.0005
R3615 GNDA.n568 GNDA.n566 16.0005
R3616 GNDA.n551 GNDA.n548 16.0005
R3617 GNDA.n552 GNDA.n551 16.0005
R3618 GNDA.n555 GNDA.n552 16.0005
R3619 GNDA.n556 GNDA.n555 16.0005
R3620 GNDA.n559 GNDA.n556 16.0005
R3621 GNDA.n560 GNDA.n559 16.0005
R3622 GNDA.n563 GNDA.n560 16.0005
R3623 GNDA.n565 GNDA.n563 16.0005
R3624 GNDA.n532 GNDA.n531 16.0005
R3625 GNDA.n535 GNDA.n532 16.0005
R3626 GNDA.n536 GNDA.n535 16.0005
R3627 GNDA.n539 GNDA.n536 16.0005
R3628 GNDA.n540 GNDA.n539 16.0005
R3629 GNDA.n544 GNDA.n543 16.0005
R3630 GNDA.n547 GNDA.n544 16.0005
R3631 GNDA.n2254 GNDA.n2253 16.0005
R3632 GNDA.n2253 GNDA.n2252 16.0005
R3633 GNDA.n2252 GNDA.n2250 16.0005
R3634 GNDA.n2250 GNDA.n2247 16.0005
R3635 GNDA.n2247 GNDA.n2246 16.0005
R3636 GNDA.n2246 GNDA.n2243 16.0005
R3637 GNDA.n2243 GNDA.n2242 16.0005
R3638 GNDA.n2242 GNDA.n2240 16.0005
R3639 GNDA.n2225 GNDA.n2222 16.0005
R3640 GNDA.n2226 GNDA.n2225 16.0005
R3641 GNDA.n2229 GNDA.n2226 16.0005
R3642 GNDA.n2230 GNDA.n2229 16.0005
R3643 GNDA.n2233 GNDA.n2230 16.0005
R3644 GNDA.n2234 GNDA.n2233 16.0005
R3645 GNDA.n2237 GNDA.n2234 16.0005
R3646 GNDA.n2239 GNDA.n2237 16.0005
R3647 GNDA.n2206 GNDA.n2157 16.0005
R3648 GNDA.n2209 GNDA.n2206 16.0005
R3649 GNDA.n2210 GNDA.n2209 16.0005
R3650 GNDA.n2213 GNDA.n2210 16.0005
R3651 GNDA.n2214 GNDA.n2213 16.0005
R3652 GNDA.n2218 GNDA.n2217 16.0005
R3653 GNDA.n2221 GNDA.n2218 16.0005
R3654 GNDA.n680 GNDA.n679 16.0005
R3655 GNDA.n717 GNDA.n679 16.0005
R3656 GNDA.n718 GNDA.n717 16.0005
R3657 GNDA.n719 GNDA.n718 16.0005
R3658 GNDA.n719 GNDA.n677 16.0005
R3659 GNDA.n677 GNDA.n676 16.0005
R3660 GNDA.n726 GNDA.n676 16.0005
R3661 GNDA.n727 GNDA.n726 16.0005
R3662 GNDA.n742 GNDA.n741 16.0005
R3663 GNDA.n741 GNDA.n740 16.0005
R3664 GNDA.n740 GNDA.n670 16.0005
R3665 GNDA.n735 GNDA.n670 16.0005
R3666 GNDA.n735 GNDA.n734 16.0005
R3667 GNDA.n734 GNDA.n733 16.0005
R3668 GNDA.n733 GNDA.n673 16.0005
R3669 GNDA.n728 GNDA.n673 16.0005
R3670 GNDA.n760 GNDA.n759 16.0005
R3671 GNDA.n759 GNDA.n665 16.0005
R3672 GNDA.n754 GNDA.n665 16.0005
R3673 GNDA.n754 GNDA.n753 16.0005
R3674 GNDA.n753 GNDA.n752 16.0005
R3675 GNDA.n748 GNDA.n747 16.0005
R3676 GNDA.n747 GNDA.n668 16.0005
R3677 GNDA.n1418 GNDA.n1417 16.0005
R3678 GNDA.n1417 GNDA.n1416 16.0005
R3679 GNDA.n1416 GNDA.n1414 16.0005
R3680 GNDA.n1414 GNDA.n1411 16.0005
R3681 GNDA.n1411 GNDA.n1410 16.0005
R3682 GNDA.n1410 GNDA.n1407 16.0005
R3683 GNDA.n1407 GNDA.n1406 16.0005
R3684 GNDA.n1406 GNDA.n1404 16.0005
R3685 GNDA.n1389 GNDA.n1386 16.0005
R3686 GNDA.n1390 GNDA.n1389 16.0005
R3687 GNDA.n1393 GNDA.n1390 16.0005
R3688 GNDA.n1394 GNDA.n1393 16.0005
R3689 GNDA.n1397 GNDA.n1394 16.0005
R3690 GNDA.n1398 GNDA.n1397 16.0005
R3691 GNDA.n1401 GNDA.n1398 16.0005
R3692 GNDA.n1403 GNDA.n1401 16.0005
R3693 GNDA.n1370 GNDA.n1369 16.0005
R3694 GNDA.n1373 GNDA.n1370 16.0005
R3695 GNDA.n1374 GNDA.n1373 16.0005
R3696 GNDA.n1377 GNDA.n1374 16.0005
R3697 GNDA.n1378 GNDA.n1377 16.0005
R3698 GNDA.n1382 GNDA.n1381 16.0005
R3699 GNDA.n1385 GNDA.n1382 16.0005
R3700 GNDA.t78 GNDA.t345 15.67
R3701 GNDA.t183 GNDA.t45 15.67
R3702 GNDA.t101 GNDA.t154 15.67
R3703 GNDA.t32 GNDA.t189 15.67
R3704 GNDA.n2297 GNDA.n380 15.5383
R3705 GNDA.n2394 GNDA.n2393 15.5383
R3706 GNDA.n414 GNDA.n370 15.5383
R3707 GNDA.n2353 GNDA.n2352 15.5383
R3708 GNDA.n1223 GNDA.n786 15.363
R3709 GNDA.n1207 GNDA.n786 15.363
R3710 GNDA.t329 GNDA.t291 14.992
R3711 GNDA.t28 GNDA.t211 14.992
R3712 GNDA.t217 GNDA.t201 14.992
R3713 GNDA.t200 GNDA.t325 14.992
R3714 GNDA.t193 GNDA.t323 14.992
R3715 GNDA.t64 GNDA.t306 14.992
R3716 GNDA.t306 GNDA.t108 14.992
R3717 GNDA.t108 GNDA.t168 14.992
R3718 GNDA.t130 GNDA.t202 14.992
R3719 GNDA.t202 GNDA.t23 14.992
R3720 GNDA.t212 GNDA.t30 14.992
R3721 GNDA.t30 GNDA.t347 14.992
R3722 GNDA.t347 GNDA.t333 14.992
R3723 GNDA.t180 GNDA.t161 14.992
R3724 GNDA.t161 GNDA.t93 14.992
R3725 GNDA.t93 GNDA.t222 14.992
R3726 GNDA.t110 GNDA.t352 14.992
R3727 GNDA.t352 GNDA.t322 14.992
R3728 GNDA.t137 GNDA.t58 14.992
R3729 GNDA.t58 GNDA.t158 14.992
R3730 GNDA.t174 GNDA.t26 14.992
R3731 GNDA.t26 GNDA.t320 14.992
R3732 GNDA.t163 GNDA.t103 14.992
R3733 GNDA.t33 GNDA.t47 14.992
R3734 GNDA.t278 GNDA.t88 14.992
R3735 GNDA.t303 GNDA.t191 14.992
R3736 GNDA.t331 GNDA.t204 14.992
R3737 GNDA.t355 GNDA.t177 14.992
R3738 GNDA.t2 GNDA.t324 14.992
R3739 GNDA.t218 GNDA.t57 14.992
R3740 GNDA.t192 GNDA.t60 14.992
R3741 GNDA.t16 GNDA.t326 14.992
R3742 GNDA.t312 GNDA.t148 14.992
R3743 GNDA.n1045 GNDA.n949 14.9411
R3744 GNDA.n1143 GNDA.n873 14.0505
R3745 GNDA.n1058 GNDA.n1057 14.0505
R3746 GNDA.n1130 GNDA.n1129 14.0193
R3747 GNDA.n427 GNDA.n375 13.9984
R3748 GNDA.n1193 GNDA.n813 13.8005
R3749 GNDA.n1090 GNDA.n1089 13.8005
R3750 GNDA.n1141 GNDA.n1140 13.8005
R3751 GNDA.n1088 GNDA.n1087 13.8005
R3752 GNDA.n1062 GNDA.n953 13.8005
R3753 GNDA.n1627 GNDA.n1626 13.7682
R3754 GNDA.n1918 GNDA.n1917 13.7682
R3755 GNDA.n2517 GNDA.n2516 13.4945
R3756 GNDA GNDA.n321 12.9783
R3757 GNDA.n1273 GNDA 12.9783
R3758 GNDA.n1750 GNDA 12.9783
R3759 GNDA.n2104 GNDA 12.9783
R3760 GNDA GNDA.n167 12.9783
R3761 GNDA.n543 GNDA 12.9783
R3762 GNDA.n2217 GNDA 12.9783
R3763 GNDA.n748 GNDA 12.9783
R3764 GNDA.n1381 GNDA 12.9783
R3765 GNDA.t86 GNDA.n1880 12.9584
R3766 GNDA.n860 GNDA.n859 12.8005
R3767 GNDA.n986 GNDA.n985 12.8005
R3768 GNDA.n1198 GNDA.n1196 12.5361
R3769 GNDA.n832 GNDA.n831 12.5361
R3770 GNDA.n1898 GNDA.n463 12.4126
R3771 GNDA.n644 GNDA.n504 12.4126
R3772 GNDA.n1630 GNDA.n1612 12.4126
R3773 GNDA.n2447 GNDA.n36 11.6369
R3774 GNDA.n2454 GNDA.n36 11.6369
R3775 GNDA.n2455 GNDA.n2454 11.6369
R3776 GNDA.n2456 GNDA.n2455 11.6369
R3777 GNDA.n2456 GNDA.n33 11.6369
R3778 GNDA.n2462 GNDA.n33 11.6369
R3779 GNDA.n2463 GNDA.n2462 11.6369
R3780 GNDA.n2464 GNDA.n2463 11.6369
R3781 GNDA.n2464 GNDA.n29 11.6369
R3782 GNDA.n1915 GNDA.n1914 11.6369
R3783 GNDA.n1914 GNDA.n1913 11.6369
R3784 GNDA.n1913 GNDA.n1888 11.6369
R3785 GNDA.n1907 GNDA.n1888 11.6369
R3786 GNDA.n1906 GNDA.n1905 11.6369
R3787 GNDA.n1905 GNDA.n1892 11.6369
R3788 GNDA.n1899 GNDA.n1892 11.6369
R3789 GNDA.n1899 GNDA.n1898 11.6369
R3790 GNDA.n1944 GNDA.n1943 11.6369
R3791 GNDA.n1945 GNDA.n1944 11.6369
R3792 GNDA.n1945 GNDA.n459 11.6369
R3793 GNDA.n1952 GNDA.n459 11.6369
R3794 GNDA.n1953 GNDA.n1952 11.6369
R3795 GNDA.n1954 GNDA.n1953 11.6369
R3796 GNDA.n1954 GNDA.n456 11.6369
R3797 GNDA.n1960 GNDA.n456 11.6369
R3798 GNDA.n1961 GNDA.n1960 11.6369
R3799 GNDA.n1963 GNDA.n1961 11.6369
R3800 GNDA.n1963 GNDA.n1962 11.6369
R3801 GNDA.n1978 GNDA.n1970 11.6369
R3802 GNDA.n1978 GNDA.n1977 11.6369
R3803 GNDA.n1977 GNDA.n1976 11.6369
R3804 GNDA.n1976 GNDA.n1971 11.6369
R3805 GNDA.n1971 GNDA.n6 11.6369
R3806 GNDA.n2509 GNDA.n7 11.6369
R3807 GNDA.n2503 GNDA.n7 11.6369
R3808 GNDA.n2503 GNDA.n2502 11.6369
R3809 GNDA.n2502 GNDA.n2501 11.6369
R3810 GNDA.n2501 GNDA.n12 11.6369
R3811 GNDA.n2488 GNDA.n20 11.6369
R3812 GNDA.n2488 GNDA.n2487 11.6369
R3813 GNDA.n2487 GNDA.n2486 11.6369
R3814 GNDA.n2486 GNDA.n21 11.6369
R3815 GNDA.n2480 GNDA.n21 11.6369
R3816 GNDA.n2480 GNDA.n2479 11.6369
R3817 GNDA.n2479 GNDA.n2478 11.6369
R3818 GNDA.n2478 GNDA.n24 11.6369
R3819 GNDA.n2472 GNDA.n24 11.6369
R3820 GNDA.n2472 GNDA.n2471 11.6369
R3821 GNDA.n2471 GNDA.n2470 11.6369
R3822 GNDA.n2304 GNDA.n2303 11.6369
R3823 GNDA.n2307 GNDA.n2304 11.6369
R3824 GNDA.n2308 GNDA.n2307 11.6369
R3825 GNDA.n2311 GNDA.n2308 11.6369
R3826 GNDA.n2312 GNDA.n2311 11.6369
R3827 GNDA.n2315 GNDA.n2312 11.6369
R3828 GNDA.n2317 GNDA.n2315 11.6369
R3829 GNDA.n2318 GNDA.n2317 11.6369
R3830 GNDA.n2320 GNDA.n2318 11.6369
R3831 GNDA.n2320 GNDA.n2319 11.6369
R3832 GNDA.n2319 GNDA.n69 11.6369
R3833 GNDA.n1868 GNDA.n1867 11.6369
R3834 GNDA.n1868 GNDA.n475 11.6369
R3835 GNDA.n1930 GNDA.n475 11.6369
R3836 GNDA.n1930 GNDA.n1929 11.6369
R3837 GNDA.n1928 GNDA.n476 11.6369
R3838 GNDA.n499 GNDA.n476 11.6369
R3839 GNDA.n503 GNDA.n499 11.6369
R3840 GNDA.n504 GNDA.n503 11.6369
R3841 GNDA.n643 GNDA.n642 11.6369
R3842 GNDA.n642 GNDA.n505 11.6369
R3843 GNDA.n601 GNDA.n505 11.6369
R3844 GNDA.n602 GNDA.n601 11.6369
R3845 GNDA.n603 GNDA.n602 11.6369
R3846 GNDA.n603 GNDA.n587 11.6369
R3847 GNDA.n623 GNDA.n587 11.6369
R3848 GNDA.n624 GNDA.n623 11.6369
R3849 GNDA.n626 GNDA.n624 11.6369
R3850 GNDA.n626 GNDA.n625 11.6369
R3851 GNDA.n625 GNDA.n409 11.6369
R3852 GNDA.n1505 GNDA.n1450 11.6369
R3853 GNDA.n1505 GNDA.n1504 11.6369
R3854 GNDA.n1504 GNDA.n1503 11.6369
R3855 GNDA.n1503 GNDA.n1455 11.6369
R3856 GNDA.n1459 GNDA.n1455 11.6369
R3857 GNDA.n1495 GNDA.n1459 11.6369
R3858 GNDA.n1495 GNDA.n1494 11.6369
R3859 GNDA.n1494 GNDA.n1493 11.6369
R3860 GNDA.n1493 GNDA.n1460 11.6369
R3861 GNDA.n1789 GNDA.n1788 11.6369
R3862 GNDA.n1792 GNDA.n1789 11.6369
R3863 GNDA.n1793 GNDA.n1792 11.6369
R3864 GNDA.n1796 GNDA.n1793 11.6369
R3865 GNDA.n1797 GNDA.n1796 11.6369
R3866 GNDA.n1800 GNDA.n1797 11.6369
R3867 GNDA.n1802 GNDA.n1800 11.6369
R3868 GNDA.n1803 GNDA.n1802 11.6369
R3869 GNDA.n1805 GNDA.n1803 11.6369
R3870 GNDA.n1805 GNDA.n1804 11.6369
R3871 GNDA.n1804 GNDA.n379 11.6369
R3872 GNDA.n1646 GNDA.n1620 11.6369
R3873 GNDA.n1646 GNDA.n1645 11.6369
R3874 GNDA.n1645 GNDA.n1644 11.6369
R3875 GNDA.n1644 GNDA.n1624 11.6369
R3876 GNDA.n1638 GNDA.n1637 11.6369
R3877 GNDA.n1637 GNDA.n1636 11.6369
R3878 GNDA.n1636 GNDA.n1631 11.6369
R3879 GNDA.n1631 GNDA.n1630 11.6369
R3880 GNDA.n2296 GNDA.n2295 11.6369
R3881 GNDA.n2295 GNDA.n381 11.6369
R3882 GNDA.n2290 GNDA.n381 11.6369
R3883 GNDA.n2290 GNDA.n2289 11.6369
R3884 GNDA.n2289 GNDA.n2288 11.6369
R3885 GNDA.n2288 GNDA.n2275 11.6369
R3886 GNDA.n2283 GNDA.n2275 11.6369
R3887 GNDA.n2283 GNDA.n2282 11.6369
R3888 GNDA.n2282 GNDA.n2281 11.6369
R3889 GNDA.n2281 GNDA.n223 11.6369
R3890 GNDA.n2354 GNDA.n223 11.6369
R3891 GNDA.n1469 GNDA.n224 11.6369
R3892 GNDA.n1470 GNDA.n1469 11.6369
R3893 GNDA.n1470 GNDA.n1465 11.6369
R3894 GNDA.n1476 GNDA.n1465 11.6369
R3895 GNDA.n1477 GNDA.n1476 11.6369
R3896 GNDA.n1478 GNDA.n1477 11.6369
R3897 GNDA.n1478 GNDA.n1463 11.6369
R3898 GNDA.n1484 GNDA.n1463 11.6369
R3899 GNDA.n1485 GNDA.n1484 11.6369
R3900 GNDA.n1486 GNDA.n1485 11.6369
R3901 GNDA.n1486 GNDA.n1461 11.6369
R3902 GNDA.n2438 GNDA.n53 11.6369
R3903 GNDA.n2432 GNDA.n53 11.6369
R3904 GNDA.n2432 GNDA.n2431 11.6369
R3905 GNDA.n2431 GNDA.n2430 11.6369
R3906 GNDA.n2430 GNDA.n57 11.6369
R3907 GNDA.n2424 GNDA.n57 11.6369
R3908 GNDA.n2424 GNDA.n2423 11.6369
R3909 GNDA.n2423 GNDA.n2422 11.6369
R3910 GNDA.n2422 GNDA.n61 11.6369
R3911 GNDA.n2395 GNDA.n67 11.6369
R3912 GNDA.n2401 GNDA.n67 11.6369
R3913 GNDA.n2402 GNDA.n2401 11.6369
R3914 GNDA.n2403 GNDA.n2402 11.6369
R3915 GNDA.n2403 GNDA.n65 11.6369
R3916 GNDA.n2409 GNDA.n65 11.6369
R3917 GNDA.n2410 GNDA.n2409 11.6369
R3918 GNDA.n2411 GNDA.n2410 11.6369
R3919 GNDA.n2411 GNDA.n63 11.6369
R3920 GNDA.n2416 GNDA.n63 11.6369
R3921 GNDA.n2417 GNDA.n2416 11.6369
R3922 GNDA.n1061 GNDA.n909 11.6255
R3923 GNDA.n1915 GNDA.n1887 11.3514
R3924 GNDA.n1867 GNDA.n1866 11.3514
R3925 GNDA.n1653 GNDA.n1620 11.3514
R3926 GNDA.n1880 GNDA.t95 11.3386
R3927 GNDA.n2447 GNDA.n2446 11.249
R3928 GNDA.n1512 GNDA.n1450 11.249
R3929 GNDA.n2439 GNDA.n2438 11.249
R3930 GNDA.t328 GNDA.n957 11.2441
R3931 GNDA.t23 GNDA.n958 11.2441
R3932 GNDA.t169 GNDA.n1134 11.2441
R3933 GNDA.n1134 GNDA.t204 11.2441
R3934 GNDA.t38 GNDA.t29 11.2441
R3935 GNDA.n932 GNDA.t143 11.2441
R3936 GNDA.t256 GNDA.n1043 11.2059
R3937 GNDA.t22 GNDA.t300 11.2059
R3938 GNDA.t49 GNDA.t105 11.2059
R3939 GNDA.t206 GNDA.t91 11.2059
R3940 GNDA.t133 GNDA.t235 11.2059
R3941 GNDA.t259 GNDA.n867 11.2059
R3942 GNDA.n1925 GNDA.n1924 10.5288
R3943 GNDA.n2510 GNDA.n2509 10.4732
R3944 GNDA GNDA.n1906 10.3439
R3945 GNDA GNDA.n1928 10.3439
R3946 GNDA.n1638 GNDA 10.3439
R3947 GNDA.n1844 GNDA.n1843 9.78488
R3948 GNDA.n814 GNDA.t216 9.6005
R3949 GNDA.n814 GNDA.t114 9.6005
R3950 GNDA.n1192 GNDA.t215 9.6005
R3951 GNDA.n1192 GNDA.t113 9.6005
R3952 GNDA.n1063 GNDA.t243 9.6005
R3953 GNDA.n1063 GNDA.t349 9.6005
R3954 GNDA.t307 GNDA.n1084 9.6005
R3955 GNDA.n1084 GNDA.t203 9.6005
R3956 GNDA.n1081 GNDA.t31 9.6005
R3957 GNDA.n1081 GNDA.t162 9.6005
R3958 GNDA.n1079 GNDA.t353 9.6005
R3959 GNDA.n1079 GNDA.t59 9.6005
R3960 GNDA.n1077 GNDA.t27 9.6005
R3961 GNDA.n1077 GNDA.t104 9.6005
R3962 GNDA.n1075 GNDA.t34 9.6005
R3963 GNDA.n1075 GNDA.t89 9.6005
R3964 GNDA.n1073 GNDA.t173 9.6005
R3965 GNDA.n1073 GNDA.t150 9.6005
R3966 GNDA.n1071 GNDA.t170 9.6005
R3967 GNDA.n1071 GNDA.t5 9.6005
R3968 GNDA.n1069 GNDA.t165 9.6005
R3969 GNDA.n1069 GNDA.t13 9.6005
R3970 GNDA.n1067 GNDA.t156 9.6005
R3971 GNDA.n1067 GNDA.t197 9.6005
R3972 GNDA.n1065 GNDA.t160 9.6005
R3973 GNDA.n1065 GNDA.t25 9.6005
R3974 GNDA.n888 GNDA.t121 9.6005
R3975 GNDA.n888 GNDA.t271 9.6005
R3976 GNDA.t79 GNDA.t183 9.40221
R3977 GNDA.t354 GNDA.t101 9.40221
R3978 GNDA.n813 GNDA.n812 9.37925
R3979 GNDA.n1115 GNDA.n1114 9.3005
R3980 GNDA.n2300 GNDA.n375 8.98697
R3981 GNDA.n1943 GNDA.n463 8.79242
R3982 GNDA.n644 GNDA.n643 8.79242
R3983 GNDA.n1788 GNDA.n1612 8.79242
R3984 GNDA.n1970 GNDA.n452 8.53383
R3985 GNDA.n20 GNDA.n16 8.53383
R3986 GNDA.n2303 GNDA.n370 8.53383
R3987 GNDA.n2297 GNDA.n2296 8.53383
R3988 GNDA.n2353 GNDA.n224 8.53383
R3989 GNDA.n2395 GNDA.n2394 8.53383
R3990 GNDA.n810 GNDA.n809 8.44175
R3991 GNDA.n250 GNDA.n247 8.35606
R3992 GNDA.n1311 GNDA.n1310 8.35606
R3993 GNDA.n1678 GNDA.n1233 8.35606
R3994 GNDA.n2062 GNDA.n2035 8.35606
R3995 GNDA.n96 GNDA.n93 8.35606
R3996 GNDA.n580 GNDA.n413 8.35606
R3997 GNDA.n2256 GNDA.n2254 8.35606
R3998 GNDA.n706 GNDA.n680 8.35606
R3999 GNDA.n1419 GNDA.n1418 8.35606
R4000 GNDA.n1835 GNDA.t225 8.20508
R4001 GNDA.n1967 GNDA.t227 8.20508
R4002 GNDA.n1843 GNDA.n786 7.71925
R4003 GNDA.n1918 GNDA.t44 7.28929
R4004 GNDA.n470 GNDA.n468 6.4005
R4005 GNDA GNDA.n2517 5.86508
R4006 GNDA.t95 GNDA.t44 5.66956
R4007 GNDA.n1129 GNDA.n1116 5.03175
R4008 GNDA.n1116 GNDA.n909 4.90675
R4009 GNDA.n1626 GNDA.t123 4.85969
R4010 GNDA.n1116 GNDA.n1115 4.7505
R4011 GNDA.n1886 GNDA.n493 4.6085
R4012 GNDA.n1865 GNDA.n652 4.6085
R4013 GNDA.n1775 GNDA.n1774 4.6085
R4014 GNDA.n1985 GNDA.n1984 4.55161
R4015 GNDA.n2495 GNDA.n2494 4.55161
R4016 GNDA.n2134 GNDA.n372 4.55161
R4017 GNDA.n2298 GNDA.n378 4.55161
R4018 GNDA.n2357 GNDA.n220 4.55161
R4019 GNDA.n2327 GNDA.n70 4.55161
R4020 GNDA.n1843 GNDA.n1842 4.5005
R4021 GNDA.n918 GNDA.n916 4.5005
R4022 GNDA.n1128 GNDA.n887 4.5005
R4023 GNDA.n1147 GNDA.n1146 4.5005
R4024 GNDA.n1962 GNDA.n452 4.39646
R4025 GNDA.n16 GNDA.n12 4.39646
R4026 GNDA.n2394 GNDA.n69 4.39646
R4027 GNDA.n409 GNDA.n370 4.39646
R4028 GNDA.n2297 GNDA.n379 4.39646
R4029 GNDA.n2354 GNDA.n2353 4.39646
R4030 GNDA.n2446 GNDA.n40 4.3013
R4031 GNDA.n2439 GNDA.n52 4.3013
R4032 GNDA.n2004 GNDA.n415 4.26717
R4033 GNDA.n2004 GNDA.n429 4.26717
R4034 GNDA.n1999 GNDA.n429 4.26717
R4035 GNDA.n1999 GNDA.n1998 4.26717
R4036 GNDA.n1998 GNDA.n1997 4.26717
R4037 GNDA.n1997 GNDA.n437 4.26717
R4038 GNDA.n1992 GNDA.n1991 4.26717
R4039 GNDA.n1991 GNDA.n1990 4.26717
R4040 GNDA.n1990 GNDA.n446 4.26717
R4041 GNDA.n1985 GNDA.n446 4.26717
R4042 GNDA.n2389 GNDA.n192 4.26717
R4043 GNDA.n195 GNDA.n192 4.26717
R4044 GNDA.n2382 GNDA.n195 4.26717
R4045 GNDA.n2382 GNDA.n2381 4.26717
R4046 GNDA.n2381 GNDA.n2380 4.26717
R4047 GNDA.n2380 GNDA.n200 4.26717
R4048 GNDA.n2375 GNDA.n2374 4.26717
R4049 GNDA.n2374 GNDA.n2373 4.26717
R4050 GNDA.n2373 GNDA.n14 4.26717
R4051 GNDA.n2495 GNDA.n14 4.26717
R4052 GNDA.n2155 GNDA.n392 4.26717
R4053 GNDA.n395 GNDA.n392 4.26717
R4054 GNDA.n2148 GNDA.n395 4.26717
R4055 GNDA.n2148 GNDA.n2147 4.26717
R4056 GNDA.n2147 GNDA.n2146 4.26717
R4057 GNDA.n2146 GNDA.n400 4.26717
R4058 GNDA.n2141 GNDA.n2140 4.26717
R4059 GNDA.n2140 GNDA.n2139 4.26717
R4060 GNDA.n2139 GNDA.n406 4.26717
R4061 GNDA.n2134 GNDA.n406 4.26717
R4062 GNDA.n1830 GNDA.n1829 4.26717
R4063 GNDA.n1829 GNDA.n1584 4.26717
R4064 GNDA.n1824 GNDA.n1584 4.26717
R4065 GNDA.n1824 GNDA.n1823 4.26717
R4066 GNDA.n1823 GNDA.n1822 4.26717
R4067 GNDA.n1822 GNDA.n1593 4.26717
R4068 GNDA.n1817 GNDA.n1816 4.26717
R4069 GNDA.n1816 GNDA.n1815 4.26717
R4070 GNDA.n1815 GNDA.n1604 4.26717
R4071 GNDA.n1604 GNDA.n378 4.26717
R4072 GNDA.n1563 GNDA.n1562 4.26717
R4073 GNDA.n1562 GNDA.n1532 4.26717
R4074 GNDA.n1557 GNDA.n1532 4.26717
R4075 GNDA.n1557 GNDA.n1556 4.26717
R4076 GNDA.n1556 GNDA.n1555 4.26717
R4077 GNDA.n1555 GNDA.n1539 4.26717
R4078 GNDA.n1550 GNDA.n1549 4.26717
R4079 GNDA.n1549 GNDA.n1548 4.26717
R4080 GNDA.n1548 GNDA.n219 4.26717
R4081 GNDA.n2357 GNDA.n219 4.26717
R4082 GNDA.n2348 GNDA.n345 4.26717
R4083 GNDA.n349 GNDA.n345 4.26717
R4084 GNDA.n2341 GNDA.n349 4.26717
R4085 GNDA.n2341 GNDA.n2340 4.26717
R4086 GNDA.n2340 GNDA.n2339 4.26717
R4087 GNDA.n2339 GNDA.n355 4.26717
R4088 GNDA.n2334 GNDA.n2333 4.26717
R4089 GNDA.n2333 GNDA.n2332 4.26717
R4090 GNDA.n2332 GNDA.n362 4.26717
R4091 GNDA.n2327 GNDA.n362 4.26717
R4092 GNDA.n1513 GNDA.n1512 4.1989
R4093 GNDA.n1842 GNDA.n813 3.813
R4094 GNDA.n1992 GNDA 3.79309
R4095 GNDA.n2375 GNDA 3.79309
R4096 GNDA.n2141 GNDA 3.79309
R4097 GNDA.n1817 GNDA 3.79309
R4098 GNDA.n1550 GNDA 3.79309
R4099 GNDA.n2334 GNDA 3.79309
R4100 GNDA.n954 GNDA.t242 3.74837
R4101 GNDA.t348 GNDA.n955 3.74837
R4102 GNDA.n960 GNDA.t28 3.74837
R4103 GNDA.t325 GNDA.n959 3.74837
R4104 GNDA.n958 GNDA.t94 3.74837
R4105 GNDA.n1111 GNDA.t297 3.74837
R4106 GNDA.n1135 GNDA.t35 3.74837
R4107 GNDA.t332 GNDA.n930 3.74837
R4108 GNDA.t29 GNDA.t332 3.74837
R4109 GNDA.n1035 GNDA.t136 3.73564
R4110 GNDA.n1034 GNDA.t350 3.73564
R4111 GNDA.t267 GNDA.t285 3.73564
R4112 GNDA.t248 GNDA.t245 3.73564
R4113 GNDA.n1129 GNDA.n1128 3.6255
R4114 GNDA.n184 GNDA.n74 3.5845
R4115 GNDA.n183 GNDA.n76 3.5845
R4116 GNDA.n106 GNDA.n104 3.5845
R4117 GNDA.n105 GNDA.n102 3.5845
R4118 GNDA.n113 GNDA.n112 3.5845
R4119 GNDA.n99 GNDA.n98 3.5845
R4120 GNDA.n121 GNDA.n119 3.5845
R4121 GNDA.n120 GNDA.n95 3.5845
R4122 GNDA.n128 GNDA.n127 3.5845
R4123 GNDA.n637 GNDA.n511 3.5845
R4124 GNDA.n595 GNDA.n594 3.5845
R4125 GNDA.n608 GNDA.n593 3.5845
R4126 GNDA.n609 GNDA.n591 3.5845
R4127 GNDA.n613 GNDA.n612 3.5845
R4128 GNDA.n619 GNDA.n614 3.5845
R4129 GNDA.n618 GNDA.n615 3.5845
R4130 GNDA.n630 GNDA.n583 3.5845
R4131 GNDA.n632 GNDA.n631 3.5845
R4132 GNDA.n2122 GNDA.n2016 3.5845
R4133 GNDA.n2121 GNDA.n2017 3.5845
R4134 GNDA.n2045 GNDA.n2043 3.5845
R4135 GNDA.n2049 GNDA.n2046 3.5845
R4136 GNDA.n2050 GNDA.n2038 3.5845
R4137 GNDA.n2055 GNDA.n2054 3.5845
R4138 GNDA.n2058 GNDA.n2037 3.5845
R4139 GNDA.n2060 GNDA.n2059 3.5845
R4140 GNDA.n2066 GNDA.n2065 3.5845
R4141 GNDA.n766 GNDA.n659 3.5845
R4142 GNDA.n765 GNDA.n660 3.5845
R4143 GNDA.n690 GNDA.n688 3.5845
R4144 GNDA.n694 GNDA.n691 3.5845
R4145 GNDA.n695 GNDA.n683 3.5845
R4146 GNDA.n700 GNDA.n699 3.5845
R4147 GNDA.n703 GNDA.n682 3.5845
R4148 GNDA.n705 GNDA.n704 3.5845
R4149 GNDA.n710 GNDA.n709 3.5845
R4150 GNDA.n2265 GNDA.n2159 3.5845
R4151 GNDA.n2186 GNDA.n2185 3.5845
R4152 GNDA.n2189 GNDA.n2184 3.5845
R4153 GNDA.n2193 GNDA.n2192 3.5845
R4154 GNDA.n2196 GNDA.n2182 3.5845
R4155 GNDA.n2200 GNDA.n2199 3.5845
R4156 GNDA.n2203 GNDA.n2181 3.5845
R4157 GNDA.n2205 GNDA.n2204 3.5845
R4158 GNDA.n2260 GNDA.n2259 3.5845
R4159 GNDA.n1523 GNDA.n1346 3.5845
R4160 GNDA.n1427 GNDA.n1426 3.5845
R4161 GNDA.n1433 GNDA.n1429 3.5845
R4162 GNDA.n1432 GNDA.n1423 3.5845
R4163 GNDA.n1439 GNDA.n1422 3.5845
R4164 GNDA.n1440 GNDA.n1421 3.5845
R4165 GNDA.n1445 GNDA.n1443 3.5845
R4166 GNDA.n1444 GNDA.n1368 3.5845
R4167 GNDA.n1518 GNDA.n1517 3.5845
R4168 GNDA.n1768 GNDA.n1659 3.5845
R4169 GNDA.n1767 GNDA.n1660 3.5845
R4170 GNDA.n1690 GNDA.n1689 3.5845
R4171 GNDA.n1695 GNDA.n1688 3.5845
R4172 GNDA.n1697 GNDA.n1696 3.5845
R4173 GNDA.n1704 GNDA.n1684 3.5845
R4174 GNDA.n1703 GNDA.n1685 3.5845
R4175 GNDA.n1710 GNDA.n1680 3.5845
R4176 GNDA.n1712 GNDA.n1711 3.5845
R4177 GNDA.n1575 GNDA.n1238 3.5845
R4178 GNDA.n1319 GNDA.n1318 3.5845
R4179 GNDA.n1325 GNDA.n1321 3.5845
R4180 GNDA.n1324 GNDA.n1315 3.5845
R4181 GNDA.n1331 GNDA.n1314 3.5845
R4182 GNDA.n1332 GNDA.n1313 3.5845
R4183 GNDA.n1337 GNDA.n1335 3.5845
R4184 GNDA.n1336 GNDA.n1260 3.5845
R4185 GNDA.n1570 GNDA.n1569 3.5845
R4186 GNDA.n338 GNDA.n228 3.5845
R4187 GNDA.n337 GNDA.n230 3.5845
R4188 GNDA.n260 GNDA.n258 3.5845
R4189 GNDA.n259 GNDA.n256 3.5845
R4190 GNDA.n267 GNDA.n266 3.5845
R4191 GNDA.n253 GNDA.n252 3.5845
R4192 GNDA.n275 GNDA.n273 3.5845
R4193 GNDA.n274 GNDA.n249 3.5845
R4194 GNDA.n282 GNDA.n281 3.5845
R4195 GNDA.n1059 GNDA.t75 3.42907
R4196 GNDA.n1059 GNDA.t50 3.42907
R4197 GNDA.n1144 GNDA.t92 3.42907
R4198 GNDA.n1144 GNDA.t73 3.42907
R4199 GNDA.n1142 GNDA.t179 3.42907
R4200 GNDA.n1142 GNDA.t199 3.42907
R4201 GNDA.n963 GNDA.t107 3.42907
R4202 GNDA.n963 GNDA.t342 3.42907
R4203 GNDA.n189 GNDA.n71 3.3797
R4204 GNDA.n96 GNDA.n40 3.3797
R4205 GNDA.n2130 GNDA.n413 3.3797
R4206 GNDA.n2129 GNDA.n2128 3.3797
R4207 GNDA.n2062 GNDA.n2061 3.3797
R4208 GNDA.n706 GNDA.n390 3.3797
R4209 GNDA.n2268 GNDA.n2156 3.3797
R4210 GNDA.n2256 GNDA.n2255 3.3797
R4211 GNDA.n1564 GNDA.n1342 3.3797
R4212 GNDA.n1513 GNDA.n1419 3.3797
R4213 GNDA.n1832 GNDA.n1233 3.3797
R4214 GNDA.n1831 GNDA.n1234 3.3797
R4215 GNDA.n1565 GNDA.n1311 3.3797
R4216 GNDA.n343 GNDA.n225 3.3797
R4217 GNDA.n250 GNDA.n52 3.3797
R4218 GNDA.n2129 GNDA.n414 3.27161
R4219 GNDA.n2393 GNDA.n71 3.27161
R4220 GNDA.n2156 GNDA.n380 3.27161
R4221 GNDA.n2352 GNDA.n225 3.27161
R4222 GNDA.n1876 GNDA.n1875 3.2005
R4223 GNDA.n1856 GNDA.n471 3.2005
R4224 GNDA.n1167 GNDA.t3 3.1344
R4225 GNDA.n1169 GNDA.t124 3.1344
R4226 GNDA.t118 GNDA.n1198 3.1344
R4227 GNDA.t337 GNDA.t288 3.1344
R4228 GNDA.n1187 GNDA.t55 3.1344
R4229 GNDA.n824 GNDA.t116 3.1344
R4230 GNDA.t129 GNDA.t229 3.1344
R4231 GNDA.n832 GNDA.t42 3.1344
R4232 GNDA.n322 GNDA 3.02272
R4233 GNDA.n1270 GNDA 3.02272
R4234 GNDA.n1754 GNDA 3.02272
R4235 GNDA.n2108 GNDA 3.02272
R4236 GNDA.n168 GNDA 3.02272
R4237 GNDA.n540 GNDA 3.02272
R4238 GNDA.n2214 GNDA 3.02272
R4239 GNDA.n752 GNDA 3.02272
R4240 GNDA.n1378 GNDA 3.02272
R4241 GNDA.n188 GNDA.n187 2.8677
R4242 GNDA.n638 GNDA.n510 2.8677
R4243 GNDA.n2015 GNDA.n416 2.8677
R4244 GNDA.n664 GNDA.n663 2.8677
R4245 GNDA.n2267 GNDA.n2266 2.8677
R4246 GNDA.n1524 GNDA.n1345 2.8677
R4247 GNDA.n1658 GNDA.n1654 2.8677
R4248 GNDA.n1576 GNDA.n1237 2.8677
R4249 GNDA.n342 GNDA.n341 2.8677
R4250 GNDA.n1147 GNDA.n887 2.5005
R4251 GNDA.n1933 GNDA.n472 2.4301
R4252 GNDA.n797 GNDA.n795 2.34425
R4253 GNDA.n805 GNDA.n803 2.34425
R4254 GNDA.n342 GNDA.n227 2.31161
R4255 GNDA.n1261 GNDA.n1237 2.31161
R4256 GNDA.n1762 GNDA.n1654 2.31161
R4257 GNDA.n2116 GNDA.n416 2.31161
R4258 GNDA.n188 GNDA.n73 2.31161
R4259 GNDA.n531 GNDA.n510 2.31161
R4260 GNDA.n2267 GNDA.n2157 2.31161
R4261 GNDA.n760 GNDA.n664 2.31161
R4262 GNDA.n1369 GNDA.n1345 2.31161
R4263 GNDA.n1146 GNDA.n1145 2.063
R4264 GNDA.n2351 GNDA.n2350 1.951
R4265 GNDA.n1580 GNDA.n1235 1.951
R4266 GNDA.n1885 GNDA.n494 1.951
R4267 GNDA.n1864 GNDA.n772 1.951
R4268 GNDA.n2008 GNDA.n373 1.951
R4269 GNDA.n2392 GNDA.n2391 1.951
R4270 GNDA.n389 GNDA.n374 1.951
R4271 GNDA.n1528 GNDA.n1343 1.951
R4272 GNDA.n1776 GNDA.n1619 1.951
R4273 GNDA.n1061 GNDA.n1060 1.813
R4274 GNDA.n1146 GNDA.n1141 1.78175
R4275 GNDA.n1062 GNDA.n1061 1.78175
R4276 GNDA.n189 GNDA.n188 1.7413
R4277 GNDA.n510 GNDA.n493 1.7413
R4278 GNDA.n2130 GNDA.n2129 1.7413
R4279 GNDA.n2128 GNDA.n416 1.7413
R4280 GNDA.n2061 GNDA.n71 1.7413
R4281 GNDA.n664 GNDA.n652 1.7413
R4282 GNDA.n2156 GNDA.n390 1.7413
R4283 GNDA.n2268 GNDA.n2267 1.7413
R4284 GNDA.n2255 GNDA.n225 1.7413
R4285 GNDA.n1345 GNDA.n1342 1.7413
R4286 GNDA.n1774 GNDA.n1654 1.7413
R4287 GNDA.n1832 GNDA.n1831 1.7413
R4288 GNDA.n1237 GNDA.n1234 1.7413
R4289 GNDA.n1565 GNDA.n1564 1.7413
R4290 GNDA.n343 GNDA.n342 1.7413
R4291 GNDA.n2516 GNDA.n2 1.73362
R4292 GNDA.n1131 GNDA.n1130 1.6005
R4293 GNDA.n2129 GNDA.n415 1.51754
R4294 GNDA.n2389 GNDA.n71 1.51754
R4295 GNDA.n2156 GNDA.n2155 1.51754
R4296 GNDA.n1831 GNDA.n1830 1.51754
R4297 GNDA.n1564 GNDA.n1563 1.51754
R4298 GNDA.n2348 GNDA.n225 1.51754
R4299 GNDA.n1907 GNDA 1.29343
R4300 GNDA.n1929 GNDA 1.29343
R4301 GNDA GNDA.n1624 1.29343
R4302 GNDA.n127 GNDA.n96 1.2293
R4303 GNDA.n631 GNDA.n413 1.2293
R4304 GNDA.n2065 GNDA.n2062 1.2293
R4305 GNDA.n709 GNDA.n706 1.2293
R4306 GNDA.n2259 GNDA.n2256 1.2293
R4307 GNDA.n1517 GNDA.n1419 1.2293
R4308 GNDA.n1711 GNDA.n1233 1.2293
R4309 GNDA.n1569 GNDA.n1311 1.2293
R4310 GNDA.n281 GNDA.n250 1.2293
R4311 GNDA.n1089 GNDA.n1088 1.21925
R4312 GNDA.n1887 GNDA.n1886 1.1781
R4313 GNDA.n1866 GNDA.n1865 1.1781
R4314 GNDA.n1775 GNDA.n1653 1.1781
R4315 GNDA.n2510 GNDA.n6 1.16414
R4316 GNDA.n187 GNDA.n74 1.0245
R4317 GNDA.n184 GNDA.n183 1.0245
R4318 GNDA.n104 GNDA.n76 1.0245
R4319 GNDA.n106 GNDA.n105 1.0245
R4320 GNDA.n113 GNDA.n102 1.0245
R4321 GNDA.n112 GNDA.n99 1.0245
R4322 GNDA.n119 GNDA.n98 1.0245
R4323 GNDA.n121 GNDA.n120 1.0245
R4324 GNDA.n128 GNDA.n95 1.0245
R4325 GNDA.n638 GNDA.n637 1.0245
R4326 GNDA.n594 GNDA.n511 1.0245
R4327 GNDA.n595 GNDA.n593 1.0245
R4328 GNDA.n609 GNDA.n608 1.0245
R4329 GNDA.n612 GNDA.n591 1.0245
R4330 GNDA.n614 GNDA.n613 1.0245
R4331 GNDA.n619 GNDA.n618 1.0245
R4332 GNDA.n615 GNDA.n583 1.0245
R4333 GNDA.n632 GNDA.n630 1.0245
R4334 GNDA.n2016 GNDA.n2015 1.0245
R4335 GNDA.n2122 GNDA.n2121 1.0245
R4336 GNDA.n2043 GNDA.n2017 1.0245
R4337 GNDA.n2046 GNDA.n2045 1.0245
R4338 GNDA.n2050 GNDA.n2049 1.0245
R4339 GNDA.n2054 GNDA.n2038 1.0245
R4340 GNDA.n2055 GNDA.n2037 1.0245
R4341 GNDA.n2059 GNDA.n2058 1.0245
R4342 GNDA.n2066 GNDA.n2060 1.0245
R4343 GNDA.n663 GNDA.n659 1.0245
R4344 GNDA.n766 GNDA.n765 1.0245
R4345 GNDA.n688 GNDA.n660 1.0245
R4346 GNDA.n691 GNDA.n690 1.0245
R4347 GNDA.n695 GNDA.n694 1.0245
R4348 GNDA.n699 GNDA.n683 1.0245
R4349 GNDA.n700 GNDA.n682 1.0245
R4350 GNDA.n704 GNDA.n703 1.0245
R4351 GNDA.n710 GNDA.n705 1.0245
R4352 GNDA.n2266 GNDA.n2265 1.0245
R4353 GNDA.n2185 GNDA.n2159 1.0245
R4354 GNDA.n2186 GNDA.n2184 1.0245
R4355 GNDA.n2192 GNDA.n2189 1.0245
R4356 GNDA.n2193 GNDA.n2182 1.0245
R4357 GNDA.n2199 GNDA.n2196 1.0245
R4358 GNDA.n2200 GNDA.n2181 1.0245
R4359 GNDA.n2204 GNDA.n2203 1.0245
R4360 GNDA.n2260 GNDA.n2205 1.0245
R4361 GNDA.n1524 GNDA.n1523 1.0245
R4362 GNDA.n1426 GNDA.n1346 1.0245
R4363 GNDA.n1429 GNDA.n1427 1.0245
R4364 GNDA.n1433 GNDA.n1432 1.0245
R4365 GNDA.n1423 GNDA.n1422 1.0245
R4366 GNDA.n1440 GNDA.n1439 1.0245
R4367 GNDA.n1443 GNDA.n1421 1.0245
R4368 GNDA.n1445 GNDA.n1444 1.0245
R4369 GNDA.n1518 GNDA.n1368 1.0245
R4370 GNDA.n1659 GNDA.n1658 1.0245
R4371 GNDA.n1768 GNDA.n1767 1.0245
R4372 GNDA.n1689 GNDA.n1660 1.0245
R4373 GNDA.n1690 GNDA.n1688 1.0245
R4374 GNDA.n1697 GNDA.n1695 1.0245
R4375 GNDA.n1696 GNDA.n1684 1.0245
R4376 GNDA.n1704 GNDA.n1703 1.0245
R4377 GNDA.n1685 GNDA.n1680 1.0245
R4378 GNDA.n1712 GNDA.n1710 1.0245
R4379 GNDA.n1576 GNDA.n1575 1.0245
R4380 GNDA.n1318 GNDA.n1238 1.0245
R4381 GNDA.n1321 GNDA.n1319 1.0245
R4382 GNDA.n1325 GNDA.n1324 1.0245
R4383 GNDA.n1315 GNDA.n1314 1.0245
R4384 GNDA.n1332 GNDA.n1331 1.0245
R4385 GNDA.n1335 GNDA.n1313 1.0245
R4386 GNDA.n1337 GNDA.n1336 1.0245
R4387 GNDA.n1570 GNDA.n1260 1.0245
R4388 GNDA.n341 GNDA.n228 1.0245
R4389 GNDA.n338 GNDA.n337 1.0245
R4390 GNDA.n258 GNDA.n230 1.0245
R4391 GNDA.n260 GNDA.n259 1.0245
R4392 GNDA.n267 GNDA.n256 1.0245
R4393 GNDA.n266 GNDA.n253 1.0245
R4394 GNDA.n273 GNDA.n252 1.0245
R4395 GNDA.n275 GNDA.n274 1.0245
R4396 GNDA.n282 GNDA.n249 1.0245
R4397 GNDA.n996 GNDA.t21 0.679512
R4398 GNDA.n1089 GNDA.n1064 0.6255
R4399 GNDA.n1019 GNDA.t19 0.578687
R4400 GNDA.n795 GNDA.n793 0.563
R4401 GNDA.n799 GNDA.n797 0.563
R4402 GNDA.n801 GNDA.n799 0.563
R4403 GNDA.n803 GNDA.n801 0.563
R4404 GNDA.n807 GNDA.n805 0.563
R4405 GNDA.n809 GNDA.n807 0.563
R4406 GNDA.n1121 GNDA.n1119 0.563
R4407 GNDA.n1123 GNDA.n1121 0.563
R4408 GNDA.n1125 GNDA.n1123 0.563
R4409 GNDA.n1127 GNDA.n1125 0.563
R4410 GNDA.n916 GNDA.n915 0.563
R4411 GNDA.n916 GNDA.n912 0.563
R4412 GNDA.n902 GNDA.n900 0.563
R4413 GNDA.n904 GNDA.n902 0.563
R4414 GNDA.n906 GNDA.n904 0.563
R4415 GNDA.n908 GNDA.n906 0.563
R4416 GNDA.n1066 GNDA.n889 0.563
R4417 GNDA.n1068 GNDA.n1066 0.563
R4418 GNDA.n1070 GNDA.n1068 0.563
R4419 GNDA.n1072 GNDA.n1070 0.563
R4420 GNDA.n1074 GNDA.n1072 0.563
R4421 GNDA.n1076 GNDA.n1074 0.563
R4422 GNDA.n1078 GNDA.n1076 0.563
R4423 GNDA.n1080 GNDA.n1078 0.563
R4424 GNDA.n1082 GNDA.n1080 0.563
R4425 GNDA.n1083 GNDA.n1082 0.563
R4426 GNDA.n1145 GNDA.n1143 0.5005
R4427 GNDA.n1060 GNDA.n1058 0.5005
R4428 GNDA GNDA.n437 0.474574
R4429 GNDA GNDA.n200 0.474574
R4430 GNDA GNDA.n400 0.474574
R4431 GNDA GNDA.n1593 0.474574
R4432 GNDA GNDA.n1539 0.474574
R4433 GNDA GNDA.n355 0.474574
R4434 GNDA.n790 GNDA.n788 0.41175
R4435 GNDA.n788 GNDA.n787 0.311875
R4436 GNDA.n1141 GNDA.n889 0.28175
R4437 GNDA.n812 GNDA.n811 0.276625
R4438 GNDA.n2517 GNDA.n1 0.276625
R4439 GNDA.n1115 GNDA.n918 0.2505
R4440 GNDA.n1088 GNDA.n1083 0.2505
R4441 GNDA.n1064 GNDA.n1062 0.2505
R4442 GNDA.n811 GNDA.n810 0.22375
R4443 GNDA.n810 GNDA.n1 0.100375
R4444 GNDA.n1984 GNDA.n452 0.0953148
R4445 GNDA.n2494 GNDA.n16 0.0953148
R4446 GNDA.n372 GNDA.n370 0.0953148
R4447 GNDA.n2298 GNDA.n2297 0.0953148
R4448 GNDA.n2353 GNDA.n220 0.0953148
R4449 GNDA.n2394 GNDA.n70 0.0953148
R4450 GNDA.n787 GNDA.n2 0.076875
R4451 a_14640_5738.t0 a_14640_5738.t1 169.905
R4452 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 345.264
R4453 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 344.7
R4454 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 344.7
R4455 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 206.052
R4456 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 205.488
R4457 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 205.488
R4458 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 205.488
R4459 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 205.488
R4460 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 122.474
R4461 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 57.7817
R4462 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 39.4005
R4463 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 39.4005
R4464 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 39.4005
R4465 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 39.4005
R4466 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 39.4005
R4467 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R4468 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R4469 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 19.7005
R4470 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 19.7005
R4471 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R4472 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 19.7005
R4473 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R4474 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 19.7005
R4475 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R4476 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R4477 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 19.7005
R4478 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 6.5005
R4479 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 6.1255
R4480 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R4481 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 0.563
R4482 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 0.563
R4483 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 0.563
R4484 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 325.473
R4485 bgr_0.V_mir2.n10 bgr_0.V_mir2.n6 325.471
R4486 bgr_0.V_mir2.n5 bgr_0.V_mir2.n1 325.471
R4487 bgr_0.V_mir2.n15 bgr_0.V_mir2.t20 310.488
R4488 bgr_0.V_mir2.n7 bgr_0.V_mir2.t22 310.488
R4489 bgr_0.V_mir2.n2 bgr_0.V_mir2.t18 310.488
R4490 bgr_0.V_mir2.n13 bgr_0.V_mir2.t1 278.312
R4491 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 228.939
R4492 bgr_0.V_mir2.n0 bgr_0.V_mir2.n11 224.439
R4493 bgr_0.V_mir2.n17 bgr_0.V_mir2.t8 184.097
R4494 bgr_0.V_mir2.n9 bgr_0.V_mir2.t14 184.097
R4495 bgr_0.V_mir2.n4 bgr_0.V_mir2.t6 184.097
R4496 bgr_0.V_mir2.n16 bgr_0.V_mir2.n15 167.094
R4497 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 167.094
R4498 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 167.094
R4499 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 152
R4500 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 152
R4501 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 152
R4502 bgr_0.V_mir2.n15 bgr_0.V_mir2.t19 120.501
R4503 bgr_0.V_mir2.n16 bgr_0.V_mir2.t4 120.501
R4504 bgr_0.V_mir2.n7 bgr_0.V_mir2.t21 120.501
R4505 bgr_0.V_mir2.n8 bgr_0.V_mir2.t10 120.501
R4506 bgr_0.V_mir2.n2 bgr_0.V_mir2.t17 120.501
R4507 bgr_0.V_mir2.n3 bgr_0.V_mir2.t12 120.501
R4508 bgr_0.V_mir2.n12 bgr_0.V_mir2.t2 48.0005
R4509 bgr_0.V_mir2.n12 bgr_0.V_mir2.t3 48.0005
R4510 bgr_0.V_mir2.n11 bgr_0.V_mir2.t0 48.0005
R4511 bgr_0.V_mir2.n11 bgr_0.V_mir2.t16 48.0005
R4512 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 40.7027
R4513 bgr_0.V_mir2.n9 bgr_0.V_mir2.n8 40.7027
R4514 bgr_0.V_mir2.n4 bgr_0.V_mir2.n3 40.7027
R4515 bgr_0.V_mir2.n6 bgr_0.V_mir2.t15 39.4005
R4516 bgr_0.V_mir2.n6 bgr_0.V_mir2.t11 39.4005
R4517 bgr_0.V_mir2.n1 bgr_0.V_mir2.t7 39.4005
R4518 bgr_0.V_mir2.n1 bgr_0.V_mir2.t13 39.4005
R4519 bgr_0.V_mir2.n19 bgr_0.V_mir2.t9 39.4005
R4520 bgr_0.V_mir2.t5 bgr_0.V_mir2.n19 39.4005
R4521 bgr_0.V_mir2.n14 bgr_0.V_mir2.n5 15.8005
R4522 bgr_0.V_mir2.n18 bgr_0.V_mir2.n14 15.8005
R4523 bgr_0.V_mir2.n0 bgr_0.V_mir2.n10 9.3005
R4524 bgr_0.V_mir2.n0 bgr_0.V_mir2.n13 5.8755
R4525 bgr_0.V_mir2.n14 bgr_0.V_mir2.n0 5.28175
R4526 bgr_0.1st_Vout_2 bgr_0.1st_Vout_2.t31 354.854
R4527 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t23 346.8
R4528 bgr_0.1st_Vout_2 bgr_0.1st_Vout_2.n11 339.522
R4529 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n4 339.522
R4530 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n6 335.022
R4531 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t10 275.909
R4532 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.n7 227.909
R4533 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n9 222.034
R4534 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t18 184.097
R4535 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t14 184.097
R4536 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t16 184.097
R4537 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t13 184.097
R4538 bgr_0.1st_Vout_2 bgr_0.1st_Vout_2.n10 166.05
R4539 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 166.05
R4540 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n2 57.7228
R4541 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t9 48.0005
R4542 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t7 48.0005
R4543 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t8 48.0005
R4544 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t6 48.0005
R4545 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t1 39.4005
R4546 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t3 39.4005
R4547 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t4 39.4005
R4548 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t5 39.4005
R4549 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t2 39.4005
R4550 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t0 39.4005
R4551 bgr_0.1st_Vout_2 bgr_0.1st_Vout_2.n0 5.6255
R4552 bgr_0.1st_Vout_2 bgr_0.1st_Vout_2.n3 5.28175
R4553 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t12 4.8295
R4554 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t29 4.8295
R4555 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t20 4.8295
R4556 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t35 4.8295
R4557 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.8295
R4558 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t28 4.8295
R4559 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.8295
R4560 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n8 4.5005
R4561 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t21 4.5005
R4562 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t27 4.5005
R4563 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t34 4.5005
R4564 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t26 4.5005
R4565 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t33 4.5005
R4566 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t15 4.5005
R4567 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.5005
R4568 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t25 4.5005
R4569 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t32 4.5005
R4570 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.5005
R4571 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t36 4.5005
R4572 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t17 4.5005
R4573 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t24 4.5005
R4574 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n1 3.8075
R4575 VDDA.n375 VDDA.n371 6600
R4576 VDDA.n375 VDDA.n372 6600
R4577 VDDA.n377 VDDA.n371 6570
R4578 VDDA.n377 VDDA.n372 6570
R4579 VDDA.n320 VDDA.n267 4710
R4580 VDDA.n320 VDDA.n268 4710
R4581 VDDA.n318 VDDA.n267 4710
R4582 VDDA.n318 VDDA.n268 4710
R4583 VDDA.n296 VDDA.n289 4710
R4584 VDDA.n298 VDDA.n289 4710
R4585 VDDA.n296 VDDA.n295 4710
R4586 VDDA.n298 VDDA.n295 4710
R4587 VDDA.n141 VDDA.n137 4605
R4588 VDDA.n141 VDDA.n138 4605
R4589 VDDA.n42 VDDA.n28 4605
R4590 VDDA.n44 VDDA.n28 4605
R4591 VDDA.n206 VDDA.n182 4590
R4592 VDDA.n208 VDDA.n182 4590
R4593 VDDA.n208 VDDA.n183 4590
R4594 VDDA.n206 VDDA.n183 4590
R4595 VDDA.n143 VDDA.n137 4575
R4596 VDDA.n143 VDDA.n138 4575
R4597 VDDA.n42 VDDA.n29 4575
R4598 VDDA.n44 VDDA.n29 4575
R4599 VDDA.n101 VDDA.n94 4020
R4600 VDDA.n103 VDDA.n94 4020
R4601 VDDA.n101 VDDA.n100 4020
R4602 VDDA.n103 VDDA.n100 4020
R4603 VDDA.n77 VDDA.n70 4020
R4604 VDDA.n79 VDDA.n70 4020
R4605 VDDA.n77 VDDA.n76 4020
R4606 VDDA.n79 VDDA.n76 4020
R4607 VDDA.n442 VDDA.n437 3420
R4608 VDDA.n440 VDDA.n437 3420
R4609 VDDA.n121 VDDA.n114 3390
R4610 VDDA.n123 VDDA.n114 3390
R4611 VDDA.n121 VDDA.n120 3390
R4612 VDDA.n123 VDDA.n120 3390
R4613 VDDA.n21 VDDA.n14 3390
R4614 VDDA.n23 VDDA.n14 3390
R4615 VDDA.n21 VDDA.n20 3390
R4616 VDDA.n23 VDDA.n20 3390
R4617 VDDA.n163 VDDA.n157 2940
R4618 VDDA.n165 VDDA.n157 2940
R4619 VDDA.n165 VDDA.n162 2940
R4620 VDDA.n163 VDDA.n162 2940
R4621 VDDA.n171 VDDA.n152 2940
R4622 VDDA.n173 VDDA.n152 2940
R4623 VDDA.n173 VDDA.n170 2940
R4624 VDDA.n171 VDDA.n170 2940
R4625 VDDA.n442 VDDA.n436 2760
R4626 VDDA.n440 VDDA.n436 2760
R4627 VDDA.n235 VDDA.n224 2415
R4628 VDDA.n235 VDDA.n225 2370
R4629 VDDA.n232 VDDA.n225 2280
R4630 VDDA.n232 VDDA.n224 2235
R4631 VDDA.n454 VDDA.n450 2145
R4632 VDDA.n457 VDDA.n450 2100
R4633 VDDA.n457 VDDA.n451 2100
R4634 VDDA.n428 VDDA.n422 2100
R4635 VDDA.n428 VDDA.n423 2100
R4636 VDDA.n426 VDDA.n422 2100
R4637 VDDA.n426 VDDA.n423 2100
R4638 VDDA.n454 VDDA.n451 2055
R4639 VDDA.n389 VDDA.n384 1770
R4640 VDDA.n391 VDDA.n384 1770
R4641 VDDA.n389 VDDA.n387 1770
R4642 VDDA.n391 VDDA.n387 1770
R4643 VDDA.n362 VDDA.n357 1770
R4644 VDDA.n364 VDDA.n357 1770
R4645 VDDA.n362 VDDA.n360 1770
R4646 VDDA.n364 VDDA.n360 1770
R4647 VDDA.n247 VDDA.n220 1575
R4648 VDDA.n246 VDDA.n220 1575
R4649 VDDA.n246 VDDA.n219 1545
R4650 VDDA.n247 VDDA.n219 1545
R4651 VDDA.n135 VDDA.t58 1216.42
R4652 VDDA.n146 VDDA.t43 1216.42
R4653 VDDA.n39 VDDA.t61 1216.42
R4654 VDDA.n47 VDDA.t89 1216.42
R4655 VDDA.n374 VDDA.n373 704
R4656 VDDA.n374 VDDA.n340 704
R4657 VDDA.n159 VDDA.t39 689.4
R4658 VDDA.n158 VDDA.t54 689.4
R4659 VDDA.n154 VDDA.t121 689.4
R4660 VDDA.n153 VDDA.t21 689.4
R4661 VDDA.n202 VDDA.t112 663.801
R4662 VDDA.n212 VDDA.t106 663.801
R4663 VDDA.n97 VDDA.t113 660.109
R4664 VDDA.n95 VDDA.t22 660.109
R4665 VDDA.n73 VDDA.t7 660.109
R4666 VDDA.n71 VDDA.t95 660.109
R4667 VDDA.n242 VDDA.t51 647.54
R4668 VDDA.n251 VDDA.t88 647.54
R4669 VDDA.n216 VDDA.n215 633.361
R4670 VDDA.n179 VDDA.n178 626.534
R4671 VDDA.n185 VDDA.n184 626.534
R4672 VDDA.n187 VDDA.n186 626.534
R4673 VDDA.n189 VDDA.n188 626.534
R4674 VDDA.n191 VDDA.n190 626.534
R4675 VDDA.n193 VDDA.n192 626.534
R4676 VDDA.n195 VDDA.n194 626.534
R4677 VDDA.n197 VDDA.n196 626.534
R4678 VDDA.n199 VDDA.n198 626.534
R4679 VDDA.n201 VDDA.n200 626.534
R4680 VDDA.n229 VDDA.t16 623.958
R4681 VDDA.n238 VDDA.t31 623.958
R4682 VDDA.t16 VDDA.n228 615.926
R4683 VDDA.n117 VDDA.t46 573.75
R4684 VDDA.n115 VDDA.t73 573.75
R4685 VDDA.n17 VDDA.t70 573.75
R4686 VDDA.n15 VDDA.t92 573.75
R4687 VDDA.n379 VDDA.n378 518.4
R4688 VDDA.n378 VDDA.n370 518.4
R4689 VDDA.n300 VDDA.n299 496
R4690 VDDA.n300 VDDA.n288 496
R4691 VDDA.n140 VDDA.n112 491.2
R4692 VDDA.n140 VDDA.n139 491.2
R4693 VDDA.n45 VDDA.n27 491.2
R4694 VDDA.n41 VDDA.n27 491.2
R4695 VDDA.n205 VDDA.n181 489.601
R4696 VDDA.n209 VDDA.n181 489.601
R4697 VDDA.n105 VDDA.n104 428.8
R4698 VDDA.n105 VDDA.n93 428.8
R4699 VDDA.n81 VDDA.n80 428.8
R4700 VDDA.n81 VDDA.n69 428.8
R4701 VDDA.n382 VDDA.t98 419.108
R4702 VDDA.n385 VDDA.t28 419.108
R4703 VDDA.n355 VDDA.t10 413.084
R4704 VDDA.n358 VDDA.t40 413.084
R4705 VDDA.n448 VDDA.t116 409.067
R4706 VDDA.n460 VDDA.t25 409.067
R4707 VDDA.n434 VDDA.t13 409.067
R4708 VDDA.n445 VDDA.t76 409.067
R4709 VDDA.n420 VDDA.t34 409.067
R4710 VDDA.n431 VDDA.t101 390.322
R4711 VDDA.t111 VDDA.n206 389.375
R4712 VDDA.n208 VDDA.t105 389.375
R4713 VDDA.t120 VDDA.n170 389.375
R4714 VDDA.t20 VDDA.n152 389.375
R4715 VDDA.n382 VDDA.t100 389.185
R4716 VDDA.n385 VDDA.t30 389.185
R4717 VDDA.n204 VDDA.n180 387.2
R4718 VDDA.n210 VDDA.n180 387.2
R4719 VDDA.n445 VDDA.t78 387.051
R4720 VDDA.n434 VDDA.t15 387.051
R4721 VDDA.n355 VDDA.t12 384.918
R4722 VDDA.n358 VDDA.t42 384.918
R4723 VDDA.n269 VDDA.t66 384.918
R4724 VDDA.n271 VDDA.t109 384.918
R4725 VDDA.n292 VDDA.t69 384.918
R4726 VDDA.n290 VDDA.t57 384.918
R4727 VDDA.t38 VDDA.n162 384.168
R4728 VDDA.t53 VDDA.n157 384.168
R4729 VDDA.n317 VDDA.n270 384
R4730 VDDA.n317 VDDA.n316 384
R4731 VDDA.n294 VDDA.n293 384
R4732 VDDA.n294 VDDA.n291 384
R4733 VDDA.n431 VDDA.t103 370.728
R4734 VDDA.n420 VDDA.t36 370.728
R4735 VDDA.n460 VDDA.t27 370.3
R4736 VDDA.n448 VDDA.t118 370.3
R4737 VDDA.n439 VDDA.n438 364.8
R4738 VDDA.n369 VDDA.t79 360.868
R4739 VDDA.n380 VDDA.t82 360.868
R4740 VDDA.n269 VDDA.t64 358.858
R4741 VDDA.n271 VDDA.t107 358.858
R4742 VDDA.n292 VDDA.t67 358.858
R4743 VDDA.n290 VDDA.t55 358.858
R4744 VDDA.n125 VDDA.n124 355.2
R4745 VDDA.n125 VDDA.n113 355.2
R4746 VDDA.n25 VDDA.n24 355.2
R4747 VDDA.n25 VDDA.n13 355.2
R4748 VDDA.t65 VDDA.n267 351.591
R4749 VDDA.t108 VDDA.n268 351.591
R4750 VDDA.t68 VDDA.n296 351.591
R4751 VDDA.n298 VDDA.t56 351.591
R4752 VDDA.t50 VDDA.n246 346.668
R4753 VDDA.n247 VDDA.t86 346.668
R4754 VDDA.n416 VDDA.n415 345.127
R4755 VDDA.n419 VDDA.n418 345.127
R4756 VDDA.n400 VDDA.n399 344.7
R4757 VDDA.n403 VDDA.n402 344.7
R4758 VDDA.t26 VDDA.n450 344.394
R4759 VDDA.t117 VDDA.n451 344.394
R4760 VDDA.t99 VDDA.n389 344.394
R4761 VDDA.n391 VDDA.t29 344.394
R4762 VDDA.t11 VDDA.n362 344.394
R4763 VDDA.n364 VDDA.t41 344.394
R4764 VDDA.n283 VDDA.n281 342.301
R4765 VDDA.n311 VDDA.n310 341.676
R4766 VDDA.n309 VDDA.n308 341.676
R4767 VDDA.n307 VDDA.n306 341.676
R4768 VDDA.n305 VDDA.n304 341.676
R4769 VDDA.n287 VDDA.n286 341.676
R4770 VDDA.n285 VDDA.n284 341.676
R4771 VDDA.n283 VDDA.n282 341.676
R4772 VDDA.t77 VDDA.n436 340.635
R4773 VDDA.t14 VDDA.n437 340.635
R4774 VDDA.t102 VDDA.n422 340.635
R4775 VDDA.t35 VDDA.n423 340.635
R4776 VDDA.n405 VDDA.n404 339.272
R4777 VDDA.n408 VDDA.n407 339.272
R4778 VDDA.n410 VDDA.n409 339.272
R4779 VDDA.n412 VDDA.n411 339.272
R4780 VDDA.n414 VDDA.n413 339.272
R4781 VDDA.n279 VDDA.n278 337.176
R4782 VDDA.n276 VDDA.n274 337.176
R4783 VDDA.n265 VDDA.n264 337.176
R4784 VDDA.n322 VDDA.n263 337.176
R4785 VDDA.n325 VDDA.n324 337.176
R4786 VDDA.n329 VDDA.n328 337.176
R4787 VDDA.n332 VDDA.n331 337.176
R4788 VDDA.n335 VDDA.n259 337.176
R4789 VDDA.n313 VDDA.n273 337.176
R4790 VDDA.n302 VDDA.n301 337.176
R4791 VDDA.n396 VDDA.n395 335.022
R4792 VDDA.n203 VDDA.t110 332.75
R4793 VDDA.n211 VDDA.t104 332.75
R4794 VDDA.n159 VDDA.t37 332.75
R4795 VDDA.n158 VDDA.t52 332.75
R4796 VDDA.n154 VDDA.t119 332.75
R4797 VDDA.n153 VDDA.t19 332.75
R4798 VDDA.n243 VDDA.t49 314.274
R4799 VDDA.n250 VDDA.t85 314.274
R4800 VDDA.n161 VDDA.n156 313.601
R4801 VDDA.n168 VDDA.n156 307.2
R4802 VDDA.n176 VDDA.n151 307.2
R4803 VDDA.n169 VDDA.n151 307.2
R4804 VDDA.n439 VDDA.n406 294.401
R4805 VDDA.t47 VDDA.n121 285.815
R4806 VDDA.n123 VDDA.t74 285.815
R4807 VDDA.t71 VDDA.n21 285.815
R4808 VDDA.n23 VDDA.t93 285.815
R4809 VDDA.t83 VDDA.n371 278.95
R4810 VDDA.t80 VDDA.n372 278.95
R4811 VDDA.n117 VDDA.t48 277.916
R4812 VDDA.n115 VDDA.t75 277.916
R4813 VDDA.n17 VDDA.t72 277.916
R4814 VDDA.n15 VDDA.t94 277.916
R4815 VDDA.n145 VDDA.n112 276.8
R4816 VDDA.n139 VDDA.n136 276.8
R4817 VDDA.n46 VDDA.n45 276.8
R4818 VDDA.n41 VDDA.n40 276.8
R4819 VDDA.n380 VDDA.t84 270.705
R4820 VDDA.n369 VDDA.t81 270.705
R4821 VDDA.n236 VDDA.n223 257.601
R4822 VDDA.n443 VDDA.n435 246.4
R4823 VDDA.t114 VDDA.n101 239.915
R4824 VDDA.n103 VDDA.t23 239.915
R4825 VDDA.t8 VDDA.n77 239.915
R4826 VDDA.n79 VDDA.t96 239.915
R4827 VDDA.n231 VDDA.n223 238.4
R4828 VDDA.n99 VDDA.n98 230.4
R4829 VDDA.n99 VDDA.n96 230.4
R4830 VDDA.n75 VDDA.n74 230.4
R4831 VDDA.n75 VDDA.n72 230.4
R4832 VDDA.n453 VDDA.n401 228.8
R4833 VDDA.n425 VDDA.n424 224
R4834 VDDA.n425 VDDA.n417 224
R4835 VDDA.n453 VDDA.n452 219.201
R4836 VDDA.n166 VDDA.n160 211.201
R4837 VDDA.n167 VDDA.n166 211.201
R4838 VDDA.n175 VDDA.n174 211.201
R4839 VDDA.n119 VDDA.n118 211.201
R4840 VDDA.n119 VDDA.n116 211.201
R4841 VDDA.n19 VDDA.n18 211.201
R4842 VDDA.n19 VDDA.n16 211.201
R4843 VDDA.n145 VDDA.n144 204.8
R4844 VDDA.n144 VDDA.n136 204.8
R4845 VDDA.n40 VDDA.n26 204.8
R4846 VDDA.n46 VDDA.n26 204.8
R4847 VDDA.n174 VDDA.n155 202.971
R4848 VDDA.n104 VDDA.n96 198.4
R4849 VDDA.n98 VDDA.n93 198.4
R4850 VDDA.n80 VDDA.n72 198.4
R4851 VDDA.n74 VDDA.n69 198.4
R4852 VDDA.n231 VDDA.n230 192
R4853 VDDA.t375 VDDA.t50 190
R4854 VDDA.t86 VDDA.t375 190
R4855 VDDA.n237 VDDA.n236 188.8
R4856 VDDA.n392 VDDA.n386 188.8
R4857 VDDA.n388 VDDA.n386 188.8
R4858 VDDA.n365 VDDA.n359 188.8
R4859 VDDA.n361 VDDA.n359 188.8
R4860 VDDA.n315 VDDA.n314 188.8
R4861 VDDA.n334 VDDA.n260 188.8
R4862 VDDA.t331 VDDA.t111 186.607
R4863 VDDA.t186 VDDA.t331 186.607
R4864 VDDA.t180 VDDA.t186 186.607
R4865 VDDA.t148 VDDA.t180 186.607
R4866 VDDA.t178 VDDA.t148 186.607
R4867 VDDA.t134 VDDA.t178 186.607
R4868 VDDA.t327 VDDA.t134 186.607
R4869 VDDA.t218 VDDA.t327 186.607
R4870 VDDA.t140 VDDA.t218 186.607
R4871 VDDA.t329 VDDA.t140 186.607
R4872 VDDA.t220 VDDA.t146 186.607
R4873 VDDA.t356 VDDA.t220 186.607
R4874 VDDA.t176 VDDA.t356 186.607
R4875 VDDA.t188 VDDA.t176 186.607
R4876 VDDA.t325 VDDA.t188 186.607
R4877 VDDA.t136 VDDA.t325 186.607
R4878 VDDA.t138 VDDA.t136 186.607
R4879 VDDA.t182 VDDA.t138 186.607
R4880 VDDA.t358 VDDA.t182 186.607
R4881 VDDA.t105 VDDA.t358 186.607
R4882 VDDA.t124 VDDA.t120 186.607
R4883 VDDA.t273 VDDA.t124 186.607
R4884 VDDA.t466 VDDA.t273 186.607
R4885 VDDA.t201 VDDA.t466 186.607
R4886 VDDA.t290 VDDA.t201 186.607
R4887 VDDA.t215 VDDA.t322 186.607
R4888 VDDA.t322 VDDA.t204 186.607
R4889 VDDA.t204 VDDA.t125 186.607
R4890 VDDA.t125 VDDA.t368 186.607
R4891 VDDA.t368 VDDA.t20 186.607
R4892 VDDA.t203 VDDA.t38 183.333
R4893 VDDA.t403 VDDA.t203 183.333
R4894 VDDA.t350 VDDA.t403 183.333
R4895 VDDA.t267 VDDA.t350 183.333
R4896 VDDA.t289 VDDA.t267 183.333
R4897 VDDA.t154 VDDA.t235 183.333
R4898 VDDA.t235 VDDA.t268 183.333
R4899 VDDA.t268 VDDA.t202 183.333
R4900 VDDA.t202 VDDA.t266 183.333
R4901 VDDA.t266 VDDA.t53 183.333
R4902 VDDA.n373 VDDA.n370 182.4
R4903 VDDA.n379 VDDA.n340 182.4
R4904 VDDA.n134 VDDA.t60 178.124
R4905 VDDA.n147 VDDA.t45 178.124
R4906 VDDA.n38 VDDA.t63 178.124
R4907 VDDA.n48 VDDA.t91 178.124
R4908 VDDA.n444 VDDA.n443 176
R4909 VDDA.n226 VDDA.n221 174.393
R4910 VDDA.t419 VDDA.t65 172.727
R4911 VDDA.t242 VDDA.t419 172.727
R4912 VDDA.t238 VDDA.t242 172.727
R4913 VDDA.t258 VDDA.t238 172.727
R4914 VDDA.t256 VDDA.t258 172.727
R4915 VDDA.t427 VDDA.t256 172.727
R4916 VDDA.t423 VDDA.t427 172.727
R4917 VDDA.t254 VDDA.t423 172.727
R4918 VDDA.t248 VDDA.t254 172.727
R4919 VDDA.t240 VDDA.t236 172.727
R4920 VDDA.t236 VDDA.t425 172.727
R4921 VDDA.t425 VDDA.t421 172.727
R4922 VDDA.t421 VDDA.t252 172.727
R4923 VDDA.t252 VDDA.t246 172.727
R4924 VDDA.t246 VDDA.t250 172.727
R4925 VDDA.t250 VDDA.t244 172.727
R4926 VDDA.t244 VDDA.t417 172.727
R4927 VDDA.t417 VDDA.t108 172.727
R4928 VDDA.t303 VDDA.t68 172.727
R4929 VDDA.t436 VDDA.t303 172.727
R4930 VDDA.t285 VDDA.t436 172.727
R4931 VDDA.t222 VDDA.t285 172.727
R4932 VDDA.t291 VDDA.t222 172.727
R4933 VDDA.t3 VDDA.t291 172.727
R4934 VDDA.t209 VDDA.t3 172.727
R4935 VDDA.t434 VDDA.t209 172.727
R4936 VDDA.t211 VDDA.t434 172.727
R4937 VDDA.t431 VDDA.t467 172.727
R4938 VDDA.t5 VDDA.t431 172.727
R4939 VDDA.t280 VDDA.t5 172.727
R4940 VDDA.t287 VDDA.t280 172.727
R4941 VDDA.t213 VDDA.t287 172.727
R4942 VDDA.t168 VDDA.t213 172.727
R4943 VDDA.t387 VDDA.t168 172.727
R4944 VDDA.t271 VDDA.t387 172.727
R4945 VDDA.t56 VDDA.t271 172.727
R4946 VDDA.t17 VDDA.n232 172.554
R4947 VDDA.n235 VDDA.t32 172.554
R4948 VDDA.n339 VDDA.n338 168.435
R4949 VDDA.n342 VDDA.n341 168.435
R4950 VDDA.n344 VDDA.n343 168.435
R4951 VDDA.n346 VDDA.n345 168.435
R4952 VDDA.n348 VDDA.n347 168.435
R4953 VDDA.n350 VDDA.n349 168.435
R4954 VDDA.n352 VDDA.n351 168.435
R4955 VDDA.n354 VDDA.n353 168.435
R4956 VDDA.n245 VDDA.n218 164.8
R4957 VDDA.n248 VDDA.n218 164.8
R4958 VDDA.t44 VDDA.n137 161.817
R4959 VDDA.t59 VDDA.n138 161.817
R4960 VDDA.t62 VDDA.n42 161.817
R4961 VDDA.n44 VDDA.t90 161.817
R4962 VDDA.n91 VDDA.n89 160.428
R4963 VDDA.n88 VDDA.n86 160.428
R4964 VDDA.n67 VDDA.n65 160.428
R4965 VDDA.n64 VDDA.n62 160.428
R4966 VDDA.t345 VDDA.t83 159.814
R4967 VDDA.t453 VDDA.t345 159.814
R4968 VDDA.t165 VDDA.t453 159.814
R4969 VDDA.t348 VDDA.t165 159.814
R4970 VDDA.t362 VDDA.t348 159.814
R4971 VDDA.t459 VDDA.t362 159.814
R4972 VDDA.t299 VDDA.t459 159.814
R4973 VDDA.t341 VDDA.t299 159.814
R4974 VDDA.t159 VDDA.t0 159.814
R4975 VDDA.t0 VDDA.t228 159.814
R4976 VDDA.t228 VDDA.t163 159.814
R4977 VDDA.t163 VDDA.t161 159.814
R4978 VDDA.t161 VDDA.t442 159.814
R4979 VDDA.t442 VDDA.t383 159.814
R4980 VDDA.t383 VDDA.t455 159.814
R4981 VDDA.t455 VDDA.t80 159.814
R4982 VDDA.n91 VDDA.n90 159.803
R4983 VDDA.n88 VDDA.n87 159.803
R4984 VDDA.n67 VDDA.n66 159.803
R4985 VDDA.n64 VDDA.n63 159.803
R4986 VDDA.t369 VDDA.t26 158.333
R4987 VDDA.t351 VDDA.t369 158.333
R4988 VDDA.t122 VDDA.t449 158.333
R4989 VDDA.t449 VDDA.t117 158.333
R4990 VDDA.t155 VDDA.t99 158.333
R4991 VDDA.t29 VDDA.t379 158.333
R4992 VDDA.t464 VDDA.t11 158.333
R4993 VDDA.t41 VDDA.t465 158.333
R4994 VDDA.t132 VDDA.t77 155.97
R4995 VDDA.t371 VDDA.t132 155.97
R4996 VDDA.t170 VDDA.t371 155.97
R4997 VDDA.t130 VDDA.t170 155.97
R4998 VDDA.t283 VDDA.t152 155.97
R4999 VDDA.t152 VDDA.t192 155.97
R5000 VDDA.t192 VDDA.t413 155.97
R5001 VDDA.t413 VDDA.t373 155.97
R5002 VDDA.t373 VDDA.t190 155.97
R5003 VDDA.t190 VDDA.t14 155.97
R5004 VDDA.t389 VDDA.t102 155.97
R5005 VDDA.t438 VDDA.t389 155.97
R5006 VDDA.t274 VDDA.t440 155.97
R5007 VDDA.t440 VDDA.t35 155.97
R5008 VDDA.n97 VDDA.t115 155.125
R5009 VDDA.n95 VDDA.t24 155.125
R5010 VDDA.n73 VDDA.t9 155.125
R5011 VDDA.n71 VDDA.t97 155.125
R5012 VDDA.n134 VDDA.n133 151.882
R5013 VDDA.n38 VDDA.n37 151.882
R5014 VDDA.n148 VDDA.n147 151.321
R5015 VDDA.n49 VDDA.n48 151.321
R5016 VDDA.n124 VDDA.n116 150.4
R5017 VDDA.n118 VDDA.n113 150.4
R5018 VDDA.n24 VDDA.n16 150.4
R5019 VDDA.n18 VDDA.n13 150.4
R5020 VDDA.n107 VDDA.n106 146.002
R5021 VDDA.n83 VDDA.n82 146.002
R5022 VDDA.n111 VDDA.n110 145.429
R5023 VDDA.n127 VDDA.n126 145.429
R5024 VDDA.n129 VDDA.n128 145.429
R5025 VDDA.n131 VDDA.n130 145.429
R5026 VDDA.n133 VDDA.n132 145.429
R5027 VDDA.n12 VDDA.n11 145.429
R5028 VDDA.n31 VDDA.n30 145.429
R5029 VDDA.n33 VDDA.n32 145.429
R5030 VDDA.n35 VDDA.n34 145.429
R5031 VDDA.n37 VDDA.n36 145.429
R5032 VDDA.n147 VDDA.n146 135.387
R5033 VDDA.n135 VDDA.n134 135.387
R5034 VDDA.n48 VDDA.n47 135.387
R5035 VDDA.n39 VDDA.n38 135.387
R5036 VDDA.t321 VDDA.t47 121.513
R5037 VDDA.t398 VDDA.t321 121.513
R5038 VDDA.t264 VDDA.t398 121.513
R5039 VDDA.t404 VDDA.t264 121.513
R5040 VDDA.t227 VDDA.t404 121.513
R5041 VDDA.t150 VDDA.t224 121.513
R5042 VDDA.t305 VDDA.t150 121.513
R5043 VDDA.t320 VDDA.t305 121.513
R5044 VDDA.t391 VDDA.t320 121.513
R5045 VDDA.t74 VDDA.t391 121.513
R5046 VDDA.t353 VDDA.t71 121.513
R5047 VDDA.t457 VDDA.t353 121.513
R5048 VDDA.t157 VDDA.t457 121.513
R5049 VDDA.t433 VDDA.t157 121.513
R5050 VDDA.t158 VDDA.t433 121.513
R5051 VDDA.t463 VDDA.t314 121.513
R5052 VDDA.t343 VDDA.t463 121.513
R5053 VDDA.t367 VDDA.t343 121.513
R5054 VDDA.t451 VDDA.t367 121.513
R5055 VDDA.t93 VDDA.t451 121.513
R5056 VDDA.n452 VDDA.n449 118.4
R5057 VDDA.n459 VDDA.n401 118.4
R5058 VDDA.n438 VDDA.n435 118.4
R5059 VDDA.n444 VDDA.n406 118.4
R5060 VDDA.n424 VDDA.n421 118.4
R5061 VDDA.n430 VDDA.n417 118.4
R5062 VDDA.n393 VDDA.n392 118.4
R5063 VDDA.n388 VDDA.n383 118.4
R5064 VDDA.n366 VDDA.n365 118.4
R5065 VDDA.n361 VDDA.n356 118.4
R5066 VDDA.n316 VDDA.n315 118.4
R5067 VDDA.n270 VDDA.n260 118.4
R5068 VDDA.n299 VDDA.n291 118.4
R5069 VDDA.n293 VDDA.n288 118.4
R5070 VDDA.n245 VDDA.n244 110.4
R5071 VDDA.n249 VDDA.n248 110.4
R5072 VDDA.n459 VDDA.n458 105.6
R5073 VDDA.n458 VDDA.n449 105.6
R5074 VDDA.n430 VDDA.n429 105.6
R5075 VDDA.n429 VDDA.n421 105.6
R5076 VDDA.t32 VDDA.t172 102.704
R5077 VDDA.n205 VDDA.n204 102.4
R5078 VDDA.n210 VDDA.n209 102.4
R5079 VDDA.n161 VDDA.n160 102.4
R5080 VDDA.n240 VDDA.n239 101.267
R5081 VDDA.t415 VDDA.t114 98.2764
R5082 VDDA.t144 VDDA.t415 98.2764
R5083 VDDA.t126 VDDA.t144 98.2764
R5084 VDDA.t297 VDDA.t126 98.2764
R5085 VDDA.t429 VDDA.t297 98.2764
R5086 VDDA.t399 VDDA.t184 98.2764
R5087 VDDA.t216 VDDA.t399 98.2764
R5088 VDDA.t196 VDDA.t216 98.2764
R5089 VDDA.t174 VDDA.t196 98.2764
R5090 VDDA.t23 VDDA.t174 98.2764
R5091 VDDA.t401 VDDA.t8 98.2764
R5092 VDDA.t335 VDDA.t401 98.2764
R5093 VDDA.t377 VDDA.t335 98.2764
R5094 VDDA.t233 VDDA.t377 98.2764
R5095 VDDA.t333 VDDA.t233 98.2764
R5096 VDDA.t407 VDDA.t194 98.2764
R5097 VDDA.t142 VDDA.t407 98.2764
R5098 VDDA.t337 VDDA.t142 98.2764
R5099 VDDA.t354 VDDA.t337 98.2764
R5100 VDDA.t96 VDDA.t354 98.2764
R5101 VDDA.n52 VDDA.n50 97.4034
R5102 VDDA.n2 VDDA.n0 97.4034
R5103 VDDA.n60 VDDA.n59 96.8409
R5104 VDDA.n58 VDDA.n57 96.8409
R5105 VDDA.n56 VDDA.n55 96.8409
R5106 VDDA.n54 VDDA.n53 96.8409
R5107 VDDA.n52 VDDA.n51 96.8409
R5108 VDDA.n10 VDDA.n9 96.8409
R5109 VDDA.n8 VDDA.n7 96.8409
R5110 VDDA.n6 VDDA.n5 96.8409
R5111 VDDA.n4 VDDA.n3 96.8409
R5112 VDDA.n2 VDDA.n1 96.8409
R5113 VDDA.n168 VDDA.n167 96.0005
R5114 VDDA.n169 VDDA.n155 96.0005
R5115 VDDA.n176 VDDA.n175 96.0005
R5116 VDDA.n207 VDDA.t329 93.3041
R5117 VDDA.t146 VDDA.n207 93.3041
R5118 VDDA.n172 VDDA.t290 93.3041
R5119 VDDA.n172 VDDA.t215 93.3041
R5120 VDDA.n219 VDDA.n218 92.5005
R5121 VDDA.t375 VDDA.n219 92.5005
R5122 VDDA.n220 VDDA.n217 92.5005
R5123 VDDA.t375 VDDA.n220 92.5005
R5124 VDDA.n224 VDDA.n223 92.5005
R5125 VDDA.n233 VDDA.n224 92.5005
R5126 VDDA.n225 VDDA.n222 92.5005
R5127 VDDA.n234 VDDA.n225 92.5005
R5128 VDDA.n206 VDDA.n205 92.5005
R5129 VDDA.n182 VDDA.n181 92.5005
R5130 VDDA.n207 VDDA.n182 92.5005
R5131 VDDA.n209 VDDA.n208 92.5005
R5132 VDDA.n183 VDDA.n180 92.5005
R5133 VDDA.n207 VDDA.n183 92.5005
R5134 VDDA.n163 VDDA.n156 92.5005
R5135 VDDA.n164 VDDA.n163 92.5005
R5136 VDDA.n162 VDDA.n161 92.5005
R5137 VDDA.n166 VDDA.n165 92.5005
R5138 VDDA.n165 VDDA.n164 92.5005
R5139 VDDA.n168 VDDA.n157 92.5005
R5140 VDDA.n171 VDDA.n151 92.5005
R5141 VDDA.n172 VDDA.n171 92.5005
R5142 VDDA.n170 VDDA.n169 92.5005
R5143 VDDA.n174 VDDA.n173 92.5005
R5144 VDDA.n173 VDDA.n172 92.5005
R5145 VDDA.n176 VDDA.n152 92.5005
R5146 VDDA.n124 VDDA.n123 92.5005
R5147 VDDA.n120 VDDA.n119 92.5005
R5148 VDDA.n122 VDDA.n120 92.5005
R5149 VDDA.n121 VDDA.n113 92.5005
R5150 VDDA.n125 VDDA.n114 92.5005
R5151 VDDA.n122 VDDA.n114 92.5005
R5152 VDDA.n144 VDDA.n143 92.5005
R5153 VDDA.n143 VDDA.n142 92.5005
R5154 VDDA.n141 VDDA.n140 92.5005
R5155 VDDA.n142 VDDA.n141 92.5005
R5156 VDDA.n104 VDDA.n103 92.5005
R5157 VDDA.n100 VDDA.n99 92.5005
R5158 VDDA.n102 VDDA.n100 92.5005
R5159 VDDA.n101 VDDA.n93 92.5005
R5160 VDDA.n105 VDDA.n94 92.5005
R5161 VDDA.n102 VDDA.n94 92.5005
R5162 VDDA.n80 VDDA.n79 92.5005
R5163 VDDA.n76 VDDA.n75 92.5005
R5164 VDDA.n78 VDDA.n76 92.5005
R5165 VDDA.n77 VDDA.n69 92.5005
R5166 VDDA.n81 VDDA.n70 92.5005
R5167 VDDA.n78 VDDA.n70 92.5005
R5168 VDDA.n24 VDDA.n23 92.5005
R5169 VDDA.n20 VDDA.n19 92.5005
R5170 VDDA.n22 VDDA.n20 92.5005
R5171 VDDA.n21 VDDA.n13 92.5005
R5172 VDDA.n25 VDDA.n14 92.5005
R5173 VDDA.n22 VDDA.n14 92.5005
R5174 VDDA.n29 VDDA.n26 92.5005
R5175 VDDA.n43 VDDA.n29 92.5005
R5176 VDDA.n28 VDDA.n27 92.5005
R5177 VDDA.n43 VDDA.n28 92.5005
R5178 VDDA.n452 VDDA.n451 92.5005
R5179 VDDA.n454 VDDA.n453 92.5005
R5180 VDDA.n455 VDDA.n454 92.5005
R5181 VDDA.n450 VDDA.n401 92.5005
R5182 VDDA.n458 VDDA.n457 92.5005
R5183 VDDA.n457 VDDA.n456 92.5005
R5184 VDDA.n438 VDDA.n437 92.5005
R5185 VDDA.n440 VDDA.n439 92.5005
R5186 VDDA.n441 VDDA.n440 92.5005
R5187 VDDA.n436 VDDA.n406 92.5005
R5188 VDDA.n443 VDDA.n442 92.5005
R5189 VDDA.n442 VDDA.n441 92.5005
R5190 VDDA.n424 VDDA.n423 92.5005
R5191 VDDA.n426 VDDA.n425 92.5005
R5192 VDDA.n427 VDDA.n426 92.5005
R5193 VDDA.n422 VDDA.n417 92.5005
R5194 VDDA.n429 VDDA.n428 92.5005
R5195 VDDA.n428 VDDA.n427 92.5005
R5196 VDDA.n392 VDDA.n391 92.5005
R5197 VDDA.n387 VDDA.n386 92.5005
R5198 VDDA.n390 VDDA.n387 92.5005
R5199 VDDA.n389 VDDA.n388 92.5005
R5200 VDDA.n394 VDDA.n384 92.5005
R5201 VDDA.n390 VDDA.n384 92.5005
R5202 VDDA.n373 VDDA.n372 92.5005
R5203 VDDA.n375 VDDA.n374 92.5005
R5204 VDDA.n376 VDDA.n375 92.5005
R5205 VDDA.n371 VDDA.n340 92.5005
R5206 VDDA.n378 VDDA.n377 92.5005
R5207 VDDA.n377 VDDA.n376 92.5005
R5208 VDDA.n365 VDDA.n364 92.5005
R5209 VDDA.n360 VDDA.n359 92.5005
R5210 VDDA.n363 VDDA.n360 92.5005
R5211 VDDA.n362 VDDA.n361 92.5005
R5212 VDDA.n367 VDDA.n357 92.5005
R5213 VDDA.n363 VDDA.n357 92.5005
R5214 VDDA.n315 VDDA.n268 92.5005
R5215 VDDA.n318 VDDA.n317 92.5005
R5216 VDDA.n319 VDDA.n318 92.5005
R5217 VDDA.n267 VDDA.n260 92.5005
R5218 VDDA.n321 VDDA.n320 92.5005
R5219 VDDA.n320 VDDA.n319 92.5005
R5220 VDDA.n299 VDDA.n298 92.5005
R5221 VDDA.n295 VDDA.n294 92.5005
R5222 VDDA.n297 VDDA.n295 92.5005
R5223 VDDA.n296 VDDA.n288 92.5005
R5224 VDDA.n300 VDDA.n289 92.5005
R5225 VDDA.n297 VDDA.n289 92.5005
R5226 VDDA.n164 VDDA.t289 91.6672
R5227 VDDA.n164 VDDA.t154 91.6672
R5228 VDDA.n228 VDDA.n227 87.4672
R5229 VDDA.n319 VDDA.t248 86.3641
R5230 VDDA.n319 VDDA.t240 86.3641
R5231 VDDA.n297 VDDA.t211 86.3641
R5232 VDDA.t467 VDDA.n297 86.3641
R5233 VDDA.n227 VDDA.t18 85.438
R5234 VDDA.n239 VDDA.t33 85.438
R5235 VDDA.n233 VDDA.t17 81.3068
R5236 VDDA.n239 VDDA.n238 81.0672
R5237 VDDA.n229 VDDA.n227 81.0672
R5238 VDDA.n376 VDDA.t341 79.907
R5239 VDDA.n376 VDDA.t159 79.907
R5240 VDDA.n456 VDDA.t351 79.1672
R5241 VDDA.n390 VDDA.t155 79.1672
R5242 VDDA.t379 VDDA.n390 79.1672
R5243 VDDA.n363 VDDA.t464 79.1672
R5244 VDDA.t465 VDDA.n363 79.1672
R5245 VDDA.n178 VDDA.t183 78.8005
R5246 VDDA.n178 VDDA.t359 78.8005
R5247 VDDA.n184 VDDA.t137 78.8005
R5248 VDDA.n184 VDDA.t139 78.8005
R5249 VDDA.n186 VDDA.t189 78.8005
R5250 VDDA.n186 VDDA.t326 78.8005
R5251 VDDA.n188 VDDA.t357 78.8005
R5252 VDDA.n188 VDDA.t177 78.8005
R5253 VDDA.n190 VDDA.t147 78.8005
R5254 VDDA.n190 VDDA.t221 78.8005
R5255 VDDA.n192 VDDA.t141 78.8005
R5256 VDDA.n192 VDDA.t330 78.8005
R5257 VDDA.n194 VDDA.t328 78.8005
R5258 VDDA.n194 VDDA.t219 78.8005
R5259 VDDA.n196 VDDA.t179 78.8005
R5260 VDDA.n196 VDDA.t135 78.8005
R5261 VDDA.n198 VDDA.t181 78.8005
R5262 VDDA.n198 VDDA.t149 78.8005
R5263 VDDA.n200 VDDA.t332 78.8005
R5264 VDDA.n200 VDDA.t187 78.8005
R5265 VDDA.n441 VDDA.t130 77.9856
R5266 VDDA.n441 VDDA.t283 77.9856
R5267 VDDA.n427 VDDA.t438 77.9856
R5268 VDDA.n427 VDDA.t274 77.9856
R5269 VDDA.n237 VDDA.n222 64.0005
R5270 VDDA.n367 VDDA.n366 64.0005
R5271 VDDA.n367 VDDA.n356 64.0005
R5272 VDDA.n334 VDDA.n333 64.0005
R5273 VDDA.n333 VDDA.n330 64.0005
R5274 VDDA.n330 VDDA.n261 64.0005
R5275 VDDA.n321 VDDA.n261 64.0005
R5276 VDDA.n321 VDDA.n266 64.0005
R5277 VDDA.n275 VDDA.n266 64.0005
R5278 VDDA.n275 VDDA.n272 64.0005
R5279 VDDA.n314 VDDA.n272 64.0005
R5280 VDDA.t312 VDDA.t44 62.9523
R5281 VDDA.t394 VDDA.t312 62.9523
R5282 VDDA.t317 VDDA.t394 62.9523
R5283 VDDA.t405 VDDA.t317 62.9523
R5284 VDDA.t207 VDDA.t405 62.9523
R5285 VDDA.t225 VDDA.t260 62.9523
R5286 VDDA.t260 VDDA.t306 62.9523
R5287 VDDA.t306 VDDA.t310 62.9523
R5288 VDDA.t310 VDDA.t205 62.9523
R5289 VDDA.t205 VDDA.t59 62.9523
R5290 VDDA.t293 VDDA.t62 62.9523
R5291 VDDA.t461 VDDA.t293 62.9523
R5292 VDDA.t128 VDDA.t461 62.9523
R5293 VDDA.t315 VDDA.t128 62.9523
R5294 VDDA.t323 VDDA.t315 62.9523
R5295 VDDA.t447 VDDA.t277 62.9523
R5296 VDDA.t198 VDDA.t447 62.9523
R5297 VDDA.t269 VDDA.t198 62.9523
R5298 VDDA.t365 VDDA.t269 62.9523
R5299 VDDA.t90 VDDA.t365 62.9523
R5300 VDDA.n394 VDDA.n393 62.7205
R5301 VDDA.n394 VDDA.n383 62.7205
R5302 VDDA.n215 VDDA.t376 62.5402
R5303 VDDA.n215 VDDA.t87 62.5402
R5304 VDDA.n246 VDDA.n245 61.6672
R5305 VDDA.n248 VDDA.n247 61.6672
R5306 VDDA.n137 VDDA.n112 61.6672
R5307 VDDA.n139 VDDA.n138 61.6672
R5308 VDDA.n45 VDDA.n44 61.6672
R5309 VDDA.n42 VDDA.n41 61.6672
R5310 VDDA.n122 VDDA.t227 60.7563
R5311 VDDA.t224 VDDA.n122 60.7563
R5312 VDDA.n22 VDDA.t158 60.7563
R5313 VDDA.t314 VDDA.n22 60.7563
R5314 VDDA.n254 VDDA.t470 59.5681
R5315 VDDA.n255 VDDA.t471 59.5681
R5316 VDDA.n244 VDDA.n217 57.6005
R5317 VDDA.n249 VDDA.n217 57.6005
R5318 VDDA.n455 VDDA.t122 57.5763
R5319 VDDA.n254 VDDA.t472 51.8887
R5320 VDDA.n230 VDDA.n222 51.2005
R5321 VDDA.n102 VDDA.t429 49.1384
R5322 VDDA.t184 VDDA.n102 49.1384
R5323 VDDA.n78 VDDA.t333 49.1384
R5324 VDDA.t194 VDDA.n78 49.1384
R5325 VDDA.n256 VDDA.t469 48.9557
R5326 VDDA.n252 VDDA.n251 48.3605
R5327 VDDA.n242 VDDA.n241 43.8605
R5328 VDDA.n202 VDDA.n201 42.0963
R5329 VDDA.n213 VDDA.n212 41.5338
R5330 VDDA.n399 VDDA.t370 39.4005
R5331 VDDA.n399 VDDA.t352 39.4005
R5332 VDDA.n402 VDDA.t123 39.4005
R5333 VDDA.n402 VDDA.t450 39.4005
R5334 VDDA.n404 VDDA.t133 39.4005
R5335 VDDA.n404 VDDA.t372 39.4005
R5336 VDDA.n407 VDDA.t171 39.4005
R5337 VDDA.n407 VDDA.t131 39.4005
R5338 VDDA.n409 VDDA.t284 39.4005
R5339 VDDA.n409 VDDA.t153 39.4005
R5340 VDDA.n411 VDDA.t193 39.4005
R5341 VDDA.n411 VDDA.t414 39.4005
R5342 VDDA.n413 VDDA.t374 39.4005
R5343 VDDA.n413 VDDA.t191 39.4005
R5344 VDDA.n415 VDDA.t390 39.4005
R5345 VDDA.n415 VDDA.t439 39.4005
R5346 VDDA.n418 VDDA.t275 39.4005
R5347 VDDA.n418 VDDA.t441 39.4005
R5348 VDDA.n395 VDDA.t156 39.4005
R5349 VDDA.n395 VDDA.t380 39.4005
R5350 VDDA.n278 VDDA.t247 39.4005
R5351 VDDA.n278 VDDA.t251 39.4005
R5352 VDDA.n274 VDDA.t422 39.4005
R5353 VDDA.n274 VDDA.t253 39.4005
R5354 VDDA.n264 VDDA.t237 39.4005
R5355 VDDA.n264 VDDA.t426 39.4005
R5356 VDDA.n263 VDDA.t249 39.4005
R5357 VDDA.n263 VDDA.t241 39.4005
R5358 VDDA.n324 VDDA.t424 39.4005
R5359 VDDA.n324 VDDA.t255 39.4005
R5360 VDDA.n328 VDDA.t257 39.4005
R5361 VDDA.n328 VDDA.t428 39.4005
R5362 VDDA.n331 VDDA.t239 39.4005
R5363 VDDA.n331 VDDA.t259 39.4005
R5364 VDDA.n259 VDDA.t420 39.4005
R5365 VDDA.n259 VDDA.t243 39.4005
R5366 VDDA.n273 VDDA.t245 39.4005
R5367 VDDA.n273 VDDA.t418 39.4005
R5368 VDDA.n310 VDDA.t304 39.4005
R5369 VDDA.n310 VDDA.t437 39.4005
R5370 VDDA.n308 VDDA.t286 39.4005
R5371 VDDA.n308 VDDA.t223 39.4005
R5372 VDDA.n306 VDDA.t292 39.4005
R5373 VDDA.n306 VDDA.t4 39.4005
R5374 VDDA.n304 VDDA.t210 39.4005
R5375 VDDA.n304 VDDA.t435 39.4005
R5376 VDDA.n301 VDDA.t212 39.4005
R5377 VDDA.n301 VDDA.t468 39.4005
R5378 VDDA.n286 VDDA.t432 39.4005
R5379 VDDA.n286 VDDA.t6 39.4005
R5380 VDDA.n284 VDDA.t281 39.4005
R5381 VDDA.n284 VDDA.t288 39.4005
R5382 VDDA.n282 VDDA.t214 39.4005
R5383 VDDA.n282 VDDA.t169 39.4005
R5384 VDDA.n281 VDDA.t388 39.4005
R5385 VDDA.n281 VDDA.t272 39.4005
R5386 VDDA.n142 VDDA.t207 31.4764
R5387 VDDA.n142 VDDA.t225 31.4764
R5388 VDDA.n43 VDDA.t323 31.4764
R5389 VDDA.t277 VDDA.n43 31.4764
R5390 VDDA.n169 VDDA.n168 28.663
R5391 VDDA.n468 VDDA.n257 28.3337
R5392 VDDA.n251 VDDA.n250 25.6005
R5393 VDDA.n243 VDDA.n242 25.6005
R5394 VDDA.n212 VDDA.n211 25.6005
R5395 VDDA.n203 VDDA.n202 25.6005
R5396 VDDA.n250 VDDA.n249 24.5338
R5397 VDDA.n244 VDDA.n243 24.5338
R5398 VDDA.n238 VDDA.n237 24.5338
R5399 VDDA.n230 VDDA.n229 24.5338
R5400 VDDA VDDA.n253 22.2202
R5401 VDDA.n456 VDDA.n455 21.5914
R5402 VDDA.n211 VDDA.n210 21.3338
R5403 VDDA.n204 VDDA.n203 21.3338
R5404 VDDA.n160 VDDA.n159 21.3338
R5405 VDDA.n167 VDDA.n158 21.3338
R5406 VDDA.n155 VDDA.n154 21.3338
R5407 VDDA.n175 VDDA.n153 21.3338
R5408 VDDA.n118 VDDA.n117 21.3338
R5409 VDDA.n116 VDDA.n115 21.3338
R5410 VDDA.n146 VDDA.n145 21.3338
R5411 VDDA.n136 VDDA.n135 21.3338
R5412 VDDA.n98 VDDA.n97 21.3338
R5413 VDDA.n96 VDDA.n95 21.3338
R5414 VDDA.n74 VDDA.n73 21.3338
R5415 VDDA.n72 VDDA.n71 21.3338
R5416 VDDA.n18 VDDA.n17 21.3338
R5417 VDDA.n16 VDDA.n15 21.3338
R5418 VDDA.n47 VDDA.n46 21.3338
R5419 VDDA.n40 VDDA.n39 21.3338
R5420 VDDA.n383 VDDA.n382 21.3338
R5421 VDDA.n393 VDDA.n385 21.3338
R5422 VDDA.n356 VDDA.n355 21.3338
R5423 VDDA.n366 VDDA.n358 21.3338
R5424 VDDA.n270 VDDA.n269 21.3338
R5425 VDDA.n316 VDDA.n271 21.3338
R5426 VDDA.n293 VDDA.n292 21.3338
R5427 VDDA.n291 VDDA.n290 21.3338
R5428 VDDA.n61 VDDA.n60 21.1567
R5429 VDDA.n177 VDDA.n176 19.5505
R5430 VDDA.n144 VDDA.n125 19.538
R5431 VDDA.n26 VDDA.n25 19.538
R5432 VDDA.n107 VDDA.n105 19.2005
R5433 VDDA.n83 VDDA.n81 19.2005
R5434 VDDA.n460 VDDA.n459 19.2005
R5435 VDDA.n449 VDDA.n448 19.2005
R5436 VDDA.n445 VDDA.n444 19.2005
R5437 VDDA.n435 VDDA.n434 19.2005
R5438 VDDA.n431 VDDA.n430 19.2005
R5439 VDDA.n421 VDDA.n420 19.2005
R5440 VDDA.n380 VDDA.n379 19.2005
R5441 VDDA.n370 VDDA.n369 19.2005
R5442 VDDA.n232 VDDA.n231 18.5005
R5443 VDDA.n236 VDDA.n235 18.5005
R5444 VDDA.t172 VDDA.n234 17.1176
R5445 VDDA.n150 VDDA.n10 16.8443
R5446 VDDA.n368 VDDA.n367 16.363
R5447 VDDA.n467 VDDA.t446 15.0181
R5448 VDDA.n420 VDDA.n419 14.363
R5449 VDDA.n228 VDDA.n221 14.0505
R5450 VDDA.n448 VDDA.n447 13.8005
R5451 VDDA.n434 VDDA.n433 13.8005
R5452 VDDA.n432 VDDA.n431 13.8005
R5453 VDDA.n446 VDDA.n445 13.8005
R5454 VDDA.n461 VDDA.n460 13.8005
R5455 VDDA.n369 VDDA.n368 13.8005
R5456 VDDA.n381 VDDA.n380 13.8005
R5457 VDDA.n338 VDDA.t346 13.1338
R5458 VDDA.n338 VDDA.t454 13.1338
R5459 VDDA.n341 VDDA.t166 13.1338
R5460 VDDA.n341 VDDA.t349 13.1338
R5461 VDDA.n343 VDDA.t363 13.1338
R5462 VDDA.n343 VDDA.t460 13.1338
R5463 VDDA.n345 VDDA.t300 13.1338
R5464 VDDA.n345 VDDA.t342 13.1338
R5465 VDDA.n347 VDDA.t160 13.1338
R5466 VDDA.n347 VDDA.t1 13.1338
R5467 VDDA.n349 VDDA.t229 13.1338
R5468 VDDA.n349 VDDA.t164 13.1338
R5469 VDDA.n351 VDDA.t162 13.1338
R5470 VDDA.n351 VDDA.t443 13.1338
R5471 VDDA.n353 VDDA.t384 13.1338
R5472 VDDA.n353 VDDA.t456 13.1338
R5473 VDDA.t18 VDDA.n226 12.313
R5474 VDDA.n226 VDDA.t173 12.313
R5475 VDDA.n106 VDDA.t430 11.2576
R5476 VDDA.n106 VDDA.t185 11.2576
R5477 VDDA.n90 VDDA.t400 11.2576
R5478 VDDA.n90 VDDA.t217 11.2576
R5479 VDDA.n89 VDDA.t197 11.2576
R5480 VDDA.n89 VDDA.t175 11.2576
R5481 VDDA.n87 VDDA.t127 11.2576
R5482 VDDA.n87 VDDA.t298 11.2576
R5483 VDDA.n86 VDDA.t416 11.2576
R5484 VDDA.n86 VDDA.t145 11.2576
R5485 VDDA.n82 VDDA.t334 11.2576
R5486 VDDA.n82 VDDA.t195 11.2576
R5487 VDDA.n66 VDDA.t408 11.2576
R5488 VDDA.n66 VDDA.t143 11.2576
R5489 VDDA.n65 VDDA.t338 11.2576
R5490 VDDA.n65 VDDA.t355 11.2576
R5491 VDDA.n63 VDDA.t378 11.2576
R5492 VDDA.n63 VDDA.t234 11.2576
R5493 VDDA.n62 VDDA.t402 11.2576
R5494 VDDA.n62 VDDA.t336 11.2576
R5495 VDDA.n108 VDDA.n107 9.3005
R5496 VDDA.n84 VDDA.n83 9.3005
R5497 VDDA.n396 VDDA.n394 9.3005
R5498 VDDA.n335 VDDA.n334 9.3005
R5499 VDDA.n333 VDDA.n332 9.3005
R5500 VDDA.n330 VDDA.n329 9.3005
R5501 VDDA.n325 VDDA.n261 9.3005
R5502 VDDA.n322 VDDA.n321 9.3005
R5503 VDDA.n266 VDDA.n265 9.3005
R5504 VDDA.n276 VDDA.n275 9.3005
R5505 VDDA.n279 VDDA.n272 9.3005
R5506 VDDA.n314 VDDA.n313 9.3005
R5507 VDDA.n302 VDDA.n300 9.3005
R5508 VDDA.n241 VDDA.n240 8.53175
R5509 VDDA.n257 VDDA.n256 8.03219
R5510 VDDA.n59 VDDA.t381 8.0005
R5511 VDDA.n59 VDDA.t412 8.0005
R5512 VDDA.n57 VDDA.t276 8.0005
R5513 VDDA.n57 VDDA.t282 8.0005
R5514 VDDA.n55 VDDA.t452 8.0005
R5515 VDDA.n55 VDDA.t279 8.0005
R5516 VDDA.n53 VDDA.t265 8.0005
R5517 VDDA.n53 VDDA.t302 8.0005
R5518 VDDA.n51 VDDA.t167 8.0005
R5519 VDDA.n51 VDDA.t200 8.0005
R5520 VDDA.n50 VDDA.t410 8.0005
R5521 VDDA.n50 VDDA.t339 8.0005
R5522 VDDA.n9 VDDA.t409 8.0005
R5523 VDDA.n9 VDDA.t308 8.0005
R5524 VDDA.n7 VDDA.t392 8.0005
R5525 VDDA.n7 VDDA.t309 8.0005
R5526 VDDA.n5 VDDA.t393 8.0005
R5527 VDDA.n5 VDDA.t262 8.0005
R5528 VDDA.n3 VDDA.t397 8.0005
R5529 VDDA.n3 VDDA.t263 8.0005
R5530 VDDA.n1 VDDA.t396 8.0005
R5531 VDDA.n1 VDDA.t319 8.0005
R5532 VDDA.n0 VDDA.t151 8.0005
R5533 VDDA.n0 VDDA.t411 8.0005
R5534 VDDA.n462 VDDA.n461 7.44175
R5535 VDDA.n214 VDDA.n213 7.438
R5536 VDDA.n110 VDDA.t313 6.56717
R5537 VDDA.n110 VDDA.t395 6.56717
R5538 VDDA.n126 VDDA.t318 6.56717
R5539 VDDA.n126 VDDA.t406 6.56717
R5540 VDDA.n128 VDDA.t208 6.56717
R5541 VDDA.n128 VDDA.t226 6.56717
R5542 VDDA.n130 VDDA.t261 6.56717
R5543 VDDA.n130 VDDA.t307 6.56717
R5544 VDDA.n132 VDDA.t311 6.56717
R5545 VDDA.n132 VDDA.t206 6.56717
R5546 VDDA.n11 VDDA.t270 6.56717
R5547 VDDA.n11 VDDA.t366 6.56717
R5548 VDDA.n30 VDDA.t448 6.56717
R5549 VDDA.n30 VDDA.t199 6.56717
R5550 VDDA.n32 VDDA.t324 6.56717
R5551 VDDA.n32 VDDA.t278 6.56717
R5552 VDDA.n34 VDDA.t129 6.56717
R5553 VDDA.n34 VDDA.t316 6.56717
R5554 VDDA.n36 VDDA.t294 6.56717
R5555 VDDA.n36 VDDA.t462 6.56717
R5556 VDDA.n109 VDDA.n85 6.313
R5557 VDDA.n398 VDDA.n397 6.13371
R5558 VDDA.n337 VDDA.n336 6.098
R5559 VDDA.n253 VDDA.n252 6.0005
R5560 VDDA.n468 VDDA.n467 5.16125
R5561 VDDA.n241 VDDA.n216 5.1255
R5562 VDDA.n109 VDDA.n108 5.063
R5563 VDDA.n85 VDDA.n84 5.063
R5564 VDDA.n108 VDDA.n92 4.5005
R5565 VDDA.n84 VDDA.n68 4.5005
R5566 VDDA.n150 VDDA.n149 4.5005
R5567 VDDA.n397 VDDA.n396 4.5005
R5568 VDDA.n303 VDDA.n302 4.5005
R5569 VDDA.n313 VDDA.n312 4.5005
R5570 VDDA.n280 VDDA.n279 4.5005
R5571 VDDA.n277 VDDA.n276 4.5005
R5572 VDDA.n265 VDDA.n262 4.5005
R5573 VDDA.n323 VDDA.n322 4.5005
R5574 VDDA.n326 VDDA.n325 4.5005
R5575 VDDA.n329 VDDA.n327 4.5005
R5576 VDDA.n332 VDDA.n258 4.5005
R5577 VDDA.n336 VDDA.n335 4.5005
R5578 VDDA.n234 VDDA.n233 4.27978
R5579 VDDA.n255 VDDA.n254 4.12334
R5580 VDDA.n85 VDDA.n61 3.688
R5581 VDDA.n149 VDDA.n109 3.5005
R5582 VDDA.n312 VDDA.n311 3.3755
R5583 VDDA.n256 VDDA.n255 2.93377
R5584 VDDA.n214 VDDA.n177 2.813
R5585 VDDA.n253 VDDA.n214 2.563
R5586 VDDA.n447 VDDA.n446 2.5005
R5587 VDDA.n397 VDDA.n381 2.47371
R5588 VDDA.n433 VDDA.n432 1.813
R5589 VDDA.n177 VDDA.n150 1.46925
R5590 VDDA.n368 VDDA.n354 1.0005
R5591 VDDA.n354 VDDA.n352 1.0005
R5592 VDDA.n352 VDDA.n350 1.0005
R5593 VDDA.n350 VDDA.n348 1.0005
R5594 VDDA.n348 VDDA.n346 1.0005
R5595 VDDA.n346 VDDA.n344 1.0005
R5596 VDDA.n344 VDDA.n342 1.0005
R5597 VDDA.n342 VDDA.n339 1.0005
R5598 VDDA.n381 VDDA.n339 1.0005
R5599 VDDA.n149 VDDA.n148 0.938
R5600 VDDA.n337 VDDA.n257 0.840625
R5601 VDDA.n61 VDDA.n49 0.7505
R5602 VDDA.n398 VDDA.n337 0.74075
R5603 VDDA.n240 VDDA.n221 0.6255
R5604 VDDA.n92 VDDA.n91 0.6255
R5605 VDDA.n92 VDDA.n88 0.6255
R5606 VDDA.n68 VDDA.n67 0.6255
R5607 VDDA.n68 VDDA.n64 0.6255
R5608 VDDA.n285 VDDA.n283 0.6255
R5609 VDDA.n287 VDDA.n285 0.6255
R5610 VDDA.n303 VDDA.n287 0.6255
R5611 VDDA.n305 VDDA.n303 0.6255
R5612 VDDA.n307 VDDA.n305 0.6255
R5613 VDDA.n309 VDDA.n307 0.6255
R5614 VDDA.n311 VDDA.n309 0.6255
R5615 VDDA.n312 VDDA.n280 0.6255
R5616 VDDA.n280 VDDA.n277 0.6255
R5617 VDDA.n277 VDDA.n262 0.6255
R5618 VDDA.n323 VDDA.n262 0.6255
R5619 VDDA.n326 VDDA.n323 0.6255
R5620 VDDA.n327 VDDA.n326 0.6255
R5621 VDDA.n327 VDDA.n258 0.6255
R5622 VDDA.n336 VDDA.n258 0.6255
R5623 VDDA.n201 VDDA.n199 0.563
R5624 VDDA.n199 VDDA.n197 0.563
R5625 VDDA.n197 VDDA.n195 0.563
R5626 VDDA.n195 VDDA.n193 0.563
R5627 VDDA.n193 VDDA.n191 0.563
R5628 VDDA.n191 VDDA.n189 0.563
R5629 VDDA.n189 VDDA.n187 0.563
R5630 VDDA.n187 VDDA.n185 0.563
R5631 VDDA.n185 VDDA.n179 0.563
R5632 VDDA.n213 VDDA.n179 0.563
R5633 VDDA.n133 VDDA.n131 0.563
R5634 VDDA.n131 VDDA.n129 0.563
R5635 VDDA.n129 VDDA.n127 0.563
R5636 VDDA.n127 VDDA.n111 0.563
R5637 VDDA.n148 VDDA.n111 0.563
R5638 VDDA.n54 VDDA.n52 0.563
R5639 VDDA.n56 VDDA.n54 0.563
R5640 VDDA.n58 VDDA.n56 0.563
R5641 VDDA.n60 VDDA.n58 0.563
R5642 VDDA.n37 VDDA.n35 0.563
R5643 VDDA.n35 VDDA.n33 0.563
R5644 VDDA.n33 VDDA.n31 0.563
R5645 VDDA.n31 VDDA.n12 0.563
R5646 VDDA.n49 VDDA.n12 0.563
R5647 VDDA.n4 VDDA.n2 0.563
R5648 VDDA.n6 VDDA.n4 0.563
R5649 VDDA.n8 VDDA.n6 0.563
R5650 VDDA.n10 VDDA.n8 0.563
R5651 VDDA.n419 VDDA.n416 0.563
R5652 VDDA.n432 VDDA.n416 0.563
R5653 VDDA.n433 VDDA.n414 0.563
R5654 VDDA.n414 VDDA.n412 0.563
R5655 VDDA.n412 VDDA.n410 0.563
R5656 VDDA.n410 VDDA.n408 0.563
R5657 VDDA.n408 VDDA.n405 0.563
R5658 VDDA.n446 VDDA.n405 0.563
R5659 VDDA.n447 VDDA.n403 0.563
R5660 VDDA.n403 VDDA.n400 0.563
R5661 VDDA.n461 VDDA.n400 0.563
R5662 VDDA.n462 VDDA.n398 0.546875
R5663 VDDA.n467 VDDA.n462 0.370625
R5664 VDDA.n252 VDDA.n216 0.2505
R5665 VDDA.t385 VDDA.t444 0.1603
R5666 VDDA.t232 VDDA.t445 0.1603
R5667 VDDA.t230 VDDA.t295 0.1603
R5668 VDDA.t2 VDDA.t347 0.1603
R5669 VDDA.t296 VDDA.t231 0.1603
R5670 VDDA.t458 VDDA.t360 0.1603
R5671 VDDA.t382 VDDA.t301 0.1603
R5672 VDDA.t361 VDDA.t340 0.1603
R5673 VDDA.n464 VDDA.t364 0.159278
R5674 VDDA.n465 VDDA.t344 0.159278
R5675 VDDA.n466 VDDA.t386 0.159278
R5676 VDDA.n466 VDDA.t385 0.1368
R5677 VDDA.n466 VDDA.t232 0.1368
R5678 VDDA.n465 VDDA.t230 0.1368
R5679 VDDA.n465 VDDA.t2 0.1368
R5680 VDDA.n464 VDDA.t296 0.1368
R5681 VDDA.n464 VDDA.t458 0.1368
R5682 VDDA.n463 VDDA.t382 0.1368
R5683 VDDA.n463 VDDA.t361 0.1368
R5684 VDDA VDDA.n468 0.024
R5685 VDDA.t364 VDDA.n463 0.00152174
R5686 VDDA.t344 VDDA.n464 0.00152174
R5687 VDDA.t386 VDDA.n465 0.00152174
R5688 VDDA.t446 VDDA.n466 0.00152174
R5689 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 394.166
R5690 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t2 384.967
R5691 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t19 369.534
R5692 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t9 369.534
R5693 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t18 369.534
R5694 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t8 369.534
R5695 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t23 369.534
R5696 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.n18 369.534
R5697 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t5 192.8
R5698 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t15 192.8
R5699 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t7 192.8
R5700 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t17 192.8
R5701 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t10 192.8
R5702 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t21 192.8
R5703 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t12 192.8
R5704 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t16 192.8
R5705 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t11 192.8
R5706 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t22 192.8
R5707 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 192.8
R5708 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t14 192.8
R5709 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t6 192.8
R5710 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t20 192.8
R5711 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R5712 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R5713 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R5714 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R5715 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R5716 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R5717 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R5718 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R5719 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R5720 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R5721 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R5722 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.n19 126.876
R5723 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R5724 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R5725 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R5726 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R5727 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R5728 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R5729 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t1 39.4005
R5730 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t0 39.4005
R5731 bgr_0.NFET_GATE_10uA.t3 bgr_0.NFET_GATE_10uA.n20 24.0005
R5732 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 24.0005
R5733 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 144.827
R5734 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 134.577
R5735 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 120.66
R5736 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 97.4009
R5737 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 96.8384
R5738 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 96.8384
R5739 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 96.8384
R5740 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 96.8384
R5741 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 64.5005
R5742 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 24.0005
R5743 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 24.0005
R5744 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R5745 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 24.0005
R5746 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R5747 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 8.0005
R5748 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R5749 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 8.0005
R5750 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R5751 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 8.0005
R5752 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R5753 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 8.0005
R5754 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R5755 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R5756 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 5.813
R5757 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 0.563
R5758 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 0.563
R5759 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.563
R5760 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 114.719
R5761 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5762 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5763 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 114.156
R5764 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5765 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5766 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5767 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5768 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5769 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5770 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5771 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5772 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5773 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5774 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5775 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5776 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5777 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5778 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5779 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5780 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5781 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5782 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5783 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5784 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5785 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5786 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5787 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5788 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5789 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5790 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5791 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5792 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5793 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5794 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5795 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5796 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5797 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5798 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5799 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5800 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n8 0.563
R5801 VOUT-.n14 VOUT-.n6 145.989
R5802 VOUT-.n9 VOUT-.n7 145.989
R5803 VOUT-.n13 VOUT-.n12 145.427
R5804 VOUT-.n11 VOUT-.n10 145.427
R5805 VOUT-.n9 VOUT-.n8 145.427
R5806 VOUT-.n16 VOUT-.n15 140.927
R5807 VOUT-.n5 VOUT-.t4 113.192
R5808 VOUT-.n2 VOUT-.n0 95.7303
R5809 VOUT-.n4 VOUT-.n3 94.6053
R5810 VOUT-.n2 VOUT-.n1 94.6053
R5811 VOUT-.n100 VOUT-.n16 20.5943
R5812 VOUT-.n100 VOUT-.n99 11.7059
R5813 VOUT- VOUT-.n100 7.813
R5814 VOUT-.n15 VOUT-.t15 6.56717
R5815 VOUT-.n15 VOUT-.t12 6.56717
R5816 VOUT-.n12 VOUT-.t16 6.56717
R5817 VOUT-.n12 VOUT-.t3 6.56717
R5818 VOUT-.n10 VOUT-.t5 6.56717
R5819 VOUT-.n10 VOUT-.t7 6.56717
R5820 VOUT-.n8 VOUT-.t9 6.56717
R5821 VOUT-.n8 VOUT-.t10 6.56717
R5822 VOUT-.n7 VOUT-.t2 6.56717
R5823 VOUT-.n7 VOUT-.t1 6.56717
R5824 VOUT-.n6 VOUT-.t0 6.56717
R5825 VOUT-.n6 VOUT-.t11 6.56717
R5826 VOUT-.n46 VOUT-.t83 4.8295
R5827 VOUT-.n48 VOUT-.t90 4.8295
R5828 VOUT-.n51 VOUT-.t128 4.8295
R5829 VOUT-.n54 VOUT-.t26 4.8295
R5830 VOUT-.n57 VOUT-.t74 4.8295
R5831 VOUT-.n70 VOUT-.t39 4.8295
R5832 VOUT-.n72 VOUT-.t34 4.8295
R5833 VOUT-.n73 VOUT-.t136 4.8295
R5834 VOUT-.n75 VOUT-.t68 4.8295
R5835 VOUT-.n76 VOUT-.t36 4.8295
R5836 VOUT-.n78 VOUT-.t94 4.8295
R5837 VOUT-.n79 VOUT-.t64 4.8295
R5838 VOUT-.n81 VOUT-.t54 4.8295
R5839 VOUT-.n82 VOUT-.t29 4.8295
R5840 VOUT-.n84 VOUT-.t89 4.8295
R5841 VOUT-.n85 VOUT-.t57 4.8295
R5842 VOUT-.n87 VOUT-.t48 4.8295
R5843 VOUT-.n88 VOUT-.t20 4.8295
R5844 VOUT-.n90 VOUT-.t148 4.8295
R5845 VOUT-.n91 VOUT-.t121 4.8295
R5846 VOUT-.n93 VOUT-.t43 4.8295
R5847 VOUT-.n94 VOUT-.t152 4.8295
R5848 VOUT-.n17 VOUT-.t107 4.8295
R5849 VOUT-.n29 VOUT-.t28 4.8295
R5850 VOUT-.n31 VOUT-.t24 4.8295
R5851 VOUT-.n32 VOUT-.t129 4.8295
R5852 VOUT-.n34 VOUT-.t59 4.8295
R5853 VOUT-.n35 VOUT-.t32 4.8295
R5854 VOUT-.n37 VOUT-.t99 4.8295
R5855 VOUT-.n38 VOUT-.t69 4.8295
R5856 VOUT-.n40 VOUT-.t67 4.8295
R5857 VOUT-.n41 VOUT-.t35 4.8295
R5858 VOUT-.n43 VOUT-.t104 4.8295
R5859 VOUT-.n44 VOUT-.t76 4.8295
R5860 VOUT-.n96 VOUT-.t115 4.8295
R5861 VOUT-.n69 VOUT-.t132 4.806
R5862 VOUT-.n68 VOUT-.t114 4.806
R5863 VOUT-.n67 VOUT-.t146 4.806
R5864 VOUT-.n66 VOUT-.t45 4.806
R5865 VOUT-.n65 VOUT-.t85 4.806
R5866 VOUT-.n64 VOUT-.t63 4.806
R5867 VOUT-.n63 VOUT-.t101 4.806
R5868 VOUT-.n62 VOUT-.t134 4.806
R5869 VOUT-.n61 VOUT-.t119 4.806
R5870 VOUT-.n60 VOUT-.t155 4.806
R5871 VOUT-.n28 VOUT-.t47 4.806
R5872 VOUT-.n27 VOUT-.t91 4.806
R5873 VOUT-.n26 VOUT-.t41 4.806
R5874 VOUT-.n25 VOUT-.t130 4.806
R5875 VOUT-.n24 VOUT-.t82 4.806
R5876 VOUT-.n23 VOUT-.t124 4.806
R5877 VOUT-.n22 VOUT-.t72 4.806
R5878 VOUT-.n21 VOUT-.t23 4.806
R5879 VOUT-.n20 VOUT-.t62 4.806
R5880 VOUT-.n19 VOUT-.t150 4.806
R5881 VOUT-.n47 VOUT-.t95 4.5005
R5882 VOUT-.n46 VOUT-.t56 4.5005
R5883 VOUT-.n48 VOUT-.t131 4.5005
R5884 VOUT-.n49 VOUT-.t103 4.5005
R5885 VOUT-.n50 VOUT-.t71 4.5005
R5886 VOUT-.n51 VOUT-.t31 4.5005
R5887 VOUT-.n52 VOUT-.t138 4.5005
R5888 VOUT-.n53 VOUT-.t106 4.5005
R5889 VOUT-.n54 VOUT-.t60 4.5005
R5890 VOUT-.n55 VOUT-.t40 4.5005
R5891 VOUT-.n56 VOUT-.t143 4.5005
R5892 VOUT-.n57 VOUT-.t113 4.5005
R5893 VOUT-.n58 VOUT-.t21 4.5005
R5894 VOUT-.n59 VOUT-.t125 4.5005
R5895 VOUT-.n60 VOUT-.t118 4.5005
R5896 VOUT-.n61 VOUT-.t80 4.5005
R5897 VOUT-.n62 VOUT-.t96 4.5005
R5898 VOUT-.n63 VOUT-.t61 4.5005
R5899 VOUT-.n64 VOUT-.t27 4.5005
R5900 VOUT-.n65 VOUT-.t44 4.5005
R5901 VOUT-.n66 VOUT-.t144 4.5005
R5902 VOUT-.n67 VOUT-.t111 4.5005
R5903 VOUT-.n68 VOUT-.t75 4.5005
R5904 VOUT-.n69 VOUT-.t92 4.5005
R5905 VOUT-.n71 VOUT-.t55 4.5005
R5906 VOUT-.n70 VOUT-.t19 4.5005
R5907 VOUT-.n72 VOUT-.t51 4.5005
R5908 VOUT-.n74 VOUT-.t156 4.5005
R5909 VOUT-.n73 VOUT-.t120 4.5005
R5910 VOUT-.n75 VOUT-.t87 4.5005
R5911 VOUT-.n77 VOUT-.t49 4.5005
R5912 VOUT-.n76 VOUT-.t151 4.5005
R5913 VOUT-.n78 VOUT-.t42 4.5005
R5914 VOUT-.n80 VOUT-.t145 4.5005
R5915 VOUT-.n79 VOUT-.t117 4.5005
R5916 VOUT-.n81 VOUT-.t141 4.5005
R5917 VOUT-.n83 VOUT-.t110 4.5005
R5918 VOUT-.n82 VOUT-.t79 4.5005
R5919 VOUT-.n84 VOUT-.t38 4.5005
R5920 VOUT-.n86 VOUT-.t139 4.5005
R5921 VOUT-.n85 VOUT-.t108 4.5005
R5922 VOUT-.n87 VOUT-.t135 4.5005
R5923 VOUT-.n89 VOUT-.t102 4.5005
R5924 VOUT-.n88 VOUT-.t70 4.5005
R5925 VOUT-.n90 VOUT-.t98 4.5005
R5926 VOUT-.n92 VOUT-.t66 4.5005
R5927 VOUT-.n91 VOUT-.t33 4.5005
R5928 VOUT-.n93 VOUT-.t133 4.5005
R5929 VOUT-.n95 VOUT-.t97 4.5005
R5930 VOUT-.n94 VOUT-.t65 4.5005
R5931 VOUT-.n18 VOUT-.t100 4.5005
R5932 VOUT-.n17 VOUT-.t149 4.5005
R5933 VOUT-.n19 VOUT-.t86 4.5005
R5934 VOUT-.n20 VOUT-.t50 4.5005
R5935 VOUT-.n21 VOUT-.t137 4.5005
R5936 VOUT-.n22 VOUT-.t105 4.5005
R5937 VOUT-.n23 VOUT-.t73 4.5005
R5938 VOUT-.n24 VOUT-.t25 4.5005
R5939 VOUT-.n25 VOUT-.t127 4.5005
R5940 VOUT-.n26 VOUT-.t88 4.5005
R5941 VOUT-.n27 VOUT-.t53 4.5005
R5942 VOUT-.n28 VOUT-.t140 4.5005
R5943 VOUT-.n30 VOUT-.t109 4.5005
R5944 VOUT-.n29 VOUT-.t78 4.5005
R5945 VOUT-.n31 VOUT-.t112 4.5005
R5946 VOUT-.n33 VOUT-.t77 4.5005
R5947 VOUT-.n32 VOUT-.t37 4.5005
R5948 VOUT-.n34 VOUT-.t147 4.5005
R5949 VOUT-.n36 VOUT-.t116 4.5005
R5950 VOUT-.n35 VOUT-.t81 4.5005
R5951 VOUT-.n37 VOUT-.t46 4.5005
R5952 VOUT-.n39 VOUT-.t153 4.5005
R5953 VOUT-.n38 VOUT-.t122 4.5005
R5954 VOUT-.n40 VOUT-.t154 4.5005
R5955 VOUT-.n42 VOUT-.t123 4.5005
R5956 VOUT-.n41 VOUT-.t84 4.5005
R5957 VOUT-.n43 VOUT-.t52 4.5005
R5958 VOUT-.n45 VOUT-.t22 4.5005
R5959 VOUT-.n44 VOUT-.t126 4.5005
R5960 VOUT-.n99 VOUT-.t142 4.5005
R5961 VOUT-.n98 VOUT-.t93 4.5005
R5962 VOUT-.n97 VOUT-.t58 4.5005
R5963 VOUT-.n96 VOUT-.t30 4.5005
R5964 VOUT-.n16 VOUT-.n14 4.5005
R5965 VOUT-.n3 VOUT-.t14 3.42907
R5966 VOUT-.n3 VOUT-.t17 3.42907
R5967 VOUT-.n1 VOUT-.t6 3.42907
R5968 VOUT-.n1 VOUT-.t13 3.42907
R5969 VOUT-.n0 VOUT-.t18 3.42907
R5970 VOUT-.n0 VOUT-.t8 3.42907
R5971 VOUT- VOUT-.n5 2.84425
R5972 VOUT-.n5 VOUT-.n4 2.03175
R5973 VOUT-.n4 VOUT-.n2 1.1255
R5974 VOUT-.n11 VOUT-.n9 0.563
R5975 VOUT-.n13 VOUT-.n11 0.563
R5976 VOUT-.n14 VOUT-.n13 0.563
R5977 VOUT-.n47 VOUT-.n46 0.3295
R5978 VOUT-.n50 VOUT-.n49 0.3295
R5979 VOUT-.n49 VOUT-.n48 0.3295
R5980 VOUT-.n53 VOUT-.n52 0.3295
R5981 VOUT-.n52 VOUT-.n51 0.3295
R5982 VOUT-.n56 VOUT-.n55 0.3295
R5983 VOUT-.n55 VOUT-.n54 0.3295
R5984 VOUT-.n59 VOUT-.n58 0.3295
R5985 VOUT-.n58 VOUT-.n57 0.3295
R5986 VOUT-.n61 VOUT-.n60 0.3295
R5987 VOUT-.n62 VOUT-.n61 0.3295
R5988 VOUT-.n63 VOUT-.n62 0.3295
R5989 VOUT-.n64 VOUT-.n63 0.3295
R5990 VOUT-.n65 VOUT-.n64 0.3295
R5991 VOUT-.n66 VOUT-.n65 0.3295
R5992 VOUT-.n67 VOUT-.n66 0.3295
R5993 VOUT-.n68 VOUT-.n67 0.3295
R5994 VOUT-.n69 VOUT-.n68 0.3295
R5995 VOUT-.n71 VOUT-.n69 0.3295
R5996 VOUT-.n71 VOUT-.n70 0.3295
R5997 VOUT-.n74 VOUT-.n72 0.3295
R5998 VOUT-.n74 VOUT-.n73 0.3295
R5999 VOUT-.n77 VOUT-.n75 0.3295
R6000 VOUT-.n77 VOUT-.n76 0.3295
R6001 VOUT-.n80 VOUT-.n78 0.3295
R6002 VOUT-.n80 VOUT-.n79 0.3295
R6003 VOUT-.n83 VOUT-.n81 0.3295
R6004 VOUT-.n83 VOUT-.n82 0.3295
R6005 VOUT-.n86 VOUT-.n84 0.3295
R6006 VOUT-.n86 VOUT-.n85 0.3295
R6007 VOUT-.n89 VOUT-.n87 0.3295
R6008 VOUT-.n89 VOUT-.n88 0.3295
R6009 VOUT-.n92 VOUT-.n90 0.3295
R6010 VOUT-.n92 VOUT-.n91 0.3295
R6011 VOUT-.n95 VOUT-.n93 0.3295
R6012 VOUT-.n95 VOUT-.n94 0.3295
R6013 VOUT-.n18 VOUT-.n17 0.3295
R6014 VOUT-.n20 VOUT-.n19 0.3295
R6015 VOUT-.n21 VOUT-.n20 0.3295
R6016 VOUT-.n22 VOUT-.n21 0.3295
R6017 VOUT-.n23 VOUT-.n22 0.3295
R6018 VOUT-.n24 VOUT-.n23 0.3295
R6019 VOUT-.n25 VOUT-.n24 0.3295
R6020 VOUT-.n26 VOUT-.n25 0.3295
R6021 VOUT-.n27 VOUT-.n26 0.3295
R6022 VOUT-.n28 VOUT-.n27 0.3295
R6023 VOUT-.n30 VOUT-.n28 0.3295
R6024 VOUT-.n30 VOUT-.n29 0.3295
R6025 VOUT-.n33 VOUT-.n31 0.3295
R6026 VOUT-.n33 VOUT-.n32 0.3295
R6027 VOUT-.n36 VOUT-.n34 0.3295
R6028 VOUT-.n36 VOUT-.n35 0.3295
R6029 VOUT-.n39 VOUT-.n37 0.3295
R6030 VOUT-.n39 VOUT-.n38 0.3295
R6031 VOUT-.n42 VOUT-.n40 0.3295
R6032 VOUT-.n42 VOUT-.n41 0.3295
R6033 VOUT-.n45 VOUT-.n43 0.3295
R6034 VOUT-.n45 VOUT-.n44 0.3295
R6035 VOUT-.n99 VOUT-.n98 0.3295
R6036 VOUT-.n98 VOUT-.n97 0.3295
R6037 VOUT-.n97 VOUT-.n96 0.3295
R6038 VOUT-.n67 VOUT-.n50 0.306
R6039 VOUT-.n66 VOUT-.n53 0.306
R6040 VOUT-.n65 VOUT-.n56 0.306
R6041 VOUT-.n64 VOUT-.n59 0.306
R6042 VOUT-.n71 VOUT-.n47 0.2825
R6043 VOUT-.n74 VOUT-.n71 0.2825
R6044 VOUT-.n77 VOUT-.n74 0.2825
R6045 VOUT-.n80 VOUT-.n77 0.2825
R6046 VOUT-.n83 VOUT-.n80 0.2825
R6047 VOUT-.n86 VOUT-.n83 0.2825
R6048 VOUT-.n89 VOUT-.n86 0.2825
R6049 VOUT-.n92 VOUT-.n89 0.2825
R6050 VOUT-.n95 VOUT-.n92 0.2825
R6051 VOUT-.n30 VOUT-.n18 0.2825
R6052 VOUT-.n33 VOUT-.n30 0.2825
R6053 VOUT-.n36 VOUT-.n33 0.2825
R6054 VOUT-.n39 VOUT-.n36 0.2825
R6055 VOUT-.n42 VOUT-.n39 0.2825
R6056 VOUT-.n45 VOUT-.n42 0.2825
R6057 VOUT-.n97 VOUT-.n45 0.2825
R6058 VOUT-.n97 VOUT-.n95 0.2825
R6059 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.083
R6060 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1603
R6061 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1603
R6062 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R6063 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R6064 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R6065 two_stage_opamp_dummy_magic_0.cap_res_X.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R6066 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R6067 two_stage_opamp_dummy_magic_0.cap_res_X.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1603
R6068 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R6069 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.1603
R6070 two_stage_opamp_dummy_magic_0.cap_res_X.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1603
R6071 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1603
R6072 two_stage_opamp_dummy_magic_0.cap_res_X.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R6073 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1603
R6074 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R6075 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1603
R6076 two_stage_opamp_dummy_magic_0.cap_res_X.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1603
R6077 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R6078 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1603
R6079 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1603
R6080 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R6081 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R6082 two_stage_opamp_dummy_magic_0.cap_res_X.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R6083 two_stage_opamp_dummy_magic_0.cap_res_X.t3 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R6084 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R6085 two_stage_opamp_dummy_magic_0.cap_res_X.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R6086 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R6087 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R6088 two_stage_opamp_dummy_magic_0.cap_res_X.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1603
R6089 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1603
R6090 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R6091 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.1603
R6092 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R6093 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R6094 two_stage_opamp_dummy_magic_0.cap_res_X.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R6095 two_stage_opamp_dummy_magic_0.cap_res_X.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.1603
R6096 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.1603
R6097 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1603
R6098 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R6099 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R6100 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1603
R6101 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R6102 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.1603
R6103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R6104 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1603
R6105 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R6106 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R6107 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1603
R6108 two_stage_opamp_dummy_magic_0.cap_res_X.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R6109 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R6110 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R6111 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R6112 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1603
R6113 two_stage_opamp_dummy_magic_0.cap_res_X.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R6114 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R6115 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R6116 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R6117 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.1603
R6118 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.159278
R6119 two_stage_opamp_dummy_magic_0.cap_res_X.t48 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R6120 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R6121 two_stage_opamp_dummy_magic_0.cap_res_X.t41 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R6122 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R6123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R6124 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R6125 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R6126 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R6127 two_stage_opamp_dummy_magic_0.cap_res_X.t91 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R6128 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R6129 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.159278
R6130 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.159278
R6131 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.159278
R6132 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.159278
R6133 two_stage_opamp_dummy_magic_0.cap_res_X.t1 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.159278
R6134 two_stage_opamp_dummy_magic_0.cap_res_X.t102 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.159278
R6135 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.159278
R6136 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.159278
R6137 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.159278
R6138 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.159278
R6139 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.159278
R6140 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.159278
R6141 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.159278
R6142 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.159278
R6143 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.159278
R6144 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.159278
R6145 two_stage_opamp_dummy_magic_0.cap_res_X.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.137822
R6146 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1368
R6147 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.1368
R6148 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.1368
R6149 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1368
R6150 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.1368
R6151 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1368
R6152 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1368
R6153 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R6154 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R6155 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1368
R6156 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R6157 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1368
R6158 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R6159 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R6160 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1368
R6161 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1368
R6162 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R6163 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R6164 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.1368
R6165 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R6166 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R6167 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1368
R6168 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1368
R6169 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1368
R6170 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1368
R6171 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R6172 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1368
R6173 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1368
R6174 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1368
R6175 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R6176 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R6177 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.118
R6178 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.114322
R6179 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R6180 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R6181 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R6182 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.1133
R6183 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.1133
R6184 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.1133
R6185 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.1133
R6186 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.1133
R6187 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.1133
R6188 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R6189 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R6190 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R6191 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R6192 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R6193 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R6194 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R6195 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R6196 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R6197 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R6198 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.00152174
R6199 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.00152174
R6200 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.00152174
R6201 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.00152174
R6202 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R6203 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R6204 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.00152174
R6205 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.00152174
R6206 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R6207 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.00152174
R6208 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.00152174
R6209 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R6210 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.00152174
R6211 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R6212 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.00152174
R6213 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.00152174
R6214 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R6215 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R6216 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.00152174
R6217 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.00152174
R6218 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R6219 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R6220 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R6221 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.00152174
R6222 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R6223 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.00152174
R6224 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.00152174
R6225 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R6226 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R6227 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.00152174
R6228 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.00152174
R6229 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.00152174
R6230 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R6231 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R6232 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.00152174
R6233 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R6234 bgr_0.cap_res2.t0 bgr_0.cap_res2.t17 188.573
R6235 bgr_0.cap_res2.t12 bgr_0.cap_res2.t13 0.1603
R6236 bgr_0.cap_res2.t1 bgr_0.cap_res2.t6 0.1603
R6237 bgr_0.cap_res2.t5 bgr_0.cap_res2.t8 0.1603
R6238 bgr_0.cap_res2.t16 bgr_0.cap_res2.t20 0.1603
R6239 bgr_0.cap_res2.t18 bgr_0.cap_res2.t2 0.1603
R6240 bgr_0.cap_res2.t10 bgr_0.cap_res2.t15 0.1603
R6241 bgr_0.cap_res2.t3 bgr_0.cap_res2.t7 0.1603
R6242 bgr_0.cap_res2.t14 bgr_0.cap_res2.t19 0.1603
R6243 bgr_0.cap_res2.n1 bgr_0.cap_res2.t9 0.159278
R6244 bgr_0.cap_res2.n2 bgr_0.cap_res2.t4 0.159278
R6245 bgr_0.cap_res2.n3 bgr_0.cap_res2.t11 0.159278
R6246 bgr_0.cap_res2.n3 bgr_0.cap_res2.t12 0.1368
R6247 bgr_0.cap_res2.n3 bgr_0.cap_res2.t1 0.1368
R6248 bgr_0.cap_res2.n2 bgr_0.cap_res2.t5 0.1368
R6249 bgr_0.cap_res2.n2 bgr_0.cap_res2.t16 0.1368
R6250 bgr_0.cap_res2.n1 bgr_0.cap_res2.t18 0.1368
R6251 bgr_0.cap_res2.n1 bgr_0.cap_res2.t10 0.1368
R6252 bgr_0.cap_res2.n0 bgr_0.cap_res2.t3 0.1368
R6253 bgr_0.cap_res2.n0 bgr_0.cap_res2.t14 0.1368
R6254 bgr_0.cap_res2.t9 bgr_0.cap_res2.n0 0.00152174
R6255 bgr_0.cap_res2.t4 bgr_0.cap_res2.n1 0.00152174
R6256 bgr_0.cap_res2.t11 bgr_0.cap_res2.n2 0.00152174
R6257 bgr_0.cap_res2.t17 bgr_0.cap_res2.n3 0.00152174
R6258 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 688.859
R6259 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 514.134
R6260 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 323.491
R6261 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 322.692
R6262 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6263 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6264 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 270.591
R6265 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 270.591
R6266 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 233.374
R6267 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 233.374
R6268 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 233.374
R6269 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 233.374
R6270 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 208.838
R6271 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 197.964
R6272 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 174.726
R6273 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6274 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 174.726
R6275 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 174.726
R6276 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 169.215
R6277 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 169.215
R6278 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 169.215
R6279 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 129.24
R6280 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 129.24
R6281 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6282 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6283 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 128.534
R6284 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 128.534
R6285 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 16.8443
R6286 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6287 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 13.1338
R6288 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6289 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6290 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6291 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6292 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 4.3755
R6293 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 4.3755
R6294 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 3.688
R6295 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 3.2505
R6296 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 3.1255
R6297 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 1.2755
R6298 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 1.2755
R6299 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 0.8005
R6300 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 632.186
R6301 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6302 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6303 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 630.264
R6304 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 628.003
R6305 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 628.003
R6306 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 626.753
R6307 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 626.753
R6308 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 625.756
R6309 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 622.231
R6310 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6311 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6312 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6313 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6314 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6315 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6316 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6317 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6318 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6319 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6320 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6321 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6322 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6323 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6324 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6325 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6326 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6327 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6328 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6329 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6330 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 7.94147
R6331 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 6.188
R6332 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 630.857
R6333 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 626.784
R6334 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n28 626.784
R6335 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n29 626.784
R6336 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n5 626.784
R6337 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.n25 585
R6338 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6339 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6340 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 176.733
R6341 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6342 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6343 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6344 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6345 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6346 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6347 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6348 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6349 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6350 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6351 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6352 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6353 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6354 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6355 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.n20 176.733
R6356 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n24 162.214
R6357 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n3 135.827
R6358 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6359 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6360 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6361 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6362 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6363 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6364 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6365 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6366 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6367 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6368 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6369 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6370 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6371 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6372 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6373 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6374 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6375 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6376 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6377 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6378 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6379 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R6380 two_stage_opamp_dummy_magic_0.V_err_gate.n29 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6381 two_stage_opamp_dummy_magic_0.V_err_gate.n29 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6382 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6383 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6384 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6385 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6386 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6387 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6388 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n2 68.0561
R6389 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n23 49.8072
R6390 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n21 49.8072
R6391 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 41.7838
R6392 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6393 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t6 24.0005
R6394 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t5 24.0005
R6395 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 1.1255
R6396 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n1 1.11856
R6397 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R6398 bgr_0.V_mir1.n9 bgr_0.V_mir1.n5 325.471
R6399 bgr_0.V_mir1.n4 bgr_0.V_mir1.n0 325.471
R6400 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R6401 bgr_0.V_mir1.n6 bgr_0.V_mir1.t22 310.488
R6402 bgr_0.V_mir1.n1 bgr_0.V_mir1.t17 310.488
R6403 bgr_0.V_mir1.n12 bgr_0.V_mir1.t14 278.312
R6404 bgr_0.V_mir1.n12 bgr_0.V_mir1.n11 228.939
R6405 bgr_0.V_mir1.n13 bgr_0.V_mir1.n10 224.439
R6406 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R6407 bgr_0.V_mir1.n8 bgr_0.V_mir1.t2 184.097
R6408 bgr_0.V_mir1.n3 bgr_0.V_mir1.t4 184.097
R6409 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R6410 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 167.094
R6411 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 167.094
R6412 bgr_0.V_mir1.n9 bgr_0.V_mir1.n8 152
R6413 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 152
R6414 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R6415 bgr_0.V_mir1.n16 bgr_0.V_mir1.t21 120.501
R6416 bgr_0.V_mir1.n17 bgr_0.V_mir1.t12 120.501
R6417 bgr_0.V_mir1.n6 bgr_0.V_mir1.t20 120.501
R6418 bgr_0.V_mir1.n7 bgr_0.V_mir1.t6 120.501
R6419 bgr_0.V_mir1.n1 bgr_0.V_mir1.t18 120.501
R6420 bgr_0.V_mir1.n2 bgr_0.V_mir1.t8 120.501
R6421 bgr_0.V_mir1.n11 bgr_0.V_mir1.t16 48.0005
R6422 bgr_0.V_mir1.n11 bgr_0.V_mir1.t0 48.0005
R6423 bgr_0.V_mir1.n10 bgr_0.V_mir1.t1 48.0005
R6424 bgr_0.V_mir1.n10 bgr_0.V_mir1.t15 48.0005
R6425 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R6426 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 40.7027
R6427 bgr_0.V_mir1.n3 bgr_0.V_mir1.n2 40.7027
R6428 bgr_0.V_mir1.n5 bgr_0.V_mir1.t7 39.4005
R6429 bgr_0.V_mir1.n5 bgr_0.V_mir1.t3 39.4005
R6430 bgr_0.V_mir1.n0 bgr_0.V_mir1.t9 39.4005
R6431 bgr_0.V_mir1.n0 bgr_0.V_mir1.t5 39.4005
R6432 bgr_0.V_mir1.t13 bgr_0.V_mir1.n20 39.4005
R6433 bgr_0.V_mir1.n20 bgr_0.V_mir1.t11 39.4005
R6434 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R6435 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R6436 bgr_0.V_mir1.n14 bgr_0.V_mir1.n9 9.3005
R6437 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 5.8755
R6438 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R6439 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 0.78175
R6440 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t26 1172.87
R6441 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t35 1172.87
R6442 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.t45 996.134
R6443 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t34 996.134
R6444 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t48 996.134
R6445 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t38 996.134
R6446 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t51 996.134
R6447 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t27 996.134
R6448 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t43 996.134
R6449 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t30 996.134
R6450 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t29 690.867
R6451 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t40 690.867
R6452 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t54 530.201
R6453 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t33 530.201
R6454 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t39 514.134
R6455 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t49 514.134
R6456 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t36 514.134
R6457 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t46 514.134
R6458 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t31 514.134
R6459 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 514.134
R6460 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t41 514.134
R6461 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t52 514.134
R6462 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6463 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.t50 353.467
R6464 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t25 353.467
R6465 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t42 353.467
R6466 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t28 353.467
R6467 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t44 353.467
R6468 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t32 353.467
R6469 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t47 353.467
R6470 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 176.733
R6471 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R6472 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R6473 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R6474 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R6475 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.n47 176.733
R6476 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 176.733
R6477 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 176.733
R6478 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 176.733
R6479 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R6480 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6481 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6482 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 176.733
R6483 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6484 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R6485 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6486 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6487 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6488 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 166.436
R6489 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n31 161.875
R6490 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n40 161.686
R6491 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n0 160.427
R6492 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 159.802
R6493 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 159.802
R6494 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 159.802
R6495 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n1 159.802
R6496 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 155.302
R6497 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n13 114.689
R6498 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n12 114.689
R6499 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 114.126
R6500 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 114.126
R6501 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 114.126
R6502 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n11 109.626
R6503 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 51.9494
R6504 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R6505 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 51.9494
R6506 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n23 51.9494
R6507 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R6508 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n32 51.9494
R6509 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.X.n52 49.3036
R6510 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t20 16.0005
R6511 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t24 16.0005
R6512 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t0 16.0005
R6513 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R6514 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t8 16.0005
R6515 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R6516 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R6517 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t19 16.0005
R6518 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t18 16.0005
R6519 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t7 16.0005
R6520 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t23 16.0005
R6521 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R6522 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n42 15.7193
R6523 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t13 11.2576
R6524 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R6525 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R6526 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t21 11.2576
R6527 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t22 11.2576
R6528 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t11 11.2576
R6529 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t12 11.2576
R6530 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t2 11.2576
R6531 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t10 11.2576
R6532 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R6533 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t9 11.2576
R6534 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t16 11.2576
R6535 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n22 10.188
R6536 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 6.188
R6537 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n8 5.1255
R6538 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n20 4.5005
R6539 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 0.6255
R6540 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.6255
R6541 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.6255
R6542 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n15 0.563
R6543 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n17 0.563
R6544 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 0.563
R6545 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n10 0.5005
R6546 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 0.438
R6547 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 344.837
R6548 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 344.274
R6549 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 292.5
R6550 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 206.052
R6551 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 205.488
R6552 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 205.488
R6553 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 205.488
R6554 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 205.488
R6555 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 122.504
R6556 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 72.5626
R6557 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 52.3363
R6558 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R6559 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 39.4005
R6560 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R6561 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 39.4005
R6562 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R6563 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R6564 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 33.3443
R6565 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R6566 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R6567 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R6568 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R6569 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 19.7005
R6570 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R6571 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R6572 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R6573 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R6574 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R6575 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 6.09425
R6576 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 0.563
R6577 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 0.563
R6578 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 0.563
R6579 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t52 1172.87
R6580 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t27 1172.87
R6581 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t44 996.134
R6582 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6583 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t49 996.134
R6584 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t37 996.134
R6585 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R6586 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t36 996.134
R6587 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t42 996.134
R6588 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.t29 996.134
R6589 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t25 690.867
R6590 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t30 690.867
R6591 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t51 530.201
R6592 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t26 530.201
R6593 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t39 514.134
R6594 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t53 514.134
R6595 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t40 514.134
R6596 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R6597 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t38 514.134
R6598 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t50 514.134
R6599 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R6600 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 514.134
R6601 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t34 353.467
R6602 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R6603 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t28 353.467
R6604 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t43 353.467
R6605 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t31 353.467
R6606 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R6607 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t35 353.467
R6608 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t46 353.467
R6609 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R6610 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R6611 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R6612 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R6613 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R6614 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 176.733
R6615 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R6616 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6617 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6618 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6619 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R6620 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R6621 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R6622 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R6623 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R6624 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R6625 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R6626 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R6627 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 166.375
R6628 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.875
R6629 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.686
R6630 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n0 160.427
R6631 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n7 159.802
R6632 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 159.802
R6633 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 159.802
R6634 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n1 159.802
R6635 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 155.302
R6636 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 114.689
R6637 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n12 114.689
R6638 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 114.126
R6639 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n15 114.126
R6640 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 114.126
R6641 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n11 109.626
R6642 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R6643 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n42 51.9494
R6644 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R6645 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n28 51.9494
R6646 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R6647 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n37 51.9494
R6648 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t2 49.2412
R6649 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R6650 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t20 16.0005
R6651 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t3 16.0005
R6652 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t23 16.0005
R6653 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t13 16.0005
R6654 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t8 16.0005
R6655 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t17 16.0005
R6656 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R6657 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t19 16.0005
R6658 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t16 16.0005
R6659 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R6660 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t21 16.0005
R6661 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 15.6567
R6662 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t22 11.2576
R6663 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t18 11.2576
R6664 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t5 11.2576
R6665 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t1 11.2576
R6666 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t7 11.2576
R6667 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t0 11.2576
R6668 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t9 11.2576
R6669 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t12 11.2576
R6670 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t14 11.2576
R6671 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t10 11.2576
R6672 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t24 11.2576
R6673 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t4 11.2576
R6674 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n51 10.313
R6675 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n40 6.063
R6676 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n8 5.1255
R6677 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 4.5005
R6678 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n2 0.6255
R6679 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n4 0.6255
R6680 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n6 0.6255
R6681 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n14 0.563
R6682 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n16 0.563
R6683 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n18 0.563
R6684 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n10 0.5005
R6685 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n21 0.438
R6686 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 144.827
R6687 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 134.577
R6688 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 120.629
R6689 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 101.376
R6690 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 97.4009
R6691 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 96.8384
R6692 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 96.8384
R6693 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 96.8384
R6694 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 96.8384
R6695 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 24.0005
R6696 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 24.0005
R6697 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 24.0005
R6698 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R6699 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R6700 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 8.0005
R6701 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R6702 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 8.0005
R6703 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R6704 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 8.0005
R6705 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R6706 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 8.0005
R6707 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R6708 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R6709 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 5.84425
R6710 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 1.46925
R6711 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 0.563
R6712 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 0.563
R6713 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.563
R6714 bgr_0.V_p_2.n1 bgr_0.V_p_2.n4 229.562
R6715 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R6716 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R6717 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 228.939
R6718 bgr_0.V_p_2.n6 bgr_0.V_p_2.n0 228.938
R6719 bgr_0.V_p_2.n0 bgr_0.V_p_2.t0 98.2282
R6720 bgr_0.V_p_2.n5 bgr_0.V_p_2.t5 48.0005
R6721 bgr_0.V_p_2.n5 bgr_0.V_p_2.t8 48.0005
R6722 bgr_0.V_p_2.n4 bgr_0.V_p_2.t1 48.0005
R6723 bgr_0.V_p_2.n4 bgr_0.V_p_2.t3 48.0005
R6724 bgr_0.V_p_2.n3 bgr_0.V_p_2.t2 48.0005
R6725 bgr_0.V_p_2.n3 bgr_0.V_p_2.t9 48.0005
R6726 bgr_0.V_p_2.n2 bgr_0.V_p_2.t10 48.0005
R6727 bgr_0.V_p_2.n2 bgr_0.V_p_2.t4 48.0005
R6728 bgr_0.V_p_2.n6 bgr_0.V_p_2.t7 48.0005
R6729 bgr_0.V_p_2.t6 bgr_0.V_p_2.n6 48.0005
R6730 bgr_0.V_p_2.n0 bgr_0.V_p_2.n1 1.8755
R6731 VOUT+.n2 VOUT+.n0 145.989
R6732 VOUT+.n8 VOUT+.n7 145.989
R6733 VOUT+.n6 VOUT+.n5 145.427
R6734 VOUT+.n4 VOUT+.n3 145.427
R6735 VOUT+.n2 VOUT+.n1 145.427
R6736 VOUT+.n10 VOUT+.n9 140.927
R6737 VOUT+.n100 VOUT+.t3 113.192
R6738 VOUT+.n97 VOUT+.n95 95.7303
R6739 VOUT+.n99 VOUT+.n98 94.6053
R6740 VOUT+.n97 VOUT+.n96 94.6053
R6741 VOUT+.n94 VOUT+.n10 20.5943
R6742 VOUT+.n94 VOUT+.n93 11.7059
R6743 VOUT+ VOUT+.n94 7.813
R6744 VOUT+.n9 VOUT+.t8 6.56717
R6745 VOUT+.n9 VOUT+.t12 6.56717
R6746 VOUT+.n7 VOUT+.t6 6.56717
R6747 VOUT+.n7 VOUT+.t1 6.56717
R6748 VOUT+.n5 VOUT+.t7 6.56717
R6749 VOUT+.n5 VOUT+.t11 6.56717
R6750 VOUT+.n3 VOUT+.t9 6.56717
R6751 VOUT+.n3 VOUT+.t13 6.56717
R6752 VOUT+.n1 VOUT+.t10 6.56717
R6753 VOUT+.n1 VOUT+.t14 6.56717
R6754 VOUT+.n0 VOUT+.t0 6.56717
R6755 VOUT+.n0 VOUT+.t15 6.56717
R6756 VOUT+.n40 VOUT+.t108 4.8295
R6757 VOUT+.n52 VOUT+.t25 4.8295
R6758 VOUT+.n49 VOUT+.t76 4.8295
R6759 VOUT+.n46 VOUT+.t113 4.8295
R6760 VOUT+.n43 VOUT+.t145 4.8295
R6761 VOUT+.n42 VOUT+.t68 4.8295
R6762 VOUT+.n66 VOUT+.t28 4.8295
R6763 VOUT+.n67 VOUT+.t77 4.8295
R6764 VOUT+.n69 VOUT+.t63 4.8295
R6765 VOUT+.n70 VOUT+.t111 4.8295
R6766 VOUT+.n72 VOUT+.t114 4.8295
R6767 VOUT+.n73 VOUT+.t99 4.8295
R6768 VOUT+.n75 VOUT+.t74 4.8295
R6769 VOUT+.n76 VOUT+.t56 4.8295
R6770 VOUT+.n78 VOUT+.t109 4.8295
R6771 VOUT+.n79 VOUT+.t92 4.8295
R6772 VOUT+.n81 VOUT+.t69 4.8295
R6773 VOUT+.n82 VOUT+.t53 4.8295
R6774 VOUT+.n84 VOUT+.t30 4.8295
R6775 VOUT+.n85 VOUT+.t153 4.8295
R6776 VOUT+.n87 VOUT+.t64 4.8295
R6777 VOUT+.n88 VOUT+.t47 4.8295
R6778 VOUT+.n11 VOUT+.t117 4.8295
R6779 VOUT+.n13 VOUT+.t72 4.8295
R6780 VOUT+.n25 VOUT+.t38 4.8295
R6781 VOUT+.n26 VOUT+.t20 4.8295
R6782 VOUT+.n28 VOUT+.t80 4.8295
R6783 VOUT+.n29 VOUT+.t61 4.8295
R6784 VOUT+.n31 VOUT+.t121 4.8295
R6785 VOUT+.n32 VOUT+.t104 4.8295
R6786 VOUT+.n34 VOUT+.t85 4.8295
R6787 VOUT+.n35 VOUT+.t67 4.8295
R6788 VOUT+.n37 VOUT+.t123 4.8295
R6789 VOUT+.n38 VOUT+.t107 4.8295
R6790 VOUT+.n90 VOUT+.t22 4.8295
R6791 VOUT+.n55 VOUT+.t33 4.806
R6792 VOUT+.n56 VOUT+.t150 4.806
R6793 VOUT+.n57 VOUT+.t51 4.806
R6794 VOUT+.n58 VOUT+.t88 4.806
R6795 VOUT+.n59 VOUT+.t125 4.806
R6796 VOUT+.n60 VOUT+.t105 4.806
R6797 VOUT+.n61 VOUT+.t140 4.806
R6798 VOUT+.n62 VOUT+.t37 4.806
R6799 VOUT+.n63 VOUT+.t156 4.806
R6800 VOUT+.n64 VOUT+.t54 4.806
R6801 VOUT+.n14 VOUT+.t73 4.806
R6802 VOUT+.n15 VOUT+.t116 4.806
R6803 VOUT+.n16 VOUT+.t65 4.806
R6804 VOUT+.n17 VOUT+.t154 4.806
R6805 VOUT+.n18 VOUT+.t106 4.806
R6806 VOUT+.n19 VOUT+.t143 4.806
R6807 VOUT+.n20 VOUT+.t96 4.806
R6808 VOUT+.n21 VOUT+.t43 4.806
R6809 VOUT+.n22 VOUT+.t87 4.806
R6810 VOUT+.n23 VOUT+.t35 4.806
R6811 VOUT+.n40 VOUT+.t70 4.5005
R6812 VOUT+.n41 VOUT+.t91 4.5005
R6813 VOUT+.n52 VOUT+.t66 4.5005
R6814 VOUT+.n53 VOUT+.t81 4.5005
R6815 VOUT+.n54 VOUT+.t44 4.5005
R6816 VOUT+.n49 VOUT+.t118 4.5005
R6817 VOUT+.n50 VOUT+.t57 4.5005
R6818 VOUT+.n51 VOUT+.t21 4.5005
R6819 VOUT+.n46 VOUT+.t151 4.5005
R6820 VOUT+.n47 VOUT+.t98 4.5005
R6821 VOUT+.n48 VOUT+.t60 4.5005
R6822 VOUT+.n43 VOUT+.t45 4.5005
R6823 VOUT+.n44 VOUT+.t136 4.5005
R6824 VOUT+.n45 VOUT+.t101 4.5005
R6825 VOUT+.n42 VOUT+.t31 4.5005
R6826 VOUT+.n65 VOUT+.t52 4.5005
R6827 VOUT+.n64 VOUT+.t155 4.5005
R6828 VOUT+.n63 VOUT+.t119 4.5005
R6829 VOUT+.n62 VOUT+.t139 4.5005
R6830 VOUT+.n61 VOUT+.t102 4.5005
R6831 VOUT+.n60 VOUT+.t62 4.5005
R6832 VOUT+.n59 VOUT+.t86 4.5005
R6833 VOUT+.n58 VOUT+.t46 4.5005
R6834 VOUT+.n57 VOUT+.t147 4.5005
R6835 VOUT+.n56 VOUT+.t110 4.5005
R6836 VOUT+.n55 VOUT+.t134 4.5005
R6837 VOUT+.n66 VOUT+.t130 4.5005
R6838 VOUT+.n68 VOUT+.t152 4.5005
R6839 VOUT+.n67 VOUT+.t115 4.5005
R6840 VOUT+.n69 VOUT+.t23 4.5005
R6841 VOUT+.n71 VOUT+.t48 4.5005
R6842 VOUT+.n70 VOUT+.t148 4.5005
R6843 VOUT+.n72 VOUT+.t79 4.5005
R6844 VOUT+.n74 VOUT+.t27 4.5005
R6845 VOUT+.n73 VOUT+.t132 4.5005
R6846 VOUT+.n75 VOUT+.t40 4.5005
R6847 VOUT+.n77 VOUT+.t128 4.5005
R6848 VOUT+.n76 VOUT+.t93 4.5005
R6849 VOUT+.n78 VOUT+.t71 4.5005
R6850 VOUT+.n80 VOUT+.t19 4.5005
R6851 VOUT+.n79 VOUT+.t126 4.5005
R6852 VOUT+.n81 VOUT+.t34 4.5005
R6853 VOUT+.n83 VOUT+.t122 4.5005
R6854 VOUT+.n82 VOUT+.t89 4.5005
R6855 VOUT+.n84 VOUT+.t135 4.5005
R6856 VOUT+.n86 VOUT+.t83 4.5005
R6857 VOUT+.n85 VOUT+.t49 4.5005
R6858 VOUT+.n87 VOUT+.t29 4.5005
R6859 VOUT+.n89 VOUT+.t120 4.5005
R6860 VOUT+.n88 VOUT+.t82 4.5005
R6861 VOUT+.n11 VOUT+.t26 4.5005
R6862 VOUT+.n12 VOUT+.t124 4.5005
R6863 VOUT+.n13 VOUT+.t39 4.5005
R6864 VOUT+.n24 VOUT+.t127 4.5005
R6865 VOUT+.n23 VOUT+.t95 4.5005
R6866 VOUT+.n22 VOUT+.t55 4.5005
R6867 VOUT+.n21 VOUT+.t144 4.5005
R6868 VOUT+.n20 VOUT+.t112 4.5005
R6869 VOUT+.n19 VOUT+.t75 4.5005
R6870 VOUT+.n18 VOUT+.t24 4.5005
R6871 VOUT+.n17 VOUT+.t131 4.5005
R6872 VOUT+.n16 VOUT+.t97 4.5005
R6873 VOUT+.n15 VOUT+.t59 4.5005
R6874 VOUT+.n14 VOUT+.t149 4.5005
R6875 VOUT+.n25 VOUT+.t142 4.5005
R6876 VOUT+.n27 VOUT+.t94 4.5005
R6877 VOUT+.n26 VOUT+.t58 4.5005
R6878 VOUT+.n28 VOUT+.t42 4.5005
R6879 VOUT+.n30 VOUT+.t133 4.5005
R6880 VOUT+.n29 VOUT+.t100 4.5005
R6881 VOUT+.n31 VOUT+.t84 4.5005
R6882 VOUT+.n33 VOUT+.t32 4.5005
R6883 VOUT+.n32 VOUT+.t137 4.5005
R6884 VOUT+.n34 VOUT+.t50 4.5005
R6885 VOUT+.n36 VOUT+.t138 4.5005
R6886 VOUT+.n35 VOUT+.t103 4.5005
R6887 VOUT+.n37 VOUT+.t90 4.5005
R6888 VOUT+.n39 VOUT+.t36 4.5005
R6889 VOUT+.n38 VOUT+.t141 4.5005
R6890 VOUT+.n90 VOUT+.t129 4.5005
R6891 VOUT+.n91 VOUT+.t78 4.5005
R6892 VOUT+.n92 VOUT+.t41 4.5005
R6893 VOUT+.n93 VOUT+.t146 4.5005
R6894 VOUT+.n10 VOUT+.n8 4.5005
R6895 VOUT+.n98 VOUT+.t17 3.42907
R6896 VOUT+.n98 VOUT+.t5 3.42907
R6897 VOUT+.n96 VOUT+.t18 3.42907
R6898 VOUT+.n96 VOUT+.t4 3.42907
R6899 VOUT+.n95 VOUT+.t2 3.42907
R6900 VOUT+.n95 VOUT+.t16 3.42907
R6901 VOUT+ VOUT+.n100 2.84425
R6902 VOUT+.n100 VOUT+.n99 2.03175
R6903 VOUT+.n99 VOUT+.n97 1.1255
R6904 VOUT+.n4 VOUT+.n2 0.563
R6905 VOUT+.n6 VOUT+.n4 0.563
R6906 VOUT+.n8 VOUT+.n6 0.563
R6907 VOUT+.n41 VOUT+.n40 0.3295
R6908 VOUT+.n54 VOUT+.n53 0.3295
R6909 VOUT+.n53 VOUT+.n52 0.3295
R6910 VOUT+.n51 VOUT+.n50 0.3295
R6911 VOUT+.n50 VOUT+.n49 0.3295
R6912 VOUT+.n48 VOUT+.n47 0.3295
R6913 VOUT+.n47 VOUT+.n46 0.3295
R6914 VOUT+.n45 VOUT+.n44 0.3295
R6915 VOUT+.n44 VOUT+.n43 0.3295
R6916 VOUT+.n65 VOUT+.n42 0.3295
R6917 VOUT+.n65 VOUT+.n64 0.3295
R6918 VOUT+.n64 VOUT+.n63 0.3295
R6919 VOUT+.n63 VOUT+.n62 0.3295
R6920 VOUT+.n62 VOUT+.n61 0.3295
R6921 VOUT+.n61 VOUT+.n60 0.3295
R6922 VOUT+.n60 VOUT+.n59 0.3295
R6923 VOUT+.n59 VOUT+.n58 0.3295
R6924 VOUT+.n58 VOUT+.n57 0.3295
R6925 VOUT+.n57 VOUT+.n56 0.3295
R6926 VOUT+.n56 VOUT+.n55 0.3295
R6927 VOUT+.n68 VOUT+.n66 0.3295
R6928 VOUT+.n68 VOUT+.n67 0.3295
R6929 VOUT+.n71 VOUT+.n69 0.3295
R6930 VOUT+.n71 VOUT+.n70 0.3295
R6931 VOUT+.n74 VOUT+.n72 0.3295
R6932 VOUT+.n74 VOUT+.n73 0.3295
R6933 VOUT+.n77 VOUT+.n75 0.3295
R6934 VOUT+.n77 VOUT+.n76 0.3295
R6935 VOUT+.n80 VOUT+.n78 0.3295
R6936 VOUT+.n80 VOUT+.n79 0.3295
R6937 VOUT+.n83 VOUT+.n81 0.3295
R6938 VOUT+.n83 VOUT+.n82 0.3295
R6939 VOUT+.n86 VOUT+.n84 0.3295
R6940 VOUT+.n86 VOUT+.n85 0.3295
R6941 VOUT+.n89 VOUT+.n87 0.3295
R6942 VOUT+.n89 VOUT+.n88 0.3295
R6943 VOUT+.n12 VOUT+.n11 0.3295
R6944 VOUT+.n24 VOUT+.n13 0.3295
R6945 VOUT+.n24 VOUT+.n23 0.3295
R6946 VOUT+.n23 VOUT+.n22 0.3295
R6947 VOUT+.n22 VOUT+.n21 0.3295
R6948 VOUT+.n21 VOUT+.n20 0.3295
R6949 VOUT+.n20 VOUT+.n19 0.3295
R6950 VOUT+.n19 VOUT+.n18 0.3295
R6951 VOUT+.n18 VOUT+.n17 0.3295
R6952 VOUT+.n17 VOUT+.n16 0.3295
R6953 VOUT+.n16 VOUT+.n15 0.3295
R6954 VOUT+.n15 VOUT+.n14 0.3295
R6955 VOUT+.n27 VOUT+.n25 0.3295
R6956 VOUT+.n27 VOUT+.n26 0.3295
R6957 VOUT+.n30 VOUT+.n28 0.3295
R6958 VOUT+.n30 VOUT+.n29 0.3295
R6959 VOUT+.n33 VOUT+.n31 0.3295
R6960 VOUT+.n33 VOUT+.n32 0.3295
R6961 VOUT+.n36 VOUT+.n34 0.3295
R6962 VOUT+.n36 VOUT+.n35 0.3295
R6963 VOUT+.n39 VOUT+.n37 0.3295
R6964 VOUT+.n39 VOUT+.n38 0.3295
R6965 VOUT+.n91 VOUT+.n90 0.3295
R6966 VOUT+.n92 VOUT+.n91 0.3295
R6967 VOUT+.n93 VOUT+.n92 0.3295
R6968 VOUT+.n59 VOUT+.n54 0.306
R6969 VOUT+.n60 VOUT+.n51 0.306
R6970 VOUT+.n61 VOUT+.n48 0.306
R6971 VOUT+.n62 VOUT+.n45 0.306
R6972 VOUT+.n65 VOUT+.n41 0.2825
R6973 VOUT+.n68 VOUT+.n65 0.2825
R6974 VOUT+.n71 VOUT+.n68 0.2825
R6975 VOUT+.n74 VOUT+.n71 0.2825
R6976 VOUT+.n77 VOUT+.n74 0.2825
R6977 VOUT+.n80 VOUT+.n77 0.2825
R6978 VOUT+.n83 VOUT+.n80 0.2825
R6979 VOUT+.n86 VOUT+.n83 0.2825
R6980 VOUT+.n89 VOUT+.n86 0.2825
R6981 VOUT+.n24 VOUT+.n12 0.2825
R6982 VOUT+.n27 VOUT+.n24 0.2825
R6983 VOUT+.n30 VOUT+.n27 0.2825
R6984 VOUT+.n33 VOUT+.n30 0.2825
R6985 VOUT+.n36 VOUT+.n33 0.2825
R6986 VOUT+.n39 VOUT+.n36 0.2825
R6987 VOUT+.n91 VOUT+.n39 0.2825
R6988 VOUT+.n91 VOUT+.n89 0.2825
R6989 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 49.2006
R6990 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.1603
R6991 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R6992 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R6993 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R6994 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.1603
R6995 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R6996 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1603
R6997 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R6998 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R6999 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R7000 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R7001 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1603
R7002 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.1603
R7003 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.1603
R7004 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1603
R7005 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1603
R7006 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R7007 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R7008 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1603
R7009 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R7010 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1603
R7011 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R7012 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1603
R7013 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1603
R7014 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.1603
R7015 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R7016 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1603
R7017 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R7018 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R7019 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1603
R7020 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R7021 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1603
R7022 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1603
R7023 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1603
R7024 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.1603
R7025 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1603
R7026 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R7027 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1603
R7028 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R7029 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1603
R7030 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R7031 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1603
R7032 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1603
R7033 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R7034 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.1603
R7035 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1603
R7036 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.1603
R7037 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1603
R7038 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1603
R7039 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R7040 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R7041 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.1603
R7042 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1603
R7043 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1603
R7044 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R7045 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R7046 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.1603
R7047 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1603
R7048 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.159278
R7049 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.159278
R7050 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.159278
R7051 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.159278
R7052 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.159278
R7053 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.159278
R7054 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.159278
R7055 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.159278
R7056 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.159278
R7057 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.159278
R7058 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.159278
R7059 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.159278
R7060 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.159278
R7061 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R7062 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R7063 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R7064 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7065 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7066 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7067 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7068 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7069 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7070 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7071 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.159278
R7072 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.159278
R7073 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.159278
R7074 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.159278
R7075 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.137822
R7076 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1368
R7077 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1368
R7078 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1368
R7079 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1368
R7080 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1368
R7081 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.1368
R7082 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1368
R7083 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.1368
R7084 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7085 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1368
R7086 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1368
R7087 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1368
R7088 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1368
R7089 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1368
R7090 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.1368
R7091 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1368
R7092 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1368
R7093 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1368
R7094 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.1368
R7095 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.1368
R7096 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.1368
R7097 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.1368
R7098 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.1368
R7099 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1368
R7100 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1368
R7101 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R7102 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1368
R7103 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1368
R7104 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R7105 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R7106 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1368
R7107 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.114322
R7108 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.1133
R7109 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.1133
R7110 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7111 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7112 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7113 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7114 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7115 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7116 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7117 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7118 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7119 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7120 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7121 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7122 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.1133
R7123 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.1133
R7124 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.1133
R7125 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.1133
R7126 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R7127 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.00152174
R7128 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.00152174
R7129 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.00152174
R7130 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.00152174
R7131 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.00152174
R7132 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.00152174
R7133 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.00152174
R7134 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R7135 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.00152174
R7136 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.00152174
R7137 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.00152174
R7138 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.00152174
R7139 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.00152174
R7140 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.00152174
R7141 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.00152174
R7142 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.00152174
R7143 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.00152174
R7144 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.00152174
R7145 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.00152174
R7146 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.00152174
R7147 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R7148 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.00152174
R7149 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.00152174
R7150 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R7151 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.00152174
R7152 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.00152174
R7153 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.00152174
R7154 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R7155 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.00152174
R7156 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.00152174
R7157 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.00152174
R7158 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.00152174
R7159 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.00152174
R7160 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R7161 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R7162 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R7163 bgr_0.Vbe2.n102 bgr_0.Vbe2.t0 162.458
R7164 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 83.5719
R7165 bgr_0.Vbe2.n115 bgr_0.Vbe2.n9 83.5719
R7166 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 83.5719
R7167 bgr_0.Vbe2.n105 bgr_0.Vbe2.n12 83.5719
R7168 bgr_0.Vbe2.n97 bgr_0.Vbe2.n13 83.5719
R7169 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 83.5719
R7170 bgr_0.Vbe2.n91 bgr_0.Vbe2.n17 83.5719
R7171 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 83.5719
R7172 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 83.5719
R7173 bgr_0.Vbe2.n77 bgr_0.Vbe2.n76 83.5719
R7174 bgr_0.Vbe2.n38 bgr_0.Vbe2.n37 83.5719
R7175 bgr_0.Vbe2.n36 bgr_0.Vbe2.n34 83.5719
R7176 bgr_0.Vbe2.n44 bgr_0.Vbe2.n33 83.5719
R7177 bgr_0.Vbe2.n52 bgr_0.Vbe2.n51 83.5719
R7178 bgr_0.Vbe2.n31 bgr_0.Vbe2.n29 83.5719
R7179 bgr_0.Vbe2.n57 bgr_0.Vbe2.n28 83.5719
R7180 bgr_0.Vbe2.n65 bgr_0.Vbe2.n64 83.5719
R7181 bgr_0.Vbe2.n130 bgr_0.Vbe2.n0 83.5719
R7182 bgr_0.Vbe2.n132 bgr_0.Vbe2.n131 83.5719
R7183 bgr_0.Vbe2.n134 bgr_0.Vbe2.n133 83.5719
R7184 bgr_0.Vbe2.n116 bgr_0.Vbe2.n8 73.682
R7185 bgr_0.Vbe2.n37 bgr_0.Vbe2.n35 73.682
R7186 bgr_0.Vbe2.n114 bgr_0.Vbe2.n10 73.3165
R7187 bgr_0.Vbe2.n98 bgr_0.Vbe2.n96 73.3165
R7188 bgr_0.Vbe2.n77 bgr_0.Vbe2.n24 73.3165
R7189 bgr_0.Vbe2.n46 bgr_0.Vbe2.n33 73.3165
R7190 bgr_0.Vbe2.n59 bgr_0.Vbe2.n28 73.3165
R7191 bgr_0.Vbe2.n135 bgr_0.Vbe2.n134 73.3165
R7192 bgr_0.Vbe2.n107 bgr_0.Vbe2.n12 73.19
R7193 bgr_0.Vbe2.n93 bgr_0.Vbe2.n17 73.19
R7194 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 73.19
R7195 bgr_0.Vbe2.n51 bgr_0.Vbe2.n50 73.19
R7196 bgr_0.Vbe2.n64 bgr_0.Vbe2.n63 73.19
R7197 bgr_0.Vbe2.n130 bgr_0.Vbe2.n4 73.19
R7198 bgr_0.Vbe2.n18 bgr_0.Vbe2.t3 36.6632
R7199 bgr_0.Vbe2.t6 bgr_0.Vbe2.n25 36.6632
R7200 bgr_0.Vbe2.n115 bgr_0.Vbe2.n114 26.074
R7201 bgr_0.Vbe2.n98 bgr_0.Vbe2.n97 26.074
R7202 bgr_0.Vbe2.n79 bgr_0.Vbe2.n77 26.074
R7203 bgr_0.Vbe2.n36 bgr_0.Vbe2.n33 26.074
R7204 bgr_0.Vbe2.n31 bgr_0.Vbe2.n28 26.074
R7205 bgr_0.Vbe2.n134 bgr_0.Vbe2.n132 26.074
R7206 bgr_0.Vbe2.n116 bgr_0.Vbe2.t7 25.7843
R7207 bgr_0.Vbe2.t2 bgr_0.Vbe2.n12 25.7843
R7208 bgr_0.Vbe2.t3 bgr_0.Vbe2.n17 25.7843
R7209 bgr_0.Vbe2.n81 bgr_0.Vbe2.t4 25.7843
R7210 bgr_0.Vbe2.n37 bgr_0.Vbe2.t1 25.7843
R7211 bgr_0.Vbe2.n51 bgr_0.Vbe2.t5 25.7843
R7212 bgr_0.Vbe2.n64 bgr_0.Vbe2.t6 25.7843
R7213 bgr_0.Vbe2.t8 bgr_0.Vbe2.n130 25.7843
R7214 bgr_0.Vbe2.n138 bgr_0.Vbe2.n3 9.3005
R7215 bgr_0.Vbe2.n124 bgr_0.Vbe2.n3 9.3005
R7216 bgr_0.Vbe2.n129 bgr_0.Vbe2.n3 9.3005
R7217 bgr_0.Vbe2.n136 bgr_0.Vbe2.n3 9.3005
R7218 bgr_0.Vbe2.n138 bgr_0.Vbe2.n5 9.3005
R7219 bgr_0.Vbe2.n124 bgr_0.Vbe2.n5 9.3005
R7220 bgr_0.Vbe2.n129 bgr_0.Vbe2.n5 9.3005
R7221 bgr_0.Vbe2.n136 bgr_0.Vbe2.n5 9.3005
R7222 bgr_0.Vbe2.n138 bgr_0.Vbe2.n2 9.3005
R7223 bgr_0.Vbe2.n124 bgr_0.Vbe2.n2 9.3005
R7224 bgr_0.Vbe2.n129 bgr_0.Vbe2.n2 9.3005
R7225 bgr_0.Vbe2.n136 bgr_0.Vbe2.n2 9.3005
R7226 bgr_0.Vbe2.n138 bgr_0.Vbe2.n6 9.3005
R7227 bgr_0.Vbe2.n124 bgr_0.Vbe2.n6 9.3005
R7228 bgr_0.Vbe2.n129 bgr_0.Vbe2.n6 9.3005
R7229 bgr_0.Vbe2.n136 bgr_0.Vbe2.n6 9.3005
R7230 bgr_0.Vbe2.n138 bgr_0.Vbe2.n1 9.3005
R7231 bgr_0.Vbe2.n124 bgr_0.Vbe2.n1 9.3005
R7232 bgr_0.Vbe2.n129 bgr_0.Vbe2.n1 9.3005
R7233 bgr_0.Vbe2.n123 bgr_0.Vbe2.n1 9.3005
R7234 bgr_0.Vbe2.n136 bgr_0.Vbe2.n1 9.3005
R7235 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 9.3005
R7236 bgr_0.Vbe2.n137 bgr_0.Vbe2.n124 9.3005
R7237 bgr_0.Vbe2.n137 bgr_0.Vbe2.n129 9.3005
R7238 bgr_0.Vbe2.n137 bgr_0.Vbe2.n123 9.3005
R7239 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 9.3005
R7240 bgr_0.Vbe2.n71 bgr_0.Vbe2.n22 9.3005
R7241 bgr_0.Vbe2.n71 bgr_0.Vbe2.n20 9.3005
R7242 bgr_0.Vbe2.n71 bgr_0.Vbe2.n23 9.3005
R7243 bgr_0.Vbe2.n86 bgr_0.Vbe2.n71 9.3005
R7244 bgr_0.Vbe2.n73 bgr_0.Vbe2.n22 9.3005
R7245 bgr_0.Vbe2.n73 bgr_0.Vbe2.n20 9.3005
R7246 bgr_0.Vbe2.n73 bgr_0.Vbe2.n23 9.3005
R7247 bgr_0.Vbe2.n86 bgr_0.Vbe2.n73 9.3005
R7248 bgr_0.Vbe2.n70 bgr_0.Vbe2.n22 9.3005
R7249 bgr_0.Vbe2.n70 bgr_0.Vbe2.n20 9.3005
R7250 bgr_0.Vbe2.n70 bgr_0.Vbe2.n23 9.3005
R7251 bgr_0.Vbe2.n86 bgr_0.Vbe2.n70 9.3005
R7252 bgr_0.Vbe2.n85 bgr_0.Vbe2.n22 9.3005
R7253 bgr_0.Vbe2.n85 bgr_0.Vbe2.n20 9.3005
R7254 bgr_0.Vbe2.n85 bgr_0.Vbe2.n23 9.3005
R7255 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 9.3005
R7256 bgr_0.Vbe2.n69 bgr_0.Vbe2.n22 9.3005
R7257 bgr_0.Vbe2.n69 bgr_0.Vbe2.n20 9.3005
R7258 bgr_0.Vbe2.n69 bgr_0.Vbe2.n23 9.3005
R7259 bgr_0.Vbe2.n69 bgr_0.Vbe2.n19 9.3005
R7260 bgr_0.Vbe2.n86 bgr_0.Vbe2.n69 9.3005
R7261 bgr_0.Vbe2.n87 bgr_0.Vbe2.n22 9.3005
R7262 bgr_0.Vbe2.n87 bgr_0.Vbe2.n20 9.3005
R7263 bgr_0.Vbe2.n87 bgr_0.Vbe2.n23 9.3005
R7264 bgr_0.Vbe2.n87 bgr_0.Vbe2.n19 9.3005
R7265 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 9.3005
R7266 bgr_0.Vbe2.n123 bgr_0.Vbe2.n121 4.64654
R7267 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 4.64654
R7268 bgr_0.Vbe2.n123 bgr_0.Vbe2.n122 4.64654
R7269 bgr_0.Vbe2.n127 bgr_0.Vbe2.n125 4.64654
R7270 bgr_0.Vbe2.n128 bgr_0.Vbe2.n127 4.64654
R7271 bgr_0.Vbe2.n72 bgr_0.Vbe2.n19 4.64654
R7272 bgr_0.Vbe2.n83 bgr_0.Vbe2.n75 4.64654
R7273 bgr_0.Vbe2.n74 bgr_0.Vbe2.n19 4.64654
R7274 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 4.64654
R7275 bgr_0.Vbe2.n83 bgr_0.Vbe2.n21 4.64654
R7276 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 2.36206
R7277 bgr_0.Vbe2.n94 bgr_0.Vbe2.n93 2.36206
R7278 bgr_0.Vbe2.n50 bgr_0.Vbe2.n48 2.36206
R7279 bgr_0.Vbe2.n63 bgr_0.Vbe2.n61 2.36206
R7280 bgr_0.Vbe2.n109 bgr_0.Vbe2.n10 2.19742
R7281 bgr_0.Vbe2.n96 bgr_0.Vbe2.n95 2.19742
R7282 bgr_0.Vbe2.n47 bgr_0.Vbe2.n46 2.19742
R7283 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 2.19742
R7284 bgr_0.Vbe2.n90 bgr_0.Vbe2.n18 1.80777
R7285 bgr_0.Vbe2.n66 bgr_0.Vbe2.n25 1.80777
R7286 bgr_0.Vbe2.n62 bgr_0.Vbe2.n26 1.5505
R7287 bgr_0.Vbe2.n67 bgr_0.Vbe2.n66 1.5505
R7288 bgr_0.Vbe2.n49 bgr_0.Vbe2.n30 1.5505
R7289 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 1.5505
R7290 bgr_0.Vbe2.n56 bgr_0.Vbe2.n55 1.5505
R7291 bgr_0.Vbe2.n58 bgr_0.Vbe2.n27 1.5505
R7292 bgr_0.Vbe2.n40 bgr_0.Vbe2.n39 1.5505
R7293 bgr_0.Vbe2.n43 bgr_0.Vbe2.n42 1.5505
R7294 bgr_0.Vbe2.n45 bgr_0.Vbe2.n32 1.5505
R7295 bgr_0.Vbe2.n92 bgr_0.Vbe2.n16 1.5505
R7296 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 1.5505
R7297 bgr_0.Vbe2.n106 bgr_0.Vbe2.n11 1.5505
R7298 bgr_0.Vbe2.n104 bgr_0.Vbe2.n103 1.5505
R7299 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 1.5505
R7300 bgr_0.Vbe2.n15 bgr_0.Vbe2.n14 1.5505
R7301 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 1.5505
R7302 bgr_0.Vbe2.n112 bgr_0.Vbe2.n7 1.5505
R7303 bgr_0.Vbe2.n111 bgr_0.Vbe2.n110 1.5505
R7304 bgr_0.Vbe2.n111 bgr_0.Vbe2.n10 1.19225
R7305 bgr_0.Vbe2.n96 bgr_0.Vbe2.n15 1.19225
R7306 bgr_0.Vbe2.n24 bgr_0.Vbe2.n19 1.19225
R7307 bgr_0.Vbe2.n46 bgr_0.Vbe2.n45 1.19225
R7308 bgr_0.Vbe2.n59 bgr_0.Vbe2.n58 1.19225
R7309 bgr_0.Vbe2.n135 bgr_0.Vbe2.n123 1.19225
R7310 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14.Emitter bgr_0.Vbe2.n8 1.07742
R7311 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12.Emitter bgr_0.Vbe2.n35 1.07742
R7312 bgr_0.Vbe2.n118 bgr_0.Vbe2.n9 1.07024
R7313 bgr_0.Vbe2.n104 bgr_0.Vbe2.n13 1.07024
R7314 bgr_0.Vbe2.n78 bgr_0.Vbe2.n20 1.07024
R7315 bgr_0.Vbe2.n39 bgr_0.Vbe2.n34 1.07024
R7316 bgr_0.Vbe2.n53 bgr_0.Vbe2.n29 1.07024
R7317 bgr_0.Vbe2.n131 bgr_0.Vbe2.n124 1.07024
R7318 bgr_0.Vbe2.n68 bgr_0.Vbe2.n25 1.04793
R7319 bgr_0.Vbe2.n88 bgr_0.Vbe2.n18 1.04793
R7320 bgr_0.Vbe2.n107 bgr_0.Vbe2.n106 1.0237
R7321 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 1.0237
R7322 bgr_0.Vbe2.n82 bgr_0.Vbe2.n22 1.0237
R7323 bgr_0.Vbe2.n50 bgr_0.Vbe2.n49 1.0237
R7324 bgr_0.Vbe2.n63 bgr_0.Vbe2.n62 1.0237
R7325 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 1.0237
R7326 bgr_0.Vbe2.n113 bgr_0.Vbe2.n111 0.959578
R7327 bgr_0.Vbe2.n99 bgr_0.Vbe2.n15 0.959578
R7328 bgr_0.Vbe2.n76 bgr_0.Vbe2.n19 0.959578
R7329 bgr_0.Vbe2.n45 bgr_0.Vbe2.n44 0.959578
R7330 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 0.959578
R7331 bgr_0.Vbe2.n133 bgr_0.Vbe2.n123 0.959578
R7332 bgr_0.Vbe2.n113 bgr_0.Vbe2.n112 0.885803
R7333 bgr_0.Vbe2.n100 bgr_0.Vbe2.n99 0.885803
R7334 bgr_0.Vbe2.n76 bgr_0.Vbe2.n23 0.885803
R7335 bgr_0.Vbe2.n44 bgr_0.Vbe2.n43 0.885803
R7336 bgr_0.Vbe2.n57 bgr_0.Vbe2.n56 0.885803
R7337 bgr_0.Vbe2.n133 bgr_0.Vbe2.n129 0.885803
R7338 bgr_0.Vbe2.n83 bgr_0.Vbe2.n82 0.812055
R7339 bgr_0.Vbe2.n127 bgr_0.Vbe2.n4 0.812055
R7340 bgr_0.Vbe2.n112 bgr_0.Vbe2.n9 0.77514
R7341 bgr_0.Vbe2.n100 bgr_0.Vbe2.n13 0.77514
R7342 bgr_0.Vbe2.n78 bgr_0.Vbe2.n23 0.77514
R7343 bgr_0.Vbe2.n43 bgr_0.Vbe2.n34 0.77514
R7344 bgr_0.Vbe2.n56 bgr_0.Vbe2.n29 0.77514
R7345 bgr_0.Vbe2.n131 bgr_0.Vbe2.n129 0.77514
R7346 bgr_0.Vbe2.n40 bgr_0.Vbe2.n35 0.763532
R7347 bgr_0.Vbe2.n119 bgr_0.Vbe2.n8 0.763532
R7348 bgr_0.Vbe2.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16.Emitter 0.756696
R7349 bgr_0.Vbe2.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11.Emitter 0.756696
R7350 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9.Emitter bgr_0.Vbe2.n22 0.756696
R7351 bgr_0.Vbe2.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15.Emitter 0.756696
R7352 bgr_0.Vbe2.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10.Emitter 0.756696
R7353 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13.Emitter bgr_0.Vbe2.n138 0.756696
R7354 bgr_0.Vbe2.n86 bgr_0.Vbe2.n24 0.647417
R7355 bgr_0.Vbe2.n136 bgr_0.Vbe2.n135 0.647417
R7356 bgr_0.Vbe2.n118 bgr_0.Vbe2.n117 0.590702
R7357 bgr_0.Vbe2.n105 bgr_0.Vbe2.n104 0.590702
R7358 bgr_0.Vbe2.n91 bgr_0.Vbe2.n90 0.590702
R7359 bgr_0.Vbe2.n80 bgr_0.Vbe2.n20 0.590702
R7360 bgr_0.Vbe2.n39 bgr_0.Vbe2.n38 0.590702
R7361 bgr_0.Vbe2.n53 bgr_0.Vbe2.n52 0.590702
R7362 bgr_0.Vbe2.n66 bgr_0.Vbe2.n65 0.590702
R7363 bgr_0.Vbe2.n124 bgr_0.Vbe2.n0 0.590702
R7364 bgr_0.Vbe2.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14.Emitter 0.498483
R7365 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16.Emitter bgr_0.Vbe2.n105 0.498483
R7366 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11.Emitter bgr_0.Vbe2.n91 0.498483
R7367 bgr_0.Vbe2.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9.Emitter 0.498483
R7368 bgr_0.Vbe2.n38 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12.Emitter 0.498483
R7369 bgr_0.Vbe2.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15.Emitter 0.498483
R7370 bgr_0.Vbe2.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10.Emitter 0.498483
R7371 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13.Emitter bgr_0.Vbe2.n0 0.498483
R7372 bgr_0.Vbe2.t7 bgr_0.Vbe2.n115 0.290206
R7373 bgr_0.Vbe2.n97 bgr_0.Vbe2.t2 0.290206
R7374 bgr_0.Vbe2.t4 bgr_0.Vbe2.n79 0.290206
R7375 bgr_0.Vbe2.t1 bgr_0.Vbe2.n36 0.290206
R7376 bgr_0.Vbe2.t5 bgr_0.Vbe2.n31 0.290206
R7377 bgr_0.Vbe2.n132 bgr_0.Vbe2.t8 0.290206
R7378 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 0.154071
R7379 bgr_0.Vbe2.n48 bgr_0.Vbe2.n47 0.154071
R7380 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.154071
R7381 bgr_0.Vbe2.n109 bgr_0.Vbe2.n108 0.154071
R7382 bgr_0.Vbe2.n137 bgr_0.Vbe2.n120 0.137464
R7383 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 0.137464
R7384 bgr_0.Vbe2.n41 bgr_0.Vbe2.n1 0.134964
R7385 bgr_0.Vbe2.n69 bgr_0.Vbe2.n68 0.134964
R7386 bgr_0.Vbe2.n67 bgr_0.Vbe2.n26 0.0183571
R7387 bgr_0.Vbe2.n61 bgr_0.Vbe2.n26 0.0183571
R7388 bgr_0.Vbe2.n60 bgr_0.Vbe2.n27 0.0183571
R7389 bgr_0.Vbe2.n55 bgr_0.Vbe2.n27 0.0183571
R7390 bgr_0.Vbe2.n55 bgr_0.Vbe2.n54 0.0183571
R7391 bgr_0.Vbe2.n54 bgr_0.Vbe2.n30 0.0183571
R7392 bgr_0.Vbe2.n48 bgr_0.Vbe2.n30 0.0183571
R7393 bgr_0.Vbe2.n47 bgr_0.Vbe2.n32 0.0183571
R7394 bgr_0.Vbe2.n42 bgr_0.Vbe2.n32 0.0183571
R7395 bgr_0.Vbe2.n89 bgr_0.Vbe2.n16 0.0183571
R7396 bgr_0.Vbe2.n94 bgr_0.Vbe2.n16 0.0183571
R7397 bgr_0.Vbe2.n95 bgr_0.Vbe2.n14 0.0183571
R7398 bgr_0.Vbe2.n101 bgr_0.Vbe2.n14 0.0183571
R7399 bgr_0.Vbe2.n103 bgr_0.Vbe2.n11 0.0183571
R7400 bgr_0.Vbe2.n108 bgr_0.Vbe2.n11 0.0183571
R7401 bgr_0.Vbe2.n110 bgr_0.Vbe2.n109 0.0183571
R7402 bgr_0.Vbe2.n110 bgr_0.Vbe2.n7 0.0183571
R7403 bgr_0.Vbe2.n68 bgr_0.Vbe2.n67 0.0106786
R7404 bgr_0.Vbe2.n41 bgr_0.Vbe2.n40 0.0106786
R7405 bgr_0.Vbe2.n89 bgr_0.Vbe2.n88 0.0106786
R7406 bgr_0.Vbe2.n120 bgr_0.Vbe2.n119 0.0106786
R7407 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 0.00996429
R7408 bgr_0.Vbe2.n137 bgr_0.Vbe2.n128 0.00992001
R7409 bgr_0.Vbe2.n121 bgr_0.Vbe2.n5 0.00992001
R7410 bgr_0.Vbe2.n126 bgr_0.Vbe2.n2 0.00992001
R7411 bgr_0.Vbe2.n122 bgr_0.Vbe2.n6 0.00992001
R7412 bgr_0.Vbe2.n125 bgr_0.Vbe2.n1 0.00992001
R7413 bgr_0.Vbe2.n128 bgr_0.Vbe2.n3 0.00992001
R7414 bgr_0.Vbe2.n121 bgr_0.Vbe2.n3 0.00992001
R7415 bgr_0.Vbe2.n126 bgr_0.Vbe2.n5 0.00992001
R7416 bgr_0.Vbe2.n122 bgr_0.Vbe2.n2 0.00992001
R7417 bgr_0.Vbe2.n125 bgr_0.Vbe2.n6 0.00992001
R7418 bgr_0.Vbe2.n87 bgr_0.Vbe2.n21 0.00992001
R7419 bgr_0.Vbe2.n73 bgr_0.Vbe2.n72 0.00992001
R7420 bgr_0.Vbe2.n75 bgr_0.Vbe2.n70 0.00992001
R7421 bgr_0.Vbe2.n85 bgr_0.Vbe2.n74 0.00992001
R7422 bgr_0.Vbe2.n84 bgr_0.Vbe2.n69 0.00992001
R7423 bgr_0.Vbe2.n71 bgr_0.Vbe2.n21 0.00992001
R7424 bgr_0.Vbe2.n72 bgr_0.Vbe2.n71 0.00992001
R7425 bgr_0.Vbe2.n75 bgr_0.Vbe2.n73 0.00992001
R7426 bgr_0.Vbe2.n74 bgr_0.Vbe2.n70 0.00992001
R7427 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 0.00992001
R7428 bgr_0.Vbe2.n103 bgr_0.Vbe2.n102 0.00889286
R7429 bgr_0.Vbe2.n42 bgr_0.Vbe2.n41 0.00817857
R7430 bgr_0.Vbe2.n120 bgr_0.Vbe2.n7 0.00817857
R7431 bgr_0.V_TOP.n0 bgr_0.V_TOP.t15 369.534
R7432 bgr_0.V_TOP.n10 bgr_0.V_TOP.n8 339.959
R7433 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R7434 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R7435 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R7436 bgr_0.V_TOP.n10 bgr_0.V_TOP.n9 339.272
R7437 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 334.772
R7438 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R7439 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R7440 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R7441 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R7442 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R7443 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R7444 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R7445 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R7446 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R7447 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R7448 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R7449 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R7450 bgr_0.V_TOP bgr_0.V_TOP.t47 214.222
R7451 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R7452 bgr_0.V_TOP.n7 bgr_0.V_TOP.t9 176.114
R7453 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R7454 bgr_0.V_TOP.n0 bgr_0.V_TOP.t49 144.601
R7455 bgr_0.V_TOP.n1 bgr_0.V_TOP.t42 144.601
R7456 bgr_0.V_TOP.n2 bgr_0.V_TOP.t37 144.601
R7457 bgr_0.V_TOP.n3 bgr_0.V_TOP.t24 144.601
R7458 bgr_0.V_TOP.n4 bgr_0.V_TOP.t44 144.601
R7459 bgr_0.V_TOP.n5 bgr_0.V_TOP.t38 144.601
R7460 bgr_0.V_TOP.n27 bgr_0.V_TOP.t14 144.601
R7461 bgr_0.V_TOP.n26 bgr_0.V_TOP.t25 144.601
R7462 bgr_0.V_TOP.n25 bgr_0.V_TOP.t29 144.601
R7463 bgr_0.V_TOP.n24 bgr_0.V_TOP.t34 144.601
R7464 bgr_0.V_TOP.n23 bgr_0.V_TOP.t17 144.601
R7465 bgr_0.V_TOP.n22 bgr_0.V_TOP.t20 144.601
R7466 bgr_0.V_TOP.n21 bgr_0.V_TOP.t31 144.601
R7467 bgr_0.V_TOP.n20 bgr_0.V_TOP.t36 144.601
R7468 bgr_0.V_TOP.n18 bgr_0.V_TOP.t6 95.447
R7469 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R7470 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R7471 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R7472 bgr_0.V_TOP.n6 bgr_0.V_TOP.t8 39.4005
R7473 bgr_0.V_TOP.n6 bgr_0.V_TOP.t4 39.4005
R7474 bgr_0.V_TOP.n11 bgr_0.V_TOP.t1 39.4005
R7475 bgr_0.V_TOP.n11 bgr_0.V_TOP.t10 39.4005
R7476 bgr_0.V_TOP.n9 bgr_0.V_TOP.t2 39.4005
R7477 bgr_0.V_TOP.n9 bgr_0.V_TOP.t12 39.4005
R7478 bgr_0.V_TOP.n8 bgr_0.V_TOP.t13 39.4005
R7479 bgr_0.V_TOP.n8 bgr_0.V_TOP.t3 39.4005
R7480 bgr_0.V_TOP.n14 bgr_0.V_TOP.t0 39.4005
R7481 bgr_0.V_TOP.n14 bgr_0.V_TOP.t7 39.4005
R7482 bgr_0.V_TOP.n16 bgr_0.V_TOP.t5 39.4005
R7483 bgr_0.V_TOP.n16 bgr_0.V_TOP.t11 39.4005
R7484 bgr_0.V_TOP.n12 bgr_0.V_TOP.n10 8.313
R7485 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R7486 bgr_0.V_TOP.n28 bgr_0.V_TOP.t30 4.8295
R7487 bgr_0.V_TOP.n29 bgr_0.V_TOP.t21 4.8295
R7488 bgr_0.V_TOP.n31 bgr_0.V_TOP.t40 4.8295
R7489 bgr_0.V_TOP.n32 bgr_0.V_TOP.t26 4.8295
R7490 bgr_0.V_TOP.n34 bgr_0.V_TOP.t28 4.8295
R7491 bgr_0.V_TOP.n35 bgr_0.V_TOP.t18 4.8295
R7492 bgr_0.V_TOP.n37 bgr_0.V_TOP.t43 4.8295
R7493 bgr_0.V_TOP.n28 bgr_0.V_TOP.t41 4.5005
R7494 bgr_0.V_TOP.n30 bgr_0.V_TOP.t35 4.5005
R7495 bgr_0.V_TOP.n29 bgr_0.V_TOP.t48 4.5005
R7496 bgr_0.V_TOP.n31 bgr_0.V_TOP.t16 4.5005
R7497 bgr_0.V_TOP.n33 bgr_0.V_TOP.t46 4.5005
R7498 bgr_0.V_TOP.n32 bgr_0.V_TOP.t19 4.5005
R7499 bgr_0.V_TOP.n34 bgr_0.V_TOP.t39 4.5005
R7500 bgr_0.V_TOP.n36 bgr_0.V_TOP.t33 4.5005
R7501 bgr_0.V_TOP.n35 bgr_0.V_TOP.t45 4.5005
R7502 bgr_0.V_TOP.n40 bgr_0.V_TOP.t22 4.5005
R7503 bgr_0.V_TOP.n39 bgr_0.V_TOP.t27 4.5005
R7504 bgr_0.V_TOP.n38 bgr_0.V_TOP.t23 4.5005
R7505 bgr_0.V_TOP.n37 bgr_0.V_TOP.t32 4.5005
R7506 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R7507 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R7508 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R7509 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R7510 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R7511 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R7512 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R7513 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R7514 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R7515 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R7516 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R7517 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R7518 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R7519 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R7520 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R7521 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R7522 bgr_0.START_UP.n1 bgr_0.START_UP.t7 238.322
R7523 bgr_0.START_UP.n1 bgr_0.START_UP.t6 238.322
R7524 bgr_0.START_UP.n5 bgr_0.START_UP.n4 175.558
R7525 bgr_0.START_UP.n4 bgr_0.START_UP.n3 168.935
R7526 bgr_0.START_UP.n2 bgr_0.START_UP.n1 166.925
R7527 bgr_0.START_UP.n0 bgr_0.START_UP.t5 130.001
R7528 bgr_0.START_UP.n0 bgr_0.START_UP.t4 81.7084
R7529 bgr_0.START_UP.n2 bgr_0.START_UP.n0 53.0427
R7530 bgr_0.START_UP.n3 bgr_0.START_UP.t1 13.1338
R7531 bgr_0.START_UP.n3 bgr_0.START_UP.t0 13.1338
R7532 bgr_0.START_UP.t3 bgr_0.START_UP.n5 13.1338
R7533 bgr_0.START_UP.n5 bgr_0.START_UP.t2 13.1338
R7534 bgr_0.START_UP.n4 bgr_0.START_UP.n2 4.21925
R7535 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 525.38
R7536 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 525.38
R7537 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 366.856
R7538 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 366.856
R7539 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7540 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 281.168
R7541 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 281.168
R7542 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 281.168
R7543 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7544 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7545 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7546 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7547 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7548 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7549 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7550 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7551 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 39.5005
R7552 a_5750_2946.t0 a_5750_2946.t1 169.905
R7553 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7554 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7555 bgr_0.Vin+.n0 bgr_0.Vin+.t9 303.259
R7556 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R7557 bgr_0.Vin+.n0 bgr_0.Vin+.t8 174.726
R7558 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R7559 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R7560 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R7561 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R7562 bgr_0.Vin+.n8 bgr_0.Vin+.t5 158.796
R7563 bgr_0.Vin+.t4 bgr_0.Vin+.n8 147.981
R7564 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7565 bgr_0.Vin+.n3 bgr_0.Vin+.t10 96.4005
R7566 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R7567 bgr_0.Vin+.n5 bgr_0.Vin+.t1 13.1338
R7568 bgr_0.Vin+.n5 bgr_0.Vin+.t0 13.1338
R7569 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R7570 bgr_0.Vin+.n4 bgr_0.Vin+.t2 13.1338
R7571 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R7572 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.t27 355.293
R7573 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t20 346.8
R7574 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.n7 339.522
R7575 bgr_0.1st_Vout_1.n21 bgr_0.1st_Vout_1.n20 339.522
R7576 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n11 335.022
R7577 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.t3 275.909
R7578 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n12 227.909
R7579 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 222.034
R7580 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.t28 184.097
R7581 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.t24 184.097
R7582 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t30 184.097
R7583 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t25 184.097
R7584 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.n18 166.05
R7585 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.n9 166.05
R7586 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t2 48.0005
R7587 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t0 48.0005
R7588 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t1 48.0005
R7589 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t4 48.0005
R7590 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t5 39.4005
R7591 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t7 39.4005
R7592 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t8 39.4005
R7593 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t6 39.4005
R7594 bgr_0.1st_Vout_1.t10 bgr_0.1st_Vout_1.n21 39.4005
R7595 bgr_0.1st_Vout_1.n21 bgr_0.1st_Vout_1.t9 39.4005
R7596 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.n4 33.1711
R7597 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t36 4.8295
R7598 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t15 4.8295
R7599 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t17 4.8295
R7600 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t21 4.8295
R7601 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t35 4.8295
R7602 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t13 4.8295
R7603 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t31 4.8295
R7604 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n13 4.5005
R7605 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t18 4.5005
R7606 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t12 4.5005
R7607 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t33 4.5005
R7608 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t22 4.5005
R7609 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t19 4.5005
R7610 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t14 4.5005
R7611 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t16 4.5005
R7612 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t11 4.5005
R7613 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t32 4.5005
R7614 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t26 4.5005
R7615 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t34 4.5005
R7616 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t29 4.5005
R7617 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t23 4.5005
R7618 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.n16 4.5005
R7619 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.n10 1.3755
R7620 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 1.3755
R7621 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.n6 1.188
R7622 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.9875
R7623 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n0 0.8935
R7624 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n15 0.78175
R7625 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.6585
R7626 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n1 0.6585
R7627 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.n8 0.6255
R7628 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.n17 0.6255
R7629 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 0.6115
R7630 bgr_0.V_p_1.n1 bgr_0.V_p_1.n2 229.562
R7631 bgr_0.V_p_1.n0 bgr_0.V_p_1.n5 228.939
R7632 bgr_0.V_p_1.n0 bgr_0.V_p_1.n4 228.939
R7633 bgr_0.V_p_1.n1 bgr_0.V_p_1.n3 228.939
R7634 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 228.938
R7635 bgr_0.V_p_1.n0 bgr_0.V_p_1.t0 98.2282
R7636 bgr_0.V_p_1.n5 bgr_0.V_p_1.t6 48.0005
R7637 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R7638 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R7639 bgr_0.V_p_1.n4 bgr_0.V_p_1.t3 48.0005
R7640 bgr_0.V_p_1.n3 bgr_0.V_p_1.t5 48.0005
R7641 bgr_0.V_p_1.n3 bgr_0.V_p_1.t10 48.0005
R7642 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R7643 bgr_0.V_p_1.n2 bgr_0.V_p_1.t4 48.0005
R7644 bgr_0.V_p_1.n6 bgr_0.V_p_1.t1 48.0005
R7645 bgr_0.V_p_1.t7 bgr_0.V_p_1.n6 48.0005
R7646 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R7647 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7648 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7649 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7650 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7651 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t23 660.109
R7652 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t20 660.109
R7653 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n14 428.8
R7654 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n15 428.8
R7655 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.VD3.n16 239.915
R7656 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.VD3.n17 239.915
R7657 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n19 230.4
R7658 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n21 230.4
R7659 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n14 198.4
R7660 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n15 198.4
R7661 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n11 160.428
R7662 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 160.427
R7663 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 160.427
R7664 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 160.053
R7665 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 159.803
R7666 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 159.803
R7667 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 159.802
R7668 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n3 159.802
R7669 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 159.802
R7670 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 155.302
R7671 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t22 155.125
R7672 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t25 155.125
R7673 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n27 146.002
R7674 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t24 98.2764
R7675 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t10 98.2764
R7676 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.t3 98.2764
R7677 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.t34 98.2764
R7678 two_stage_opamp_dummy_magic_0.VD3.t26 two_stage_opamp_dummy_magic_0.VD3.t36 98.2764
R7679 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.VD3.t5 98.2764
R7680 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.VD3.t17 98.2764
R7681 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t8 98.2764
R7682 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t14 98.2764
R7683 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.t21 98.2764
R7684 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.n14 92.5005
R7685 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n25 92.5005
R7686 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 92.5005
R7687 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 92.5005
R7688 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 92.5005
R7689 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.n23 92.5005
R7690 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t26 49.1384
R7691 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t28 49.1384
R7692 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 21.3338
R7693 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 21.3338
R7694 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n26 19.2005
R7695 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n28 13.8005
R7696 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t6 11.2576
R7697 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t18 11.2576
R7698 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t19 11.2576
R7699 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t16 11.2576
R7700 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t12 11.2576
R7701 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t0 11.2576
R7702 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R7703 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R7704 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R7705 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t33 11.2576
R7706 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R7707 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t2 11.2576
R7708 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R7709 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t32 11.2576
R7710 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R7711 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R7712 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t35 11.2576
R7713 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R7714 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R7715 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t4 11.2576
R7716 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R7717 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R7718 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n33 5.40675
R7719 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n8 4.5005
R7720 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n10 0.78175
R7721 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R7722 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R7723 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n6 0.6255
R7724 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n29 0.6255
R7725 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n13 0.6255
R7726 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n31 0.2505
R7727 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 628.034
R7728 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 626.784
R7729 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 626.784
R7730 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 289.2
R7731 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 289.2
R7732 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 228.252
R7733 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 212.733
R7734 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 212.733
R7735 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 176.733
R7736 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 176.733
R7737 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R7738 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 176.733
R7739 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 176.733
R7740 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 152
R7741 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 152
R7742 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R7743 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R7744 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 112.468
R7745 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 112.468
R7746 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R7747 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R7748 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 112.468
R7749 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 112.468
R7750 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 78.8005
R7751 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 78.8005
R7752 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R7753 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R7754 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R7755 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R7756 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 48.0005
R7757 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 48.0005
R7758 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 48.0005
R7759 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 48.0005
R7760 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 48.0005
R7761 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 48.0005
R7762 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 45.5227
R7763 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 45.5227
R7764 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 45.5227
R7765 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R7766 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 33.8443
R7767 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 14.2693
R7768 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 14.2693
R7769 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 1.2505
R7770 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 1.2505
R7771 bgr_0.cap_res1.t0 bgr_0.cap_res1.t7 178.633
R7772 bgr_0.cap_res1.t9 bgr_0.cap_res1.t6 0.1603
R7773 bgr_0.cap_res1.t3 bgr_0.cap_res1.t8 0.1603
R7774 bgr_0.cap_res1.t5 bgr_0.cap_res1.t18 0.1603
R7775 bgr_0.cap_res1.t15 bgr_0.cap_res1.t2 0.1603
R7776 bgr_0.cap_res1.t17 bgr_0.cap_res1.t11 0.1603
R7777 bgr_0.cap_res1.t10 bgr_0.cap_res1.t14 0.1603
R7778 bgr_0.cap_res1.t4 bgr_0.cap_res1.t16 0.1603
R7779 bgr_0.cap_res1.t13 bgr_0.cap_res1.t1 0.1603
R7780 bgr_0.cap_res1.n1 bgr_0.cap_res1.t19 0.159278
R7781 bgr_0.cap_res1.n2 bgr_0.cap_res1.t12 0.159278
R7782 bgr_0.cap_res1.n3 bgr_0.cap_res1.t20 0.159278
R7783 bgr_0.cap_res1.n3 bgr_0.cap_res1.t9 0.1368
R7784 bgr_0.cap_res1.n3 bgr_0.cap_res1.t3 0.1368
R7785 bgr_0.cap_res1.n2 bgr_0.cap_res1.t5 0.1368
R7786 bgr_0.cap_res1.n2 bgr_0.cap_res1.t15 0.1368
R7787 bgr_0.cap_res1.n1 bgr_0.cap_res1.t17 0.1368
R7788 bgr_0.cap_res1.n1 bgr_0.cap_res1.t10 0.1368
R7789 bgr_0.cap_res1.n0 bgr_0.cap_res1.t4 0.1368
R7790 bgr_0.cap_res1.n0 bgr_0.cap_res1.t13 0.1368
R7791 bgr_0.cap_res1.t19 bgr_0.cap_res1.n0 0.00152174
R7792 bgr_0.cap_res1.t12 bgr_0.cap_res1.n1 0.00152174
R7793 bgr_0.cap_res1.t20 bgr_0.cap_res1.n2 0.00152174
R7794 bgr_0.cap_res1.t7 bgr_0.cap_res1.n3 0.00152174
R7795 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t16 623.701
R7796 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t23 611.739
R7797 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R7798 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t17 611.739
R7799 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.t26 611.739
R7800 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R7801 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R7802 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R7803 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R7804 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R7805 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R7806 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R7807 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R7808 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R7809 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t20 421.75
R7810 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t25 421.75
R7811 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t12 421.75
R7812 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R7813 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R7814 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R7815 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R7816 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 176.964
R7817 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n12 172.436
R7818 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.n17 167.094
R7819 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R7820 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R7821 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n13 167.094
R7822 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R7823 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R7824 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.n8 167.094
R7825 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R7826 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R7827 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.n4 167.094
R7828 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R7829 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R7830 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 166.25
R7831 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n0 139.638
R7832 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 139.638
R7833 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n1 134.577
R7834 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 74.1567
R7835 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 47.1294
R7836 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n16 47.1294
R7837 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 47.1294
R7838 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n7 47.1294
R7839 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R7840 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R7841 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R7842 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R7843 two_stage_opamp_dummy_magic_0.Vb3.t5 two_stage_opamp_dummy_magic_0.Vb3.n26 24.0005
R7844 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R7845 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 16.8755
R7846 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t7 10.9449
R7847 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t0 10.9449
R7848 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n3 10.9067
R7849 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n24 4.5005
R7850 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7851 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7852 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t14 449.868
R7853 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t18 449.868
R7854 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n21 339.961
R7855 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 339.272
R7856 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7857 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7858 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7859 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R7860 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7861 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7862 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7863 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7864 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7865 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7866 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7867 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7868 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R7869 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7870 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7871 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7872 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t1 184.625
R7873 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R7874 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.n15 176.733
R7875 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7876 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 176.733
R7877 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n11 176.733
R7878 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 176.733
R7879 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R7880 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.n6 176.733
R7881 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7882 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 176.733
R7883 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.n2 176.733
R7884 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R7885 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n9 170.269
R7886 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 165.8
R7887 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t0 61.1914
R7888 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 56.2338
R7889 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n13 56.2338
R7890 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 56.2338
R7891 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n4 56.2338
R7892 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n20 54.4067
R7893 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7894 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.t2 39.4005
R7895 two_stage_opamp_dummy_magic_0.Vb1.t3 two_stage_opamp_dummy_magic_0.Vb1.n23 39.4005
R7896 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7897 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 22.3599
R7898 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n0 6.81097
R7899 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n7 114.719
R7900 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7901 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n8 114.156
R7902 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7903 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7904 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7905 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7906 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7907 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7908 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7909 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7910 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7911 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7912 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7913 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7914 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7915 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7916 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7917 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7918 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7919 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7920 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7921 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7922 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7923 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7924 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7925 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7926 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7927 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7928 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7929 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7930 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7931 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7932 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7933 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7934 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7935 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7936 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7937 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7938 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 0.563
R7939 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7940 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7941 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7942 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7943 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7944 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7945 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7946 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7947 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7948 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7949 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7950 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7951 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7952 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7953 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7954 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7955 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7956 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7957 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7958 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7959 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7960 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7961 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7962 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7963 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7964 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7965 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7966 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7967 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7968 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7969 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7970 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7971 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7972 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7973 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7974 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7975 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7976 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.3272
R7977 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R7978 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R7979 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R7980 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7981 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7982 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R7983 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R7984 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R7985 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R7986 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R7987 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R7988 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R7989 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.n0 165.8
R7990 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R7991 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R7992 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R7993 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R7994 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R7995 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R7996 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t3 117.591
R7997 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t2 117.591
R7998 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t1 108.424
R7999 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 108.424
R8000 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 42.6121
R8001 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 21.2996
R8002 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n8 17.0005
R8003 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 3.31612
R8004 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 1.26612
R8005 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.2505
R8006 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n4 1.15363
R8007 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t20 369.534
R8008 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t16 369.534
R8009 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.t15 369.534
R8010 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t27 369.534
R8011 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R8012 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t14 369.534
R8013 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.n4 341.397
R8014 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R8015 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.n5 339.272
R8016 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 334.772
R8017 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t18 238.322
R8018 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t29 238.322
R8019 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t3 194.895
R8020 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t23 192.8
R8021 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t13 192.8
R8022 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t26 192.8
R8023 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t17 192.8
R8024 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t10 192.8
R8025 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t22 192.8
R8026 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t12 192.8
R8027 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t25 192.8
R8028 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.t28 192.8
R8029 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t19 192.8
R8030 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t11 192.8
R8031 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t24 192.8
R8032 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R8033 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R8034 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.n22 176.733
R8035 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R8036 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R8037 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R8038 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 171.321
R8039 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n3 169.394
R8040 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n2 168.166
R8041 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R8042 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t2 100.635
R8043 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R8044 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n20 56.2338
R8045 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 56.2338
R8046 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n15 56.2338
R8047 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R8048 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R8049 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.t4 39.4005
R8050 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.t1 39.4005
R8051 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t8 39.4005
R8052 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t6 39.4005
R8053 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.t9 39.4005
R8054 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.t7 39.4005
R8055 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t0 39.4005
R8056 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t5 39.4005
R8057 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 26.9067
R8058 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.n11 5.15675
R8059 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n9 4.5005
R8060 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 4.188
R8061 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n14 3.03175
R8062 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 2.1255
R8063 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.n8 2.1255
R8064 VIN-.n4 VIN-.t8 485.021
R8065 VIN-.n1 VIN-.t6 484.159
R8066 VIN-.n5 VIN-.t7 483.358
R8067 VIN-.n8 VIN-.t10 431.536
R8068 VIN-.n2 VIN-.t9 431.536
R8069 VIN-.n6 VIN-.t1 431.257
R8070 VIN-.n0 VIN-.t0 431.257
R8071 VIN-.n6 VIN-.t2 289.908
R8072 VIN-.n0 VIN-.t5 289.908
R8073 VIN-.n8 VIN-.t4 279.183
R8074 VIN-.n2 VIN-.t3 279.183
R8075 VIN-.n7 VIN-.n6 233.374
R8076 VIN-.n1 VIN-.n0 233.374
R8077 VIN-.n9 VIN-.n8 188.989
R8078 VIN-.n3 VIN-.n2 188.989
R8079 VIN-.n4 VIN-.n3 2.463
R8080 VIN- VIN-.n9 2.03175
R8081 VIN-.n5 VIN-.n4 1.563
R8082 VIN-.n3 VIN-.n1 1.2755
R8083 VIN-.n9 VIN-.n7 1.2755
R8084 VIN-.n7 VIN-.n5 0.8005
R8085 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t0 202.595
R8086 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n3 118.168
R8087 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n0 117.831
R8088 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n35 117.269
R8089 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n10 117.269
R8090 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.n8 117.269
R8091 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n6 117.269
R8092 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n4 117.269
R8093 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n1 117.269
R8094 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.n37 117.267
R8095 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n12 113.136
R8096 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n13 101.335
R8097 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n14 99.647
R8098 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.n28 99.0845
R8099 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.n26 99.0845
R8100 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n24 99.0845
R8101 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n22 99.0845
R8102 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n17 99.0845
R8103 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n15 99.0845
R8104 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n31 94.5845
R8105 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.n19 94.5845
R8106 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.t31 16.0005
R8107 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.t16 16.0005
R8108 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t11 16.0005
R8109 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t38 16.0005
R8110 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t12 16.0005
R8111 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t27 16.0005
R8112 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t32 16.0005
R8113 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t17 16.0005
R8114 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t18 16.0005
R8115 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t7 16.0005
R8116 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t34 16.0005
R8117 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t15 16.0005
R8118 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t10 16.0005
R8119 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t35 16.0005
R8120 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t37 16.0005
R8121 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t14 16.0005
R8122 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t13 16.0005
R8123 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t36 16.0005
R8124 two_stage_opamp_dummy_magic_0.V_p.t19 two_stage_opamp_dummy_magic_0.V_p.n38 16.0005
R8125 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.t33 16.0005
R8126 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t29 9.6005
R8127 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t4 9.6005
R8128 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.t23 9.6005
R8129 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.t40 9.6005
R8130 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t6 9.6005
R8131 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t3 9.6005
R8132 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t9 9.6005
R8133 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t5 9.6005
R8134 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t8 9.6005
R8135 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t26 9.6005
R8136 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t20 9.6005
R8137 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t25 9.6005
R8138 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.t1 9.6005
R8139 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.t24 9.6005
R8140 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t2 9.6005
R8141 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t21 9.6005
R8142 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t28 9.6005
R8143 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t22 9.6005
R8144 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t39 9.6005
R8145 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t30 9.6005
R8146 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n20 4.5005
R8147 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n30 4.5005
R8148 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n33 4.5005
R8149 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n11 3.65675
R8150 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n32 1.28175
R8151 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n16 0.563
R8152 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n18 0.563
R8153 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n21 0.563
R8154 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n23 0.563
R8155 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.n25 0.563
R8156 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.n27 0.563
R8157 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n29 0.563
R8158 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n5 0.563
R8159 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.n7 0.563
R8160 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n9 0.563
R8161 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n36 0.563
R8162 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n2 0.563
R8163 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n34 0.53175
R8164 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t16 681.128
R8165 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 619.134
R8166 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t24 611.739
R8167 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t12 611.739
R8168 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t18 611.739
R8169 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t27 611.739
R8170 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t28 421.75
R8171 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R8172 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R8173 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R8174 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t31 421.75
R8175 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R8176 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R8177 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R8178 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R8179 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R8180 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R8181 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R8182 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t22 421.75
R8183 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R8184 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R8185 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R8186 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t1 288.166
R8187 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 169.125
R8188 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n18 169.125
R8189 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n23 167.094
R8190 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 167.094
R8191 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.n25 167.094
R8192 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 167.094
R8193 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 167.094
R8194 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 167.094
R8195 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.n14 167.094
R8196 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R8197 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R8198 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.n10 167.094
R8199 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R8200 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R8201 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n3 140.546
R8202 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n0 140.546
R8203 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n1 139.296
R8204 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 139.296
R8205 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 73.938
R8206 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t0 62.5402
R8207 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t2 62.5402
R8208 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n26 47.1294
R8209 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n22 47.1294
R8210 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 47.1294
R8211 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n13 47.1294
R8212 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 32.5005
R8213 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R8214 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t10 24.0005
R8215 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R8216 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R8217 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R8218 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R8219 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R8220 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t8 24.0005
R8221 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 14.6443
R8222 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n9 6.15675
R8223 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n6 5.6255
R8224 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n2 3.71925
R8225 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n5 3.71925
R8226 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1.t1 178.194
R8227 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 610.534
R8228 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 610.534
R8229 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R8230 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R8231 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R8232 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R8233 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R8234 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R8235 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R8236 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R8237 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R8238 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R8239 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 433.8
R8240 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R8241 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R8242 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R8243 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R8244 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R8245 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R8246 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 433.8
R8247 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.836
R8248 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 339.834
R8249 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R8250 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 334.772
R8251 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 221.293
R8252 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R8253 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R8254 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R8255 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R8256 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R8257 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R8258 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 176.733
R8259 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 176.733
R8260 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R8261 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R8262 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 176.733
R8263 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 176.733
R8264 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R8265 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R8266 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R8267 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R8268 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 118.45
R8269 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 78.2817
R8270 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 64.5795
R8271 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 56.2338
R8272 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 56.2338
R8273 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 53.2453
R8274 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R8275 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 39.4005
R8276 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R8277 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R8278 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R8279 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R8280 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R8281 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 39.4005
R8282 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R8283 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R8284 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R8285 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 16.0005
R8286 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 4.5005
R8287 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R8288 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R8289 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R8290 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t4 303.259
R8291 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R8292 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R8293 bgr_0.V_CUR_REF_REG.t2 bgr_0.V_CUR_REF_REG.n5 245.284
R8294 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t5 174.726
R8295 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t7 174.726
R8296 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R8297 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R8298 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t3 96.4005
R8299 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t0 39.4005
R8300 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t1 39.4005
R8301 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8302 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8303 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8304 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8305 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t32 660.109
R8306 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t35 660.109
R8307 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 428.8
R8308 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n0 428.8
R8309 two_stage_opamp_dummy_magic_0.VD4.t33 two_stage_opamp_dummy_magic_0.VD4.n8 239.915
R8310 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t36 239.915
R8311 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 230.4
R8312 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n3 230.4
R8313 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 198.4
R8314 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n0 198.4
R8315 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n28 160.428
R8316 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 160.427
R8317 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n14 160.427
R8318 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n13 160.053
R8319 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n29 159.803
R8320 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.803
R8321 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 159.802
R8322 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 159.802
R8323 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 159.802
R8324 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n23 155.302
R8325 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t34 155.125
R8326 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t37 155.125
R8327 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 146.004
R8328 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t33 98.2764
R8329 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t12 98.2764
R8330 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t18 98.2764
R8331 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.VD4.t26 98.2764
R8332 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.VD4.t22 98.2764
R8333 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t30 98.2764
R8334 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t14 98.2764
R8335 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.VD4.t20 98.2764
R8336 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t16 98.2764
R8337 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.VD4.t24 98.2764
R8338 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R8339 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.n6 92.5005
R8340 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n7 92.5005
R8341 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n0 92.5005
R8342 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8343 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8344 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t28 49.1384
R8345 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.VD4.n9 49.1384
R8346 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n4 21.3338
R8347 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.n2 21.3338
R8348 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n12 19.2005
R8349 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 13.8005
R8350 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R8351 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R8352 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R8353 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R8354 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R8355 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R8356 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t5 11.2576
R8357 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R8358 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8359 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R8360 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R8361 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t3 11.2576
R8362 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R8363 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t4 11.2576
R8364 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R8365 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R8366 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R8367 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t2 11.2576
R8368 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R8369 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R8370 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R8371 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.VD4.n33 11.2576
R8372 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 6.188
R8373 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n22 4.5005
R8374 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 0.6255
R8375 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n17 0.6255
R8376 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n19 0.6255
R8377 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 0.6255
R8378 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n27 0.6255
R8379 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.2505
R8380 VIN+.n9 VIN+.t5 485.127
R8381 VIN+.n4 VIN+.t3 485.127
R8382 VIN+.n3 VIN+.t4 485.127
R8383 VIN+.n7 VIN+.t9 318.656
R8384 VIN+.n7 VIN+.t2 318.656
R8385 VIN+.n5 VIN+.t7 318.656
R8386 VIN+.n5 VIN+.t1 318.656
R8387 VIN+.n1 VIN+.t8 318.656
R8388 VIN+.n1 VIN+.t6 318.656
R8389 VIN+.n0 VIN+.t10 318.656
R8390 VIN+.n0 VIN+.t0 318.656
R8391 VIN+.n2 VIN+.n0 167.05
R8392 VIN+.n8 VIN+.n7 165.8
R8393 VIN+.n6 VIN+.n5 165.8
R8394 VIN+.n2 VIN+.n1 165.8
R8395 VIN+.n6 VIN+.n4 2.34425
R8396 VIN+.n4 VIN+.n3 1.3005
R8397 VIN+.n8 VIN+.n6 1.2505
R8398 VIN+ VIN+.n9 1.213
R8399 VIN+.n3 VIN+.n2 1.15675
R8400 VIN+.n9 VIN+.n8 1.15675
R8401 a_n9700_9790.t0 a_n9700_9790.t1 258.591
R8402 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t12 650.729
R8403 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n6 630.607
R8404 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 627.128
R8405 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n10 627.128
R8406 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 227.784
R8407 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 226.534
R8408 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n3 226.534
R8409 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8410 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t10 78.8005
R8411 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t7 78.8005
R8412 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t9 78.8005
R8413 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t6 78.8005
R8414 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t8 78.8005
R8415 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t2 48.0005
R8416 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t4 48.0005
R8417 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t1 48.0005
R8418 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t3 48.0005
R8419 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t11 48.0005
R8420 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t5 48.0005
R8421 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n5 21.1255
R8422 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.n4 10.8755
R8423 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n7 1.3755
R8424 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.2505
R8425 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 1.2505
R8426 a_5230_5758.t0 a_5230_5758.t1 294.339
R8427 a_14520_5738.t0 a_14520_5738.t1 294.339
R8428 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2655
R8429 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 2595
R8430 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2280
R8431 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 2250
R8432 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 672.159
R8433 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 672.159
R8434 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 276.8
R8435 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 240
R8436 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 206.4
R8437 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 204.8
R8438 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 180.904
R8439 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 170.3
R8440 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 160.517
R8441 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 160.517
R8442 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 110.425
R8443 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 110.05
R8444 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 95.7988
R8445 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8446 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8447 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 92.5005
R8448 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8449 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 89.6005
R8450 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 89.6005
R8451 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 76.8005
R8452 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 75.9449
R8453 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 75.9449
R8454 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 47.8997
R8455 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 47.8997
R8456 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 38.4005
R8457 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 24.5338
R8458 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 24.5338
R8459 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 16.8187
R8460 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 16.8187
R8461 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 12.313
R8462 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 12.313
R8463 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 10.9449
R8464 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 10.9449
R8465 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8466 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 4.5005
R8467 bgr_0.Vin-.n11 bgr_0.Vin-.t9 688.859
R8468 bgr_0.Vin-.n13 bgr_0.Vin-.n12 514.134
R8469 bgr_0.Vin-.n9 bgr_0.Vin-.n8 345.116
R8470 bgr_0.Vin-.n15 bgr_0.Vin-.n14 214.713
R8471 bgr_0.Vin-.n11 bgr_0.Vin-.t11 174.726
R8472 bgr_0.Vin-.n12 bgr_0.Vin-.t12 174.726
R8473 bgr_0.Vin-.n13 bgr_0.Vin-.t8 174.726
R8474 bgr_0.Vin-.n14 bgr_0.Vin-.t10 174.726
R8475 bgr_0.Vin-.n7 bgr_0.Vin-.n5 173.029
R8476 bgr_0.Vin-.n7 bgr_0.Vin-.n6 168.654
R8477 bgr_0.Vin-.n9 bgr_0.Vin-.t4 162.921
R8478 bgr_0.Vin-.n12 bgr_0.Vin-.n11 128.534
R8479 bgr_0.Vin-.n14 bgr_0.Vin-.n13 128.534
R8480 bgr_0.Vin-.n1 bgr_0.Vin-.n0 83.5719
R8481 bgr_0.Vin-.n22 bgr_0.Vin-.n21 83.5719
R8482 bgr_0.Vin-.n20 bgr_0.Vin-.n19 83.5719
R8483 bgr_0.Vin-.n25 bgr_0.Vin-.n1 73.682
R8484 bgr_0.Vin-.n20 bgr_0.Vin-.n4 73.3165
R8485 bgr_0.Vin-.n8 bgr_0.Vin-.t6 39.4005
R8486 bgr_0.Vin-.n8 bgr_0.Vin-.t5 39.4005
R8487 bgr_0.Vin-.n21 bgr_0.Vin-.n20 26.074
R8488 bgr_0.Vin-.t7 bgr_0.Vin-.n1 25.7843
R8489 bgr_0.Vin-.n16 bgr_0.Vin-.n15 17.526
R8490 bgr_0.Vin-.n6 bgr_0.Vin-.t3 13.1338
R8491 bgr_0.Vin-.n6 bgr_0.Vin-.t0 13.1338
R8492 bgr_0.Vin-.n5 bgr_0.Vin-.t2 13.1338
R8493 bgr_0.Vin-.n5 bgr_0.Vin-.t1 13.1338
R8494 bgr_0.Vin-.n15 bgr_0.Vin-.n10 12.5317
R8495 bgr_0.Vin-.n10 bgr_0.Vin-.n9 6.40675
R8496 bgr_0.Vin-.n10 bgr_0.Vin-.n7 3.8755
R8497 bgr_0.Vin-.n16 bgr_0.Vin-.n4 2.19742
R8498 bgr_0.Vin-.n24 bgr_0.Vin-.n23 1.5505
R8499 bgr_0.Vin-.n3 bgr_0.Vin-.n2 1.5505
R8500 bgr_0.Vin-.n18 bgr_0.Vin-.n17 1.5505
R8501 bgr_0.Vin-.n18 bgr_0.Vin-.n4 1.19225
R8502 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n25 1.07742
R8503 bgr_0.Vin-.n23 bgr_0.Vin-.n22 1.07024
R8504 bgr_0.Vin-.n19 bgr_0.Vin-.n18 0.959578
R8505 bgr_0.Vin-.n19 bgr_0.Vin-.n3 0.885803
R8506 bgr_0.Vin-.n22 bgr_0.Vin-.n3 0.77514
R8507 bgr_0.Vin-.n25 bgr_0.Vin-.n24 0.763532
R8508 bgr_0.Vin-.n23 bgr_0.Vin-.n0 0.590702
R8509 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.498483
R8510 bgr_0.Vin-.n21 bgr_0.Vin-.t7 0.290206
R8511 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.0183571
R8512 bgr_0.Vin-.n17 bgr_0.Vin-.n2 0.0183571
R8513 bgr_0.Vin-.n24 bgr_0.Vin-.n2 0.0183571
R8514 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 220.678
R8515 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R8516 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R8517 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R8518 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t1 9.6005
R8519 a_5350_5758.t0 a_5350_5758.t1 169.905
R8520 a_14240_2946.t0 a_14240_2946.t1 169.905
R8521 a_n8798_9040.t0 a_n8798_9040.t1 376.99
R8522 a_n7190_9400.t0 a_n7190_9400.t1 258.591
R8523 a_n9760_9260.t0 a_n9760_9260.t1 258.591
C0 VOUT- two_stage_opamp_dummy_magic_0.V_err_gate 0.068595f
C1 VDDA bgr_0.1st_Vout_2 2.79809f
C2 bgr_0.V_TOP bgr_0.PFET_GATE_10uA 2.47368f
C3 m2_n4150_7140# bgr_0.V_TOP 0.012f
C4 VIN- VIN+ 0.555219f
C5 VOUT- two_stage_opamp_dummy_magic_0.cap_res_X 50.7533f
C6 VDDA li_n2700_10430# 0.021911f
C7 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_gate 4.78237f
C8 VDDA bgr_0.PFET_GATE_10uA 10.3925f
C9 m2_n4150_7140# VDDA 0.010446f
C10 VDDA bgr_0.V_TOP 16.1354f
C11 VDDA two_stage_opamp_dummy_magic_0.VD3 3.70112f
C12 VDDA two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.963643f
C13 VOUT+ two_stage_opamp_dummy_magic_0.cap_res_X 0.020189f
C14 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.cap_res_X 1.25369f
C15 li_n4800_10220# bgr_0.1st_Vout_2 0.020658f
C16 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.1st_Vout_2 1.24865f
C17 m2_n2790_7140# bgr_0.1st_Vout_2 0.075543f
C18 VDDA two_stage_opamp_dummy_magic_0.err_amp_out 1.00936f
C19 VDDA two_stage_opamp_dummy_magic_0.Y 4.15025f
C20 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.cap_res_X 0.356357f
C21 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.VD1 0.017583f
C22 VOUT+ two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.059472f
C23 VDDA VOUT- 6.78335f
C24 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.VD1 1.06369f
C25 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.PFET_GATE_10uA 2.46518f
C26 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.V_TOP 1.13839f
C27 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.Y 0.040365f
C28 VDDA VOUT+ 6.69232f
C29 m2_n2790_7140# bgr_0.PFET_GATE_10uA 0.012f
C30 bgr_0.V_TOP li_n1300_10330# 0.020062f
C31 VDDA two_stage_opamp_dummy_magic_0.V_err_amp_ref 3.85441f
C32 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.V_err_gate 0.01134f
C33 VOUT+ two_stage_opamp_dummy_magic_0.Y 2.10995f
C34 m2_n2790_7140# VDDA 0.010446f
C35 VIN- two_stage_opamp_dummy_magic_0.VD1 0.881219f
C36 VOUT- VOUT+ 0.210644f
C37 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.err_amp_out 0.406563f
C38 VDDA two_stage_opamp_dummy_magic_0.V_err_gate 3.57771f
C39 VIN+ two_stage_opamp_dummy_magic_0.VD1 0.057219f
C40 VOUT- two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.068695f
C41 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.cap_res_X 0.04831f
C42 bgr_0.1st_Vout_2 bgr_0.PFET_GATE_10uA 1.24195f
C43 bgr_0.V_TOP bgr_0.1st_Vout_2 1.46737f
C44 VDDA two_stage_opamp_dummy_magic_0.cap_res_X 1.05846f
C45 VIN+ GNDA 2.09083f
C46 VIN- GNDA 2.156752f
C47 VOUT+ GNDA 17.60256f
C48 VOUT- GNDA 17.193665f
C49 VDDA GNDA 0.156674p
C50 li_n4800_10220# GNDA 0.043891f $ **FLOATING
C51 li_n6200_10220# GNDA 0.049096f $ **FLOATING
C52 li_n1300_10330# GNDA 0.047034f $ **FLOATING
C53 li_n8300_10330# GNDA 0.049721f $ **FLOATING
C54 li_n9700_10330# GNDA 0.050514f $ **FLOATING
C55 li_n2700_10430# GNDA 0.050654f $ **FLOATING
C56 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.38758f
C57 two_stage_opamp_dummy_magic_0.Y GNDA 4.963086f
C58 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 32.13635f
C59 bgr_0.1st_Vout_2 GNDA 5.078303f
C60 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.945237f
C61 bgr_0.V_TOP GNDA 6.845387f
C62 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 8.815428f
C63 bgr_0.PFET_GATE_10uA GNDA 5.13248f
C64 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 9.47159f
C65 two_stage_opamp_dummy_magic_0.VD3 GNDA 6.535289f
C66 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.61725f
C67 bgr_0.Vin-.n0 GNDA 0.048818f
C68 bgr_0.Vin-.n1 GNDA 0.333648f
C69 bgr_0.Vin-.n2 GNDA 0.166915f
C70 bgr_0.Vin-.n3 GNDA 0.074468f
C71 bgr_0.Vin-.n4 GNDA 0.338979f
C72 bgr_0.Vin-.t2 GNDA 0.028614f
C73 bgr_0.Vin-.t1 GNDA 0.028614f
C74 bgr_0.Vin-.n5 GNDA 0.099613f
C75 bgr_0.Vin-.t3 GNDA 0.028614f
C76 bgr_0.Vin-.t0 GNDA 0.028614f
C77 bgr_0.Vin-.n6 GNDA 0.095121f
C78 bgr_0.Vin-.n7 GNDA 0.408067f
C79 bgr_0.Vin-.t4 GNDA 0.098662f
C80 bgr_0.Vin-.n8 GNDA 0.025702f
C81 bgr_0.Vin-.n9 GNDA 0.469862f
C82 bgr_0.Vin-.n10 GNDA 0.222852f
C83 bgr_0.Vin-.t9 GNDA 0.023594f
C84 bgr_0.Vin-.n11 GNDA 0.027673f
C85 bgr_0.Vin-.n12 GNDA 0.022653f
C86 bgr_0.Vin-.n13 GNDA 0.022653f
C87 bgr_0.Vin-.n14 GNDA 0.040466f
C88 bgr_0.Vin-.n15 GNDA 0.524007f
C89 bgr_0.Vin-.n16 GNDA 0.461299f
C90 bgr_0.Vin-.n17 GNDA 0.166915f
C91 bgr_0.Vin-.n18 GNDA 0.10855f
C92 bgr_0.Vin-.n19 GNDA 0.082742f
C93 bgr_0.Vin-.n20 GNDA 0.331333f
C94 bgr_0.Vin-.t7 GNDA 0.072966f
C95 bgr_0.Vin-.n21 GNDA 0.073776f
C96 bgr_0.Vin-.n22 GNDA 0.082742f
C97 bgr_0.Vin-.n23 GNDA 0.074468f
C98 bgr_0.Vin-.n24 GNDA 0.656866f
C99 bgr_0.Vin-.n25 GNDA 0.389111f
C100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.086659f
C101 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA 0.013381f
C102 two_stage_opamp_dummy_magic_0.err_amp_out.t3 GNDA 0.013381f
C103 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.038511f
C104 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA 0.013381f
C105 two_stage_opamp_dummy_magic_0.err_amp_out.t4 GNDA 0.013381f
C106 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.037365f
C107 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.464702f
C108 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA 0.013381f
C109 two_stage_opamp_dummy_magic_0.err_amp_out.t5 GNDA 0.013381f
C110 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.037365f
C111 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.496077f
C112 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.095614f
C113 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 1.60863f
C114 two_stage_opamp_dummy_magic_0.err_amp_out.t0 GNDA 0.013381f
C115 two_stage_opamp_dummy_magic_0.err_amp_out.t10 GNDA 0.013381f
C116 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 0.031078f
C117 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.918238f
C118 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA 0.013381f
C119 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA 0.013381f
C120 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.031328f
C121 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.351359f
C122 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA 0.013381f
C123 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA 0.013381f
C124 two_stage_opamp_dummy_magic_0.err_amp_out.n10 GNDA 0.031328f
C125 VIN+.t0 GNDA 0.041803f
C126 VIN+.t10 GNDA 0.041803f
C127 VIN+.n0 GNDA 0.086391f
C128 VIN+.t6 GNDA 0.041803f
C129 VIN+.t8 GNDA 0.041803f
C130 VIN+.n1 GNDA 0.085194f
C131 VIN+.n2 GNDA 0.359761f
C132 VIN+.t4 GNDA 0.058811f
C133 VIN+.n3 GNDA 0.215335f
C134 VIN+.t3 GNDA 0.058811f
C135 VIN+.n4 GNDA 0.262589f
C136 VIN+.t1 GNDA 0.041803f
C137 VIN+.t7 GNDA 0.041803f
C138 VIN+.n5 GNDA 0.085194f
C139 VIN+.n6 GNDA 0.248358f
C140 VIN+.t2 GNDA 0.041803f
C141 VIN+.t9 GNDA 0.041803f
C142 VIN+.n7 GNDA 0.085194f
C143 VIN+.n8 GNDA 0.200956f
C144 VIN+.t5 GNDA 0.058811f
C145 VIN+.n9 GNDA 0.211601f
C146 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.024416f
C147 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.069509f
C148 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.094519f
C149 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.120449f
C150 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.042516f
C151 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.078578f
C152 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.050655f
C153 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.120449f
C154 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.042516f
C155 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.078578f
C156 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.050655f
C157 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.050227f
C158 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.094519f
C159 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.281683f
C160 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.420453f
C161 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.242764f
C162 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.242764f
C163 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.242764f
C164 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.242764f
C165 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.182073f
C166 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.121382f
C167 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.182073f
C168 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.242764f
C169 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.242764f
C170 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.242764f
C171 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.242764f
C172 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.420453f
C173 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.281683f
C174 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.069509f
C175 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.097309f
C176 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.024416f
C177 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.024416f
C178 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.084727f
C179 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.024416f
C180 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.024416f
C181 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.084913f
C182 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.024416f
C183 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.024416f
C184 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.084913f
C185 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.024416f
C186 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.024416f
C187 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.084613f
C188 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.15974f
C189 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.024416f
C190 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.024416f
C191 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.084613f
C192 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.082811f
C193 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.024416f
C194 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.024416f
C195 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.084613f
C196 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.082811f
C197 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.099252f
C198 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.024416f
C199 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.024416f
C200 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.08286f
C201 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.100481f
C202 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.094683f
C203 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.024416f
C204 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.024416f
C205 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.084612f
C206 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.078625f
C207 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.024416f
C208 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.024416f
C209 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.084913f
C210 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.024416f
C211 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.024416f
C212 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.084612f
C213 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.15974f
C214 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.029845f
C215 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.057972f
C216 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.079606f
C217 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.024416f
C218 bgr_0.V_CUR_REF_REG.t4 GNDA 0.014208f
C219 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C220 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C221 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C222 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C223 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C224 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C225 bgr_0.V_CUR_REF_REG.t2 GNDA 0.42777f
C226 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.021072f
C227 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.021072f
C228 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.021072f
C229 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.052748f
C230 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.021072f
C231 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.021072f
C232 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.052748f
C233 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.021072f
C234 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.021072f
C235 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.052465f
C236 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.356252f
C237 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.233824f
C238 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.031607f
C239 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.031607f
C240 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.114383f
C241 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.056103f
C242 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.056103f
C243 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.056103f
C244 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.056103f
C245 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.056103f
C246 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.056103f
C247 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.056103f
C248 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.065481f
C249 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.061738f
C250 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.038719f
C251 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.038719f
C252 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.038719f
C253 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.038719f
C254 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.038719f
C255 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.034599f
C256 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.056103f
C257 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.056103f
C258 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.056103f
C259 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.056103f
C260 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.056103f
C261 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.056103f
C262 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.056103f
C263 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.056103f
C264 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.056103f
C265 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.056103f
C266 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.056103f
C267 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.065481f
C268 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.061738f
C269 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.038719f
C270 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.038719f
C271 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.038719f
C272 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.038719f
C273 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.038719f
C274 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.038719f
C275 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.038719f
C276 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.038719f
C277 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.038719f
C278 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.034599f
C279 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.086466f
C280 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.031607f
C281 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.031607f
C282 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.063214f
C283 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.245032f
C284 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 2.43922f
C285 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 2.08227f
C286 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 0.05082f
C287 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.021072f
C288 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.027982f
C289 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.027982f
C290 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.093821f
C291 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.027982f
C292 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.027982f
C293 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.091248f
C294 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.736953f
C295 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.027982f
C296 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.027982f
C297 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.093821f
C298 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.027982f
C299 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.027982f
C300 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.091248f
C301 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.736953f
C302 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.384386f
C303 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.174317f
C304 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.017629f
C305 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.017629f
C306 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.038202f
C307 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.05475f
C308 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.185713f
C309 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 1.22899f
C310 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.138513f
C311 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.138513f
C312 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.138513f
C313 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.138513f
C314 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.159843f
C315 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.129775f
C316 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.07975f
C317 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.07975f
C318 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.074675f
C319 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.138513f
C320 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.138513f
C321 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.138513f
C322 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.138513f
C323 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.159843f
C324 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.129775f
C325 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.07975f
C326 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.07975f
C327 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.074675f
C328 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.049949f
C329 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.138513f
C330 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.138513f
C331 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.138513f
C332 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.138513f
C333 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.159843f
C334 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.129775f
C335 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.07975f
C336 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.07975f
C337 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 0.074675f
C338 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.138513f
C339 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.138513f
C340 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.138513f
C341 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.138513f
C342 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.159843f
C343 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.129775f
C344 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.07975f
C345 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.07975f
C346 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.074675f
C347 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.049949f
C348 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 1.68217f
C349 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 3.89317f
C350 bgr_0.VB2_CUR_BIAS GNDA 2.74386f
C351 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA 0.014624f
C352 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA 0.014624f
C353 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA 0.014624f
C354 two_stage_opamp_dummy_magic_0.V_p.n0 GNDA 0.052539f
C355 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA 0.014624f
C356 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA 0.014624f
C357 two_stage_opamp_dummy_magic_0.V_p.n1 GNDA 0.052133f
C358 two_stage_opamp_dummy_magic_0.V_p.n2 GNDA 0.176305f
C359 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA 0.014624f
C360 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA 0.014624f
C361 two_stage_opamp_dummy_magic_0.V_p.n3 GNDA 0.052516f
C362 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA 0.014624f
C363 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA 0.014624f
C364 two_stage_opamp_dummy_magic_0.V_p.n4 GNDA 0.052133f
C365 two_stage_opamp_dummy_magic_0.V_p.n5 GNDA 0.174572f
C366 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA 0.014624f
C367 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA 0.014624f
C368 two_stage_opamp_dummy_magic_0.V_p.n6 GNDA 0.052133f
C369 two_stage_opamp_dummy_magic_0.V_p.n7 GNDA 0.091767f
C370 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA 0.014624f
C371 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA 0.014624f
C372 two_stage_opamp_dummy_magic_0.V_p.n8 GNDA 0.052133f
C373 two_stage_opamp_dummy_magic_0.V_p.n9 GNDA 0.091767f
C374 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA 0.014624f
C375 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA 0.014624f
C376 two_stage_opamp_dummy_magic_0.V_p.n10 GNDA 0.052133f
C377 two_stage_opamp_dummy_magic_0.V_p.n11 GNDA 0.140027f
C378 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA 0.014624f
C379 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA 0.014624f
C380 two_stage_opamp_dummy_magic_0.V_p.n12 GNDA 0.049685f
C381 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA 0.024373f
C382 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA 0.024373f
C383 two_stage_opamp_dummy_magic_0.V_p.n13 GNDA 0.099127f
C384 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA 0.024373f
C385 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA 0.024373f
C386 two_stage_opamp_dummy_magic_0.V_p.n14 GNDA 0.097223f
C387 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA 0.024373f
C388 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA 0.024373f
C389 two_stage_opamp_dummy_magic_0.V_p.n15 GNDA 0.096773f
C390 two_stage_opamp_dummy_magic_0.V_p.n16 GNDA 0.165755f
C391 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA 0.024373f
C392 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA 0.024373f
C393 two_stage_opamp_dummy_magic_0.V_p.n17 GNDA 0.096773f
C394 two_stage_opamp_dummy_magic_0.V_p.n18 GNDA 0.086515f
C395 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA 0.085877f
C396 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA 0.024373f
C397 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA 0.024373f
C398 two_stage_opamp_dummy_magic_0.V_p.n19 GNDA 0.094049f
C399 two_stage_opamp_dummy_magic_0.V_p.n20 GNDA 0.56785f
C400 two_stage_opamp_dummy_magic_0.V_p.n21 GNDA 0.029248f
C401 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA 0.024373f
C402 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA 0.024373f
C403 two_stage_opamp_dummy_magic_0.V_p.n22 GNDA 0.096773f
C404 two_stage_opamp_dummy_magic_0.V_p.n23 GNDA 0.086515f
C405 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA 0.024373f
C406 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA 0.024373f
C407 two_stage_opamp_dummy_magic_0.V_p.n24 GNDA 0.096773f
C408 two_stage_opamp_dummy_magic_0.V_p.n25 GNDA 0.086515f
C409 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA 0.024373f
C410 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA 0.024373f
C411 two_stage_opamp_dummy_magic_0.V_p.n26 GNDA 0.096773f
C412 two_stage_opamp_dummy_magic_0.V_p.n27 GNDA 0.086515f
C413 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA 0.024373f
C414 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA 0.024373f
C415 two_stage_opamp_dummy_magic_0.V_p.n28 GNDA 0.096773f
C416 two_stage_opamp_dummy_magic_0.V_p.n29 GNDA 0.086515f
C417 two_stage_opamp_dummy_magic_0.V_p.n30 GNDA 0.159231f
C418 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA 0.024373f
C419 two_stage_opamp_dummy_magic_0.V_p.t4 GNDA 0.024373f
C420 two_stage_opamp_dummy_magic_0.V_p.n31 GNDA 0.094049f
C421 two_stage_opamp_dummy_magic_0.V_p.n32 GNDA 0.078027f
C422 two_stage_opamp_dummy_magic_0.V_p.n33 GNDA 0.082224f
C423 two_stage_opamp_dummy_magic_0.V_p.n34 GNDA 0.07702f
C424 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA 0.014624f
C425 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA 0.014624f
C426 two_stage_opamp_dummy_magic_0.V_p.n35 GNDA 0.052133f
C427 two_stage_opamp_dummy_magic_0.V_p.n36 GNDA 0.09128f
C428 two_stage_opamp_dummy_magic_0.V_p.n37 GNDA 0.091767f
C429 two_stage_opamp_dummy_magic_0.V_p.n38 GNDA 0.052133f
C430 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA 0.014624f
C431 VIN-.t6 GNDA 0.050642f
C432 VIN-.t5 GNDA 0.033412f
C433 VIN-.t0 GNDA 0.041251f
C434 VIN-.n0 GNDA 0.059274f
C435 VIN-.n1 GNDA 0.280478f
C436 VIN-.t3 GNDA 0.032863f
C437 VIN-.t9 GNDA 0.041265f
C438 VIN-.n2 GNDA 0.064892f
C439 VIN-.n3 GNDA 0.200879f
C440 VIN-.t8 GNDA 0.050078f
C441 VIN-.n4 GNDA 0.236241f
C442 VIN-.t7 GNDA 0.050425f
C443 VIN-.n5 GNDA 0.180621f
C444 VIN-.t2 GNDA 0.033412f
C445 VIN-.t1 GNDA 0.041251f
C446 VIN-.n6 GNDA 0.059274f
C447 VIN-.n7 GNDA 0.149629f
C448 VIN-.t4 GNDA 0.032863f
C449 VIN-.t10 GNDA 0.041265f
C450 VIN-.n8 GNDA 0.064892f
C451 VIN-.n9 GNDA 0.186141f
C452 bgr_0.PFET_GATE_10uA.t24 GNDA 0.039179f
C453 bgr_0.PFET_GATE_10uA.t14 GNDA 0.057916f
C454 bgr_0.PFET_GATE_10uA.n0 GNDA 0.063817f
C455 bgr_0.PFET_GATE_10uA.t11 GNDA 0.039179f
C456 bgr_0.PFET_GATE_10uA.t21 GNDA 0.057916f
C457 bgr_0.PFET_GATE_10uA.n1 GNDA 0.063817f
C458 bgr_0.PFET_GATE_10uA.n2 GNDA 0.064022f
C459 bgr_0.PFET_GATE_10uA.t29 GNDA 0.045299f
C460 bgr_0.PFET_GATE_10uA.t18 GNDA 0.045299f
C461 bgr_0.PFET_GATE_10uA.n3 GNDA 0.137138f
C462 bgr_0.PFET_GATE_10uA.t3 GNDA 0.781422f
C463 bgr_0.PFET_GATE_10uA.t0 GNDA 0.040183f
C464 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040183f
C465 bgr_0.PFET_GATE_10uA.n4 GNDA 0.102705f
C466 bgr_0.PFET_GATE_10uA.t9 GNDA 0.040183f
C467 bgr_0.PFET_GATE_10uA.t7 GNDA 0.040183f
C468 bgr_0.PFET_GATE_10uA.n5 GNDA 0.100051f
C469 bgr_0.PFET_GATE_10uA.n6 GNDA 0.978629f
C470 bgr_0.PFET_GATE_10uA.t8 GNDA 0.040183f
C471 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040183f
C472 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100051f
C473 bgr_0.PFET_GATE_10uA.n8 GNDA 0.554934f
C474 bgr_0.PFET_GATE_10uA.t2 GNDA 0.586977f
C475 bgr_0.PFET_GATE_10uA.n9 GNDA 1.13286f
C476 bgr_0.PFET_GATE_10uA.t4 GNDA 0.040183f
C477 bgr_0.PFET_GATE_10uA.t1 GNDA 0.040183f
C478 bgr_0.PFET_GATE_10uA.n10 GNDA 0.096913f
C479 bgr_0.PFET_GATE_10uA.n11 GNDA 0.356682f
C480 bgr_0.PFET_GATE_10uA.n12 GNDA 3.84996f
C481 bgr_0.PFET_GATE_10uA.n13 GNDA 1.78858f
C482 bgr_0.PFET_GATE_10uA.n14 GNDA 1.41725f
C483 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039179f
C484 bgr_0.PFET_GATE_10uA.t27 GNDA 0.057916f
C485 bgr_0.PFET_GATE_10uA.n15 GNDA 0.063817f
C486 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039179f
C487 bgr_0.PFET_GATE_10uA.t15 GNDA 0.057916f
C488 bgr_0.PFET_GATE_10uA.n16 GNDA 0.063817f
C489 bgr_0.PFET_GATE_10uA.n17 GNDA 0.076791f
C490 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039179f
C491 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039179f
C492 bgr_0.PFET_GATE_10uA.t25 GNDA 0.039179f
C493 bgr_0.PFET_GATE_10uA.t16 GNDA 0.057916f
C494 bgr_0.PFET_GATE_10uA.n18 GNDA 0.071675f
C495 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051234f
C496 bgr_0.PFET_GATE_10uA.n20 GNDA 0.043376f
C497 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039179f
C498 bgr_0.PFET_GATE_10uA.t17 GNDA 0.039179f
C499 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039179f
C500 bgr_0.PFET_GATE_10uA.t13 GNDA 0.039179f
C501 bgr_0.PFET_GATE_10uA.t23 GNDA 0.039179f
C502 bgr_0.PFET_GATE_10uA.t20 GNDA 0.057916f
C503 bgr_0.PFET_GATE_10uA.n21 GNDA 0.071675f
C504 bgr_0.PFET_GATE_10uA.n22 GNDA 0.051234f
C505 bgr_0.PFET_GATE_10uA.n23 GNDA 0.051234f
C506 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051234f
C507 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043376f
C508 bgr_0.PFET_GATE_10uA.n26 GNDA 0.05954f
C509 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.098962f
C510 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.011218f
C511 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.018267f
C512 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.106822f
C513 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.021464f
C514 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.095301f
C515 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.011144f
C516 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.091464f
C517 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.021464f
C518 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.066547f
C519 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.021464f
C520 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.204094f
C521 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.098951f
C522 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.092891f
C523 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.321853f
C524 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 0.772935f
C525 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.513063f
C526 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.092891f
C527 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.02127f
C528 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020358f
C529 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020407f
C530 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021244f
C531 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.021116f
C532 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.299998f
C533 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.021116f
C534 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.156484f
C535 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.021116f
C536 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.190977f
C537 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.153542f
C538 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.133374f
C539 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.242929f
C540 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.02127f
C541 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020976f
C542 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.328367f
C543 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020976f
C544 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.180843f
C545 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.180843f
C546 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020976f
C547 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.030602f
C548 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.030602f
C549 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.030602f
C550 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.098572f
C551 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.030602f
C552 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.030602f
C553 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.092431f
C554 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.110167f
C555 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.110167f
C556 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.405846f
C557 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.175527f
C558 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 1.31573f
C559 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.15148f
C560 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.15148f
C561 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.15148f
C562 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.15148f
C563 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.174807f
C564 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.141924f
C565 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.087216f
C566 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.087216f
C567 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.081666f
C568 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.15148f
C569 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.15148f
C570 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.15148f
C571 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.15148f
C572 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.174807f
C573 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.141924f
C574 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.087216f
C575 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.087216f
C576 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.081666f
C577 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.067093f
C578 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.15148f
C579 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.15148f
C580 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.15148f
C581 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.15148f
C582 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.174807f
C583 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.141924f
C584 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.087216f
C585 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.087216f
C586 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.081666f
C587 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.15148f
C588 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.15148f
C589 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.15148f
C590 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.15148f
C591 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.174807f
C592 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.141924f
C593 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.087216f
C594 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.087216f
C595 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.081666f
C596 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.049314f
C597 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 1.55338f
C598 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 3.93468f
C599 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 3.04649f
C600 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.543425f
C601 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 0.098572f
C602 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.030602f
C603 bgr_0.cap_res1.t8 GNDA 0.417173f
C604 bgr_0.cap_res1.t3 GNDA 0.418684f
C605 bgr_0.cap_res1.t6 GNDA 0.417173f
C606 bgr_0.cap_res1.t9 GNDA 0.418684f
C607 bgr_0.cap_res1.t2 GNDA 0.417173f
C608 bgr_0.cap_res1.t15 GNDA 0.418684f
C609 bgr_0.cap_res1.t18 GNDA 0.417173f
C610 bgr_0.cap_res1.t5 GNDA 0.418684f
C611 bgr_0.cap_res1.t14 GNDA 0.417173f
C612 bgr_0.cap_res1.t10 GNDA 0.418684f
C613 bgr_0.cap_res1.t11 GNDA 0.417173f
C614 bgr_0.cap_res1.t17 GNDA 0.418684f
C615 bgr_0.cap_res1.t1 GNDA 0.417173f
C616 bgr_0.cap_res1.t13 GNDA 0.418684f
C617 bgr_0.cap_res1.t16 GNDA 0.417173f
C618 bgr_0.cap_res1.t4 GNDA 0.418684f
C619 bgr_0.cap_res1.n0 GNDA 0.279631f
C620 bgr_0.cap_res1.t19 GNDA 0.222685f
C621 bgr_0.cap_res1.n1 GNDA 0.303406f
C622 bgr_0.cap_res1.t12 GNDA 0.222685f
C623 bgr_0.cap_res1.n2 GNDA 0.303406f
C624 bgr_0.cap_res1.t20 GNDA 0.222685f
C625 bgr_0.cap_res1.n3 GNDA 0.303406f
C626 bgr_0.cap_res1.t7 GNDA 0.649059f
C627 bgr_0.cap_res1.t0 GNDA 0.10618f
C628 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA 0.020233f
C629 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 GNDA 0.020233f
C630 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 GNDA 0.020233f
C631 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 GNDA 0.047731f
C632 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA 0.020233f
C633 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 GNDA 0.020233f
C634 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 GNDA 0.046922f
C635 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 GNDA 0.884615f
C636 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA 0.020233f
C637 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA 0.020233f
C638 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 GNDA 0.046922f
C639 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 GNDA 2.10658f
C640 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 GNDA 1.98101f
C641 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA 0.020233f
C642 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA 0.020233f
C643 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 GNDA 0.04777f
C644 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA 0.016692f
C645 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA 0.016692f
C646 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA 0.016692f
C647 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA 0.016692f
C648 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA 0.016692f
C649 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA 0.036166f
C650 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 GNDA 0.051623f
C651 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA 0.020233f
C652 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA 0.020233f
C653 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 GNDA 0.04777f
C654 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 GNDA 0.17992f
C655 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 GNDA 0.05811f
C656 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 GNDA 0.039231f
C657 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 GNDA 0.044006f
C658 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 GNDA 0.044006f
C659 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 GNDA 0.039231f
C660 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA 0.016692f
C661 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 GNDA 0.016692f
C662 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA 0.016692f
C663 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA 0.036166f
C664 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 GNDA 0.056399f
C665 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 GNDA 0.044006f
C666 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 GNDA 0.039231f
C667 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 GNDA 0.05811f
C668 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 GNDA 0.17992f
C669 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 GNDA 0.746838f
C670 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 GNDA 0.061393f
C671 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA 0.020233f
C672 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.03144f
C673 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.03144f
C674 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.10934f
C675 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.03144f
C676 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.03144f
C677 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.108953f
C678 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.205692f
C679 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.03144f
C680 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.03144f
C681 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.108953f
C682 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.106633f
C683 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.03144f
C684 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.03144f
C685 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.108953f
C686 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.106633f
C687 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.03144f
C688 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.03144f
C689 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.10934f
C690 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.127804f
C691 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.03144f
C692 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.03144f
C693 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.106696f
C694 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.089361f
C695 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.03144f
C696 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.03144f
C697 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.10934f
C698 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.03144f
C699 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.03144f
C700 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.108953f
C701 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.205693f
C702 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.089505f
C703 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.089505f
C704 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.362715f
C705 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.362715f
C706 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.541405f
C707 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.3126f
C708 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.3126f
C709 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.3126f
C710 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.3126f
C711 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.23445f
C712 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.155099f
C713 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.054747f
C714 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.101182f
C715 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.065226f
C716 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.155099f
C717 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.054747f
C718 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.101182f
C719 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.065226f
C720 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.064676f
C721 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.12171f
C722 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.541405f
C723 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.3126f
C724 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.3126f
C725 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.3126f
C726 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.3126f
C727 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.23445f
C728 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.1563f
C729 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.12171f
C730 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.125303f
C731 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.03144f
C732 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.03144f
C733 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.102506f
C734 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.074649f
C735 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.038431f
C736 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.03144f
C737 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.03144f
C738 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.108953f
C739 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.101243f
C740 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.03144f
C741 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.03144f
C742 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.1091f
C743 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.116136f
C744 bgr_0.1st_Vout_1.n0 GNDA 0.96394f
C745 bgr_0.1st_Vout_1.n1 GNDA 0.23261f
C746 bgr_0.1st_Vout_1.n2 GNDA 0.23261f
C747 bgr_0.1st_Vout_1.n3 GNDA 0.96394f
C748 bgr_0.1st_Vout_1.n4 GNDA 0.588341f
C749 bgr_0.1st_Vout_1.n5 GNDA 0.23261f
C750 bgr_0.1st_Vout_1.t27 GNDA 0.020816f
C751 bgr_0.1st_Vout_1.t26 GNDA 0.346936f
C752 bgr_0.1st_Vout_1.t36 GNDA 0.352846f
C753 bgr_0.1st_Vout_1.t18 GNDA 0.346936f
C754 bgr_0.1st_Vout_1.t12 GNDA 0.346936f
C755 bgr_0.1st_Vout_1.t15 GNDA 0.352846f
C756 bgr_0.1st_Vout_1.t33 GNDA 0.346936f
C757 bgr_0.1st_Vout_1.t17 GNDA 0.352846f
C758 bgr_0.1st_Vout_1.t22 GNDA 0.346936f
C759 bgr_0.1st_Vout_1.t19 GNDA 0.346936f
C760 bgr_0.1st_Vout_1.t21 GNDA 0.352846f
C761 bgr_0.1st_Vout_1.t14 GNDA 0.346936f
C762 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C763 bgr_0.1st_Vout_1.t16 GNDA 0.346936f
C764 bgr_0.1st_Vout_1.t11 GNDA 0.346936f
C765 bgr_0.1st_Vout_1.t13 GNDA 0.352846f
C766 bgr_0.1st_Vout_1.t32 GNDA 0.346936f
C767 bgr_0.1st_Vout_1.t31 GNDA 0.352846f
C768 bgr_0.1st_Vout_1.t23 GNDA 0.346936f
C769 bgr_0.1st_Vout_1.t29 GNDA 0.346936f
C770 bgr_0.1st_Vout_1.t34 GNDA 0.346936f
C771 bgr_0.1st_Vout_1.t20 GNDA 0.022665f
C772 bgr_0.1st_Vout_1.n6 GNDA 0.389472f
C773 bgr_0.1st_Vout_1.n7 GNDA 0.021864f
C774 bgr_0.1st_Vout_1.n8 GNDA 0.103033f
C775 bgr_0.1st_Vout_1.t25 GNDA 0.013213f
C776 bgr_0.1st_Vout_1.t30 GNDA 0.013213f
C777 bgr_0.1st_Vout_1.n9 GNDA 0.029393f
C778 bgr_0.1st_Vout_1.n10 GNDA 0.081221f
C779 bgr_0.1st_Vout_1.n11 GNDA 0.020958f
C780 bgr_0.1st_Vout_1.n12 GNDA 0.012529f
C781 bgr_0.1st_Vout_1.t3 GNDA 0.018268f
C782 bgr_0.1st_Vout_1.n13 GNDA 0.189508f
C783 bgr_0.1st_Vout_1.n14 GNDA 0.011336f
C784 bgr_0.1st_Vout_1.n15 GNDA 0.048077f
C785 bgr_0.1st_Vout_1.n16 GNDA 0.077485f
C786 bgr_0.1st_Vout_1.n17 GNDA 0.038163f
C787 bgr_0.1st_Vout_1.t24 GNDA 0.013213f
C788 bgr_0.1st_Vout_1.t28 GNDA 0.013213f
C789 bgr_0.1st_Vout_1.n18 GNDA 0.029393f
C790 bgr_0.1st_Vout_1.n19 GNDA 0.081221f
C791 bgr_0.1st_Vout_1.n20 GNDA 0.166349f
C792 bgr_0.1st_Vout_1.n21 GNDA 0.021864f
C793 bgr_0.Vin+.t9 GNDA 0.020459f
C794 bgr_0.Vin+.t8 GNDA 0.013299f
C795 bgr_0.Vin+.n0 GNDA 0.04388f
C796 bgr_0.Vin+.t6 GNDA 0.013299f
C797 bgr_0.Vin+.n1 GNDA 0.034146f
C798 bgr_0.Vin+.t7 GNDA 0.013299f
C799 bgr_0.Vin+.n2 GNDA 0.034607f
C800 bgr_0.Vin+.n3 GNDA 0.074523f
C801 bgr_0.Vin+.t3 GNDA 0.043132f
C802 bgr_0.Vin+.t2 GNDA 0.043132f
C803 bgr_0.Vin+.n4 GNDA 0.144858f
C804 bgr_0.Vin+.t1 GNDA 0.043132f
C805 bgr_0.Vin+.t0 GNDA 0.043132f
C806 bgr_0.Vin+.n5 GNDA 0.142496f
C807 bgr_0.Vin+.n6 GNDA 0.656763f
C808 bgr_0.Vin+.n7 GNDA 0.71769f
C809 bgr_0.Vin+.t5 GNDA 0.137433f
C810 bgr_0.Vin+.n8 GNDA 0.446219f
C811 bgr_0.Vin+.t4 GNDA 0.125873f
C812 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.163765f
C813 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.409099f
C814 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.409099f
C815 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.485537f
C816 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.256456f
C817 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.162306f
C818 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.446073f
C819 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.149996f
C820 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.917914f
C821 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.446073f
C822 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.409099f
C823 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.409099f
C824 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.485537f
C825 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.256456f
C826 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.162306f
C827 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.149996f
C828 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.917423f
C829 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.163765f
C830 bgr_0.START_UP.t2 GNDA 0.041701f
C831 bgr_0.START_UP.t4 GNDA 1.6623f
C832 bgr_0.START_UP.t5 GNDA 0.043697f
C833 bgr_0.START_UP.n0 GNDA 1.28651f
C834 bgr_0.START_UP.t6 GNDA 0.01567f
C835 bgr_0.START_UP.t7 GNDA 0.01567f
C836 bgr_0.START_UP.n1 GNDA 0.044238f
C837 bgr_0.START_UP.n2 GNDA 0.853868f
C838 bgr_0.START_UP.t1 GNDA 0.041701f
C839 bgr_0.START_UP.t0 GNDA 0.041701f
C840 bgr_0.START_UP.n3 GNDA 0.139173f
C841 bgr_0.START_UP.n4 GNDA 0.720786f
C842 bgr_0.START_UP.n5 GNDA 0.151283f
C843 bgr_0.START_UP.t3 GNDA 0.041701f
C844 bgr_0.V_TOP.t47 GNDA 0.132572f
C845 bgr_0.V_TOP.t14 GNDA 0.115045f
C846 bgr_0.V_TOP.t25 GNDA 0.115045f
C847 bgr_0.V_TOP.t29 GNDA 0.115045f
C848 bgr_0.V_TOP.t34 GNDA 0.115045f
C849 bgr_0.V_TOP.t17 GNDA 0.115045f
C850 bgr_0.V_TOP.t20 GNDA 0.115045f
C851 bgr_0.V_TOP.t31 GNDA 0.115045f
C852 bgr_0.V_TOP.t36 GNDA 0.115045f
C853 bgr_0.V_TOP.t38 GNDA 0.115045f
C854 bgr_0.V_TOP.t44 GNDA 0.115045f
C855 bgr_0.V_TOP.t24 GNDA 0.115045f
C856 bgr_0.V_TOP.t37 GNDA 0.115045f
C857 bgr_0.V_TOP.t42 GNDA 0.115045f
C858 bgr_0.V_TOP.t49 GNDA 0.115045f
C859 bgr_0.V_TOP.t15 GNDA 0.150392f
C860 bgr_0.V_TOP.n0 GNDA 0.084081f
C861 bgr_0.V_TOP.n1 GNDA 0.061357f
C862 bgr_0.V_TOP.n2 GNDA 0.061357f
C863 bgr_0.V_TOP.n3 GNDA 0.061357f
C864 bgr_0.V_TOP.n4 GNDA 0.061357f
C865 bgr_0.V_TOP.n5 GNDA 0.057217f
C866 bgr_0.V_TOP.t6 GNDA 0.147947f
C867 bgr_0.V_TOP.t9 GNDA 0.155772f
C868 bgr_0.V_TOP.t8 GNDA 0.010957f
C869 bgr_0.V_TOP.t4 GNDA 0.010957f
C870 bgr_0.V_TOP.n6 GNDA 0.027281f
C871 bgr_0.V_TOP.n7 GNDA 0.726844f
C872 bgr_0.V_TOP.t13 GNDA 0.010957f
C873 bgr_0.V_TOP.t3 GNDA 0.010957f
C874 bgr_0.V_TOP.n8 GNDA 0.027465f
C875 bgr_0.V_TOP.t2 GNDA 0.010957f
C876 bgr_0.V_TOP.t12 GNDA 0.010957f
C877 bgr_0.V_TOP.n9 GNDA 0.027281f
C878 bgr_0.V_TOP.n10 GNDA 0.252824f
C879 bgr_0.V_TOP.t1 GNDA 0.010957f
C880 bgr_0.V_TOP.t10 GNDA 0.010957f
C881 bgr_0.V_TOP.n11 GNDA 0.026425f
C882 bgr_0.V_TOP.n12 GNDA 0.153577f
C883 bgr_0.V_TOP.n13 GNDA 0.087653f
C884 bgr_0.V_TOP.t0 GNDA 0.010957f
C885 bgr_0.V_TOP.t7 GNDA 0.010957f
C886 bgr_0.V_TOP.n14 GNDA 0.027281f
C887 bgr_0.V_TOP.n15 GNDA 0.151313f
C888 bgr_0.V_TOP.t5 GNDA 0.010957f
C889 bgr_0.V_TOP.t11 GNDA 0.010957f
C890 bgr_0.V_TOP.n16 GNDA 0.027281f
C891 bgr_0.V_TOP.n17 GNDA 0.149874f
C892 bgr_0.V_TOP.n18 GNDA 0.329448f
C893 bgr_0.V_TOP.n19 GNDA 0.023183f
C894 bgr_0.V_TOP.n20 GNDA 0.057217f
C895 bgr_0.V_TOP.n21 GNDA 0.061357f
C896 bgr_0.V_TOP.n22 GNDA 0.061357f
C897 bgr_0.V_TOP.n23 GNDA 0.061357f
C898 bgr_0.V_TOP.n24 GNDA 0.061357f
C899 bgr_0.V_TOP.n25 GNDA 0.061357f
C900 bgr_0.V_TOP.n26 GNDA 0.061357f
C901 bgr_0.V_TOP.n27 GNDA 0.057217f
C902 bgr_0.V_TOP.t22 GNDA 0.438267f
C903 bgr_0.V_TOP.t30 GNDA 0.445732f
C904 bgr_0.V_TOP.t41 GNDA 0.438267f
C905 bgr_0.V_TOP.n28 GNDA 0.293844f
C906 bgr_0.V_TOP.t35 GNDA 0.438267f
C907 bgr_0.V_TOP.t21 GNDA 0.445732f
C908 bgr_0.V_TOP.t48 GNDA 0.438267f
C909 bgr_0.V_TOP.n29 GNDA 0.293844f
C910 bgr_0.V_TOP.n30 GNDA 0.273917f
C911 bgr_0.V_TOP.t40 GNDA 0.445732f
C912 bgr_0.V_TOP.t16 GNDA 0.438267f
C913 bgr_0.V_TOP.n31 GNDA 0.293844f
C914 bgr_0.V_TOP.t46 GNDA 0.438267f
C915 bgr_0.V_TOP.t26 GNDA 0.445732f
C916 bgr_0.V_TOP.t19 GNDA 0.438267f
C917 bgr_0.V_TOP.n32 GNDA 0.293844f
C918 bgr_0.V_TOP.n33 GNDA 0.356092f
C919 bgr_0.V_TOP.t28 GNDA 0.445732f
C920 bgr_0.V_TOP.t39 GNDA 0.438267f
C921 bgr_0.V_TOP.n34 GNDA 0.293844f
C922 bgr_0.V_TOP.t33 GNDA 0.438267f
C923 bgr_0.V_TOP.t18 GNDA 0.445732f
C924 bgr_0.V_TOP.t45 GNDA 0.438267f
C925 bgr_0.V_TOP.n35 GNDA 0.293844f
C926 bgr_0.V_TOP.n36 GNDA 0.356092f
C927 bgr_0.V_TOP.t43 GNDA 0.445732f
C928 bgr_0.V_TOP.t32 GNDA 0.438267f
C929 bgr_0.V_TOP.n37 GNDA 0.293844f
C930 bgr_0.V_TOP.t23 GNDA 0.438267f
C931 bgr_0.V_TOP.n38 GNDA 0.273917f
C932 bgr_0.V_TOP.t27 GNDA 0.438267f
C933 bgr_0.V_TOP.n39 GNDA 0.191742f
C934 bgr_0.V_TOP.n40 GNDA 0.893239f
C935 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.345114f
C936 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.346365f
C937 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.345114f
C938 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.34782f
C939 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.378304f
C940 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.345114f
C941 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.346365f
C942 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.345114f
C943 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.346365f
C944 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.345114f
C945 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.346365f
C946 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.345114f
C947 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.346365f
C948 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.345114f
C949 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.346365f
C950 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.345114f
C951 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.346365f
C952 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.345114f
C953 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.346365f
C954 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.345114f
C955 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.346365f
C956 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.345114f
C957 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.346365f
C958 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.345114f
C959 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.346365f
C960 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.345114f
C961 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.346365f
C962 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.345114f
C963 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.346365f
C964 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.345114f
C965 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.346365f
C966 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.345114f
C967 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.346365f
C968 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.345114f
C969 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.346365f
C970 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.345114f
C971 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.346365f
C972 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.345114f
C973 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.346365f
C974 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.345114f
C975 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.346365f
C976 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.345114f
C977 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.346365f
C978 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.345114f
C979 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.346365f
C980 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.345114f
C981 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.346365f
C982 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.345114f
C983 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.346365f
C984 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.345114f
C985 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.346365f
C986 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.345114f
C987 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.346365f
C988 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.345114f
C989 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.346365f
C990 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.345114f
C991 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.346365f
C992 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.345114f
C993 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.346365f
C994 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.345114f
C995 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.346365f
C996 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.345114f
C997 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.346365f
C998 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.345114f
C999 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.362035f
C1000 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.345114f
C1001 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.185368f
C1002 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.198389f
C1003 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.345114f
C1004 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.185368f
C1005 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.196789f
C1006 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.345114f
C1007 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.185368f
C1008 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.196789f
C1009 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.345114f
C1010 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.185368f
C1011 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.196789f
C1012 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.345114f
C1013 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.185368f
C1014 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.196789f
C1015 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.345114f
C1016 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.185368f
C1017 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.196789f
C1018 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.345114f
C1019 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.185368f
C1020 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.196789f
C1021 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.345114f
C1022 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.185368f
C1023 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196789f
C1024 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.345114f
C1025 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.185368f
C1026 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196789f
C1027 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.345114f
C1028 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.346365f
C1029 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.166846f
C1030 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.215207f
C1031 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.18422f
C1032 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.233728f
C1033 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.18422f
C1034 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.250999f
C1035 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.18422f
C1036 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.250999f
C1037 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.18422f
C1038 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.250999f
C1039 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.18422f
C1040 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.250999f
C1041 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.18422f
C1042 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.250999f
C1043 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.18422f
C1044 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.250999f
C1045 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.18422f
C1046 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250999f
C1047 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.18422f
C1048 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250999f
C1049 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.18422f
C1050 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250999f
C1051 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.18422f
C1052 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250999f
C1053 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.18422f
C1054 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250999f
C1055 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.18422f
C1056 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250999f
C1057 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.18422f
C1058 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250999f
C1059 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.18422f
C1060 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250999f
C1061 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.18422f
C1062 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.233728f
C1063 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.343967f
C1064 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.166846f
C1065 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.216458f
C1066 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.343967f
C1067 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.166846f
C1068 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.216458f
C1069 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.343967f
C1070 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.345114f
C1071 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.363635f
C1072 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.363635f
C1073 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.363635f
C1074 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.185368f
C1075 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.216458f
C1076 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.343967f
C1077 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.166846f
C1078 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.197936f
C1079 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.343967f
C1080 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.166846f
C1081 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.216458f
C1082 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.343967f
C1083 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.166846f
C1084 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.216458f
C1085 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.343967f
C1086 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.166846f
C1087 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216458f
C1088 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.343967f
C1089 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.345114f
C1090 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.363635f
C1091 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.363635f
C1092 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.363635f
C1093 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.185368f
C1094 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216458f
C1095 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.343967f
C1096 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.345114f
C1097 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.363635f
C1098 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.363635f
C1099 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.363635f
C1100 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.185368f
C1101 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216458f
C1102 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.343967f
C1103 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216458f
C1104 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.185368f
C1105 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.363635f
C1106 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.363635f
C1107 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.363635f
C1108 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.602274f
C1109 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.298233f
C1110 VOUT+.t0 GNDA 0.043577f
C1111 VOUT+.t15 GNDA 0.043577f
C1112 VOUT+.n0 GNDA 0.175148f
C1113 VOUT+.t10 GNDA 0.043577f
C1114 VOUT+.t14 GNDA 0.043577f
C1115 VOUT+.n1 GNDA 0.174825f
C1116 VOUT+.n2 GNDA 0.172223f
C1117 VOUT+.t9 GNDA 0.043577f
C1118 VOUT+.t13 GNDA 0.043577f
C1119 VOUT+.n3 GNDA 0.174825f
C1120 VOUT+.n4 GNDA 0.088815f
C1121 VOUT+.t7 GNDA 0.043577f
C1122 VOUT+.t11 GNDA 0.043577f
C1123 VOUT+.n5 GNDA 0.174825f
C1124 VOUT+.n6 GNDA 0.088815f
C1125 VOUT+.t6 GNDA 0.043577f
C1126 VOUT+.t1 GNDA 0.043577f
C1127 VOUT+.n7 GNDA 0.175148f
C1128 VOUT+.n8 GNDA 0.105197f
C1129 VOUT+.t8 GNDA 0.043577f
C1130 VOUT+.t12 GNDA 0.043577f
C1131 VOUT+.n9 GNDA 0.172685f
C1132 VOUT+.n10 GNDA 0.210763f
C1133 VOUT+.t117 GNDA 0.295461f
C1134 VOUT+.t26 GNDA 0.290513f
C1135 VOUT+.n11 GNDA 0.194779f
C1136 VOUT+.t124 GNDA 0.290513f
C1137 VOUT+.n12 GNDA 0.127099f
C1138 VOUT+.t72 GNDA 0.295461f
C1139 VOUT+.t39 GNDA 0.290513f
C1140 VOUT+.n13 GNDA 0.194779f
C1141 VOUT+.t127 GNDA 0.290513f
C1142 VOUT+.t35 GNDA 0.294841f
C1143 VOUT+.t87 GNDA 0.294841f
C1144 VOUT+.t43 GNDA 0.294841f
C1145 VOUT+.t96 GNDA 0.294841f
C1146 VOUT+.t143 GNDA 0.294841f
C1147 VOUT+.t106 GNDA 0.294841f
C1148 VOUT+.t154 GNDA 0.294841f
C1149 VOUT+.t65 GNDA 0.294841f
C1150 VOUT+.t116 GNDA 0.294841f
C1151 VOUT+.t73 GNDA 0.294841f
C1152 VOUT+.t149 GNDA 0.290513f
C1153 VOUT+.n14 GNDA 0.195399f
C1154 VOUT+.t59 GNDA 0.290513f
C1155 VOUT+.n15 GNDA 0.24987f
C1156 VOUT+.t97 GNDA 0.290513f
C1157 VOUT+.n16 GNDA 0.24987f
C1158 VOUT+.t131 GNDA 0.290513f
C1159 VOUT+.n17 GNDA 0.24987f
C1160 VOUT+.t24 GNDA 0.290513f
C1161 VOUT+.n18 GNDA 0.24987f
C1162 VOUT+.t75 GNDA 0.290513f
C1163 VOUT+.n19 GNDA 0.24987f
C1164 VOUT+.t112 GNDA 0.290513f
C1165 VOUT+.n20 GNDA 0.24987f
C1166 VOUT+.t144 GNDA 0.290513f
C1167 VOUT+.n21 GNDA 0.24987f
C1168 VOUT+.t55 GNDA 0.290513f
C1169 VOUT+.n22 GNDA 0.24987f
C1170 VOUT+.t95 GNDA 0.290513f
C1171 VOUT+.n23 GNDA 0.24987f
C1172 VOUT+.n24 GNDA 0.236042f
C1173 VOUT+.t38 GNDA 0.295461f
C1174 VOUT+.t142 GNDA 0.290513f
C1175 VOUT+.n25 GNDA 0.194779f
C1176 VOUT+.t94 GNDA 0.290513f
C1177 VOUT+.t20 GNDA 0.295461f
C1178 VOUT+.t58 GNDA 0.290513f
C1179 VOUT+.n26 GNDA 0.194779f
C1180 VOUT+.n27 GNDA 0.236042f
C1181 VOUT+.t80 GNDA 0.295461f
C1182 VOUT+.t42 GNDA 0.290513f
C1183 VOUT+.n28 GNDA 0.194779f
C1184 VOUT+.t133 GNDA 0.290513f
C1185 VOUT+.t61 GNDA 0.295461f
C1186 VOUT+.t100 GNDA 0.290513f
C1187 VOUT+.n29 GNDA 0.194779f
C1188 VOUT+.n30 GNDA 0.236042f
C1189 VOUT+.t121 GNDA 0.295461f
C1190 VOUT+.t84 GNDA 0.290513f
C1191 VOUT+.n31 GNDA 0.194779f
C1192 VOUT+.t32 GNDA 0.290513f
C1193 VOUT+.t104 GNDA 0.295461f
C1194 VOUT+.t137 GNDA 0.290513f
C1195 VOUT+.n32 GNDA 0.194779f
C1196 VOUT+.n33 GNDA 0.236042f
C1197 VOUT+.t85 GNDA 0.295461f
C1198 VOUT+.t50 GNDA 0.290513f
C1199 VOUT+.n34 GNDA 0.194779f
C1200 VOUT+.t138 GNDA 0.290513f
C1201 VOUT+.t67 GNDA 0.295461f
C1202 VOUT+.t103 GNDA 0.290513f
C1203 VOUT+.n35 GNDA 0.194779f
C1204 VOUT+.n36 GNDA 0.236042f
C1205 VOUT+.t123 GNDA 0.295461f
C1206 VOUT+.t90 GNDA 0.290513f
C1207 VOUT+.n37 GNDA 0.194779f
C1208 VOUT+.t36 GNDA 0.290513f
C1209 VOUT+.t107 GNDA 0.295337f
C1210 VOUT+.t141 GNDA 0.290513f
C1211 VOUT+.n38 GNDA 0.193087f
C1212 VOUT+.n39 GNDA 0.236042f
C1213 VOUT+.t108 GNDA 0.295461f
C1214 VOUT+.t70 GNDA 0.290513f
C1215 VOUT+.n40 GNDA 0.194779f
C1216 VOUT+.t91 GNDA 0.290513f
C1217 VOUT+.n41 GNDA 0.127099f
C1218 VOUT+.t68 GNDA 0.295461f
C1219 VOUT+.t31 GNDA 0.290513f
C1220 VOUT+.n42 GNDA 0.194779f
C1221 VOUT+.t52 GNDA 0.290513f
C1222 VOUT+.t54 GNDA 0.294841f
C1223 VOUT+.t156 GNDA 0.294841f
C1224 VOUT+.t145 GNDA 0.295461f
C1225 VOUT+.t45 GNDA 0.290513f
C1226 VOUT+.n43 GNDA 0.194779f
C1227 VOUT+.t136 GNDA 0.290513f
C1228 VOUT+.n44 GNDA 0.127099f
C1229 VOUT+.t101 GNDA 0.290513f
C1230 VOUT+.n45 GNDA 0.12256f
C1231 VOUT+.t37 GNDA 0.294841f
C1232 VOUT+.t113 GNDA 0.295461f
C1233 VOUT+.t151 GNDA 0.290513f
C1234 VOUT+.n46 GNDA 0.194779f
C1235 VOUT+.t98 GNDA 0.290513f
C1236 VOUT+.n47 GNDA 0.127099f
C1237 VOUT+.t60 GNDA 0.290513f
C1238 VOUT+.n48 GNDA 0.12256f
C1239 VOUT+.t140 GNDA 0.294841f
C1240 VOUT+.t76 GNDA 0.295461f
C1241 VOUT+.t118 GNDA 0.290513f
C1242 VOUT+.n49 GNDA 0.194779f
C1243 VOUT+.t57 GNDA 0.290513f
C1244 VOUT+.n50 GNDA 0.127099f
C1245 VOUT+.t21 GNDA 0.290513f
C1246 VOUT+.n51 GNDA 0.12256f
C1247 VOUT+.t105 GNDA 0.294841f
C1248 VOUT+.t25 GNDA 0.295461f
C1249 VOUT+.t66 GNDA 0.290513f
C1250 VOUT+.n52 GNDA 0.194779f
C1251 VOUT+.t81 GNDA 0.290513f
C1252 VOUT+.n53 GNDA 0.127099f
C1253 VOUT+.t44 GNDA 0.290513f
C1254 VOUT+.n54 GNDA 0.12256f
C1255 VOUT+.t125 GNDA 0.294841f
C1256 VOUT+.t88 GNDA 0.294841f
C1257 VOUT+.t51 GNDA 0.294841f
C1258 VOUT+.t150 GNDA 0.294841f
C1259 VOUT+.t33 GNDA 0.294841f
C1260 VOUT+.t134 GNDA 0.290513f
C1261 VOUT+.n55 GNDA 0.195399f
C1262 VOUT+.t110 GNDA 0.290513f
C1263 VOUT+.n56 GNDA 0.24987f
C1264 VOUT+.t147 GNDA 0.290513f
C1265 VOUT+.n57 GNDA 0.24987f
C1266 VOUT+.t46 GNDA 0.290513f
C1267 VOUT+.n58 GNDA 0.24987f
C1268 VOUT+.t86 GNDA 0.290513f
C1269 VOUT+.n59 GNDA 0.30888f
C1270 VOUT+.t62 GNDA 0.290513f
C1271 VOUT+.n60 GNDA 0.30888f
C1272 VOUT+.t102 GNDA 0.290513f
C1273 VOUT+.n61 GNDA 0.30888f
C1274 VOUT+.t139 GNDA 0.290513f
C1275 VOUT+.n62 GNDA 0.30888f
C1276 VOUT+.t119 GNDA 0.290513f
C1277 VOUT+.n63 GNDA 0.24987f
C1278 VOUT+.t155 GNDA 0.290513f
C1279 VOUT+.n64 GNDA 0.24987f
C1280 VOUT+.n65 GNDA 0.236042f
C1281 VOUT+.t28 GNDA 0.295461f
C1282 VOUT+.t130 GNDA 0.290513f
C1283 VOUT+.n66 GNDA 0.194779f
C1284 VOUT+.t152 GNDA 0.290513f
C1285 VOUT+.t77 GNDA 0.295461f
C1286 VOUT+.t115 GNDA 0.290513f
C1287 VOUT+.n67 GNDA 0.194779f
C1288 VOUT+.n68 GNDA 0.236042f
C1289 VOUT+.t63 GNDA 0.295461f
C1290 VOUT+.t23 GNDA 0.290513f
C1291 VOUT+.n69 GNDA 0.194779f
C1292 VOUT+.t48 GNDA 0.290513f
C1293 VOUT+.t111 GNDA 0.295461f
C1294 VOUT+.t148 GNDA 0.290513f
C1295 VOUT+.n70 GNDA 0.194779f
C1296 VOUT+.n71 GNDA 0.236042f
C1297 VOUT+.t114 GNDA 0.295461f
C1298 VOUT+.t79 GNDA 0.290513f
C1299 VOUT+.n72 GNDA 0.194779f
C1300 VOUT+.t27 GNDA 0.290513f
C1301 VOUT+.t99 GNDA 0.295461f
C1302 VOUT+.t132 GNDA 0.290513f
C1303 VOUT+.n73 GNDA 0.194779f
C1304 VOUT+.n74 GNDA 0.236042f
C1305 VOUT+.t74 GNDA 0.295461f
C1306 VOUT+.t40 GNDA 0.290513f
C1307 VOUT+.n75 GNDA 0.194779f
C1308 VOUT+.t128 GNDA 0.290513f
C1309 VOUT+.t56 GNDA 0.295461f
C1310 VOUT+.t93 GNDA 0.290513f
C1311 VOUT+.n76 GNDA 0.194779f
C1312 VOUT+.n77 GNDA 0.236042f
C1313 VOUT+.t109 GNDA 0.295461f
C1314 VOUT+.t71 GNDA 0.290513f
C1315 VOUT+.n78 GNDA 0.194779f
C1316 VOUT+.t19 GNDA 0.290513f
C1317 VOUT+.t92 GNDA 0.295461f
C1318 VOUT+.t126 GNDA 0.290513f
C1319 VOUT+.n79 GNDA 0.194779f
C1320 VOUT+.n80 GNDA 0.236042f
C1321 VOUT+.t69 GNDA 0.295461f
C1322 VOUT+.t34 GNDA 0.290513f
C1323 VOUT+.n81 GNDA 0.194779f
C1324 VOUT+.t122 GNDA 0.290513f
C1325 VOUT+.t53 GNDA 0.295461f
C1326 VOUT+.t89 GNDA 0.290513f
C1327 VOUT+.n82 GNDA 0.194779f
C1328 VOUT+.n83 GNDA 0.236042f
C1329 VOUT+.t30 GNDA 0.295461f
C1330 VOUT+.t135 GNDA 0.290513f
C1331 VOUT+.n84 GNDA 0.194779f
C1332 VOUT+.t83 GNDA 0.290513f
C1333 VOUT+.t153 GNDA 0.295461f
C1334 VOUT+.t49 GNDA 0.290513f
C1335 VOUT+.n85 GNDA 0.194779f
C1336 VOUT+.n86 GNDA 0.236042f
C1337 VOUT+.t64 GNDA 0.295461f
C1338 VOUT+.t29 GNDA 0.290513f
C1339 VOUT+.n87 GNDA 0.194779f
C1340 VOUT+.t120 GNDA 0.290513f
C1341 VOUT+.t47 GNDA 0.295461f
C1342 VOUT+.t82 GNDA 0.290513f
C1343 VOUT+.n88 GNDA 0.194779f
C1344 VOUT+.n89 GNDA 0.236042f
C1345 VOUT+.t22 GNDA 0.295461f
C1346 VOUT+.t129 GNDA 0.290513f
C1347 VOUT+.n90 GNDA 0.194779f
C1348 VOUT+.t78 GNDA 0.290513f
C1349 VOUT+.n91 GNDA 0.236042f
C1350 VOUT+.t41 GNDA 0.290513f
C1351 VOUT+.n92 GNDA 0.127099f
C1352 VOUT+.t146 GNDA 0.290513f
C1353 VOUT+.n93 GNDA 0.238016f
C1354 VOUT+.n94 GNDA 0.268648f
C1355 VOUT+.t2 GNDA 0.05084f
C1356 VOUT+.t16 GNDA 0.05084f
C1357 VOUT+.n95 GNDA 0.235187f
C1358 VOUT+.t18 GNDA 0.05084f
C1359 VOUT+.t4 GNDA 0.05084f
C1360 VOUT+.n96 GNDA 0.2344f
C1361 VOUT+.n97 GNDA 0.144847f
C1362 VOUT+.t17 GNDA 0.05084f
C1363 VOUT+.t5 GNDA 0.05084f
C1364 VOUT+.n98 GNDA 0.2344f
C1365 VOUT+.n99 GNDA 0.089159f
C1366 VOUT+.t3 GNDA 0.084056f
C1367 VOUT+.n100 GNDA 0.119121f
C1368 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.017997f
C1369 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.014955f
C1370 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.09349f
C1371 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.061605f
C1372 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.014854f
C1373 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.014854f
C1374 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.061426f
C1375 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.014854f
C1376 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.014854f
C1377 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.061191f
C1378 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.084841f
C1379 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.014854f
C1380 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.014854f
C1381 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.061191f
C1382 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.044271f
C1383 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.014854f
C1384 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.014854f
C1385 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.061191f
C1386 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.044271f
C1387 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.014854f
C1388 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.014854f
C1389 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.061191f
C1390 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.063995f
C1391 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.767169f
C1392 bgr_0.V_CMFB_S4 GNDA 0.732874f
C1393 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.053187f
C1394 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.053187f
C1395 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.184972f
C1396 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.053187f
C1397 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.053187f
C1398 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.184316f
C1399 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.347971f
C1400 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.053187f
C1401 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.053187f
C1402 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.184316f
C1403 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.180392f
C1404 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.053187f
C1405 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.053187f
C1406 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.184316f
C1407 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.180392f
C1408 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.053187f
C1409 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.053187f
C1410 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.184316f
C1411 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.212415f
C1412 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.053187f
C1413 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.053187f
C1414 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.180498f
C1415 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.149147f
C1416 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.022794f
C1417 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.022794f
C1418 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.076959f
C1419 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.022794f
C1420 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.022794f
C1421 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.082252f
C1422 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.022794f
C1423 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.022794f
C1424 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.081534f
C1425 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.302737f
C1426 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.022794f
C1427 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.022794f
C1428 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.081534f
C1429 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.157046f
C1430 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.022794f
C1431 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.022794f
C1432 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.081534f
C1433 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.157046f
C1434 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.022794f
C1435 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.022794f
C1436 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.082252f
C1437 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.191279f
C1438 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.123631f
C1439 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.031912f
C1440 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.031912f
C1441 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.031912f
C1442 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.031912f
C1443 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.031912f
C1444 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.031912f
C1445 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.031912f
C1446 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.03875f
C1447 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.03875f
C1448 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.025074f
C1449 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.025074f
C1450 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.025074f
C1451 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.025074f
C1452 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.025074f
C1453 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.022459f
C1454 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.031912f
C1455 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.03875f
C1456 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.036135f
C1457 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.022101f
C1458 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.049008f
C1459 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.049008f
C1460 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.049008f
C1461 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.049008f
C1462 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.049008f
C1463 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.049008f
C1464 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.049008f
C1465 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.055713f
C1466 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.05028f
C1467 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.030772f
C1468 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.030772f
C1469 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.030772f
C1470 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.030772f
C1471 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.030772f
C1472 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.028157f
C1473 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.049008f
C1474 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.055713f
C1475 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.047665f
C1476 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.022031f
C1477 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.153015f
C1478 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.741299f
C1479 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.100295f
C1480 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.100295f
C1481 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.106821f
C1482 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.084651f
C1483 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.045253f
C1484 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.100295f
C1485 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.100295f
C1486 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.100295f
C1487 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.100295f
C1488 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.100295f
C1489 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.100295f
C1490 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.106821f
C1491 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.084651f
C1492 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.047868f
C1493 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.047868f
C1494 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.047868f
C1495 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.047868f
C1496 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.045253f
C1497 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.024415f
C1498 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 1.03694f
C1499 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.458663f
C1500 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.183453f
C1501 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.028649f
C1502 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.028649f
C1503 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.084054f
C1504 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.028649f
C1505 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.028649f
C1506 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.083672f
C1507 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.28922f
C1508 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.028649f
C1509 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.028649f
C1510 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.083672f
C1511 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.149814f
C1512 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.028649f
C1513 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.028649f
C1514 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.083672f
C1515 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.149814f
C1516 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.028649f
C1517 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.028649f
C1518 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.083672f
C1519 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.215233f
C1520 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 1.07185f
C1521 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.014324f
C1522 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.014324f
C1523 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.035906f
C1524 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.014324f
C1525 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.014324f
C1526 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.035717f
C1527 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.31745f
C1528 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.014324f
C1529 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.014324f
C1530 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.028649f
C1531 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 0.173365f
C1532 bgr_0.V_CMFB_S1 GNDA 1.45835f
C1533 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.052601f
C1534 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.052601f
C1535 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.182935f
C1536 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.052601f
C1537 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.052601f
C1538 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.182287f
C1539 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.344139f
C1540 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.052601f
C1541 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.052601f
C1542 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.182287f
C1543 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.178405f
C1544 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.052601f
C1545 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.052601f
C1546 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.182287f
C1547 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.178405f
C1548 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.052601f
C1549 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.052601f
C1550 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.182287f
C1551 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.210076f
C1552 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.052601f
C1553 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.052601f
C1554 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.178511f
C1555 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.147505f
C1556 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.022543f
C1557 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.022543f
C1558 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.076111f
C1559 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.022543f
C1560 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.022543f
C1561 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.081346f
C1562 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.022543f
C1563 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.022543f
C1564 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.081346f
C1565 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.022543f
C1566 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.022543f
C1567 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.080636f
C1568 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.299403f
C1569 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.022543f
C1570 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.022543f
C1571 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.080636f
C1572 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.155317f
C1573 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.022543f
C1574 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.022543f
C1575 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.080636f
C1576 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.155317f
C1577 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.189173f
C1578 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.122269f
C1579 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.128676f
C1580 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.03156f
C1581 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.038324f
C1582 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.035737f
C1583 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.03156f
C1584 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.03156f
C1585 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.03156f
C1586 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.03156f
C1587 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.03156f
C1588 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.03156f
C1589 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.03156f
C1590 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.038324f
C1591 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.038324f
C1592 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.024798f
C1593 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.024798f
C1594 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.024798f
C1595 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.024798f
C1596 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.024798f
C1597 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.022211f
C1598 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.021857f
C1599 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.048468f
C1600 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.0551f
C1601 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.04714f
C1602 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.048468f
C1603 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.048468f
C1604 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.048468f
C1605 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.048468f
C1606 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.048468f
C1607 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.048468f
C1608 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.048468f
C1609 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.0551f
C1610 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.049726f
C1611 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.030433f
C1612 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.030433f
C1613 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.030433f
C1614 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.030433f
C1615 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.030433f
C1616 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.027847f
C1617 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.021789f
C1618 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.153028f
C1619 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.454714f
C1620 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.09919f
C1621 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.09919f
C1622 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.09919f
C1623 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.09919f
C1624 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.09919f
C1625 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.09919f
C1626 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.105644f
C1627 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.083719f
C1628 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.047341f
C1629 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.047341f
C1630 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.047341f
C1631 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.047341f
C1632 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.044755f
C1633 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.09919f
C1634 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.09919f
C1635 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.105644f
C1636 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.083719f
C1637 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.044755f
C1638 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.024251f
C1639 two_stage_opamp_dummy_magic_0.X.n52 GNDA 1.03308f
C1640 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.734227f
C1641 bgr_0.V_mir1.t9 GNDA 0.03537f
C1642 bgr_0.V_mir1.t5 GNDA 0.03537f
C1643 bgr_0.V_mir1.n0 GNDA 0.08097f
C1644 bgr_0.V_mir1.t8 GNDA 0.042444f
C1645 bgr_0.V_mir1.t18 GNDA 0.042444f
C1646 bgr_0.V_mir1.t17 GNDA 0.06851f
C1647 bgr_0.V_mir1.n1 GNDA 0.076506f
C1648 bgr_0.V_mir1.n2 GNDA 0.052264f
C1649 bgr_0.V_mir1.t4 GNDA 0.053881f
C1650 bgr_0.V_mir1.n3 GNDA 0.081315f
C1651 bgr_0.V_mir1.n4 GNDA 0.201563f
C1652 bgr_0.V_mir1.t7 GNDA 0.03537f
C1653 bgr_0.V_mir1.t3 GNDA 0.03537f
C1654 bgr_0.V_mir1.n5 GNDA 0.08097f
C1655 bgr_0.V_mir1.t6 GNDA 0.042444f
C1656 bgr_0.V_mir1.t20 GNDA 0.042444f
C1657 bgr_0.V_mir1.t22 GNDA 0.06851f
C1658 bgr_0.V_mir1.n6 GNDA 0.076506f
C1659 bgr_0.V_mir1.n7 GNDA 0.052264f
C1660 bgr_0.V_mir1.t2 GNDA 0.053881f
C1661 bgr_0.V_mir1.n8 GNDA 0.081315f
C1662 bgr_0.V_mir1.n9 GNDA 0.156007f
C1663 bgr_0.V_mir1.t1 GNDA 0.017685f
C1664 bgr_0.V_mir1.t15 GNDA 0.017685f
C1665 bgr_0.V_mir1.n10 GNDA 0.046242f
C1666 bgr_0.V_mir1.t14 GNDA 0.075466f
C1667 bgr_0.V_mir1.t16 GNDA 0.017685f
C1668 bgr_0.V_mir1.t0 GNDA 0.017685f
C1669 bgr_0.V_mir1.n11 GNDA 0.050199f
C1670 bgr_0.V_mir1.n12 GNDA 0.827814f
C1671 bgr_0.V_mir1.n13 GNDA 0.268286f
C1672 bgr_0.V_mir1.n14 GNDA 0.09373f
C1673 bgr_0.V_mir1.n15 GNDA 0.699157f
C1674 bgr_0.V_mir1.t12 GNDA 0.042444f
C1675 bgr_0.V_mir1.t21 GNDA 0.042444f
C1676 bgr_0.V_mir1.t19 GNDA 0.06851f
C1677 bgr_0.V_mir1.n16 GNDA 0.076506f
C1678 bgr_0.V_mir1.n17 GNDA 0.052264f
C1679 bgr_0.V_mir1.t10 GNDA 0.053881f
C1680 bgr_0.V_mir1.n18 GNDA 0.081315f
C1681 bgr_0.V_mir1.n19 GNDA 0.203577f
C1682 bgr_0.V_mir1.t11 GNDA 0.03537f
C1683 bgr_0.V_mir1.n20 GNDA 0.08097f
C1684 bgr_0.V_mir1.t13 GNDA 0.03537f
C1685 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 0.809844f
C1686 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 0.783855f
C1687 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 5.36727f
C1688 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.045982f
C1689 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.045982f
C1690 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.141876f
C1691 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.022991f
C1692 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.022991f
C1693 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.053263f
C1694 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.022991f
C1695 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.022991f
C1696 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.053319f
C1697 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.018968f
C1698 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.018968f
C1699 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.018968f
C1700 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.018968f
C1701 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.018968f
C1702 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.018968f
C1703 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.018968f
C1704 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.018968f
C1705 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.018968f
C1706 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.018968f
C1707 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.018968f
C1708 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.018968f
C1709 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.018968f
C1710 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.018968f
C1711 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.018968f
C1712 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.018968f
C1713 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.041097f
C1714 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.064088f
C1715 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.050006f
C1716 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.050006f
C1717 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.050006f
C1718 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.050006f
C1719 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.050006f
C1720 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.050006f
C1721 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.050006f
C1722 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.050006f
C1723 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.050006f
C1724 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.050006f
C1725 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.050006f
C1726 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.050006f
C1727 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.050006f
C1728 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.050006f
C1729 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.042791f
C1730 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.018968f
C1731 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.018968f
C1732 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.041097f
C1733 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.064088f
C1734 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.042791f
C1735 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.068952f
C1736 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.022991f
C1737 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.022991f
C1738 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.045982f
C1739 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.136971f
C1740 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.022991f
C1741 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.022991f
C1742 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.053319f
C1743 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.022991f
C1744 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.022991f
C1745 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.053319f
C1746 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.022991f
C1747 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.022991f
C1748 two_stage_opamp_dummy_magic_0.V_err_gate.n29 GNDA 0.053319f
C1749 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.047121f
C1750 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.014801f
C1751 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.027621f
C1752 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.065943f
C1753 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.412331f
C1754 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.014801f
C1755 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.027621f
C1756 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.065943f
C1757 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.380897f
C1758 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.04667f
C1759 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.370881f
C1760 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.014801f
C1761 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.027621f
C1762 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 0.065943f
C1763 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.230305f
C1764 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.014801f
C1765 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.027621f
C1766 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.065943f
C1767 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.357959f
C1768 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.080632f
C1769 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.030151f
C1770 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 0.09457f
C1771 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.030151f
C1772 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.077415f
C1773 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.030151f
C1774 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.077415f
C1775 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.030151f
C1776 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.118769f
C1777 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.769974f
C1778 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.097787f
C1779 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.097787f
C1780 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.327687f
C1781 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 3.69228f
C1782 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.097787f
C1783 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.097787f
C1784 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.327687f
C1785 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.884875f
C1786 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.097787f
C1787 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.097787f
C1788 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.327687f
C1789 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 1.26508f
C1790 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 1.10047f
C1791 bgr_0.cap_res2.t6 GNDA 0.406156f
C1792 bgr_0.cap_res2.t1 GNDA 0.407628f
C1793 bgr_0.cap_res2.t13 GNDA 0.406156f
C1794 bgr_0.cap_res2.t12 GNDA 0.407628f
C1795 bgr_0.cap_res2.t20 GNDA 0.406156f
C1796 bgr_0.cap_res2.t16 GNDA 0.407628f
C1797 bgr_0.cap_res2.t8 GNDA 0.406156f
C1798 bgr_0.cap_res2.t5 GNDA 0.407628f
C1799 bgr_0.cap_res2.t15 GNDA 0.406156f
C1800 bgr_0.cap_res2.t10 GNDA 0.407628f
C1801 bgr_0.cap_res2.t2 GNDA 0.406156f
C1802 bgr_0.cap_res2.t18 GNDA 0.407628f
C1803 bgr_0.cap_res2.t19 GNDA 0.406156f
C1804 bgr_0.cap_res2.t14 GNDA 0.407628f
C1805 bgr_0.cap_res2.t7 GNDA 0.406156f
C1806 bgr_0.cap_res2.t3 GNDA 0.407628f
C1807 bgr_0.cap_res2.n0 GNDA 0.272247f
C1808 bgr_0.cap_res2.t9 GNDA 0.216805f
C1809 bgr_0.cap_res2.n1 GNDA 0.295394f
C1810 bgr_0.cap_res2.t4 GNDA 0.216805f
C1811 bgr_0.cap_res2.n2 GNDA 0.295394f
C1812 bgr_0.cap_res2.t11 GNDA 0.216805f
C1813 bgr_0.cap_res2.n3 GNDA 0.295394f
C1814 bgr_0.cap_res2.t17 GNDA 0.846971f
C1815 bgr_0.cap_res2.t0 GNDA 0.133907f
C1816 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.344645f
C1817 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.167175f
C1818 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.198327f
C1819 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.344645f
C1820 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.167175f
C1821 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.216884f
C1822 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.344645f
C1823 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.167175f
C1824 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.216884f
C1825 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.344645f
C1826 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.167175f
C1827 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.216884f
C1828 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344645f
C1829 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.345795f
C1830 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.364353f
C1831 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.364353f
C1832 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.364353f
C1833 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.185733f
C1834 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.216884f
C1835 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344645f
C1836 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.345795f
C1837 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.364353f
C1838 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.364353f
C1839 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.364353f
C1840 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.185733f
C1841 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.216884f
C1842 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345795f
C1843 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.347048f
C1844 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345795f
C1845 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.348506f
C1846 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.37905f
C1847 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.345795f
C1848 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.347048f
C1849 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.345795f
C1850 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.347048f
C1851 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.345795f
C1852 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.347048f
C1853 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.345795f
C1854 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.347048f
C1855 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.345795f
C1856 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.347048f
C1857 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.345795f
C1858 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.347048f
C1859 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.345795f
C1860 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.347048f
C1861 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.345795f
C1862 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.347048f
C1863 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345795f
C1864 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.347048f
C1865 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.345795f
C1866 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.347048f
C1867 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.345795f
C1868 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.347048f
C1869 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.345795f
C1870 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.347048f
C1871 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.345795f
C1872 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.347048f
C1873 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.345795f
C1874 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.347048f
C1875 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.345795f
C1876 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.347048f
C1877 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.345795f
C1878 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.347048f
C1879 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.345795f
C1880 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.347048f
C1881 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.345795f
C1882 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.347048f
C1883 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.345795f
C1884 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.347048f
C1885 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.345795f
C1886 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.347048f
C1887 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.345795f
C1888 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.347048f
C1889 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.345795f
C1890 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.347048f
C1891 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.345795f
C1892 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.347048f
C1893 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.345795f
C1894 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.347048f
C1895 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.345795f
C1896 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.347048f
C1897 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.345795f
C1898 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.347048f
C1899 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.345795f
C1900 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.347048f
C1901 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.345795f
C1902 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.347048f
C1903 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.345795f
C1904 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.362749f
C1905 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.345795f
C1906 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.185733f
C1907 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.198781f
C1908 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.345795f
C1909 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.185733f
C1910 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.197177f
C1911 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.345795f
C1912 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.185733f
C1913 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.197177f
C1914 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.345795f
C1915 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.185733f
C1916 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.197177f
C1917 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.345795f
C1918 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185733f
C1919 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.197177f
C1920 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.345795f
C1921 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.185733f
C1922 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.197177f
C1923 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.345795f
C1924 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.185733f
C1925 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.197177f
C1926 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.345795f
C1927 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.185733f
C1928 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.197177f
C1929 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.345795f
C1930 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185733f
C1931 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.197177f
C1932 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.345795f
C1933 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.347048f
C1934 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.345795f
C1935 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.347048f
C1936 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.167175f
C1937 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.215631f
C1938 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.184584f
C1939 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.234189f
C1940 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.184584f
C1941 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.251494f
C1942 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.184584f
C1943 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.251494f
C1944 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.184584f
C1945 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.251494f
C1946 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.184584f
C1947 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.251494f
C1948 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.184584f
C1949 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.251494f
C1950 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.184584f
C1951 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.251494f
C1952 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.184584f
C1953 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.251494f
C1954 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.184584f
C1955 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.251494f
C1956 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.184584f
C1957 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.251494f
C1958 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.184584f
C1959 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.251494f
C1960 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.184584f
C1961 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.251494f
C1962 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.184584f
C1963 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.251494f
C1964 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.184584f
C1965 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.251494f
C1966 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.184584f
C1967 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.251494f
C1968 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.184584f
C1969 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.234189f
C1970 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.344645f
C1971 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.167175f
C1972 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216884f
C1973 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C1974 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.167175f
C1975 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216884f
C1976 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344645f
C1977 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.345795f
C1978 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.364353f
C1979 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.364353f
C1980 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.364353f
C1981 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185733f
C1982 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216884f
C1983 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.344645f
C1984 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216884f
C1985 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185733f
C1986 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.364353f
C1987 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.364353f
C1988 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.364353f
C1989 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.337351f
C1990 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.298183f
C1991 VOUT-.t18 GNDA 0.051003f
C1992 VOUT-.t8 GNDA 0.051003f
C1993 VOUT-.n0 GNDA 0.235943f
C1994 VOUT-.t6 GNDA 0.051003f
C1995 VOUT-.t13 GNDA 0.051003f
C1996 VOUT-.n1 GNDA 0.235153f
C1997 VOUT-.n2 GNDA 0.145313f
C1998 VOUT-.t14 GNDA 0.051003f
C1999 VOUT-.t17 GNDA 0.051003f
C2000 VOUT-.n3 GNDA 0.235153f
C2001 VOUT-.n4 GNDA 0.089445f
C2002 VOUT-.t4 GNDA 0.084326f
C2003 VOUT-.n5 GNDA 0.119504f
C2004 VOUT-.t0 GNDA 0.043717f
C2005 VOUT-.t11 GNDA 0.043717f
C2006 VOUT-.n6 GNDA 0.175711f
C2007 VOUT-.t2 GNDA 0.043717f
C2008 VOUT-.t1 GNDA 0.043717f
C2009 VOUT-.n7 GNDA 0.17571f
C2010 VOUT-.t9 GNDA 0.043717f
C2011 VOUT-.t10 GNDA 0.043717f
C2012 VOUT-.n8 GNDA 0.175387f
C2013 VOUT-.n9 GNDA 0.172777f
C2014 VOUT-.t5 GNDA 0.043717f
C2015 VOUT-.t7 GNDA 0.043717f
C2016 VOUT-.n10 GNDA 0.175387f
C2017 VOUT-.n11 GNDA 0.0891f
C2018 VOUT-.t16 GNDA 0.043717f
C2019 VOUT-.t3 GNDA 0.043717f
C2020 VOUT-.n12 GNDA 0.175387f
C2021 VOUT-.n13 GNDA 0.0891f
C2022 VOUT-.n14 GNDA 0.105535f
C2023 VOUT-.t15 GNDA 0.043717f
C2024 VOUT-.t12 GNDA 0.043717f
C2025 VOUT-.n15 GNDA 0.17324f
C2026 VOUT-.n16 GNDA 0.211953f
C2027 VOUT-.t100 GNDA 0.291446f
C2028 VOUT-.t107 GNDA 0.29641f
C2029 VOUT-.t149 GNDA 0.291446f
C2030 VOUT-.n17 GNDA 0.195405f
C2031 VOUT-.n18 GNDA 0.127508f
C2032 VOUT-.t47 GNDA 0.295788f
C2033 VOUT-.t91 GNDA 0.295788f
C2034 VOUT-.t41 GNDA 0.295788f
C2035 VOUT-.t130 GNDA 0.295788f
C2036 VOUT-.t82 GNDA 0.295788f
C2037 VOUT-.t124 GNDA 0.295788f
C2038 VOUT-.t72 GNDA 0.295788f
C2039 VOUT-.t23 GNDA 0.295788f
C2040 VOUT-.t62 GNDA 0.295788f
C2041 VOUT-.t150 GNDA 0.295788f
C2042 VOUT-.t86 GNDA 0.291446f
C2043 VOUT-.n19 GNDA 0.196026f
C2044 VOUT-.t50 GNDA 0.291446f
C2045 VOUT-.n20 GNDA 0.250673f
C2046 VOUT-.t137 GNDA 0.291446f
C2047 VOUT-.n21 GNDA 0.250673f
C2048 VOUT-.t105 GNDA 0.291446f
C2049 VOUT-.n22 GNDA 0.250673f
C2050 VOUT-.t73 GNDA 0.291446f
C2051 VOUT-.n23 GNDA 0.250673f
C2052 VOUT-.t25 GNDA 0.291446f
C2053 VOUT-.n24 GNDA 0.250673f
C2054 VOUT-.t127 GNDA 0.291446f
C2055 VOUT-.n25 GNDA 0.250673f
C2056 VOUT-.t88 GNDA 0.291446f
C2057 VOUT-.n26 GNDA 0.250673f
C2058 VOUT-.t53 GNDA 0.291446f
C2059 VOUT-.n27 GNDA 0.250673f
C2060 VOUT-.t140 GNDA 0.291446f
C2061 VOUT-.n28 GNDA 0.250673f
C2062 VOUT-.t109 GNDA 0.291446f
C2063 VOUT-.t28 GNDA 0.29641f
C2064 VOUT-.t78 GNDA 0.291446f
C2065 VOUT-.n29 GNDA 0.195405f
C2066 VOUT-.n30 GNDA 0.2368f
C2067 VOUT-.t24 GNDA 0.29641f
C2068 VOUT-.t112 GNDA 0.291446f
C2069 VOUT-.n31 GNDA 0.195405f
C2070 VOUT-.t77 GNDA 0.291446f
C2071 VOUT-.t129 GNDA 0.29641f
C2072 VOUT-.t37 GNDA 0.291446f
C2073 VOUT-.n32 GNDA 0.195405f
C2074 VOUT-.n33 GNDA 0.2368f
C2075 VOUT-.t59 GNDA 0.29641f
C2076 VOUT-.t147 GNDA 0.291446f
C2077 VOUT-.n34 GNDA 0.195405f
C2078 VOUT-.t116 GNDA 0.291446f
C2079 VOUT-.t32 GNDA 0.29641f
C2080 VOUT-.t81 GNDA 0.291446f
C2081 VOUT-.n35 GNDA 0.195405f
C2082 VOUT-.n36 GNDA 0.2368f
C2083 VOUT-.t99 GNDA 0.29641f
C2084 VOUT-.t46 GNDA 0.291446f
C2085 VOUT-.n37 GNDA 0.195405f
C2086 VOUT-.t153 GNDA 0.291446f
C2087 VOUT-.t69 GNDA 0.29641f
C2088 VOUT-.t122 GNDA 0.291446f
C2089 VOUT-.n38 GNDA 0.195405f
C2090 VOUT-.n39 GNDA 0.2368f
C2091 VOUT-.t67 GNDA 0.29641f
C2092 VOUT-.t154 GNDA 0.291446f
C2093 VOUT-.n40 GNDA 0.195405f
C2094 VOUT-.t123 GNDA 0.291446f
C2095 VOUT-.t35 GNDA 0.29641f
C2096 VOUT-.t84 GNDA 0.291446f
C2097 VOUT-.n41 GNDA 0.195405f
C2098 VOUT-.n42 GNDA 0.2368f
C2099 VOUT-.t104 GNDA 0.29641f
C2100 VOUT-.t52 GNDA 0.291446f
C2101 VOUT-.n43 GNDA 0.195405f
C2102 VOUT-.t22 GNDA 0.291446f
C2103 VOUT-.t76 GNDA 0.29641f
C2104 VOUT-.t126 GNDA 0.291446f
C2105 VOUT-.n44 GNDA 0.195405f
C2106 VOUT-.n45 GNDA 0.2368f
C2107 VOUT-.t95 GNDA 0.291446f
C2108 VOUT-.t83 GNDA 0.29641f
C2109 VOUT-.t56 GNDA 0.291446f
C2110 VOUT-.n46 GNDA 0.195405f
C2111 VOUT-.n47 GNDA 0.127508f
C2112 VOUT-.t132 GNDA 0.295788f
C2113 VOUT-.t114 GNDA 0.295788f
C2114 VOUT-.t90 GNDA 0.29641f
C2115 VOUT-.t131 GNDA 0.291446f
C2116 VOUT-.n48 GNDA 0.195405f
C2117 VOUT-.t103 GNDA 0.291446f
C2118 VOUT-.n49 GNDA 0.127508f
C2119 VOUT-.t71 GNDA 0.291446f
C2120 VOUT-.n50 GNDA 0.122954f
C2121 VOUT-.t146 GNDA 0.295788f
C2122 VOUT-.t128 GNDA 0.29641f
C2123 VOUT-.t31 GNDA 0.291446f
C2124 VOUT-.n51 GNDA 0.195405f
C2125 VOUT-.t138 GNDA 0.291446f
C2126 VOUT-.n52 GNDA 0.127508f
C2127 VOUT-.t106 GNDA 0.291446f
C2128 VOUT-.n53 GNDA 0.122954f
C2129 VOUT-.t45 GNDA 0.295788f
C2130 VOUT-.t26 GNDA 0.29641f
C2131 VOUT-.t60 GNDA 0.291446f
C2132 VOUT-.n54 GNDA 0.195405f
C2133 VOUT-.t40 GNDA 0.291446f
C2134 VOUT-.n55 GNDA 0.127508f
C2135 VOUT-.t143 GNDA 0.291446f
C2136 VOUT-.n56 GNDA 0.122954f
C2137 VOUT-.t85 GNDA 0.295788f
C2138 VOUT-.t74 GNDA 0.29641f
C2139 VOUT-.t113 GNDA 0.291446f
C2140 VOUT-.n57 GNDA 0.195405f
C2141 VOUT-.t21 GNDA 0.291446f
C2142 VOUT-.n58 GNDA 0.127508f
C2143 VOUT-.t125 GNDA 0.291446f
C2144 VOUT-.n59 GNDA 0.122954f
C2145 VOUT-.t63 GNDA 0.295788f
C2146 VOUT-.t101 GNDA 0.295788f
C2147 VOUT-.t134 GNDA 0.295788f
C2148 VOUT-.t119 GNDA 0.295788f
C2149 VOUT-.t155 GNDA 0.295788f
C2150 VOUT-.t118 GNDA 0.291446f
C2151 VOUT-.n60 GNDA 0.196026f
C2152 VOUT-.t80 GNDA 0.291446f
C2153 VOUT-.n61 GNDA 0.250673f
C2154 VOUT-.t96 GNDA 0.291446f
C2155 VOUT-.n62 GNDA 0.250673f
C2156 VOUT-.t61 GNDA 0.291446f
C2157 VOUT-.n63 GNDA 0.250673f
C2158 VOUT-.t27 GNDA 0.291446f
C2159 VOUT-.n64 GNDA 0.309873f
C2160 VOUT-.t44 GNDA 0.291446f
C2161 VOUT-.n65 GNDA 0.309873f
C2162 VOUT-.t144 GNDA 0.291446f
C2163 VOUT-.n66 GNDA 0.309873f
C2164 VOUT-.t111 GNDA 0.291446f
C2165 VOUT-.n67 GNDA 0.309873f
C2166 VOUT-.t75 GNDA 0.291446f
C2167 VOUT-.n68 GNDA 0.250673f
C2168 VOUT-.t92 GNDA 0.291446f
C2169 VOUT-.n69 GNDA 0.250673f
C2170 VOUT-.t55 GNDA 0.291446f
C2171 VOUT-.t39 GNDA 0.29641f
C2172 VOUT-.t19 GNDA 0.291446f
C2173 VOUT-.n70 GNDA 0.195405f
C2174 VOUT-.n71 GNDA 0.2368f
C2175 VOUT-.t34 GNDA 0.29641f
C2176 VOUT-.t51 GNDA 0.291446f
C2177 VOUT-.n72 GNDA 0.195405f
C2178 VOUT-.t156 GNDA 0.291446f
C2179 VOUT-.t136 GNDA 0.29641f
C2180 VOUT-.t120 GNDA 0.291446f
C2181 VOUT-.n73 GNDA 0.195405f
C2182 VOUT-.n74 GNDA 0.2368f
C2183 VOUT-.t68 GNDA 0.29641f
C2184 VOUT-.t87 GNDA 0.291446f
C2185 VOUT-.n75 GNDA 0.195405f
C2186 VOUT-.t49 GNDA 0.291446f
C2187 VOUT-.t36 GNDA 0.29641f
C2188 VOUT-.t151 GNDA 0.291446f
C2189 VOUT-.n76 GNDA 0.195405f
C2190 VOUT-.n77 GNDA 0.2368f
C2191 VOUT-.t94 GNDA 0.29641f
C2192 VOUT-.t42 GNDA 0.291446f
C2193 VOUT-.n78 GNDA 0.195405f
C2194 VOUT-.t145 GNDA 0.291446f
C2195 VOUT-.t64 GNDA 0.29641f
C2196 VOUT-.t117 GNDA 0.291446f
C2197 VOUT-.n79 GNDA 0.195405f
C2198 VOUT-.n80 GNDA 0.2368f
C2199 VOUT-.t54 GNDA 0.29641f
C2200 VOUT-.t141 GNDA 0.291446f
C2201 VOUT-.n81 GNDA 0.195405f
C2202 VOUT-.t110 GNDA 0.291446f
C2203 VOUT-.t29 GNDA 0.29641f
C2204 VOUT-.t79 GNDA 0.291446f
C2205 VOUT-.n82 GNDA 0.195405f
C2206 VOUT-.n83 GNDA 0.2368f
C2207 VOUT-.t89 GNDA 0.29641f
C2208 VOUT-.t38 GNDA 0.291446f
C2209 VOUT-.n84 GNDA 0.195405f
C2210 VOUT-.t139 GNDA 0.291446f
C2211 VOUT-.t57 GNDA 0.29641f
C2212 VOUT-.t108 GNDA 0.291446f
C2213 VOUT-.n85 GNDA 0.195405f
C2214 VOUT-.n86 GNDA 0.2368f
C2215 VOUT-.t48 GNDA 0.29641f
C2216 VOUT-.t135 GNDA 0.291446f
C2217 VOUT-.n87 GNDA 0.195405f
C2218 VOUT-.t102 GNDA 0.291446f
C2219 VOUT-.t20 GNDA 0.29641f
C2220 VOUT-.t70 GNDA 0.291446f
C2221 VOUT-.n88 GNDA 0.195405f
C2222 VOUT-.n89 GNDA 0.2368f
C2223 VOUT-.t148 GNDA 0.29641f
C2224 VOUT-.t98 GNDA 0.291446f
C2225 VOUT-.n90 GNDA 0.195405f
C2226 VOUT-.t66 GNDA 0.291446f
C2227 VOUT-.t121 GNDA 0.29641f
C2228 VOUT-.t33 GNDA 0.291446f
C2229 VOUT-.n91 GNDA 0.195405f
C2230 VOUT-.n92 GNDA 0.2368f
C2231 VOUT-.t43 GNDA 0.29641f
C2232 VOUT-.t133 GNDA 0.291446f
C2233 VOUT-.n93 GNDA 0.195405f
C2234 VOUT-.t97 GNDA 0.291446f
C2235 VOUT-.t152 GNDA 0.29641f
C2236 VOUT-.t65 GNDA 0.291446f
C2237 VOUT-.n94 GNDA 0.195405f
C2238 VOUT-.n95 GNDA 0.2368f
C2239 VOUT-.t115 GNDA 0.29641f
C2240 VOUT-.t30 GNDA 0.291446f
C2241 VOUT-.n96 GNDA 0.195405f
C2242 VOUT-.t58 GNDA 0.291446f
C2243 VOUT-.n97 GNDA 0.2368f
C2244 VOUT-.t93 GNDA 0.291446f
C2245 VOUT-.n98 GNDA 0.127508f
C2246 VOUT-.t142 GNDA 0.291446f
C2247 VOUT-.n99 GNDA 0.23878f
C2248 VOUT-.n100 GNDA 0.268998f
C2249 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2250 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2251 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2252 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2253 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2254 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2255 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2256 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2257 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2258 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2259 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2260 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2261 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2262 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2263 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2264 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2265 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2266 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2267 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2268 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2269 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.04969f
C2270 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.186051f
C2271 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2272 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2273 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.050131f
C2274 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2275 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2276 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2277 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.186051f
C2278 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.027755f
C2279 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2280 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2281 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2282 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2283 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2284 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2285 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2286 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2287 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2288 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2289 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2290 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2291 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.026104f
C2292 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.021692f
C2293 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.722672f
C2294 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.021546f
C2295 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.021546f
C2296 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.089099f
C2297 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.021546f
C2298 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.021546f
C2299 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.088757f
C2300 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.123062f
C2301 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.021546f
C2302 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.021546f
C2303 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.088757f
C2304 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.064216f
C2305 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.021546f
C2306 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.021546f
C2307 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.088757f
C2308 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.064216f
C2309 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.021546f
C2310 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.021546f
C2311 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.088757f
C2312 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.092294f
C2313 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.708017f
C2314 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.089418f
C2315 VDDA.t151 GNDA 0.019611f
C2316 VDDA.t411 GNDA 0.019611f
C2317 VDDA.n0 GNDA 0.081102f
C2318 VDDA.t396 GNDA 0.019611f
C2319 VDDA.t319 GNDA 0.019611f
C2320 VDDA.n1 GNDA 0.080791f
C2321 VDDA.n2 GNDA 0.112012f
C2322 VDDA.t397 GNDA 0.019611f
C2323 VDDA.t263 GNDA 0.019611f
C2324 VDDA.n3 GNDA 0.080791f
C2325 VDDA.n4 GNDA 0.05845f
C2326 VDDA.t393 GNDA 0.019611f
C2327 VDDA.t262 GNDA 0.019611f
C2328 VDDA.n5 GNDA 0.080791f
C2329 VDDA.n6 GNDA 0.05845f
C2330 VDDA.t392 GNDA 0.019611f
C2331 VDDA.t309 GNDA 0.019611f
C2332 VDDA.n7 GNDA 0.080791f
C2333 VDDA.n8 GNDA 0.05845f
C2334 VDDA.t409 GNDA 0.019611f
C2335 VDDA.t308 GNDA 0.019611f
C2336 VDDA.n9 GNDA 0.080791f
C2337 VDDA.n10 GNDA 0.168808f
C2338 VDDA.t270 GNDA 0.039223f
C2339 VDDA.t366 GNDA 0.039223f
C2340 VDDA.n11 GNDA 0.157356f
C2341 VDDA.n12 GNDA 0.079941f
C2342 VDDA.t91 GNDA 0.039072f
C2343 VDDA.n13 GNDA 0.052907f
C2344 VDDA.n14 GNDA 0.074679f
C2345 VDDA.t94 GNDA 0.043394f
C2346 VDDA.t92 GNDA 0.019003f
C2347 VDDA.n15 GNDA 0.068836f
C2348 VDDA.n16 GNDA 0.040523f
C2349 VDDA.t72 GNDA 0.043394f
C2350 VDDA.t70 GNDA 0.019003f
C2351 VDDA.n17 GNDA 0.068836f
C2352 VDDA.n18 GNDA 0.040523f
C2353 VDDA.n19 GNDA 0.043145f
C2354 VDDA.n20 GNDA 0.074679f
C2355 VDDA.n21 GNDA 0.21589f
C2356 VDDA.t71 GNDA 0.267373f
C2357 VDDA.t353 GNDA 0.154602f
C2358 VDDA.t457 GNDA 0.154602f
C2359 VDDA.t157 GNDA 0.154602f
C2360 VDDA.t433 GNDA 0.154602f
C2361 VDDA.t158 GNDA 0.115952f
C2362 VDDA.n22 GNDA 0.077301f
C2363 VDDA.t314 GNDA 0.115952f
C2364 VDDA.t463 GNDA 0.154602f
C2365 VDDA.t343 GNDA 0.154602f
C2366 VDDA.t367 GNDA 0.154602f
C2367 VDDA.t451 GNDA 0.154602f
C2368 VDDA.t93 GNDA 0.267373f
C2369 VDDA.n23 GNDA 0.21589f
C2370 VDDA.n24 GNDA 0.052907f
C2371 VDDA.n25 GNDA 0.100118f
C2372 VDDA.n26 GNDA 0.068517f
C2373 VDDA.n27 GNDA 0.101631f
C2374 VDDA.n28 GNDA 0.101631f
C2375 VDDA.n29 GNDA 0.100968f
C2376 VDDA.t63 GNDA 0.039072f
C2377 VDDA.t448 GNDA 0.039223f
C2378 VDDA.t199 GNDA 0.039223f
C2379 VDDA.n30 GNDA 0.157356f
C2380 VDDA.n31 GNDA 0.079941f
C2381 VDDA.t324 GNDA 0.039223f
C2382 VDDA.t278 GNDA 0.039223f
C2383 VDDA.n32 GNDA 0.157356f
C2384 VDDA.n33 GNDA 0.079941f
C2385 VDDA.t129 GNDA 0.039223f
C2386 VDDA.t316 GNDA 0.039223f
C2387 VDDA.n34 GNDA 0.157356f
C2388 VDDA.n35 GNDA 0.079941f
C2389 VDDA.t294 GNDA 0.039223f
C2390 VDDA.t462 GNDA 0.039223f
C2391 VDDA.n36 GNDA 0.157356f
C2392 VDDA.n37 GNDA 0.167984f
C2393 VDDA.n38 GNDA 0.126831f
C2394 VDDA.t61 GNDA 0.047409f
C2395 VDDA.n39 GNDA 0.090707f
C2396 VDDA.n40 GNDA 0.052994f
C2397 VDDA.n41 GNDA 0.079291f
C2398 VDDA.n42 GNDA 0.34901f
C2399 VDDA.t62 GNDA 0.539081f
C2400 VDDA.t293 GNDA 0.298419f
C2401 VDDA.t461 GNDA 0.298419f
C2402 VDDA.t128 GNDA 0.298419f
C2403 VDDA.t315 GNDA 0.298419f
C2404 VDDA.t323 GNDA 0.223814f
C2405 VDDA.n43 GNDA 0.149209f
C2406 VDDA.t277 GNDA 0.223814f
C2407 VDDA.t447 GNDA 0.298419f
C2408 VDDA.t198 GNDA 0.298419f
C2409 VDDA.t269 GNDA 0.298419f
C2410 VDDA.t365 GNDA 0.298419f
C2411 VDDA.t90 GNDA 0.539081f
C2412 VDDA.n44 GNDA 0.34901f
C2413 VDDA.n45 GNDA 0.079291f
C2414 VDDA.n46 GNDA 0.052994f
C2415 VDDA.t89 GNDA 0.047409f
C2416 VDDA.n47 GNDA 0.090707f
C2417 VDDA.n48 GNDA 0.126504f
C2418 VDDA.n49 GNDA 0.094908f
C2419 VDDA.t410 GNDA 0.019611f
C2420 VDDA.t339 GNDA 0.019611f
C2421 VDDA.n50 GNDA 0.081102f
C2422 VDDA.t167 GNDA 0.019611f
C2423 VDDA.t200 GNDA 0.019611f
C2424 VDDA.n51 GNDA 0.080791f
C2425 VDDA.n52 GNDA 0.112012f
C2426 VDDA.t265 GNDA 0.019611f
C2427 VDDA.t302 GNDA 0.019611f
C2428 VDDA.n53 GNDA 0.080791f
C2429 VDDA.n54 GNDA 0.05845f
C2430 VDDA.t452 GNDA 0.019611f
C2431 VDDA.t279 GNDA 0.019611f
C2432 VDDA.n55 GNDA 0.080791f
C2433 VDDA.n56 GNDA 0.05845f
C2434 VDDA.t276 GNDA 0.019611f
C2435 VDDA.t282 GNDA 0.019611f
C2436 VDDA.n57 GNDA 0.080791f
C2437 VDDA.n58 GNDA 0.05845f
C2438 VDDA.t381 GNDA 0.019611f
C2439 VDDA.t412 GNDA 0.019611f
C2440 VDDA.n59 GNDA 0.080791f
C2441 VDDA.n60 GNDA 0.201937f
C2442 VDDA.n61 GNDA 0.186636f
C2443 VDDA.t402 GNDA 0.02288f
C2444 VDDA.t336 GNDA 0.02288f
C2445 VDDA.n62 GNDA 0.079571f
C2446 VDDA.t378 GNDA 0.02288f
C2447 VDDA.t234 GNDA 0.02288f
C2448 VDDA.n63 GNDA 0.079289f
C2449 VDDA.n64 GNDA 0.149691f
C2450 VDDA.t338 GNDA 0.02288f
C2451 VDDA.t355 GNDA 0.02288f
C2452 VDDA.n65 GNDA 0.079571f
C2453 VDDA.t408 GNDA 0.02288f
C2454 VDDA.t143 GNDA 0.02288f
C2455 VDDA.n66 GNDA 0.079289f
C2456 VDDA.n67 GNDA 0.149691f
C2457 VDDA.n68 GNDA 0.020919f
C2458 VDDA.n69 GNDA 0.065136f
C2459 VDDA.n70 GNDA 0.088573f
C2460 VDDA.t97 GNDA 0.112871f
C2461 VDDA.t95 GNDA 0.039842f
C2462 VDDA.n71 GNDA 0.073634f
C2463 VDDA.n72 GNDA 0.047468f
C2464 VDDA.t9 GNDA 0.112871f
C2465 VDDA.t7 GNDA 0.039842f
C2466 VDDA.n73 GNDA 0.073634f
C2467 VDDA.n74 GNDA 0.047468f
C2468 VDDA.n75 GNDA 0.047067f
C2469 VDDA.n76 GNDA 0.088573f
C2470 VDDA.n77 GNDA 0.263962f
C2471 VDDA.t8 GNDA 0.394002f
C2472 VDDA.t401 GNDA 0.227491f
C2473 VDDA.t335 GNDA 0.227491f
C2474 VDDA.t377 GNDA 0.227491f
C2475 VDDA.t233 GNDA 0.227491f
C2476 VDDA.t333 GNDA 0.170618f
C2477 VDDA.n78 GNDA 0.113746f
C2478 VDDA.t194 GNDA 0.170618f
C2479 VDDA.t407 GNDA 0.227491f
C2480 VDDA.t142 GNDA 0.227491f
C2481 VDDA.t337 GNDA 0.227491f
C2482 VDDA.t354 GNDA 0.227491f
C2483 VDDA.t96 GNDA 0.394002f
C2484 VDDA.n79 GNDA 0.263962f
C2485 VDDA.n80 GNDA 0.065136f
C2486 VDDA.n81 GNDA 0.091188f
C2487 VDDA.t334 GNDA 0.02288f
C2488 VDDA.t195 GNDA 0.02288f
C2489 VDDA.n82 GNDA 0.074598f
C2490 VDDA.n83 GNDA 0.050914f
C2491 VDDA.n84 GNDA 0.0284f
C2492 VDDA.n85 GNDA 0.114109f
C2493 VDDA.t416 GNDA 0.02288f
C2494 VDDA.t145 GNDA 0.02288f
C2495 VDDA.n86 GNDA 0.079571f
C2496 VDDA.t127 GNDA 0.02288f
C2497 VDDA.t298 GNDA 0.02288f
C2498 VDDA.n87 GNDA 0.079289f
C2499 VDDA.n88 GNDA 0.149691f
C2500 VDDA.t197 GNDA 0.02288f
C2501 VDDA.t175 GNDA 0.02288f
C2502 VDDA.n89 GNDA 0.079571f
C2503 VDDA.t400 GNDA 0.02288f
C2504 VDDA.t217 GNDA 0.02288f
C2505 VDDA.n90 GNDA 0.079289f
C2506 VDDA.n91 GNDA 0.149691f
C2507 VDDA.n92 GNDA 0.020919f
C2508 VDDA.n93 GNDA 0.065136f
C2509 VDDA.n94 GNDA 0.088573f
C2510 VDDA.t24 GNDA 0.112871f
C2511 VDDA.t22 GNDA 0.039842f
C2512 VDDA.n95 GNDA 0.073634f
C2513 VDDA.n96 GNDA 0.047468f
C2514 VDDA.t115 GNDA 0.112871f
C2515 VDDA.t113 GNDA 0.039842f
C2516 VDDA.n97 GNDA 0.073634f
C2517 VDDA.n98 GNDA 0.047468f
C2518 VDDA.n99 GNDA 0.047067f
C2519 VDDA.n100 GNDA 0.088573f
C2520 VDDA.n101 GNDA 0.263962f
C2521 VDDA.t114 GNDA 0.394002f
C2522 VDDA.t415 GNDA 0.227491f
C2523 VDDA.t144 GNDA 0.227491f
C2524 VDDA.t126 GNDA 0.227491f
C2525 VDDA.t297 GNDA 0.227491f
C2526 VDDA.t429 GNDA 0.170618f
C2527 VDDA.n102 GNDA 0.113746f
C2528 VDDA.t184 GNDA 0.170618f
C2529 VDDA.t399 GNDA 0.227491f
C2530 VDDA.t216 GNDA 0.227491f
C2531 VDDA.t196 GNDA 0.227491f
C2532 VDDA.t174 GNDA 0.227491f
C2533 VDDA.t23 GNDA 0.394002f
C2534 VDDA.n103 GNDA 0.263962f
C2535 VDDA.n104 GNDA 0.065136f
C2536 VDDA.n105 GNDA 0.091188f
C2537 VDDA.t430 GNDA 0.02288f
C2538 VDDA.t185 GNDA 0.02288f
C2539 VDDA.n106 GNDA 0.074598f
C2540 VDDA.n107 GNDA 0.050914f
C2541 VDDA.n108 GNDA 0.0284f
C2542 VDDA.n109 GNDA 0.112148f
C2543 VDDA.t313 GNDA 0.039223f
C2544 VDDA.t395 GNDA 0.039223f
C2545 VDDA.n110 GNDA 0.157356f
C2546 VDDA.n111 GNDA 0.079941f
C2547 VDDA.t45 GNDA 0.039072f
C2548 VDDA.n112 GNDA 0.079291f
C2549 VDDA.n113 GNDA 0.052907f
C2550 VDDA.n114 GNDA 0.074679f
C2551 VDDA.t75 GNDA 0.043394f
C2552 VDDA.t73 GNDA 0.019003f
C2553 VDDA.n115 GNDA 0.068836f
C2554 VDDA.n116 GNDA 0.040523f
C2555 VDDA.t48 GNDA 0.043394f
C2556 VDDA.t46 GNDA 0.019003f
C2557 VDDA.n117 GNDA 0.068836f
C2558 VDDA.n118 GNDA 0.040523f
C2559 VDDA.n119 GNDA 0.043145f
C2560 VDDA.n120 GNDA 0.074679f
C2561 VDDA.n121 GNDA 0.21589f
C2562 VDDA.t47 GNDA 0.267373f
C2563 VDDA.t321 GNDA 0.154602f
C2564 VDDA.t398 GNDA 0.154602f
C2565 VDDA.t264 GNDA 0.154602f
C2566 VDDA.t404 GNDA 0.154602f
C2567 VDDA.t227 GNDA 0.115952f
C2568 VDDA.n122 GNDA 0.077301f
C2569 VDDA.t224 GNDA 0.115952f
C2570 VDDA.t150 GNDA 0.154602f
C2571 VDDA.t305 GNDA 0.154602f
C2572 VDDA.t320 GNDA 0.154602f
C2573 VDDA.t391 GNDA 0.154602f
C2574 VDDA.t74 GNDA 0.267373f
C2575 VDDA.n123 GNDA 0.21589f
C2576 VDDA.n124 GNDA 0.052907f
C2577 VDDA.n125 GNDA 0.100118f
C2578 VDDA.t60 GNDA 0.039072f
C2579 VDDA.t318 GNDA 0.039223f
C2580 VDDA.t406 GNDA 0.039223f
C2581 VDDA.n126 GNDA 0.157356f
C2582 VDDA.n127 GNDA 0.079941f
C2583 VDDA.t208 GNDA 0.039223f
C2584 VDDA.t226 GNDA 0.039223f
C2585 VDDA.n128 GNDA 0.157356f
C2586 VDDA.n129 GNDA 0.079941f
C2587 VDDA.t261 GNDA 0.039223f
C2588 VDDA.t307 GNDA 0.039223f
C2589 VDDA.n130 GNDA 0.157356f
C2590 VDDA.n131 GNDA 0.079941f
C2591 VDDA.t311 GNDA 0.039223f
C2592 VDDA.t206 GNDA 0.039223f
C2593 VDDA.n132 GNDA 0.157356f
C2594 VDDA.n133 GNDA 0.167984f
C2595 VDDA.n134 GNDA 0.126831f
C2596 VDDA.t58 GNDA 0.047409f
C2597 VDDA.n135 GNDA 0.090707f
C2598 VDDA.n136 GNDA 0.052994f
C2599 VDDA.n137 GNDA 0.34901f
C2600 VDDA.n138 GNDA 0.34901f
C2601 VDDA.t44 GNDA 0.539081f
C2602 VDDA.t312 GNDA 0.298419f
C2603 VDDA.t394 GNDA 0.298419f
C2604 VDDA.t317 GNDA 0.298419f
C2605 VDDA.t405 GNDA 0.298419f
C2606 VDDA.t207 GNDA 0.223814f
C2607 VDDA.n139 GNDA 0.079291f
C2608 VDDA.n140 GNDA 0.101631f
C2609 VDDA.n141 GNDA 0.101631f
C2610 VDDA.t59 GNDA 0.539081f
C2611 VDDA.t205 GNDA 0.298419f
C2612 VDDA.t310 GNDA 0.298419f
C2613 VDDA.t306 GNDA 0.298419f
C2614 VDDA.t260 GNDA 0.298419f
C2615 VDDA.t225 GNDA 0.223814f
C2616 VDDA.n142 GNDA 0.149209f
C2617 VDDA.n143 GNDA 0.100968f
C2618 VDDA.n144 GNDA 0.068517f
C2619 VDDA.n145 GNDA 0.052994f
C2620 VDDA.t43 GNDA 0.047409f
C2621 VDDA.n146 GNDA 0.090707f
C2622 VDDA.n147 GNDA 0.126504f
C2623 VDDA.n148 GNDA 0.096869f
C2624 VDDA.n149 GNDA 0.054258f
C2625 VDDA.n150 GNDA 0.183484f
C2626 VDDA.n151 GNDA 0.063328f
C2627 VDDA.n152 GNDA 0.169067f
C2628 VDDA.t21 GNDA 0.012318f
C2629 VDDA.n153 GNDA 0.026209f
C2630 VDDA.t121 GNDA 0.012318f
C2631 VDDA.n154 GNDA 0.026209f
C2632 VDDA.n155 GNDA 0.038055f
C2633 VDDA.n156 GNDA 0.063963f
C2634 VDDA.n157 GNDA 0.170463f
C2635 VDDA.t54 GNDA 0.012318f
C2636 VDDA.n158 GNDA 0.026209f
C2637 VDDA.t39 GNDA 0.012318f
C2638 VDDA.n159 GNDA 0.026209f
C2639 VDDA.n160 GNDA 0.035464f
C2640 VDDA.n161 GNDA 0.044022f
C2641 VDDA.n162 GNDA 0.170463f
C2642 VDDA.t38 GNDA 0.165828f
C2643 VDDA.t203 GNDA 0.102469f
C2644 VDDA.t403 GNDA 0.102469f
C2645 VDDA.t350 GNDA 0.102469f
C2646 VDDA.t267 GNDA 0.102469f
C2647 VDDA.t289 GNDA 0.076852f
C2648 VDDA.t53 GNDA 0.165828f
C2649 VDDA.t266 GNDA 0.102469f
C2650 VDDA.t202 GNDA 0.102469f
C2651 VDDA.t268 GNDA 0.102469f
C2652 VDDA.t235 GNDA 0.102469f
C2653 VDDA.t154 GNDA 0.076852f
C2654 VDDA.n163 GNDA 0.064597f
C2655 VDDA.n164 GNDA 0.051235f
C2656 VDDA.n165 GNDA 0.064597f
C2657 VDDA.n166 GNDA 0.043145f
C2658 VDDA.n167 GNDA 0.034908f
C2659 VDDA.n168 GNDA 0.081166f
C2660 VDDA.n169 GNDA 0.081166f
C2661 VDDA.n170 GNDA 0.169067f
C2662 VDDA.t120 GNDA 0.162484f
C2663 VDDA.t124 GNDA 0.100671f
C2664 VDDA.t273 GNDA 0.100671f
C2665 VDDA.t466 GNDA 0.100671f
C2666 VDDA.t201 GNDA 0.100671f
C2667 VDDA.t290 GNDA 0.075504f
C2668 VDDA.t20 GNDA 0.162484f
C2669 VDDA.t368 GNDA 0.100671f
C2670 VDDA.t125 GNDA 0.100671f
C2671 VDDA.t204 GNDA 0.100671f
C2672 VDDA.t322 GNDA 0.100671f
C2673 VDDA.t215 GNDA 0.075504f
C2674 VDDA.n171 GNDA 0.064597f
C2675 VDDA.n172 GNDA 0.050336f
C2676 VDDA.n173 GNDA 0.064597f
C2677 VDDA.n174 GNDA 0.042939f
C2678 VDDA.n175 GNDA 0.034908f
C2679 VDDA.n176 GNDA 0.067579f
C2680 VDDA.n177 GNDA 0.090398f
C2681 VDDA.n179 GNDA 0.050053f
C2682 VDDA.n180 GNDA 0.079099f
C2683 VDDA.n181 GNDA 0.100359f
C2684 VDDA.n182 GNDA 0.100359f
C2685 VDDA.n183 GNDA 0.100359f
C2686 VDDA.n185 GNDA 0.050053f
C2687 VDDA.n187 GNDA 0.050053f
C2688 VDDA.n189 GNDA 0.050053f
C2689 VDDA.n191 GNDA 0.050053f
C2690 VDDA.n193 GNDA 0.050053f
C2691 VDDA.n195 GNDA 0.050053f
C2692 VDDA.n197 GNDA 0.050053f
C2693 VDDA.n199 GNDA 0.050053f
C2694 VDDA.n201 GNDA 0.081907f
C2695 VDDA.t112 GNDA 0.01191f
C2696 VDDA.n202 GNDA 0.017684f
C2697 VDDA.n203 GNDA 0.015647f
C2698 VDDA.n204 GNDA 0.053441f
C2699 VDDA.n205 GNDA 0.062095f
C2700 VDDA.n206 GNDA 0.205213f
C2701 VDDA.t111 GNDA 0.162484f
C2702 VDDA.t331 GNDA 0.100671f
C2703 VDDA.t186 GNDA 0.100671f
C2704 VDDA.t180 GNDA 0.100671f
C2705 VDDA.t148 GNDA 0.100671f
C2706 VDDA.t178 GNDA 0.100671f
C2707 VDDA.t134 GNDA 0.100671f
C2708 VDDA.t327 GNDA 0.100671f
C2709 VDDA.t218 GNDA 0.100671f
C2710 VDDA.t140 GNDA 0.100671f
C2711 VDDA.t329 GNDA 0.075504f
C2712 VDDA.n207 GNDA 0.050336f
C2713 VDDA.t146 GNDA 0.075504f
C2714 VDDA.t220 GNDA 0.100671f
C2715 VDDA.t356 GNDA 0.100671f
C2716 VDDA.t176 GNDA 0.100671f
C2717 VDDA.t188 GNDA 0.100671f
C2718 VDDA.t325 GNDA 0.100671f
C2719 VDDA.t136 GNDA 0.100671f
C2720 VDDA.t138 GNDA 0.100671f
C2721 VDDA.t182 GNDA 0.100671f
C2722 VDDA.t358 GNDA 0.100671f
C2723 VDDA.t105 GNDA 0.162484f
C2724 VDDA.n208 GNDA 0.205213f
C2725 VDDA.n209 GNDA 0.062095f
C2726 VDDA.n210 GNDA 0.053441f
C2727 VDDA.n211 GNDA 0.015647f
C2728 VDDA.t106 GNDA 0.01191f
C2729 VDDA.n212 GNDA 0.017253f
C2730 VDDA.n213 GNDA 0.08583f
C2731 VDDA.n214 GNDA 0.079813f
C2732 VDDA.n216 GNDA 0.063787f
C2733 VDDA.n217 GNDA 0.011767f
C2734 VDDA.n218 GNDA 0.034758f
C2735 VDDA.n219 GNDA 0.034758f
C2736 VDDA.n220 GNDA 0.03544f
C2737 VDDA.n221 GNDA 0.089052f
C2738 VDDA.n222 GNDA 0.011767f
C2739 VDDA.n223 GNDA 0.052267f
C2740 VDDA.n224 GNDA 0.052267f
C2741 VDDA.n225 GNDA 0.052266f
C2742 VDDA.t173 GNDA 0.020919f
C2743 VDDA.n226 GNDA 0.072591f
C2744 VDDA.t18 GNDA 0.09555f
C2745 VDDA.n227 GNDA 0.047382f
C2746 VDDA.n228 GNDA 0.045486f
C2747 VDDA.t16 GNDA 0.036306f
C2748 VDDA.n229 GNDA 0.038438f
C2749 VDDA.n230 GNDA 0.028772f
C2750 VDDA.n231 GNDA 0.044706f
C2751 VDDA.n232 GNDA 0.29309f
C2752 VDDA.t17 GNDA 0.278605f
C2753 VDDA.n233 GNDA 0.090702f
C2754 VDDA.n234 GNDA 0.022676f
C2755 VDDA.t172 GNDA 0.126983f
C2756 VDDA.t32 GNDA 0.30128f
C2757 VDDA.n235 GNDA 0.296124f
C2758 VDDA.n236 GNDA 0.04639f
C2759 VDDA.n237 GNDA 0.029748f
C2760 VDDA.t31 GNDA 0.036959f
C2761 VDDA.n238 GNDA 0.038438f
C2762 VDDA.t33 GNDA 0.074631f
C2763 VDDA.n239 GNDA 0.051218f
C2764 VDDA.n240 GNDA 0.101927f
C2765 VDDA.n241 GNDA 0.067804f
C2766 VDDA.t51 GNDA 0.01528f
C2767 VDDA.n242 GNDA 0.0166f
C2768 VDDA.t49 GNDA 0.012819f
C2769 VDDA.n243 GNDA 0.01623f
C2770 VDDA.n244 GNDA 0.020897f
C2771 VDDA.n245 GNDA 0.029326f
C2772 VDDA.n246 GNDA 0.156422f
C2773 VDDA.t50 GNDA 0.173249f
C2774 VDDA.t375 GNDA 0.117668f
C2775 VDDA.t86 GNDA 0.173249f
C2776 VDDA.n247 GNDA 0.156422f
C2777 VDDA.n248 GNDA 0.029326f
C2778 VDDA.n249 GNDA 0.020897f
C2779 VDDA.t85 GNDA 0.012819f
C2780 VDDA.n250 GNDA 0.01623f
C2781 VDDA.t88 GNDA 0.01528f
C2782 VDDA.n251 GNDA 0.01853f
C2783 VDDA.n252 GNDA 0.063592f
C2784 VDDA.n253 GNDA 0.492776f
C2785 VDDA.t469 GNDA 0.722704f
C2786 VDDA.t472 GNDA 0.738614f
C2787 VDDA.t470 GNDA 0.770264f
C2788 VDDA.n254 GNDA 0.51631f
C2789 VDDA.t471 GNDA 0.770264f
C2790 VDDA.n255 GNDA 0.250668f
C2791 VDDA.n256 GNDA 0.321372f
C2792 VDDA.n257 GNDA 2.58933f
C2793 VDDA.n258 GNDA 0.020919f
C2794 VDDA.n259 GNDA 0.015833f
C2795 VDDA.n260 GNDA 0.032622f
C2796 VDDA.n261 GNDA 0.020919f
C2797 VDDA.n262 GNDA 0.020919f
C2798 VDDA.n263 GNDA 0.015833f
C2799 VDDA.n264 GNDA 0.015833f
C2800 VDDA.n265 GNDA 0.04627f
C2801 VDDA.n266 GNDA 0.020919f
C2802 VDDA.n267 GNDA 0.224058f
C2803 VDDA.n268 GNDA 0.224058f
C2804 VDDA.t65 GNDA 0.204359f
C2805 VDDA.t419 GNDA 0.129435f
C2806 VDDA.t242 GNDA 0.129435f
C2807 VDDA.t238 GNDA 0.129435f
C2808 VDDA.t258 GNDA 0.129435f
C2809 VDDA.t256 GNDA 0.129435f
C2810 VDDA.t427 GNDA 0.129435f
C2811 VDDA.t423 GNDA 0.129435f
C2812 VDDA.t254 GNDA 0.129435f
C2813 VDDA.t248 GNDA 0.097076f
C2814 VDDA.t66 GNDA 0.024557f
C2815 VDDA.t64 GNDA 0.016182f
C2816 VDDA.n269 GNDA 0.038524f
C2817 VDDA.n270 GNDA 0.054814f
C2818 VDDA.t109 GNDA 0.024557f
C2819 VDDA.t107 GNDA 0.016182f
C2820 VDDA.n271 GNDA 0.038524f
C2821 VDDA.n272 GNDA 0.020919f
C2822 VDDA.n273 GNDA 0.015833f
C2823 VDDA.n274 GNDA 0.015833f
C2824 VDDA.n275 GNDA 0.020919f
C2825 VDDA.n276 GNDA 0.04627f
C2826 VDDA.n277 GNDA 0.020919f
C2827 VDDA.n278 GNDA 0.015833f
C2828 VDDA.n279 GNDA 0.04627f
C2829 VDDA.n280 GNDA 0.020919f
C2830 VDDA.n281 GNDA 0.016554f
C2831 VDDA.n282 GNDA 0.016442f
C2832 VDDA.n283 GNDA 0.127816f
C2833 VDDA.n284 GNDA 0.016442f
C2834 VDDA.n285 GNDA 0.066579f
C2835 VDDA.n286 GNDA 0.016442f
C2836 VDDA.n287 GNDA 0.066579f
C2837 VDDA.n288 GNDA 0.064302f
C2838 VDDA.n289 GNDA 0.103049f
C2839 VDDA.t57 GNDA 0.024557f
C2840 VDDA.t55 GNDA 0.016182f
C2841 VDDA.n290 GNDA 0.038524f
C2842 VDDA.n291 GNDA 0.054814f
C2843 VDDA.t69 GNDA 0.024557f
C2844 VDDA.t67 GNDA 0.016182f
C2845 VDDA.n292 GNDA 0.038524f
C2846 VDDA.n293 GNDA 0.054814f
C2847 VDDA.n294 GNDA 0.078445f
C2848 VDDA.n295 GNDA 0.103049f
C2849 VDDA.n296 GNDA 0.224058f
C2850 VDDA.t68 GNDA 0.204359f
C2851 VDDA.t303 GNDA 0.129435f
C2852 VDDA.t436 GNDA 0.129435f
C2853 VDDA.t285 GNDA 0.129435f
C2854 VDDA.t222 GNDA 0.129435f
C2855 VDDA.t291 GNDA 0.129435f
C2856 VDDA.t3 GNDA 0.129435f
C2857 VDDA.t209 GNDA 0.129435f
C2858 VDDA.t434 GNDA 0.129435f
C2859 VDDA.t211 GNDA 0.097076f
C2860 VDDA.n297 GNDA 0.064717f
C2861 VDDA.t467 GNDA 0.097076f
C2862 VDDA.t431 GNDA 0.129435f
C2863 VDDA.t5 GNDA 0.129435f
C2864 VDDA.t280 GNDA 0.129435f
C2865 VDDA.t287 GNDA 0.129435f
C2866 VDDA.t213 GNDA 0.129435f
C2867 VDDA.t168 GNDA 0.129435f
C2868 VDDA.t387 GNDA 0.129435f
C2869 VDDA.t271 GNDA 0.129435f
C2870 VDDA.t56 GNDA 0.204359f
C2871 VDDA.n298 GNDA 0.224058f
C2872 VDDA.n299 GNDA 0.064302f
C2873 VDDA.n300 GNDA 0.109541f
C2874 VDDA.n301 GNDA 0.015833f
C2875 VDDA.n302 GNDA 0.04627f
C2876 VDDA.n303 GNDA 0.020919f
C2877 VDDA.n304 GNDA 0.016442f
C2878 VDDA.n305 GNDA 0.066579f
C2879 VDDA.n306 GNDA 0.016442f
C2880 VDDA.n307 GNDA 0.066579f
C2881 VDDA.n308 GNDA 0.016442f
C2882 VDDA.n309 GNDA 0.066579f
C2883 VDDA.n310 GNDA 0.016442f
C2884 VDDA.n311 GNDA 0.095342f
C2885 VDDA.n312 GNDA 0.049682f
C2886 VDDA.n313 GNDA 0.04627f
C2887 VDDA.n314 GNDA 0.034154f
C2888 VDDA.n315 GNDA 0.032622f
C2889 VDDA.n316 GNDA 0.054814f
C2890 VDDA.n317 GNDA 0.078445f
C2891 VDDA.n318 GNDA 0.103049f
C2892 VDDA.t108 GNDA 0.204359f
C2893 VDDA.t417 GNDA 0.129435f
C2894 VDDA.t244 GNDA 0.129435f
C2895 VDDA.t250 GNDA 0.129435f
C2896 VDDA.t246 GNDA 0.129435f
C2897 VDDA.t252 GNDA 0.129435f
C2898 VDDA.t421 GNDA 0.129435f
C2899 VDDA.t425 GNDA 0.129435f
C2900 VDDA.t236 GNDA 0.129435f
C2901 VDDA.t240 GNDA 0.097076f
C2902 VDDA.n319 GNDA 0.064717f
C2903 VDDA.n320 GNDA 0.103049f
C2904 VDDA.n321 GNDA 0.020919f
C2905 VDDA.n322 GNDA 0.04627f
C2906 VDDA.n323 GNDA 0.020919f
C2907 VDDA.n324 GNDA 0.015833f
C2908 VDDA.n325 GNDA 0.04627f
C2909 VDDA.n326 GNDA 0.020919f
C2910 VDDA.n327 GNDA 0.020919f
C2911 VDDA.n328 GNDA 0.015833f
C2912 VDDA.n329 GNDA 0.04627f
C2913 VDDA.n330 GNDA 0.020919f
C2914 VDDA.n331 GNDA 0.015833f
C2915 VDDA.n332 GNDA 0.04627f
C2916 VDDA.n333 GNDA 0.020919f
C2917 VDDA.n334 GNDA 0.034154f
C2918 VDDA.n335 GNDA 0.04627f
C2919 VDDA.n336 GNDA 0.063329f
C2920 VDDA.n337 GNDA 0.192271f
C2921 VDDA.t346 GNDA 0.019611f
C2922 VDDA.t454 GNDA 0.019611f
C2923 VDDA.n338 GNDA 0.06479f
C2924 VDDA.n339 GNDA 0.083603f
C2925 VDDA.n340 GNDA 0.091848f
C2926 VDDA.t79 GNDA 0.093515f
C2927 VDDA.t81 GNDA 0.060101f
C2928 VDDA.t166 GNDA 0.019611f
C2929 VDDA.t349 GNDA 0.019611f
C2930 VDDA.n341 GNDA 0.06479f
C2931 VDDA.n342 GNDA 0.083603f
C2932 VDDA.t363 GNDA 0.019611f
C2933 VDDA.t460 GNDA 0.019611f
C2934 VDDA.n343 GNDA 0.06479f
C2935 VDDA.n344 GNDA 0.083603f
C2936 VDDA.t300 GNDA 0.019611f
C2937 VDDA.t342 GNDA 0.019611f
C2938 VDDA.n345 GNDA 0.06479f
C2939 VDDA.n346 GNDA 0.083603f
C2940 VDDA.t160 GNDA 0.019611f
C2941 VDDA.t1 GNDA 0.019611f
C2942 VDDA.n347 GNDA 0.06479f
C2943 VDDA.n348 GNDA 0.083603f
C2944 VDDA.t229 GNDA 0.019611f
C2945 VDDA.t164 GNDA 0.019611f
C2946 VDDA.n349 GNDA 0.06479f
C2947 VDDA.n350 GNDA 0.083603f
C2948 VDDA.t162 GNDA 0.019611f
C2949 VDDA.t443 GNDA 0.019611f
C2950 VDDA.n351 GNDA 0.06479f
C2951 VDDA.n352 GNDA 0.083603f
C2952 VDDA.t384 GNDA 0.019611f
C2953 VDDA.t456 GNDA 0.019611f
C2954 VDDA.n353 GNDA 0.06479f
C2955 VDDA.n354 GNDA 0.083603f
C2956 VDDA.t12 GNDA 0.024557f
C2957 VDDA.t10 GNDA 0.012393f
C2958 VDDA.n355 GNDA 0.038717f
C2959 VDDA.n356 GNDA 0.022325f
C2960 VDDA.n357 GNDA 0.039677f
C2961 VDDA.t42 GNDA 0.024557f
C2962 VDDA.t40 GNDA 0.012393f
C2963 VDDA.n358 GNDA 0.038717f
C2964 VDDA.n359 GNDA 0.039677f
C2965 VDDA.n360 GNDA 0.039677f
C2966 VDDA.n361 GNDA 0.032556f
C2967 VDDA.n362 GNDA 0.16433f
C2968 VDDA.t11 GNDA 0.199332f
C2969 VDDA.t464 GNDA 0.088986f
C2970 VDDA.n363 GNDA 0.059324f
C2971 VDDA.t465 GNDA 0.088986f
C2972 VDDA.t41 GNDA 0.196435f
C2973 VDDA.n364 GNDA 0.156441f
C2974 VDDA.n365 GNDA 0.032556f
C2975 VDDA.n366 GNDA 0.022325f
C2976 VDDA.n367 GNDA 0.031364f
C2977 VDDA.n368 GNDA 0.092307f
C2978 VDDA.n369 GNDA 0.111606f
C2979 VDDA.n370 GNDA 0.075228f
C2980 VDDA.n371 GNDA 0.338416f
C2981 VDDA.n372 GNDA 0.338416f
C2982 VDDA.t83 GNDA 0.436669f
C2983 VDDA.t345 GNDA 0.314762f
C2984 VDDA.t453 GNDA 0.314762f
C2985 VDDA.t165 GNDA 0.314762f
C2986 VDDA.t348 GNDA 0.314762f
C2987 VDDA.t362 GNDA 0.314762f
C2988 VDDA.t459 GNDA 0.314762f
C2989 VDDA.t299 GNDA 0.314762f
C2990 VDDA.t341 GNDA 0.236071f
C2991 VDDA.n373 GNDA 0.091848f
C2992 VDDA.n374 GNDA 0.144363f
C2993 VDDA.n375 GNDA 0.144363f
C2994 VDDA.t80 GNDA 0.436669f
C2995 VDDA.t455 GNDA 0.314762f
C2996 VDDA.t383 GNDA 0.314762f
C2997 VDDA.t442 GNDA 0.314762f
C2998 VDDA.t161 GNDA 0.314762f
C2999 VDDA.t163 GNDA 0.314762f
C3000 VDDA.t228 GNDA 0.314762f
C3001 VDDA.t0 GNDA 0.314762f
C3002 VDDA.t159 GNDA 0.236071f
C3003 VDDA.n376 GNDA 0.157381f
C3004 VDDA.n377 GNDA 0.1437f
C3005 VDDA.n378 GNDA 0.105901f
C3006 VDDA.n379 GNDA 0.075228f
C3007 VDDA.t84 GNDA 0.060101f
C3008 VDDA.t82 GNDA 0.093515f
C3009 VDDA.n380 GNDA 0.111606f
C3010 VDDA.n381 GNDA 0.051232f
C3011 VDDA.t100 GNDA 0.024739f
C3012 VDDA.t98 GNDA 0.012072f
C3013 VDDA.n382 GNDA 0.037058f
C3014 VDDA.n383 GNDA 0.022222f
C3015 VDDA.n384 GNDA 0.039677f
C3016 VDDA.t30 GNDA 0.024739f
C3017 VDDA.t28 GNDA 0.012072f
C3018 VDDA.n385 GNDA 0.037058f
C3019 VDDA.n386 GNDA 0.039677f
C3020 VDDA.n387 GNDA 0.039677f
C3021 VDDA.n388 GNDA 0.032556f
C3022 VDDA.n389 GNDA 0.156441f
C3023 VDDA.t99 GNDA 0.196435f
C3024 VDDA.t155 GNDA 0.088986f
C3025 VDDA.n390 GNDA 0.059324f
C3026 VDDA.t379 GNDA 0.088986f
C3027 VDDA.t29 GNDA 0.196435f
C3028 VDDA.n391 GNDA 0.156441f
C3029 VDDA.n392 GNDA 0.032556f
C3030 VDDA.n393 GNDA 0.022222f
C3031 VDDA.n394 GNDA 0.023347f
C3032 VDDA.n395 GNDA 0.015788f
C3033 VDDA.n396 GNDA 0.0437f
C3034 VDDA.n397 GNDA 0.09207f
C3035 VDDA.n398 GNDA 0.159877f
C3036 VDDA.n399 GNDA 0.016307f
C3037 VDDA.n400 GNDA 0.057562f
C3038 VDDA.n401 GNDA 0.036738f
C3039 VDDA.t116 GNDA 0.012874f
C3040 VDDA.t118 GNDA 0.025799f
C3041 VDDA.n402 GNDA 0.016307f
C3042 VDDA.n403 GNDA 0.057562f
C3043 VDDA.n404 GNDA 0.016277f
C3044 VDDA.n405 GNDA 0.057593f
C3045 VDDA.n406 GNDA 0.043541f
C3046 VDDA.t13 GNDA 0.012874f
C3047 VDDA.t15 GNDA 0.02462f
C3048 VDDA.n407 GNDA 0.016277f
C3049 VDDA.n408 GNDA 0.057593f
C3050 VDDA.n409 GNDA 0.016277f
C3051 VDDA.n410 GNDA 0.057593f
C3052 VDDA.n411 GNDA 0.016277f
C3053 VDDA.n412 GNDA 0.057593f
C3054 VDDA.n413 GNDA 0.016277f
C3055 VDDA.n414 GNDA 0.057593f
C3056 VDDA.n415 GNDA 0.016314f
C3057 VDDA.n416 GNDA 0.057556f
C3058 VDDA.n417 GNDA 0.036238f
C3059 VDDA.t34 GNDA 0.012874f
C3060 VDDA.t36 GNDA 0.025809f
C3061 VDDA.n418 GNDA 0.016314f
C3062 VDDA.n419 GNDA 0.078775f
C3063 VDDA.n420 GNDA 0.044201f
C3064 VDDA.n421 GNDA 0.026378f
C3065 VDDA.n422 GNDA 0.16509f
C3066 VDDA.n423 GNDA 0.16509f
C3067 VDDA.t102 GNDA 0.19989f
C3068 VDDA.t389 GNDA 0.120446f
C3069 VDDA.t438 GNDA 0.090335f
C3070 VDDA.n424 GNDA 0.036238f
C3071 VDDA.n425 GNDA 0.046694f
C3072 VDDA.n426 GNDA 0.046694f
C3073 VDDA.t35 GNDA 0.19989f
C3074 VDDA.t440 GNDA 0.120446f
C3075 VDDA.t274 GNDA 0.090335f
C3076 VDDA.n427 GNDA 0.060223f
C3077 VDDA.n428 GNDA 0.046694f
C3078 VDDA.n429 GNDA 0.021572f
C3079 VDDA.n430 GNDA 0.026378f
C3080 VDDA.t103 GNDA 0.025809f
C3081 VDDA.t101 GNDA 0.013282f
C3082 VDDA.n431 GNDA 0.043745f
C3083 VDDA.n432 GNDA 0.039734f
C3084 VDDA.n433 GNDA 0.039734f
C3085 VDDA.n434 GNDA 0.044526f
C3086 VDDA.n435 GNDA 0.04076f
C3087 VDDA.n436 GNDA 0.179695f
C3088 VDDA.n437 GNDA 0.194214f
C3089 VDDA.t77 GNDA 0.19989f
C3090 VDDA.t132 GNDA 0.120446f
C3091 VDDA.t371 GNDA 0.120446f
C3092 VDDA.t170 GNDA 0.120446f
C3093 VDDA.t130 GNDA 0.090335f
C3094 VDDA.n438 GNDA 0.0508f
C3095 VDDA.n439 GNDA 0.067974f
C3096 VDDA.n440 GNDA 0.067974f
C3097 VDDA.t14 GNDA 0.19989f
C3098 VDDA.t190 GNDA 0.120446f
C3099 VDDA.t373 GNDA 0.120446f
C3100 VDDA.t413 GNDA 0.120446f
C3101 VDDA.t192 GNDA 0.120446f
C3102 VDDA.t152 GNDA 0.120446f
C3103 VDDA.t283 GNDA 0.090335f
C3104 VDDA.n441 GNDA 0.060223f
C3105 VDDA.n442 GNDA 0.067974f
C3106 VDDA.n443 GNDA 0.043145f
C3107 VDDA.n444 GNDA 0.033569f
C3108 VDDA.t78 GNDA 0.02462f
C3109 VDDA.t76 GNDA 0.012874f
C3110 VDDA.n445 GNDA 0.044526f
C3111 VDDA.n446 GNDA 0.046925f
C3112 VDDA.n447 GNDA 0.046925f
C3113 VDDA.n448 GNDA 0.043347f
C3114 VDDA.n449 GNDA 0.026378f
C3115 VDDA.n450 GNDA 0.164306f
C3116 VDDA.n451 GNDA 0.163305f
C3117 VDDA.t26 GNDA 0.196435f
C3118 VDDA.t369 GNDA 0.118648f
C3119 VDDA.t351 GNDA 0.088986f
C3120 VDDA.t117 GNDA 0.196435f
C3121 VDDA.t449 GNDA 0.118648f
C3122 VDDA.t122 GNDA 0.080897f
C3123 VDDA.n452 GNDA 0.035737f
C3124 VDDA.n453 GNDA 0.046694f
C3125 VDDA.n454 GNDA 0.046694f
C3126 VDDA.n455 GNDA 0.029662f
C3127 VDDA.n456 GNDA 0.037752f
C3128 VDDA.n457 GNDA 0.046694f
C3129 VDDA.n458 GNDA 0.021572f
C3130 VDDA.n459 GNDA 0.026378f
C3131 VDDA.t27 GNDA 0.025799f
C3132 VDDA.t25 GNDA 0.012874f
C3133 VDDA.n460 GNDA 0.043347f
C3134 VDDA.n461 GNDA 0.086457f
C3135 VDDA.n462 GNDA 0.129779f
C3136 VDDA.t445 GNDA 0.365424f
C3137 VDDA.t232 GNDA 0.366748f
C3138 VDDA.t444 GNDA 0.365424f
C3139 VDDA.t385 GNDA 0.366748f
C3140 VDDA.t347 GNDA 0.365424f
C3141 VDDA.t2 GNDA 0.366748f
C3142 VDDA.t295 GNDA 0.365424f
C3143 VDDA.t230 GNDA 0.366748f
C3144 VDDA.t360 GNDA 0.365424f
C3145 VDDA.t458 GNDA 0.366748f
C3146 VDDA.t231 GNDA 0.365424f
C3147 VDDA.t296 GNDA 0.366748f
C3148 VDDA.t340 GNDA 0.365424f
C3149 VDDA.t361 GNDA 0.366748f
C3150 VDDA.t301 GNDA 0.365424f
C3151 VDDA.t382 GNDA 0.366748f
C3152 VDDA.n463 GNDA 0.244944f
C3153 VDDA.t364 GNDA 0.195062f
C3154 VDDA.n464 GNDA 0.26577f
C3155 VDDA.t344 GNDA 0.195062f
C3156 VDDA.n465 GNDA 0.26577f
C3157 VDDA.t386 GNDA 0.195062f
C3158 VDDA.n466 GNDA 0.26577f
C3159 VDDA.t446 GNDA 0.291072f
C3160 VDDA.n467 GNDA 0.457313f
C3161 VDDA.n468 GNDA 3.08441f
C3162 bgr_0.1st_Vout_2.n0 GNDA 0.706398f
C3163 bgr_0.1st_Vout_2.n1 GNDA 1.47663f
C3164 bgr_0.1st_Vout_2.n2 GNDA 2.04197f
C3165 bgr_0.1st_Vout_2.n3 GNDA 0.129733f
C3166 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C3167 bgr_0.1st_Vout_2.t12 GNDA 0.364565f
C3168 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C3169 bgr_0.1st_Vout_2.t27 GNDA 0.358459f
C3170 bgr_0.1st_Vout_2.t29 GNDA 0.364565f
C3171 bgr_0.1st_Vout_2.t34 GNDA 0.358459f
C3172 bgr_0.1st_Vout_2.t20 GNDA 0.364565f
C3173 bgr_0.1st_Vout_2.t26 GNDA 0.358459f
C3174 bgr_0.1st_Vout_2.t33 GNDA 0.358459f
C3175 bgr_0.1st_Vout_2.t35 GNDA 0.364565f
C3176 bgr_0.1st_Vout_2.t15 GNDA 0.358459f
C3177 bgr_0.1st_Vout_2.t11 GNDA 0.364565f
C3178 bgr_0.1st_Vout_2.t19 GNDA 0.358459f
C3179 bgr_0.1st_Vout_2.t25 GNDA 0.358459f
C3180 bgr_0.1st_Vout_2.t28 GNDA 0.364565f
C3181 bgr_0.1st_Vout_2.t32 GNDA 0.358459f
C3182 bgr_0.1st_Vout_2.t22 GNDA 0.364565f
C3183 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C3184 bgr_0.1st_Vout_2.t17 GNDA 0.358459f
C3185 bgr_0.1st_Vout_2.t36 GNDA 0.358459f
C3186 bgr_0.1st_Vout_2.t23 GNDA 0.023417f
C3187 bgr_0.1st_Vout_2.n4 GNDA 0.02259f
C3188 bgr_0.1st_Vout_2.t13 GNDA 0.013652f
C3189 bgr_0.1st_Vout_2.t16 GNDA 0.013652f
C3190 bgr_0.1st_Vout_2.n5 GNDA 0.03037f
C3191 bgr_0.1st_Vout_2.n6 GNDA 0.021654f
C3192 bgr_0.1st_Vout_2.t10 GNDA 0.018875f
C3193 bgr_0.1st_Vout_2.n7 GNDA 0.012945f
C3194 bgr_0.1st_Vout_2.n8 GNDA 0.195802f
C3195 bgr_0.1st_Vout_2.n9 GNDA 0.011712f
C3196 bgr_0.1st_Vout_2.t14 GNDA 0.013652f
C3197 bgr_0.1st_Vout_2.t18 GNDA 0.013652f
C3198 bgr_0.1st_Vout_2.n10 GNDA 0.03037f
C3199 bgr_0.1st_Vout_2.n11 GNDA 0.02259f
C3200 bgr_0.1st_Vout_2.t31 GNDA 0.021427f
C3201 bgr_0.V_mir2.n0 GNDA 0.362016f
C3202 bgr_0.V_mir2.t9 GNDA 0.03537f
C3203 bgr_0.V_mir2.t7 GNDA 0.03537f
C3204 bgr_0.V_mir2.t13 GNDA 0.03537f
C3205 bgr_0.V_mir2.n1 GNDA 0.08097f
C3206 bgr_0.V_mir2.t6 GNDA 0.053881f
C3207 bgr_0.V_mir2.t12 GNDA 0.042444f
C3208 bgr_0.V_mir2.t17 GNDA 0.042444f
C3209 bgr_0.V_mir2.t18 GNDA 0.06851f
C3210 bgr_0.V_mir2.n2 GNDA 0.076506f
C3211 bgr_0.V_mir2.n3 GNDA 0.052264f
C3212 bgr_0.V_mir2.n4 GNDA 0.081315f
C3213 bgr_0.V_mir2.n5 GNDA 0.203577f
C3214 bgr_0.V_mir2.t15 GNDA 0.03537f
C3215 bgr_0.V_mir2.t11 GNDA 0.03537f
C3216 bgr_0.V_mir2.n6 GNDA 0.08097f
C3217 bgr_0.V_mir2.t14 GNDA 0.053881f
C3218 bgr_0.V_mir2.t10 GNDA 0.042444f
C3219 bgr_0.V_mir2.t21 GNDA 0.042444f
C3220 bgr_0.V_mir2.t22 GNDA 0.06851f
C3221 bgr_0.V_mir2.n7 GNDA 0.076506f
C3222 bgr_0.V_mir2.n8 GNDA 0.052264f
C3223 bgr_0.V_mir2.n9 GNDA 0.081315f
C3224 bgr_0.V_mir2.n10 GNDA 0.156007f
C3225 bgr_0.V_mir2.t0 GNDA 0.017685f
C3226 bgr_0.V_mir2.t16 GNDA 0.017685f
C3227 bgr_0.V_mir2.n11 GNDA 0.046242f
C3228 bgr_0.V_mir2.t1 GNDA 0.075466f
C3229 bgr_0.V_mir2.t2 GNDA 0.017685f
C3230 bgr_0.V_mir2.t3 GNDA 0.017685f
C3231 bgr_0.V_mir2.n12 GNDA 0.050199f
C3232 bgr_0.V_mir2.n13 GNDA 0.827814f
C3233 bgr_0.V_mir2.n14 GNDA 0.699157f
C3234 bgr_0.V_mir2.t8 GNDA 0.053881f
C3235 bgr_0.V_mir2.t4 GNDA 0.042444f
C3236 bgr_0.V_mir2.t19 GNDA 0.042444f
C3237 bgr_0.V_mir2.t20 GNDA 0.06851f
C3238 bgr_0.V_mir2.n15 GNDA 0.076506f
C3239 bgr_0.V_mir2.n16 GNDA 0.052264f
C3240 bgr_0.V_mir2.n17 GNDA 0.081315f
C3241 bgr_0.V_mir2.n18 GNDA 0.201563f
C3242 bgr_0.V_mir2.n19 GNDA 0.08097f
C3243 bgr_0.V_mir2.t5 GNDA 0.03537f
C3244 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.081131f
C3245 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.012679f
C3246 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.012679f
C3247 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.0372f
C3248 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.012679f
C3249 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.012679f
C3250 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.037031f
C3251 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.128001f
C3252 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.012679f
C3253 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.012679f
C3254 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.037031f
C3255 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.066304f
C3256 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.012679f
C3257 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.012679f
C3258 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.037031f
C3259 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.066304f
C3260 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.012679f
C3261 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.012679f
C3262 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.037031f
C3263 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.095712f
C3264 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.706057f
C3265 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.015898f
C3266 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.015814f
C3267 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.107124f
C3268 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.015814f
C3269 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 0.11603f
C3270 bgr_0.V_CMFB_S3 GNDA 0.635658f
.ends

