magic
tech sky130A
timestamp 1752660866
<< nwell >>
rect -30 2305 310 2695
rect 440 2305 780 2525
rect 910 2305 1250 2695
rect 1380 2305 1720 2695
rect -1225 1730 -345 2120
rect -100 1730 780 2120
rect 910 1730 1790 2120
rect 2035 1730 2915 2120
rect -900 1725 -750 1730
rect 2440 1725 2590 1730
rect -1195 815 -375 1455
rect 395 1215 1295 1505
rect 2065 815 2885 1455
rect -1195 400 -375 640
rect 2065 400 2885 640
<< nmos >>
rect -65 700 -50 850
rect -10 700 5 850
rect 45 700 60 850
rect 100 700 115 850
rect 155 700 170 850
rect 210 700 225 850
rect 265 700 280 850
rect 320 700 335 850
rect 375 700 390 850
rect 430 700 445 850
rect 485 700 500 850
rect 540 700 555 850
rect 755 625 770 875
rect 810 625 825 875
rect 865 625 880 875
rect 920 625 935 875
rect 1135 700 1150 850
rect 1190 700 1205 850
rect 1245 700 1260 850
rect 1300 700 1315 850
rect 1355 700 1370 850
rect 1410 700 1425 850
rect 1465 700 1480 850
rect 1520 700 1535 850
rect 1575 700 1590 850
rect 1630 700 1645 850
rect 1685 700 1700 850
rect 1740 700 1755 850
rect -65 305 -50 455
rect -10 305 5 455
rect 45 305 60 455
rect 100 305 115 455
rect 155 305 170 455
rect 210 305 225 455
rect 265 305 280 455
rect 320 305 335 455
rect 375 305 390 455
rect 430 305 445 455
rect 485 305 500 455
rect 540 305 555 455
rect 755 305 770 455
rect 810 305 825 455
rect 865 305 880 455
rect 920 305 935 455
rect 1135 305 1150 455
rect 1190 305 1205 455
rect 1245 305 1260 455
rect 1300 305 1315 455
rect 1355 305 1370 455
rect 1410 305 1425 455
rect 1465 305 1480 455
rect 1520 305 1535 455
rect 1575 305 1590 455
rect 1630 305 1645 455
rect 1685 305 1700 455
rect 1740 305 1755 455
rect -1095 -70 -1080 230
rect -1040 -70 -1025 230
rect -985 -70 -970 230
rect -930 -70 -915 230
rect -875 -70 -860 230
rect -820 -70 -805 230
rect -765 -70 -750 230
rect -710 -70 -695 230
rect -655 -70 -640 230
rect -600 -70 -585 230
rect -545 -70 -530 230
rect -490 -70 -475 230
rect 755 -290 770 -40
rect 810 -290 825 -40
rect 865 -290 880 -40
rect 920 -290 935 -40
rect 2165 -70 2180 230
rect 2220 -70 2235 230
rect 2275 -70 2290 230
rect 2330 -70 2345 230
rect 2385 -70 2400 230
rect 2440 -70 2455 230
rect 2495 -70 2510 230
rect 2550 -70 2565 230
rect 2605 -70 2620 230
rect 2660 -70 2675 230
rect 2715 -70 2730 230
rect 2770 -70 2785 230
rect -1065 -1055 -1005 -355
rect -965 -1055 -905 -355
rect -865 -1055 -805 -355
rect -765 -1055 -705 -355
rect -665 -1055 -605 -355
rect -565 -1055 -505 -355
rect 315 -785 330 -535
rect 370 -785 385 -535
rect 425 -785 440 -535
rect 480 -785 495 -535
rect 535 -785 550 -535
rect 590 -785 605 -535
rect 645 -785 660 -535
rect 700 -785 715 -535
rect 755 -785 770 -535
rect 810 -785 825 -535
rect 865 -785 880 -535
rect 920 -785 935 -535
rect 975 -785 990 -535
rect 1030 -785 1045 -535
rect 1085 -785 1100 -535
rect 1140 -785 1155 -535
rect 1195 -785 1210 -535
rect 1250 -785 1265 -535
rect 1305 -785 1320 -535
rect 1360 -785 1375 -535
rect 1415 -785 1430 -535
rect 535 -1100 550 -950
rect 590 -1100 605 -950
rect 645 -1100 660 -950
rect 700 -1100 715 -950
rect 755 -1100 770 -950
rect 810 -1100 825 -950
rect 1000 -1100 1300 -950
rect 2195 -1055 2255 -355
rect 2295 -1055 2355 -355
rect 2395 -1055 2455 -355
rect 2495 -1055 2555 -355
rect 2595 -1055 2655 -355
rect 2695 -1055 2755 -355
<< pmos >>
rect 70 2325 90 2675
rect 130 2325 150 2675
rect 190 2325 210 2675
rect 540 2325 560 2505
rect 600 2325 620 2505
rect 660 2325 680 2505
rect 1010 2325 1030 2675
rect 1070 2325 1090 2675
rect 1130 2325 1150 2675
rect 1480 2325 1500 2675
rect 1540 2325 1560 2675
rect 1600 2325 1620 2675
rect -1125 1750 -1105 2100
rect -1065 1750 -1045 2100
rect -1005 1750 -985 2100
rect -945 1750 -925 2100
rect -885 1750 -865 2100
rect -825 1750 -805 2100
rect -765 1750 -745 2100
rect -705 1750 -685 2100
rect -645 1750 -625 2100
rect -585 1750 -565 2100
rect -525 1750 -505 2100
rect -465 1750 -445 2100
rect 0 1750 20 2100
rect 60 1750 80 2100
rect 120 1750 140 2100
rect 180 1750 200 2100
rect 240 1750 260 2100
rect 300 1750 320 2100
rect 360 1750 380 2100
rect 420 1750 440 2100
rect 480 1750 500 2100
rect 540 1750 560 2100
rect 600 1750 620 2100
rect 660 1750 680 2100
rect 1010 1750 1030 2100
rect 1070 1750 1090 2100
rect 1130 1750 1150 2100
rect 1190 1750 1210 2100
rect 1250 1750 1270 2100
rect 1310 1750 1330 2100
rect 1370 1750 1390 2100
rect 1430 1750 1450 2100
rect 1490 1750 1510 2100
rect 1550 1750 1570 2100
rect 1610 1750 1630 2100
rect 1670 1750 1690 2100
rect 2135 1750 2155 2100
rect 2195 1750 2215 2100
rect 2255 1750 2275 2100
rect 2315 1750 2335 2100
rect 2375 1750 2395 2100
rect 2435 1750 2455 2100
rect 2495 1750 2515 2100
rect 2555 1750 2575 2100
rect 2615 1750 2635 2100
rect 2675 1750 2695 2100
rect 2735 1750 2755 2100
rect 2795 1750 2815 2100
rect -1095 835 -1080 1435
rect -1040 835 -1025 1435
rect -985 835 -970 1435
rect -930 835 -915 1435
rect -875 835 -860 1435
rect -820 835 -805 1435
rect -765 835 -750 1435
rect -710 835 -695 1435
rect -655 835 -640 1435
rect -600 835 -585 1435
rect -545 835 -530 1435
rect -490 835 -475 1435
rect 495 1235 510 1485
rect 550 1235 565 1485
rect 605 1235 620 1485
rect 660 1235 675 1485
rect 715 1235 730 1485
rect 770 1235 785 1485
rect 905 1235 920 1485
rect 960 1235 975 1485
rect 1015 1235 1030 1485
rect 1070 1235 1085 1485
rect 1125 1235 1140 1485
rect 1180 1235 1195 1485
rect 2165 835 2180 1435
rect 2220 835 2235 1435
rect 2275 835 2290 1435
rect 2330 835 2345 1435
rect 2385 835 2400 1435
rect 2440 835 2455 1435
rect 2495 835 2510 1435
rect 2550 835 2565 1435
rect 2605 835 2620 1435
rect 2660 835 2675 1435
rect 2715 835 2730 1435
rect 2770 835 2785 1435
rect -1095 420 -1080 620
rect -1040 420 -1025 620
rect -985 420 -970 620
rect -930 420 -915 620
rect -875 420 -860 620
rect -820 420 -805 620
rect -765 420 -750 620
rect -710 420 -695 620
rect -655 420 -640 620
rect -600 420 -585 620
rect -545 420 -530 620
rect -490 420 -475 620
rect 2165 420 2180 620
rect 2220 420 2235 620
rect 2275 420 2290 620
rect 2330 420 2345 620
rect 2385 420 2400 620
rect 2440 420 2455 620
rect 2495 420 2510 620
rect 2550 420 2565 620
rect 2605 420 2620 620
rect 2660 420 2675 620
rect 2715 420 2730 620
rect 2770 420 2785 620
<< ndiff >>
rect 715 860 755 875
rect -105 835 -65 850
rect -105 715 -95 835
rect -75 715 -65 835
rect -105 700 -65 715
rect -50 835 -10 850
rect -50 715 -40 835
rect -20 715 -10 835
rect -50 700 -10 715
rect 5 835 45 850
rect 5 715 15 835
rect 35 715 45 835
rect 5 700 45 715
rect 60 835 100 850
rect 60 715 70 835
rect 90 715 100 835
rect 60 700 100 715
rect 115 835 155 850
rect 115 715 125 835
rect 145 715 155 835
rect 115 700 155 715
rect 170 835 210 850
rect 170 715 180 835
rect 200 715 210 835
rect 170 700 210 715
rect 225 835 265 850
rect 225 715 235 835
rect 255 715 265 835
rect 225 700 265 715
rect 280 835 320 850
rect 280 715 290 835
rect 310 715 320 835
rect 280 700 320 715
rect 335 835 375 850
rect 335 715 345 835
rect 365 715 375 835
rect 335 700 375 715
rect 390 835 430 850
rect 390 715 400 835
rect 420 715 430 835
rect 390 700 430 715
rect 445 835 485 850
rect 445 715 455 835
rect 475 715 485 835
rect 445 700 485 715
rect 500 835 540 850
rect 500 715 510 835
rect 530 715 540 835
rect 500 700 540 715
rect 555 835 595 850
rect 555 715 565 835
rect 585 715 595 835
rect 555 700 595 715
rect 715 640 725 860
rect 745 640 755 860
rect 715 625 755 640
rect 770 860 810 875
rect 770 640 780 860
rect 800 640 810 860
rect 770 625 810 640
rect 825 860 865 875
rect 825 640 835 860
rect 855 640 865 860
rect 825 625 865 640
rect 880 860 920 875
rect 880 640 890 860
rect 910 640 920 860
rect 880 625 920 640
rect 935 860 975 875
rect 935 640 945 860
rect 965 640 975 860
rect 1095 835 1135 850
rect 1095 715 1105 835
rect 1125 715 1135 835
rect 1095 700 1135 715
rect 1150 835 1190 850
rect 1150 715 1160 835
rect 1180 715 1190 835
rect 1150 700 1190 715
rect 1205 835 1245 850
rect 1205 715 1215 835
rect 1235 715 1245 835
rect 1205 700 1245 715
rect 1260 835 1300 850
rect 1260 715 1270 835
rect 1290 715 1300 835
rect 1260 700 1300 715
rect 1315 835 1355 850
rect 1315 715 1325 835
rect 1345 715 1355 835
rect 1315 700 1355 715
rect 1370 835 1410 850
rect 1370 715 1380 835
rect 1400 715 1410 835
rect 1370 700 1410 715
rect 1425 835 1465 850
rect 1425 715 1435 835
rect 1455 715 1465 835
rect 1425 700 1465 715
rect 1480 835 1520 850
rect 1480 715 1490 835
rect 1510 715 1520 835
rect 1480 700 1520 715
rect 1535 835 1575 850
rect 1535 715 1545 835
rect 1565 715 1575 835
rect 1535 700 1575 715
rect 1590 835 1630 850
rect 1590 715 1600 835
rect 1620 715 1630 835
rect 1590 700 1630 715
rect 1645 835 1685 850
rect 1645 715 1655 835
rect 1675 715 1685 835
rect 1645 700 1685 715
rect 1700 835 1740 850
rect 1700 715 1710 835
rect 1730 715 1740 835
rect 1700 700 1740 715
rect 1755 835 1795 850
rect 1755 715 1765 835
rect 1785 715 1795 835
rect 1755 700 1795 715
rect 935 625 975 640
rect -105 440 -65 455
rect -105 320 -95 440
rect -75 320 -65 440
rect -105 305 -65 320
rect -50 440 -10 455
rect -50 320 -40 440
rect -20 320 -10 440
rect -50 305 -10 320
rect 5 440 45 455
rect 5 320 15 440
rect 35 320 45 440
rect 5 305 45 320
rect 60 440 100 455
rect 60 320 70 440
rect 90 320 100 440
rect 60 305 100 320
rect 115 440 155 455
rect 115 320 125 440
rect 145 320 155 440
rect 115 305 155 320
rect 170 440 210 455
rect 170 320 180 440
rect 200 320 210 440
rect 170 305 210 320
rect 225 440 265 455
rect 225 320 235 440
rect 255 320 265 440
rect 225 305 265 320
rect 280 440 320 455
rect 280 320 290 440
rect 310 320 320 440
rect 280 305 320 320
rect 335 440 375 455
rect 335 320 345 440
rect 365 320 375 440
rect 335 305 375 320
rect 390 440 430 455
rect 390 320 400 440
rect 420 320 430 440
rect 390 305 430 320
rect 445 440 485 455
rect 445 320 455 440
rect 475 320 485 440
rect 445 305 485 320
rect 500 440 540 455
rect 500 320 510 440
rect 530 320 540 440
rect 500 305 540 320
rect 555 440 595 455
rect 555 320 565 440
rect 585 320 595 440
rect 555 305 595 320
rect 715 440 755 455
rect 715 320 725 440
rect 745 320 755 440
rect 715 305 755 320
rect 770 440 810 455
rect 770 320 780 440
rect 800 320 810 440
rect 770 305 810 320
rect 825 440 865 455
rect 825 320 835 440
rect 855 320 865 440
rect 825 305 865 320
rect 880 440 920 455
rect 880 320 890 440
rect 910 320 920 440
rect 880 305 920 320
rect 935 440 975 455
rect 935 320 945 440
rect 965 320 975 440
rect 935 305 975 320
rect 1095 440 1135 455
rect 1095 320 1105 440
rect 1125 320 1135 440
rect 1095 305 1135 320
rect 1150 440 1190 455
rect 1150 320 1160 440
rect 1180 320 1190 440
rect 1150 305 1190 320
rect 1205 440 1245 455
rect 1205 320 1215 440
rect 1235 320 1245 440
rect 1205 305 1245 320
rect 1260 440 1300 455
rect 1260 320 1270 440
rect 1290 320 1300 440
rect 1260 305 1300 320
rect 1315 440 1355 455
rect 1315 320 1325 440
rect 1345 320 1355 440
rect 1315 305 1355 320
rect 1370 440 1410 455
rect 1370 320 1380 440
rect 1400 320 1410 440
rect 1370 305 1410 320
rect 1425 440 1465 455
rect 1425 320 1435 440
rect 1455 320 1465 440
rect 1425 305 1465 320
rect 1480 440 1520 455
rect 1480 320 1490 440
rect 1510 320 1520 440
rect 1480 305 1520 320
rect 1535 440 1575 455
rect 1535 320 1545 440
rect 1565 320 1575 440
rect 1535 305 1575 320
rect 1590 440 1630 455
rect 1590 320 1600 440
rect 1620 320 1630 440
rect 1590 305 1630 320
rect 1645 440 1685 455
rect 1645 320 1655 440
rect 1675 320 1685 440
rect 1645 305 1685 320
rect 1700 440 1740 455
rect 1700 320 1710 440
rect 1730 320 1740 440
rect 1700 305 1740 320
rect 1755 440 1795 455
rect 1755 320 1765 440
rect 1785 320 1795 440
rect 1755 305 1795 320
rect -1135 215 -1095 230
rect -1135 -55 -1125 215
rect -1105 -55 -1095 215
rect -1135 -70 -1095 -55
rect -1080 215 -1040 230
rect -1080 -55 -1070 215
rect -1050 -55 -1040 215
rect -1080 -70 -1040 -55
rect -1025 215 -985 230
rect -1025 -55 -1015 215
rect -995 -55 -985 215
rect -1025 -70 -985 -55
rect -970 215 -930 230
rect -970 -55 -960 215
rect -940 -55 -930 215
rect -970 -70 -930 -55
rect -915 215 -875 230
rect -915 -55 -905 215
rect -885 -55 -875 215
rect -915 -70 -875 -55
rect -860 215 -820 230
rect -860 -55 -850 215
rect -830 -55 -820 215
rect -860 -70 -820 -55
rect -805 215 -765 230
rect -805 -55 -795 215
rect -775 -55 -765 215
rect -805 -70 -765 -55
rect -750 215 -710 230
rect -750 -55 -740 215
rect -720 -55 -710 215
rect -750 -70 -710 -55
rect -695 215 -655 230
rect -695 -55 -685 215
rect -665 -55 -655 215
rect -695 -70 -655 -55
rect -640 215 -600 230
rect -640 -55 -630 215
rect -610 -55 -600 215
rect -640 -70 -600 -55
rect -585 215 -545 230
rect -585 -55 -575 215
rect -555 -55 -545 215
rect -585 -70 -545 -55
rect -530 215 -490 230
rect -530 -55 -520 215
rect -500 -55 -490 215
rect -530 -70 -490 -55
rect -475 215 -435 230
rect -475 -55 -465 215
rect -445 -55 -435 215
rect 2125 215 2165 230
rect -475 -70 -435 -55
rect 715 -55 755 -40
rect 715 -275 725 -55
rect 745 -275 755 -55
rect 715 -290 755 -275
rect 770 -55 810 -40
rect 770 -275 780 -55
rect 800 -275 810 -55
rect 770 -290 810 -275
rect 825 -55 865 -40
rect 825 -275 835 -55
rect 855 -275 865 -55
rect 825 -290 865 -275
rect 880 -55 920 -40
rect 880 -275 890 -55
rect 910 -275 920 -55
rect 880 -290 920 -275
rect 935 -55 975 -40
rect 935 -275 945 -55
rect 965 -275 975 -55
rect 2125 -55 2135 215
rect 2155 -55 2165 215
rect 2125 -70 2165 -55
rect 2180 215 2220 230
rect 2180 -55 2190 215
rect 2210 -55 2220 215
rect 2180 -70 2220 -55
rect 2235 215 2275 230
rect 2235 -55 2245 215
rect 2265 -55 2275 215
rect 2235 -70 2275 -55
rect 2290 215 2330 230
rect 2290 -55 2300 215
rect 2320 -55 2330 215
rect 2290 -70 2330 -55
rect 2345 215 2385 230
rect 2345 -55 2355 215
rect 2375 -55 2385 215
rect 2345 -70 2385 -55
rect 2400 215 2440 230
rect 2400 -55 2410 215
rect 2430 -55 2440 215
rect 2400 -70 2440 -55
rect 2455 215 2495 230
rect 2455 -55 2465 215
rect 2485 -55 2495 215
rect 2455 -70 2495 -55
rect 2510 215 2550 230
rect 2510 -55 2520 215
rect 2540 -55 2550 215
rect 2510 -70 2550 -55
rect 2565 215 2605 230
rect 2565 -55 2575 215
rect 2595 -55 2605 215
rect 2565 -70 2605 -55
rect 2620 215 2660 230
rect 2620 -55 2630 215
rect 2650 -55 2660 215
rect 2620 -70 2660 -55
rect 2675 215 2715 230
rect 2675 -55 2685 215
rect 2705 -55 2715 215
rect 2675 -70 2715 -55
rect 2730 215 2770 230
rect 2730 -55 2740 215
rect 2760 -55 2770 215
rect 2730 -70 2770 -55
rect 2785 215 2825 230
rect 2785 -55 2795 215
rect 2815 -55 2825 215
rect 2785 -70 2825 -55
rect 935 -290 975 -275
rect -1105 -370 -1065 -355
rect -1105 -1040 -1095 -370
rect -1075 -1040 -1065 -370
rect -1105 -1055 -1065 -1040
rect -1005 -370 -965 -355
rect -1005 -1040 -995 -370
rect -975 -1040 -965 -370
rect -1005 -1055 -965 -1040
rect -905 -370 -865 -355
rect -905 -1040 -895 -370
rect -875 -1040 -865 -370
rect -905 -1055 -865 -1040
rect -805 -370 -765 -355
rect -805 -1040 -795 -370
rect -775 -1040 -765 -370
rect -805 -1055 -765 -1040
rect -705 -370 -665 -355
rect -705 -1040 -695 -370
rect -675 -1040 -665 -370
rect -705 -1055 -665 -1040
rect -605 -370 -565 -355
rect -605 -1040 -595 -370
rect -575 -1040 -565 -370
rect -605 -1055 -565 -1040
rect -505 -370 -465 -355
rect -505 -1040 -495 -370
rect -475 -1040 -465 -370
rect 2155 -370 2195 -355
rect 275 -550 315 -535
rect 275 -770 285 -550
rect 305 -770 315 -550
rect 275 -785 315 -770
rect 330 -550 370 -535
rect 330 -770 340 -550
rect 360 -770 370 -550
rect 330 -785 370 -770
rect 385 -550 425 -535
rect 385 -770 395 -550
rect 415 -770 425 -550
rect 385 -785 425 -770
rect 440 -550 480 -535
rect 440 -770 450 -550
rect 470 -770 480 -550
rect 440 -785 480 -770
rect 495 -550 535 -535
rect 495 -770 505 -550
rect 525 -770 535 -550
rect 495 -785 535 -770
rect 550 -550 590 -535
rect 550 -770 560 -550
rect 580 -770 590 -550
rect 550 -785 590 -770
rect 605 -550 645 -535
rect 605 -770 615 -550
rect 635 -770 645 -550
rect 605 -785 645 -770
rect 660 -550 700 -535
rect 660 -770 670 -550
rect 690 -770 700 -550
rect 660 -785 700 -770
rect 715 -550 755 -535
rect 715 -770 725 -550
rect 745 -770 755 -550
rect 715 -785 755 -770
rect 770 -550 810 -535
rect 770 -770 780 -550
rect 800 -770 810 -550
rect 770 -785 810 -770
rect 825 -550 865 -535
rect 825 -770 835 -550
rect 855 -770 865 -550
rect 825 -785 865 -770
rect 880 -550 920 -535
rect 880 -770 890 -550
rect 910 -770 920 -550
rect 880 -785 920 -770
rect 935 -550 975 -535
rect 935 -770 945 -550
rect 965 -770 975 -550
rect 935 -785 975 -770
rect 990 -550 1030 -535
rect 990 -770 1000 -550
rect 1020 -770 1030 -550
rect 990 -785 1030 -770
rect 1045 -550 1085 -535
rect 1045 -770 1055 -550
rect 1075 -770 1085 -550
rect 1045 -785 1085 -770
rect 1100 -550 1140 -535
rect 1100 -770 1110 -550
rect 1130 -770 1140 -550
rect 1100 -785 1140 -770
rect 1155 -550 1195 -535
rect 1155 -770 1165 -550
rect 1185 -770 1195 -550
rect 1155 -785 1195 -770
rect 1210 -550 1250 -535
rect 1210 -770 1220 -550
rect 1240 -770 1250 -550
rect 1210 -785 1250 -770
rect 1265 -550 1305 -535
rect 1265 -770 1275 -550
rect 1295 -770 1305 -550
rect 1265 -785 1305 -770
rect 1320 -550 1360 -535
rect 1320 -770 1330 -550
rect 1350 -770 1360 -550
rect 1320 -785 1360 -770
rect 1375 -550 1415 -535
rect 1375 -770 1385 -550
rect 1405 -770 1415 -550
rect 1375 -785 1415 -770
rect 1430 -550 1470 -535
rect 1430 -770 1440 -550
rect 1460 -770 1470 -550
rect 1430 -785 1470 -770
rect -505 -1055 -465 -1040
rect 495 -965 535 -950
rect 495 -1085 505 -965
rect 525 -1085 535 -965
rect 495 -1100 535 -1085
rect 550 -965 590 -950
rect 550 -1085 560 -965
rect 580 -1085 590 -965
rect 550 -1100 590 -1085
rect 605 -965 645 -950
rect 605 -1085 615 -965
rect 635 -1085 645 -965
rect 605 -1100 645 -1085
rect 660 -965 700 -950
rect 660 -1085 670 -965
rect 690 -1085 700 -965
rect 660 -1100 700 -1085
rect 715 -965 755 -950
rect 715 -1085 725 -965
rect 745 -1085 755 -965
rect 715 -1100 755 -1085
rect 770 -965 810 -950
rect 770 -1085 780 -965
rect 800 -1085 810 -965
rect 770 -1100 810 -1085
rect 825 -965 865 -950
rect 825 -1085 835 -965
rect 855 -1085 865 -965
rect 825 -1100 865 -1085
rect 960 -965 1000 -950
rect 960 -1085 970 -965
rect 990 -1085 1000 -965
rect 960 -1100 1000 -1085
rect 1300 -965 1340 -950
rect 1300 -1085 1310 -965
rect 1330 -1085 1340 -965
rect 2155 -1040 2165 -370
rect 2185 -1040 2195 -370
rect 2155 -1055 2195 -1040
rect 2255 -370 2295 -355
rect 2255 -1040 2265 -370
rect 2285 -1040 2295 -370
rect 2255 -1055 2295 -1040
rect 2355 -370 2395 -355
rect 2355 -1040 2365 -370
rect 2385 -1040 2395 -370
rect 2355 -1055 2395 -1040
rect 2455 -370 2495 -355
rect 2455 -1040 2465 -370
rect 2485 -1040 2495 -370
rect 2455 -1055 2495 -1040
rect 2555 -370 2595 -355
rect 2555 -1040 2565 -370
rect 2585 -1040 2595 -370
rect 2555 -1055 2595 -1040
rect 2655 -370 2695 -355
rect 2655 -1040 2665 -370
rect 2685 -1040 2695 -370
rect 2655 -1055 2695 -1040
rect 2755 -370 2795 -355
rect 2755 -1040 2765 -370
rect 2785 -1040 2795 -370
rect 2755 -1055 2795 -1040
rect 1300 -1100 1340 -1085
<< pdiff >>
rect 30 2660 70 2675
rect 30 2340 40 2660
rect 60 2340 70 2660
rect 30 2325 70 2340
rect 90 2660 130 2675
rect 90 2340 100 2660
rect 120 2340 130 2660
rect 90 2325 130 2340
rect 150 2660 190 2675
rect 150 2340 160 2660
rect 180 2340 190 2660
rect 150 2325 190 2340
rect 210 2660 250 2675
rect 210 2340 220 2660
rect 240 2340 250 2660
rect 970 2660 1010 2675
rect 210 2325 250 2340
rect 500 2490 540 2505
rect 500 2340 510 2490
rect 530 2340 540 2490
rect 500 2325 540 2340
rect 560 2490 600 2505
rect 560 2340 570 2490
rect 590 2340 600 2490
rect 560 2325 600 2340
rect 620 2490 660 2505
rect 620 2340 630 2490
rect 650 2340 660 2490
rect 620 2325 660 2340
rect 680 2490 720 2505
rect 680 2340 690 2490
rect 710 2340 720 2490
rect 680 2325 720 2340
rect 970 2340 980 2660
rect 1000 2340 1010 2660
rect 970 2325 1010 2340
rect 1030 2660 1070 2675
rect 1030 2340 1040 2660
rect 1060 2340 1070 2660
rect 1030 2325 1070 2340
rect 1090 2660 1130 2675
rect 1090 2340 1100 2660
rect 1120 2340 1130 2660
rect 1090 2325 1130 2340
rect 1150 2660 1190 2675
rect 1150 2340 1160 2660
rect 1180 2340 1190 2660
rect 1150 2325 1190 2340
rect 1440 2660 1480 2675
rect 1440 2340 1450 2660
rect 1470 2340 1480 2660
rect 1440 2325 1480 2340
rect 1500 2660 1540 2675
rect 1500 2340 1510 2660
rect 1530 2340 1540 2660
rect 1500 2325 1540 2340
rect 1560 2660 1600 2675
rect 1560 2340 1570 2660
rect 1590 2340 1600 2660
rect 1560 2325 1600 2340
rect 1620 2660 1660 2675
rect 1620 2340 1630 2660
rect 1650 2340 1660 2660
rect 1620 2325 1660 2340
rect -1165 2085 -1125 2100
rect -1165 1765 -1155 2085
rect -1135 1765 -1125 2085
rect -1165 1750 -1125 1765
rect -1105 2085 -1065 2100
rect -1105 1765 -1095 2085
rect -1075 1765 -1065 2085
rect -1105 1750 -1065 1765
rect -1045 2085 -1005 2100
rect -1045 1765 -1035 2085
rect -1015 1765 -1005 2085
rect -1045 1750 -1005 1765
rect -985 2085 -945 2100
rect -985 1765 -975 2085
rect -955 1765 -945 2085
rect -985 1750 -945 1765
rect -925 2085 -885 2100
rect -925 1765 -915 2085
rect -895 1765 -885 2085
rect -925 1750 -885 1765
rect -865 2085 -825 2100
rect -865 1765 -855 2085
rect -835 1765 -825 2085
rect -865 1750 -825 1765
rect -805 2085 -765 2100
rect -805 1765 -795 2085
rect -775 1765 -765 2085
rect -805 1750 -765 1765
rect -745 2085 -705 2100
rect -745 1765 -735 2085
rect -715 1765 -705 2085
rect -745 1750 -705 1765
rect -685 2085 -645 2100
rect -685 1765 -675 2085
rect -655 1765 -645 2085
rect -685 1750 -645 1765
rect -625 2085 -585 2100
rect -625 1765 -615 2085
rect -595 1765 -585 2085
rect -625 1750 -585 1765
rect -565 2085 -525 2100
rect -565 1765 -555 2085
rect -535 1765 -525 2085
rect -565 1750 -525 1765
rect -505 2085 -465 2100
rect -505 1765 -495 2085
rect -475 1765 -465 2085
rect -505 1750 -465 1765
rect -445 2085 -405 2100
rect -445 1765 -435 2085
rect -415 1765 -405 2085
rect -445 1750 -405 1765
rect -40 2085 0 2100
rect -40 1765 -30 2085
rect -10 1765 0 2085
rect -40 1750 0 1765
rect 20 2085 60 2100
rect 20 1765 30 2085
rect 50 1765 60 2085
rect 20 1750 60 1765
rect 80 2085 120 2100
rect 80 1765 90 2085
rect 110 1765 120 2085
rect 80 1750 120 1765
rect 140 2085 180 2100
rect 140 1765 150 2085
rect 170 1765 180 2085
rect 140 1750 180 1765
rect 200 2085 240 2100
rect 200 1765 210 2085
rect 230 1765 240 2085
rect 200 1750 240 1765
rect 260 2085 300 2100
rect 260 1765 270 2085
rect 290 1765 300 2085
rect 260 1750 300 1765
rect 320 2085 360 2100
rect 320 1765 330 2085
rect 350 1765 360 2085
rect 320 1750 360 1765
rect 380 2085 420 2100
rect 380 1765 390 2085
rect 410 1765 420 2085
rect 380 1750 420 1765
rect 440 2085 480 2100
rect 440 1765 450 2085
rect 470 1765 480 2085
rect 440 1750 480 1765
rect 500 2085 540 2100
rect 500 1765 510 2085
rect 530 1765 540 2085
rect 500 1750 540 1765
rect 560 2085 600 2100
rect 560 1765 570 2085
rect 590 1765 600 2085
rect 560 1750 600 1765
rect 620 2085 660 2100
rect 620 1765 630 2085
rect 650 1765 660 2085
rect 620 1750 660 1765
rect 680 2085 720 2100
rect 680 1765 690 2085
rect 710 1765 720 2085
rect 680 1750 720 1765
rect 970 2085 1010 2100
rect 970 1765 980 2085
rect 1000 1765 1010 2085
rect 970 1750 1010 1765
rect 1030 2085 1070 2100
rect 1030 1765 1040 2085
rect 1060 1765 1070 2085
rect 1030 1750 1070 1765
rect 1090 2085 1130 2100
rect 1090 1765 1100 2085
rect 1120 1765 1130 2085
rect 1090 1750 1130 1765
rect 1150 2085 1190 2100
rect 1150 1765 1160 2085
rect 1180 1765 1190 2085
rect 1150 1750 1190 1765
rect 1210 2085 1250 2100
rect 1210 1765 1220 2085
rect 1240 1765 1250 2085
rect 1210 1750 1250 1765
rect 1270 2085 1310 2100
rect 1270 1765 1280 2085
rect 1300 1765 1310 2085
rect 1270 1750 1310 1765
rect 1330 2085 1370 2100
rect 1330 1765 1340 2085
rect 1360 1765 1370 2085
rect 1330 1750 1370 1765
rect 1390 2085 1430 2100
rect 1390 1765 1400 2085
rect 1420 1765 1430 2085
rect 1390 1750 1430 1765
rect 1450 2085 1490 2100
rect 1450 1765 1460 2085
rect 1480 1765 1490 2085
rect 1450 1750 1490 1765
rect 1510 2085 1550 2100
rect 1510 1765 1520 2085
rect 1540 1765 1550 2085
rect 1510 1750 1550 1765
rect 1570 2085 1610 2100
rect 1570 1765 1580 2085
rect 1600 1765 1610 2085
rect 1570 1750 1610 1765
rect 1630 2085 1670 2100
rect 1630 1765 1640 2085
rect 1660 1765 1670 2085
rect 1630 1750 1670 1765
rect 1690 2085 1730 2100
rect 1690 1765 1700 2085
rect 1720 1765 1730 2085
rect 1690 1750 1730 1765
rect 2095 2085 2135 2100
rect 2095 1765 2105 2085
rect 2125 1765 2135 2085
rect 2095 1750 2135 1765
rect 2155 2085 2195 2100
rect 2155 1765 2165 2085
rect 2185 1765 2195 2085
rect 2155 1750 2195 1765
rect 2215 2085 2255 2100
rect 2215 1765 2225 2085
rect 2245 1765 2255 2085
rect 2215 1750 2255 1765
rect 2275 2085 2315 2100
rect 2275 1765 2285 2085
rect 2305 1765 2315 2085
rect 2275 1750 2315 1765
rect 2335 2085 2375 2100
rect 2335 1765 2345 2085
rect 2365 1765 2375 2085
rect 2335 1750 2375 1765
rect 2395 2085 2435 2100
rect 2395 1765 2405 2085
rect 2425 1765 2435 2085
rect 2395 1750 2435 1765
rect 2455 2085 2495 2100
rect 2455 1765 2465 2085
rect 2485 1765 2495 2085
rect 2455 1750 2495 1765
rect 2515 2085 2555 2100
rect 2515 1765 2525 2085
rect 2545 1765 2555 2085
rect 2515 1750 2555 1765
rect 2575 2085 2615 2100
rect 2575 1765 2585 2085
rect 2605 1765 2615 2085
rect 2575 1750 2615 1765
rect 2635 2085 2675 2100
rect 2635 1765 2645 2085
rect 2665 1765 2675 2085
rect 2635 1750 2675 1765
rect 2695 2085 2735 2100
rect 2695 1765 2705 2085
rect 2725 1765 2735 2085
rect 2695 1750 2735 1765
rect 2755 2085 2795 2100
rect 2755 1765 2765 2085
rect 2785 1765 2795 2085
rect 2755 1750 2795 1765
rect 2815 2085 2855 2100
rect 2815 1765 2825 2085
rect 2845 1765 2855 2085
rect 2815 1750 2855 1765
rect 455 1470 495 1485
rect -1135 1420 -1095 1435
rect -1135 850 -1125 1420
rect -1105 850 -1095 1420
rect -1135 835 -1095 850
rect -1080 1420 -1040 1435
rect -1080 850 -1070 1420
rect -1050 850 -1040 1420
rect -1080 835 -1040 850
rect -1025 1420 -985 1435
rect -1025 850 -1015 1420
rect -995 850 -985 1420
rect -1025 835 -985 850
rect -970 1420 -930 1435
rect -970 850 -960 1420
rect -940 850 -930 1420
rect -970 835 -930 850
rect -915 1420 -875 1435
rect -915 850 -905 1420
rect -885 850 -875 1420
rect -915 835 -875 850
rect -860 1420 -820 1435
rect -860 850 -850 1420
rect -830 850 -820 1420
rect -860 835 -820 850
rect -805 1420 -765 1435
rect -805 850 -795 1420
rect -775 850 -765 1420
rect -805 835 -765 850
rect -750 1420 -710 1435
rect -750 850 -740 1420
rect -720 850 -710 1420
rect -750 835 -710 850
rect -695 1420 -655 1435
rect -695 850 -685 1420
rect -665 850 -655 1420
rect -695 835 -655 850
rect -640 1420 -600 1435
rect -640 850 -630 1420
rect -610 850 -600 1420
rect -640 835 -600 850
rect -585 1420 -545 1435
rect -585 850 -575 1420
rect -555 850 -545 1420
rect -585 835 -545 850
rect -530 1420 -490 1435
rect -530 850 -520 1420
rect -500 850 -490 1420
rect -530 835 -490 850
rect -475 1420 -435 1435
rect -475 850 -465 1420
rect -445 850 -435 1420
rect 455 1250 465 1470
rect 485 1250 495 1470
rect 455 1235 495 1250
rect 510 1470 550 1485
rect 510 1250 520 1470
rect 540 1250 550 1470
rect 510 1235 550 1250
rect 565 1470 605 1485
rect 565 1250 575 1470
rect 595 1250 605 1470
rect 565 1235 605 1250
rect 620 1470 660 1485
rect 620 1250 630 1470
rect 650 1250 660 1470
rect 620 1235 660 1250
rect 675 1470 715 1485
rect 675 1250 685 1470
rect 705 1250 715 1470
rect 675 1235 715 1250
rect 730 1470 770 1485
rect 730 1250 740 1470
rect 760 1250 770 1470
rect 730 1235 770 1250
rect 785 1470 825 1485
rect 865 1470 905 1485
rect 785 1250 795 1470
rect 815 1250 825 1470
rect 865 1250 875 1470
rect 895 1250 905 1470
rect 785 1235 825 1250
rect 865 1235 905 1250
rect 920 1470 960 1485
rect 920 1250 930 1470
rect 950 1250 960 1470
rect 920 1235 960 1250
rect 975 1470 1015 1485
rect 975 1250 985 1470
rect 1005 1250 1015 1470
rect 975 1235 1015 1250
rect 1030 1470 1070 1485
rect 1030 1250 1040 1470
rect 1060 1250 1070 1470
rect 1030 1235 1070 1250
rect 1085 1470 1125 1485
rect 1085 1250 1095 1470
rect 1115 1250 1125 1470
rect 1085 1235 1125 1250
rect 1140 1470 1180 1485
rect 1140 1250 1150 1470
rect 1170 1250 1180 1470
rect 1140 1235 1180 1250
rect 1195 1470 1235 1485
rect 1195 1250 1205 1470
rect 1225 1250 1235 1470
rect 1195 1235 1235 1250
rect 2125 1420 2165 1435
rect -475 835 -435 850
rect 2125 850 2135 1420
rect 2155 850 2165 1420
rect 2125 835 2165 850
rect 2180 1420 2220 1435
rect 2180 850 2190 1420
rect 2210 850 2220 1420
rect 2180 835 2220 850
rect 2235 1420 2275 1435
rect 2235 850 2245 1420
rect 2265 850 2275 1420
rect 2235 835 2275 850
rect 2290 1420 2330 1435
rect 2290 850 2300 1420
rect 2320 850 2330 1420
rect 2290 835 2330 850
rect 2345 1420 2385 1435
rect 2345 850 2355 1420
rect 2375 850 2385 1420
rect 2345 835 2385 850
rect 2400 1420 2440 1435
rect 2400 850 2410 1420
rect 2430 850 2440 1420
rect 2400 835 2440 850
rect 2455 1420 2495 1435
rect 2455 850 2465 1420
rect 2485 850 2495 1420
rect 2455 835 2495 850
rect 2510 1420 2550 1435
rect 2510 850 2520 1420
rect 2540 850 2550 1420
rect 2510 835 2550 850
rect 2565 1420 2605 1435
rect 2565 850 2575 1420
rect 2595 850 2605 1420
rect 2565 835 2605 850
rect 2620 1420 2660 1435
rect 2620 850 2630 1420
rect 2650 850 2660 1420
rect 2620 835 2660 850
rect 2675 1420 2715 1435
rect 2675 850 2685 1420
rect 2705 850 2715 1420
rect 2675 835 2715 850
rect 2730 1420 2770 1435
rect 2730 850 2740 1420
rect 2760 850 2770 1420
rect 2730 835 2770 850
rect 2785 1420 2825 1435
rect 2785 850 2795 1420
rect 2815 850 2825 1420
rect 2785 835 2825 850
rect -1135 605 -1095 620
rect -1135 435 -1125 605
rect -1105 435 -1095 605
rect -1135 420 -1095 435
rect -1080 605 -1040 620
rect -1080 435 -1070 605
rect -1050 435 -1040 605
rect -1080 420 -1040 435
rect -1025 605 -985 620
rect -1025 435 -1015 605
rect -995 435 -985 605
rect -1025 420 -985 435
rect -970 605 -930 620
rect -970 435 -960 605
rect -940 435 -930 605
rect -970 420 -930 435
rect -915 605 -875 620
rect -915 435 -905 605
rect -885 435 -875 605
rect -915 420 -875 435
rect -860 605 -820 620
rect -860 435 -850 605
rect -830 435 -820 605
rect -860 420 -820 435
rect -805 605 -765 620
rect -805 435 -795 605
rect -775 435 -765 605
rect -805 420 -765 435
rect -750 605 -710 620
rect -750 435 -740 605
rect -720 435 -710 605
rect -750 420 -710 435
rect -695 605 -655 620
rect -695 435 -685 605
rect -665 435 -655 605
rect -695 420 -655 435
rect -640 605 -600 620
rect -640 435 -630 605
rect -610 435 -600 605
rect -640 420 -600 435
rect -585 605 -545 620
rect -585 435 -575 605
rect -555 435 -545 605
rect -585 420 -545 435
rect -530 605 -490 620
rect -530 435 -520 605
rect -500 435 -490 605
rect -530 420 -490 435
rect -475 605 -435 620
rect -475 435 -465 605
rect -445 435 -435 605
rect 2125 605 2165 620
rect -475 420 -435 435
rect 2125 435 2135 605
rect 2155 435 2165 605
rect 2125 420 2165 435
rect 2180 605 2220 620
rect 2180 435 2190 605
rect 2210 435 2220 605
rect 2180 420 2220 435
rect 2235 605 2275 620
rect 2235 435 2245 605
rect 2265 435 2275 605
rect 2235 420 2275 435
rect 2290 605 2330 620
rect 2290 435 2300 605
rect 2320 435 2330 605
rect 2290 420 2330 435
rect 2345 605 2385 620
rect 2345 435 2355 605
rect 2375 435 2385 605
rect 2345 420 2385 435
rect 2400 605 2440 620
rect 2400 435 2410 605
rect 2430 435 2440 605
rect 2400 420 2440 435
rect 2455 605 2495 620
rect 2455 435 2465 605
rect 2485 435 2495 605
rect 2455 420 2495 435
rect 2510 605 2550 620
rect 2510 435 2520 605
rect 2540 435 2550 605
rect 2510 420 2550 435
rect 2565 605 2605 620
rect 2565 435 2575 605
rect 2595 435 2605 605
rect 2565 420 2605 435
rect 2620 605 2660 620
rect 2620 435 2630 605
rect 2650 435 2660 605
rect 2620 420 2660 435
rect 2675 605 2715 620
rect 2675 435 2685 605
rect 2705 435 2715 605
rect 2675 420 2715 435
rect 2730 605 2770 620
rect 2730 435 2740 605
rect 2760 435 2770 605
rect 2730 420 2770 435
rect 2785 605 2825 620
rect 2785 435 2795 605
rect 2815 435 2825 605
rect 2785 420 2825 435
<< ndiffc >>
rect -95 715 -75 835
rect -40 715 -20 835
rect 15 715 35 835
rect 70 715 90 835
rect 125 715 145 835
rect 180 715 200 835
rect 235 715 255 835
rect 290 715 310 835
rect 345 715 365 835
rect 400 715 420 835
rect 455 715 475 835
rect 510 715 530 835
rect 565 715 585 835
rect 725 640 745 860
rect 780 640 800 860
rect 835 640 855 860
rect 890 640 910 860
rect 945 640 965 860
rect 1105 715 1125 835
rect 1160 715 1180 835
rect 1215 715 1235 835
rect 1270 715 1290 835
rect 1325 715 1345 835
rect 1380 715 1400 835
rect 1435 715 1455 835
rect 1490 715 1510 835
rect 1545 715 1565 835
rect 1600 715 1620 835
rect 1655 715 1675 835
rect 1710 715 1730 835
rect 1765 715 1785 835
rect -95 320 -75 440
rect -40 320 -20 440
rect 15 320 35 440
rect 70 320 90 440
rect 125 320 145 440
rect 180 320 200 440
rect 235 320 255 440
rect 290 320 310 440
rect 345 320 365 440
rect 400 320 420 440
rect 455 320 475 440
rect 510 320 530 440
rect 565 320 585 440
rect 725 320 745 440
rect 780 320 800 440
rect 835 320 855 440
rect 890 320 910 440
rect 945 320 965 440
rect 1105 320 1125 440
rect 1160 320 1180 440
rect 1215 320 1235 440
rect 1270 320 1290 440
rect 1325 320 1345 440
rect 1380 320 1400 440
rect 1435 320 1455 440
rect 1490 320 1510 440
rect 1545 320 1565 440
rect 1600 320 1620 440
rect 1655 320 1675 440
rect 1710 320 1730 440
rect 1765 320 1785 440
rect -1125 -55 -1105 215
rect -1070 -55 -1050 215
rect -1015 -55 -995 215
rect -960 -55 -940 215
rect -905 -55 -885 215
rect -850 -55 -830 215
rect -795 -55 -775 215
rect -740 -55 -720 215
rect -685 -55 -665 215
rect -630 -55 -610 215
rect -575 -55 -555 215
rect -520 -55 -500 215
rect -465 -55 -445 215
rect 725 -275 745 -55
rect 780 -275 800 -55
rect 835 -275 855 -55
rect 890 -275 910 -55
rect 945 -275 965 -55
rect 2135 -55 2155 215
rect 2190 -55 2210 215
rect 2245 -55 2265 215
rect 2300 -55 2320 215
rect 2355 -55 2375 215
rect 2410 -55 2430 215
rect 2465 -55 2485 215
rect 2520 -55 2540 215
rect 2575 -55 2595 215
rect 2630 -55 2650 215
rect 2685 -55 2705 215
rect 2740 -55 2760 215
rect 2795 -55 2815 215
rect -1095 -1040 -1075 -370
rect -995 -1040 -975 -370
rect -895 -1040 -875 -370
rect -795 -1040 -775 -370
rect -695 -1040 -675 -370
rect -595 -1040 -575 -370
rect -495 -1040 -475 -370
rect 285 -770 305 -550
rect 340 -770 360 -550
rect 395 -770 415 -550
rect 450 -770 470 -550
rect 505 -770 525 -550
rect 560 -770 580 -550
rect 615 -770 635 -550
rect 670 -770 690 -550
rect 725 -770 745 -550
rect 780 -770 800 -550
rect 835 -770 855 -550
rect 890 -770 910 -550
rect 945 -770 965 -550
rect 1000 -770 1020 -550
rect 1055 -770 1075 -550
rect 1110 -770 1130 -550
rect 1165 -770 1185 -550
rect 1220 -770 1240 -550
rect 1275 -770 1295 -550
rect 1330 -770 1350 -550
rect 1385 -770 1405 -550
rect 1440 -770 1460 -550
rect 505 -1085 525 -965
rect 560 -1085 580 -965
rect 615 -1085 635 -965
rect 670 -1085 690 -965
rect 725 -1085 745 -965
rect 780 -1085 800 -965
rect 835 -1085 855 -965
rect 970 -1085 990 -965
rect 1310 -1085 1330 -965
rect 2165 -1040 2185 -370
rect 2265 -1040 2285 -370
rect 2365 -1040 2385 -370
rect 2465 -1040 2485 -370
rect 2565 -1040 2585 -370
rect 2665 -1040 2685 -370
rect 2765 -1040 2785 -370
<< pdiffc >>
rect 40 2340 60 2660
rect 100 2340 120 2660
rect 160 2340 180 2660
rect 220 2340 240 2660
rect 510 2340 530 2490
rect 570 2340 590 2490
rect 630 2340 650 2490
rect 690 2340 710 2490
rect 980 2340 1000 2660
rect 1040 2340 1060 2660
rect 1100 2340 1120 2660
rect 1160 2340 1180 2660
rect 1450 2340 1470 2660
rect 1510 2340 1530 2660
rect 1570 2340 1590 2660
rect 1630 2340 1650 2660
rect -1155 1765 -1135 2085
rect -1095 1765 -1075 2085
rect -1035 1765 -1015 2085
rect -975 1765 -955 2085
rect -915 1765 -895 2085
rect -855 1765 -835 2085
rect -795 1765 -775 2085
rect -735 1765 -715 2085
rect -675 1765 -655 2085
rect -615 1765 -595 2085
rect -555 1765 -535 2085
rect -495 1765 -475 2085
rect -435 1765 -415 2085
rect -30 1765 -10 2085
rect 30 1765 50 2085
rect 90 1765 110 2085
rect 150 1765 170 2085
rect 210 1765 230 2085
rect 270 1765 290 2085
rect 330 1765 350 2085
rect 390 1765 410 2085
rect 450 1765 470 2085
rect 510 1765 530 2085
rect 570 1765 590 2085
rect 630 1765 650 2085
rect 690 1765 710 2085
rect 980 1765 1000 2085
rect 1040 1765 1060 2085
rect 1100 1765 1120 2085
rect 1160 1765 1180 2085
rect 1220 1765 1240 2085
rect 1280 1765 1300 2085
rect 1340 1765 1360 2085
rect 1400 1765 1420 2085
rect 1460 1765 1480 2085
rect 1520 1765 1540 2085
rect 1580 1765 1600 2085
rect 1640 1765 1660 2085
rect 1700 1765 1720 2085
rect 2105 1765 2125 2085
rect 2165 1765 2185 2085
rect 2225 1765 2245 2085
rect 2285 1765 2305 2085
rect 2345 1765 2365 2085
rect 2405 1765 2425 2085
rect 2465 1765 2485 2085
rect 2525 1765 2545 2085
rect 2585 1765 2605 2085
rect 2645 1765 2665 2085
rect 2705 1765 2725 2085
rect 2765 1765 2785 2085
rect 2825 1765 2845 2085
rect -1125 850 -1105 1420
rect -1070 850 -1050 1420
rect -1015 850 -995 1420
rect -960 850 -940 1420
rect -905 850 -885 1420
rect -850 850 -830 1420
rect -795 850 -775 1420
rect -740 850 -720 1420
rect -685 850 -665 1420
rect -630 850 -610 1420
rect -575 850 -555 1420
rect -520 850 -500 1420
rect -465 850 -445 1420
rect 465 1250 485 1470
rect 520 1250 540 1470
rect 575 1250 595 1470
rect 630 1250 650 1470
rect 685 1250 705 1470
rect 740 1250 760 1470
rect 795 1250 815 1470
rect 875 1250 895 1470
rect 930 1250 950 1470
rect 985 1250 1005 1470
rect 1040 1250 1060 1470
rect 1095 1250 1115 1470
rect 1150 1250 1170 1470
rect 1205 1250 1225 1470
rect 2135 850 2155 1420
rect 2190 850 2210 1420
rect 2245 850 2265 1420
rect 2300 850 2320 1420
rect 2355 850 2375 1420
rect 2410 850 2430 1420
rect 2465 850 2485 1420
rect 2520 850 2540 1420
rect 2575 850 2595 1420
rect 2630 850 2650 1420
rect 2685 850 2705 1420
rect 2740 850 2760 1420
rect 2795 850 2815 1420
rect -1125 435 -1105 605
rect -1070 435 -1050 605
rect -1015 435 -995 605
rect -960 435 -940 605
rect -905 435 -885 605
rect -850 435 -830 605
rect -795 435 -775 605
rect -740 435 -720 605
rect -685 435 -665 605
rect -630 435 -610 605
rect -575 435 -555 605
rect -520 435 -500 605
rect -465 435 -445 605
rect 2135 435 2155 605
rect 2190 435 2210 605
rect 2245 435 2265 605
rect 2300 435 2320 605
rect 2355 435 2375 605
rect 2410 435 2430 605
rect 2465 435 2485 605
rect 2520 435 2540 605
rect 2575 435 2595 605
rect 2630 435 2650 605
rect 2685 435 2705 605
rect 2740 435 2760 605
rect 2795 435 2815 605
<< psubdiff >>
rect 675 860 715 875
rect -145 835 -105 850
rect -145 715 -135 835
rect -115 715 -105 835
rect -145 700 -105 715
rect 595 835 635 850
rect 595 715 605 835
rect 625 715 635 835
rect 595 700 635 715
rect 675 640 685 860
rect 705 640 715 860
rect 675 625 715 640
rect 975 860 1015 875
rect 975 640 985 860
rect 1005 640 1015 860
rect 1055 835 1095 850
rect 1055 715 1065 835
rect 1085 715 1095 835
rect 1055 700 1095 715
rect 1795 835 1835 850
rect 1795 715 1805 835
rect 1825 715 1835 835
rect 1795 700 1835 715
rect 975 625 1015 640
rect -145 440 -105 455
rect -145 320 -135 440
rect -115 320 -105 440
rect -145 305 -105 320
rect 595 440 635 455
rect 595 320 605 440
rect 625 320 635 440
rect 595 305 635 320
rect 675 440 715 455
rect 675 320 685 440
rect 705 320 715 440
rect 675 305 715 320
rect 975 440 1015 455
rect 975 320 985 440
rect 1005 320 1015 440
rect 975 305 1015 320
rect 1055 440 1095 455
rect 1055 320 1065 440
rect 1085 320 1095 440
rect 1055 305 1095 320
rect 1795 440 1835 455
rect 1795 320 1805 440
rect 1825 320 1835 440
rect 1795 305 1835 320
rect -1175 215 -1135 230
rect -1175 -55 -1165 215
rect -1145 -55 -1135 215
rect -1175 -70 -1135 -55
rect -435 215 -395 230
rect -435 -55 -425 215
rect -405 -55 -395 215
rect 2085 215 2125 230
rect -435 -70 -395 -55
rect 675 -55 715 -40
rect 675 -275 685 -55
rect 705 -275 715 -55
rect 675 -290 715 -275
rect 975 -55 1015 -40
rect 975 -275 985 -55
rect 1005 -275 1015 -55
rect 2085 -55 2095 215
rect 2115 -55 2125 215
rect 2085 -70 2125 -55
rect 2825 215 2865 230
rect 2825 -55 2835 215
rect 2855 -55 2865 215
rect 2825 -70 2865 -55
rect 975 -290 1015 -275
rect -1145 -370 -1105 -355
rect -1145 -1040 -1135 -370
rect -1115 -1040 -1105 -370
rect -1145 -1055 -1105 -1040
rect -465 -370 -425 -355
rect -465 -1040 -455 -370
rect -435 -1040 -425 -370
rect 2115 -370 2155 -355
rect 235 -550 275 -535
rect 235 -770 245 -550
rect 265 -770 275 -550
rect 235 -785 275 -770
rect 1470 -550 1510 -535
rect 1470 -770 1480 -550
rect 1500 -770 1510 -550
rect 1470 -785 1510 -770
rect -465 -1055 -425 -1040
rect 455 -965 495 -950
rect 455 -1085 465 -965
rect 485 -1085 495 -965
rect 455 -1100 495 -1085
rect 865 -965 905 -950
rect 865 -1085 875 -965
rect 895 -1085 905 -965
rect 865 -1100 905 -1085
rect 2115 -1040 2125 -370
rect 2145 -1040 2155 -370
rect 2115 -1055 2155 -1040
rect 2795 -370 2835 -355
rect 2795 -1040 2805 -370
rect 2825 -1040 2835 -370
rect 2795 -1055 2835 -1040
<< nsubdiff >>
rect -10 2660 30 2675
rect -10 2340 0 2660
rect 20 2340 30 2660
rect -10 2325 30 2340
rect 250 2660 290 2675
rect 250 2340 260 2660
rect 280 2340 290 2660
rect 930 2660 970 2675
rect 250 2325 290 2340
rect 460 2490 500 2505
rect 460 2340 470 2490
rect 490 2340 500 2490
rect 460 2325 500 2340
rect 720 2490 760 2505
rect 720 2340 730 2490
rect 750 2340 760 2490
rect 720 2325 760 2340
rect 930 2340 940 2660
rect 960 2340 970 2660
rect 930 2325 970 2340
rect 1190 2660 1230 2675
rect 1190 2340 1200 2660
rect 1220 2340 1230 2660
rect 1190 2325 1230 2340
rect 1400 2660 1440 2675
rect 1400 2340 1410 2660
rect 1430 2340 1440 2660
rect 1400 2325 1440 2340
rect 1660 2660 1700 2675
rect 1660 2340 1670 2660
rect 1690 2340 1700 2660
rect 1660 2325 1700 2340
rect -1205 2085 -1165 2100
rect -1205 1765 -1195 2085
rect -1175 1765 -1165 2085
rect -1205 1750 -1165 1765
rect -405 2085 -365 2100
rect -405 1765 -395 2085
rect -375 1765 -365 2085
rect -405 1750 -365 1765
rect -80 2085 -40 2100
rect -80 1765 -70 2085
rect -50 1765 -40 2085
rect -80 1750 -40 1765
rect 720 2085 760 2100
rect 720 1765 730 2085
rect 750 1765 760 2085
rect 720 1750 760 1765
rect 930 2085 970 2100
rect 930 1765 940 2085
rect 960 1765 970 2085
rect 930 1750 970 1765
rect 1730 2085 1770 2100
rect 1730 1765 1740 2085
rect 1760 1765 1770 2085
rect 1730 1750 1770 1765
rect 2055 2085 2095 2100
rect 2055 1765 2065 2085
rect 2085 1765 2095 2085
rect 2055 1750 2095 1765
rect 2855 2085 2895 2100
rect 2855 1765 2865 2085
rect 2885 1765 2895 2085
rect 2855 1750 2895 1765
rect 415 1470 455 1485
rect -1175 1420 -1135 1435
rect -1175 850 -1165 1420
rect -1145 850 -1135 1420
rect -1175 835 -1135 850
rect -435 1420 -395 1435
rect -435 850 -425 1420
rect -405 850 -395 1420
rect 415 1250 425 1470
rect 445 1250 455 1470
rect 415 1235 455 1250
rect 825 1470 865 1485
rect 825 1250 835 1470
rect 855 1250 865 1470
rect 825 1235 865 1250
rect 1235 1470 1275 1485
rect 1235 1250 1245 1470
rect 1265 1250 1275 1470
rect 1235 1235 1275 1250
rect 2085 1420 2125 1435
rect -435 835 -395 850
rect 2085 850 2095 1420
rect 2115 850 2125 1420
rect 2085 835 2125 850
rect 2825 1420 2865 1435
rect 2825 850 2835 1420
rect 2855 850 2865 1420
rect 2825 835 2865 850
rect -1175 605 -1135 620
rect -1175 435 -1165 605
rect -1145 435 -1135 605
rect -1175 420 -1135 435
rect -435 605 -395 620
rect -435 435 -425 605
rect -405 435 -395 605
rect 2085 605 2125 620
rect -435 420 -395 435
rect 2085 435 2095 605
rect 2115 435 2125 605
rect 2085 420 2125 435
rect 2825 605 2865 620
rect 2825 435 2835 605
rect 2855 435 2865 605
rect 2825 420 2865 435
<< psubdiffcont >>
rect -135 715 -115 835
rect 605 715 625 835
rect 685 640 705 860
rect 985 640 1005 860
rect 1065 715 1085 835
rect 1805 715 1825 835
rect -135 320 -115 440
rect 605 320 625 440
rect 685 320 705 440
rect 985 320 1005 440
rect 1065 320 1085 440
rect 1805 320 1825 440
rect -1165 -55 -1145 215
rect -425 -55 -405 215
rect 685 -275 705 -55
rect 985 -275 1005 -55
rect 2095 -55 2115 215
rect 2835 -55 2855 215
rect -1135 -1040 -1115 -370
rect -455 -1040 -435 -370
rect 245 -770 265 -550
rect 1480 -770 1500 -550
rect 465 -1085 485 -965
rect 875 -1085 895 -965
rect 2125 -1040 2145 -370
rect 2805 -1040 2825 -370
<< nsubdiffcont >>
rect 0 2340 20 2660
rect 260 2340 280 2660
rect 470 2340 490 2490
rect 730 2340 750 2490
rect 940 2340 960 2660
rect 1200 2340 1220 2660
rect 1410 2340 1430 2660
rect 1670 2340 1690 2660
rect -1195 1765 -1175 2085
rect -395 1765 -375 2085
rect -70 1765 -50 2085
rect 730 1765 750 2085
rect 940 1765 960 2085
rect 1740 1765 1760 2085
rect 2065 1765 2085 2085
rect 2865 1765 2885 2085
rect -1165 850 -1145 1420
rect -425 850 -405 1420
rect 425 1250 445 1470
rect 835 1250 855 1470
rect 1245 1250 1265 1470
rect 2095 850 2115 1420
rect 2835 850 2855 1420
rect -1165 435 -1145 605
rect -425 435 -405 605
rect 2095 435 2115 605
rect 2835 435 2855 605
<< poly >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2705 70 2720
rect 210 2720 250 2730
rect 210 2705 220 2720
rect 60 2700 90 2705
rect 30 2690 90 2700
rect 190 2700 220 2705
rect 240 2700 250 2720
rect 190 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2705 1010 2720
rect 1150 2720 1190 2730
rect 1150 2705 1160 2720
rect 1000 2700 1030 2705
rect 970 2690 1030 2700
rect 1130 2700 1160 2705
rect 1180 2700 1190 2720
rect 1130 2690 1190 2700
rect 1440 2720 1480 2730
rect 1440 2700 1450 2720
rect 1470 2705 1480 2720
rect 1620 2720 1660 2730
rect 1620 2705 1630 2720
rect 1470 2700 1500 2705
rect 1440 2690 1500 2700
rect 1600 2700 1630 2705
rect 1650 2700 1660 2720
rect 1600 2690 1660 2700
rect 70 2675 90 2690
rect 130 2675 150 2690
rect 190 2675 210 2690
rect 1010 2675 1030 2690
rect 1070 2675 1090 2690
rect 1130 2675 1150 2690
rect 1480 2675 1500 2690
rect 1540 2675 1560 2690
rect 1600 2675 1620 2690
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2535 540 2550
rect 680 2550 720 2560
rect 680 2535 690 2550
rect 530 2530 560 2535
rect 500 2520 560 2530
rect 660 2530 690 2535
rect 710 2530 720 2550
rect 660 2520 720 2530
rect 540 2505 560 2520
rect 600 2505 620 2520
rect 660 2505 680 2520
rect 70 2310 90 2325
rect 130 2310 150 2325
rect 190 2310 210 2325
rect 540 2310 560 2325
rect 600 2310 620 2325
rect 660 2310 680 2325
rect 1010 2310 1030 2325
rect 1070 2310 1090 2325
rect 1130 2310 1150 2325
rect 1480 2310 1500 2325
rect 1540 2310 1560 2325
rect 1600 2310 1620 2325
rect 130 2300 169 2310
rect 130 2295 144 2300
rect 139 2280 144 2295
rect 164 2280 169 2300
rect 600 2300 639 2310
rect 600 2295 614 2300
rect 139 2270 169 2280
rect 609 2280 614 2295
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1090 2310
rect 1051 2280 1056 2300
rect 1076 2295 1090 2300
rect 1521 2300 1560 2310
rect 1076 2280 1081 2295
rect 1051 2270 1081 2280
rect 1521 2280 1526 2300
rect 1546 2295 1560 2300
rect 1546 2280 1551 2295
rect 1521 2270 1551 2280
rect -1165 2145 -1125 2155
rect -1165 2125 -1155 2145
rect -1135 2130 -1125 2145
rect -445 2145 -405 2155
rect -445 2130 -435 2145
rect -1135 2125 -1105 2130
rect -1165 2115 -1105 2125
rect -465 2125 -435 2130
rect -415 2125 -405 2145
rect -465 2115 -405 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2130 0 2145
rect 680 2145 720 2155
rect 680 2130 690 2145
rect -10 2125 20 2130
rect -40 2115 20 2125
rect 660 2125 690 2130
rect 710 2125 720 2145
rect 660 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2130 1010 2145
rect 1690 2145 1730 2155
rect 1690 2130 1700 2145
rect 1000 2125 1030 2130
rect 970 2115 1030 2125
rect 1670 2125 1700 2130
rect 1720 2125 1730 2145
rect 1670 2115 1730 2125
rect 2095 2145 2135 2155
rect 2095 2125 2105 2145
rect 2125 2130 2135 2145
rect 2815 2145 2855 2155
rect 2815 2130 2825 2145
rect 2125 2125 2155 2130
rect 2095 2115 2155 2125
rect 2795 2125 2825 2130
rect 2845 2125 2855 2145
rect 2795 2115 2855 2125
rect -1125 2100 -1105 2115
rect -1065 2100 -1045 2115
rect -1005 2100 -985 2115
rect -945 2100 -925 2115
rect -885 2100 -865 2115
rect -825 2100 -805 2115
rect -765 2100 -745 2115
rect -705 2100 -685 2115
rect -645 2100 -625 2115
rect -585 2100 -565 2115
rect -525 2100 -505 2115
rect -465 2100 -445 2115
rect 0 2100 20 2115
rect 60 2100 80 2115
rect 120 2100 140 2115
rect 180 2100 200 2115
rect 240 2100 260 2115
rect 300 2100 320 2115
rect 360 2100 380 2115
rect 420 2100 440 2115
rect 480 2100 500 2115
rect 540 2100 560 2115
rect 600 2100 620 2115
rect 660 2100 680 2115
rect 1010 2100 1030 2115
rect 1070 2100 1090 2115
rect 1130 2100 1150 2115
rect 1190 2100 1210 2115
rect 1250 2100 1270 2115
rect 1310 2100 1330 2115
rect 1370 2100 1390 2115
rect 1430 2100 1450 2115
rect 1490 2100 1510 2115
rect 1550 2100 1570 2115
rect 1610 2100 1630 2115
rect 1670 2100 1690 2115
rect 2135 2100 2155 2115
rect 2195 2100 2215 2115
rect 2255 2100 2275 2115
rect 2315 2100 2335 2115
rect 2375 2100 2395 2115
rect 2435 2100 2455 2115
rect 2495 2100 2515 2115
rect 2555 2100 2575 2115
rect 2615 2100 2635 2115
rect 2675 2100 2695 2115
rect 2735 2100 2755 2115
rect 2795 2100 2815 2115
rect -1125 1735 -1105 1750
rect -1065 1740 -1045 1750
rect -1005 1740 -985 1750
rect -945 1740 -925 1750
rect -885 1740 -865 1750
rect -825 1740 -805 1750
rect -765 1740 -745 1750
rect -705 1740 -685 1750
rect -645 1740 -625 1750
rect -585 1740 -565 1750
rect -525 1740 -505 1750
rect -1065 1725 -505 1740
rect -465 1735 -445 1750
rect 0 1735 20 1750
rect 60 1740 80 1750
rect 120 1740 140 1750
rect 180 1740 200 1750
rect 240 1740 260 1750
rect 300 1740 320 1750
rect 360 1740 380 1750
rect 420 1740 440 1750
rect 480 1740 500 1750
rect 540 1740 560 1750
rect 600 1740 620 1750
rect 60 1725 620 1740
rect 660 1735 680 1750
rect 1010 1735 1030 1750
rect 1070 1740 1090 1750
rect 1130 1740 1150 1750
rect 1190 1740 1210 1750
rect 1250 1740 1270 1750
rect 1310 1740 1330 1750
rect 1370 1740 1390 1750
rect 1430 1740 1450 1750
rect 1490 1740 1510 1750
rect 1550 1740 1570 1750
rect 1610 1740 1630 1750
rect 1070 1725 1630 1740
rect 1670 1735 1690 1750
rect 2135 1735 2155 1750
rect 2195 1740 2215 1750
rect 2255 1740 2275 1750
rect 2315 1740 2335 1750
rect 2375 1740 2395 1750
rect 2435 1740 2455 1750
rect 2495 1740 2515 1750
rect 2555 1740 2575 1750
rect 2615 1740 2635 1750
rect 2675 1740 2695 1750
rect 2735 1740 2755 1750
rect 2195 1725 2755 1740
rect 2795 1735 2815 1750
rect -705 1630 -685 1725
rect 420 1675 440 1725
rect 1250 1675 1270 1725
rect 410 1665 450 1675
rect 410 1645 420 1665
rect 440 1645 450 1665
rect 410 1635 450 1645
rect 1240 1665 1280 1675
rect 1240 1645 1250 1665
rect 1270 1645 1280 1665
rect 1240 1635 1280 1645
rect 2375 1630 2395 1725
rect -715 1620 -675 1630
rect -715 1600 -705 1620
rect -685 1600 -675 1620
rect -715 1590 -675 1600
rect 2365 1620 2405 1630
rect 2365 1600 2375 1620
rect 2395 1600 2405 1620
rect 2365 1590 2405 1600
rect 455 1570 495 1580
rect 455 1550 465 1570
rect 485 1555 495 1570
rect 785 1570 825 1580
rect 785 1555 795 1570
rect 485 1550 510 1555
rect 455 1540 510 1550
rect -1135 1480 -1095 1490
rect -1135 1460 -1125 1480
rect -1105 1465 -1095 1480
rect -475 1480 -435 1490
rect 495 1485 510 1540
rect 770 1550 795 1555
rect 815 1550 825 1570
rect 770 1540 825 1550
rect 865 1570 905 1580
rect 865 1550 875 1570
rect 895 1555 905 1570
rect 1195 1570 1235 1580
rect 1195 1555 1205 1570
rect 895 1550 920 1555
rect 865 1540 920 1550
rect 550 1485 565 1500
rect 605 1485 620 1500
rect 660 1485 675 1500
rect 715 1485 730 1500
rect 770 1485 785 1540
rect 905 1485 920 1540
rect 1180 1550 1205 1555
rect 1225 1550 1235 1570
rect 1180 1540 1235 1550
rect 960 1485 975 1500
rect 1015 1485 1030 1500
rect 1070 1485 1085 1500
rect 1125 1485 1140 1500
rect 1180 1485 1195 1540
rect -475 1465 -465 1480
rect -1105 1460 -1080 1465
rect -1135 1450 -1080 1460
rect -490 1460 -465 1465
rect -445 1460 -435 1480
rect -490 1450 -435 1460
rect -1095 1435 -1080 1450
rect -1040 1435 -1025 1450
rect -985 1435 -970 1450
rect -930 1435 -915 1450
rect -875 1435 -860 1450
rect -820 1435 -805 1450
rect -765 1435 -750 1450
rect -710 1435 -695 1450
rect -655 1435 -640 1450
rect -600 1435 -585 1450
rect -545 1435 -530 1450
rect -490 1435 -475 1450
rect 2125 1480 2165 1490
rect 2125 1460 2135 1480
rect 2155 1465 2165 1480
rect 2785 1480 2825 1490
rect 2785 1465 2795 1480
rect 2155 1460 2180 1465
rect 2125 1450 2180 1460
rect 2770 1460 2795 1465
rect 2815 1460 2825 1480
rect 2770 1450 2825 1460
rect 2165 1435 2180 1450
rect 2220 1435 2235 1450
rect 2275 1435 2290 1450
rect 2330 1435 2345 1450
rect 2385 1435 2400 1450
rect 2440 1435 2455 1450
rect 2495 1435 2510 1450
rect 2550 1435 2565 1450
rect 2605 1435 2620 1450
rect 2660 1435 2675 1450
rect 2715 1435 2730 1450
rect 2770 1435 2785 1450
rect 495 1220 510 1235
rect 550 1220 565 1235
rect 605 1225 620 1235
rect 660 1225 675 1235
rect 550 1210 582 1220
rect 605 1210 675 1225
rect 715 1220 730 1235
rect 770 1220 785 1235
rect 905 1220 920 1235
rect 960 1220 975 1235
rect 1015 1225 1030 1235
rect 1070 1225 1085 1235
rect 698 1210 730 1220
rect 960 1210 992 1220
rect 1015 1210 1085 1225
rect 1125 1220 1140 1235
rect 1180 1220 1195 1235
rect 1108 1210 1140 1220
rect 552 1190 557 1210
rect 577 1190 582 1210
rect 552 1180 582 1190
rect 620 1190 630 1210
rect 650 1190 660 1210
rect 620 1180 660 1190
rect 698 1190 703 1210
rect 723 1190 728 1210
rect 698 1180 728 1190
rect 962 1190 967 1210
rect 987 1190 992 1210
rect 962 1180 992 1190
rect 1030 1190 1040 1210
rect 1060 1190 1070 1210
rect 1030 1180 1070 1190
rect 1108 1190 1113 1210
rect 1133 1190 1138 1210
rect 1108 1180 1138 1190
rect 145 945 175 955
rect 145 925 150 945
rect 170 925 175 945
rect 1515 945 1545 955
rect 145 915 175 925
rect 795 920 835 930
rect 155 875 170 915
rect 795 900 805 920
rect 825 900 835 920
rect 1515 925 1520 945
rect 1540 925 1545 945
rect 1515 915 1545 925
rect 755 875 770 890
rect 795 885 880 900
rect 810 875 825 885
rect 865 875 880 885
rect 920 875 935 890
rect 1520 875 1535 915
rect -65 850 -50 865
rect -10 860 500 875
rect -10 850 5 860
rect 45 850 60 860
rect 100 850 115 860
rect 155 850 170 860
rect 210 850 225 860
rect 265 850 280 860
rect 320 850 335 860
rect 375 850 390 860
rect 430 850 445 860
rect 485 850 500 860
rect 540 850 555 865
rect -1095 820 -1080 835
rect -1040 825 -1025 835
rect -985 825 -970 835
rect -930 825 -915 835
rect -875 825 -860 835
rect -820 825 -805 835
rect -765 825 -750 835
rect -710 825 -695 835
rect -655 825 -640 835
rect -600 825 -585 835
rect -545 825 -530 835
rect -1040 810 -530 825
rect -490 820 -475 835
rect -795 720 -775 810
rect -805 710 -765 720
rect -805 690 -795 710
rect -775 690 -765 710
rect -805 680 -765 690
rect -65 685 -50 700
rect -10 685 5 700
rect 45 685 60 700
rect 100 685 115 700
rect 155 685 170 700
rect 210 685 225 700
rect 265 685 280 700
rect 320 685 335 700
rect 375 685 390 700
rect 430 685 445 700
rect 485 685 500 700
rect 540 685 555 700
rect -100 675 -50 685
rect -1145 665 -1105 675
rect -1145 645 -1135 665
rect -1115 650 -1105 665
rect -465 665 -425 675
rect -465 650 -455 665
rect -1115 645 -1080 650
rect -1145 635 -1080 645
rect -490 645 -455 650
rect -435 645 -425 665
rect -100 655 -95 675
rect -75 670 -50 675
rect 540 675 590 685
rect 540 670 565 675
rect -75 655 -70 670
rect -100 645 -70 655
rect 560 655 565 670
rect 585 655 590 675
rect 560 645 590 655
rect -490 635 -425 645
rect -1095 620 -1080 635
rect -1040 620 -1025 635
rect -985 620 -970 635
rect -930 620 -915 635
rect -875 620 -860 635
rect -820 620 -805 635
rect -765 620 -750 635
rect -710 620 -695 635
rect -655 620 -640 635
rect -600 620 -585 635
rect -545 620 -530 635
rect -490 620 -475 635
rect 1135 850 1150 865
rect 1190 860 1700 875
rect 1190 850 1205 860
rect 1245 850 1260 860
rect 1300 850 1315 860
rect 1355 850 1370 860
rect 1410 850 1425 860
rect 1465 850 1480 860
rect 1520 850 1535 860
rect 1575 850 1590 860
rect 1630 850 1645 860
rect 1685 850 1700 860
rect 1740 850 1755 865
rect 2165 820 2180 835
rect 2220 825 2235 835
rect 2275 825 2290 835
rect 2330 825 2345 835
rect 2385 825 2400 835
rect 2440 825 2455 835
rect 2495 825 2510 835
rect 2550 825 2565 835
rect 2605 825 2620 835
rect 2660 825 2675 835
rect 2715 825 2730 835
rect 2220 810 2730 825
rect 2770 820 2785 835
rect 2465 720 2485 810
rect 2455 710 2495 720
rect 1135 685 1150 700
rect 1190 685 1205 700
rect 1245 685 1260 700
rect 1300 685 1315 700
rect 1355 685 1370 700
rect 1410 685 1425 700
rect 1465 685 1480 700
rect 1520 685 1535 700
rect 1575 685 1590 700
rect 1630 685 1645 700
rect 1685 685 1700 700
rect 1740 685 1755 700
rect 2455 690 2465 710
rect 2485 690 2495 710
rect 1100 675 1150 685
rect 1100 655 1105 675
rect 1125 670 1150 675
rect 1740 675 1790 685
rect 2455 680 2495 690
rect 1740 670 1765 675
rect 1125 655 1130 670
rect 1100 645 1130 655
rect 1760 655 1765 670
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 2115 665 2155 675
rect 2115 645 2125 665
rect 2145 650 2155 665
rect 2795 665 2835 675
rect 2795 650 2805 665
rect 2145 645 2180 650
rect 2115 635 2180 645
rect 2770 645 2805 650
rect 2825 645 2835 665
rect 2770 635 2835 645
rect 755 610 770 625
rect 810 610 825 625
rect 865 610 880 625
rect 920 610 935 625
rect 2165 620 2180 635
rect 2220 620 2235 635
rect 2275 620 2290 635
rect 2330 620 2345 635
rect 2385 620 2400 635
rect 2440 620 2455 635
rect 2495 620 2510 635
rect 2550 620 2565 635
rect 2605 620 2620 635
rect 2660 620 2675 635
rect 2715 620 2730 635
rect 2770 620 2785 635
rect 715 600 770 610
rect 715 580 725 600
rect 745 595 770 600
rect 920 600 975 610
rect 920 595 945 600
rect 745 580 755 595
rect 715 570 755 580
rect 935 580 945 595
rect 965 580 975 600
rect 935 570 975 580
rect 145 545 175 555
rect 145 525 150 545
rect 170 525 175 545
rect 145 515 175 525
rect 795 545 825 555
rect 795 525 800 545
rect 820 525 825 545
rect 795 515 825 525
rect 155 480 170 515
rect 715 500 755 510
rect 715 480 725 500
rect 745 485 755 500
rect 745 480 770 485
rect -65 455 -50 470
rect -10 465 500 480
rect 715 470 770 480
rect -10 455 5 465
rect 45 455 60 465
rect 100 455 115 465
rect 155 455 170 465
rect 210 455 225 465
rect 265 455 280 465
rect 320 455 335 465
rect 375 455 390 465
rect 430 455 445 465
rect 485 455 500 465
rect 540 455 555 470
rect 755 455 770 470
rect 810 455 825 515
rect 865 545 895 555
rect 865 525 870 545
rect 890 525 895 545
rect 865 515 895 525
rect 1515 545 1545 555
rect 1515 525 1520 545
rect 1540 525 1545 545
rect 1515 515 1545 525
rect 865 455 880 515
rect 935 500 975 510
rect 935 485 945 500
rect 920 480 945 485
rect 965 480 975 500
rect 1520 480 1535 515
rect 920 470 975 480
rect 920 455 935 470
rect 1135 455 1150 470
rect 1190 465 1700 480
rect 1190 455 1205 465
rect 1245 455 1260 465
rect 1300 455 1315 465
rect 1355 455 1370 465
rect 1410 455 1425 465
rect 1465 455 1480 465
rect 1520 455 1535 465
rect 1575 455 1590 465
rect 1630 455 1645 465
rect 1685 455 1700 465
rect 1740 455 1755 470
rect -1095 405 -1080 420
rect -1040 410 -1025 420
rect -985 410 -970 420
rect -930 410 -915 420
rect -875 410 -860 420
rect -820 410 -805 420
rect -765 410 -750 420
rect -710 410 -695 420
rect -655 410 -640 420
rect -600 410 -585 420
rect -545 410 -530 420
rect -1040 395 -530 410
rect -490 405 -475 420
rect -740 345 -720 395
rect -750 335 -710 345
rect -750 315 -740 335
rect -720 315 -710 335
rect -750 305 -710 315
rect 2165 405 2180 420
rect 2220 410 2235 420
rect 2275 410 2290 420
rect 2330 410 2345 420
rect 2385 410 2400 420
rect 2440 410 2455 420
rect 2495 410 2510 420
rect 2550 410 2565 420
rect 2605 410 2620 420
rect 2660 410 2675 420
rect 2715 410 2730 420
rect 2220 395 2730 410
rect 2770 405 2785 420
rect 2410 345 2430 395
rect 2400 335 2440 345
rect 2400 315 2410 335
rect 2430 315 2440 335
rect 2400 305 2440 315
rect -740 255 -720 305
rect -65 290 -50 305
rect -10 290 5 305
rect 45 290 60 305
rect 100 290 115 305
rect 155 290 170 305
rect 210 290 225 305
rect 265 290 280 305
rect 320 290 335 305
rect 375 290 390 305
rect 430 290 445 305
rect 485 290 500 305
rect 540 290 555 305
rect 755 290 770 305
rect 810 290 825 305
rect 865 290 880 305
rect 920 290 935 305
rect 1135 290 1150 305
rect 1190 290 1205 305
rect 1245 290 1260 305
rect 1300 290 1315 305
rect 1355 290 1370 305
rect 1410 290 1425 305
rect 1465 290 1480 305
rect 1520 290 1535 305
rect 1575 290 1590 305
rect 1630 290 1645 305
rect 1685 290 1700 305
rect 1740 290 1755 305
rect -100 280 -50 290
rect -100 260 -95 280
rect -75 275 -50 280
rect 540 280 630 290
rect 540 275 605 280
rect -75 260 -70 275
rect -1095 230 -1080 245
rect -1040 240 -530 255
rect -100 250 -70 260
rect 600 260 605 275
rect 625 260 630 280
rect 600 250 630 260
rect 1060 280 1150 290
rect 1060 260 1065 280
rect 1085 275 1150 280
rect 1740 280 1790 290
rect 1740 275 1765 280
rect 1085 260 1090 275
rect 1060 250 1090 260
rect 1760 260 1765 275
rect 1785 260 1790 280
rect 1760 250 1790 260
rect 2410 255 2430 305
rect -1040 230 -1025 240
rect -985 230 -970 240
rect -930 230 -915 240
rect -875 230 -860 240
rect -820 230 -805 240
rect -765 230 -750 240
rect -710 230 -695 240
rect -655 230 -640 240
rect -600 230 -585 240
rect -545 230 -530 240
rect -490 230 -475 245
rect 2165 230 2180 245
rect 2220 240 2730 255
rect 2220 230 2235 240
rect 2275 230 2290 240
rect 2330 230 2345 240
rect 2385 230 2400 240
rect 2440 230 2455 240
rect 2495 230 2510 240
rect 2550 230 2565 240
rect 2605 230 2620 240
rect 2660 230 2675 240
rect 2715 230 2730 240
rect 2770 230 2785 245
rect 830 10 860 20
rect 830 -10 835 10
rect 855 -10 860 10
rect 830 -15 860 -10
rect 755 -40 770 -25
rect 810 -30 880 -15
rect 810 -40 825 -30
rect 865 -40 880 -30
rect 920 -40 935 -25
rect -1095 -85 -1080 -70
rect -1040 -85 -1025 -70
rect -985 -85 -970 -70
rect -930 -85 -915 -70
rect -875 -85 -860 -70
rect -820 -85 -805 -70
rect -765 -85 -750 -70
rect -710 -85 -695 -70
rect -655 -85 -640 -70
rect -600 -85 -585 -70
rect -545 -85 -530 -70
rect -490 -85 -475 -70
rect -1145 -95 -1080 -85
rect -1145 -115 -1135 -95
rect -1115 -100 -1080 -95
rect -490 -95 -425 -85
rect -490 -100 -455 -95
rect -1115 -115 -1105 -100
rect -1145 -125 -1105 -115
rect -465 -115 -455 -100
rect -435 -115 -425 -95
rect -465 -125 -425 -115
rect -805 -250 -765 -240
rect -805 -270 -795 -250
rect -775 -270 -765 -250
rect -805 -280 -765 -270
rect -795 -330 -775 -280
rect 2165 -85 2180 -70
rect 2220 -85 2235 -70
rect 2275 -85 2290 -70
rect 2330 -85 2345 -70
rect 2385 -85 2400 -70
rect 2440 -85 2455 -70
rect 2495 -85 2510 -70
rect 2550 -85 2565 -70
rect 2605 -85 2620 -70
rect 2660 -85 2675 -70
rect 2715 -85 2730 -70
rect 2770 -85 2785 -70
rect 2115 -95 2180 -85
rect 2115 -115 2125 -95
rect 2145 -100 2180 -95
rect 2770 -95 2835 -85
rect 2770 -100 2805 -95
rect 2145 -115 2155 -100
rect 2115 -125 2155 -115
rect 2795 -115 2805 -100
rect 2825 -115 2835 -95
rect 2795 -125 2835 -115
rect 2455 -250 2495 -240
rect 2455 -270 2465 -250
rect 2485 -270 2495 -250
rect 2455 -280 2495 -270
rect 755 -305 770 -290
rect 810 -305 825 -290
rect 865 -305 880 -290
rect 920 -305 935 -290
rect 715 -315 770 -305
rect -1065 -355 -1005 -340
rect -965 -345 -605 -330
rect 715 -335 725 -315
rect 745 -320 770 -315
rect 920 -315 975 -305
rect 920 -320 945 -315
rect 745 -335 755 -320
rect -965 -355 -905 -345
rect -865 -355 -805 -345
rect -765 -355 -705 -345
rect -665 -355 -605 -345
rect -565 -355 -505 -340
rect 715 -345 755 -335
rect 935 -335 945 -320
rect 965 -335 975 -315
rect 2465 -330 2485 -280
rect 935 -345 975 -335
rect 2195 -355 2255 -340
rect 2295 -345 2655 -330
rect 2295 -355 2355 -345
rect 2395 -355 2455 -345
rect 2495 -355 2555 -345
rect 2595 -355 2655 -345
rect 2695 -355 2755 -340
rect 1350 -430 1390 -420
rect 445 -440 475 -430
rect 445 -460 450 -440
rect 470 -460 475 -440
rect 1350 -450 1360 -430
rect 1380 -450 1390 -430
rect 1350 -460 1390 -450
rect 445 -470 475 -460
rect 450 -510 470 -470
rect 315 -535 330 -520
rect 370 -525 1320 -510
rect 370 -535 385 -525
rect 425 -535 440 -525
rect 480 -535 495 -525
rect 535 -535 550 -525
rect 590 -535 605 -525
rect 645 -535 660 -525
rect 700 -535 715 -525
rect 755 -535 770 -525
rect 810 -535 825 -525
rect 865 -535 880 -525
rect 920 -535 935 -525
rect 975 -535 990 -525
rect 1030 -535 1045 -525
rect 1085 -535 1100 -525
rect 1140 -535 1155 -525
rect 1195 -535 1210 -525
rect 1250 -535 1265 -525
rect 1305 -535 1320 -525
rect 1360 -535 1375 -460
rect 1415 -535 1430 -520
rect 315 -800 330 -785
rect 370 -800 385 -785
rect 425 -800 440 -785
rect 480 -800 495 -785
rect 535 -800 550 -785
rect 590 -800 605 -785
rect 645 -800 660 -785
rect 700 -800 715 -785
rect 755 -800 770 -785
rect 810 -800 825 -785
rect 865 -800 880 -785
rect 920 -800 935 -785
rect 975 -800 990 -785
rect 1030 -800 1045 -785
rect 1085 -800 1100 -785
rect 1140 -800 1155 -785
rect 1195 -800 1210 -785
rect 1250 -800 1265 -785
rect 1305 -800 1320 -785
rect 1360 -800 1375 -785
rect 1415 -800 1430 -785
rect 265 -810 330 -800
rect 265 -830 275 -810
rect 295 -815 330 -810
rect 1415 -810 1470 -800
rect 1415 -815 1440 -810
rect 295 -830 305 -815
rect 265 -840 305 -830
rect 1430 -830 1440 -815
rect 1460 -830 1470 -810
rect 1430 -840 1470 -830
rect 660 -905 700 -895
rect 660 -925 670 -905
rect 690 -925 700 -905
rect 1130 -905 1170 -895
rect 1130 -925 1140 -905
rect 1160 -925 1170 -905
rect 535 -950 550 -935
rect 590 -940 770 -925
rect 1130 -935 1170 -925
rect 590 -950 605 -940
rect 645 -950 660 -940
rect 700 -950 715 -940
rect 755 -950 770 -940
rect 810 -950 825 -935
rect 1000 -950 1300 -935
rect -1065 -1070 -1005 -1055
rect -965 -1070 -905 -1055
rect -865 -1070 -805 -1055
rect -765 -1070 -705 -1055
rect -665 -1070 -605 -1055
rect -565 -1070 -505 -1055
rect -1105 -1080 -1005 -1070
rect -1105 -1100 -1095 -1080
rect -1075 -1085 -1005 -1080
rect -565 -1080 -465 -1070
rect -565 -1085 -495 -1080
rect -1075 -1100 -1065 -1085
rect -1105 -1110 -1065 -1100
rect -505 -1100 -495 -1085
rect -475 -1100 -465 -1080
rect 2195 -1070 2255 -1055
rect 2295 -1070 2355 -1055
rect 2395 -1070 2455 -1055
rect 2495 -1070 2555 -1055
rect 2595 -1070 2655 -1055
rect 2695 -1070 2755 -1055
rect 2155 -1080 2255 -1070
rect 2155 -1100 2165 -1080
rect 2185 -1085 2255 -1080
rect 2695 -1080 2795 -1070
rect 2695 -1085 2765 -1080
rect 2185 -1100 2195 -1085
rect -505 -1110 -465 -1100
rect 535 -1115 550 -1100
rect 590 -1115 605 -1100
rect 645 -1115 660 -1100
rect 700 -1115 715 -1100
rect 755 -1115 770 -1100
rect 810 -1115 825 -1100
rect 1000 -1115 1300 -1100
rect 2155 -1110 2195 -1100
rect 2755 -1100 2765 -1085
rect 2785 -1100 2795 -1080
rect 2755 -1110 2795 -1100
rect 500 -1125 550 -1115
rect 500 -1145 505 -1125
rect 525 -1130 550 -1125
rect 810 -1125 860 -1115
rect 810 -1130 835 -1125
rect 525 -1145 530 -1130
rect 500 -1155 530 -1145
rect 830 -1145 835 -1130
rect 855 -1145 860 -1125
rect 830 -1155 860 -1145
<< polycont >>
rect 40 2700 60 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1160 2700 1180 2720
rect 1450 2700 1470 2720
rect 1630 2700 1650 2720
rect 510 2530 530 2550
rect 690 2530 710 2550
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1526 2280 1546 2300
rect -1155 2125 -1135 2145
rect -435 2125 -415 2145
rect -30 2125 -10 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1700 2125 1720 2145
rect 2105 2125 2125 2145
rect 2825 2125 2845 2145
rect 420 1645 440 1665
rect 1250 1645 1270 1665
rect -705 1600 -685 1620
rect 2375 1600 2395 1620
rect 465 1550 485 1570
rect -1125 1460 -1105 1480
rect 795 1550 815 1570
rect 875 1550 895 1570
rect 1205 1550 1225 1570
rect -465 1460 -445 1480
rect 2135 1460 2155 1480
rect 2795 1460 2815 1480
rect 557 1190 577 1210
rect 630 1190 650 1210
rect 703 1190 723 1210
rect 967 1190 987 1210
rect 1040 1190 1060 1210
rect 1113 1190 1133 1210
rect 150 925 170 945
rect 805 900 825 920
rect 1520 925 1540 945
rect -795 690 -775 710
rect -1135 645 -1115 665
rect -455 645 -435 665
rect -95 655 -75 675
rect 565 655 585 675
rect 2465 690 2485 710
rect 1105 655 1125 675
rect 1765 655 1785 675
rect 2125 645 2145 665
rect 2805 645 2825 665
rect 725 580 745 600
rect 945 580 965 600
rect 150 525 170 545
rect 800 525 820 545
rect 725 480 745 500
rect 870 525 890 545
rect 1520 525 1540 545
rect 945 480 965 500
rect -740 315 -720 335
rect 2410 315 2430 335
rect -95 260 -75 280
rect 605 260 625 280
rect 1065 260 1085 280
rect 1765 260 1785 280
rect 835 -10 855 10
rect -1135 -115 -1115 -95
rect -455 -115 -435 -95
rect -795 -270 -775 -250
rect 2125 -115 2145 -95
rect 2805 -115 2825 -95
rect 2465 -270 2485 -250
rect 725 -335 745 -315
rect 945 -335 965 -315
rect 450 -460 470 -440
rect 1360 -450 1380 -430
rect 275 -830 295 -810
rect 1440 -830 1460 -810
rect 670 -925 690 -905
rect 1140 -925 1160 -905
rect -1095 -1100 -1075 -1080
rect -495 -1100 -475 -1080
rect 2165 -1100 2185 -1080
rect 2765 -1100 2785 -1080
rect 505 -1145 525 -1125
rect 835 -1145 855 -1125
<< xpolycontact >>
rect -1501 1170 -1360 1390
rect -1501 825 -1360 1045
rect 3050 1170 3191 1390
rect 3050 825 3191 1045
rect -1490 297 -1455 517
rect -1490 -85 -1455 138
rect -1430 297 -1395 517
rect -1430 -85 -1395 138
rect -1370 297 -1335 517
rect -1370 -85 -1335 138
rect -1310 297 -1275 517
rect 2965 297 3000 517
rect -1310 -85 -1275 138
rect 2965 -85 3000 138
rect 3025 297 3060 517
rect 3025 -85 3060 138
rect 3085 297 3120 517
rect 3085 -85 3120 138
rect 3145 297 3180 517
rect 3145 -85 3180 138
rect -1290 -638 -1255 -415
rect -1290 -1105 -1255 -885
rect -1230 -638 -1195 -415
rect -1230 -1105 -1195 -885
rect 2885 -638 2920 -415
rect 2885 -1105 2920 -885
rect 2945 -638 2980 -415
rect 2945 -1105 2980 -885
<< ppolyres >>
rect -1501 1045 -1360 1170
rect 3050 1045 3191 1170
<< xpolyres >>
rect -1490 138 -1455 297
rect -1430 138 -1395 297
rect -1370 138 -1335 297
rect -1310 138 -1275 297
rect 2965 138 3000 297
rect 3025 138 3060 297
rect 3085 138 3120 297
rect 3145 138 3180 297
rect -1290 -885 -1255 -638
rect -1230 -885 -1195 -638
rect 2885 -885 2920 -638
rect 2945 -885 2980 -638
<< locali >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2710 70 2720
rect 210 2720 250 2730
rect 210 2710 220 2720
rect 60 2700 220 2710
rect 240 2700 250 2720
rect 30 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2700 1010 2720
rect 970 2690 1010 2700
rect 1035 2720 1065 2730
rect 1035 2700 1040 2720
rect 1060 2700 1065 2720
rect 35 2670 65 2690
rect -5 2660 65 2670
rect -5 2340 0 2660
rect 20 2340 40 2660
rect 60 2340 65 2660
rect -5 2330 65 2340
rect 95 2660 125 2670
rect 95 2340 100 2660
rect 120 2340 125 2660
rect 95 2330 125 2340
rect 155 2660 185 2690
rect 155 2340 160 2660
rect 180 2340 185 2660
rect 155 2330 185 2340
rect 215 2670 245 2690
rect 975 2670 1005 2690
rect 215 2660 285 2670
rect 215 2340 220 2660
rect 240 2340 260 2660
rect 280 2340 285 2660
rect 935 2660 1005 2670
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2530 540 2550
rect 500 2520 540 2530
rect 560 2550 600 2560
rect 560 2530 570 2550
rect 590 2530 600 2550
rect 560 2520 600 2530
rect 625 2550 655 2560
rect 625 2530 630 2550
rect 650 2530 655 2550
rect 505 2500 535 2520
rect 215 2330 285 2340
rect 465 2490 535 2500
rect 465 2340 470 2490
rect 490 2340 510 2490
rect 530 2340 535 2490
rect 465 2330 535 2340
rect 565 2490 595 2520
rect 565 2340 570 2490
rect 590 2340 595 2490
rect 565 2330 595 2340
rect 625 2490 655 2530
rect 680 2550 720 2560
rect 680 2530 690 2550
rect 710 2530 720 2550
rect 680 2520 720 2530
rect 625 2340 630 2490
rect 650 2340 655 2490
rect 625 2330 655 2340
rect 685 2500 715 2520
rect 685 2490 755 2500
rect 685 2340 690 2490
rect 710 2340 730 2490
rect 750 2340 755 2490
rect 685 2330 755 2340
rect 935 2340 940 2660
rect 960 2340 980 2660
rect 1000 2340 1005 2660
rect 935 2330 1005 2340
rect 1035 2660 1065 2700
rect 1090 2720 1130 2730
rect 1090 2700 1100 2720
rect 1120 2700 1130 2720
rect 1090 2690 1130 2700
rect 1150 2720 1190 2730
rect 1150 2700 1160 2720
rect 1180 2700 1190 2720
rect 1150 2690 1190 2700
rect 1440 2720 1480 2730
rect 1440 2700 1450 2720
rect 1470 2710 1480 2720
rect 1620 2720 1660 2730
rect 1620 2710 1630 2720
rect 1470 2700 1630 2710
rect 1650 2700 1660 2720
rect 1440 2690 1660 2700
rect 1035 2340 1040 2660
rect 1060 2340 1065 2660
rect 1035 2330 1065 2340
rect 1095 2660 1125 2690
rect 1095 2340 1100 2660
rect 1120 2340 1125 2660
rect 1095 2330 1125 2340
rect 1155 2670 1185 2690
rect 1445 2670 1475 2690
rect 1155 2660 1225 2670
rect 1155 2340 1160 2660
rect 1180 2340 1200 2660
rect 1220 2340 1225 2660
rect 1155 2330 1225 2340
rect 1405 2660 1475 2670
rect 1405 2340 1410 2660
rect 1430 2340 1450 2660
rect 1470 2340 1475 2660
rect 1405 2330 1475 2340
rect 1505 2660 1535 2690
rect 1625 2670 1655 2690
rect 1505 2340 1510 2660
rect 1530 2340 1535 2660
rect 1505 2330 1535 2340
rect 1565 2660 1595 2670
rect 1565 2340 1570 2660
rect 1590 2340 1595 2660
rect 1565 2330 1595 2340
rect 1625 2660 1695 2670
rect 1625 2340 1630 2660
rect 1650 2340 1670 2660
rect 1690 2340 1695 2660
rect 1625 2330 1695 2340
rect 95 2310 115 2330
rect 1575 2310 1595 2330
rect 75 2300 115 2310
rect 75 2280 85 2300
rect 105 2280 115 2300
rect 75 2270 115 2280
rect 139 2300 169 2310
rect 139 2280 144 2300
rect 164 2280 169 2300
rect 139 2270 169 2280
rect 609 2300 639 2310
rect 609 2280 614 2300
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1521 2300 1551 2310
rect 1521 2280 1526 2300
rect 1546 2280 1551 2300
rect 1521 2270 1551 2280
rect 1575 2300 1615 2310
rect 1575 2280 1585 2300
rect 1605 2280 1615 2300
rect 1575 2270 1615 2280
rect -1165 2145 -1125 2155
rect -1165 2125 -1155 2145
rect -1135 2135 -1125 2145
rect -800 2145 -770 2155
rect -800 2135 -795 2145
rect -1135 2125 -795 2135
rect -775 2135 -770 2145
rect -445 2145 -405 2155
rect -445 2135 -435 2145
rect -775 2125 -435 2135
rect -415 2125 -405 2145
rect -1165 2115 -405 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2135 0 2145
rect 680 2145 720 2155
rect 680 2135 690 2145
rect -10 2125 690 2135
rect 710 2125 720 2145
rect -40 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2135 1010 2145
rect 1690 2145 1730 2155
rect 1690 2135 1700 2145
rect 1000 2125 1700 2135
rect 1720 2125 1730 2145
rect 970 2115 1730 2125
rect 2095 2145 2135 2155
rect 2095 2125 2105 2145
rect 2125 2135 2135 2145
rect 2460 2145 2490 2155
rect 2460 2135 2465 2145
rect 2125 2125 2465 2135
rect 2485 2135 2490 2145
rect 2815 2145 2855 2155
rect 2815 2135 2825 2145
rect 2485 2125 2825 2135
rect 2845 2125 2855 2145
rect 2095 2115 2855 2125
rect -1160 2095 -1130 2115
rect -1200 2085 -1130 2095
rect -1200 1765 -1195 2085
rect -1175 1765 -1155 2085
rect -1135 1765 -1130 2085
rect -1200 1755 -1130 1765
rect -1100 2085 -1070 2095
rect -1100 1765 -1095 2085
rect -1075 1765 -1070 2085
rect -1100 1740 -1070 1765
rect -1040 2085 -1010 2115
rect -1040 1765 -1035 2085
rect -1015 1765 -1010 2085
rect -1040 1755 -1010 1765
rect -980 2085 -950 2095
rect -980 1765 -975 2085
rect -955 1765 -950 2085
rect -1100 1735 -1065 1740
rect -980 1735 -950 1765
rect -920 2085 -890 2115
rect -920 1765 -915 2085
rect -895 1765 -890 2085
rect -920 1755 -890 1765
rect -860 2085 -830 2095
rect -860 1765 -855 2085
rect -835 1765 -830 2085
rect -860 1735 -830 1765
rect -800 2085 -770 2115
rect -800 1765 -795 2085
rect -775 1765 -770 2085
rect -800 1755 -770 1765
rect -740 2085 -710 2095
rect -740 1765 -735 2085
rect -715 1765 -710 2085
rect -740 1735 -710 1765
rect -680 2085 -650 2115
rect -680 1765 -675 2085
rect -655 1765 -650 2085
rect -680 1755 -650 1765
rect -620 2085 -590 2095
rect -620 1765 -615 2085
rect -595 1765 -590 2085
rect -620 1735 -590 1765
rect -560 2085 -530 2115
rect -440 2095 -410 2115
rect -35 2095 -5 2115
rect -560 1765 -555 2085
rect -535 1765 -530 2085
rect -560 1755 -530 1765
rect -500 2085 -470 2095
rect -500 1765 -495 2085
rect -475 1765 -470 2085
rect -500 1735 -470 1765
rect -440 2085 -370 2095
rect -440 1765 -435 2085
rect -415 1765 -395 2085
rect -375 1765 -370 2085
rect -440 1755 -370 1765
rect -75 2085 -5 2095
rect -75 1765 -70 2085
rect -50 1765 -30 2085
rect -10 1765 -5 2085
rect -75 1755 -5 1765
rect 25 2085 55 2095
rect 25 1765 30 2085
rect 50 1765 55 2085
rect 25 1740 55 1765
rect 85 2085 115 2115
rect 85 1765 90 2085
rect 110 1765 115 2085
rect 85 1755 115 1765
rect 145 2085 175 2095
rect 145 1765 150 2085
rect 170 1765 175 2085
rect 25 1735 60 1740
rect 145 1735 175 1765
rect 205 2085 235 2115
rect 205 1765 210 2085
rect 230 1765 235 2085
rect 205 1755 235 1765
rect 265 2085 295 2095
rect 265 1765 270 2085
rect 290 1765 295 2085
rect 265 1735 295 1765
rect 325 2085 355 2115
rect 325 1765 330 2085
rect 350 1765 355 2085
rect 325 1755 355 1765
rect 385 2085 415 2095
rect 385 1765 390 2085
rect 410 1765 415 2085
rect 385 1735 415 1765
rect 445 2085 475 2115
rect 445 1765 450 2085
rect 470 1765 475 2085
rect 445 1755 475 1765
rect 505 2085 535 2095
rect 505 1765 510 2085
rect 530 1765 535 2085
rect 505 1735 535 1765
rect 565 2085 595 2115
rect 685 2095 715 2115
rect 975 2095 1005 2115
rect 565 1765 570 2085
rect 590 1765 595 2085
rect 565 1755 595 1765
rect 625 2085 655 2095
rect 625 1765 630 2085
rect 650 1765 655 2085
rect 625 1735 655 1765
rect 685 2085 755 2095
rect 685 1765 690 2085
rect 710 1765 730 2085
rect 750 1765 755 2085
rect 685 1755 755 1765
rect 935 2085 1005 2095
rect 935 1765 940 2085
rect 960 1765 980 2085
rect 1000 1765 1005 2085
rect 935 1755 1005 1765
rect 1035 2085 1065 2095
rect 1035 1765 1040 2085
rect 1060 1765 1065 2085
rect -1100 1725 -465 1735
rect -1100 1715 -495 1725
rect -505 1705 -495 1715
rect -475 1705 -465 1725
rect 25 1725 655 1735
rect 25 1715 330 1725
rect -505 1695 -465 1705
rect 325 1705 330 1715
rect 350 1715 655 1725
rect 1035 1735 1065 1765
rect 1095 2085 1125 2115
rect 1095 1765 1100 2085
rect 1120 1765 1125 2085
rect 1095 1755 1125 1765
rect 1155 2085 1185 2095
rect 1155 1765 1160 2085
rect 1180 1765 1185 2085
rect 1155 1735 1185 1765
rect 1215 2085 1245 2115
rect 1215 1765 1220 2085
rect 1240 1765 1245 2085
rect 1215 1755 1245 1765
rect 1275 2085 1305 2095
rect 1275 1765 1280 2085
rect 1300 1765 1305 2085
rect 1275 1735 1305 1765
rect 1335 2085 1365 2115
rect 1335 1765 1340 2085
rect 1360 1765 1365 2085
rect 1335 1755 1365 1765
rect 1395 2085 1425 2095
rect 1395 1765 1400 2085
rect 1420 1765 1425 2085
rect 1395 1735 1425 1765
rect 1455 2085 1485 2115
rect 1455 1765 1460 2085
rect 1480 1765 1485 2085
rect 1455 1755 1485 1765
rect 1515 2085 1545 2095
rect 1515 1765 1520 2085
rect 1540 1765 1545 2085
rect 1515 1735 1545 1765
rect 1575 2085 1605 2115
rect 1695 2095 1725 2115
rect 2100 2095 2130 2115
rect 1575 1765 1580 2085
rect 1600 1765 1605 2085
rect 1575 1755 1605 1765
rect 1635 2085 1665 2095
rect 1635 1765 1640 2085
rect 1660 1765 1665 2085
rect 1635 1740 1665 1765
rect 1695 2085 1765 2095
rect 1695 1765 1700 2085
rect 1720 1765 1740 2085
rect 1760 1765 1765 2085
rect 1695 1755 1765 1765
rect 2060 2085 2130 2095
rect 2060 1765 2065 2085
rect 2085 1765 2105 2085
rect 2125 1765 2130 2085
rect 2060 1755 2130 1765
rect 2160 2085 2190 2095
rect 2160 1765 2165 2085
rect 2185 1765 2190 2085
rect 1630 1735 1665 1740
rect 2160 1735 2190 1765
rect 2220 2085 2250 2115
rect 2220 1765 2225 2085
rect 2245 1765 2250 2085
rect 2220 1755 2250 1765
rect 2280 2085 2310 2095
rect 2280 1765 2285 2085
rect 2305 1765 2310 2085
rect 2280 1735 2310 1765
rect 2340 2085 2370 2115
rect 2340 1765 2345 2085
rect 2365 1765 2370 2085
rect 2340 1755 2370 1765
rect 2400 2085 2430 2095
rect 2400 1765 2405 2085
rect 2425 1765 2430 2085
rect 2400 1735 2430 1765
rect 2460 2085 2490 2115
rect 2460 1765 2465 2085
rect 2485 1765 2490 2085
rect 2460 1755 2490 1765
rect 2520 2085 2550 2095
rect 2520 1765 2525 2085
rect 2545 1765 2550 2085
rect 2520 1735 2550 1765
rect 2580 2085 2610 2115
rect 2580 1765 2585 2085
rect 2605 1765 2610 2085
rect 2580 1755 2610 1765
rect 2640 2085 2670 2095
rect 2640 1765 2645 2085
rect 2665 1765 2670 2085
rect 2640 1735 2670 1765
rect 2700 2085 2730 2115
rect 2820 2095 2850 2115
rect 2700 1765 2705 2085
rect 2725 1765 2730 2085
rect 2700 1755 2730 1765
rect 2760 2085 2790 2095
rect 2760 1765 2765 2085
rect 2785 1765 2790 2085
rect 2760 1740 2790 1765
rect 2820 2085 2890 2095
rect 2820 1765 2825 2085
rect 2845 1765 2865 2085
rect 2885 1765 2890 2085
rect 2820 1755 2890 1765
rect 2755 1735 2790 1740
rect 1035 1725 1665 1735
rect 1035 1715 1340 1725
rect 350 1705 355 1715
rect 325 1695 355 1705
rect 1335 1705 1340 1715
rect 1360 1715 1665 1725
rect 2155 1725 2790 1735
rect 1360 1705 1365 1715
rect 1335 1695 1365 1705
rect 2155 1705 2165 1725
rect 2185 1715 2790 1725
rect 2185 1705 2195 1715
rect 2155 1695 2195 1705
rect 410 1665 450 1675
rect 410 1645 420 1665
rect 440 1645 450 1665
rect 410 1635 450 1645
rect 1240 1665 1280 1675
rect 1240 1645 1250 1665
rect 1270 1645 1280 1665
rect 1240 1635 1280 1645
rect -715 1620 -675 1630
rect -715 1600 -705 1620
rect -685 1600 -675 1620
rect -715 1590 -675 1600
rect 2365 1620 2405 1630
rect 2365 1600 2375 1620
rect 2395 1600 2405 1620
rect 2365 1590 2405 1600
rect 455 1570 1235 1580
rect 455 1550 465 1570
rect 485 1560 795 1570
rect 485 1550 495 1560
rect 455 1540 495 1550
rect -1135 1480 -1095 1490
rect -1135 1460 -1125 1480
rect -1105 1470 -1095 1480
rect -475 1480 -435 1490
rect 465 1480 485 1540
rect 565 1530 605 1540
rect 565 1510 575 1530
rect 595 1510 605 1530
rect 565 1500 605 1510
rect 575 1480 595 1500
rect 630 1480 650 1560
rect 785 1550 795 1560
rect 815 1560 875 1570
rect 815 1550 825 1560
rect 785 1540 825 1550
rect 865 1550 875 1560
rect 895 1560 1205 1570
rect 895 1550 905 1560
rect 865 1540 905 1550
rect 675 1530 715 1540
rect 675 1510 685 1530
rect 705 1510 715 1530
rect 675 1500 715 1510
rect 685 1480 705 1500
rect 795 1480 815 1540
rect 875 1480 895 1540
rect 975 1530 1015 1540
rect 975 1510 985 1530
rect 1005 1510 1015 1530
rect 975 1500 1015 1510
rect 985 1480 1005 1500
rect 1040 1480 1060 1560
rect 1195 1550 1205 1560
rect 1225 1550 1235 1570
rect 1195 1540 1235 1550
rect 1085 1530 1125 1540
rect 1085 1510 1095 1530
rect 1115 1510 1125 1530
rect 1085 1500 1125 1510
rect 1095 1480 1115 1500
rect 1205 1480 1225 1540
rect 2125 1480 2165 1490
rect -475 1470 -465 1480
rect -1105 1460 -465 1470
rect -445 1460 -435 1480
rect -1135 1450 -435 1460
rect 420 1470 490 1480
rect -1130 1430 -1100 1450
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -1170 1420 -1100 1430
rect -1170 850 -1165 1420
rect -1145 850 -1125 1420
rect -1105 850 -1100 1420
rect -1170 840 -1100 850
rect -1075 1420 -1045 1430
rect -1075 850 -1070 1420
rect -1050 850 -1045 1420
rect -1501 815 -1360 825
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1075 820 -1045 850
rect -1020 1420 -990 1450
rect -1020 850 -1015 1420
rect -995 850 -990 1420
rect -1020 840 -990 850
rect -965 1420 -935 1430
rect -965 850 -960 1420
rect -940 850 -935 1420
rect -965 820 -935 850
rect -910 1420 -880 1450
rect -910 850 -905 1420
rect -885 850 -880 1420
rect -910 840 -880 850
rect -855 1420 -825 1430
rect -855 850 -850 1420
rect -830 850 -825 1420
rect -855 820 -825 850
rect -800 1420 -770 1450
rect -800 850 -795 1420
rect -775 850 -770 1420
rect -800 840 -770 850
rect -745 1420 -715 1430
rect -745 850 -740 1420
rect -720 850 -715 1420
rect -745 820 -715 850
rect -690 1420 -660 1450
rect -690 850 -685 1420
rect -665 850 -660 1420
rect -690 840 -660 850
rect -635 1420 -605 1430
rect -635 850 -630 1420
rect -610 850 -605 1420
rect -635 820 -605 850
rect -580 1420 -550 1450
rect -470 1430 -440 1450
rect -580 850 -575 1420
rect -555 850 -550 1420
rect -580 840 -550 850
rect -525 1420 -495 1430
rect -525 850 -520 1420
rect -500 850 -495 1420
rect -525 820 -495 850
rect -470 1420 -400 1430
rect -470 850 -465 1420
rect -445 850 -425 1420
rect -405 850 -400 1420
rect 420 1250 425 1470
rect 445 1250 465 1470
rect 485 1250 490 1470
rect 420 1240 490 1250
rect 515 1470 545 1480
rect 515 1250 520 1470
rect 540 1250 545 1470
rect 515 1240 545 1250
rect 570 1470 600 1480
rect 570 1250 575 1470
rect 595 1250 600 1470
rect 570 1240 600 1250
rect 625 1470 655 1480
rect 625 1250 630 1470
rect 650 1250 655 1470
rect 625 1240 655 1250
rect 680 1470 710 1480
rect 680 1250 685 1470
rect 705 1250 710 1470
rect 680 1240 710 1250
rect 735 1470 765 1480
rect 735 1250 740 1470
rect 760 1250 765 1470
rect 735 1240 765 1250
rect 790 1470 900 1480
rect 790 1250 795 1470
rect 815 1250 835 1470
rect 855 1250 875 1470
rect 895 1250 900 1470
rect 790 1240 900 1250
rect 925 1470 955 1480
rect 925 1250 930 1470
rect 950 1250 955 1470
rect 925 1240 955 1250
rect 980 1470 1010 1480
rect 980 1250 985 1470
rect 1005 1250 1010 1470
rect 980 1240 1010 1250
rect 1035 1470 1065 1480
rect 1035 1250 1040 1470
rect 1060 1250 1065 1470
rect 1035 1240 1065 1250
rect 1090 1470 1120 1480
rect 1090 1250 1095 1470
rect 1115 1250 1120 1470
rect 1090 1240 1120 1250
rect 1145 1470 1175 1480
rect 1145 1250 1150 1470
rect 1170 1250 1175 1470
rect 1145 1240 1175 1250
rect 1200 1470 1270 1480
rect 1200 1250 1205 1470
rect 1225 1250 1245 1470
rect 1265 1250 1270 1470
rect 2125 1460 2135 1480
rect 2155 1470 2165 1480
rect 2785 1480 2825 1490
rect 2785 1470 2795 1480
rect 2155 1460 2795 1470
rect 2815 1460 2825 1480
rect 2125 1450 2825 1460
rect 2130 1430 2160 1450
rect 1200 1240 1270 1250
rect 2090 1420 2160 1430
rect 515 1230 535 1240
rect 505 1220 535 1230
rect 745 1230 765 1240
rect 925 1230 945 1240
rect 745 1220 775 1230
rect 505 1200 510 1220
rect 530 1200 535 1220
rect 505 1190 535 1200
rect 552 1210 582 1220
rect 552 1190 557 1210
rect 577 1190 582 1210
rect 552 1180 582 1190
rect 620 1210 660 1220
rect 620 1190 630 1210
rect 650 1190 660 1210
rect 620 1180 660 1190
rect 698 1210 728 1220
rect 698 1190 703 1210
rect 723 1190 728 1210
rect 745 1200 750 1220
rect 770 1200 775 1220
rect 745 1190 775 1200
rect 915 1220 945 1230
rect 1155 1230 1175 1240
rect 1155 1220 1185 1230
rect 915 1200 920 1220
rect 940 1200 945 1220
rect 915 1190 945 1200
rect 962 1210 992 1220
rect 962 1190 967 1210
rect 987 1190 992 1210
rect 698 1180 728 1190
rect 962 1180 992 1190
rect 1030 1210 1070 1220
rect 1030 1190 1040 1210
rect 1060 1190 1070 1210
rect 1030 1180 1070 1190
rect 1108 1210 1138 1220
rect 1108 1190 1113 1210
rect 1133 1190 1138 1210
rect 1155 1200 1160 1220
rect 1180 1200 1185 1220
rect 1155 1190 1185 1200
rect 1108 1180 1138 1190
rect 545 1150 585 1160
rect 545 1130 555 1150
rect 575 1130 585 1150
rect 545 1120 585 1130
rect 1105 1150 1145 1160
rect 1105 1130 1115 1150
rect 1135 1130 1145 1150
rect 1105 1120 1145 1130
rect 145 945 175 955
rect 145 925 150 945
rect 170 925 175 945
rect 1515 945 1545 955
rect 145 915 175 925
rect 780 920 835 930
rect 225 895 265 905
rect 225 885 235 895
rect -470 840 -400 850
rect -45 875 235 885
rect 255 885 265 895
rect 780 900 805 920
rect 825 900 835 920
rect 780 890 835 900
rect 880 920 920 930
rect 880 900 890 920
rect 910 900 920 920
rect 1515 925 1520 945
rect 1540 925 1545 945
rect 1515 915 1545 925
rect 880 890 920 900
rect 1425 895 1465 905
rect 255 875 535 885
rect -45 865 535 875
rect 780 870 800 890
rect 890 870 910 890
rect 1425 885 1435 895
rect 1155 875 1435 885
rect 1455 885 1465 895
rect 1455 875 1735 885
rect -1075 810 -495 820
rect -1075 800 -960 810
rect -1501 785 -1360 795
rect -965 790 -960 800
rect -940 800 -495 810
rect -140 835 -70 845
rect -940 790 -935 800
rect -965 780 -935 790
rect -805 710 -765 720
rect -805 690 -795 710
rect -775 690 -765 710
rect -140 715 -135 835
rect -115 715 -95 835
rect -75 715 -70 835
rect -140 705 -70 715
rect -45 835 -15 865
rect -45 715 -40 835
rect -20 715 -15 835
rect -45 705 -15 715
rect 10 835 40 845
rect 10 715 15 835
rect 35 715 40 835
rect -805 680 -765 690
rect -95 685 -75 705
rect 10 685 40 715
rect 65 835 95 865
rect 65 715 70 835
rect 90 715 95 835
rect 65 705 95 715
rect 120 835 150 845
rect 120 715 125 835
rect 145 715 150 835
rect 120 685 150 715
rect 175 835 205 865
rect 175 715 180 835
rect 200 715 205 835
rect 175 705 205 715
rect 230 835 260 845
rect 230 715 235 835
rect 255 715 260 835
rect 230 685 260 715
rect 285 835 315 865
rect 285 715 290 835
rect 310 715 315 835
rect 285 705 315 715
rect 340 835 370 845
rect 340 715 345 835
rect 365 715 370 835
rect 340 685 370 715
rect 395 835 425 865
rect 395 715 400 835
rect 420 715 425 835
rect 395 705 425 715
rect 450 835 480 845
rect 450 715 455 835
rect 475 715 480 835
rect 450 685 480 715
rect 505 835 535 865
rect 680 860 750 870
rect 505 715 510 835
rect 530 715 535 835
rect 505 705 535 715
rect 560 835 630 845
rect 560 715 565 835
rect 585 715 605 835
rect 625 715 630 835
rect 560 705 630 715
rect 565 685 585 705
rect -100 675 -70 685
rect -1145 665 -1105 675
rect -1145 645 -1135 665
rect -1115 645 -1105 665
rect -530 665 -490 675
rect -530 655 -520 665
rect -1145 635 -1105 645
rect -1125 615 -1105 635
rect -1070 645 -520 655
rect -500 645 -490 665
rect -1070 635 -490 645
rect -465 665 -425 675
rect -465 645 -455 665
rect -435 645 -425 665
rect -100 655 -95 675
rect -75 655 -70 675
rect 10 675 480 685
rect 10 665 235 675
rect -100 645 -70 655
rect 230 655 235 665
rect 255 665 480 675
rect 560 675 590 685
rect 255 655 260 665
rect 230 645 260 655
rect 560 655 565 675
rect 585 655 590 675
rect 560 645 590 655
rect -465 635 -425 645
rect 680 640 685 860
rect 705 640 725 860
rect 745 640 750 860
rect -1070 615 -1050 635
rect -960 615 -940 635
rect -850 615 -830 635
rect -740 615 -720 635
rect -630 615 -610 635
rect -520 615 -500 635
rect -465 615 -445 635
rect 680 630 750 640
rect 775 860 805 870
rect 775 640 780 860
rect 800 640 805 860
rect 775 630 805 640
rect 830 860 860 870
rect 830 640 835 860
rect 855 640 860 860
rect -1170 605 -1100 615
rect -1490 537 -1275 572
rect -1490 517 -1455 537
rect -1310 517 -1275 537
rect -1395 467 -1370 517
rect -1170 435 -1165 605
rect -1145 435 -1125 605
rect -1105 435 -1100 605
rect -1170 425 -1100 435
rect -1075 605 -1045 615
rect -1075 435 -1070 605
rect -1050 435 -1045 605
rect -1075 425 -1045 435
rect -1020 605 -990 615
rect -1020 435 -1015 605
rect -995 435 -990 605
rect -1020 405 -990 435
rect -965 605 -935 615
rect -965 435 -960 605
rect -940 435 -935 605
rect -965 425 -935 435
rect -910 605 -880 615
rect -910 435 -905 605
rect -885 435 -880 605
rect -910 405 -880 435
rect -855 605 -825 615
rect -855 435 -850 605
rect -830 435 -825 605
rect -855 425 -825 435
rect -800 605 -770 615
rect -800 435 -795 605
rect -775 435 -770 605
rect -800 405 -770 435
rect -745 605 -715 615
rect -745 435 -740 605
rect -720 435 -715 605
rect -745 425 -715 435
rect -690 605 -660 615
rect -690 435 -685 605
rect -665 435 -660 605
rect -690 405 -660 435
rect -635 605 -605 615
rect -635 435 -630 605
rect -610 435 -605 605
rect -635 425 -605 435
rect -580 605 -550 615
rect -580 435 -575 605
rect -555 435 -550 605
rect -580 405 -550 435
rect -525 605 -495 615
rect -525 435 -520 605
rect -500 435 -495 605
rect -525 425 -495 435
rect -470 605 -400 615
rect 720 610 750 630
rect 830 610 860 640
rect 885 860 915 870
rect 885 640 890 860
rect 910 640 915 860
rect 885 630 915 640
rect 940 860 1010 870
rect 940 640 945 860
rect 965 640 985 860
rect 1005 640 1010 860
rect 1155 865 1735 875
rect 1060 835 1130 845
rect 1060 715 1065 835
rect 1085 715 1105 835
rect 1125 715 1130 835
rect 1060 705 1130 715
rect 1155 835 1185 865
rect 1155 715 1160 835
rect 1180 715 1185 835
rect 1155 705 1185 715
rect 1210 835 1240 845
rect 1210 715 1215 835
rect 1235 715 1240 835
rect 1105 685 1125 705
rect 1210 685 1240 715
rect 1265 835 1295 865
rect 1265 715 1270 835
rect 1290 715 1295 835
rect 1265 705 1295 715
rect 1320 835 1350 845
rect 1320 715 1325 835
rect 1345 715 1350 835
rect 1320 685 1350 715
rect 1375 835 1405 865
rect 1375 715 1380 835
rect 1400 715 1405 835
rect 1375 705 1405 715
rect 1430 835 1460 845
rect 1430 715 1435 835
rect 1455 715 1460 835
rect 1430 685 1460 715
rect 1485 835 1515 865
rect 1485 715 1490 835
rect 1510 715 1515 835
rect 1485 705 1515 715
rect 1540 835 1570 845
rect 1540 715 1545 835
rect 1565 715 1570 835
rect 1540 685 1570 715
rect 1595 835 1625 865
rect 1595 715 1600 835
rect 1620 715 1625 835
rect 1595 705 1625 715
rect 1650 835 1680 845
rect 1650 715 1655 835
rect 1675 715 1680 835
rect 1650 685 1680 715
rect 1705 835 1735 865
rect 2090 850 2095 1420
rect 2115 850 2135 1420
rect 2155 850 2160 1420
rect 1705 715 1710 835
rect 1730 715 1735 835
rect 1705 705 1735 715
rect 1760 835 1830 845
rect 2090 840 2160 850
rect 2185 1420 2215 1430
rect 2185 850 2190 1420
rect 2210 850 2215 1420
rect 1760 715 1765 835
rect 1785 715 1805 835
rect 1825 715 1830 835
rect 2185 820 2215 850
rect 2240 1420 2270 1450
rect 2240 850 2245 1420
rect 2265 850 2270 1420
rect 2240 840 2270 850
rect 2295 1420 2325 1430
rect 2295 850 2300 1420
rect 2320 850 2325 1420
rect 2295 820 2325 850
rect 2350 1420 2380 1450
rect 2350 850 2355 1420
rect 2375 850 2380 1420
rect 2350 840 2380 850
rect 2405 1420 2435 1430
rect 2405 850 2410 1420
rect 2430 850 2435 1420
rect 2405 820 2435 850
rect 2460 1420 2490 1450
rect 2460 850 2465 1420
rect 2485 850 2490 1420
rect 2460 840 2490 850
rect 2515 1420 2545 1430
rect 2515 850 2520 1420
rect 2540 850 2545 1420
rect 2515 820 2545 850
rect 2570 1420 2600 1450
rect 2570 850 2575 1420
rect 2595 850 2600 1420
rect 2570 840 2600 850
rect 2625 1420 2655 1430
rect 2625 850 2630 1420
rect 2650 850 2655 1420
rect 2625 820 2655 850
rect 2680 1420 2710 1450
rect 2790 1430 2820 1450
rect 2680 850 2685 1420
rect 2705 850 2710 1420
rect 2680 840 2710 850
rect 2735 1420 2765 1430
rect 2735 850 2740 1420
rect 2760 850 2765 1420
rect 2735 820 2765 850
rect 2790 1420 2860 1430
rect 2790 850 2795 1420
rect 2815 850 2835 1420
rect 2855 850 2860 1420
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2790 840 2860 850
rect 2185 810 2765 820
rect 2185 800 2630 810
rect 2625 790 2630 800
rect 2650 800 2765 810
rect 3050 815 3191 825
rect 2650 790 2655 800
rect 2625 780 2655 790
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 1760 705 1830 715
rect 2455 710 2495 720
rect 1765 685 1785 705
rect 2455 690 2465 710
rect 2485 690 2495 710
rect 1100 675 1130 685
rect 1100 655 1105 675
rect 1125 655 1130 675
rect 1210 675 1680 685
rect 1210 665 1435 675
rect 1100 645 1130 655
rect 1430 655 1435 665
rect 1455 665 1680 675
rect 1760 675 1790 685
rect 2455 680 2495 690
rect 1455 655 1460 665
rect 1430 645 1460 655
rect 1760 655 1765 675
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 2115 665 2155 675
rect 2115 645 2125 665
rect 2145 645 2155 665
rect 940 630 1010 640
rect 2115 635 2155 645
rect 2180 665 2220 675
rect 2180 645 2190 665
rect 2210 655 2220 665
rect 2795 665 2835 675
rect 2210 645 2760 655
rect 2180 635 2760 645
rect 940 610 970 630
rect 2135 615 2155 635
rect 2190 615 2210 635
rect 2300 615 2320 635
rect 2410 615 2430 635
rect 2520 615 2540 635
rect 2630 615 2650 635
rect 2740 615 2760 635
rect 2795 645 2805 665
rect 2825 645 2835 665
rect 2795 635 2835 645
rect 2795 615 2815 635
rect -470 435 -465 605
rect -445 435 -425 605
rect -405 435 -400 605
rect 715 600 975 610
rect 715 580 725 600
rect 745 590 945 600
rect 745 580 755 590
rect 715 570 755 580
rect 935 580 945 590
rect 965 580 975 600
rect 935 570 975 580
rect 2090 605 2160 615
rect 145 545 175 555
rect 145 525 150 545
rect 170 525 175 545
rect 145 515 175 525
rect 795 545 825 555
rect 795 525 800 545
rect 820 525 825 545
rect 795 515 825 525
rect 865 545 895 555
rect 865 525 870 545
rect 890 525 895 545
rect 865 515 895 525
rect 1515 545 1545 555
rect 1515 525 1520 545
rect 1540 525 1545 545
rect 1515 515 1545 525
rect 230 500 260 510
rect 230 490 235 500
rect -45 480 235 490
rect 255 490 260 500
rect 715 500 755 510
rect 255 480 535 490
rect -45 470 535 480
rect 715 480 725 500
rect 745 480 755 500
rect 715 470 755 480
rect 935 500 975 510
rect 935 480 945 500
rect 965 480 975 500
rect 1430 500 1460 510
rect 1430 490 1435 500
rect 935 470 975 480
rect 1155 480 1435 490
rect 1455 490 1460 500
rect 1455 480 1735 490
rect 1155 470 1735 480
rect -470 425 -400 435
rect -140 440 -70 450
rect -1025 395 -550 405
rect -1025 375 -1015 395
rect -995 385 -550 395
rect -995 375 -985 385
rect -1025 365 -985 375
rect -750 335 -710 345
rect -750 315 -740 335
rect -720 315 -710 335
rect -750 305 -710 315
rect -140 320 -135 440
rect -115 320 -95 440
rect -75 320 -70 440
rect -140 310 -70 320
rect -45 440 -15 470
rect -45 320 -40 440
rect -20 320 -15 440
rect -45 310 -15 320
rect 10 440 40 450
rect 10 320 15 440
rect 35 320 40 440
rect -95 290 -75 310
rect 10 290 40 320
rect 65 440 95 470
rect 65 320 70 440
rect 90 320 95 440
rect 65 310 95 320
rect 120 440 150 450
rect 120 320 125 440
rect 145 320 150 440
rect 120 290 150 320
rect 175 440 205 470
rect 175 320 180 440
rect 200 320 205 440
rect 175 310 205 320
rect 230 440 260 450
rect 230 320 235 440
rect 255 320 260 440
rect 230 290 260 320
rect 285 440 315 470
rect 285 320 290 440
rect 310 320 315 440
rect 285 310 315 320
rect 340 440 370 450
rect 340 320 345 440
rect 365 320 370 440
rect 340 290 370 320
rect 395 440 425 470
rect 395 320 400 440
rect 420 320 425 440
rect 395 310 425 320
rect 450 440 480 450
rect 450 320 455 440
rect 475 320 480 440
rect 450 290 480 320
rect 505 440 535 470
rect 725 450 745 470
rect 945 450 965 470
rect 505 320 510 440
rect 530 320 535 440
rect 505 310 535 320
rect 560 440 630 450
rect 560 320 565 440
rect 585 320 605 440
rect 625 320 630 440
rect 560 310 630 320
rect 680 440 750 450
rect 680 320 685 440
rect 705 320 725 440
rect 745 320 750 440
rect 680 310 750 320
rect 775 440 805 450
rect 775 320 780 440
rect 800 320 805 440
rect 775 310 805 320
rect 830 440 860 450
rect 830 320 835 440
rect 855 320 860 440
rect 830 310 860 320
rect 885 440 915 450
rect 885 320 890 440
rect 910 320 915 440
rect 885 310 915 320
rect 940 440 1010 450
rect 940 320 945 440
rect 965 320 985 440
rect 1005 320 1010 440
rect 940 310 1010 320
rect 1060 440 1130 450
rect 1060 320 1065 440
rect 1085 320 1105 440
rect 1125 320 1130 440
rect 1060 310 1130 320
rect 1155 440 1185 470
rect 1155 320 1160 440
rect 1180 320 1185 440
rect 1155 310 1185 320
rect 1210 440 1240 450
rect 1210 320 1215 440
rect 1235 320 1240 440
rect 605 290 625 310
rect 780 290 800 310
rect 835 290 855 310
rect 890 290 910 310
rect 1065 290 1085 310
rect 1210 290 1240 320
rect 1265 440 1295 470
rect 1265 320 1270 440
rect 1290 320 1295 440
rect 1265 310 1295 320
rect 1320 440 1350 450
rect 1320 320 1325 440
rect 1345 320 1350 440
rect 1320 290 1350 320
rect 1375 440 1405 470
rect 1375 320 1380 440
rect 1400 320 1405 440
rect 1375 310 1405 320
rect 1430 440 1460 450
rect 1430 320 1435 440
rect 1455 320 1460 440
rect 1430 290 1460 320
rect 1485 440 1515 470
rect 1485 320 1490 440
rect 1510 320 1515 440
rect 1485 310 1515 320
rect 1540 440 1570 450
rect 1540 320 1545 440
rect 1565 320 1570 440
rect 1540 290 1570 320
rect 1595 440 1625 470
rect 1595 320 1600 440
rect 1620 320 1625 440
rect 1595 310 1625 320
rect 1650 440 1680 450
rect 1650 320 1655 440
rect 1675 320 1680 440
rect 1650 290 1680 320
rect 1705 440 1735 470
rect 1705 320 1710 440
rect 1730 320 1735 440
rect 1705 310 1735 320
rect 1760 440 1830 450
rect 1760 320 1765 440
rect 1785 320 1805 440
rect 1825 320 1830 440
rect 2090 435 2095 605
rect 2115 435 2135 605
rect 2155 435 2160 605
rect 2090 425 2160 435
rect 2185 605 2215 615
rect 2185 435 2190 605
rect 2210 435 2215 605
rect 2185 425 2215 435
rect 2240 605 2270 615
rect 2240 435 2245 605
rect 2265 435 2270 605
rect 2240 405 2270 435
rect 2295 605 2325 615
rect 2295 435 2300 605
rect 2320 435 2325 605
rect 2295 425 2325 435
rect 2350 605 2380 615
rect 2350 435 2355 605
rect 2375 435 2380 605
rect 2350 405 2380 435
rect 2405 605 2435 615
rect 2405 435 2410 605
rect 2430 435 2435 605
rect 2405 425 2435 435
rect 2460 605 2490 615
rect 2460 435 2465 605
rect 2485 435 2490 605
rect 2460 405 2490 435
rect 2515 605 2545 615
rect 2515 435 2520 605
rect 2540 435 2545 605
rect 2515 425 2545 435
rect 2570 605 2600 615
rect 2570 435 2575 605
rect 2595 435 2600 605
rect 2570 405 2600 435
rect 2625 605 2655 615
rect 2625 435 2630 605
rect 2650 435 2655 605
rect 2625 425 2655 435
rect 2680 605 2710 615
rect 2680 435 2685 605
rect 2705 435 2710 605
rect 2680 405 2710 435
rect 2735 605 2765 615
rect 2735 435 2740 605
rect 2760 435 2765 605
rect 2735 425 2765 435
rect 2790 605 2860 615
rect 2790 435 2795 605
rect 2815 435 2835 605
rect 2855 435 2860 605
rect 2790 425 2860 435
rect 2965 537 3180 572
rect 2965 517 3000 537
rect 3145 517 3180 537
rect 2240 395 2715 405
rect 2240 385 2685 395
rect 2675 375 2685 385
rect 2705 375 2715 395
rect 2675 365 2715 375
rect 1760 310 1830 320
rect 2400 335 2440 345
rect 2400 315 2410 335
rect 2430 315 2440 335
rect 1765 290 1785 310
rect 2400 305 2440 315
rect 3060 467 3085 517
rect -1025 275 -985 285
rect -1025 255 -1015 275
rect -995 265 -985 275
rect -100 280 -70 290
rect -995 255 -550 265
rect -1025 245 -550 255
rect -100 260 -95 280
rect -75 260 -70 280
rect 10 280 485 290
rect 10 270 455 280
rect -100 250 -70 260
rect 445 260 455 270
rect 475 260 485 280
rect 445 250 485 260
rect 600 280 630 290
rect 600 260 605 280
rect 625 260 630 280
rect 600 250 630 260
rect 775 280 805 290
rect 775 260 780 280
rect 800 260 805 280
rect 775 250 805 260
rect 830 280 860 290
rect 830 260 835 280
rect 855 260 860 280
rect 830 250 860 260
rect 885 280 915 290
rect 885 260 890 280
rect 910 260 915 280
rect 885 250 915 260
rect 1060 280 1090 290
rect 1060 260 1065 280
rect 1085 260 1090 280
rect 1060 250 1090 260
rect 1205 280 1680 290
rect 1205 260 1215 280
rect 1235 270 1680 280
rect 1760 280 1790 290
rect 1235 260 1245 270
rect 1205 250 1245 260
rect 1760 260 1765 280
rect 1785 260 1790 280
rect 2675 275 2715 285
rect 2675 265 2685 275
rect 1760 250 1790 260
rect 2240 255 2685 265
rect 2705 255 2715 275
rect -1170 215 -1100 225
rect -1490 -93 -1455 -85
rect -1490 -113 -1485 -93
rect -1460 -113 -1455 -93
rect -1490 -120 -1455 -113
rect -1430 -93 -1395 -85
rect -1430 -113 -1425 -93
rect -1400 -113 -1395 -93
rect -1430 -120 -1395 -113
rect -1370 -93 -1335 -85
rect -1370 -113 -1365 -93
rect -1340 -113 -1335 -93
rect -1370 -120 -1335 -113
rect -1170 -55 -1165 215
rect -1145 -55 -1125 215
rect -1105 -55 -1100 215
rect -1170 -65 -1100 -55
rect -1130 -85 -1100 -65
rect -1075 215 -1045 225
rect -1075 -55 -1070 215
rect -1050 -55 -1045 215
rect -1075 -85 -1045 -55
rect -1020 215 -990 245
rect -1020 -55 -1015 215
rect -995 -55 -990 215
rect -1020 -65 -990 -55
rect -965 215 -935 225
rect -965 -55 -960 215
rect -940 -55 -935 215
rect -965 -85 -935 -55
rect -910 215 -880 245
rect -910 -55 -905 215
rect -885 -55 -880 215
rect -910 -65 -880 -55
rect -855 215 -825 225
rect -855 -55 -850 215
rect -830 -55 -825 215
rect -855 -85 -825 -55
rect -800 215 -770 245
rect -800 -55 -795 215
rect -775 -55 -770 215
rect -800 -65 -770 -55
rect -745 215 -715 225
rect -745 -55 -740 215
rect -720 -55 -715 215
rect -745 -85 -715 -55
rect -690 215 -660 245
rect -690 -55 -685 215
rect -665 -55 -660 215
rect -690 -65 -660 -55
rect -635 215 -605 225
rect -635 -55 -630 215
rect -610 -55 -605 215
rect -635 -85 -605 -55
rect -580 215 -550 245
rect 2240 245 2715 255
rect -580 -55 -575 215
rect -555 -55 -550 215
rect -580 -65 -550 -55
rect -525 215 -495 225
rect -525 -55 -520 215
rect -500 -55 -495 215
rect -525 -85 -495 -55
rect -470 215 -400 225
rect -470 -55 -465 215
rect -445 -55 -425 215
rect -405 -55 -400 215
rect 2090 215 2160 225
rect 775 5 805 15
rect 775 -15 780 5
rect 800 -15 805 5
rect 775 -25 805 -15
rect 830 10 860 20
rect 830 -10 835 10
rect 855 -10 860 10
rect 830 -20 860 -10
rect 885 5 915 15
rect 885 -15 890 5
rect 910 -15 915 5
rect 885 -25 915 -15
rect 780 -45 800 -25
rect 890 -45 910 -25
rect -470 -65 -400 -55
rect 680 -55 750 -45
rect -470 -85 -440 -65
rect -1310 -93 -1275 -85
rect -1310 -113 -1305 -93
rect -1280 -113 -1275 -93
rect -1310 -120 -1275 -113
rect -1145 -95 -1105 -85
rect -1145 -115 -1135 -95
rect -1115 -115 -1105 -95
rect -1075 -95 -495 -85
rect -1075 -105 -795 -95
rect -1145 -125 -1105 -115
rect -805 -115 -795 -105
rect -775 -105 -495 -95
rect -465 -95 -425 -85
rect -775 -115 -765 -105
rect -805 -125 -765 -115
rect -465 -115 -455 -95
rect -435 -115 -425 -95
rect -465 -125 -425 -115
rect -805 -250 -765 -240
rect -805 -270 -795 -250
rect -775 -270 -765 -250
rect -805 -280 -765 -270
rect 680 -275 685 -55
rect 705 -275 725 -55
rect 745 -275 750 -55
rect 680 -285 750 -275
rect 775 -55 805 -45
rect 775 -275 780 -55
rect 800 -275 805 -55
rect 775 -285 805 -275
rect 830 -55 860 -45
rect 830 -275 835 -55
rect 855 -275 860 -55
rect -1005 -310 -965 -300
rect 720 -305 750 -285
rect 830 -305 860 -275
rect 885 -55 915 -45
rect 885 -275 890 -55
rect 910 -275 915 -55
rect 885 -285 915 -275
rect 940 -55 1010 -45
rect 940 -275 945 -55
rect 965 -275 985 -55
rect 1005 -275 1010 -55
rect 2090 -55 2095 215
rect 2115 -55 2135 215
rect 2155 -55 2160 215
rect 2090 -65 2160 -55
rect 2130 -85 2160 -65
rect 2185 215 2215 225
rect 2185 -55 2190 215
rect 2210 -55 2215 215
rect 2185 -85 2215 -55
rect 2240 215 2270 245
rect 2240 -55 2245 215
rect 2265 -55 2270 215
rect 2240 -65 2270 -55
rect 2295 215 2325 225
rect 2295 -55 2300 215
rect 2320 -55 2325 215
rect 2295 -85 2325 -55
rect 2350 215 2380 245
rect 2350 -55 2355 215
rect 2375 -55 2380 215
rect 2350 -65 2380 -55
rect 2405 215 2435 225
rect 2405 -55 2410 215
rect 2430 -55 2435 215
rect 2405 -85 2435 -55
rect 2460 215 2490 245
rect 2460 -55 2465 215
rect 2485 -55 2490 215
rect 2460 -65 2490 -55
rect 2515 215 2545 225
rect 2515 -55 2520 215
rect 2540 -55 2545 215
rect 2515 -85 2545 -55
rect 2570 215 2600 245
rect 2570 -55 2575 215
rect 2595 -55 2600 215
rect 2570 -65 2600 -55
rect 2625 215 2655 225
rect 2625 -55 2630 215
rect 2650 -55 2655 215
rect 2625 -85 2655 -55
rect 2680 215 2710 245
rect 2680 -55 2685 215
rect 2705 -55 2710 215
rect 2680 -65 2710 -55
rect 2735 215 2765 225
rect 2735 -55 2740 215
rect 2760 -55 2765 215
rect 2735 -85 2765 -55
rect 2790 215 2860 225
rect 2790 -55 2795 215
rect 2815 -55 2835 215
rect 2855 -55 2860 215
rect 2790 -65 2860 -55
rect 2790 -85 2820 -65
rect 2115 -95 2155 -85
rect 2115 -115 2125 -95
rect 2145 -115 2155 -95
rect 2185 -95 2765 -85
rect 2185 -105 2465 -95
rect 2115 -125 2155 -115
rect 2455 -115 2465 -105
rect 2485 -105 2765 -95
rect 2795 -95 2835 -85
rect 2485 -115 2495 -105
rect 2455 -125 2495 -115
rect 2795 -115 2805 -95
rect 2825 -115 2835 -95
rect 2795 -125 2835 -115
rect 2965 -93 3000 -85
rect 2965 -113 2970 -93
rect 2995 -113 3000 -93
rect 2965 -120 3000 -113
rect 3025 -93 3060 -85
rect 3025 -113 3030 -93
rect 3055 -113 3060 -93
rect 3025 -120 3060 -113
rect 3085 -93 3120 -85
rect 3085 -113 3090 -93
rect 3115 -113 3120 -93
rect 3085 -120 3120 -113
rect 3145 -93 3180 -85
rect 3145 -113 3150 -93
rect 3175 -113 3180 -93
rect 3145 -120 3180 -113
rect 940 -285 1010 -275
rect 2455 -250 2495 -240
rect 2455 -270 2465 -250
rect 2485 -270 2495 -250
rect 2455 -280 2495 -270
rect 940 -305 970 -285
rect -1005 -330 -995 -310
rect -975 -320 -965 -310
rect 715 -315 975 -305
rect -975 -330 -570 -320
rect -1005 -340 -570 -330
rect -1140 -370 -1070 -360
rect -1290 -387 -1255 -380
rect -1290 -407 -1285 -387
rect -1260 -407 -1255 -387
rect -1290 -415 -1255 -407
rect -1230 -387 -1195 -380
rect -1230 -407 -1225 -387
rect -1200 -407 -1195 -387
rect -1230 -415 -1195 -407
rect -1255 -1105 -1230 -1055
rect -1140 -1040 -1135 -370
rect -1115 -1040 -1095 -370
rect -1075 -1040 -1070 -370
rect -1140 -1050 -1070 -1040
rect -1000 -370 -970 -340
rect -1000 -1040 -995 -370
rect -975 -1040 -970 -370
rect -1000 -1050 -970 -1040
rect -900 -370 -870 -360
rect -900 -1040 -895 -370
rect -875 -1040 -870 -370
rect -1100 -1070 -1070 -1050
rect -900 -1070 -870 -1040
rect -800 -370 -770 -340
rect -800 -1040 -795 -370
rect -775 -1040 -770 -370
rect -800 -1050 -770 -1040
rect -700 -370 -670 -360
rect -700 -1040 -695 -370
rect -675 -1040 -670 -370
rect -700 -1070 -670 -1040
rect -600 -370 -570 -340
rect 715 -335 725 -315
rect 745 -325 835 -315
rect 745 -335 755 -325
rect 715 -345 755 -335
rect 825 -335 835 -325
rect 855 -325 945 -315
rect 855 -335 865 -325
rect 825 -345 865 -335
rect 935 -335 945 -325
rect 965 -335 975 -315
rect 2655 -310 2695 -300
rect 2655 -320 2665 -310
rect 935 -345 975 -335
rect 2260 -330 2665 -320
rect 2685 -330 2695 -310
rect 2260 -340 2695 -330
rect -600 -1040 -595 -370
rect -575 -1040 -570 -370
rect -600 -1050 -570 -1040
rect -500 -370 -430 -360
rect -500 -1040 -495 -370
rect -475 -1040 -455 -370
rect -435 -1040 -430 -370
rect 2120 -370 2190 -360
rect 1350 -430 1390 -420
rect 445 -440 475 -430
rect 445 -460 450 -440
rect 470 -460 475 -440
rect 1350 -450 1360 -430
rect 1380 -450 1390 -430
rect 1350 -460 1390 -450
rect 445 -470 475 -460
rect 1210 -490 1250 -480
rect 390 -510 1220 -490
rect 1240 -510 1410 -490
rect 240 -550 310 -540
rect 240 -770 245 -550
rect 265 -770 285 -550
rect 305 -770 310 -550
rect 240 -780 310 -770
rect 335 -550 365 -540
rect 335 -770 340 -550
rect 360 -770 365 -550
rect 285 -800 305 -780
rect 335 -800 365 -770
rect 390 -550 420 -510
rect 390 -770 395 -550
rect 415 -770 420 -550
rect 390 -780 420 -770
rect 445 -550 475 -540
rect 445 -770 450 -550
rect 470 -770 475 -550
rect 445 -800 475 -770
rect 500 -550 530 -510
rect 500 -770 505 -550
rect 525 -770 530 -550
rect 500 -780 530 -770
rect 555 -550 585 -540
rect 555 -770 560 -550
rect 580 -770 585 -550
rect 555 -800 585 -770
rect 610 -550 640 -510
rect 610 -770 615 -550
rect 635 -770 640 -550
rect 610 -780 640 -770
rect 665 -550 695 -540
rect 665 -770 670 -550
rect 690 -770 695 -550
rect 665 -800 695 -770
rect 720 -550 750 -510
rect 720 -770 725 -550
rect 745 -770 750 -550
rect 720 -780 750 -770
rect 775 -550 805 -540
rect 775 -770 780 -550
rect 800 -770 805 -550
rect 775 -800 805 -770
rect 830 -550 860 -510
rect 830 -770 835 -550
rect 855 -770 860 -550
rect 830 -780 860 -770
rect 885 -550 915 -540
rect 885 -770 890 -550
rect 910 -770 915 -550
rect 885 -800 915 -770
rect 940 -550 970 -510
rect 940 -770 945 -550
rect 965 -770 970 -550
rect 940 -780 970 -770
rect 995 -550 1025 -540
rect 995 -770 1000 -550
rect 1020 -770 1025 -550
rect 995 -800 1025 -770
rect 1050 -550 1080 -510
rect 1050 -770 1055 -550
rect 1075 -770 1080 -550
rect 1050 -780 1080 -770
rect 1105 -550 1135 -540
rect 1105 -770 1110 -550
rect 1130 -770 1135 -550
rect 1105 -800 1135 -770
rect 1160 -550 1190 -510
rect 1210 -520 1250 -510
rect 1160 -770 1165 -550
rect 1185 -770 1190 -550
rect 1160 -780 1190 -770
rect 1215 -550 1245 -540
rect 1215 -770 1220 -550
rect 1240 -770 1245 -550
rect 1215 -800 1245 -770
rect 1270 -550 1300 -510
rect 1270 -770 1275 -550
rect 1295 -770 1300 -550
rect 1270 -780 1300 -770
rect 1325 -550 1355 -540
rect 1325 -770 1330 -550
rect 1350 -770 1355 -550
rect 1325 -800 1355 -770
rect 1380 -550 1410 -510
rect 1380 -770 1385 -550
rect 1405 -770 1410 -550
rect 1380 -780 1410 -770
rect 1435 -550 1505 -540
rect 1435 -770 1440 -550
rect 1460 -770 1480 -550
rect 1500 -770 1505 -550
rect 1435 -780 1505 -770
rect 1440 -800 1460 -780
rect 265 -810 1470 -800
rect 265 -830 275 -810
rect 295 -820 1440 -810
rect 295 -830 305 -820
rect 265 -840 305 -830
rect 1430 -830 1440 -820
rect 1460 -830 1470 -810
rect 1430 -840 1470 -830
rect 660 -905 700 -895
rect 660 -925 670 -905
rect 690 -925 700 -905
rect 660 -935 700 -925
rect 1130 -905 1170 -895
rect 1130 -925 1140 -905
rect 1160 -925 1170 -905
rect 1130 -935 1170 -925
rect 1305 -910 1345 -900
rect 1305 -930 1315 -910
rect 1335 -930 1345 -910
rect 1305 -940 1345 -930
rect -500 -1050 -430 -1040
rect 460 -965 530 -955
rect -500 -1070 -470 -1050
rect -1105 -1080 -465 -1070
rect -1105 -1100 -1095 -1080
rect -1075 -1090 -795 -1080
rect -1075 -1100 -1065 -1090
rect -1105 -1110 -1065 -1100
rect -805 -1100 -795 -1090
rect -775 -1090 -495 -1080
rect -775 -1100 -765 -1090
rect -805 -1110 -765 -1100
rect -505 -1100 -495 -1090
rect -475 -1100 -465 -1080
rect 460 -1085 465 -965
rect 485 -1085 505 -965
rect 525 -1085 530 -965
rect 460 -1095 530 -1085
rect 555 -965 585 -955
rect 555 -1085 560 -965
rect 580 -1085 585 -965
rect 555 -1095 585 -1085
rect 610 -965 640 -955
rect 610 -1085 615 -965
rect 635 -1085 640 -965
rect 610 -1095 640 -1085
rect 665 -965 695 -955
rect 665 -1085 670 -965
rect 690 -1085 695 -965
rect 665 -1095 695 -1085
rect 720 -965 750 -955
rect 720 -1085 725 -965
rect 745 -1085 750 -965
rect 720 -1095 750 -1085
rect 775 -965 805 -955
rect 775 -1085 780 -965
rect 800 -1085 805 -965
rect 775 -1095 805 -1085
rect 830 -965 900 -955
rect 830 -1085 835 -965
rect 855 -1085 875 -965
rect 895 -1085 900 -965
rect 965 -965 995 -955
rect 965 -1005 970 -965
rect 925 -1015 970 -1005
rect 925 -1035 935 -1015
rect 955 -1035 970 -1015
rect 925 -1045 970 -1035
rect 830 -1095 900 -1085
rect 965 -1085 970 -1045
rect 990 -1085 995 -965
rect 965 -1095 995 -1085
rect 1305 -965 1335 -940
rect 1305 -1085 1310 -965
rect 1330 -1085 1335 -965
rect 2120 -1040 2125 -370
rect 2145 -1040 2165 -370
rect 2185 -1040 2190 -370
rect 2120 -1050 2190 -1040
rect 2260 -370 2290 -340
rect 2260 -1040 2265 -370
rect 2285 -1040 2290 -370
rect 2260 -1050 2290 -1040
rect 2360 -370 2390 -360
rect 2360 -1040 2365 -370
rect 2385 -1040 2390 -370
rect 2160 -1070 2190 -1050
rect 2360 -1070 2390 -1040
rect 2460 -370 2490 -340
rect 2460 -1040 2465 -370
rect 2485 -1040 2490 -370
rect 2460 -1050 2490 -1040
rect 2560 -370 2590 -360
rect 2560 -1040 2565 -370
rect 2585 -1040 2590 -370
rect 2560 -1070 2590 -1040
rect 2660 -370 2690 -340
rect 2660 -1040 2665 -370
rect 2685 -1040 2690 -370
rect 2660 -1050 2690 -1040
rect 2760 -370 2830 -360
rect 2760 -1040 2765 -370
rect 2785 -1040 2805 -370
rect 2825 -1040 2830 -370
rect 2885 -387 2920 -380
rect 2885 -407 2890 -387
rect 2915 -407 2920 -387
rect 2885 -415 2920 -407
rect 2945 -387 2980 -380
rect 2945 -407 2950 -387
rect 2975 -407 2980 -387
rect 2945 -415 2980 -407
rect 2760 -1050 2830 -1040
rect 2760 -1070 2790 -1050
rect 1305 -1095 1335 -1085
rect 2155 -1080 2795 -1070
rect -505 -1110 -465 -1100
rect 500 -1125 530 -1095
rect 500 -1145 505 -1125
rect 525 -1145 530 -1125
rect 500 -1155 530 -1145
rect 830 -1125 860 -1095
rect 2155 -1100 2165 -1080
rect 2185 -1090 2465 -1080
rect 2185 -1100 2195 -1090
rect 2155 -1110 2195 -1100
rect 2455 -1100 2465 -1090
rect 2485 -1090 2765 -1080
rect 2485 -1100 2495 -1090
rect 2455 -1110 2495 -1100
rect 2755 -1100 2765 -1090
rect 2785 -1100 2795 -1080
rect 2755 -1110 2795 -1100
rect 2920 -1105 2945 -1055
rect 830 -1145 835 -1125
rect 855 -1145 860 -1125
rect 830 -1155 860 -1145
<< viali >>
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1040 2700 1060 2720
rect 510 2530 530 2550
rect 570 2530 590 2550
rect 630 2530 650 2550
rect 690 2530 710 2550
rect 1100 2700 1120 2720
rect 1160 2700 1180 2720
rect 1450 2700 1470 2720
rect 85 2280 105 2300
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1526 2280 1546 2300
rect 1585 2280 1605 2300
rect -795 2125 -775 2145
rect -435 2125 -415 2145
rect -30 2125 -10 2145
rect 1700 2125 1720 2145
rect 2105 2125 2125 2145
rect 2465 2125 2485 2145
rect -495 1705 -475 1725
rect 330 1705 350 1725
rect 1340 1705 1360 1725
rect 2165 1705 2185 1725
rect 420 1645 440 1665
rect 1250 1645 1270 1665
rect -705 1600 -685 1620
rect 2375 1600 2395 1620
rect 575 1510 595 1530
rect 685 1510 705 1530
rect 985 1510 1005 1530
rect 1205 1550 1225 1570
rect 1095 1510 1115 1530
rect -465 1460 -445 1480
rect -1495 1400 -1475 1420
rect -1440 1400 -1420 1420
rect -1385 1400 -1365 1420
rect -1495 795 -1475 815
rect -1440 795 -1420 815
rect -1385 795 -1365 815
rect 2135 1460 2155 1480
rect 510 1200 530 1220
rect 557 1190 577 1210
rect 630 1190 650 1210
rect 703 1190 723 1210
rect 750 1200 770 1220
rect 920 1200 940 1220
rect 967 1190 987 1210
rect 1040 1190 1060 1210
rect 1113 1190 1133 1210
rect 1160 1200 1180 1220
rect 555 1130 575 1150
rect 1115 1130 1135 1150
rect 150 925 170 945
rect 235 875 255 895
rect 805 900 825 920
rect 890 900 910 920
rect 1520 925 1540 945
rect 1435 875 1455 895
rect -960 790 -940 810
rect -795 690 -775 710
rect -1135 645 -1115 665
rect -520 645 -500 665
rect -455 645 -435 665
rect -95 655 -75 675
rect 235 655 255 675
rect 565 655 585 675
rect 3055 1400 3075 1420
rect 3110 1400 3130 1420
rect 3165 1400 3185 1420
rect 2630 790 2650 810
rect 3055 795 3075 815
rect 3110 795 3130 815
rect 3165 795 3185 815
rect 2465 690 2485 710
rect 1105 655 1125 675
rect 1435 655 1455 675
rect 1765 655 1785 675
rect 2125 645 2145 665
rect 2190 645 2210 665
rect 2805 645 2825 665
rect 725 580 745 600
rect 945 580 965 600
rect 150 525 170 545
rect 800 525 820 545
rect 870 525 890 545
rect 1520 525 1540 545
rect 235 480 255 500
rect 725 480 745 500
rect 945 480 965 500
rect 1435 480 1455 500
rect -1015 375 -995 395
rect -740 315 -720 335
rect 2685 375 2705 395
rect 2410 315 2430 335
rect -1015 255 -995 275
rect -95 260 -75 280
rect 455 260 475 280
rect 605 260 625 280
rect 780 260 800 280
rect 835 260 855 280
rect 890 260 910 280
rect 1065 260 1085 280
rect 1215 260 1235 280
rect 1765 260 1785 280
rect 2685 255 2705 275
rect -1485 -113 -1460 -93
rect -1425 -113 -1400 -93
rect -1365 -113 -1340 -93
rect 780 -15 800 5
rect 835 -10 855 10
rect 890 -15 910 5
rect -1305 -113 -1280 -93
rect -1135 -115 -1115 -95
rect -795 -115 -775 -95
rect -455 -115 -435 -95
rect -795 -270 -775 -250
rect 2125 -115 2145 -95
rect 2465 -115 2485 -95
rect 2805 -115 2825 -95
rect 2970 -113 2995 -93
rect 3030 -113 3055 -93
rect 3090 -113 3115 -93
rect 3150 -113 3175 -93
rect 2465 -270 2485 -250
rect -995 -330 -975 -310
rect -1285 -407 -1260 -387
rect -1225 -407 -1200 -387
rect 835 -335 855 -315
rect 2665 -330 2685 -310
rect 450 -460 470 -440
rect 1360 -450 1380 -430
rect 1220 -510 1240 -490
rect 275 -830 295 -810
rect 1440 -830 1460 -810
rect 670 -925 690 -905
rect 1140 -925 1160 -905
rect 1315 -930 1335 -910
rect -795 -1100 -775 -1080
rect 560 -1085 580 -965
rect 615 -1085 635 -965
rect 670 -1085 690 -965
rect 725 -1085 745 -965
rect 780 -1085 800 -965
rect 935 -1035 955 -1015
rect 2890 -407 2915 -387
rect 2950 -407 2975 -387
rect 505 -1145 525 -1125
rect 2465 -1100 2485 -1080
rect 835 -1145 855 -1125
<< metal1 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 210 2780 250 2785
rect 210 2750 215 2780
rect 245 2750 250 2780
rect 210 2725 250 2750
rect 620 2780 660 2785
rect 620 2750 625 2780
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 210 2695 215 2725
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 630 2560 650 2745
rect 835 2730 855 4240
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2750 1070 2780
rect 1030 2745 1070 2750
rect 1440 2780 1480 2785
rect 1440 2750 1445 2780
rect 1475 2750 1480 2780
rect 1040 2730 1060 2745
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2695 865 2725
rect 825 2690 865 2695
rect 970 2725 1010 2730
rect 970 2695 975 2725
rect 1005 2695 1010 2725
rect 970 2690 1010 2695
rect 1035 2720 1065 2730
rect 1035 2700 1040 2720
rect 1060 2700 1065 2720
rect 1035 2690 1065 2700
rect 1090 2725 1130 2730
rect 1090 2695 1095 2725
rect 1125 2695 1130 2725
rect 1090 2690 1130 2695
rect 1150 2725 1190 2730
rect 1150 2695 1155 2725
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1440 2725 1480 2750
rect 1440 2695 1445 2725
rect 1475 2695 1480 2725
rect 1440 2690 1480 2695
rect 835 2560 855 2690
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2525 540 2555
rect 500 2520 540 2525
rect 560 2555 600 2560
rect 560 2525 565 2555
rect 595 2525 600 2555
rect 560 2520 600 2525
rect 625 2550 655 2560
rect 625 2530 630 2550
rect 650 2530 655 2550
rect 625 2520 655 2530
rect 680 2555 720 2560
rect 680 2525 685 2555
rect 715 2525 720 2555
rect 680 2520 720 2525
rect 825 2555 865 2560
rect 825 2525 830 2555
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2275 115 2305
rect 75 2270 115 2275
rect 139 2305 169 2310
rect 139 2270 169 2275
rect 609 2305 639 2310
rect 609 2270 639 2275
rect 770 2305 810 2310
rect 770 2275 775 2305
rect 805 2275 810 2305
rect 770 2270 810 2275
rect -805 2205 -765 2210
rect -805 2175 -800 2205
rect -770 2175 -765 2205
rect -805 2170 -765 2175
rect -235 2205 -195 2210
rect -235 2175 -230 2205
rect -200 2175 -195 2205
rect -235 2170 -195 2175
rect -800 2145 -770 2170
rect -800 2125 -795 2145
rect -775 2125 -770 2145
rect -800 2115 -770 2125
rect -445 2150 -405 2155
rect -445 2120 -440 2150
rect -410 2120 -405 2150
rect -445 2115 -405 2120
rect -280 2150 -240 2155
rect -280 2120 -275 2150
rect -245 2120 -240 2150
rect -280 2115 -240 2120
rect -270 1735 -250 2115
rect -505 1730 -465 1735
rect -505 1700 -500 1730
rect -470 1700 -465 1730
rect -505 1695 -465 1700
rect -280 1730 -240 1735
rect -280 1700 -275 1730
rect -245 1700 -240 1730
rect -280 1695 -240 1700
rect -370 1670 -330 1675
rect -370 1640 -365 1670
rect -335 1640 -330 1670
rect -370 1635 -330 1640
rect -715 1625 -675 1630
rect -715 1595 -710 1625
rect -680 1595 -675 1625
rect -715 1590 -675 1595
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -1440 1430 -1420 1505
rect -475 1485 -435 1490
rect -475 1455 -470 1485
rect -440 1455 -435 1485
rect -475 1450 -435 1455
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -360 905 -340 1635
rect -225 1490 -205 2170
rect -40 2150 0 2155
rect -40 2120 -35 2150
rect -5 2120 0 2150
rect -40 2115 0 2120
rect 325 1725 355 1735
rect 325 1705 330 1725
rect 350 1705 355 1725
rect 325 1695 355 1705
rect 330 1675 350 1695
rect 790 1675 810 2270
rect 835 2210 855 2520
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1521 2305 1551 2310
rect 1521 2270 1551 2275
rect 1575 2300 1615 2310
rect 1575 2280 1585 2300
rect 1605 2280 1615 2300
rect 1575 2270 1615 2280
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2230 920 2260
rect 1055 2255 1075 2270
rect 1585 2255 1605 2270
rect 880 2225 920 2230
rect 1045 2250 1085 2255
rect 825 2205 865 2210
rect 825 2175 830 2205
rect 860 2175 865 2205
rect 825 2170 865 2175
rect 320 1670 360 1675
rect 320 1640 325 1670
rect 355 1640 360 1670
rect 320 1635 360 1640
rect 410 1670 450 1675
rect 410 1640 415 1670
rect 445 1640 450 1670
rect 410 1635 450 1640
rect 780 1670 820 1675
rect 780 1640 785 1670
rect 815 1640 820 1670
rect 780 1635 820 1640
rect 880 1630 900 2225
rect 1045 2220 1050 2250
rect 1080 2220 1085 2250
rect 1045 2215 1085 2220
rect 1575 2250 1615 2255
rect 1575 2220 1580 2250
rect 1610 2220 1615 2250
rect 1575 2215 1615 2220
rect 1885 2205 1925 2210
rect 1885 2175 1890 2205
rect 1920 2175 1925 2205
rect 1885 2170 1925 2175
rect 2455 2205 2495 2210
rect 2455 2175 2460 2205
rect 2490 2175 2495 2205
rect 2455 2170 2495 2175
rect 1690 2150 1730 2155
rect 1690 2120 1695 2150
rect 1725 2120 1730 2150
rect 1690 2115 1730 2120
rect 1335 1725 1365 1735
rect 1335 1705 1340 1725
rect 1360 1705 1365 1725
rect 1335 1695 1365 1705
rect 1340 1675 1360 1695
rect 1240 1670 1280 1675
rect 1240 1640 1245 1670
rect 1275 1640 1280 1670
rect 1240 1635 1280 1640
rect 1330 1670 1370 1675
rect 1330 1640 1335 1670
rect 1365 1640 1370 1670
rect 1330 1635 1370 1640
rect 870 1600 875 1630
rect 905 1600 910 1630
rect 1895 1580 1915 2170
rect 1930 2150 1970 2155
rect 1930 2120 1935 2150
rect 1965 2120 1970 2150
rect 1930 2115 1970 2120
rect 2095 2150 2135 2155
rect 2095 2120 2100 2150
rect 2130 2120 2135 2150
rect 2095 2115 2135 2120
rect 2460 2145 2490 2170
rect 2460 2125 2465 2145
rect 2485 2125 2490 2145
rect 2460 2115 2490 2125
rect 1940 1735 1960 2115
rect 1930 1730 1970 1735
rect 1930 1700 1935 1730
rect 1965 1700 1970 1730
rect 1930 1695 1970 1700
rect 2155 1730 2195 1735
rect 2155 1700 2160 1730
rect 2190 1700 2195 1730
rect 2155 1695 2195 1700
rect 2020 1670 2060 1675
rect 2020 1640 2025 1670
rect 2055 1640 2060 1670
rect 2020 1635 2060 1640
rect 1195 1575 1235 1580
rect 1195 1545 1200 1575
rect 1230 1545 1235 1575
rect 1195 1540 1235 1545
rect 1885 1575 1925 1580
rect 1885 1545 1890 1575
rect 1920 1545 1925 1575
rect 1885 1540 1925 1545
rect 565 1535 605 1540
rect 565 1505 570 1535
rect 600 1505 605 1535
rect 565 1500 605 1505
rect 675 1535 715 1540
rect 675 1505 680 1535
rect 710 1505 715 1535
rect 675 1500 715 1505
rect 975 1535 1015 1540
rect 975 1505 980 1535
rect 1010 1505 1015 1535
rect 975 1500 1015 1505
rect 1085 1535 1125 1540
rect 1085 1505 1090 1535
rect 1120 1505 1125 1535
rect 1085 1500 1125 1505
rect 1895 1490 1915 1540
rect -235 1485 -195 1490
rect -235 1455 -230 1485
rect -200 1455 -195 1485
rect -235 1450 -195 1455
rect 1885 1485 1925 1490
rect 1885 1455 1890 1485
rect 1920 1455 1925 1485
rect 1885 1450 1925 1455
rect -325 1105 -285 1110
rect -325 1075 -320 1105
rect -290 1075 -285 1105
rect -325 1070 -285 1075
rect -370 900 -330 905
rect -370 870 -365 900
rect -335 870 -330 900
rect -370 865 -330 870
rect -1501 815 -1360 825
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -965 810 -935 820
rect -965 790 -960 810
rect -940 790 -935 810
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 730 -1500 760
rect -1540 725 -1500 730
rect -1530 360 -1510 725
rect -1440 720 -1420 785
rect -965 780 -935 790
rect -960 760 -940 780
rect -530 760 -490 765
rect -970 730 -965 760
rect -935 730 -930 760
rect -530 730 -525 760
rect -495 730 -490 760
rect -530 725 -490 730
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 685 -1410 715
rect -1450 680 -1410 685
rect -805 715 -765 720
rect -805 685 -800 715
rect -770 685 -765 715
rect -805 680 -765 685
rect -520 675 -500 725
rect -360 720 -340 865
rect -370 715 -330 720
rect -370 685 -365 715
rect -335 685 -330 715
rect -370 680 -330 685
rect -1145 670 -1105 675
rect -1145 640 -1140 670
rect -1110 640 -1105 670
rect -1145 635 -1105 640
rect -530 670 -490 675
rect -530 640 -525 670
rect -495 640 -490 670
rect -530 635 -490 640
rect -465 670 -425 675
rect -465 640 -460 670
rect -430 640 -425 670
rect -465 635 -425 640
rect -1270 400 -1230 405
rect -1270 370 -1265 400
rect -1235 370 -1230 400
rect -1270 365 -1230 370
rect -1025 400 -985 405
rect -1025 370 -1020 400
rect -990 370 -985 400
rect -1025 365 -985 370
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect -1545 310 -1495 320
rect -1530 -300 -1510 310
rect -1490 -120 -1486 -85
rect -1459 -120 -1455 -85
rect -1430 -120 -1426 -85
rect -1399 -120 -1395 -85
rect -1370 -120 -1366 -85
rect -1339 -120 -1335 -85
rect -1310 -120 -1306 -85
rect -1279 -120 -1275 -85
rect -1485 -185 -1460 -120
rect -1370 -145 -1335 -120
rect -1260 -140 -1240 365
rect -360 345 -340 680
rect -750 340 -710 345
rect -750 310 -745 340
rect -715 310 -710 340
rect -750 305 -710 310
rect -370 340 -330 345
rect -370 310 -365 340
rect -335 310 -330 340
rect -370 305 -330 310
rect -1225 280 -1185 285
rect -1225 250 -1220 280
rect -1190 250 -1185 280
rect -1225 245 -1185 250
rect -1025 280 -985 285
rect -1025 250 -1020 280
rect -990 250 -985 280
rect -1025 245 -985 250
rect -1215 -85 -1195 245
rect -1225 -90 -1185 -85
rect -1225 -120 -1220 -90
rect -1190 -120 -1185 -90
rect -1225 -125 -1185 -120
rect -1145 -95 -1105 -85
rect -1145 -115 -1135 -95
rect -1115 -115 -1105 -95
rect -1145 -125 -1105 -115
rect -805 -90 -765 -85
rect -805 -120 -800 -90
rect -770 -120 -765 -90
rect -805 -125 -765 -120
rect -465 -95 -425 -85
rect -465 -115 -455 -95
rect -435 -115 -425 -95
rect -465 -125 -425 -115
rect -1135 -140 -1115 -125
rect -455 -140 -435 -125
rect -1370 -180 -1335 -175
rect -1270 -145 -1230 -140
rect -1270 -175 -1265 -145
rect -1235 -175 -1230 -145
rect -1270 -180 -1230 -175
rect -1145 -145 -1105 -140
rect -1145 -175 -1140 -145
rect -1110 -175 -1105 -145
rect -1145 -180 -1105 -175
rect -465 -145 -425 -140
rect -465 -175 -460 -145
rect -430 -175 -425 -145
rect -465 -180 -425 -175
rect -1490 -190 -1455 -185
rect -315 -190 -295 1070
rect -280 770 -240 775
rect -280 740 -275 770
rect -245 740 -240 770
rect -280 735 -240 740
rect -270 -140 -250 735
rect -225 675 -205 1450
rect 505 1225 535 1230
rect 745 1225 775 1230
rect 505 1190 535 1195
rect 552 1210 582 1220
rect 552 1190 557 1210
rect 577 1190 582 1210
rect 552 1180 582 1190
rect 620 1215 660 1220
rect 620 1185 625 1215
rect 655 1185 660 1215
rect 620 1180 660 1185
rect 698 1210 728 1220
rect 698 1190 703 1210
rect 723 1190 728 1210
rect 745 1190 775 1195
rect 915 1220 945 1230
rect 1155 1220 1185 1230
rect 915 1200 920 1220
rect 940 1200 945 1220
rect 915 1190 945 1200
rect 962 1210 992 1220
rect 962 1190 967 1210
rect 987 1190 992 1210
rect 698 1180 728 1190
rect 555 1160 575 1180
rect 545 1155 585 1160
rect 545 1125 550 1155
rect 580 1125 585 1155
rect 545 1120 585 1125
rect 705 1110 725 1180
rect 690 1105 730 1110
rect 690 1075 695 1105
rect 725 1075 730 1105
rect 690 1070 730 1075
rect 915 1065 935 1190
rect 962 1180 992 1190
rect 1030 1215 1070 1220
rect 1030 1185 1035 1215
rect 1065 1185 1070 1215
rect 1030 1180 1070 1185
rect 1108 1210 1138 1220
rect 1108 1190 1113 1210
rect 1133 1190 1138 1210
rect 1155 1200 1160 1220
rect 1180 1200 1185 1220
rect 1155 1190 1185 1200
rect 1108 1180 1138 1190
rect 965 1110 985 1180
rect 1115 1160 1135 1180
rect 1105 1155 1145 1160
rect 1105 1125 1110 1155
rect 1140 1125 1145 1155
rect 1105 1120 1145 1125
rect 960 1105 1000 1110
rect 960 1075 965 1105
rect 995 1075 1000 1105
rect 960 1070 1000 1075
rect 795 1060 835 1065
rect 795 1030 800 1060
rect 830 1030 835 1060
rect 795 1025 835 1030
rect 905 1060 945 1065
rect 905 1030 910 1060
rect 940 1030 945 1060
rect 905 1025 945 1030
rect 805 1010 825 1025
rect 1165 1015 1185 1190
rect 1155 1010 1195 1015
rect 795 1005 835 1010
rect 795 975 800 1005
rect 830 975 835 1005
rect 795 970 835 975
rect 880 1005 920 1010
rect 880 975 885 1005
rect 915 975 920 1005
rect 1155 980 1160 1010
rect 1190 980 1195 1010
rect 1155 975 1195 980
rect 1840 1010 1880 1015
rect 1840 980 1845 1010
rect 1875 980 1880 1010
rect 1840 975 1880 980
rect 880 970 920 975
rect -190 950 -150 955
rect -190 920 -185 950
rect -155 920 -150 950
rect -190 915 -150 920
rect 145 950 175 955
rect 805 930 825 970
rect 890 930 910 970
rect 1515 950 1545 955
rect 145 915 175 920
rect 795 920 835 930
rect -235 670 -195 675
rect -235 640 -230 670
rect -200 640 -195 670
rect -235 635 -195 640
rect -225 -85 -205 635
rect -235 -90 -195 -85
rect -235 -120 -230 -90
rect -200 -120 -195 -90
rect -235 -125 -195 -120
rect -280 -145 -240 -140
rect -280 -175 -275 -145
rect -245 -175 -240 -145
rect -1490 -225 -1455 -220
rect -325 -220 -320 -190
rect -290 -220 -285 -190
rect -325 -225 -285 -220
rect -1290 -245 -1255 -240
rect -1290 -280 -1255 -275
rect -805 -245 -765 -240
rect -805 -275 -800 -245
rect -770 -275 -765 -245
rect -805 -280 -765 -275
rect -1540 -305 -1500 -300
rect -1540 -335 -1535 -305
rect -1505 -335 -1500 -305
rect -1540 -340 -1500 -335
rect -1285 -380 -1260 -280
rect -1230 -305 -1195 -300
rect -1230 -340 -1195 -335
rect -1005 -305 -965 -300
rect -1005 -335 -1000 -305
rect -970 -335 -965 -305
rect -1005 -340 -965 -335
rect -1225 -380 -1200 -340
rect -1290 -415 -1286 -380
rect -1259 -415 -1255 -380
rect -1230 -415 -1226 -380
rect -1199 -415 -1195 -380
rect -805 -1075 -765 -1070
rect -805 -1105 -800 -1075
rect -770 -1105 -765 -1075
rect -805 -1110 -765 -1105
rect -795 -1170 -775 -1110
rect -270 -1170 -250 -175
rect -235 -245 -195 -240
rect -235 -275 -230 -245
rect -200 -275 -195 -245
rect -235 -280 -195 -275
rect -225 -360 -205 -280
rect -235 -365 -195 -360
rect -235 -395 -230 -365
rect -200 -395 -195 -365
rect -235 -400 -195 -395
rect -180 -895 -160 915
rect 225 900 265 905
rect 225 870 230 900
rect 260 870 265 900
rect 795 900 805 920
rect 825 900 835 920
rect 795 890 835 900
rect 880 920 920 930
rect 880 900 890 920
rect 910 900 920 920
rect 1515 915 1545 920
rect 880 890 920 900
rect 1425 900 1465 905
rect 225 865 265 870
rect 1425 870 1430 900
rect 1460 870 1465 900
rect 1425 865 1465 870
rect -100 675 -70 685
rect -100 655 -95 675
rect -75 655 -70 675
rect -100 645 -70 655
rect 230 675 260 685
rect 230 655 235 675
rect 255 655 260 675
rect -95 630 -75 645
rect -105 625 -65 630
rect -105 595 -100 625
rect -70 595 -65 625
rect -105 590 -65 595
rect 145 550 175 555
rect 145 515 175 520
rect 230 500 260 655
rect 560 675 590 685
rect 560 655 565 675
rect 585 655 590 675
rect 560 645 590 655
rect 1100 675 1130 685
rect 1100 655 1105 675
rect 1125 655 1130 675
rect 1100 645 1130 655
rect 1430 675 1460 685
rect 1430 655 1435 675
rect 1455 655 1460 675
rect 565 630 585 645
rect 1105 630 1125 645
rect 555 625 595 630
rect 555 595 560 625
rect 590 595 595 625
rect 1095 625 1135 630
rect 555 590 595 595
rect 715 605 755 610
rect 715 575 720 605
rect 750 575 755 605
rect 715 570 755 575
rect 935 605 975 610
rect 935 575 940 605
rect 970 575 975 605
rect 1095 595 1100 625
rect 1130 595 1135 625
rect 1095 590 1135 595
rect 935 570 975 575
rect 725 510 745 570
rect 795 550 825 555
rect 795 515 825 520
rect 865 550 895 555
rect 865 515 895 520
rect 945 510 965 570
rect 230 480 235 500
rect 255 480 260 500
rect 230 470 260 480
rect 715 500 755 510
rect 715 480 725 500
rect 745 480 755 500
rect 715 470 755 480
rect 935 500 975 510
rect 935 480 945 500
rect 965 480 975 500
rect 935 470 975 480
rect 1430 500 1460 655
rect 1760 675 1790 685
rect 1760 655 1765 675
rect 1785 655 1790 675
rect 1760 645 1790 655
rect 1765 630 1785 645
rect 1755 625 1795 630
rect 1755 595 1760 625
rect 1790 595 1795 625
rect 1755 590 1795 595
rect 1515 550 1545 555
rect 1515 515 1545 520
rect 1430 480 1435 500
rect 1455 480 1460 500
rect 1430 470 1460 480
rect -100 280 -70 290
rect -100 260 -95 280
rect -75 260 -70 280
rect -100 250 -70 260
rect 445 285 485 290
rect 445 255 450 285
rect 480 255 485 285
rect 445 250 485 255
rect 600 280 630 290
rect 600 260 605 280
rect 625 260 630 280
rect 600 250 630 260
rect 775 280 805 290
rect 775 260 780 280
rect 800 260 805 280
rect 775 250 805 260
rect 830 280 860 290
rect 830 260 835 280
rect 855 260 860 280
rect 830 250 860 260
rect 885 280 915 290
rect 885 260 890 280
rect 910 260 915 280
rect 885 250 915 260
rect 1060 280 1090 290
rect 1060 260 1065 280
rect 1085 260 1090 280
rect 1060 250 1090 260
rect 1205 285 1245 290
rect 1205 255 1210 285
rect 1240 255 1245 285
rect 1205 250 1245 255
rect 1760 280 1790 290
rect 1760 260 1765 280
rect 1785 260 1790 280
rect 1760 250 1790 260
rect -95 -305 -75 250
rect 440 15 480 20
rect 440 -15 445 15
rect 475 -15 480 15
rect 440 -20 480 -15
rect -105 -310 -65 -305
rect -105 -340 -100 -310
rect -70 -340 -65 -310
rect -105 -345 -65 -340
rect 450 -430 470 -20
rect 605 -305 625 250
rect 780 235 800 250
rect 780 230 820 235
rect 780 200 785 230
rect 815 200 820 230
rect 780 195 820 200
rect 795 125 815 195
rect 835 180 855 250
rect 890 235 910 250
rect 870 230 910 235
rect 870 200 875 230
rect 905 200 910 230
rect 870 195 910 200
rect 835 175 895 180
rect 835 145 860 175
rect 890 145 895 175
rect 835 140 895 145
rect 795 120 855 125
rect 795 90 800 120
rect 830 90 855 120
rect 795 85 855 90
rect 780 65 820 70
rect 780 35 785 65
rect 815 35 820 65
rect 780 30 820 35
rect 780 15 800 30
rect 835 20 855 85
rect 875 70 895 140
rect 870 65 910 70
rect 870 35 875 65
rect 905 35 910 65
rect 870 30 910 35
rect 830 15 860 20
rect 890 15 910 30
rect 775 5 805 15
rect 775 -15 780 5
rect 800 -15 805 5
rect 775 -25 805 -15
rect 830 -20 860 -15
rect 885 5 915 15
rect 885 -15 890 5
rect 910 -15 915 5
rect 885 -25 915 -15
rect 1065 -305 1085 250
rect 595 -310 635 -305
rect 595 -340 600 -310
rect 630 -340 635 -310
rect 595 -345 635 -340
rect 825 -310 865 -305
rect 825 -340 830 -310
rect 860 -340 865 -310
rect 825 -345 865 -340
rect 1065 -310 1105 -305
rect 1065 -340 1070 -310
rect 1100 -340 1105 -310
rect 1065 -345 1105 -340
rect 445 -440 475 -430
rect 445 -460 450 -440
rect 470 -460 475 -440
rect 445 -470 475 -460
rect 1215 -480 1235 250
rect 1760 -305 1780 250
rect 1750 -310 1790 -305
rect 1750 -340 1755 -310
rect 1785 -340 1790 -310
rect 1750 -345 1790 -340
rect 1850 -420 1870 975
rect 1895 675 1915 1450
rect 1975 1105 2015 1110
rect 1975 1075 1980 1105
rect 2010 1075 2015 1105
rect 1975 1070 2015 1075
rect 1930 760 1970 765
rect 1930 730 1935 760
rect 1965 730 1970 760
rect 1930 725 1970 730
rect 1885 670 1925 675
rect 1885 640 1890 670
rect 1920 640 1925 670
rect 1885 635 1925 640
rect 1895 -85 1915 635
rect 1940 620 1960 725
rect 1930 615 1970 620
rect 1930 585 1935 615
rect 1965 585 1970 615
rect 1930 580 1970 585
rect 1885 -90 1925 -85
rect 1885 -120 1890 -90
rect 1920 -120 1925 -90
rect 1885 -125 1925 -120
rect 1940 -140 1960 580
rect 1930 -145 1970 -140
rect 1930 -175 1935 -145
rect 1965 -175 1970 -145
rect 1885 -245 1925 -240
rect 1885 -275 1890 -245
rect 1920 -275 1925 -245
rect 1885 -280 1925 -275
rect 1895 -360 1915 -280
rect 1940 -305 1960 -175
rect 1985 -190 2005 1070
rect 2030 905 2050 1635
rect 2365 1625 2405 1630
rect 2365 1595 2370 1625
rect 2400 1595 2405 1625
rect 2365 1590 2405 1595
rect 3100 1490 3140 1495
rect 2125 1485 2165 1490
rect 2125 1455 2130 1485
rect 2160 1455 2165 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2125 1450 2165 1455
rect 3110 1430 3130 1455
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2020 900 2060 905
rect 2020 870 2025 900
rect 2055 870 2060 900
rect 2020 865 2060 870
rect 2030 720 2050 865
rect 2625 810 2655 820
rect 2625 790 2630 810
rect 2650 790 2655 810
rect 2625 780 2655 790
rect 3050 815 3191 825
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 2180 760 2220 765
rect 2630 760 2650 780
rect 2180 730 2185 760
rect 2215 730 2220 760
rect 2620 730 2625 760
rect 2655 730 2660 760
rect 2180 725 2220 730
rect 2020 715 2060 720
rect 2020 685 2025 715
rect 2055 685 2060 715
rect 2020 680 2060 685
rect 2030 345 2050 680
rect 2190 675 2210 725
rect 3110 720 3130 785
rect 3190 760 3230 765
rect 3190 730 3195 760
rect 3225 730 3230 760
rect 3190 725 3230 730
rect 2455 715 2495 720
rect 2455 685 2460 715
rect 2490 685 2495 715
rect 2455 680 2495 685
rect 3100 715 3140 720
rect 3100 685 3105 715
rect 3135 685 3140 715
rect 3100 680 3140 685
rect 2115 670 2155 675
rect 2115 640 2120 670
rect 2150 640 2155 670
rect 2115 635 2155 640
rect 2180 670 2220 675
rect 2180 640 2185 670
rect 2215 640 2220 670
rect 2180 635 2220 640
rect 2795 670 2835 675
rect 2795 640 2800 670
rect 2830 640 2835 670
rect 2795 635 2835 640
rect 2675 400 2715 405
rect 2675 370 2680 400
rect 2710 370 2715 400
rect 2675 365 2715 370
rect 2920 400 2960 405
rect 2920 370 2925 400
rect 2955 370 2960 400
rect 2920 365 2960 370
rect 2020 340 2060 345
rect 2020 310 2025 340
rect 2055 310 2060 340
rect 2020 305 2060 310
rect 2400 340 2440 345
rect 2400 310 2405 340
rect 2435 310 2440 340
rect 2400 305 2440 310
rect 2675 280 2715 285
rect 2675 250 2680 280
rect 2710 250 2715 280
rect 2675 245 2715 250
rect 2875 280 2915 285
rect 2875 250 2880 280
rect 2910 250 2915 280
rect 2875 245 2915 250
rect 2885 -85 2905 245
rect 2115 -95 2155 -85
rect 2115 -115 2125 -95
rect 2145 -115 2155 -95
rect 2115 -125 2155 -115
rect 2455 -90 2495 -85
rect 2455 -120 2460 -90
rect 2490 -120 2495 -90
rect 2455 -125 2495 -120
rect 2795 -95 2835 -85
rect 2795 -115 2805 -95
rect 2825 -115 2835 -95
rect 2795 -125 2835 -115
rect 2875 -90 2915 -85
rect 2875 -120 2880 -90
rect 2910 -120 2915 -90
rect 2875 -125 2915 -120
rect 2125 -140 2145 -125
rect 2805 -140 2825 -125
rect 2930 -140 2950 365
rect 3200 360 3220 725
rect 3185 350 3235 360
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2965 -120 2969 -85
rect 2996 -120 3000 -85
rect 3025 -120 3029 -85
rect 3056 -120 3060 -85
rect 3085 -120 3089 -85
rect 3116 -120 3120 -85
rect 3145 -120 3149 -85
rect 3176 -120 3180 -85
rect 2115 -145 2155 -140
rect 2115 -175 2120 -145
rect 2150 -175 2155 -145
rect 2115 -180 2155 -175
rect 2795 -145 2835 -140
rect 2795 -175 2800 -145
rect 2830 -175 2835 -145
rect 2795 -180 2835 -175
rect 2920 -145 2960 -140
rect 2920 -175 2925 -145
rect 2955 -175 2960 -145
rect 2920 -180 2960 -175
rect 3025 -145 3060 -120
rect 3025 -180 3060 -175
rect 3150 -185 3175 -120
rect 3145 -190 3180 -185
rect 1975 -220 1980 -190
rect 2010 -220 2015 -190
rect 1975 -225 2015 -220
rect 3145 -225 3180 -220
rect 2455 -245 2495 -240
rect 2455 -275 2460 -245
rect 2490 -275 2495 -245
rect 2455 -280 2495 -275
rect 2945 -245 2980 -240
rect 2945 -280 2980 -275
rect 2655 -305 2695 -300
rect 1930 -310 1970 -305
rect 1930 -340 1935 -310
rect 1965 -340 1970 -310
rect 2655 -335 2660 -305
rect 2690 -335 2695 -305
rect 2655 -340 2695 -335
rect 2885 -305 2920 -300
rect 2885 -340 2920 -335
rect 1930 -345 1970 -340
rect 1885 -365 1925 -360
rect 1885 -395 1890 -365
rect 1920 -395 1925 -365
rect 1885 -400 1925 -395
rect 1350 -425 1390 -420
rect 1350 -455 1355 -425
rect 1385 -455 1390 -425
rect 1350 -460 1390 -455
rect 1840 -425 1880 -420
rect 1840 -455 1845 -425
rect 1875 -455 1880 -425
rect 1840 -460 1880 -455
rect 1210 -485 1250 -480
rect 1210 -515 1215 -485
rect 1245 -515 1250 -485
rect 1210 -520 1250 -515
rect 1690 -485 1730 -480
rect 1690 -515 1695 -485
rect 1725 -515 1730 -485
rect 1690 -520 1730 -515
rect 265 -805 305 -800
rect 265 -835 270 -805
rect 300 -835 305 -805
rect 265 -840 305 -835
rect 1430 -805 1470 -800
rect 1430 -835 1435 -805
rect 1465 -835 1470 -805
rect 1430 -840 1470 -835
rect -190 -900 -150 -895
rect -190 -930 -185 -900
rect -155 -930 -150 -900
rect -190 -935 -150 -930
rect 550 -900 590 -895
rect 550 -930 555 -900
rect 585 -930 590 -900
rect 550 -935 590 -930
rect 660 -900 700 -895
rect 660 -930 665 -900
rect 695 -930 700 -900
rect 660 -935 700 -930
rect 770 -900 810 -895
rect 770 -930 775 -900
rect 805 -930 810 -900
rect 770 -935 810 -930
rect 1130 -900 1170 -895
rect 1700 -900 1720 -520
rect 1940 -800 1960 -345
rect 2890 -380 2915 -340
rect 2950 -380 2975 -280
rect 3200 -300 3220 310
rect 3190 -305 3230 -300
rect 3190 -335 3195 -305
rect 3225 -335 3230 -305
rect 3190 -340 3230 -335
rect 2885 -415 2889 -380
rect 2916 -415 2920 -380
rect 2945 -415 2949 -380
rect 2976 -415 2980 -380
rect 1930 -805 1970 -800
rect 1930 -835 1935 -805
rect 1965 -835 1970 -805
rect 1930 -840 1970 -835
rect 1130 -930 1135 -900
rect 1165 -930 1170 -900
rect 1130 -935 1170 -930
rect 1305 -905 1345 -900
rect 1305 -935 1310 -905
rect 1340 -935 1345 -905
rect 555 -965 585 -935
rect 555 -1085 560 -965
rect 580 -1085 585 -965
rect 555 -1095 585 -1085
rect 610 -965 640 -955
rect 610 -1085 615 -965
rect 635 -1085 640 -965
rect 610 -1115 640 -1085
rect 665 -965 695 -935
rect 665 -1085 670 -965
rect 690 -1085 695 -965
rect 665 -1095 695 -1085
rect 720 -965 750 -955
rect 720 -1085 725 -965
rect 745 -1085 750 -965
rect 720 -1115 750 -1085
rect 775 -965 805 -935
rect 1305 -940 1345 -935
rect 1690 -905 1730 -900
rect 1690 -935 1695 -905
rect 1725 -935 1730 -905
rect 1690 -940 1730 -935
rect 775 -1085 780 -965
rect 800 -1085 805 -965
rect 925 -1010 965 -1005
rect 925 -1040 930 -1010
rect 960 -1040 965 -1010
rect 925 -1045 965 -1040
rect 775 -1095 805 -1085
rect 935 -1115 955 -1045
rect 500 -1125 530 -1115
rect 500 -1145 505 -1125
rect 525 -1145 530 -1125
rect 500 -1170 530 -1145
rect 605 -1120 645 -1115
rect 605 -1150 610 -1120
rect 640 -1150 645 -1120
rect 605 -1155 645 -1150
rect 715 -1120 755 -1115
rect 715 -1150 720 -1120
rect 750 -1150 755 -1120
rect 715 -1155 755 -1150
rect 830 -1125 860 -1115
rect 830 -1145 835 -1125
rect 855 -1145 860 -1125
rect 830 -1170 860 -1145
rect 925 -1120 965 -1115
rect 925 -1150 930 -1120
rect 960 -1150 965 -1120
rect 925 -1155 965 -1150
rect 1940 -1170 1960 -840
rect 2455 -1075 2495 -1070
rect 2455 -1105 2460 -1075
rect 2490 -1105 2495 -1075
rect 2455 -1110 2495 -1105
rect 2465 -1170 2485 -1110
rect -805 -1175 -765 -1170
rect -805 -1205 -800 -1175
rect -770 -1205 -765 -1175
rect -805 -1210 -765 -1205
rect -280 -1175 -240 -1170
rect -280 -1205 -275 -1175
rect -245 -1205 -240 -1175
rect -280 -1210 -240 -1205
rect 495 -1175 535 -1170
rect 495 -1205 500 -1175
rect 530 -1205 535 -1175
rect 495 -1210 535 -1205
rect 825 -1175 865 -1170
rect 825 -1205 830 -1175
rect 860 -1205 865 -1175
rect 825 -1210 865 -1205
rect 1930 -1175 1970 -1170
rect 1930 -1205 1935 -1175
rect 1965 -1205 1970 -1175
rect 1930 -1210 1970 -1205
rect 2455 -1175 2495 -1170
rect 2455 -1205 2460 -1175
rect 2490 -1205 2495 -1175
rect 2455 -1210 2495 -1205
rect 835 -2420 855 -1210
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via1 >>
rect 830 4245 860 4275
rect 215 2750 245 2780
rect 625 2750 655 2780
rect 215 2720 245 2725
rect 215 2700 220 2720
rect 220 2700 240 2720
rect 240 2700 245 2720
rect 215 2695 245 2700
rect 1035 2750 1065 2780
rect 1445 2750 1475 2780
rect 830 2695 860 2725
rect 975 2720 1005 2725
rect 975 2700 980 2720
rect 980 2700 1000 2720
rect 1000 2700 1005 2720
rect 975 2695 1005 2700
rect 1095 2720 1125 2725
rect 1095 2700 1100 2720
rect 1100 2700 1120 2720
rect 1120 2700 1125 2720
rect 1095 2695 1125 2700
rect 1155 2720 1185 2725
rect 1155 2700 1160 2720
rect 1160 2700 1180 2720
rect 1180 2700 1185 2720
rect 1155 2695 1185 2700
rect 1445 2720 1475 2725
rect 1445 2700 1450 2720
rect 1450 2700 1470 2720
rect 1470 2700 1475 2720
rect 1445 2695 1475 2700
rect 505 2550 535 2555
rect 505 2530 510 2550
rect 510 2530 530 2550
rect 530 2530 535 2550
rect 505 2525 535 2530
rect 565 2550 595 2555
rect 565 2530 570 2550
rect 570 2530 590 2550
rect 590 2530 595 2550
rect 565 2525 595 2530
rect 685 2550 715 2555
rect 685 2530 690 2550
rect 690 2530 710 2550
rect 710 2530 715 2550
rect 685 2525 715 2530
rect 830 2525 860 2555
rect 80 2300 110 2305
rect 80 2280 85 2300
rect 85 2280 105 2300
rect 105 2280 110 2300
rect 80 2275 110 2280
rect 139 2300 169 2305
rect 139 2280 144 2300
rect 144 2280 164 2300
rect 164 2280 169 2300
rect 139 2275 169 2280
rect 609 2300 639 2305
rect 609 2280 614 2300
rect 614 2280 634 2300
rect 634 2280 639 2300
rect 609 2275 639 2280
rect 775 2275 805 2305
rect -800 2175 -770 2205
rect -230 2175 -200 2205
rect -440 2145 -410 2150
rect -440 2125 -435 2145
rect -435 2125 -415 2145
rect -415 2125 -410 2145
rect -440 2120 -410 2125
rect -275 2120 -245 2150
rect -500 1725 -470 1730
rect -500 1705 -495 1725
rect -495 1705 -475 1725
rect -475 1705 -470 1725
rect -500 1700 -470 1705
rect -275 1700 -245 1730
rect -365 1640 -335 1670
rect -710 1620 -680 1625
rect -710 1600 -705 1620
rect -705 1600 -685 1620
rect -685 1600 -680 1620
rect -710 1595 -680 1600
rect -1445 1510 -1415 1540
rect -470 1480 -440 1485
rect -470 1460 -465 1480
rect -465 1460 -445 1480
rect -445 1460 -440 1480
rect -470 1455 -440 1460
rect -35 2145 -5 2150
rect -35 2125 -30 2145
rect -30 2125 -10 2145
rect -10 2125 -5 2145
rect -35 2120 -5 2125
rect 1521 2300 1551 2305
rect 1521 2280 1526 2300
rect 1526 2280 1546 2300
rect 1546 2280 1551 2300
rect 1521 2275 1551 2280
rect 885 2230 915 2260
rect 830 2175 860 2205
rect 325 1640 355 1670
rect 415 1665 445 1670
rect 415 1645 420 1665
rect 420 1645 440 1665
rect 440 1645 445 1665
rect 415 1640 445 1645
rect 785 1640 815 1670
rect 1050 2220 1080 2250
rect 1580 2220 1610 2250
rect 1890 2175 1920 2205
rect 2460 2175 2490 2205
rect 1695 2145 1725 2150
rect 1695 2125 1700 2145
rect 1700 2125 1720 2145
rect 1720 2125 1725 2145
rect 1695 2120 1725 2125
rect 1245 1665 1275 1670
rect 1245 1645 1250 1665
rect 1250 1645 1270 1665
rect 1270 1645 1275 1665
rect 1245 1640 1275 1645
rect 1335 1640 1365 1670
rect 875 1600 905 1630
rect 1935 2120 1965 2150
rect 2100 2145 2130 2150
rect 2100 2125 2105 2145
rect 2105 2125 2125 2145
rect 2125 2125 2130 2145
rect 2100 2120 2130 2125
rect 1935 1700 1965 1730
rect 2160 1725 2190 1730
rect 2160 1705 2165 1725
rect 2165 1705 2185 1725
rect 2185 1705 2190 1725
rect 2160 1700 2190 1705
rect 2025 1640 2055 1670
rect 1200 1570 1230 1575
rect 1200 1550 1205 1570
rect 1205 1550 1225 1570
rect 1225 1550 1230 1570
rect 1200 1545 1230 1550
rect 1890 1545 1920 1575
rect 570 1530 600 1535
rect 570 1510 575 1530
rect 575 1510 595 1530
rect 595 1510 600 1530
rect 570 1505 600 1510
rect 680 1530 710 1535
rect 680 1510 685 1530
rect 685 1510 705 1530
rect 705 1510 710 1530
rect 680 1505 710 1510
rect 980 1530 1010 1535
rect 980 1510 985 1530
rect 985 1510 1005 1530
rect 1005 1510 1010 1530
rect 980 1505 1010 1510
rect 1090 1530 1120 1535
rect 1090 1510 1095 1530
rect 1095 1510 1115 1530
rect 1115 1510 1120 1530
rect 1090 1505 1120 1510
rect -230 1455 -200 1485
rect 1890 1455 1920 1485
rect -320 1075 -290 1105
rect -365 870 -335 900
rect -1535 730 -1505 760
rect -965 730 -935 760
rect -525 730 -495 760
rect -1445 685 -1415 715
rect -800 710 -770 715
rect -800 690 -795 710
rect -795 690 -775 710
rect -775 690 -770 710
rect -800 685 -770 690
rect -365 685 -335 715
rect -1140 665 -1110 670
rect -1140 645 -1135 665
rect -1135 645 -1115 665
rect -1115 645 -1110 665
rect -1140 640 -1110 645
rect -525 665 -495 670
rect -525 645 -520 665
rect -520 645 -500 665
rect -500 645 -495 665
rect -525 640 -495 645
rect -460 665 -430 670
rect -460 645 -455 665
rect -455 645 -435 665
rect -435 645 -430 665
rect -460 640 -430 645
rect -1265 370 -1235 400
rect -1020 395 -990 400
rect -1020 375 -1015 395
rect -1015 375 -995 395
rect -995 375 -990 395
rect -1020 370 -990 375
rect -1535 320 -1505 350
rect -1486 -93 -1459 -85
rect -1486 -113 -1485 -93
rect -1485 -113 -1460 -93
rect -1460 -113 -1459 -93
rect -1486 -120 -1459 -113
rect -1426 -93 -1399 -85
rect -1426 -113 -1425 -93
rect -1425 -113 -1400 -93
rect -1400 -113 -1399 -93
rect -1426 -120 -1399 -113
rect -1366 -93 -1339 -85
rect -1366 -113 -1365 -93
rect -1365 -113 -1340 -93
rect -1340 -113 -1339 -93
rect -1366 -120 -1339 -113
rect -1306 -93 -1279 -85
rect -1306 -113 -1305 -93
rect -1305 -113 -1280 -93
rect -1280 -113 -1279 -93
rect -1306 -120 -1279 -113
rect -745 335 -715 340
rect -745 315 -740 335
rect -740 315 -720 335
rect -720 315 -715 335
rect -745 310 -715 315
rect -365 310 -335 340
rect -1220 250 -1190 280
rect -1020 275 -990 280
rect -1020 255 -1015 275
rect -1015 255 -995 275
rect -995 255 -990 275
rect -1020 250 -990 255
rect -1220 -120 -1190 -90
rect -800 -95 -770 -90
rect -800 -115 -795 -95
rect -795 -115 -775 -95
rect -775 -115 -770 -95
rect -800 -120 -770 -115
rect -1370 -175 -1335 -145
rect -1265 -175 -1235 -145
rect -1140 -175 -1110 -145
rect -460 -175 -430 -145
rect -275 740 -245 770
rect 505 1220 535 1225
rect 745 1220 775 1225
rect 505 1200 510 1220
rect 510 1200 530 1220
rect 530 1200 535 1220
rect 505 1195 535 1200
rect 625 1210 655 1215
rect 625 1190 630 1210
rect 630 1190 650 1210
rect 650 1190 655 1210
rect 625 1185 655 1190
rect 745 1200 750 1220
rect 750 1200 770 1220
rect 770 1200 775 1220
rect 745 1195 775 1200
rect 550 1150 580 1155
rect 550 1130 555 1150
rect 555 1130 575 1150
rect 575 1130 580 1150
rect 550 1125 580 1130
rect 695 1075 725 1105
rect 1035 1210 1065 1215
rect 1035 1190 1040 1210
rect 1040 1190 1060 1210
rect 1060 1190 1065 1210
rect 1035 1185 1065 1190
rect 1110 1150 1140 1155
rect 1110 1130 1115 1150
rect 1115 1130 1135 1150
rect 1135 1130 1140 1150
rect 1110 1125 1140 1130
rect 965 1075 995 1105
rect 800 1030 830 1060
rect 910 1030 940 1060
rect 800 975 830 1005
rect 885 975 915 1005
rect 1160 980 1190 1010
rect 1845 980 1875 1010
rect -185 920 -155 950
rect 145 945 175 950
rect 145 925 150 945
rect 150 925 170 945
rect 170 925 175 945
rect 1515 945 1545 950
rect 145 920 175 925
rect -230 640 -200 670
rect -230 -120 -200 -90
rect -275 -175 -245 -145
rect -1490 -220 -1455 -190
rect -320 -220 -290 -190
rect -1290 -275 -1255 -245
rect -800 -250 -770 -245
rect -800 -270 -795 -250
rect -795 -270 -775 -250
rect -775 -270 -770 -250
rect -800 -275 -770 -270
rect -1535 -335 -1505 -305
rect -1230 -335 -1195 -305
rect -1000 -310 -970 -305
rect -1000 -330 -995 -310
rect -995 -330 -975 -310
rect -975 -330 -970 -310
rect -1000 -335 -970 -330
rect -1286 -387 -1259 -380
rect -1286 -407 -1285 -387
rect -1285 -407 -1260 -387
rect -1260 -407 -1259 -387
rect -1286 -415 -1259 -407
rect -1226 -387 -1199 -380
rect -1226 -407 -1225 -387
rect -1225 -407 -1200 -387
rect -1200 -407 -1199 -387
rect -1226 -415 -1199 -407
rect -800 -1080 -770 -1075
rect -800 -1100 -795 -1080
rect -795 -1100 -775 -1080
rect -775 -1100 -770 -1080
rect -800 -1105 -770 -1100
rect -230 -275 -200 -245
rect -230 -395 -200 -365
rect 230 895 260 900
rect 230 875 235 895
rect 235 875 255 895
rect 255 875 260 895
rect 230 870 260 875
rect 1515 925 1520 945
rect 1520 925 1540 945
rect 1540 925 1545 945
rect 1515 920 1545 925
rect 1430 895 1460 900
rect 1430 875 1435 895
rect 1435 875 1455 895
rect 1455 875 1460 895
rect 1430 870 1460 875
rect -100 595 -70 625
rect 145 545 175 550
rect 145 525 150 545
rect 150 525 170 545
rect 170 525 175 545
rect 145 520 175 525
rect 560 595 590 625
rect 720 600 750 605
rect 720 580 725 600
rect 725 580 745 600
rect 745 580 750 600
rect 720 575 750 580
rect 940 600 970 605
rect 940 580 945 600
rect 945 580 965 600
rect 965 580 970 600
rect 940 575 970 580
rect 1100 595 1130 625
rect 795 545 825 550
rect 795 525 800 545
rect 800 525 820 545
rect 820 525 825 545
rect 795 520 825 525
rect 865 545 895 550
rect 865 525 870 545
rect 870 525 890 545
rect 890 525 895 545
rect 865 520 895 525
rect 1760 595 1790 625
rect 1515 545 1545 550
rect 1515 525 1520 545
rect 1520 525 1540 545
rect 1540 525 1545 545
rect 1515 520 1545 525
rect 450 280 480 285
rect 450 260 455 280
rect 455 260 475 280
rect 475 260 480 280
rect 450 255 480 260
rect 1210 280 1240 285
rect 1210 260 1215 280
rect 1215 260 1235 280
rect 1235 260 1240 280
rect 1210 255 1240 260
rect 445 -15 475 15
rect -100 -340 -70 -310
rect 785 200 815 230
rect 875 200 905 230
rect 860 145 890 175
rect 800 90 830 120
rect 785 35 815 65
rect 875 35 905 65
rect 830 10 860 15
rect 830 -10 835 10
rect 835 -10 855 10
rect 855 -10 860 10
rect 830 -15 860 -10
rect 600 -340 630 -310
rect 830 -315 860 -310
rect 830 -335 835 -315
rect 835 -335 855 -315
rect 855 -335 860 -315
rect 830 -340 860 -335
rect 1070 -340 1100 -310
rect 1755 -340 1785 -310
rect 1980 1075 2010 1105
rect 1935 730 1965 760
rect 1890 640 1920 670
rect 1935 585 1965 615
rect 1890 -120 1920 -90
rect 1935 -175 1965 -145
rect 1890 -275 1920 -245
rect 2370 1620 2400 1625
rect 2370 1600 2375 1620
rect 2375 1600 2395 1620
rect 2395 1600 2400 1620
rect 2370 1595 2400 1600
rect 2130 1480 2160 1485
rect 2130 1460 2135 1480
rect 2135 1460 2155 1480
rect 2155 1460 2160 1480
rect 2130 1455 2160 1460
rect 3105 1460 3135 1490
rect 2025 870 2055 900
rect 2185 730 2215 760
rect 2625 730 2655 760
rect 2025 685 2055 715
rect 3195 730 3225 760
rect 2460 710 2490 715
rect 2460 690 2465 710
rect 2465 690 2485 710
rect 2485 690 2490 710
rect 2460 685 2490 690
rect 3105 685 3135 715
rect 2120 665 2150 670
rect 2120 645 2125 665
rect 2125 645 2145 665
rect 2145 645 2150 665
rect 2120 640 2150 645
rect 2185 665 2215 670
rect 2185 645 2190 665
rect 2190 645 2210 665
rect 2210 645 2215 665
rect 2185 640 2215 645
rect 2800 665 2830 670
rect 2800 645 2805 665
rect 2805 645 2825 665
rect 2825 645 2830 665
rect 2800 640 2830 645
rect 2680 395 2710 400
rect 2680 375 2685 395
rect 2685 375 2705 395
rect 2705 375 2710 395
rect 2680 370 2710 375
rect 2925 370 2955 400
rect 2025 310 2055 340
rect 2405 335 2435 340
rect 2405 315 2410 335
rect 2410 315 2430 335
rect 2430 315 2435 335
rect 2405 310 2435 315
rect 2680 275 2710 280
rect 2680 255 2685 275
rect 2685 255 2705 275
rect 2705 255 2710 275
rect 2680 250 2710 255
rect 2880 250 2910 280
rect 2460 -95 2490 -90
rect 2460 -115 2465 -95
rect 2465 -115 2485 -95
rect 2485 -115 2490 -95
rect 2460 -120 2490 -115
rect 2880 -120 2910 -90
rect 3195 320 3225 350
rect 2969 -93 2996 -85
rect 2969 -113 2970 -93
rect 2970 -113 2995 -93
rect 2995 -113 2996 -93
rect 2969 -120 2996 -113
rect 3029 -93 3056 -85
rect 3029 -113 3030 -93
rect 3030 -113 3055 -93
rect 3055 -113 3056 -93
rect 3029 -120 3056 -113
rect 3089 -93 3116 -85
rect 3089 -113 3090 -93
rect 3090 -113 3115 -93
rect 3115 -113 3116 -93
rect 3089 -120 3116 -113
rect 3149 -93 3176 -85
rect 3149 -113 3150 -93
rect 3150 -113 3175 -93
rect 3175 -113 3176 -93
rect 3149 -120 3176 -113
rect 2120 -175 2150 -145
rect 2800 -175 2830 -145
rect 2925 -175 2955 -145
rect 3025 -175 3060 -145
rect 1980 -220 2010 -190
rect 3145 -220 3180 -190
rect 2460 -250 2490 -245
rect 2460 -270 2465 -250
rect 2465 -270 2485 -250
rect 2485 -270 2490 -250
rect 2460 -275 2490 -270
rect 2945 -275 2980 -245
rect 1935 -340 1965 -310
rect 2660 -310 2690 -305
rect 2660 -330 2665 -310
rect 2665 -330 2685 -310
rect 2685 -330 2690 -310
rect 2660 -335 2690 -330
rect 2885 -335 2920 -305
rect 1890 -395 1920 -365
rect 1355 -430 1385 -425
rect 1355 -450 1360 -430
rect 1360 -450 1380 -430
rect 1380 -450 1385 -430
rect 1355 -455 1385 -450
rect 1845 -455 1875 -425
rect 1215 -490 1245 -485
rect 1215 -510 1220 -490
rect 1220 -510 1240 -490
rect 1240 -510 1245 -490
rect 1215 -515 1245 -510
rect 1695 -515 1725 -485
rect 270 -810 300 -805
rect 270 -830 275 -810
rect 275 -830 295 -810
rect 295 -830 300 -810
rect 270 -835 300 -830
rect 1435 -810 1465 -805
rect 1435 -830 1440 -810
rect 1440 -830 1460 -810
rect 1460 -830 1465 -810
rect 1435 -835 1465 -830
rect -185 -930 -155 -900
rect 555 -930 585 -900
rect 665 -905 695 -900
rect 665 -925 670 -905
rect 670 -925 690 -905
rect 690 -925 695 -905
rect 665 -930 695 -925
rect 775 -930 805 -900
rect 3195 -335 3225 -305
rect 2889 -387 2916 -380
rect 2889 -407 2890 -387
rect 2890 -407 2915 -387
rect 2915 -407 2916 -387
rect 2889 -415 2916 -407
rect 2949 -387 2976 -380
rect 2949 -407 2950 -387
rect 2950 -407 2975 -387
rect 2975 -407 2976 -387
rect 2949 -415 2976 -407
rect 1935 -835 1965 -805
rect 1135 -905 1165 -900
rect 1135 -925 1140 -905
rect 1140 -925 1160 -905
rect 1160 -925 1165 -905
rect 1135 -930 1165 -925
rect 1310 -910 1340 -905
rect 1310 -930 1315 -910
rect 1315 -930 1335 -910
rect 1335 -930 1340 -910
rect 1310 -935 1340 -930
rect 1695 -935 1725 -905
rect 930 -1015 960 -1010
rect 930 -1035 935 -1015
rect 935 -1035 955 -1015
rect 955 -1035 960 -1015
rect 930 -1040 960 -1035
rect 610 -1150 640 -1120
rect 720 -1150 750 -1120
rect 930 -1150 960 -1120
rect 2460 -1080 2490 -1075
rect 2460 -1100 2465 -1080
rect 2465 -1100 2485 -1080
rect 2485 -1100 2490 -1080
rect 2460 -1105 2490 -1100
rect -800 -1205 -770 -1175
rect -275 -1205 -245 -1175
rect 500 -1205 530 -1175
rect 830 -1205 860 -1175
rect 1935 -1205 1965 -1175
rect 2460 -1205 2490 -1175
rect 830 -2455 860 -2425
<< metal2 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 210 2780 250 2785
rect 210 2750 215 2780
rect 245 2775 250 2780
rect 620 2780 660 2785
rect 620 2775 625 2780
rect 245 2755 625 2775
rect 245 2750 250 2755
rect 210 2745 250 2750
rect 620 2750 625 2755
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2775 1070 2780
rect 1440 2780 1480 2785
rect 1440 2775 1445 2780
rect 1065 2755 1445 2775
rect 1065 2750 1070 2755
rect 1030 2745 1070 2750
rect 1440 2750 1445 2755
rect 1475 2750 1480 2780
rect 1440 2745 1480 2750
rect 210 2725 250 2730
rect 210 2695 215 2725
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2720 865 2725
rect 970 2725 1010 2730
rect 970 2720 975 2725
rect 860 2700 975 2720
rect 860 2695 865 2700
rect 825 2690 865 2695
rect 970 2695 975 2700
rect 1005 2720 1010 2725
rect 1090 2725 1130 2730
rect 1090 2720 1095 2725
rect 1005 2700 1095 2720
rect 1005 2695 1010 2700
rect 970 2690 1010 2695
rect 1090 2695 1095 2700
rect 1125 2720 1130 2725
rect 1150 2725 1190 2730
rect 1150 2720 1155 2725
rect 1125 2700 1155 2720
rect 1125 2695 1130 2700
rect 1090 2690 1130 2695
rect 1150 2695 1155 2700
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1440 2725 1480 2730
rect 1440 2695 1445 2725
rect 1475 2695 1480 2725
rect 1440 2690 1480 2695
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2550 540 2555
rect 560 2555 600 2560
rect 560 2550 565 2555
rect 535 2530 565 2550
rect 535 2525 540 2530
rect 500 2520 540 2525
rect 560 2525 565 2530
rect 595 2550 600 2555
rect 680 2555 720 2560
rect 680 2550 685 2555
rect 595 2530 685 2550
rect 595 2525 600 2530
rect 560 2520 600 2525
rect 680 2525 685 2530
rect 715 2550 720 2555
rect 825 2555 865 2560
rect 825 2550 830 2555
rect 715 2530 830 2550
rect 715 2525 720 2530
rect 680 2520 720 2525
rect 825 2525 830 2530
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2300 115 2305
rect 139 2305 169 2310
rect 110 2280 139 2300
rect 110 2275 115 2280
rect 75 2270 115 2275
rect 609 2305 639 2310
rect 169 2280 609 2300
rect 139 2270 169 2275
rect 770 2305 810 2310
rect 770 2300 775 2305
rect 639 2280 775 2300
rect 609 2270 639 2275
rect 770 2275 775 2280
rect 805 2300 810 2305
rect 1521 2305 1551 2310
rect 805 2280 1521 2300
rect 805 2275 810 2280
rect 770 2270 810 2275
rect 1521 2270 1551 2275
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2245 920 2260
rect 1045 2250 1085 2255
rect 1045 2245 1050 2250
rect 915 2230 1050 2245
rect 880 2225 1050 2230
rect 1045 2220 1050 2225
rect 1080 2245 1085 2250
rect 1575 2250 1615 2255
rect 1575 2245 1580 2250
rect 1080 2225 1580 2245
rect 1080 2220 1085 2225
rect 1045 2215 1085 2220
rect 1575 2220 1580 2225
rect 1610 2220 1615 2250
rect 1575 2215 1615 2220
rect -805 2205 -765 2210
rect -805 2175 -800 2205
rect -770 2200 -765 2205
rect -235 2205 -195 2210
rect -235 2200 -230 2205
rect -770 2180 -230 2200
rect -770 2175 -765 2180
rect -805 2170 -765 2175
rect -235 2175 -230 2180
rect -200 2200 -195 2205
rect 825 2205 865 2210
rect 825 2200 830 2205
rect -200 2180 830 2200
rect -200 2175 -195 2180
rect -235 2170 -195 2175
rect 825 2175 830 2180
rect 860 2200 865 2205
rect 1885 2205 1925 2210
rect 1885 2200 1890 2205
rect 860 2180 1890 2200
rect 860 2175 865 2180
rect 825 2170 865 2175
rect 1885 2175 1890 2180
rect 1920 2200 1925 2205
rect 2455 2205 2495 2210
rect 2455 2200 2460 2205
rect 1920 2180 2460 2200
rect 1920 2175 1925 2180
rect 1885 2170 1925 2175
rect 2455 2175 2460 2180
rect 2490 2175 2495 2205
rect 2455 2170 2495 2175
rect -445 2150 -405 2155
rect -445 2120 -440 2150
rect -410 2120 -405 2150
rect -445 2115 -405 2120
rect -280 2150 -240 2155
rect -280 2120 -275 2150
rect -245 2145 -240 2150
rect -40 2150 0 2155
rect -40 2145 -35 2150
rect -245 2125 -35 2145
rect -245 2120 -240 2125
rect -280 2115 -240 2120
rect -40 2120 -35 2125
rect -5 2120 0 2150
rect -40 2115 0 2120
rect 1690 2150 1730 2155
rect 1690 2120 1695 2150
rect 1725 2145 1730 2150
rect 1930 2150 1970 2155
rect 1930 2145 1935 2150
rect 1725 2125 1935 2145
rect 1725 2120 1730 2125
rect 1690 2115 1730 2120
rect 1930 2120 1935 2125
rect 1965 2120 1970 2150
rect 1930 2115 1970 2120
rect 2095 2150 2135 2155
rect 2095 2120 2100 2150
rect 2130 2120 2135 2150
rect 2095 2115 2135 2120
rect -505 1730 -465 1735
rect -505 1700 -500 1730
rect -470 1725 -465 1730
rect -280 1730 -240 1735
rect -280 1725 -275 1730
rect -470 1705 -275 1725
rect -470 1700 -465 1705
rect -505 1695 -465 1700
rect -280 1700 -275 1705
rect -245 1700 -240 1730
rect -280 1695 -240 1700
rect 1930 1730 1970 1735
rect 1930 1700 1935 1730
rect 1965 1725 1970 1730
rect 2155 1730 2195 1735
rect 2155 1725 2160 1730
rect 1965 1705 2160 1725
rect 1965 1700 1970 1705
rect 1930 1695 1970 1700
rect 2155 1700 2160 1705
rect 2190 1700 2195 1730
rect 2155 1695 2195 1700
rect -370 1670 -330 1675
rect -370 1640 -365 1670
rect -335 1665 -330 1670
rect 320 1670 360 1675
rect 320 1665 325 1670
rect -335 1645 325 1665
rect -335 1640 -330 1645
rect -370 1635 -330 1640
rect 320 1640 325 1645
rect 355 1640 360 1670
rect 320 1635 360 1640
rect 410 1670 450 1675
rect 410 1640 415 1670
rect 445 1665 450 1670
rect 780 1670 820 1675
rect 780 1665 785 1670
rect 445 1645 785 1665
rect 445 1640 450 1645
rect 410 1635 450 1640
rect 780 1640 785 1645
rect 815 1665 820 1670
rect 1240 1670 1280 1675
rect 1240 1665 1245 1670
rect 815 1645 1245 1665
rect 815 1640 820 1645
rect 780 1635 820 1640
rect 1240 1640 1245 1645
rect 1275 1640 1280 1670
rect 1240 1635 1280 1640
rect 1330 1670 1370 1675
rect 1330 1640 1335 1670
rect 1365 1665 1370 1670
rect 2020 1670 2060 1675
rect 2020 1665 2025 1670
rect 1365 1645 2025 1665
rect 1365 1640 1370 1645
rect 1330 1635 1370 1640
rect 2020 1640 2025 1645
rect 2055 1640 2060 1670
rect 2020 1635 2060 1640
rect -715 1625 -675 1630
rect -715 1595 -710 1625
rect -680 1620 -675 1625
rect 870 1620 875 1630
rect -680 1600 875 1620
rect 905 1620 910 1630
rect 2365 1625 2405 1630
rect 2365 1620 2370 1625
rect 905 1600 2370 1620
rect -680 1595 -675 1600
rect -715 1590 -675 1595
rect 2365 1595 2370 1600
rect 2400 1595 2405 1625
rect 2365 1590 2405 1595
rect 1195 1575 1235 1580
rect 1195 1545 1200 1575
rect 1230 1570 1235 1575
rect 1885 1575 1925 1580
rect 1885 1570 1890 1575
rect 1230 1550 1890 1570
rect 1230 1545 1235 1550
rect -1450 1540 -1410 1545
rect 1195 1540 1235 1545
rect 1885 1545 1890 1550
rect 1920 1545 1925 1575
rect 1885 1540 1925 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect 565 1535 605 1540
rect 565 1505 570 1535
rect 600 1530 605 1535
rect 675 1535 715 1540
rect 675 1530 680 1535
rect 600 1510 680 1530
rect 600 1505 605 1510
rect 565 1500 605 1505
rect 675 1505 680 1510
rect 710 1505 715 1535
rect 675 1500 715 1505
rect 975 1535 1015 1540
rect 975 1505 980 1535
rect 1010 1530 1015 1535
rect 1085 1535 1125 1540
rect 1085 1530 1090 1535
rect 1010 1510 1090 1530
rect 1010 1505 1015 1510
rect 975 1500 1015 1505
rect 1085 1505 1090 1510
rect 1120 1505 1125 1535
rect 1085 1500 1125 1505
rect 3100 1490 3140 1495
rect -475 1485 -435 1490
rect -475 1455 -470 1485
rect -440 1480 -435 1485
rect -235 1485 -195 1490
rect -235 1480 -230 1485
rect -440 1460 -230 1480
rect -440 1455 -435 1460
rect -475 1450 -435 1455
rect -235 1455 -230 1460
rect -200 1455 -195 1485
rect -235 1450 -195 1455
rect 1885 1485 1925 1490
rect 1885 1455 1890 1485
rect 1920 1480 1925 1485
rect 2125 1485 2165 1490
rect 2125 1480 2130 1485
rect 1920 1460 2130 1480
rect 1920 1455 1925 1460
rect 1885 1450 1925 1455
rect 2125 1455 2130 1460
rect 2160 1455 2165 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2125 1450 2165 1455
rect 505 1225 535 1230
rect 745 1225 775 1230
rect 620 1215 660 1220
rect 620 1210 625 1215
rect 535 1195 625 1210
rect 505 1190 625 1195
rect 620 1185 625 1190
rect 655 1210 660 1215
rect 655 1195 745 1210
rect 1030 1215 1070 1220
rect 1030 1210 1035 1215
rect 775 1195 1035 1210
rect 655 1190 1035 1195
rect 655 1185 660 1190
rect 620 1180 660 1185
rect 1030 1185 1035 1190
rect 1065 1210 1070 1215
rect 1065 1190 1075 1210
rect 1065 1185 1070 1190
rect 1030 1180 1070 1185
rect 545 1155 585 1160
rect 545 1150 550 1155
rect 310 1130 550 1150
rect 545 1125 550 1130
rect 580 1150 585 1155
rect 1105 1155 1145 1160
rect 1105 1150 1110 1155
rect 580 1130 1110 1150
rect 580 1125 585 1130
rect 545 1120 585 1125
rect 1105 1125 1110 1130
rect 1140 1125 1145 1155
rect 1105 1120 1145 1125
rect -325 1105 -285 1110
rect -325 1075 -320 1105
rect -290 1100 -285 1105
rect 690 1105 730 1110
rect 690 1100 695 1105
rect -290 1080 695 1100
rect -290 1075 -285 1080
rect -325 1070 -285 1075
rect 690 1075 695 1080
rect 725 1100 730 1105
rect 960 1105 1000 1110
rect 960 1100 965 1105
rect 725 1080 965 1100
rect 725 1075 730 1080
rect 690 1070 730 1075
rect 960 1075 965 1080
rect 995 1100 1000 1105
rect 1975 1105 2015 1110
rect 1975 1100 1980 1105
rect 995 1080 1980 1100
rect 995 1075 1000 1080
rect 960 1070 1000 1075
rect 1975 1075 1980 1080
rect 2010 1075 2015 1105
rect 1975 1070 2015 1075
rect 795 1060 835 1065
rect 795 1030 800 1060
rect 830 1055 835 1060
rect 905 1060 945 1065
rect 905 1055 910 1060
rect 830 1035 910 1055
rect 830 1030 835 1035
rect 795 1025 835 1030
rect 905 1030 910 1035
rect 940 1030 945 1060
rect 905 1025 945 1030
rect 1155 1010 1195 1015
rect 795 1005 835 1010
rect 795 975 800 1005
rect 830 975 835 1005
rect 795 970 835 975
rect 880 1005 920 1010
rect 880 975 885 1005
rect 915 1000 920 1005
rect 1155 1000 1160 1010
rect 915 980 1160 1000
rect 1190 1005 1195 1010
rect 1840 1010 1880 1015
rect 1840 1005 1845 1010
rect 1190 985 1845 1005
rect 1190 980 1195 985
rect 915 975 920 980
rect 1155 975 1195 980
rect 1840 980 1845 985
rect 1875 980 1880 1010
rect 1840 975 1880 980
rect 880 970 920 975
rect -190 950 -150 955
rect -190 920 -185 950
rect -155 945 -150 950
rect 145 950 175 955
rect -155 925 145 945
rect -155 920 -150 925
rect -190 915 -150 920
rect 1515 950 1545 955
rect 175 925 1515 945
rect 145 915 175 920
rect 1515 915 1545 920
rect -370 900 -330 905
rect -370 870 -365 900
rect -335 895 -330 900
rect 225 900 265 905
rect 225 895 230 900
rect -335 875 230 895
rect -335 870 -330 875
rect -370 865 -330 870
rect 225 870 230 875
rect 260 870 265 900
rect 225 865 265 870
rect 1425 900 1465 905
rect 1425 870 1430 900
rect 1460 895 1465 900
rect 2020 900 2060 905
rect 2020 895 2025 900
rect 1460 875 2025 895
rect 1460 870 1465 875
rect 1425 865 1465 870
rect 2020 870 2025 875
rect 2055 870 2060 900
rect 2020 865 2060 870
rect -280 770 -240 775
rect -1540 760 -1500 765
rect -530 760 -490 765
rect -1540 730 -1535 760
rect -1505 755 -1500 760
rect -970 755 -965 760
rect -1505 735 -965 755
rect -1505 730 -1500 735
rect -970 730 -965 735
rect -935 730 -930 760
rect -530 730 -525 760
rect -495 755 -490 760
rect -280 755 -275 770
rect -495 740 -275 755
rect -245 740 -240 770
rect -495 735 -240 740
rect 1930 760 1970 765
rect -495 730 -490 735
rect -1540 725 -1500 730
rect -530 725 -490 730
rect 1930 730 1935 760
rect 1965 755 1970 760
rect 2180 760 2220 765
rect 3190 760 3230 765
rect 2180 755 2185 760
rect 1965 735 2185 755
rect 1965 730 1970 735
rect 1930 725 1970 730
rect 2180 730 2185 735
rect 2215 730 2220 760
rect 2620 730 2625 760
rect 2655 755 2660 760
rect 3190 755 3195 760
rect 2655 735 3195 755
rect 2655 730 2660 735
rect 3190 730 3195 735
rect 3225 730 3230 760
rect 2180 725 2220 730
rect 3190 725 3230 730
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 710 -1410 715
rect -805 715 -765 720
rect -805 710 -800 715
rect -1415 690 -800 710
rect -1415 685 -1410 690
rect -1450 680 -1410 685
rect -805 685 -800 690
rect -770 710 -765 715
rect -370 715 -330 720
rect -370 710 -365 715
rect -770 690 -365 710
rect -770 685 -765 690
rect -805 680 -765 685
rect -370 685 -365 690
rect -335 685 -330 715
rect -370 680 -330 685
rect 2020 715 2060 720
rect 2020 685 2025 715
rect 2055 710 2060 715
rect 2455 715 2495 720
rect 2455 710 2460 715
rect 2055 690 2460 710
rect 2055 685 2060 690
rect 2020 680 2060 685
rect 2455 685 2460 690
rect 2490 710 2495 715
rect 3100 715 3140 720
rect 3100 710 3105 715
rect 2490 690 3105 710
rect 2490 685 2495 690
rect 2455 680 2495 685
rect 3100 685 3105 690
rect 3135 685 3140 715
rect 3100 680 3140 685
rect -1145 670 -1105 675
rect -1145 640 -1140 670
rect -1110 640 -1105 670
rect -1145 635 -1105 640
rect -530 670 -490 675
rect -530 640 -525 670
rect -495 640 -490 670
rect -530 635 -490 640
rect -465 670 -425 675
rect -465 640 -460 670
rect -430 665 -425 670
rect -235 670 -195 675
rect -235 665 -230 670
rect -430 645 -230 665
rect -430 640 -425 645
rect -465 635 -425 640
rect -235 640 -230 645
rect -200 640 -195 670
rect -235 635 -195 640
rect 1885 670 1925 675
rect 1885 640 1890 670
rect 1920 665 1925 670
rect 2115 670 2155 675
rect 2115 665 2120 670
rect 1920 645 2120 665
rect 1920 640 1925 645
rect 1885 635 1925 640
rect 2115 640 2120 645
rect 2150 640 2155 670
rect 2115 635 2155 640
rect 2180 670 2220 675
rect 2180 640 2185 670
rect 2215 640 2220 670
rect 2180 635 2220 640
rect 2795 670 2835 675
rect 2795 640 2800 670
rect 2830 640 2835 670
rect 2795 635 2835 640
rect -105 625 -65 630
rect -105 595 -100 625
rect -70 610 -65 625
rect 555 625 595 630
rect 555 610 560 625
rect -70 595 560 610
rect 590 610 595 625
rect 1095 625 1135 630
rect 1095 610 1100 625
rect 590 605 755 610
rect 590 595 720 605
rect -105 590 720 595
rect 715 575 720 590
rect 750 575 755 605
rect 715 570 755 575
rect 935 605 1100 610
rect 935 575 940 605
rect 970 595 1100 605
rect 1130 610 1135 625
rect 1755 625 1795 630
rect 1755 610 1760 625
rect 1130 595 1760 610
rect 1790 620 1795 625
rect 1790 615 1970 620
rect 1790 600 1935 615
rect 1790 595 1795 600
rect 970 590 1795 595
rect 970 575 975 590
rect 1930 585 1935 600
rect 1965 585 1970 615
rect 1930 580 1970 585
rect 935 570 975 575
rect 145 550 175 555
rect -105 525 145 545
rect 795 550 825 555
rect 175 525 795 545
rect 145 515 175 520
rect 795 515 825 520
rect 865 550 895 555
rect 1515 550 1545 555
rect 895 525 1515 545
rect 865 515 895 520
rect 1545 525 1795 545
rect 1515 515 1545 520
rect -1270 400 -1230 405
rect -1270 370 -1265 400
rect -1235 395 -1230 400
rect -1025 400 -985 405
rect -1025 395 -1020 400
rect -1235 375 -1020 395
rect -1235 370 -1230 375
rect -1270 365 -1230 370
rect -1025 370 -1020 375
rect -990 370 -985 400
rect -1025 365 -985 370
rect 2675 400 2715 405
rect 2675 370 2680 400
rect 2710 395 2715 400
rect 2920 400 2960 405
rect 2920 395 2925 400
rect 2710 375 2925 395
rect 2710 370 2715 375
rect 2675 365 2715 370
rect 2920 370 2925 375
rect 2955 370 2960 400
rect 2920 365 2960 370
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect 3185 350 3235 360
rect -1545 310 -1495 320
rect -750 340 -710 345
rect -750 310 -745 340
rect -715 335 -710 340
rect -370 340 -330 345
rect -370 335 -365 340
rect -715 315 -365 335
rect -715 310 -710 315
rect -750 305 -710 310
rect -370 310 -365 315
rect -335 310 -330 340
rect -370 305 -330 310
rect 2020 340 2060 345
rect 2020 310 2025 340
rect 2055 335 2060 340
rect 2400 340 2440 345
rect 2400 335 2405 340
rect 2055 315 2405 335
rect 2055 310 2060 315
rect 2020 305 2060 310
rect 2400 310 2405 315
rect 2435 310 2440 340
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2400 305 2440 310
rect 445 285 485 290
rect -1225 280 -1185 285
rect -1225 250 -1220 280
rect -1190 275 -1185 280
rect -1025 280 -985 285
rect -1025 275 -1020 280
rect -1190 255 -1020 275
rect -1190 250 -1185 255
rect -1225 245 -1185 250
rect -1025 250 -1020 255
rect -990 250 -985 280
rect 445 255 450 285
rect 480 280 485 285
rect 1205 285 1245 290
rect 1205 280 1210 285
rect 480 260 1210 280
rect 480 255 485 260
rect 445 250 485 255
rect 1205 255 1210 260
rect 1240 255 1245 285
rect 1205 250 1245 255
rect 2675 280 2715 285
rect 2675 250 2680 280
rect 2710 275 2715 280
rect 2875 280 2915 285
rect 2875 275 2880 280
rect 2710 255 2880 275
rect 2710 250 2715 255
rect -1025 245 -985 250
rect 2675 245 2715 250
rect 2875 250 2880 255
rect 2910 250 2915 280
rect 2875 245 2915 250
rect 780 230 820 235
rect 780 200 785 230
rect 815 225 820 230
rect 870 230 910 235
rect 870 225 875 230
rect 815 205 875 225
rect 815 200 820 205
rect 780 195 820 200
rect 870 200 875 205
rect 905 200 910 230
rect 870 195 910 200
rect 855 175 895 180
rect 855 145 860 175
rect 890 145 895 175
rect 855 140 895 145
rect 795 120 835 125
rect 795 90 800 120
rect 830 90 835 120
rect 795 85 835 90
rect 780 65 820 70
rect 780 35 785 65
rect 815 60 820 65
rect 870 65 910 70
rect 870 60 875 65
rect 815 40 875 60
rect 815 35 820 40
rect 780 30 820 35
rect 870 35 875 40
rect 905 35 910 65
rect 870 30 910 35
rect 440 15 480 20
rect 440 -15 445 15
rect 475 10 480 15
rect 830 15 860 20
rect 475 -10 830 10
rect 475 -15 480 -10
rect 440 -20 480 -15
rect 830 -20 860 -15
rect -1490 -120 -1486 -85
rect -1459 -120 -1426 -85
rect -1399 -120 -1395 -85
rect -1370 -120 -1366 -85
rect -1339 -120 -1335 -85
rect -1310 -120 -1306 -85
rect -1279 -95 -1275 -85
rect -1225 -90 -1185 -85
rect -1225 -95 -1220 -90
rect -1279 -115 -1220 -95
rect -1279 -120 -1275 -115
rect -1225 -120 -1220 -115
rect -1190 -120 -1185 -90
rect -1225 -125 -1185 -120
rect -805 -90 -765 -85
rect -805 -120 -800 -90
rect -770 -95 -765 -90
rect -235 -90 -195 -85
rect -235 -95 -230 -90
rect -770 -115 -230 -95
rect -770 -120 -765 -115
rect -805 -125 -765 -120
rect -235 -120 -230 -115
rect -200 -120 -195 -90
rect -235 -125 -195 -120
rect 1885 -90 1925 -85
rect 1885 -120 1890 -90
rect 1920 -95 1925 -90
rect 2455 -90 2495 -85
rect 2455 -95 2460 -90
rect 1920 -115 2460 -95
rect 1920 -120 1925 -115
rect 1885 -125 1925 -120
rect 2455 -120 2460 -115
rect 2490 -120 2495 -90
rect 2455 -125 2495 -120
rect 2875 -90 2915 -85
rect 2875 -120 2880 -90
rect 2910 -95 2915 -90
rect 2965 -95 2969 -85
rect 2910 -115 2969 -95
rect 2910 -120 2915 -115
rect 2965 -120 2969 -115
rect 2996 -120 3000 -85
rect 3025 -120 3029 -85
rect 3056 -120 3060 -85
rect 3085 -120 3089 -85
rect 3116 -120 3149 -85
rect 3176 -120 3180 -85
rect 2875 -125 2915 -120
rect -1370 -145 -1335 -140
rect -1270 -145 -1230 -140
rect -1270 -150 -1265 -145
rect -1335 -170 -1265 -150
rect -1370 -180 -1335 -175
rect -1270 -175 -1265 -170
rect -1235 -175 -1230 -145
rect -1270 -180 -1230 -175
rect -1145 -145 -1105 -140
rect -1145 -175 -1140 -145
rect -1110 -150 -1105 -145
rect -465 -145 -425 -140
rect -465 -150 -460 -145
rect -1110 -170 -460 -150
rect -1110 -175 -1105 -170
rect -1145 -180 -1105 -175
rect -465 -175 -460 -170
rect -430 -150 -425 -145
rect -280 -145 -240 -140
rect -280 -150 -275 -145
rect -430 -170 -275 -150
rect -430 -175 -425 -170
rect -280 -175 -275 -170
rect -245 -175 -240 -145
rect 1930 -145 1970 -140
rect 1930 -175 1935 -145
rect 1965 -150 1970 -145
rect 2115 -145 2155 -140
rect 2115 -150 2120 -145
rect 1965 -170 2120 -150
rect 1965 -175 1970 -170
rect 2115 -175 2120 -170
rect 2150 -150 2155 -145
rect 2795 -145 2835 -140
rect 2795 -150 2800 -145
rect 2150 -170 2800 -150
rect 2150 -175 2155 -170
rect -465 -180 -425 -175
rect 2115 -180 2155 -175
rect 2795 -175 2800 -170
rect 2830 -175 2835 -145
rect 2795 -180 2835 -175
rect 2920 -145 2960 -140
rect 2920 -175 2925 -145
rect 2955 -150 2960 -145
rect 3025 -145 3060 -140
rect 2955 -170 3025 -150
rect 2955 -175 2960 -170
rect 2920 -180 2960 -175
rect 3025 -180 3060 -175
rect -1490 -190 -1455 -185
rect 3145 -190 3180 -185
rect -325 -195 -320 -190
rect -1455 -215 -320 -195
rect -1490 -225 -1455 -220
rect -325 -220 -320 -215
rect -290 -220 -285 -190
rect -325 -225 -285 -220
rect 1975 -220 1980 -190
rect 2010 -195 2015 -190
rect 2010 -215 3145 -195
rect 2010 -220 2015 -215
rect 1975 -225 2015 -220
rect 3145 -225 3180 -220
rect -1290 -245 -1255 -240
rect -805 -245 -765 -240
rect -805 -250 -800 -245
rect -1255 -270 -800 -250
rect -1290 -280 -1255 -275
rect -805 -275 -800 -270
rect -770 -250 -765 -245
rect -235 -245 -195 -240
rect -235 -250 -230 -245
rect -770 -270 -230 -250
rect -770 -275 -765 -270
rect -805 -280 -765 -275
rect -235 -275 -230 -270
rect -200 -275 -195 -245
rect -235 -280 -195 -275
rect 1885 -245 1925 -240
rect 1885 -275 1890 -245
rect 1920 -250 1925 -245
rect 2455 -245 2495 -240
rect 2455 -250 2460 -245
rect 1920 -270 2460 -250
rect 1920 -275 1925 -270
rect 1885 -280 1925 -275
rect 2455 -275 2460 -270
rect 2490 -250 2495 -245
rect 2945 -245 2980 -240
rect 2490 -270 2945 -250
rect 2490 -275 2495 -270
rect 2455 -280 2495 -275
rect 2945 -280 2980 -275
rect -1540 -305 -1500 -300
rect -1540 -335 -1535 -305
rect -1505 -310 -1500 -305
rect -1230 -305 -1195 -300
rect -1505 -330 -1230 -310
rect -1505 -335 -1500 -330
rect -1540 -340 -1500 -335
rect -1005 -305 -965 -300
rect 2655 -305 2695 -300
rect -1005 -310 -1000 -305
rect -1195 -330 -1000 -310
rect -1230 -340 -1195 -335
rect -1005 -335 -1000 -330
rect -970 -335 -965 -305
rect -1005 -340 -965 -335
rect -105 -310 -65 -305
rect -105 -340 -100 -310
rect -70 -315 -65 -310
rect 595 -310 635 -305
rect 595 -315 600 -310
rect -70 -335 600 -315
rect -70 -340 -65 -335
rect -105 -345 -65 -340
rect 595 -340 600 -335
rect 630 -315 635 -310
rect 825 -310 865 -305
rect 825 -315 830 -310
rect 630 -335 830 -315
rect 630 -340 635 -335
rect 595 -345 635 -340
rect 825 -340 830 -335
rect 860 -315 865 -310
rect 1065 -310 1105 -305
rect 1065 -315 1070 -310
rect 860 -335 1070 -315
rect 860 -340 865 -335
rect 825 -345 865 -340
rect 1065 -340 1070 -335
rect 1100 -315 1105 -310
rect 1750 -310 1790 -305
rect 1750 -315 1755 -310
rect 1100 -335 1755 -315
rect 1100 -340 1105 -335
rect 1065 -345 1105 -340
rect 1750 -340 1755 -335
rect 1785 -315 1790 -310
rect 1930 -310 1970 -305
rect 1930 -315 1935 -310
rect 1785 -335 1935 -315
rect 1785 -340 1790 -335
rect 1750 -345 1790 -340
rect 1930 -340 1935 -335
rect 1965 -340 1970 -310
rect 2655 -335 2660 -305
rect 2690 -310 2695 -305
rect 2885 -305 2920 -300
rect 2690 -330 2885 -310
rect 2690 -335 2695 -330
rect 2655 -340 2695 -335
rect 3190 -305 3230 -300
rect 3190 -310 3195 -305
rect 2920 -330 3195 -310
rect 2885 -340 2920 -335
rect 3190 -335 3195 -330
rect 3225 -335 3230 -305
rect 3190 -340 3230 -335
rect 1930 -345 1970 -340
rect -235 -365 -195 -360
rect -1290 -415 -1286 -380
rect -1259 -415 -1255 -380
rect -1230 -415 -1226 -380
rect -1199 -415 -1195 -380
rect -235 -395 -230 -365
rect -200 -370 -195 -365
rect 1885 -365 1925 -360
rect 1885 -370 1890 -365
rect -200 -390 1890 -370
rect -200 -395 -195 -390
rect -235 -400 -195 -395
rect 1885 -395 1890 -390
rect 1920 -395 1925 -365
rect 1885 -400 1925 -395
rect 2885 -415 2889 -380
rect 2916 -415 2920 -380
rect 2945 -415 2949 -380
rect 2976 -415 2980 -380
rect 1350 -425 1390 -420
rect 1350 -455 1355 -425
rect 1385 -430 1390 -425
rect 1840 -425 1880 -420
rect 1840 -430 1845 -425
rect 1385 -450 1845 -430
rect 1385 -455 1390 -450
rect 1350 -460 1390 -455
rect 1840 -455 1845 -450
rect 1875 -455 1880 -425
rect 1840 -460 1880 -455
rect 1210 -485 1250 -480
rect 1210 -515 1215 -485
rect 1245 -490 1250 -485
rect 1690 -485 1730 -480
rect 1690 -490 1695 -485
rect 1245 -510 1695 -490
rect 1245 -515 1250 -510
rect 1210 -520 1250 -515
rect 1690 -515 1695 -510
rect 1725 -515 1730 -485
rect 1690 -520 1730 -515
rect 265 -805 305 -800
rect 265 -835 270 -805
rect 300 -810 305 -805
rect 1430 -805 1470 -800
rect 1430 -810 1435 -805
rect 300 -830 1435 -810
rect 300 -835 305 -830
rect 265 -840 305 -835
rect 1430 -835 1435 -830
rect 1465 -810 1470 -805
rect 1930 -805 1970 -800
rect 1930 -810 1935 -805
rect 1465 -830 1935 -810
rect 1465 -835 1470 -830
rect 1430 -840 1470 -835
rect 1930 -835 1935 -830
rect 1965 -835 1970 -805
rect 1930 -840 1970 -835
rect -190 -900 -150 -895
rect -190 -930 -185 -900
rect -155 -905 -150 -900
rect 550 -900 590 -895
rect 550 -905 555 -900
rect -155 -925 555 -905
rect -155 -930 -150 -925
rect -190 -935 -150 -930
rect 550 -930 555 -925
rect 585 -905 590 -900
rect 660 -900 700 -895
rect 660 -905 665 -900
rect 585 -925 665 -905
rect 585 -930 590 -925
rect 550 -935 590 -930
rect 660 -930 665 -925
rect 695 -905 700 -900
rect 770 -900 810 -895
rect 770 -905 775 -900
rect 695 -925 775 -905
rect 695 -930 700 -925
rect 660 -935 700 -930
rect 770 -930 775 -925
rect 805 -905 810 -900
rect 1130 -900 1170 -895
rect 1130 -905 1135 -900
rect 805 -925 1135 -905
rect 805 -930 810 -925
rect 770 -935 810 -930
rect 1130 -930 1135 -925
rect 1165 -930 1170 -900
rect 1130 -935 1170 -930
rect 1305 -905 1345 -900
rect 1305 -935 1310 -905
rect 1340 -910 1345 -905
rect 1690 -905 1730 -900
rect 1690 -910 1695 -905
rect 1340 -930 1695 -910
rect 1340 -935 1345 -930
rect 1305 -940 1345 -935
rect 1690 -935 1695 -930
rect 1725 -935 1730 -905
rect 1690 -940 1730 -935
rect 925 -1010 965 -1005
rect 925 -1040 930 -1010
rect 960 -1040 965 -1010
rect 925 -1045 965 -1040
rect -805 -1075 -765 -1070
rect -805 -1105 -800 -1075
rect -770 -1105 -765 -1075
rect -805 -1110 -765 -1105
rect 2455 -1075 2495 -1070
rect 2455 -1105 2460 -1075
rect 2490 -1105 2495 -1075
rect 2455 -1110 2495 -1105
rect 605 -1120 645 -1115
rect 605 -1150 610 -1120
rect 640 -1125 645 -1120
rect 715 -1120 755 -1115
rect 715 -1125 720 -1120
rect 640 -1145 720 -1125
rect 640 -1150 645 -1145
rect 605 -1155 645 -1150
rect 715 -1150 720 -1145
rect 750 -1125 755 -1120
rect 830 -1125 860 -1115
rect 925 -1120 965 -1115
rect 925 -1125 930 -1120
rect 750 -1145 930 -1125
rect 750 -1150 755 -1145
rect 715 -1155 755 -1150
rect 830 -1155 860 -1145
rect 925 -1150 930 -1145
rect 960 -1150 965 -1120
rect 925 -1155 965 -1150
rect -805 -1175 -765 -1170
rect -805 -1205 -800 -1175
rect -770 -1180 -765 -1175
rect -280 -1175 -240 -1170
rect -280 -1180 -275 -1175
rect -770 -1200 -275 -1180
rect -770 -1205 -765 -1200
rect -805 -1210 -765 -1205
rect -280 -1205 -275 -1200
rect -245 -1180 -240 -1175
rect 495 -1175 535 -1170
rect 495 -1180 500 -1175
rect -245 -1200 500 -1180
rect -245 -1205 -240 -1200
rect -280 -1210 -240 -1205
rect 495 -1205 500 -1200
rect 530 -1180 535 -1175
rect 825 -1175 865 -1170
rect 825 -1180 830 -1175
rect 530 -1200 830 -1180
rect 530 -1205 535 -1200
rect 495 -1210 535 -1205
rect 825 -1205 830 -1200
rect 860 -1180 865 -1175
rect 1930 -1175 1970 -1170
rect 1930 -1180 1935 -1175
rect 860 -1200 1935 -1180
rect 860 -1205 865 -1200
rect 825 -1210 865 -1205
rect 1930 -1205 1935 -1200
rect 1965 -1180 1970 -1175
rect 2455 -1175 2495 -1170
rect 2455 -1180 2460 -1175
rect 1965 -1200 2460 -1180
rect 1965 -1205 1970 -1200
rect 1930 -1210 1970 -1205
rect 2455 -1205 2460 -1200
rect 2490 -1205 2495 -1175
rect 2455 -1210 2495 -1205
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via2 >>
rect 830 4245 860 4275
rect -1445 1510 -1415 1540
rect 3105 1460 3135 1490
rect -1535 320 -1505 350
rect 3195 320 3225 350
rect 830 -2455 860 -2425
<< metal3 >>
rect 820 4280 870 4285
rect 820 4240 825 4280
rect 865 4240 870 4280
rect 820 4235 870 4240
rect -3295 3860 -3065 3945
rect -2945 3860 -2715 3945
rect -2595 3860 -2365 3945
rect -3295 3810 -2365 3860
rect -3295 3715 -3065 3810
rect -2945 3715 -2715 3810
rect -2595 3715 -2365 3810
rect -2245 3715 -2015 3945
rect -1895 3715 -1665 3945
rect -1545 3715 -1315 3945
rect -1195 3715 -965 3945
rect -845 3715 -615 3945
rect -495 3715 -265 3945
rect -145 3715 85 3945
rect 205 3715 435 3945
rect 555 3715 785 3945
rect 905 3715 1135 3945
rect 1255 3715 1485 3945
rect 1605 3715 1835 3945
rect 1955 3715 2185 3945
rect 2305 3715 2535 3945
rect 2655 3715 2885 3945
rect 3005 3715 3235 3945
rect 3355 3715 3585 3945
rect 3705 3715 3935 3945
rect 4055 3860 4285 3945
rect 4405 3860 4635 3945
rect 4755 3860 4985 3945
rect 4055 3810 4985 3860
rect 4055 3715 4285 3810
rect 4405 3715 4635 3810
rect 4755 3715 4985 3810
rect -2505 3595 -2455 3715
rect -2155 3595 -2105 3715
rect -1805 3595 -1755 3715
rect -1455 3595 -1405 3715
rect -1105 3595 -1055 3715
rect -755 3595 -705 3715
rect -405 3595 -355 3715
rect -55 3595 -5 3715
rect 295 3595 345 3715
rect 645 3595 695 3715
rect 995 3595 1045 3715
rect 1345 3595 1395 3715
rect 1695 3595 1745 3715
rect 2045 3595 2095 3715
rect 2395 3595 2445 3715
rect 2745 3595 2795 3715
rect 3095 3595 3145 3715
rect 3445 3595 3495 3715
rect 3795 3595 3845 3715
rect 4145 3595 4195 3715
rect -3295 3510 -3065 3595
rect -2945 3510 -2715 3595
rect -2595 3510 -2365 3595
rect -2245 3510 -2015 3595
rect -1895 3510 -1665 3595
rect -1545 3510 -1315 3595
rect -1195 3510 -965 3595
rect -845 3510 -615 3595
rect -495 3510 -265 3595
rect -145 3510 85 3595
rect 205 3510 435 3595
rect 555 3510 785 3595
rect -3295 3460 785 3510
rect -3295 3365 -3065 3460
rect -2945 3365 -2715 3460
rect -2595 3365 -2365 3460
rect -2245 3365 -2015 3460
rect -1895 3365 -1665 3460
rect -1545 3365 -1315 3460
rect -1195 3365 -965 3460
rect -845 3365 -615 3460
rect -495 3365 -265 3460
rect -145 3365 85 3460
rect 205 3365 435 3460
rect 555 3365 785 3460
rect 905 3510 1135 3595
rect 1255 3510 1485 3595
rect 1605 3510 1835 3595
rect 1955 3510 2185 3595
rect 2305 3510 2535 3595
rect 2655 3510 2885 3595
rect 3005 3510 3235 3595
rect 3355 3510 3585 3595
rect 3705 3510 3935 3595
rect 4055 3510 4285 3595
rect 4405 3510 4635 3595
rect 4755 3510 4985 3595
rect 905 3460 4985 3510
rect 905 3365 1135 3460
rect 1255 3365 1485 3460
rect 1605 3365 1835 3460
rect 1955 3365 2185 3460
rect 2305 3365 2535 3460
rect 2655 3365 2885 3460
rect 3005 3365 3235 3460
rect 3355 3365 3585 3460
rect 3705 3365 3935 3460
rect 4055 3365 4285 3460
rect 4405 3365 4635 3460
rect 4755 3365 4985 3460
rect -2505 3245 -2455 3365
rect -1805 3245 -1755 3365
rect -1455 3245 -1405 3365
rect -1105 3245 -1055 3365
rect -755 3245 -705 3365
rect -405 3245 -355 3365
rect -55 3245 -5 3365
rect 295 3245 345 3365
rect 645 3245 695 3365
rect 995 3245 1045 3365
rect 1345 3245 1395 3365
rect 1695 3245 1745 3365
rect 2045 3245 2095 3365
rect 2395 3245 2445 3365
rect 2745 3245 2795 3365
rect 3095 3245 3145 3365
rect 3445 3245 3495 3365
rect 4145 3245 4195 3365
rect -3295 3160 -3065 3245
rect -2945 3160 -2715 3245
rect -2595 3160 -2365 3245
rect -2245 3160 -2015 3245
rect -3295 3110 -2015 3160
rect -3295 3015 -3065 3110
rect -2945 3015 -2715 3110
rect -2595 3015 -2365 3110
rect -2245 3015 -2015 3110
rect -1895 3015 -1665 3245
rect -1545 3015 -1315 3245
rect -1195 3015 -965 3245
rect -845 3015 -615 3245
rect -495 3015 -265 3245
rect -145 3015 85 3245
rect 205 3015 435 3245
rect 555 3015 785 3245
rect 905 3015 1135 3245
rect 1255 3015 1485 3245
rect 1605 3015 1835 3245
rect 1955 3015 2185 3245
rect 2305 3015 2535 3245
rect 2655 3015 2885 3245
rect 3005 3015 3235 3245
rect 3355 3015 3585 3245
rect 3705 3160 3935 3245
rect 4055 3160 4285 3245
rect 4405 3160 4635 3245
rect 4755 3160 4985 3245
rect 3705 3110 4985 3160
rect 3705 3015 3935 3110
rect 4055 3015 4285 3110
rect 4405 3015 4635 3110
rect 4755 3015 4985 3110
rect -2505 2895 -2455 3015
rect -1805 2895 -1755 3015
rect -1455 2895 -1405 3015
rect -1105 2895 -1055 3015
rect -755 2895 -705 3015
rect 2395 2895 2445 3015
rect 2745 2895 2795 3015
rect 3095 2895 3145 3015
rect 3445 2895 3495 3015
rect 4145 2895 4195 3015
rect -3295 2810 -3065 2895
rect -2945 2810 -2715 2895
rect -2595 2810 -2365 2895
rect -2245 2810 -2015 2895
rect -3295 2760 -2015 2810
rect -3295 2665 -3065 2760
rect -2945 2665 -2715 2760
rect -2595 2665 -2365 2760
rect -2245 2665 -2015 2760
rect -1895 2665 -1665 2895
rect -1545 2665 -1315 2895
rect -1195 2665 -965 2895
rect -845 2665 -615 2895
rect 2305 2665 2535 2895
rect 2655 2665 2885 2895
rect 3005 2665 3235 2895
rect 3355 2665 3585 2895
rect 3705 2810 3935 2895
rect 4055 2810 4285 2895
rect 4405 2810 4635 2895
rect 4755 2810 4985 2895
rect 3705 2760 4985 2810
rect 3705 2665 3935 2760
rect 4055 2665 4285 2760
rect 4405 2665 4635 2760
rect 4755 2665 4985 2760
rect -2505 2545 -2455 2665
rect -1455 2545 -1405 2665
rect -1105 2545 -1055 2665
rect -755 2545 -705 2665
rect 2395 2545 2445 2665
rect 2745 2545 2795 2665
rect 3095 2545 3145 2665
rect 4145 2545 4195 2665
rect -3295 2460 -3065 2545
rect -2945 2460 -2715 2545
rect -2595 2460 -2365 2545
rect -2245 2460 -2015 2545
rect -1895 2460 -1665 2545
rect -3295 2410 -1665 2460
rect -3295 2315 -3065 2410
rect -2945 2315 -2715 2410
rect -2595 2315 -2365 2410
rect -2245 2315 -2015 2410
rect -1895 2315 -1665 2410
rect -1545 2315 -1315 2545
rect -1195 2315 -965 2545
rect -845 2315 -615 2545
rect 2305 2315 2535 2545
rect 2655 2315 2885 2545
rect 3005 2315 3235 2545
rect 3355 2460 3585 2545
rect 3705 2460 3935 2545
rect 4055 2460 4285 2545
rect 4405 2460 4635 2545
rect 4755 2460 4985 2545
rect 3355 2410 4985 2460
rect 3355 2315 3585 2410
rect 3705 2315 3935 2410
rect 4055 2315 4285 2410
rect 4405 2315 4635 2410
rect 4755 2315 4985 2410
rect -2505 2195 -2455 2315
rect -3295 2110 -3065 2195
rect -2945 2110 -2715 2195
rect -2595 2110 -2365 2195
rect -2245 2110 -2015 2195
rect -1895 2110 -1665 2195
rect -3295 2060 -1665 2110
rect -3295 1965 -3065 2060
rect -2945 1965 -2715 2060
rect -2595 1965 -2365 2060
rect -2245 1965 -2015 2060
rect -1895 1965 -1665 2060
rect -2505 1845 -2455 1965
rect -3295 1760 -3065 1845
rect -2945 1760 -2715 1845
rect -2595 1760 -2365 1845
rect -2245 1760 -2015 1845
rect -1895 1760 -1665 1845
rect -3295 1710 -1665 1760
rect -3295 1615 -3065 1710
rect -2945 1615 -2715 1710
rect -2595 1615 -2365 1710
rect -2245 1615 -2015 1710
rect -1895 1615 -1665 1710
rect -2505 1495 -2455 1615
rect -1450 1540 -1410 2315
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -3295 1410 -3065 1495
rect -2945 1410 -2715 1495
rect -2595 1410 -2365 1495
rect -2245 1410 -2015 1495
rect -1895 1410 -1665 1495
rect 3100 1490 3140 2315
rect 4145 2195 4195 2315
rect 3355 2110 3585 2195
rect 3705 2110 3935 2195
rect 4055 2110 4285 2195
rect 4405 2110 4635 2195
rect 4755 2110 4985 2195
rect 3355 2060 4985 2110
rect 3355 1965 3585 2060
rect 3705 1965 3935 2060
rect 4055 1965 4285 2060
rect 4405 1965 4635 2060
rect 4755 1965 4985 2060
rect 4145 1845 4195 1965
rect 3355 1760 3585 1845
rect 3705 1760 3935 1845
rect 4055 1760 4285 1845
rect 4405 1760 4635 1845
rect 4755 1760 4985 1845
rect 3355 1710 4985 1760
rect 3355 1615 3585 1710
rect 3705 1615 3935 1710
rect 4055 1615 4285 1710
rect 4405 1615 4635 1710
rect 4755 1615 4985 1710
rect 4145 1495 4195 1615
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect -3295 1360 -1665 1410
rect -3295 1265 -3065 1360
rect -2945 1265 -2715 1360
rect -2595 1265 -2365 1360
rect -2245 1265 -2015 1360
rect -1895 1265 -1665 1360
rect 3355 1410 3585 1495
rect 3705 1410 3935 1495
rect 4055 1410 4285 1495
rect 4405 1410 4635 1495
rect 4755 1410 4985 1495
rect 3355 1360 4985 1410
rect 3355 1265 3585 1360
rect 3705 1265 3935 1360
rect 4055 1265 4285 1360
rect 4405 1265 4635 1360
rect 4755 1265 4985 1360
rect -2505 1145 -2455 1265
rect 4145 1145 4195 1265
rect -3295 1060 -3065 1145
rect -2945 1060 -2715 1145
rect -2595 1060 -2365 1145
rect -2245 1060 -2015 1145
rect -1895 1060 -1665 1145
rect -3295 1010 -1665 1060
rect -3295 915 -3065 1010
rect -2945 915 -2715 1010
rect -2595 915 -2365 1010
rect -2245 915 -2015 1010
rect -1895 915 -1665 1010
rect 3355 1060 3585 1145
rect 3705 1060 3935 1145
rect 4055 1060 4285 1145
rect 4405 1060 4635 1145
rect 4755 1060 4985 1145
rect 3355 1010 4985 1060
rect 3355 915 3585 1010
rect 3705 915 3935 1010
rect 4055 915 4285 1010
rect 4405 915 4635 1010
rect 4755 915 4985 1010
rect -2505 795 -2455 915
rect 4145 795 4195 915
rect -3295 710 -3065 795
rect -2945 710 -2715 795
rect -2595 710 -2365 795
rect -2245 710 -2015 795
rect -1895 710 -1665 795
rect -3295 660 -1665 710
rect -3295 565 -3065 660
rect -2945 565 -2715 660
rect -2595 565 -2365 660
rect -2245 565 -2015 660
rect -1895 565 -1665 660
rect 3355 710 3585 795
rect 3705 710 3935 795
rect 4055 710 4285 795
rect 4405 710 4635 795
rect 4755 710 4985 795
rect 3355 660 4985 710
rect 3355 565 3585 660
rect 3705 565 3935 660
rect 4055 565 4285 660
rect 4405 565 4635 660
rect 4755 565 4985 660
rect -2505 445 -2455 565
rect 4145 445 4195 565
rect -3295 360 -3065 445
rect -2945 360 -2715 445
rect -2595 360 -2365 445
rect -2245 360 -2015 445
rect -1895 360 -1665 445
rect 3355 360 3585 445
rect 3705 360 3935 445
rect 4055 360 4285 445
rect 4405 360 4635 445
rect 4755 360 4985 445
rect -3295 310 -1665 360
rect -1545 355 -1495 360
rect -1545 315 -1540 355
rect -1500 315 -1495 355
rect -1545 310 -1495 315
rect 3185 355 3235 360
rect 3185 315 3190 355
rect 3230 315 3235 355
rect 3185 310 3235 315
rect 3355 310 4985 360
rect -3295 215 -3065 310
rect -2945 215 -2715 310
rect -2595 215 -2365 310
rect -2245 215 -2015 310
rect -1895 215 -1665 310
rect 3355 215 3585 310
rect 3705 215 3935 310
rect 4055 215 4285 310
rect 4405 215 4635 310
rect 4755 215 4985 310
rect -2505 95 -2455 215
rect 4145 95 4195 215
rect -3295 10 -3065 95
rect -2945 10 -2715 95
rect -2595 10 -2365 95
rect -2245 10 -2015 95
rect -1895 10 -1665 95
rect -3295 -40 -1665 10
rect -3295 -135 -3065 -40
rect -2945 -135 -2715 -40
rect -2595 -135 -2365 -40
rect -2245 -135 -2015 -40
rect -1895 -135 -1665 -40
rect 3355 10 3585 95
rect 3705 10 3935 95
rect 4055 10 4285 95
rect 4405 10 4635 95
rect 4755 10 4985 95
rect 3355 -40 4985 10
rect 3355 -135 3585 -40
rect 3705 -135 3935 -40
rect 4055 -135 4285 -40
rect 4405 -135 4635 -40
rect 4755 -135 4985 -40
rect -2505 -255 -2455 -135
rect 4145 -255 4195 -135
rect -3295 -340 -3065 -255
rect -2945 -340 -2715 -255
rect -2595 -340 -2365 -255
rect -2245 -340 -2015 -255
rect -1895 -340 -1665 -255
rect -3295 -390 -1665 -340
rect -3295 -485 -3065 -390
rect -2945 -485 -2715 -390
rect -2595 -485 -2365 -390
rect -2245 -485 -2015 -390
rect -1895 -485 -1665 -390
rect 3355 -340 3585 -255
rect 3705 -340 3935 -255
rect 4055 -340 4285 -255
rect 4405 -340 4635 -255
rect 4755 -340 4985 -255
rect 3355 -390 4985 -340
rect 3355 -485 3585 -390
rect 3705 -485 3935 -390
rect 4055 -485 4285 -390
rect 4405 -485 4635 -390
rect 4755 -485 4985 -390
rect -2505 -605 -2455 -485
rect 4145 -605 4195 -485
rect -3295 -690 -3065 -605
rect -2945 -690 -2715 -605
rect -2595 -690 -2365 -605
rect -2245 -690 -2015 -605
rect -1895 -690 -1665 -605
rect -3295 -740 -1665 -690
rect -3295 -835 -3065 -740
rect -2945 -835 -2715 -740
rect -2595 -835 -2365 -740
rect -2245 -835 -2015 -740
rect -1895 -835 -1665 -740
rect 3355 -690 3585 -605
rect 3705 -690 3935 -605
rect 4055 -690 4285 -605
rect 4405 -690 4635 -605
rect 4755 -690 4985 -605
rect 3355 -740 4985 -690
rect 3355 -835 3585 -740
rect 3705 -835 3935 -740
rect 4055 -835 4285 -740
rect 4405 -835 4635 -740
rect 4755 -835 4985 -740
rect -2505 -955 -2455 -835
rect 4145 -955 4195 -835
rect -3295 -1040 -3065 -955
rect -2945 -1040 -2715 -955
rect -2595 -1040 -2365 -955
rect -2245 -1040 -2015 -955
rect -1895 -1040 -1665 -955
rect -3295 -1090 -1665 -1040
rect -3295 -1185 -3065 -1090
rect -2945 -1185 -2715 -1090
rect -2595 -1185 -2365 -1090
rect -2245 -1185 -2015 -1090
rect -1895 -1185 -1665 -1090
rect 3355 -1040 3585 -955
rect 3705 -1040 3935 -955
rect 4055 -1040 4285 -955
rect 4405 -1040 4635 -955
rect 4755 -1040 4985 -955
rect 3355 -1090 4985 -1040
rect 3355 -1185 3585 -1090
rect 3705 -1185 3935 -1090
rect 4055 -1185 4285 -1090
rect 4405 -1185 4635 -1090
rect 4755 -1185 4985 -1090
rect -2505 -1305 -2455 -1185
rect 4145 -1305 4195 -1185
rect -3295 -1390 -3065 -1305
rect -2945 -1390 -2715 -1305
rect -2595 -1390 -2365 -1305
rect -2245 -1390 -2015 -1305
rect -1895 -1390 -1665 -1305
rect -3295 -1440 -1665 -1390
rect -3295 -1535 -3065 -1440
rect -2945 -1535 -2715 -1440
rect -2595 -1535 -2365 -1440
rect -2245 -1535 -2015 -1440
rect -1895 -1535 -1665 -1440
rect -1545 -1535 -1315 -1305
rect -1195 -1535 -965 -1305
rect -845 -1535 -615 -1305
rect -495 -1535 -265 -1305
rect -145 -1535 85 -1305
rect 205 -1535 435 -1305
rect 555 -1535 785 -1305
rect 905 -1535 1135 -1305
rect 1255 -1535 1485 -1305
rect 1605 -1535 1835 -1305
rect 1955 -1535 2185 -1305
rect 2305 -1535 2535 -1305
rect 2655 -1535 2885 -1305
rect 3005 -1535 3235 -1305
rect 3355 -1390 3585 -1305
rect 3705 -1390 3935 -1305
rect 4055 -1390 4285 -1305
rect 4405 -1390 4635 -1305
rect 4755 -1390 4985 -1305
rect 3355 -1440 4985 -1390
rect 3355 -1535 3585 -1440
rect 3705 -1535 3935 -1440
rect 4055 -1535 4285 -1440
rect 4405 -1535 4635 -1440
rect 4755 -1535 4985 -1440
rect -2505 -1655 -2455 -1535
rect -1455 -1655 -1405 -1535
rect -1105 -1655 -1055 -1535
rect -755 -1655 -705 -1535
rect -405 -1655 -355 -1535
rect -55 -1655 -5 -1535
rect 295 -1655 345 -1535
rect 645 -1655 695 -1535
rect 995 -1655 1045 -1535
rect 1345 -1655 1395 -1535
rect 1695 -1655 1745 -1535
rect 2045 -1655 2095 -1535
rect 2395 -1655 2445 -1535
rect 2745 -1655 2795 -1535
rect 3095 -1655 3145 -1535
rect 4145 -1655 4195 -1535
rect -3295 -1740 -3065 -1655
rect -2945 -1740 -2715 -1655
rect -2595 -1740 -2365 -1655
rect -2245 -1740 -2015 -1655
rect -1895 -1740 -1665 -1655
rect -1545 -1740 -1315 -1655
rect -1195 -1740 -965 -1655
rect -845 -1740 -615 -1655
rect -495 -1740 -265 -1655
rect -145 -1740 85 -1655
rect 205 -1740 435 -1655
rect 555 -1740 785 -1655
rect -3295 -1790 785 -1740
rect -3295 -1885 -3065 -1790
rect -2945 -1885 -2715 -1790
rect -2595 -1885 -2365 -1790
rect -2245 -1885 -2015 -1790
rect -1895 -1885 -1665 -1790
rect -1545 -1885 -1315 -1790
rect -1195 -1885 -965 -1790
rect -845 -1885 -615 -1790
rect -495 -1885 -265 -1790
rect -145 -1885 85 -1790
rect 205 -1885 435 -1790
rect 555 -1885 785 -1790
rect 905 -1740 1135 -1655
rect 1255 -1740 1485 -1655
rect 1605 -1740 1835 -1655
rect 1955 -1740 2185 -1655
rect 2305 -1740 2535 -1655
rect 2655 -1740 2885 -1655
rect 3005 -1740 3235 -1655
rect 3355 -1740 3585 -1655
rect 3705 -1740 3935 -1655
rect 4055 -1740 4285 -1655
rect 4405 -1740 4635 -1655
rect 4755 -1740 4985 -1655
rect 905 -1790 4985 -1740
rect 905 -1885 1135 -1790
rect 1255 -1885 1485 -1790
rect 1605 -1885 1835 -1790
rect 1955 -1885 2185 -1790
rect 2305 -1885 2535 -1790
rect 2655 -1885 2885 -1790
rect 3005 -1885 3235 -1790
rect 3355 -1885 3585 -1790
rect 3705 -1885 3935 -1790
rect 4055 -1885 4285 -1790
rect 4405 -1885 4635 -1790
rect 4755 -1885 4985 -1790
rect -2505 -2005 -2455 -1885
rect -2155 -2005 -2105 -1885
rect -1805 -2005 -1755 -1885
rect -1455 -2005 -1405 -1885
rect -1105 -2005 -1055 -1885
rect -755 -2005 -705 -1885
rect -405 -2005 -355 -1885
rect -55 -2005 -5 -1885
rect 295 -2005 345 -1885
rect 645 -2005 695 -1885
rect 995 -2005 1045 -1885
rect 1345 -2005 1395 -1885
rect 1695 -2005 1745 -1885
rect 2045 -2005 2095 -1885
rect 2395 -2005 2445 -1885
rect 2745 -2005 2795 -1885
rect 3095 -2005 3145 -1885
rect 3445 -2005 3495 -1885
rect 3795 -2005 3845 -1885
rect 4145 -2005 4195 -1885
rect -3295 -2090 -3065 -2005
rect -2945 -2090 -2715 -2005
rect -2595 -2090 -2365 -2005
rect -3295 -2140 -2365 -2090
rect -3295 -2235 -3065 -2140
rect -2945 -2235 -2715 -2140
rect -2595 -2235 -2365 -2140
rect -2245 -2235 -2015 -2005
rect -1895 -2235 -1665 -2005
rect -1545 -2235 -1315 -2005
rect -1195 -2235 -965 -2005
rect -845 -2235 -615 -2005
rect -495 -2235 -265 -2005
rect -145 -2235 85 -2005
rect 205 -2235 435 -2005
rect 555 -2235 785 -2005
rect 905 -2235 1135 -2005
rect 1255 -2235 1485 -2005
rect 1605 -2235 1835 -2005
rect 1955 -2235 2185 -2005
rect 2305 -2235 2535 -2005
rect 2655 -2235 2885 -2005
rect 3005 -2235 3235 -2005
rect 3355 -2235 3585 -2005
rect 3705 -2235 3935 -2005
rect 4055 -2090 4285 -2005
rect 4405 -2090 4635 -2005
rect 4755 -2090 4985 -2005
rect 4055 -2140 4985 -2090
rect 4055 -2235 4285 -2140
rect 4405 -2235 4635 -2140
rect 4755 -2235 4985 -2140
rect 820 -2420 870 -2415
rect 820 -2460 825 -2420
rect 865 -2460 870 -2420
rect 820 -2465 870 -2460
<< via3 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 830 4245 860 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect -1540 350 -1500 355
rect -1540 320 -1535 350
rect -1535 320 -1505 350
rect -1505 320 -1500 350
rect -1540 315 -1500 320
rect 3190 350 3230 355
rect 3190 320 3195 350
rect 3195 320 3225 350
rect 3225 320 3230 350
rect 3190 315 3230 320
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 830 -2455 860 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< mimcap >>
rect -3280 3855 -3080 3930
rect -3280 3815 -3200 3855
rect -3160 3815 -3080 3855
rect -3280 3730 -3080 3815
rect -2930 3855 -2730 3930
rect -2930 3815 -2850 3855
rect -2810 3815 -2730 3855
rect -2930 3730 -2730 3815
rect -2580 3855 -2380 3930
rect -2580 3815 -2500 3855
rect -2460 3815 -2380 3855
rect -2580 3730 -2380 3815
rect -2230 3855 -2030 3930
rect -2230 3815 -2150 3855
rect -2110 3815 -2030 3855
rect -2230 3730 -2030 3815
rect -1880 3855 -1680 3930
rect -1880 3815 -1800 3855
rect -1760 3815 -1680 3855
rect -1880 3730 -1680 3815
rect -1530 3855 -1330 3930
rect -1530 3815 -1450 3855
rect -1410 3815 -1330 3855
rect -1530 3730 -1330 3815
rect -1180 3855 -980 3930
rect -1180 3815 -1100 3855
rect -1060 3815 -980 3855
rect -1180 3730 -980 3815
rect -830 3855 -630 3930
rect -830 3815 -750 3855
rect -710 3815 -630 3855
rect -830 3730 -630 3815
rect -480 3855 -280 3930
rect -480 3815 -400 3855
rect -360 3815 -280 3855
rect -480 3730 -280 3815
rect -130 3855 70 3930
rect -130 3815 -50 3855
rect -10 3815 70 3855
rect -130 3730 70 3815
rect 220 3855 420 3930
rect 220 3815 300 3855
rect 340 3815 420 3855
rect 220 3730 420 3815
rect 570 3855 770 3930
rect 570 3815 650 3855
rect 690 3815 770 3855
rect 570 3730 770 3815
rect 920 3855 1120 3930
rect 920 3815 1000 3855
rect 1040 3815 1120 3855
rect 920 3730 1120 3815
rect 1270 3855 1470 3930
rect 1270 3815 1350 3855
rect 1390 3815 1470 3855
rect 1270 3730 1470 3815
rect 1620 3855 1820 3930
rect 1620 3815 1700 3855
rect 1740 3815 1820 3855
rect 1620 3730 1820 3815
rect 1970 3855 2170 3930
rect 1970 3815 2050 3855
rect 2090 3815 2170 3855
rect 1970 3730 2170 3815
rect 2320 3855 2520 3930
rect 2320 3815 2400 3855
rect 2440 3815 2520 3855
rect 2320 3730 2520 3815
rect 2670 3855 2870 3930
rect 2670 3815 2750 3855
rect 2790 3815 2870 3855
rect 2670 3730 2870 3815
rect 3020 3855 3220 3930
rect 3020 3815 3100 3855
rect 3140 3815 3220 3855
rect 3020 3730 3220 3815
rect 3370 3855 3570 3930
rect 3370 3815 3450 3855
rect 3490 3815 3570 3855
rect 3370 3730 3570 3815
rect 3720 3855 3920 3930
rect 3720 3815 3800 3855
rect 3840 3815 3920 3855
rect 3720 3730 3920 3815
rect 4070 3855 4270 3930
rect 4070 3815 4150 3855
rect 4190 3815 4270 3855
rect 4070 3730 4270 3815
rect 4420 3855 4620 3930
rect 4420 3815 4500 3855
rect 4540 3815 4620 3855
rect 4420 3730 4620 3815
rect 4770 3855 4970 3930
rect 4770 3815 4850 3855
rect 4890 3815 4970 3855
rect 4770 3730 4970 3815
rect -3280 3505 -3080 3580
rect -3280 3465 -3200 3505
rect -3160 3465 -3080 3505
rect -3280 3380 -3080 3465
rect -2930 3505 -2730 3580
rect -2930 3465 -2850 3505
rect -2810 3465 -2730 3505
rect -2930 3380 -2730 3465
rect -2580 3505 -2380 3580
rect -2580 3465 -2500 3505
rect -2460 3465 -2380 3505
rect -2580 3380 -2380 3465
rect -2230 3505 -2030 3580
rect -2230 3465 -2150 3505
rect -2110 3465 -2030 3505
rect -2230 3380 -2030 3465
rect -1880 3505 -1680 3580
rect -1880 3465 -1800 3505
rect -1760 3465 -1680 3505
rect -1880 3380 -1680 3465
rect -1530 3505 -1330 3580
rect -1530 3465 -1450 3505
rect -1410 3465 -1330 3505
rect -1530 3380 -1330 3465
rect -1180 3505 -980 3580
rect -1180 3465 -1100 3505
rect -1060 3465 -980 3505
rect -1180 3380 -980 3465
rect -830 3505 -630 3580
rect -830 3465 -750 3505
rect -710 3465 -630 3505
rect -830 3380 -630 3465
rect -480 3505 -280 3580
rect -480 3465 -400 3505
rect -360 3465 -280 3505
rect -480 3380 -280 3465
rect -130 3505 70 3580
rect -130 3465 -50 3505
rect -10 3465 70 3505
rect -130 3380 70 3465
rect 220 3505 420 3580
rect 220 3465 300 3505
rect 340 3465 420 3505
rect 220 3380 420 3465
rect 570 3505 770 3580
rect 570 3465 650 3505
rect 690 3465 770 3505
rect 570 3380 770 3465
rect 920 3505 1120 3580
rect 920 3465 1000 3505
rect 1040 3465 1120 3505
rect 920 3380 1120 3465
rect 1270 3505 1470 3580
rect 1270 3465 1350 3505
rect 1390 3465 1470 3505
rect 1270 3380 1470 3465
rect 1620 3505 1820 3580
rect 1620 3465 1700 3505
rect 1740 3465 1820 3505
rect 1620 3380 1820 3465
rect 1970 3505 2170 3580
rect 1970 3465 2050 3505
rect 2090 3465 2170 3505
rect 1970 3380 2170 3465
rect 2320 3505 2520 3580
rect 2320 3465 2400 3505
rect 2440 3465 2520 3505
rect 2320 3380 2520 3465
rect 2670 3505 2870 3580
rect 2670 3465 2750 3505
rect 2790 3465 2870 3505
rect 2670 3380 2870 3465
rect 3020 3505 3220 3580
rect 3020 3465 3100 3505
rect 3140 3465 3220 3505
rect 3020 3380 3220 3465
rect 3370 3505 3570 3580
rect 3370 3465 3450 3505
rect 3490 3465 3570 3505
rect 3370 3380 3570 3465
rect 3720 3505 3920 3580
rect 3720 3465 3800 3505
rect 3840 3465 3920 3505
rect 3720 3380 3920 3465
rect 4070 3505 4270 3580
rect 4070 3465 4150 3505
rect 4190 3465 4270 3505
rect 4070 3380 4270 3465
rect 4420 3505 4620 3580
rect 4420 3465 4500 3505
rect 4540 3465 4620 3505
rect 4420 3380 4620 3465
rect 4770 3505 4970 3580
rect 4770 3465 4850 3505
rect 4890 3465 4970 3505
rect 4770 3380 4970 3465
rect -3280 3155 -3080 3230
rect -3280 3115 -3200 3155
rect -3160 3115 -3080 3155
rect -3280 3030 -3080 3115
rect -2930 3155 -2730 3230
rect -2930 3115 -2850 3155
rect -2810 3115 -2730 3155
rect -2930 3030 -2730 3115
rect -2580 3155 -2380 3230
rect -2580 3115 -2500 3155
rect -2460 3115 -2380 3155
rect -2580 3030 -2380 3115
rect -2230 3155 -2030 3230
rect -2230 3115 -2150 3155
rect -2110 3115 -2030 3155
rect -2230 3030 -2030 3115
rect -1880 3155 -1680 3230
rect -1880 3115 -1800 3155
rect -1760 3115 -1680 3155
rect -1880 3030 -1680 3115
rect -1530 3155 -1330 3230
rect -1530 3115 -1450 3155
rect -1410 3115 -1330 3155
rect -1530 3030 -1330 3115
rect -1180 3155 -980 3230
rect -1180 3115 -1100 3155
rect -1060 3115 -980 3155
rect -1180 3030 -980 3115
rect -830 3155 -630 3230
rect -830 3115 -750 3155
rect -710 3115 -630 3155
rect -830 3030 -630 3115
rect -480 3155 -280 3230
rect -480 3115 -400 3155
rect -360 3115 -280 3155
rect -480 3030 -280 3115
rect -130 3145 70 3230
rect -130 3105 -50 3145
rect -10 3105 70 3145
rect -130 3030 70 3105
rect 220 3145 420 3230
rect 220 3105 300 3145
rect 340 3105 420 3145
rect 220 3030 420 3105
rect 570 3145 770 3230
rect 570 3105 650 3145
rect 690 3105 770 3145
rect 570 3030 770 3105
rect 920 3145 1120 3230
rect 920 3105 1000 3145
rect 1040 3105 1120 3145
rect 920 3030 1120 3105
rect 1270 3145 1470 3230
rect 1270 3105 1350 3145
rect 1390 3105 1470 3145
rect 1270 3030 1470 3105
rect 1620 3145 1820 3230
rect 1620 3105 1700 3145
rect 1740 3105 1820 3145
rect 1620 3030 1820 3105
rect 1970 3155 2170 3230
rect 1970 3115 2050 3155
rect 2090 3115 2170 3155
rect 1970 3030 2170 3115
rect 2320 3155 2520 3230
rect 2320 3115 2400 3155
rect 2440 3115 2520 3155
rect 2320 3030 2520 3115
rect 2670 3155 2870 3230
rect 2670 3115 2750 3155
rect 2790 3115 2870 3155
rect 2670 3030 2870 3115
rect 3020 3155 3220 3230
rect 3020 3115 3100 3155
rect 3140 3115 3220 3155
rect 3020 3030 3220 3115
rect 3370 3155 3570 3230
rect 3370 3115 3450 3155
rect 3490 3115 3570 3155
rect 3370 3030 3570 3115
rect 3720 3155 3920 3230
rect 3720 3115 3800 3155
rect 3840 3115 3920 3155
rect 3720 3030 3920 3115
rect 4070 3155 4270 3230
rect 4070 3115 4150 3155
rect 4190 3115 4270 3155
rect 4070 3030 4270 3115
rect 4420 3155 4620 3230
rect 4420 3115 4500 3155
rect 4540 3115 4620 3155
rect 4420 3030 4620 3115
rect 4770 3155 4970 3230
rect 4770 3115 4850 3155
rect 4890 3115 4970 3155
rect 4770 3030 4970 3115
rect -3280 2805 -3080 2880
rect -3280 2765 -3200 2805
rect -3160 2765 -3080 2805
rect -3280 2680 -3080 2765
rect -2930 2805 -2730 2880
rect -2930 2765 -2850 2805
rect -2810 2765 -2730 2805
rect -2930 2680 -2730 2765
rect -2580 2805 -2380 2880
rect -2580 2765 -2500 2805
rect -2460 2765 -2380 2805
rect -2580 2680 -2380 2765
rect -2230 2805 -2030 2880
rect -2230 2765 -2150 2805
rect -2110 2765 -2030 2805
rect -2230 2680 -2030 2765
rect -1880 2805 -1680 2880
rect -1880 2765 -1800 2805
rect -1760 2765 -1680 2805
rect -1880 2680 -1680 2765
rect -1530 2805 -1330 2880
rect -1530 2765 -1450 2805
rect -1410 2765 -1330 2805
rect -1530 2680 -1330 2765
rect -1180 2805 -980 2880
rect -1180 2765 -1100 2805
rect -1060 2765 -980 2805
rect -1180 2680 -980 2765
rect -830 2805 -630 2880
rect -830 2765 -750 2805
rect -710 2765 -630 2805
rect -830 2680 -630 2765
rect 2320 2805 2520 2880
rect 2320 2765 2400 2805
rect 2440 2765 2520 2805
rect 2320 2680 2520 2765
rect 2670 2805 2870 2880
rect 2670 2765 2750 2805
rect 2790 2765 2870 2805
rect 2670 2680 2870 2765
rect 3020 2805 3220 2880
rect 3020 2765 3100 2805
rect 3140 2765 3220 2805
rect 3020 2680 3220 2765
rect 3370 2805 3570 2880
rect 3370 2765 3450 2805
rect 3490 2765 3570 2805
rect 3370 2680 3570 2765
rect 3720 2805 3920 2880
rect 3720 2765 3800 2805
rect 3840 2765 3920 2805
rect 3720 2680 3920 2765
rect 4070 2805 4270 2880
rect 4070 2765 4150 2805
rect 4190 2765 4270 2805
rect 4070 2680 4270 2765
rect 4420 2805 4620 2880
rect 4420 2765 4500 2805
rect 4540 2765 4620 2805
rect 4420 2680 4620 2765
rect 4770 2805 4970 2880
rect 4770 2765 4850 2805
rect 4890 2765 4970 2805
rect 4770 2680 4970 2765
rect -3280 2455 -3080 2530
rect -3280 2415 -3200 2455
rect -3160 2415 -3080 2455
rect -3280 2330 -3080 2415
rect -2930 2455 -2730 2530
rect -2930 2415 -2850 2455
rect -2810 2415 -2730 2455
rect -2930 2330 -2730 2415
rect -2580 2455 -2380 2530
rect -2580 2415 -2500 2455
rect -2460 2415 -2380 2455
rect -2580 2330 -2380 2415
rect -2230 2455 -2030 2530
rect -2230 2415 -2150 2455
rect -2110 2415 -2030 2455
rect -2230 2330 -2030 2415
rect -1880 2455 -1680 2530
rect -1880 2415 -1800 2455
rect -1760 2415 -1680 2455
rect -1880 2330 -1680 2415
rect -1530 2455 -1330 2530
rect -1530 2415 -1450 2455
rect -1410 2415 -1330 2455
rect -1530 2330 -1330 2415
rect -1180 2455 -980 2530
rect -1180 2415 -1100 2455
rect -1060 2415 -980 2455
rect -1180 2330 -980 2415
rect -830 2455 -630 2530
rect -830 2415 -750 2455
rect -710 2415 -630 2455
rect -830 2330 -630 2415
rect 2320 2455 2520 2530
rect 2320 2415 2400 2455
rect 2440 2415 2520 2455
rect 2320 2330 2520 2415
rect 2670 2455 2870 2530
rect 2670 2415 2750 2455
rect 2790 2415 2870 2455
rect 2670 2330 2870 2415
rect 3020 2455 3220 2530
rect 3020 2415 3100 2455
rect 3140 2415 3220 2455
rect 3020 2330 3220 2415
rect 3370 2455 3570 2530
rect 3370 2415 3450 2455
rect 3490 2415 3570 2455
rect 3370 2330 3570 2415
rect 3720 2455 3920 2530
rect 3720 2415 3800 2455
rect 3840 2415 3920 2455
rect 3720 2330 3920 2415
rect 4070 2455 4270 2530
rect 4070 2415 4150 2455
rect 4190 2415 4270 2455
rect 4070 2330 4270 2415
rect 4420 2455 4620 2530
rect 4420 2415 4500 2455
rect 4540 2415 4620 2455
rect 4420 2330 4620 2415
rect 4770 2455 4970 2530
rect 4770 2415 4850 2455
rect 4890 2415 4970 2455
rect 4770 2330 4970 2415
rect -3280 2105 -3080 2180
rect -3280 2065 -3200 2105
rect -3160 2065 -3080 2105
rect -3280 1980 -3080 2065
rect -2930 2105 -2730 2180
rect -2930 2065 -2850 2105
rect -2810 2065 -2730 2105
rect -2930 1980 -2730 2065
rect -2580 2105 -2380 2180
rect -2580 2065 -2500 2105
rect -2460 2065 -2380 2105
rect -2580 1980 -2380 2065
rect -2230 2105 -2030 2180
rect -2230 2065 -2150 2105
rect -2110 2065 -2030 2105
rect -2230 1980 -2030 2065
rect -1880 2105 -1680 2180
rect -1880 2065 -1800 2105
rect -1760 2065 -1680 2105
rect -1880 1980 -1680 2065
rect 3370 2105 3570 2180
rect 3370 2065 3450 2105
rect 3490 2065 3570 2105
rect 3370 1980 3570 2065
rect 3720 2105 3920 2180
rect 3720 2065 3800 2105
rect 3840 2065 3920 2105
rect 3720 1980 3920 2065
rect 4070 2105 4270 2180
rect 4070 2065 4150 2105
rect 4190 2065 4270 2105
rect 4070 1980 4270 2065
rect 4420 2105 4620 2180
rect 4420 2065 4500 2105
rect 4540 2065 4620 2105
rect 4420 1980 4620 2065
rect 4770 2105 4970 2180
rect 4770 2065 4850 2105
rect 4890 2065 4970 2105
rect 4770 1980 4970 2065
rect -3280 1755 -3080 1830
rect -3280 1715 -3200 1755
rect -3160 1715 -3080 1755
rect -3280 1630 -3080 1715
rect -2930 1755 -2730 1830
rect -2930 1715 -2850 1755
rect -2810 1715 -2730 1755
rect -2930 1630 -2730 1715
rect -2580 1755 -2380 1830
rect -2580 1715 -2500 1755
rect -2460 1715 -2380 1755
rect -2580 1630 -2380 1715
rect -2230 1755 -2030 1830
rect -2230 1715 -2150 1755
rect -2110 1715 -2030 1755
rect -2230 1630 -2030 1715
rect -1880 1755 -1680 1830
rect -1880 1715 -1800 1755
rect -1760 1715 -1680 1755
rect -1880 1630 -1680 1715
rect 3370 1755 3570 1830
rect 3370 1715 3450 1755
rect 3490 1715 3570 1755
rect 3370 1630 3570 1715
rect 3720 1755 3920 1830
rect 3720 1715 3800 1755
rect 3840 1715 3920 1755
rect 3720 1630 3920 1715
rect 4070 1755 4270 1830
rect 4070 1715 4150 1755
rect 4190 1715 4270 1755
rect 4070 1630 4270 1715
rect 4420 1755 4620 1830
rect 4420 1715 4500 1755
rect 4540 1715 4620 1755
rect 4420 1630 4620 1715
rect 4770 1755 4970 1830
rect 4770 1715 4850 1755
rect 4890 1715 4970 1755
rect 4770 1630 4970 1715
rect -3280 1405 -3080 1480
rect -3280 1365 -3200 1405
rect -3160 1365 -3080 1405
rect -3280 1280 -3080 1365
rect -2930 1405 -2730 1480
rect -2930 1365 -2850 1405
rect -2810 1365 -2730 1405
rect -2930 1280 -2730 1365
rect -2580 1405 -2380 1480
rect -2580 1365 -2500 1405
rect -2460 1365 -2380 1405
rect -2580 1280 -2380 1365
rect -2230 1405 -2030 1480
rect -2230 1365 -2150 1405
rect -2110 1365 -2030 1405
rect -2230 1280 -2030 1365
rect -1880 1405 -1680 1480
rect -1880 1365 -1800 1405
rect -1760 1365 -1680 1405
rect -1880 1280 -1680 1365
rect 3370 1405 3570 1480
rect 3370 1365 3450 1405
rect 3490 1365 3570 1405
rect 3370 1280 3570 1365
rect 3720 1405 3920 1480
rect 3720 1365 3800 1405
rect 3840 1365 3920 1405
rect 3720 1280 3920 1365
rect 4070 1405 4270 1480
rect 4070 1365 4150 1405
rect 4190 1365 4270 1405
rect 4070 1280 4270 1365
rect 4420 1405 4620 1480
rect 4420 1365 4500 1405
rect 4540 1365 4620 1405
rect 4420 1280 4620 1365
rect 4770 1405 4970 1480
rect 4770 1365 4850 1405
rect 4890 1365 4970 1405
rect 4770 1280 4970 1365
rect -3280 1055 -3080 1130
rect -3280 1015 -3200 1055
rect -3160 1015 -3080 1055
rect -3280 930 -3080 1015
rect -2930 1055 -2730 1130
rect -2930 1015 -2850 1055
rect -2810 1015 -2730 1055
rect -2930 930 -2730 1015
rect -2580 1055 -2380 1130
rect -2580 1015 -2500 1055
rect -2460 1015 -2380 1055
rect -2580 930 -2380 1015
rect -2230 1055 -2030 1130
rect -2230 1015 -2150 1055
rect -2110 1015 -2030 1055
rect -2230 930 -2030 1015
rect -1880 1055 -1680 1130
rect -1880 1015 -1800 1055
rect -1760 1015 -1680 1055
rect -1880 930 -1680 1015
rect 3370 1055 3570 1130
rect 3370 1015 3450 1055
rect 3490 1015 3570 1055
rect 3370 930 3570 1015
rect 3720 1055 3920 1130
rect 3720 1015 3800 1055
rect 3840 1015 3920 1055
rect 3720 930 3920 1015
rect 4070 1055 4270 1130
rect 4070 1015 4150 1055
rect 4190 1015 4270 1055
rect 4070 930 4270 1015
rect 4420 1055 4620 1130
rect 4420 1015 4500 1055
rect 4540 1015 4620 1055
rect 4420 930 4620 1015
rect 4770 1055 4970 1130
rect 4770 1015 4850 1055
rect 4890 1015 4970 1055
rect 4770 930 4970 1015
rect -3280 705 -3080 780
rect -3280 665 -3200 705
rect -3160 665 -3080 705
rect -3280 580 -3080 665
rect -2930 705 -2730 780
rect -2930 665 -2850 705
rect -2810 665 -2730 705
rect -2930 580 -2730 665
rect -2580 705 -2380 780
rect -2580 665 -2500 705
rect -2460 665 -2380 705
rect -2580 580 -2380 665
rect -2230 705 -2030 780
rect -2230 665 -2150 705
rect -2110 665 -2030 705
rect -2230 580 -2030 665
rect -1880 705 -1680 780
rect -1880 665 -1800 705
rect -1760 665 -1680 705
rect -1880 580 -1680 665
rect 3370 705 3570 780
rect 3370 665 3450 705
rect 3490 665 3570 705
rect 3370 580 3570 665
rect 3720 705 3920 780
rect 3720 665 3800 705
rect 3840 665 3920 705
rect 3720 580 3920 665
rect 4070 705 4270 780
rect 4070 665 4150 705
rect 4190 665 4270 705
rect 4070 580 4270 665
rect 4420 705 4620 780
rect 4420 665 4500 705
rect 4540 665 4620 705
rect 4420 580 4620 665
rect 4770 705 4970 780
rect 4770 665 4850 705
rect 4890 665 4970 705
rect 4770 580 4970 665
rect -3280 355 -3080 430
rect -3280 315 -3200 355
rect -3160 315 -3080 355
rect -3280 230 -3080 315
rect -2930 355 -2730 430
rect -2930 315 -2850 355
rect -2810 315 -2730 355
rect -2930 230 -2730 315
rect -2580 355 -2380 430
rect -2580 315 -2500 355
rect -2460 315 -2380 355
rect -2580 230 -2380 315
rect -2230 355 -2030 430
rect -2230 315 -2150 355
rect -2110 315 -2030 355
rect -2230 230 -2030 315
rect -1880 355 -1680 430
rect -1880 315 -1800 355
rect -1760 315 -1680 355
rect -1880 230 -1680 315
rect 3370 355 3570 430
rect 3370 315 3450 355
rect 3490 315 3570 355
rect 3370 230 3570 315
rect 3720 355 3920 430
rect 3720 315 3800 355
rect 3840 315 3920 355
rect 3720 230 3920 315
rect 4070 355 4270 430
rect 4070 315 4150 355
rect 4190 315 4270 355
rect 4070 230 4270 315
rect 4420 355 4620 430
rect 4420 315 4500 355
rect 4540 315 4620 355
rect 4420 230 4620 315
rect 4770 355 4970 430
rect 4770 315 4850 355
rect 4890 315 4970 355
rect 4770 230 4970 315
rect -3280 5 -3080 80
rect -3280 -35 -3200 5
rect -3160 -35 -3080 5
rect -3280 -120 -3080 -35
rect -2930 5 -2730 80
rect -2930 -35 -2850 5
rect -2810 -35 -2730 5
rect -2930 -120 -2730 -35
rect -2580 5 -2380 80
rect -2580 -35 -2500 5
rect -2460 -35 -2380 5
rect -2580 -120 -2380 -35
rect -2230 5 -2030 80
rect -2230 -35 -2150 5
rect -2110 -35 -2030 5
rect -2230 -120 -2030 -35
rect -1880 5 -1680 80
rect -1880 -35 -1800 5
rect -1760 -35 -1680 5
rect -1880 -120 -1680 -35
rect 3370 5 3570 80
rect 3370 -35 3450 5
rect 3490 -35 3570 5
rect 3370 -120 3570 -35
rect 3720 5 3920 80
rect 3720 -35 3800 5
rect 3840 -35 3920 5
rect 3720 -120 3920 -35
rect 4070 5 4270 80
rect 4070 -35 4150 5
rect 4190 -35 4270 5
rect 4070 -120 4270 -35
rect 4420 5 4620 80
rect 4420 -35 4500 5
rect 4540 -35 4620 5
rect 4420 -120 4620 -35
rect 4770 5 4970 80
rect 4770 -35 4850 5
rect 4890 -35 4970 5
rect 4770 -120 4970 -35
rect -3280 -345 -3080 -270
rect -3280 -385 -3200 -345
rect -3160 -385 -3080 -345
rect -3280 -470 -3080 -385
rect -2930 -345 -2730 -270
rect -2930 -385 -2850 -345
rect -2810 -385 -2730 -345
rect -2930 -470 -2730 -385
rect -2580 -345 -2380 -270
rect -2580 -385 -2500 -345
rect -2460 -385 -2380 -345
rect -2580 -470 -2380 -385
rect -2230 -345 -2030 -270
rect -2230 -385 -2150 -345
rect -2110 -385 -2030 -345
rect -2230 -470 -2030 -385
rect -1880 -345 -1680 -270
rect -1880 -385 -1800 -345
rect -1760 -385 -1680 -345
rect -1880 -470 -1680 -385
rect 3370 -345 3570 -270
rect 3370 -385 3450 -345
rect 3490 -385 3570 -345
rect 3370 -470 3570 -385
rect 3720 -345 3920 -270
rect 3720 -385 3800 -345
rect 3840 -385 3920 -345
rect 3720 -470 3920 -385
rect 4070 -345 4270 -270
rect 4070 -385 4150 -345
rect 4190 -385 4270 -345
rect 4070 -470 4270 -385
rect 4420 -345 4620 -270
rect 4420 -385 4500 -345
rect 4540 -385 4620 -345
rect 4420 -470 4620 -385
rect 4770 -345 4970 -270
rect 4770 -385 4850 -345
rect 4890 -385 4970 -345
rect 4770 -470 4970 -385
rect -3280 -695 -3080 -620
rect -3280 -735 -3200 -695
rect -3160 -735 -3080 -695
rect -3280 -820 -3080 -735
rect -2930 -695 -2730 -620
rect -2930 -735 -2850 -695
rect -2810 -735 -2730 -695
rect -2930 -820 -2730 -735
rect -2580 -695 -2380 -620
rect -2580 -735 -2500 -695
rect -2460 -735 -2380 -695
rect -2580 -820 -2380 -735
rect -2230 -695 -2030 -620
rect -2230 -735 -2150 -695
rect -2110 -735 -2030 -695
rect -2230 -820 -2030 -735
rect -1880 -695 -1680 -620
rect -1880 -735 -1800 -695
rect -1760 -735 -1680 -695
rect -1880 -820 -1680 -735
rect 3370 -695 3570 -620
rect 3370 -735 3450 -695
rect 3490 -735 3570 -695
rect 3370 -820 3570 -735
rect 3720 -695 3920 -620
rect 3720 -735 3800 -695
rect 3840 -735 3920 -695
rect 3720 -820 3920 -735
rect 4070 -695 4270 -620
rect 4070 -735 4150 -695
rect 4190 -735 4270 -695
rect 4070 -820 4270 -735
rect 4420 -695 4620 -620
rect 4420 -735 4500 -695
rect 4540 -735 4620 -695
rect 4420 -820 4620 -735
rect 4770 -695 4970 -620
rect 4770 -735 4850 -695
rect 4890 -735 4970 -695
rect 4770 -820 4970 -735
rect -3280 -1045 -3080 -970
rect -3280 -1085 -3200 -1045
rect -3160 -1085 -3080 -1045
rect -3280 -1170 -3080 -1085
rect -2930 -1045 -2730 -970
rect -2930 -1085 -2850 -1045
rect -2810 -1085 -2730 -1045
rect -2930 -1170 -2730 -1085
rect -2580 -1045 -2380 -970
rect -2580 -1085 -2500 -1045
rect -2460 -1085 -2380 -1045
rect -2580 -1170 -2380 -1085
rect -2230 -1045 -2030 -970
rect -2230 -1085 -2150 -1045
rect -2110 -1085 -2030 -1045
rect -2230 -1170 -2030 -1085
rect -1880 -1045 -1680 -970
rect -1880 -1085 -1800 -1045
rect -1760 -1085 -1680 -1045
rect -1880 -1170 -1680 -1085
rect 3370 -1045 3570 -970
rect 3370 -1085 3450 -1045
rect 3490 -1085 3570 -1045
rect 3370 -1170 3570 -1085
rect 3720 -1045 3920 -970
rect 3720 -1085 3800 -1045
rect 3840 -1085 3920 -1045
rect 3720 -1170 3920 -1085
rect 4070 -1045 4270 -970
rect 4070 -1085 4150 -1045
rect 4190 -1085 4270 -1045
rect 4070 -1170 4270 -1085
rect 4420 -1045 4620 -970
rect 4420 -1085 4500 -1045
rect 4540 -1085 4620 -1045
rect 4420 -1170 4620 -1085
rect 4770 -1045 4970 -970
rect 4770 -1085 4850 -1045
rect 4890 -1085 4970 -1045
rect 4770 -1170 4970 -1085
rect -3280 -1395 -3080 -1320
rect -3280 -1435 -3200 -1395
rect -3160 -1435 -3080 -1395
rect -3280 -1520 -3080 -1435
rect -2930 -1395 -2730 -1320
rect -2930 -1435 -2850 -1395
rect -2810 -1435 -2730 -1395
rect -2930 -1520 -2730 -1435
rect -2580 -1395 -2380 -1320
rect -2580 -1435 -2500 -1395
rect -2460 -1435 -2380 -1395
rect -2580 -1520 -2380 -1435
rect -2230 -1395 -2030 -1320
rect -2230 -1435 -2150 -1395
rect -2110 -1435 -2030 -1395
rect -2230 -1520 -2030 -1435
rect -1880 -1395 -1680 -1320
rect -1880 -1435 -1800 -1395
rect -1760 -1435 -1680 -1395
rect -1880 -1520 -1680 -1435
rect -1530 -1395 -1330 -1320
rect -1530 -1435 -1450 -1395
rect -1410 -1435 -1330 -1395
rect -1530 -1520 -1330 -1435
rect -1180 -1395 -980 -1320
rect -1180 -1435 -1100 -1395
rect -1060 -1435 -980 -1395
rect -1180 -1520 -980 -1435
rect -830 -1395 -630 -1320
rect -830 -1435 -750 -1395
rect -710 -1435 -630 -1395
rect -830 -1520 -630 -1435
rect -480 -1395 -280 -1320
rect -480 -1435 -400 -1395
rect -360 -1435 -280 -1395
rect -480 -1520 -280 -1435
rect -130 -1395 70 -1320
rect -130 -1435 -50 -1395
rect -10 -1435 70 -1395
rect -130 -1520 70 -1435
rect 220 -1395 420 -1320
rect 220 -1435 300 -1395
rect 340 -1435 420 -1395
rect 220 -1520 420 -1435
rect 570 -1395 770 -1320
rect 570 -1435 650 -1395
rect 690 -1435 770 -1395
rect 570 -1520 770 -1435
rect 920 -1395 1120 -1320
rect 920 -1435 1000 -1395
rect 1040 -1435 1120 -1395
rect 920 -1520 1120 -1435
rect 1270 -1395 1470 -1320
rect 1270 -1435 1350 -1395
rect 1390 -1435 1470 -1395
rect 1270 -1520 1470 -1435
rect 1620 -1395 1820 -1320
rect 1620 -1435 1700 -1395
rect 1740 -1435 1820 -1395
rect 1620 -1520 1820 -1435
rect 1970 -1395 2170 -1320
rect 1970 -1435 2050 -1395
rect 2090 -1435 2170 -1395
rect 1970 -1520 2170 -1435
rect 2320 -1395 2520 -1320
rect 2320 -1435 2400 -1395
rect 2440 -1435 2520 -1395
rect 2320 -1520 2520 -1435
rect 2670 -1395 2870 -1320
rect 2670 -1435 2750 -1395
rect 2790 -1435 2870 -1395
rect 2670 -1520 2870 -1435
rect 3020 -1395 3220 -1320
rect 3020 -1435 3100 -1395
rect 3140 -1435 3220 -1395
rect 3020 -1520 3220 -1435
rect 3370 -1395 3570 -1320
rect 3370 -1435 3450 -1395
rect 3490 -1435 3570 -1395
rect 3370 -1520 3570 -1435
rect 3720 -1395 3920 -1320
rect 3720 -1435 3800 -1395
rect 3840 -1435 3920 -1395
rect 3720 -1520 3920 -1435
rect 4070 -1395 4270 -1320
rect 4070 -1435 4150 -1395
rect 4190 -1435 4270 -1395
rect 4070 -1520 4270 -1435
rect 4420 -1395 4620 -1320
rect 4420 -1435 4500 -1395
rect 4540 -1435 4620 -1395
rect 4420 -1520 4620 -1435
rect 4770 -1395 4970 -1320
rect 4770 -1435 4850 -1395
rect 4890 -1435 4970 -1395
rect 4770 -1520 4970 -1435
rect -3280 -1745 -3080 -1670
rect -3280 -1785 -3200 -1745
rect -3160 -1785 -3080 -1745
rect -3280 -1870 -3080 -1785
rect -2930 -1745 -2730 -1670
rect -2930 -1785 -2850 -1745
rect -2810 -1785 -2730 -1745
rect -2930 -1870 -2730 -1785
rect -2580 -1745 -2380 -1670
rect -2580 -1785 -2500 -1745
rect -2460 -1785 -2380 -1745
rect -2580 -1870 -2380 -1785
rect -2230 -1745 -2030 -1670
rect -2230 -1785 -2150 -1745
rect -2110 -1785 -2030 -1745
rect -2230 -1870 -2030 -1785
rect -1880 -1745 -1680 -1670
rect -1880 -1785 -1800 -1745
rect -1760 -1785 -1680 -1745
rect -1880 -1870 -1680 -1785
rect -1530 -1745 -1330 -1670
rect -1530 -1785 -1450 -1745
rect -1410 -1785 -1330 -1745
rect -1530 -1870 -1330 -1785
rect -1180 -1745 -980 -1670
rect -1180 -1785 -1100 -1745
rect -1060 -1785 -980 -1745
rect -1180 -1870 -980 -1785
rect -830 -1745 -630 -1670
rect -830 -1785 -750 -1745
rect -710 -1785 -630 -1745
rect -830 -1870 -630 -1785
rect -480 -1745 -280 -1670
rect -480 -1785 -400 -1745
rect -360 -1785 -280 -1745
rect -480 -1870 -280 -1785
rect -130 -1745 70 -1670
rect -130 -1785 -50 -1745
rect -10 -1785 70 -1745
rect -130 -1870 70 -1785
rect 220 -1745 420 -1670
rect 220 -1785 300 -1745
rect 340 -1785 420 -1745
rect 220 -1870 420 -1785
rect 570 -1745 770 -1670
rect 570 -1785 650 -1745
rect 690 -1785 770 -1745
rect 570 -1870 770 -1785
rect 920 -1745 1120 -1670
rect 920 -1785 1000 -1745
rect 1040 -1785 1120 -1745
rect 920 -1870 1120 -1785
rect 1270 -1745 1470 -1670
rect 1270 -1785 1350 -1745
rect 1390 -1785 1470 -1745
rect 1270 -1870 1470 -1785
rect 1620 -1745 1820 -1670
rect 1620 -1785 1700 -1745
rect 1740 -1785 1820 -1745
rect 1620 -1870 1820 -1785
rect 1970 -1745 2170 -1670
rect 1970 -1785 2050 -1745
rect 2090 -1785 2170 -1745
rect 1970 -1870 2170 -1785
rect 2320 -1745 2520 -1670
rect 2320 -1785 2400 -1745
rect 2440 -1785 2520 -1745
rect 2320 -1870 2520 -1785
rect 2670 -1745 2870 -1670
rect 2670 -1785 2750 -1745
rect 2790 -1785 2870 -1745
rect 2670 -1870 2870 -1785
rect 3020 -1745 3220 -1670
rect 3020 -1785 3100 -1745
rect 3140 -1785 3220 -1745
rect 3020 -1870 3220 -1785
rect 3370 -1745 3570 -1670
rect 3370 -1785 3450 -1745
rect 3490 -1785 3570 -1745
rect 3370 -1870 3570 -1785
rect 3720 -1745 3920 -1670
rect 3720 -1785 3800 -1745
rect 3840 -1785 3920 -1745
rect 3720 -1870 3920 -1785
rect 4070 -1745 4270 -1670
rect 4070 -1785 4150 -1745
rect 4190 -1785 4270 -1745
rect 4070 -1870 4270 -1785
rect 4420 -1745 4620 -1670
rect 4420 -1785 4500 -1745
rect 4540 -1785 4620 -1745
rect 4420 -1870 4620 -1785
rect 4770 -1745 4970 -1670
rect 4770 -1785 4850 -1745
rect 4890 -1785 4970 -1745
rect 4770 -1870 4970 -1785
rect -3280 -2095 -3080 -2020
rect -3280 -2135 -3200 -2095
rect -3160 -2135 -3080 -2095
rect -3280 -2220 -3080 -2135
rect -2930 -2095 -2730 -2020
rect -2930 -2135 -2850 -2095
rect -2810 -2135 -2730 -2095
rect -2930 -2220 -2730 -2135
rect -2580 -2095 -2380 -2020
rect -2580 -2135 -2500 -2095
rect -2460 -2135 -2380 -2095
rect -2580 -2220 -2380 -2135
rect -2230 -2095 -2030 -2020
rect -2230 -2135 -2150 -2095
rect -2110 -2135 -2030 -2095
rect -2230 -2220 -2030 -2135
rect -1880 -2095 -1680 -2020
rect -1880 -2135 -1800 -2095
rect -1760 -2135 -1680 -2095
rect -1880 -2220 -1680 -2135
rect -1530 -2095 -1330 -2020
rect -1530 -2135 -1450 -2095
rect -1410 -2135 -1330 -2095
rect -1530 -2220 -1330 -2135
rect -1180 -2095 -980 -2020
rect -1180 -2135 -1100 -2095
rect -1060 -2135 -980 -2095
rect -1180 -2220 -980 -2135
rect -830 -2095 -630 -2020
rect -830 -2135 -750 -2095
rect -710 -2135 -630 -2095
rect -830 -2220 -630 -2135
rect -480 -2095 -280 -2020
rect -480 -2135 -400 -2095
rect -360 -2135 -280 -2095
rect -480 -2220 -280 -2135
rect -130 -2095 70 -2020
rect -130 -2135 -50 -2095
rect -10 -2135 70 -2095
rect -130 -2220 70 -2135
rect 220 -2095 420 -2020
rect 220 -2135 300 -2095
rect 340 -2135 420 -2095
rect 220 -2220 420 -2135
rect 570 -2095 770 -2020
rect 570 -2135 650 -2095
rect 690 -2135 770 -2095
rect 570 -2220 770 -2135
rect 920 -2095 1120 -2020
rect 920 -2135 1000 -2095
rect 1040 -2135 1120 -2095
rect 920 -2220 1120 -2135
rect 1270 -2095 1470 -2020
rect 1270 -2135 1350 -2095
rect 1390 -2135 1470 -2095
rect 1270 -2220 1470 -2135
rect 1620 -2095 1820 -2020
rect 1620 -2135 1700 -2095
rect 1740 -2135 1820 -2095
rect 1620 -2220 1820 -2135
rect 1970 -2095 2170 -2020
rect 1970 -2135 2050 -2095
rect 2090 -2135 2170 -2095
rect 1970 -2220 2170 -2135
rect 2320 -2095 2520 -2020
rect 2320 -2135 2400 -2095
rect 2440 -2135 2520 -2095
rect 2320 -2220 2520 -2135
rect 2670 -2095 2870 -2020
rect 2670 -2135 2750 -2095
rect 2790 -2135 2870 -2095
rect 2670 -2220 2870 -2135
rect 3020 -2095 3220 -2020
rect 3020 -2135 3100 -2095
rect 3140 -2135 3220 -2095
rect 3020 -2220 3220 -2135
rect 3370 -2095 3570 -2020
rect 3370 -2135 3450 -2095
rect 3490 -2135 3570 -2095
rect 3370 -2220 3570 -2135
rect 3720 -2095 3920 -2020
rect 3720 -2135 3800 -2095
rect 3840 -2135 3920 -2095
rect 3720 -2220 3920 -2135
rect 4070 -2095 4270 -2020
rect 4070 -2135 4150 -2095
rect 4190 -2135 4270 -2095
rect 4070 -2220 4270 -2135
rect 4420 -2095 4620 -2020
rect 4420 -2135 4500 -2095
rect 4540 -2135 4620 -2095
rect 4420 -2220 4620 -2135
rect 4770 -2095 4970 -2020
rect 4770 -2135 4850 -2095
rect 4890 -2135 4970 -2095
rect 4770 -2220 4970 -2135
<< mimcapcontact >>
rect -3200 3815 -3160 3855
rect -2850 3815 -2810 3855
rect -2500 3815 -2460 3855
rect -2150 3815 -2110 3855
rect -1800 3815 -1760 3855
rect -1450 3815 -1410 3855
rect -1100 3815 -1060 3855
rect -750 3815 -710 3855
rect -400 3815 -360 3855
rect -50 3815 -10 3855
rect 300 3815 340 3855
rect 650 3815 690 3855
rect 1000 3815 1040 3855
rect 1350 3815 1390 3855
rect 1700 3815 1740 3855
rect 2050 3815 2090 3855
rect 2400 3815 2440 3855
rect 2750 3815 2790 3855
rect 3100 3815 3140 3855
rect 3450 3815 3490 3855
rect 3800 3815 3840 3855
rect 4150 3815 4190 3855
rect 4500 3815 4540 3855
rect 4850 3815 4890 3855
rect -3200 3465 -3160 3505
rect -2850 3465 -2810 3505
rect -2500 3465 -2460 3505
rect -2150 3465 -2110 3505
rect -1800 3465 -1760 3505
rect -1450 3465 -1410 3505
rect -1100 3465 -1060 3505
rect -750 3465 -710 3505
rect -400 3465 -360 3505
rect -50 3465 -10 3505
rect 300 3465 340 3505
rect 650 3465 690 3505
rect 1000 3465 1040 3505
rect 1350 3465 1390 3505
rect 1700 3465 1740 3505
rect 2050 3465 2090 3505
rect 2400 3465 2440 3505
rect 2750 3465 2790 3505
rect 3100 3465 3140 3505
rect 3450 3465 3490 3505
rect 3800 3465 3840 3505
rect 4150 3465 4190 3505
rect 4500 3465 4540 3505
rect 4850 3465 4890 3505
rect -3200 3115 -3160 3155
rect -2850 3115 -2810 3155
rect -2500 3115 -2460 3155
rect -2150 3115 -2110 3155
rect -1800 3115 -1760 3155
rect -1450 3115 -1410 3155
rect -1100 3115 -1060 3155
rect -750 3115 -710 3155
rect -400 3115 -360 3155
rect -50 3105 -10 3145
rect 300 3105 340 3145
rect 650 3105 690 3145
rect 1000 3105 1040 3145
rect 1350 3105 1390 3145
rect 1700 3105 1740 3145
rect 2050 3115 2090 3155
rect 2400 3115 2440 3155
rect 2750 3115 2790 3155
rect 3100 3115 3140 3155
rect 3450 3115 3490 3155
rect 3800 3115 3840 3155
rect 4150 3115 4190 3155
rect 4500 3115 4540 3155
rect 4850 3115 4890 3155
rect -3200 2765 -3160 2805
rect -2850 2765 -2810 2805
rect -2500 2765 -2460 2805
rect -2150 2765 -2110 2805
rect -1800 2765 -1760 2805
rect -1450 2765 -1410 2805
rect -1100 2765 -1060 2805
rect -750 2765 -710 2805
rect 2400 2765 2440 2805
rect 2750 2765 2790 2805
rect 3100 2765 3140 2805
rect 3450 2765 3490 2805
rect 3800 2765 3840 2805
rect 4150 2765 4190 2805
rect 4500 2765 4540 2805
rect 4850 2765 4890 2805
rect -3200 2415 -3160 2455
rect -2850 2415 -2810 2455
rect -2500 2415 -2460 2455
rect -2150 2415 -2110 2455
rect -1800 2415 -1760 2455
rect -1450 2415 -1410 2455
rect -1100 2415 -1060 2455
rect -750 2415 -710 2455
rect 2400 2415 2440 2455
rect 2750 2415 2790 2455
rect 3100 2415 3140 2455
rect 3450 2415 3490 2455
rect 3800 2415 3840 2455
rect 4150 2415 4190 2455
rect 4500 2415 4540 2455
rect 4850 2415 4890 2455
rect -3200 2065 -3160 2105
rect -2850 2065 -2810 2105
rect -2500 2065 -2460 2105
rect -2150 2065 -2110 2105
rect -1800 2065 -1760 2105
rect 3450 2065 3490 2105
rect 3800 2065 3840 2105
rect 4150 2065 4190 2105
rect 4500 2065 4540 2105
rect 4850 2065 4890 2105
rect -3200 1715 -3160 1755
rect -2850 1715 -2810 1755
rect -2500 1715 -2460 1755
rect -2150 1715 -2110 1755
rect -1800 1715 -1760 1755
rect 3450 1715 3490 1755
rect 3800 1715 3840 1755
rect 4150 1715 4190 1755
rect 4500 1715 4540 1755
rect 4850 1715 4890 1755
rect -3200 1365 -3160 1405
rect -2850 1365 -2810 1405
rect -2500 1365 -2460 1405
rect -2150 1365 -2110 1405
rect -1800 1365 -1760 1405
rect 3450 1365 3490 1405
rect 3800 1365 3840 1405
rect 4150 1365 4190 1405
rect 4500 1365 4540 1405
rect 4850 1365 4890 1405
rect -3200 1015 -3160 1055
rect -2850 1015 -2810 1055
rect -2500 1015 -2460 1055
rect -2150 1015 -2110 1055
rect -1800 1015 -1760 1055
rect 3450 1015 3490 1055
rect 3800 1015 3840 1055
rect 4150 1015 4190 1055
rect 4500 1015 4540 1055
rect 4850 1015 4890 1055
rect -3200 665 -3160 705
rect -2850 665 -2810 705
rect -2500 665 -2460 705
rect -2150 665 -2110 705
rect -1800 665 -1760 705
rect 3450 665 3490 705
rect 3800 665 3840 705
rect 4150 665 4190 705
rect 4500 665 4540 705
rect 4850 665 4890 705
rect -3200 315 -3160 355
rect -2850 315 -2810 355
rect -2500 315 -2460 355
rect -2150 315 -2110 355
rect -1800 315 -1760 355
rect 3450 315 3490 355
rect 3800 315 3840 355
rect 4150 315 4190 355
rect 4500 315 4540 355
rect 4850 315 4890 355
rect -3200 -35 -3160 5
rect -2850 -35 -2810 5
rect -2500 -35 -2460 5
rect -2150 -35 -2110 5
rect -1800 -35 -1760 5
rect 3450 -35 3490 5
rect 3800 -35 3840 5
rect 4150 -35 4190 5
rect 4500 -35 4540 5
rect 4850 -35 4890 5
rect -3200 -385 -3160 -345
rect -2850 -385 -2810 -345
rect -2500 -385 -2460 -345
rect -2150 -385 -2110 -345
rect -1800 -385 -1760 -345
rect 3450 -385 3490 -345
rect 3800 -385 3840 -345
rect 4150 -385 4190 -345
rect 4500 -385 4540 -345
rect 4850 -385 4890 -345
rect -3200 -735 -3160 -695
rect -2850 -735 -2810 -695
rect -2500 -735 -2460 -695
rect -2150 -735 -2110 -695
rect -1800 -735 -1760 -695
rect 3450 -735 3490 -695
rect 3800 -735 3840 -695
rect 4150 -735 4190 -695
rect 4500 -735 4540 -695
rect 4850 -735 4890 -695
rect -3200 -1085 -3160 -1045
rect -2850 -1085 -2810 -1045
rect -2500 -1085 -2460 -1045
rect -2150 -1085 -2110 -1045
rect -1800 -1085 -1760 -1045
rect 3450 -1085 3490 -1045
rect 3800 -1085 3840 -1045
rect 4150 -1085 4190 -1045
rect 4500 -1085 4540 -1045
rect 4850 -1085 4890 -1045
rect -3200 -1435 -3160 -1395
rect -2850 -1435 -2810 -1395
rect -2500 -1435 -2460 -1395
rect -2150 -1435 -2110 -1395
rect -1800 -1435 -1760 -1395
rect -1450 -1435 -1410 -1395
rect -1100 -1435 -1060 -1395
rect -750 -1435 -710 -1395
rect -400 -1435 -360 -1395
rect -50 -1435 -10 -1395
rect 300 -1435 340 -1395
rect 650 -1435 690 -1395
rect 1000 -1435 1040 -1395
rect 1350 -1435 1390 -1395
rect 1700 -1435 1740 -1395
rect 2050 -1435 2090 -1395
rect 2400 -1435 2440 -1395
rect 2750 -1435 2790 -1395
rect 3100 -1435 3140 -1395
rect 3450 -1435 3490 -1395
rect 3800 -1435 3840 -1395
rect 4150 -1435 4190 -1395
rect 4500 -1435 4540 -1395
rect 4850 -1435 4890 -1395
rect -3200 -1785 -3160 -1745
rect -2850 -1785 -2810 -1745
rect -2500 -1785 -2460 -1745
rect -2150 -1785 -2110 -1745
rect -1800 -1785 -1760 -1745
rect -1450 -1785 -1410 -1745
rect -1100 -1785 -1060 -1745
rect -750 -1785 -710 -1745
rect -400 -1785 -360 -1745
rect -50 -1785 -10 -1745
rect 300 -1785 340 -1745
rect 650 -1785 690 -1745
rect 1000 -1785 1040 -1745
rect 1350 -1785 1390 -1745
rect 1700 -1785 1740 -1745
rect 2050 -1785 2090 -1745
rect 2400 -1785 2440 -1745
rect 2750 -1785 2790 -1745
rect 3100 -1785 3140 -1745
rect 3450 -1785 3490 -1745
rect 3800 -1785 3840 -1745
rect 4150 -1785 4190 -1745
rect 4500 -1785 4540 -1745
rect 4850 -1785 4890 -1745
rect -3200 -2135 -3160 -2095
rect -2850 -2135 -2810 -2095
rect -2500 -2135 -2460 -2095
rect -2150 -2135 -2110 -2095
rect -1800 -2135 -1760 -2095
rect -1450 -2135 -1410 -2095
rect -1100 -2135 -1060 -2095
rect -750 -2135 -710 -2095
rect -400 -2135 -360 -2095
rect -50 -2135 -10 -2095
rect 300 -2135 340 -2095
rect 650 -2135 690 -2095
rect 1000 -2135 1040 -2095
rect 1350 -2135 1390 -2095
rect 1700 -2135 1740 -2095
rect 2050 -2135 2090 -2095
rect 2400 -2135 2440 -2095
rect 2750 -2135 2790 -2095
rect 3100 -2135 3140 -2095
rect 3450 -2135 3490 -2095
rect 3800 -2135 3840 -2095
rect 4150 -2135 4190 -2095
rect 4500 -2135 4540 -2095
rect 4850 -2135 4890 -2095
<< metal4 >>
rect -3850 4280 5140 4285
rect -3850 4240 825 4280
rect 865 4240 5140 4280
rect -3850 4235 5140 4240
rect -3205 3855 -2455 3860
rect -3205 3815 -3200 3855
rect -3160 3815 -2850 3855
rect -2810 3815 -2500 3855
rect -2460 3815 -2455 3855
rect -3205 3810 -2455 3815
rect -2505 3510 -2455 3810
rect -2155 3855 -2105 3860
rect -2155 3815 -2150 3855
rect -2110 3815 -2105 3855
rect -2155 3510 -2105 3815
rect -1805 3855 -1755 3860
rect -1805 3815 -1800 3855
rect -1760 3815 -1755 3855
rect -1805 3510 -1755 3815
rect -1455 3855 -1405 3860
rect -1455 3815 -1450 3855
rect -1410 3815 -1405 3855
rect -1455 3510 -1405 3815
rect -1105 3855 -1055 3860
rect -1105 3815 -1100 3855
rect -1060 3815 -1055 3855
rect -1105 3510 -1055 3815
rect -755 3855 -705 3860
rect -755 3815 -750 3855
rect -710 3815 -705 3855
rect -755 3510 -705 3815
rect -405 3855 -355 3860
rect -405 3815 -400 3855
rect -360 3815 -355 3855
rect -405 3510 -355 3815
rect -55 3855 -5 3860
rect -55 3815 -50 3855
rect -10 3815 -5 3855
rect -55 3510 -5 3815
rect 295 3855 345 3860
rect 295 3815 300 3855
rect 340 3815 345 3855
rect 295 3510 345 3815
rect 645 3855 695 3860
rect 645 3815 650 3855
rect 690 3815 695 3855
rect 645 3510 695 3815
rect -3205 3505 695 3510
rect -3205 3465 -3200 3505
rect -3160 3465 -2850 3505
rect -2810 3465 -2500 3505
rect -2460 3465 -2150 3505
rect -2110 3465 -1800 3505
rect -1760 3465 -1450 3505
rect -1410 3465 -1100 3505
rect -1060 3465 -750 3505
rect -710 3465 -400 3505
rect -360 3465 -50 3505
rect -10 3465 300 3505
rect 340 3465 650 3505
rect 690 3465 695 3505
rect -3205 3460 695 3465
rect -2505 3160 -2455 3460
rect -3205 3155 -2105 3160
rect -3205 3115 -3200 3155
rect -3160 3115 -2850 3155
rect -2810 3115 -2500 3155
rect -2460 3115 -2150 3155
rect -2110 3115 -2105 3155
rect -3205 3110 -2105 3115
rect -1805 3155 -1755 3460
rect -1805 3115 -1800 3155
rect -1760 3115 -1755 3155
rect -2505 2810 -2455 3110
rect -3205 2805 -2105 2810
rect -3205 2765 -3200 2805
rect -3160 2765 -2850 2805
rect -2810 2765 -2500 2805
rect -2460 2765 -2150 2805
rect -2110 2765 -2105 2805
rect -3205 2760 -2105 2765
rect -1805 2805 -1755 3115
rect -1805 2765 -1800 2805
rect -1760 2765 -1755 2805
rect -1805 2760 -1755 2765
rect -1455 3155 -1405 3460
rect -1455 3115 -1450 3155
rect -1410 3115 -1405 3155
rect -1455 2805 -1405 3115
rect -1455 2765 -1450 2805
rect -1410 2765 -1405 2805
rect -2505 2460 -2455 2760
rect -3205 2455 -1755 2460
rect -3205 2415 -3200 2455
rect -3160 2415 -2850 2455
rect -2810 2415 -2500 2455
rect -2460 2415 -2150 2455
rect -2110 2415 -1800 2455
rect -1760 2415 -1755 2455
rect -3205 2410 -1755 2415
rect -1455 2455 -1405 2765
rect -1455 2415 -1450 2455
rect -1410 2415 -1405 2455
rect -1455 2410 -1405 2415
rect -1105 3155 -1055 3460
rect -1105 3115 -1100 3155
rect -1060 3115 -1055 3155
rect -1105 2805 -1055 3115
rect -1105 2765 -1100 2805
rect -1060 2765 -1055 2805
rect -1105 2455 -1055 2765
rect -1105 2415 -1100 2455
rect -1060 2415 -1055 2455
rect -1105 2410 -1055 2415
rect -755 3155 -705 3460
rect -755 3115 -750 3155
rect -710 3115 -705 3155
rect -755 2805 -705 3115
rect -405 3155 -355 3460
rect -405 3115 -400 3155
rect -360 3115 -355 3155
rect -405 3110 -355 3115
rect -55 3145 -5 3460
rect -55 3105 -50 3145
rect -10 3105 -5 3145
rect -55 3100 -5 3105
rect 295 3145 345 3460
rect 295 3105 300 3145
rect 340 3105 345 3145
rect 295 3100 345 3105
rect 645 3145 695 3460
rect 645 3105 650 3145
rect 690 3105 695 3145
rect 645 3100 695 3105
rect 995 3855 1045 3860
rect 995 3815 1000 3855
rect 1040 3815 1045 3855
rect 995 3510 1045 3815
rect 1345 3855 1395 3860
rect 1345 3815 1350 3855
rect 1390 3815 1395 3855
rect 1345 3510 1395 3815
rect 1695 3855 1745 3860
rect 1695 3815 1700 3855
rect 1740 3815 1745 3855
rect 1695 3510 1745 3815
rect 2045 3855 2095 3860
rect 2045 3815 2050 3855
rect 2090 3815 2095 3855
rect 2045 3510 2095 3815
rect 2395 3855 2445 3860
rect 2395 3815 2400 3855
rect 2440 3815 2445 3855
rect 2395 3510 2445 3815
rect 2745 3855 2795 3860
rect 2745 3815 2750 3855
rect 2790 3815 2795 3855
rect 2745 3510 2795 3815
rect 3095 3855 3145 3860
rect 3095 3815 3100 3855
rect 3140 3815 3145 3855
rect 3095 3510 3145 3815
rect 3445 3855 3495 3860
rect 3445 3815 3450 3855
rect 3490 3815 3495 3855
rect 3445 3510 3495 3815
rect 3795 3855 3845 3860
rect 3795 3815 3800 3855
rect 3840 3815 3845 3855
rect 3795 3510 3845 3815
rect 4145 3855 4895 3860
rect 4145 3815 4150 3855
rect 4190 3815 4500 3855
rect 4540 3815 4850 3855
rect 4890 3815 4895 3855
rect 4145 3810 4895 3815
rect 4145 3510 4195 3810
rect 995 3505 4895 3510
rect 995 3465 1000 3505
rect 1040 3465 1350 3505
rect 1390 3465 1700 3505
rect 1740 3465 2050 3505
rect 2090 3465 2400 3505
rect 2440 3465 2750 3505
rect 2790 3465 3100 3505
rect 3140 3465 3450 3505
rect 3490 3465 3800 3505
rect 3840 3465 4150 3505
rect 4190 3465 4500 3505
rect 4540 3465 4850 3505
rect 4890 3465 4895 3505
rect 995 3460 4895 3465
rect 995 3145 1045 3460
rect 995 3105 1000 3145
rect 1040 3105 1045 3145
rect 995 3100 1045 3105
rect 1345 3145 1395 3460
rect 1345 3105 1350 3145
rect 1390 3105 1395 3145
rect 1345 3100 1395 3105
rect 1695 3145 1745 3460
rect 1695 3105 1700 3145
rect 1740 3105 1745 3145
rect 2045 3155 2095 3460
rect 2045 3115 2050 3155
rect 2090 3115 2095 3155
rect 2045 3110 2095 3115
rect 2395 3155 2445 3460
rect 2395 3115 2400 3155
rect 2440 3115 2445 3155
rect 1695 3100 1745 3105
rect -755 2765 -750 2805
rect -710 2765 -705 2805
rect -755 2455 -705 2765
rect -755 2415 -750 2455
rect -710 2415 -705 2455
rect -755 2410 -705 2415
rect 2395 2805 2445 3115
rect 2395 2765 2400 2805
rect 2440 2765 2445 2805
rect 2395 2455 2445 2765
rect 2395 2415 2400 2455
rect 2440 2415 2445 2455
rect 2395 2410 2445 2415
rect 2745 3155 2795 3460
rect 2745 3115 2750 3155
rect 2790 3115 2795 3155
rect 2745 2805 2795 3115
rect 2745 2765 2750 2805
rect 2790 2765 2795 2805
rect 2745 2455 2795 2765
rect 2745 2415 2750 2455
rect 2790 2415 2795 2455
rect 2745 2410 2795 2415
rect 3095 3155 3145 3460
rect 3095 3115 3100 3155
rect 3140 3115 3145 3155
rect 3095 2805 3145 3115
rect 3095 2765 3100 2805
rect 3140 2765 3145 2805
rect 3095 2455 3145 2765
rect 3445 3155 3495 3460
rect 4145 3160 4195 3460
rect 3445 3115 3450 3155
rect 3490 3115 3495 3155
rect 3445 2805 3495 3115
rect 3795 3155 4895 3160
rect 3795 3115 3800 3155
rect 3840 3115 4150 3155
rect 4190 3115 4500 3155
rect 4540 3115 4850 3155
rect 4890 3115 4895 3155
rect 3795 3110 4895 3115
rect 4145 2810 4195 3110
rect 3445 2765 3450 2805
rect 3490 2765 3495 2805
rect 3445 2760 3495 2765
rect 3795 2805 4895 2810
rect 3795 2765 3800 2805
rect 3840 2765 4150 2805
rect 4190 2765 4500 2805
rect 4540 2765 4850 2805
rect 4890 2765 4895 2805
rect 3795 2760 4895 2765
rect 4145 2460 4195 2760
rect 3095 2415 3100 2455
rect 3140 2415 3145 2455
rect 3095 2410 3145 2415
rect 3445 2455 4895 2460
rect 3445 2415 3450 2455
rect 3490 2415 3800 2455
rect 3840 2415 4150 2455
rect 4190 2415 4500 2455
rect 4540 2415 4850 2455
rect 4890 2415 4895 2455
rect 3445 2410 4895 2415
rect -2505 2110 -2455 2410
rect 4145 2110 4195 2410
rect -3205 2105 -1755 2110
rect -3205 2065 -3200 2105
rect -3160 2065 -2850 2105
rect -2810 2065 -2500 2105
rect -2460 2065 -2150 2105
rect -2110 2065 -1800 2105
rect -1760 2065 -1755 2105
rect -3205 2060 -1755 2065
rect 3445 2105 4895 2110
rect 3445 2065 3450 2105
rect 3490 2065 3800 2105
rect 3840 2065 4150 2105
rect 4190 2065 4500 2105
rect 4540 2065 4850 2105
rect 4890 2065 4895 2105
rect 3445 2060 4895 2065
rect -2505 1760 -2455 2060
rect 4145 1760 4195 2060
rect -3205 1755 -1755 1760
rect -3205 1715 -3200 1755
rect -3160 1715 -2850 1755
rect -2810 1715 -2500 1755
rect -2460 1715 -2150 1755
rect -2110 1715 -1800 1755
rect -1760 1715 -1755 1755
rect -3205 1710 -1755 1715
rect 3445 1755 4895 1760
rect 3445 1715 3450 1755
rect 3490 1715 3800 1755
rect 3840 1715 4150 1755
rect 4190 1715 4500 1755
rect 4540 1715 4850 1755
rect 4890 1715 4895 1755
rect 3445 1710 4895 1715
rect -2505 1410 -2455 1710
rect 4145 1410 4195 1710
rect -3205 1405 -1755 1410
rect -3205 1365 -3200 1405
rect -3160 1365 -2850 1405
rect -2810 1365 -2500 1405
rect -2460 1365 -2150 1405
rect -2110 1365 -1800 1405
rect -1760 1365 -1755 1405
rect -3205 1360 -1755 1365
rect 3445 1405 4895 1410
rect 3445 1365 3450 1405
rect 3490 1365 3800 1405
rect 3840 1365 4150 1405
rect 4190 1365 4500 1405
rect 4540 1365 4850 1405
rect 4890 1365 4895 1405
rect 3445 1360 4895 1365
rect -2505 1060 -2455 1360
rect 4145 1060 4195 1360
rect -3205 1055 -1755 1060
rect -3205 1015 -3200 1055
rect -3160 1015 -2850 1055
rect -2810 1015 -2500 1055
rect -2460 1015 -2150 1055
rect -2110 1015 -1800 1055
rect -1760 1015 -1755 1055
rect -3205 1010 -1755 1015
rect 3445 1055 4895 1060
rect 3445 1015 3450 1055
rect 3490 1015 3800 1055
rect 3840 1015 4150 1055
rect 4190 1015 4500 1055
rect 4540 1015 4850 1055
rect 4890 1015 4895 1055
rect 3445 1010 4895 1015
rect -2505 710 -2455 1010
rect 4145 710 4195 1010
rect -3205 705 -1755 710
rect -3205 665 -3200 705
rect -3160 665 -2850 705
rect -2810 665 -2500 705
rect -2460 665 -2150 705
rect -2110 665 -1800 705
rect -1760 665 -1755 705
rect -3205 660 -1755 665
rect 3445 705 4895 710
rect 3445 665 3450 705
rect 3490 665 3800 705
rect 3840 665 4150 705
rect 4190 665 4500 705
rect 4540 665 4850 705
rect 4890 665 4895 705
rect 3445 660 4895 665
rect -2505 360 -2455 660
rect 4145 360 4195 660
rect -3205 355 -1495 360
rect -3205 315 -3200 355
rect -3160 315 -2850 355
rect -2810 315 -2500 355
rect -2460 315 -2150 355
rect -2110 315 -1800 355
rect -1760 315 -1540 355
rect -1500 315 -1495 355
rect -3205 310 -1495 315
rect 3185 355 4895 360
rect 3185 315 3190 355
rect 3230 315 3450 355
rect 3490 315 3800 355
rect 3840 315 4150 355
rect 4190 315 4500 355
rect 4540 315 4850 355
rect 4890 315 4895 355
rect 3185 310 4895 315
rect -2505 10 -2455 310
rect 4145 10 4195 310
rect -3205 5 -1755 10
rect -3205 -35 -3200 5
rect -3160 -35 -2850 5
rect -2810 -35 -2500 5
rect -2460 -35 -2150 5
rect -2110 -35 -1800 5
rect -1760 -35 -1755 5
rect -3205 -40 -1755 -35
rect 3445 5 4895 10
rect 3445 -35 3450 5
rect 3490 -35 3800 5
rect 3840 -35 4150 5
rect 4190 -35 4500 5
rect 4540 -35 4850 5
rect 4890 -35 4895 5
rect 3445 -40 4895 -35
rect -2505 -340 -2455 -40
rect 4145 -340 4195 -40
rect -3205 -345 -1755 -340
rect -3205 -385 -3200 -345
rect -3160 -385 -2850 -345
rect -2810 -385 -2500 -345
rect -2460 -385 -2150 -345
rect -2110 -385 -1800 -345
rect -1760 -385 -1755 -345
rect -3205 -390 -1755 -385
rect 3445 -345 4895 -340
rect 3445 -385 3450 -345
rect 3490 -385 3800 -345
rect 3840 -385 4150 -345
rect 4190 -385 4500 -345
rect 4540 -385 4850 -345
rect 4890 -385 4895 -345
rect 3445 -390 4895 -385
rect -2505 -690 -2455 -390
rect 4145 -690 4195 -390
rect -3205 -695 -1755 -690
rect -3205 -735 -3200 -695
rect -3160 -735 -2850 -695
rect -2810 -735 -2500 -695
rect -2460 -735 -2150 -695
rect -2110 -735 -1800 -695
rect -1760 -735 -1755 -695
rect -3205 -740 -1755 -735
rect 3445 -695 4895 -690
rect 3445 -735 3450 -695
rect 3490 -735 3800 -695
rect 3840 -735 4150 -695
rect 4190 -735 4500 -695
rect 4540 -735 4850 -695
rect 4890 -735 4895 -695
rect 3445 -740 4895 -735
rect -2505 -1040 -2455 -740
rect 4145 -1040 4195 -740
rect -3205 -1045 -1755 -1040
rect -3205 -1085 -3200 -1045
rect -3160 -1085 -2850 -1045
rect -2810 -1085 -2500 -1045
rect -2460 -1085 -2150 -1045
rect -2110 -1085 -1800 -1045
rect -1760 -1085 -1755 -1045
rect -3205 -1090 -1755 -1085
rect 3445 -1045 4895 -1040
rect 3445 -1085 3450 -1045
rect 3490 -1085 3800 -1045
rect 3840 -1085 4150 -1045
rect 4190 -1085 4500 -1045
rect 4540 -1085 4850 -1045
rect 4890 -1085 4895 -1045
rect 3445 -1090 4895 -1085
rect -2505 -1390 -2455 -1090
rect 4145 -1390 4195 -1090
rect -3205 -1395 -1755 -1390
rect -3205 -1435 -3200 -1395
rect -3160 -1435 -2850 -1395
rect -2810 -1435 -2500 -1395
rect -2460 -1435 -2150 -1395
rect -2110 -1435 -1800 -1395
rect -1760 -1435 -1755 -1395
rect -3205 -1440 -1755 -1435
rect -1455 -1395 -1405 -1390
rect -1455 -1435 -1450 -1395
rect -1410 -1435 -1405 -1395
rect -2505 -1740 -2455 -1440
rect -1455 -1740 -1405 -1435
rect -1105 -1395 -1055 -1390
rect -1105 -1435 -1100 -1395
rect -1060 -1435 -1055 -1395
rect -1105 -1740 -1055 -1435
rect -755 -1395 -705 -1390
rect -755 -1435 -750 -1395
rect -710 -1435 -705 -1395
rect -755 -1740 -705 -1435
rect -405 -1395 -355 -1390
rect -405 -1435 -400 -1395
rect -360 -1435 -355 -1395
rect -405 -1740 -355 -1435
rect -55 -1395 -5 -1390
rect -55 -1435 -50 -1395
rect -10 -1435 -5 -1395
rect -55 -1740 -5 -1435
rect 295 -1395 345 -1390
rect 295 -1435 300 -1395
rect 340 -1435 345 -1395
rect 295 -1740 345 -1435
rect 645 -1395 695 -1390
rect 645 -1435 650 -1395
rect 690 -1435 695 -1395
rect 645 -1740 695 -1435
rect -3205 -1745 695 -1740
rect -3205 -1785 -3200 -1745
rect -3160 -1785 -2850 -1745
rect -2810 -1785 -2500 -1745
rect -2460 -1785 -2150 -1745
rect -2110 -1785 -1800 -1745
rect -1760 -1785 -1450 -1745
rect -1410 -1785 -1100 -1745
rect -1060 -1785 -750 -1745
rect -710 -1785 -400 -1745
rect -360 -1785 -50 -1745
rect -10 -1785 300 -1745
rect 340 -1785 650 -1745
rect 690 -1785 695 -1745
rect -3205 -1790 695 -1785
rect -2505 -2090 -2455 -1790
rect -3205 -2095 -2455 -2090
rect -3205 -2135 -3200 -2095
rect -3160 -2135 -2850 -2095
rect -2810 -2135 -2500 -2095
rect -2460 -2135 -2455 -2095
rect -3205 -2140 -2455 -2135
rect -2155 -2095 -2105 -1790
rect -2155 -2135 -2150 -2095
rect -2110 -2135 -2105 -2095
rect -2155 -2140 -2105 -2135
rect -1805 -2095 -1755 -1790
rect -1805 -2135 -1800 -2095
rect -1760 -2135 -1755 -2095
rect -1805 -2140 -1755 -2135
rect -1455 -2095 -1405 -1790
rect -1455 -2135 -1450 -2095
rect -1410 -2135 -1405 -2095
rect -1455 -2140 -1405 -2135
rect -1105 -2095 -1055 -1790
rect -1105 -2135 -1100 -2095
rect -1060 -2135 -1055 -2095
rect -1105 -2140 -1055 -2135
rect -755 -2095 -705 -1790
rect -755 -2135 -750 -2095
rect -710 -2135 -705 -2095
rect -755 -2140 -705 -2135
rect -405 -2095 -355 -1790
rect -405 -2135 -400 -2095
rect -360 -2135 -355 -2095
rect -405 -2140 -355 -2135
rect -55 -2095 -5 -1790
rect -55 -2135 -50 -2095
rect -10 -2135 -5 -2095
rect -55 -2140 -5 -2135
rect 295 -2095 345 -1790
rect 295 -2135 300 -2095
rect 340 -2135 345 -2095
rect 295 -2140 345 -2135
rect 645 -2095 695 -1790
rect 645 -2135 650 -2095
rect 690 -2135 695 -2095
rect 645 -2140 695 -2135
rect 995 -1395 1045 -1390
rect 995 -1435 1000 -1395
rect 1040 -1435 1045 -1395
rect 995 -1740 1045 -1435
rect 1345 -1395 1395 -1390
rect 1345 -1435 1350 -1395
rect 1390 -1435 1395 -1395
rect 1345 -1740 1395 -1435
rect 1695 -1395 1745 -1390
rect 1695 -1435 1700 -1395
rect 1740 -1435 1745 -1395
rect 1695 -1740 1745 -1435
rect 2045 -1395 2095 -1390
rect 2045 -1435 2050 -1395
rect 2090 -1435 2095 -1395
rect 2045 -1740 2095 -1435
rect 2395 -1395 2445 -1390
rect 2395 -1435 2400 -1395
rect 2440 -1435 2445 -1395
rect 2395 -1740 2445 -1435
rect 2745 -1395 2795 -1390
rect 2745 -1435 2750 -1395
rect 2790 -1435 2795 -1395
rect 2745 -1740 2795 -1435
rect 3095 -1395 3145 -1390
rect 3095 -1435 3100 -1395
rect 3140 -1435 3145 -1395
rect 3095 -1740 3145 -1435
rect 3445 -1395 4895 -1390
rect 3445 -1435 3450 -1395
rect 3490 -1435 3800 -1395
rect 3840 -1435 4150 -1395
rect 4190 -1435 4500 -1395
rect 4540 -1435 4850 -1395
rect 4890 -1435 4895 -1395
rect 3445 -1440 4895 -1435
rect 4145 -1740 4195 -1440
rect 995 -1745 4895 -1740
rect 995 -1785 1000 -1745
rect 1040 -1785 1350 -1745
rect 1390 -1785 1700 -1745
rect 1740 -1785 2050 -1745
rect 2090 -1785 2400 -1745
rect 2440 -1785 2750 -1745
rect 2790 -1785 3100 -1745
rect 3140 -1785 3450 -1745
rect 3490 -1785 3800 -1745
rect 3840 -1785 4150 -1745
rect 4190 -1785 4500 -1745
rect 4540 -1785 4850 -1745
rect 4890 -1785 4895 -1745
rect 995 -1790 4895 -1785
rect 995 -2095 1045 -1790
rect 995 -2135 1000 -2095
rect 1040 -2135 1045 -2095
rect 995 -2140 1045 -2135
rect 1345 -2095 1395 -1790
rect 1345 -2135 1350 -2095
rect 1390 -2135 1395 -2095
rect 1345 -2140 1395 -2135
rect 1695 -2095 1745 -1790
rect 1695 -2135 1700 -2095
rect 1740 -2135 1745 -2095
rect 1695 -2140 1745 -2135
rect 2045 -2095 2095 -1790
rect 2045 -2135 2050 -2095
rect 2090 -2135 2095 -2095
rect 2045 -2140 2095 -2135
rect 2395 -2095 2445 -1790
rect 2395 -2135 2400 -2095
rect 2440 -2135 2445 -2095
rect 2395 -2140 2445 -2135
rect 2745 -2095 2795 -1790
rect 2745 -2135 2750 -2095
rect 2790 -2135 2795 -2095
rect 2745 -2140 2795 -2135
rect 3095 -2095 3145 -1790
rect 3095 -2135 3100 -2095
rect 3140 -2135 3145 -2095
rect 3095 -2140 3145 -2135
rect 3445 -2095 3495 -1790
rect 3445 -2135 3450 -2095
rect 3490 -2135 3495 -2095
rect 3445 -2140 3495 -2135
rect 3795 -2095 3845 -1790
rect 3795 -2135 3800 -2095
rect 3840 -2135 3845 -2095
rect 3795 -2140 3845 -2135
rect 4145 -2090 4195 -1790
rect 4145 -2095 4895 -2090
rect 4145 -2135 4150 -2095
rect 4190 -2135 4500 -2095
rect 4540 -2135 4850 -2095
rect 4890 -2135 4895 -2095
rect 4145 -2140 4895 -2135
rect -3850 -2420 5140 -2415
rect -3850 -2460 825 -2420
rect 865 -2460 5140 -2420
rect -3850 -2465 5140 -2460
<< labels >>
flabel metal3 3100 1595 3100 1595 7 FreeSans 240 0 -80 0 cap_res_X
flabel metal3 -1410 1610 -1410 1610 3 FreeSans 240 0 80 0 cap_res_Y
flabel metal4 -3850 -2440 -3850 -2440 7 FreeSans 240 0 -80 0 GNDA
port 16 w
flabel metal2 1310 2775 1310 2775 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 400 2775 400 2775 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 1125 1520 1125 1520 3 FreeSans 240 0 80 0 V_err_p
flabel metal1 565 1520 565 1520 7 FreeSans 240 0 -80 0 V_err_mir_p
flabel metal2 310 1140 310 1140 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal2 1525 1100 1525 1100 1 FreeSans 240 0 0 160 V_tot
flabel metal2 1070 1200 1070 1200 3 FreeSans 240 0 80 0 V_err_gate
port 13 e
flabel metal2 945 1045 945 1045 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal1 -350 305 -350 305 5 FreeSans 240 0 0 -80 Y
flabel metal1 1455 580 1455 580 3 FreeSans 240 0 80 0 VD1
flabel metal1 235 580 235 580 7 FreeSans 240 0 -80 0 VD2
flabel metal1 910 50 910 50 3 FreeSans 240 0 80 0 V_p_mir
flabel metal1 1970 2135 1970 2135 3 FreeSans 240 0 80 0 VD3
flabel metal2 965 -1135 965 -1135 3 FreeSans 240 0 80 0 Vb1_2
flabel metal2 460 20 460 20 1 FreeSans 240 0 0 80 V_tail_gate
port 11 n
flabel metal1 1235 -140 1235 -140 3 FreeSans 240 0 80 0 V_source
flabel metal2 1470 1005 1470 1005 1 FreeSans 240 0 0 80 err_amp_out
flabel metal2 -105 535 -105 535 7 FreeSans 240 0 -80 0 VIN+
port 14 w
flabel metal2 1795 535 1795 535 3 FreeSans 240 0 80 0 VIN-
port 15 e
flabel metal1 -280 2135 -280 2135 7 FreeSans 240 0 -80 0 VD4
flabel metal1 2940 405 2940 405 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 2895 285 2895 285 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal1 2040 305 2040 305 5 FreeSans 240 0 0 -80 X
flabel metal1 3210 -340 3210 -340 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal2 1570 -390 1570 -390 5 FreeSans 240 0 0 -80 V_b_2nd_stage
flabel metal1 -1520 -340 -1520 -340 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal1 -1205 285 -1205 285 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal1 -1250 405 -1250 405 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal2 845 945 845 945 1 FreeSans 240 0 0 80 Vb1
port 6 n
flabel metal4 -3850 4260 -3850 4260 7 FreeSans 240 0 -80 0 VDDA
port 1 w
flabel metal2 2260 1600 2260 1600 5 FreeSans 240 0 0 -80 Vb3
port 4 s
flabel metal2 1070 1665 1070 1665 1 FreeSans 240 0 0 80 Vb2
port 5 n
<< end >>
