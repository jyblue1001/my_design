magic
tech sky130A
timestamp 1754014703
<< nwell >>
rect 16315 1110 16695 1250
rect 16825 1110 17315 1250
rect 17445 1110 18155 1250
rect 18285 1110 18775 1250
rect 16375 545 16760 685
rect 16910 445 18690 785
rect 18845 545 19170 785
rect 16360 -195 17725 -55
rect 17880 -195 19240 -55
<< pwell >>
rect 17780 -4300 17820 -4120
<< nmos >>
rect 17000 -610 17020 -360
rect 17060 -610 17080 -360
rect 18520 -610 18540 -360
rect 18580 -610 18600 -360
rect 16570 -1060 17070 -810
rect 17190 -1060 17690 -810
rect 17910 -1060 18410 -810
rect 18530 -1060 19030 -810
rect 16780 -1290 17780 -1190
rect 17820 -1290 18820 -1190
rect 16580 -1640 16595 -1540
rect 16635 -1640 16650 -1540
rect 16690 -1640 16705 -1540
rect 16745 -1640 16760 -1540
rect 16800 -1640 16815 -1540
rect 17065 -1640 17080 -1540
rect 17120 -1640 17135 -1540
rect 17175 -1640 17190 -1540
rect 17230 -1640 17245 -1540
rect 17285 -1640 17300 -1540
rect 17340 -1640 17355 -1540
rect 17395 -1640 17410 -1540
rect 17450 -1640 17465 -1540
rect 17655 -1640 17670 -1540
rect 17710 -1640 17725 -1540
rect 17765 -1640 17780 -1540
rect 17820 -1640 17835 -1540
rect 17875 -1640 17890 -1540
rect 17930 -1640 17945 -1540
rect 18135 -1640 18150 -1540
rect 18190 -1640 18205 -1540
rect 18245 -1640 18260 -1540
rect 18300 -1640 18315 -1540
rect 18355 -1640 18370 -1540
rect 18410 -1640 18425 -1540
rect 18465 -1640 18480 -1540
rect 18520 -1640 18535 -1540
<< pmos >>
rect 16415 1130 16430 1230
rect 16470 1130 16485 1230
rect 16525 1130 16540 1230
rect 16580 1130 16595 1230
rect 16925 1130 16940 1230
rect 16980 1130 16995 1230
rect 17035 1130 17050 1230
rect 17090 1130 17105 1230
rect 17145 1130 17160 1230
rect 17200 1130 17215 1230
rect 17545 1130 17560 1230
rect 17600 1130 17615 1230
rect 17655 1130 17670 1230
rect 17710 1130 17725 1230
rect 17765 1130 17780 1230
rect 17820 1130 17835 1230
rect 17875 1130 17890 1230
rect 17930 1130 17945 1230
rect 17985 1130 18000 1230
rect 18040 1130 18055 1230
rect 18385 1130 18400 1230
rect 18440 1130 18455 1230
rect 18495 1130 18510 1230
rect 18550 1130 18565 1230
rect 18605 1130 18620 1230
rect 18660 1130 18675 1230
rect 16475 565 16490 665
rect 16530 565 16545 665
rect 16585 565 16600 665
rect 16640 565 16655 665
rect 17010 465 17060 765
rect 17100 465 17150 765
rect 17190 465 17240 765
rect 17280 465 17330 765
rect 17370 465 17420 765
rect 17460 465 17510 765
rect 17550 465 17600 765
rect 17640 465 17690 765
rect 17730 465 17780 765
rect 17820 465 17870 765
rect 17910 465 17960 765
rect 18000 465 18050 765
rect 18090 465 18140 765
rect 18180 465 18230 765
rect 18270 465 18320 765
rect 18360 465 18410 765
rect 18450 465 18500 765
rect 18540 465 18590 765
rect 18945 565 18960 765
rect 19000 565 19015 765
rect 19055 565 19070 765
rect 16460 -175 16480 -75
rect 16520 -175 16540 -75
rect 16580 -175 16600 -75
rect 16640 -175 16660 -75
rect 16700 -175 16720 -75
rect 16760 -175 16780 -75
rect 16820 -175 16840 -75
rect 16880 -175 16900 -75
rect 16940 -175 16960 -75
rect 17000 -175 17020 -75
rect 17060 -175 17080 -75
rect 17120 -175 17140 -75
rect 17180 -175 17200 -75
rect 17240 -175 17260 -75
rect 17300 -175 17320 -75
rect 17360 -175 17380 -75
rect 17420 -175 17440 -75
rect 17480 -175 17500 -75
rect 17540 -175 17560 -75
rect 17600 -175 17620 -75
rect 17980 -175 18000 -75
rect 18040 -175 18060 -75
rect 18100 -175 18120 -75
rect 18160 -175 18180 -75
rect 18220 -175 18240 -75
rect 18280 -175 18300 -75
rect 18340 -175 18360 -75
rect 18400 -175 18420 -75
rect 18460 -175 18480 -75
rect 18520 -175 18540 -75
rect 18580 -175 18600 -75
rect 18640 -175 18660 -75
rect 18700 -175 18720 -75
rect 18760 -175 18780 -75
rect 18820 -175 18840 -75
rect 18880 -175 18900 -75
rect 18940 -175 18960 -75
rect 19000 -175 19020 -75
rect 19060 -175 19080 -75
rect 19120 -175 19140 -75
<< ndiff >>
rect 16960 -375 17000 -360
rect 16960 -395 16970 -375
rect 16990 -395 17000 -375
rect 16960 -425 17000 -395
rect 16960 -445 16970 -425
rect 16990 -445 17000 -425
rect 16960 -475 17000 -445
rect 16960 -495 16970 -475
rect 16990 -495 17000 -475
rect 16960 -525 17000 -495
rect 16960 -545 16970 -525
rect 16990 -545 17000 -525
rect 16960 -575 17000 -545
rect 16960 -595 16970 -575
rect 16990 -595 17000 -575
rect 16960 -610 17000 -595
rect 17020 -375 17060 -360
rect 17020 -395 17030 -375
rect 17050 -395 17060 -375
rect 17020 -425 17060 -395
rect 17020 -445 17030 -425
rect 17050 -445 17060 -425
rect 17020 -475 17060 -445
rect 17020 -495 17030 -475
rect 17050 -495 17060 -475
rect 17020 -525 17060 -495
rect 17020 -545 17030 -525
rect 17050 -545 17060 -525
rect 17020 -575 17060 -545
rect 17020 -595 17030 -575
rect 17050 -595 17060 -575
rect 17020 -610 17060 -595
rect 17080 -375 17120 -360
rect 17080 -395 17090 -375
rect 17110 -395 17120 -375
rect 17080 -425 17120 -395
rect 18480 -375 18520 -360
rect 18480 -395 18490 -375
rect 18510 -395 18520 -375
rect 17080 -445 17090 -425
rect 17110 -445 17120 -425
rect 17080 -475 17120 -445
rect 17080 -495 17090 -475
rect 17110 -495 17120 -475
rect 17080 -525 17120 -495
rect 17080 -545 17090 -525
rect 17110 -545 17120 -525
rect 17080 -575 17120 -545
rect 17080 -595 17090 -575
rect 17110 -595 17120 -575
rect 17080 -610 17120 -595
rect 18480 -425 18520 -395
rect 18480 -445 18490 -425
rect 18510 -445 18520 -425
rect 18480 -475 18520 -445
rect 18480 -495 18490 -475
rect 18510 -495 18520 -475
rect 18480 -525 18520 -495
rect 18480 -545 18490 -525
rect 18510 -545 18520 -525
rect 18480 -575 18520 -545
rect 18480 -595 18490 -575
rect 18510 -595 18520 -575
rect 18480 -610 18520 -595
rect 18540 -375 18580 -360
rect 18540 -395 18550 -375
rect 18570 -395 18580 -375
rect 18540 -425 18580 -395
rect 18540 -445 18550 -425
rect 18570 -445 18580 -425
rect 18540 -475 18580 -445
rect 18540 -495 18550 -475
rect 18570 -495 18580 -475
rect 18540 -525 18580 -495
rect 18540 -545 18550 -525
rect 18570 -545 18580 -525
rect 18540 -575 18580 -545
rect 18540 -595 18550 -575
rect 18570 -595 18580 -575
rect 18540 -610 18580 -595
rect 18600 -375 18640 -360
rect 18600 -395 18610 -375
rect 18630 -395 18640 -375
rect 18600 -425 18640 -395
rect 18600 -445 18610 -425
rect 18630 -445 18640 -425
rect 18600 -475 18640 -445
rect 18600 -495 18610 -475
rect 18630 -495 18640 -475
rect 18600 -525 18640 -495
rect 18600 -545 18610 -525
rect 18630 -545 18640 -525
rect 18600 -575 18640 -545
rect 18600 -595 18610 -575
rect 18630 -595 18640 -575
rect 18600 -610 18640 -595
rect 16530 -825 16570 -810
rect 16530 -845 16540 -825
rect 16560 -845 16570 -825
rect 16530 -875 16570 -845
rect 16530 -895 16540 -875
rect 16560 -895 16570 -875
rect 16530 -925 16570 -895
rect 16530 -945 16540 -925
rect 16560 -945 16570 -925
rect 16530 -975 16570 -945
rect 16530 -995 16540 -975
rect 16560 -995 16570 -975
rect 16530 -1025 16570 -995
rect 16530 -1045 16540 -1025
rect 16560 -1045 16570 -1025
rect 16530 -1060 16570 -1045
rect 17070 -825 17110 -810
rect 17150 -825 17190 -810
rect 17070 -845 17080 -825
rect 17100 -845 17110 -825
rect 17150 -845 17160 -825
rect 17180 -845 17190 -825
rect 17070 -875 17110 -845
rect 17150 -875 17190 -845
rect 17070 -895 17080 -875
rect 17100 -895 17110 -875
rect 17150 -895 17160 -875
rect 17180 -895 17190 -875
rect 17070 -925 17110 -895
rect 17150 -925 17190 -895
rect 17070 -945 17080 -925
rect 17100 -945 17110 -925
rect 17150 -945 17160 -925
rect 17180 -945 17190 -925
rect 17070 -975 17110 -945
rect 17150 -975 17190 -945
rect 17070 -995 17080 -975
rect 17100 -995 17110 -975
rect 17150 -995 17160 -975
rect 17180 -995 17190 -975
rect 17070 -1025 17110 -995
rect 17150 -1025 17190 -995
rect 17070 -1045 17080 -1025
rect 17100 -1045 17110 -1025
rect 17150 -1045 17160 -1025
rect 17180 -1045 17190 -1025
rect 17070 -1055 17110 -1045
rect 17150 -1055 17190 -1045
rect 17070 -1060 17190 -1055
rect 17690 -825 17730 -810
rect 17690 -845 17700 -825
rect 17720 -845 17730 -825
rect 17690 -875 17730 -845
rect 17690 -895 17700 -875
rect 17720 -895 17730 -875
rect 17690 -925 17730 -895
rect 17690 -945 17700 -925
rect 17720 -945 17730 -925
rect 17690 -975 17730 -945
rect 17690 -995 17700 -975
rect 17720 -995 17730 -975
rect 17690 -1025 17730 -995
rect 17690 -1045 17700 -1025
rect 17720 -1045 17730 -1025
rect 17690 -1060 17730 -1045
rect 17870 -825 17910 -810
rect 17870 -845 17880 -825
rect 17900 -845 17910 -825
rect 17870 -875 17910 -845
rect 17870 -895 17880 -875
rect 17900 -895 17910 -875
rect 17870 -925 17910 -895
rect 17870 -945 17880 -925
rect 17900 -945 17910 -925
rect 17870 -975 17910 -945
rect 17870 -995 17880 -975
rect 17900 -995 17910 -975
rect 17870 -1025 17910 -995
rect 17870 -1045 17880 -1025
rect 17900 -1045 17910 -1025
rect 17870 -1060 17910 -1045
rect 18410 -825 18450 -810
rect 18490 -825 18530 -810
rect 18410 -845 18420 -825
rect 18440 -845 18450 -825
rect 18490 -845 18500 -825
rect 18520 -845 18530 -825
rect 18410 -875 18450 -845
rect 18490 -875 18530 -845
rect 18410 -895 18420 -875
rect 18440 -895 18450 -875
rect 18490 -895 18500 -875
rect 18520 -895 18530 -875
rect 18410 -925 18450 -895
rect 18490 -925 18530 -895
rect 18410 -945 18420 -925
rect 18440 -945 18450 -925
rect 18490 -945 18500 -925
rect 18520 -945 18530 -925
rect 18410 -975 18450 -945
rect 18490 -975 18530 -945
rect 18410 -995 18420 -975
rect 18440 -995 18450 -975
rect 18490 -995 18500 -975
rect 18520 -995 18530 -975
rect 18410 -1025 18450 -995
rect 18490 -1025 18530 -995
rect 18410 -1045 18420 -1025
rect 18440 -1045 18450 -1025
rect 18490 -1045 18500 -1025
rect 18520 -1045 18530 -1025
rect 18410 -1060 18450 -1045
rect 18490 -1060 18530 -1045
rect 19030 -825 19070 -810
rect 19030 -845 19040 -825
rect 19060 -845 19070 -825
rect 19030 -875 19070 -845
rect 19030 -895 19040 -875
rect 19060 -895 19070 -875
rect 19030 -925 19070 -895
rect 19030 -945 19040 -925
rect 19060 -945 19070 -925
rect 19030 -975 19070 -945
rect 19030 -995 19040 -975
rect 19060 -995 19070 -975
rect 19030 -1025 19070 -995
rect 19030 -1045 19040 -1025
rect 19060 -1045 19070 -1025
rect 19030 -1060 19070 -1045
rect 16740 -1205 16780 -1190
rect 16740 -1225 16750 -1205
rect 16770 -1225 16780 -1205
rect 16740 -1255 16780 -1225
rect 16740 -1275 16750 -1255
rect 16770 -1275 16780 -1255
rect 16740 -1290 16780 -1275
rect 17780 -1205 17820 -1190
rect 17780 -1225 17790 -1205
rect 17810 -1225 17820 -1205
rect 17780 -1255 17820 -1225
rect 17780 -1275 17790 -1255
rect 17810 -1275 17820 -1255
rect 17780 -1290 17820 -1275
rect 18820 -1205 18860 -1190
rect 18820 -1225 18830 -1205
rect 18850 -1225 18860 -1205
rect 18820 -1255 18860 -1225
rect 18820 -1275 18830 -1255
rect 18850 -1275 18860 -1255
rect 18820 -1290 18860 -1275
rect 16540 -1555 16580 -1540
rect 16540 -1575 16550 -1555
rect 16570 -1575 16580 -1555
rect 16540 -1605 16580 -1575
rect 16540 -1625 16550 -1605
rect 16570 -1625 16580 -1605
rect 16540 -1640 16580 -1625
rect 16595 -1555 16635 -1540
rect 16595 -1575 16605 -1555
rect 16625 -1575 16635 -1555
rect 16595 -1605 16635 -1575
rect 16595 -1625 16605 -1605
rect 16625 -1625 16635 -1605
rect 16595 -1640 16635 -1625
rect 16650 -1555 16690 -1540
rect 16650 -1575 16660 -1555
rect 16680 -1575 16690 -1555
rect 16650 -1605 16690 -1575
rect 16650 -1625 16660 -1605
rect 16680 -1625 16690 -1605
rect 16650 -1640 16690 -1625
rect 16705 -1555 16745 -1540
rect 16705 -1575 16715 -1555
rect 16735 -1575 16745 -1555
rect 16705 -1605 16745 -1575
rect 16705 -1625 16715 -1605
rect 16735 -1625 16745 -1605
rect 16705 -1640 16745 -1625
rect 16760 -1555 16800 -1540
rect 16760 -1575 16770 -1555
rect 16790 -1575 16800 -1555
rect 16760 -1605 16800 -1575
rect 16760 -1625 16770 -1605
rect 16790 -1625 16800 -1605
rect 16760 -1640 16800 -1625
rect 16815 -1555 16855 -1540
rect 16815 -1575 16825 -1555
rect 16845 -1575 16855 -1555
rect 16815 -1605 16855 -1575
rect 16815 -1625 16825 -1605
rect 16845 -1625 16855 -1605
rect 16815 -1640 16855 -1625
rect 17025 -1555 17065 -1540
rect 17025 -1575 17035 -1555
rect 17055 -1575 17065 -1555
rect 17025 -1605 17065 -1575
rect 17025 -1625 17035 -1605
rect 17055 -1625 17065 -1605
rect 17025 -1640 17065 -1625
rect 17080 -1555 17120 -1540
rect 17080 -1575 17090 -1555
rect 17110 -1575 17120 -1555
rect 17080 -1605 17120 -1575
rect 17080 -1625 17090 -1605
rect 17110 -1625 17120 -1605
rect 17080 -1640 17120 -1625
rect 17135 -1555 17175 -1540
rect 17135 -1575 17145 -1555
rect 17165 -1575 17175 -1555
rect 17135 -1605 17175 -1575
rect 17135 -1625 17145 -1605
rect 17165 -1625 17175 -1605
rect 17135 -1640 17175 -1625
rect 17190 -1555 17230 -1540
rect 17190 -1575 17200 -1555
rect 17220 -1575 17230 -1555
rect 17190 -1605 17230 -1575
rect 17190 -1625 17200 -1605
rect 17220 -1625 17230 -1605
rect 17190 -1640 17230 -1625
rect 17245 -1555 17285 -1540
rect 17245 -1575 17255 -1555
rect 17275 -1575 17285 -1555
rect 17245 -1605 17285 -1575
rect 17245 -1625 17255 -1605
rect 17275 -1625 17285 -1605
rect 17245 -1640 17285 -1625
rect 17300 -1555 17340 -1540
rect 17300 -1575 17310 -1555
rect 17330 -1575 17340 -1555
rect 17300 -1605 17340 -1575
rect 17300 -1625 17310 -1605
rect 17330 -1625 17340 -1605
rect 17300 -1640 17340 -1625
rect 17355 -1555 17395 -1540
rect 17355 -1575 17365 -1555
rect 17385 -1575 17395 -1555
rect 17355 -1605 17395 -1575
rect 17355 -1625 17365 -1605
rect 17385 -1625 17395 -1605
rect 17355 -1640 17395 -1625
rect 17410 -1555 17450 -1540
rect 17410 -1575 17420 -1555
rect 17440 -1575 17450 -1555
rect 17410 -1605 17450 -1575
rect 17410 -1625 17420 -1605
rect 17440 -1625 17450 -1605
rect 17410 -1640 17450 -1625
rect 17465 -1555 17505 -1540
rect 17465 -1575 17475 -1555
rect 17495 -1575 17505 -1555
rect 17465 -1605 17505 -1575
rect 17465 -1625 17475 -1605
rect 17495 -1625 17505 -1605
rect 17465 -1640 17505 -1625
rect 17615 -1555 17655 -1540
rect 17615 -1575 17625 -1555
rect 17645 -1575 17655 -1555
rect 17615 -1605 17655 -1575
rect 17615 -1625 17625 -1605
rect 17645 -1625 17655 -1605
rect 17615 -1640 17655 -1625
rect 17670 -1555 17710 -1540
rect 17670 -1575 17680 -1555
rect 17700 -1575 17710 -1555
rect 17670 -1605 17710 -1575
rect 17670 -1625 17680 -1605
rect 17700 -1625 17710 -1605
rect 17670 -1640 17710 -1625
rect 17725 -1555 17765 -1540
rect 17725 -1575 17735 -1555
rect 17755 -1575 17765 -1555
rect 17725 -1605 17765 -1575
rect 17725 -1625 17735 -1605
rect 17755 -1625 17765 -1605
rect 17725 -1640 17765 -1625
rect 17780 -1555 17820 -1540
rect 17780 -1575 17790 -1555
rect 17810 -1575 17820 -1555
rect 17780 -1605 17820 -1575
rect 17780 -1625 17790 -1605
rect 17810 -1625 17820 -1605
rect 17780 -1640 17820 -1625
rect 17835 -1555 17875 -1540
rect 17835 -1575 17845 -1555
rect 17865 -1575 17875 -1555
rect 17835 -1605 17875 -1575
rect 17835 -1625 17845 -1605
rect 17865 -1625 17875 -1605
rect 17835 -1640 17875 -1625
rect 17890 -1555 17930 -1540
rect 17890 -1575 17900 -1555
rect 17920 -1575 17930 -1555
rect 17890 -1605 17930 -1575
rect 17890 -1625 17900 -1605
rect 17920 -1625 17930 -1605
rect 17890 -1640 17930 -1625
rect 17945 -1555 17985 -1540
rect 17945 -1575 17955 -1555
rect 17975 -1575 17985 -1555
rect 17945 -1605 17985 -1575
rect 17945 -1625 17955 -1605
rect 17975 -1625 17985 -1605
rect 17945 -1640 17985 -1625
rect 18095 -1555 18135 -1540
rect 18095 -1575 18105 -1555
rect 18125 -1575 18135 -1555
rect 18095 -1605 18135 -1575
rect 18095 -1625 18105 -1605
rect 18125 -1625 18135 -1605
rect 18095 -1640 18135 -1625
rect 18150 -1555 18190 -1540
rect 18150 -1575 18160 -1555
rect 18180 -1575 18190 -1555
rect 18150 -1605 18190 -1575
rect 18150 -1625 18160 -1605
rect 18180 -1625 18190 -1605
rect 18150 -1640 18190 -1625
rect 18205 -1555 18245 -1540
rect 18205 -1575 18215 -1555
rect 18235 -1575 18245 -1555
rect 18205 -1605 18245 -1575
rect 18205 -1625 18215 -1605
rect 18235 -1625 18245 -1605
rect 18205 -1640 18245 -1625
rect 18260 -1555 18300 -1540
rect 18260 -1575 18270 -1555
rect 18290 -1575 18300 -1555
rect 18260 -1605 18300 -1575
rect 18260 -1625 18270 -1605
rect 18290 -1625 18300 -1605
rect 18260 -1640 18300 -1625
rect 18315 -1555 18355 -1540
rect 18315 -1575 18325 -1555
rect 18345 -1575 18355 -1555
rect 18315 -1605 18355 -1575
rect 18315 -1625 18325 -1605
rect 18345 -1625 18355 -1605
rect 18315 -1640 18355 -1625
rect 18370 -1555 18410 -1540
rect 18370 -1575 18380 -1555
rect 18400 -1575 18410 -1555
rect 18370 -1605 18410 -1575
rect 18370 -1625 18380 -1605
rect 18400 -1625 18410 -1605
rect 18370 -1640 18410 -1625
rect 18425 -1555 18465 -1540
rect 18425 -1575 18435 -1555
rect 18455 -1575 18465 -1555
rect 18425 -1605 18465 -1575
rect 18425 -1625 18435 -1605
rect 18455 -1625 18465 -1605
rect 18425 -1640 18465 -1625
rect 18480 -1555 18520 -1540
rect 18480 -1575 18490 -1555
rect 18510 -1575 18520 -1555
rect 18480 -1605 18520 -1575
rect 18480 -1625 18490 -1605
rect 18510 -1625 18520 -1605
rect 18480 -1640 18520 -1625
rect 18535 -1555 18575 -1540
rect 18535 -1575 18545 -1555
rect 18565 -1575 18575 -1555
rect 18535 -1605 18575 -1575
rect 18535 -1625 18545 -1605
rect 18565 -1625 18575 -1605
rect 18535 -1640 18575 -1625
<< pdiff >>
rect 16375 1215 16415 1230
rect 16375 1195 16385 1215
rect 16405 1195 16415 1215
rect 16375 1165 16415 1195
rect 16375 1145 16385 1165
rect 16405 1145 16415 1165
rect 16375 1130 16415 1145
rect 16430 1215 16470 1230
rect 16430 1195 16440 1215
rect 16460 1195 16470 1215
rect 16430 1165 16470 1195
rect 16430 1145 16440 1165
rect 16460 1145 16470 1165
rect 16430 1130 16470 1145
rect 16485 1215 16525 1230
rect 16485 1195 16495 1215
rect 16515 1195 16525 1215
rect 16485 1165 16525 1195
rect 16485 1145 16495 1165
rect 16515 1145 16525 1165
rect 16485 1130 16525 1145
rect 16540 1215 16580 1230
rect 16540 1195 16550 1215
rect 16570 1195 16580 1215
rect 16540 1165 16580 1195
rect 16540 1145 16550 1165
rect 16570 1145 16580 1165
rect 16540 1130 16580 1145
rect 16595 1215 16635 1230
rect 16595 1195 16605 1215
rect 16625 1195 16635 1215
rect 16595 1165 16635 1195
rect 16595 1145 16605 1165
rect 16625 1145 16635 1165
rect 16595 1130 16635 1145
rect 16885 1215 16925 1230
rect 16885 1143 16895 1215
rect 16915 1143 16925 1215
rect 16885 1130 16925 1143
rect 16940 1215 16980 1230
rect 16940 1143 16950 1215
rect 16970 1143 16980 1215
rect 16940 1130 16980 1143
rect 16995 1215 17035 1230
rect 16995 1143 17005 1215
rect 17025 1143 17035 1215
rect 16995 1130 17035 1143
rect 17050 1215 17090 1230
rect 17050 1143 17060 1215
rect 17080 1143 17090 1215
rect 17050 1130 17090 1143
rect 17105 1215 17145 1230
rect 17105 1143 17115 1215
rect 17135 1143 17145 1215
rect 17105 1130 17145 1143
rect 17160 1215 17200 1230
rect 17160 1143 17170 1215
rect 17190 1143 17200 1215
rect 17160 1130 17200 1143
rect 17215 1215 17255 1230
rect 17215 1143 17225 1215
rect 17245 1143 17255 1215
rect 17215 1130 17255 1143
rect 17505 1215 17545 1230
rect 17505 1195 17515 1215
rect 17535 1195 17545 1215
rect 17505 1165 17545 1195
rect 17505 1145 17515 1165
rect 17535 1145 17545 1165
rect 17505 1130 17545 1145
rect 17560 1215 17600 1230
rect 17560 1195 17570 1215
rect 17590 1195 17600 1215
rect 17560 1165 17600 1195
rect 17560 1145 17570 1165
rect 17590 1145 17600 1165
rect 17560 1130 17600 1145
rect 17615 1215 17655 1230
rect 17615 1195 17625 1215
rect 17645 1195 17655 1215
rect 17615 1165 17655 1195
rect 17615 1145 17625 1165
rect 17645 1145 17655 1165
rect 17615 1130 17655 1145
rect 17670 1215 17710 1230
rect 17670 1195 17680 1215
rect 17700 1195 17710 1215
rect 17670 1165 17710 1195
rect 17670 1145 17680 1165
rect 17700 1145 17710 1165
rect 17670 1130 17710 1145
rect 17725 1215 17765 1230
rect 17725 1195 17735 1215
rect 17755 1195 17765 1215
rect 17725 1165 17765 1195
rect 17725 1145 17735 1165
rect 17755 1145 17765 1165
rect 17725 1130 17765 1145
rect 17780 1215 17820 1230
rect 17780 1195 17790 1215
rect 17810 1195 17820 1215
rect 17780 1165 17820 1195
rect 17780 1145 17790 1165
rect 17810 1145 17820 1165
rect 17780 1130 17820 1145
rect 17835 1215 17875 1230
rect 17835 1195 17845 1215
rect 17865 1195 17875 1215
rect 17835 1165 17875 1195
rect 17835 1145 17845 1165
rect 17865 1145 17875 1165
rect 17835 1130 17875 1145
rect 17890 1215 17930 1230
rect 17890 1195 17900 1215
rect 17920 1195 17930 1215
rect 17890 1165 17930 1195
rect 17890 1145 17900 1165
rect 17920 1145 17930 1165
rect 17890 1130 17930 1145
rect 17945 1215 17985 1230
rect 17945 1195 17955 1215
rect 17975 1195 17985 1215
rect 17945 1165 17985 1195
rect 17945 1145 17955 1165
rect 17975 1145 17985 1165
rect 17945 1130 17985 1145
rect 18000 1215 18040 1230
rect 18000 1195 18010 1215
rect 18030 1195 18040 1215
rect 18000 1165 18040 1195
rect 18000 1145 18010 1165
rect 18030 1145 18040 1165
rect 18000 1130 18040 1145
rect 18055 1215 18095 1230
rect 18055 1195 18065 1215
rect 18085 1195 18095 1215
rect 18055 1165 18095 1195
rect 18055 1145 18065 1165
rect 18085 1145 18095 1165
rect 18055 1130 18095 1145
rect 18345 1215 18385 1230
rect 18345 1145 18355 1215
rect 18375 1145 18385 1215
rect 18345 1130 18385 1145
rect 18400 1215 18440 1230
rect 18400 1145 18410 1215
rect 18430 1145 18440 1215
rect 18400 1130 18440 1145
rect 18455 1215 18495 1230
rect 18455 1145 18465 1215
rect 18485 1145 18495 1215
rect 18455 1130 18495 1145
rect 18510 1215 18550 1230
rect 18510 1145 18520 1215
rect 18540 1145 18550 1215
rect 18510 1130 18550 1145
rect 18565 1215 18605 1230
rect 18565 1145 18575 1215
rect 18595 1145 18605 1215
rect 18565 1130 18605 1145
rect 18620 1215 18660 1230
rect 18620 1145 18630 1215
rect 18650 1145 18660 1215
rect 18620 1130 18660 1145
rect 18675 1215 18715 1230
rect 18675 1145 18685 1215
rect 18705 1145 18715 1215
rect 18675 1130 18715 1145
rect 16970 750 17010 765
rect 16970 730 16980 750
rect 17000 730 17010 750
rect 16970 700 17010 730
rect 16970 680 16980 700
rect 17000 680 17010 700
rect 16435 650 16475 665
rect 16435 630 16445 650
rect 16465 630 16475 650
rect 16435 600 16475 630
rect 16435 580 16445 600
rect 16465 580 16475 600
rect 16435 565 16475 580
rect 16490 650 16530 665
rect 16490 630 16500 650
rect 16520 630 16530 650
rect 16490 600 16530 630
rect 16490 580 16500 600
rect 16520 580 16530 600
rect 16490 565 16530 580
rect 16545 650 16585 665
rect 16545 630 16555 650
rect 16575 630 16585 650
rect 16545 600 16585 630
rect 16545 580 16555 600
rect 16575 580 16585 600
rect 16545 565 16585 580
rect 16600 650 16640 665
rect 16600 630 16610 650
rect 16630 630 16640 650
rect 16600 600 16640 630
rect 16600 580 16610 600
rect 16630 580 16640 600
rect 16600 565 16640 580
rect 16655 650 16700 665
rect 16655 630 16665 650
rect 16685 630 16700 650
rect 16655 600 16700 630
rect 16655 580 16665 600
rect 16685 580 16700 600
rect 16655 565 16700 580
rect 16970 650 17010 680
rect 16970 630 16980 650
rect 17000 630 17010 650
rect 16970 600 17010 630
rect 16970 580 16980 600
rect 17000 580 17010 600
rect 16970 550 17010 580
rect 16970 530 16980 550
rect 17000 530 17010 550
rect 16970 500 17010 530
rect 16970 480 16980 500
rect 17000 480 17010 500
rect 16970 465 17010 480
rect 17060 750 17100 765
rect 17060 730 17070 750
rect 17090 730 17100 750
rect 17060 700 17100 730
rect 17060 680 17070 700
rect 17090 680 17100 700
rect 17060 650 17100 680
rect 17060 630 17070 650
rect 17090 630 17100 650
rect 17060 600 17100 630
rect 17060 580 17070 600
rect 17090 580 17100 600
rect 17060 550 17100 580
rect 17060 530 17070 550
rect 17090 530 17100 550
rect 17060 500 17100 530
rect 17060 480 17070 500
rect 17090 480 17100 500
rect 17060 465 17100 480
rect 17150 750 17190 765
rect 17150 730 17160 750
rect 17180 730 17190 750
rect 17150 700 17190 730
rect 17150 680 17160 700
rect 17180 680 17190 700
rect 17150 650 17190 680
rect 17150 630 17160 650
rect 17180 630 17190 650
rect 17150 600 17190 630
rect 17150 580 17160 600
rect 17180 580 17190 600
rect 17150 550 17190 580
rect 17150 530 17160 550
rect 17180 530 17190 550
rect 17150 500 17190 530
rect 17150 480 17160 500
rect 17180 480 17190 500
rect 17150 465 17190 480
rect 17240 750 17280 765
rect 17240 730 17250 750
rect 17270 730 17280 750
rect 17240 700 17280 730
rect 17240 680 17250 700
rect 17270 680 17280 700
rect 17240 650 17280 680
rect 17240 630 17250 650
rect 17270 630 17280 650
rect 17240 600 17280 630
rect 17240 580 17250 600
rect 17270 580 17280 600
rect 17240 550 17280 580
rect 17240 530 17250 550
rect 17270 530 17280 550
rect 17240 500 17280 530
rect 17240 480 17250 500
rect 17270 480 17280 500
rect 17240 465 17280 480
rect 17330 750 17370 765
rect 17330 730 17340 750
rect 17360 730 17370 750
rect 17330 700 17370 730
rect 17330 680 17340 700
rect 17360 680 17370 700
rect 17330 650 17370 680
rect 17330 630 17340 650
rect 17360 630 17370 650
rect 17330 600 17370 630
rect 17330 580 17340 600
rect 17360 580 17370 600
rect 17330 550 17370 580
rect 17330 530 17340 550
rect 17360 530 17370 550
rect 17330 500 17370 530
rect 17330 480 17340 500
rect 17360 480 17370 500
rect 17330 465 17370 480
rect 17420 750 17460 765
rect 17420 730 17430 750
rect 17450 730 17460 750
rect 17420 700 17460 730
rect 17420 680 17430 700
rect 17450 680 17460 700
rect 17420 650 17460 680
rect 17420 630 17430 650
rect 17450 630 17460 650
rect 17420 600 17460 630
rect 17420 580 17430 600
rect 17450 580 17460 600
rect 17420 550 17460 580
rect 17420 530 17430 550
rect 17450 530 17460 550
rect 17420 500 17460 530
rect 17420 480 17430 500
rect 17450 480 17460 500
rect 17420 465 17460 480
rect 17510 750 17550 765
rect 17510 730 17520 750
rect 17540 730 17550 750
rect 17510 700 17550 730
rect 17510 680 17520 700
rect 17540 680 17550 700
rect 17510 650 17550 680
rect 17510 630 17520 650
rect 17540 630 17550 650
rect 17510 600 17550 630
rect 17510 580 17520 600
rect 17540 580 17550 600
rect 17510 550 17550 580
rect 17510 530 17520 550
rect 17540 530 17550 550
rect 17510 500 17550 530
rect 17510 480 17520 500
rect 17540 480 17550 500
rect 17510 465 17550 480
rect 17600 750 17640 765
rect 17600 730 17610 750
rect 17630 730 17640 750
rect 17600 700 17640 730
rect 17600 680 17610 700
rect 17630 680 17640 700
rect 17600 650 17640 680
rect 17600 630 17610 650
rect 17630 630 17640 650
rect 17600 600 17640 630
rect 17600 580 17610 600
rect 17630 580 17640 600
rect 17600 550 17640 580
rect 17600 530 17610 550
rect 17630 530 17640 550
rect 17600 500 17640 530
rect 17600 480 17610 500
rect 17630 480 17640 500
rect 17600 465 17640 480
rect 17690 750 17730 765
rect 17690 730 17700 750
rect 17720 730 17730 750
rect 17690 700 17730 730
rect 17690 680 17700 700
rect 17720 680 17730 700
rect 17690 650 17730 680
rect 17690 630 17700 650
rect 17720 630 17730 650
rect 17690 600 17730 630
rect 17690 580 17700 600
rect 17720 580 17730 600
rect 17690 550 17730 580
rect 17690 530 17700 550
rect 17720 530 17730 550
rect 17690 500 17730 530
rect 17690 480 17700 500
rect 17720 480 17730 500
rect 17690 465 17730 480
rect 17780 750 17820 765
rect 17780 730 17790 750
rect 17810 730 17820 750
rect 17780 700 17820 730
rect 17780 680 17790 700
rect 17810 680 17820 700
rect 17780 650 17820 680
rect 17780 630 17790 650
rect 17810 630 17820 650
rect 17780 600 17820 630
rect 17780 580 17790 600
rect 17810 580 17820 600
rect 17780 550 17820 580
rect 17780 530 17790 550
rect 17810 530 17820 550
rect 17780 500 17820 530
rect 17780 480 17790 500
rect 17810 480 17820 500
rect 17780 465 17820 480
rect 17870 750 17910 765
rect 17870 730 17880 750
rect 17900 730 17910 750
rect 17870 700 17910 730
rect 17870 680 17880 700
rect 17900 680 17910 700
rect 17870 650 17910 680
rect 17870 630 17880 650
rect 17900 630 17910 650
rect 17870 600 17910 630
rect 17870 580 17880 600
rect 17900 580 17910 600
rect 17870 550 17910 580
rect 17870 530 17880 550
rect 17900 530 17910 550
rect 17870 500 17910 530
rect 17870 480 17880 500
rect 17900 480 17910 500
rect 17870 465 17910 480
rect 17960 750 18000 765
rect 17960 730 17970 750
rect 17990 730 18000 750
rect 17960 700 18000 730
rect 17960 680 17970 700
rect 17990 680 18000 700
rect 17960 650 18000 680
rect 17960 630 17970 650
rect 17990 630 18000 650
rect 17960 600 18000 630
rect 17960 580 17970 600
rect 17990 580 18000 600
rect 17960 550 18000 580
rect 17960 530 17970 550
rect 17990 530 18000 550
rect 17960 500 18000 530
rect 17960 480 17970 500
rect 17990 480 18000 500
rect 17960 465 18000 480
rect 18050 750 18090 765
rect 18050 730 18060 750
rect 18080 730 18090 750
rect 18050 700 18090 730
rect 18050 680 18060 700
rect 18080 680 18090 700
rect 18050 650 18090 680
rect 18050 630 18060 650
rect 18080 630 18090 650
rect 18050 600 18090 630
rect 18050 580 18060 600
rect 18080 580 18090 600
rect 18050 550 18090 580
rect 18050 530 18060 550
rect 18080 530 18090 550
rect 18050 500 18090 530
rect 18050 480 18060 500
rect 18080 480 18090 500
rect 18050 465 18090 480
rect 18140 750 18180 765
rect 18140 730 18150 750
rect 18170 730 18180 750
rect 18140 700 18180 730
rect 18140 680 18150 700
rect 18170 680 18180 700
rect 18140 650 18180 680
rect 18140 630 18150 650
rect 18170 630 18180 650
rect 18140 600 18180 630
rect 18140 580 18150 600
rect 18170 580 18180 600
rect 18140 550 18180 580
rect 18140 530 18150 550
rect 18170 530 18180 550
rect 18140 500 18180 530
rect 18140 480 18150 500
rect 18170 480 18180 500
rect 18140 465 18180 480
rect 18230 750 18270 765
rect 18230 730 18240 750
rect 18260 730 18270 750
rect 18230 700 18270 730
rect 18230 680 18240 700
rect 18260 680 18270 700
rect 18230 650 18270 680
rect 18230 630 18240 650
rect 18260 630 18270 650
rect 18230 600 18270 630
rect 18230 580 18240 600
rect 18260 580 18270 600
rect 18230 550 18270 580
rect 18230 530 18240 550
rect 18260 530 18270 550
rect 18230 500 18270 530
rect 18230 480 18240 500
rect 18260 480 18270 500
rect 18230 465 18270 480
rect 18320 750 18360 765
rect 18320 730 18330 750
rect 18350 730 18360 750
rect 18320 700 18360 730
rect 18320 680 18330 700
rect 18350 680 18360 700
rect 18320 650 18360 680
rect 18320 630 18330 650
rect 18350 630 18360 650
rect 18320 600 18360 630
rect 18320 580 18330 600
rect 18350 580 18360 600
rect 18320 550 18360 580
rect 18320 530 18330 550
rect 18350 530 18360 550
rect 18320 500 18360 530
rect 18320 480 18330 500
rect 18350 480 18360 500
rect 18320 465 18360 480
rect 18410 750 18450 765
rect 18410 730 18420 750
rect 18440 730 18450 750
rect 18410 700 18450 730
rect 18410 680 18420 700
rect 18440 680 18450 700
rect 18410 650 18450 680
rect 18410 630 18420 650
rect 18440 630 18450 650
rect 18410 600 18450 630
rect 18410 580 18420 600
rect 18440 580 18450 600
rect 18410 550 18450 580
rect 18410 530 18420 550
rect 18440 530 18450 550
rect 18410 500 18450 530
rect 18410 480 18420 500
rect 18440 480 18450 500
rect 18410 465 18450 480
rect 18500 750 18540 765
rect 18500 730 18510 750
rect 18530 730 18540 750
rect 18500 700 18540 730
rect 18500 680 18510 700
rect 18530 680 18540 700
rect 18500 650 18540 680
rect 18500 630 18510 650
rect 18530 630 18540 650
rect 18500 600 18540 630
rect 18500 580 18510 600
rect 18530 580 18540 600
rect 18500 550 18540 580
rect 18500 530 18510 550
rect 18530 530 18540 550
rect 18500 500 18540 530
rect 18500 480 18510 500
rect 18530 480 18540 500
rect 18500 465 18540 480
rect 18590 750 18630 765
rect 18590 730 18600 750
rect 18620 730 18630 750
rect 18590 700 18630 730
rect 18590 680 18600 700
rect 18620 680 18630 700
rect 18590 650 18630 680
rect 18590 630 18600 650
rect 18620 630 18630 650
rect 18590 600 18630 630
rect 18590 580 18600 600
rect 18620 580 18630 600
rect 18590 550 18630 580
rect 18905 750 18945 765
rect 18905 730 18915 750
rect 18935 730 18945 750
rect 18905 700 18945 730
rect 18905 680 18915 700
rect 18935 680 18945 700
rect 18905 650 18945 680
rect 18905 630 18915 650
rect 18935 630 18945 650
rect 18905 600 18945 630
rect 18905 580 18915 600
rect 18935 580 18945 600
rect 18905 565 18945 580
rect 18960 750 19000 765
rect 18960 730 18970 750
rect 18990 730 19000 750
rect 18960 700 19000 730
rect 18960 680 18970 700
rect 18990 680 19000 700
rect 18960 650 19000 680
rect 18960 630 18970 650
rect 18990 630 19000 650
rect 18960 600 19000 630
rect 18960 580 18970 600
rect 18990 580 19000 600
rect 18960 565 19000 580
rect 19015 750 19055 765
rect 19015 730 19025 750
rect 19045 730 19055 750
rect 19015 700 19055 730
rect 19015 680 19025 700
rect 19045 680 19055 700
rect 19015 650 19055 680
rect 19015 630 19025 650
rect 19045 630 19055 650
rect 19015 600 19055 630
rect 19015 580 19025 600
rect 19045 580 19055 600
rect 19015 565 19055 580
rect 19070 750 19110 765
rect 19070 730 19080 750
rect 19100 730 19110 750
rect 19070 700 19110 730
rect 19070 680 19080 700
rect 19100 680 19110 700
rect 19070 650 19110 680
rect 19070 630 19080 650
rect 19100 630 19110 650
rect 19070 600 19110 630
rect 19070 580 19080 600
rect 19100 580 19110 600
rect 19070 565 19110 580
rect 18590 530 18600 550
rect 18620 530 18630 550
rect 18590 500 18630 530
rect 18590 480 18600 500
rect 18620 480 18630 500
rect 18590 465 18630 480
rect 16420 -90 16460 -75
rect 16420 -110 16430 -90
rect 16450 -110 16460 -90
rect 16420 -140 16460 -110
rect 16420 -160 16430 -140
rect 16450 -160 16460 -140
rect 16420 -175 16460 -160
rect 16480 -90 16520 -75
rect 16480 -110 16490 -90
rect 16510 -110 16520 -90
rect 16480 -140 16520 -110
rect 16480 -160 16490 -140
rect 16510 -160 16520 -140
rect 16480 -175 16520 -160
rect 16540 -90 16580 -75
rect 16540 -110 16550 -90
rect 16570 -110 16580 -90
rect 16540 -140 16580 -110
rect 16540 -160 16550 -140
rect 16570 -160 16580 -140
rect 16540 -175 16580 -160
rect 16600 -90 16640 -75
rect 16600 -110 16610 -90
rect 16630 -110 16640 -90
rect 16600 -140 16640 -110
rect 16600 -160 16610 -140
rect 16630 -160 16640 -140
rect 16600 -175 16640 -160
rect 16660 -90 16700 -75
rect 16660 -110 16670 -90
rect 16690 -110 16700 -90
rect 16660 -140 16700 -110
rect 16660 -160 16670 -140
rect 16690 -160 16700 -140
rect 16660 -175 16700 -160
rect 16720 -90 16760 -75
rect 16720 -110 16730 -90
rect 16750 -110 16760 -90
rect 16720 -140 16760 -110
rect 16720 -160 16730 -140
rect 16750 -160 16760 -140
rect 16720 -175 16760 -160
rect 16780 -90 16820 -75
rect 16780 -110 16790 -90
rect 16810 -110 16820 -90
rect 16780 -140 16820 -110
rect 16780 -160 16790 -140
rect 16810 -160 16820 -140
rect 16780 -175 16820 -160
rect 16840 -90 16880 -75
rect 16840 -110 16850 -90
rect 16870 -110 16880 -90
rect 16840 -140 16880 -110
rect 16840 -160 16850 -140
rect 16870 -160 16880 -140
rect 16840 -175 16880 -160
rect 16900 -90 16940 -75
rect 16900 -110 16910 -90
rect 16930 -110 16940 -90
rect 16900 -140 16940 -110
rect 16900 -160 16910 -140
rect 16930 -160 16940 -140
rect 16900 -175 16940 -160
rect 16960 -90 17000 -75
rect 16960 -110 16970 -90
rect 16990 -110 17000 -90
rect 16960 -140 17000 -110
rect 16960 -160 16970 -140
rect 16990 -160 17000 -140
rect 16960 -175 17000 -160
rect 17020 -90 17060 -75
rect 17020 -110 17030 -90
rect 17050 -110 17060 -90
rect 17020 -140 17060 -110
rect 17020 -160 17030 -140
rect 17050 -160 17060 -140
rect 17020 -175 17060 -160
rect 17080 -90 17120 -75
rect 17080 -110 17090 -90
rect 17110 -110 17120 -90
rect 17080 -140 17120 -110
rect 17080 -160 17090 -140
rect 17110 -160 17120 -140
rect 17080 -175 17120 -160
rect 17140 -90 17180 -75
rect 17140 -110 17150 -90
rect 17170 -110 17180 -90
rect 17140 -140 17180 -110
rect 17140 -160 17150 -140
rect 17170 -160 17180 -140
rect 17140 -175 17180 -160
rect 17200 -90 17240 -75
rect 17200 -110 17210 -90
rect 17230 -110 17240 -90
rect 17200 -140 17240 -110
rect 17200 -160 17210 -140
rect 17230 -160 17240 -140
rect 17200 -175 17240 -160
rect 17260 -90 17300 -75
rect 17260 -110 17270 -90
rect 17290 -110 17300 -90
rect 17260 -140 17300 -110
rect 17260 -160 17270 -140
rect 17290 -160 17300 -140
rect 17260 -175 17300 -160
rect 17320 -90 17360 -75
rect 17320 -110 17330 -90
rect 17350 -110 17360 -90
rect 17320 -140 17360 -110
rect 17320 -160 17330 -140
rect 17350 -160 17360 -140
rect 17320 -175 17360 -160
rect 17380 -90 17420 -75
rect 17380 -110 17390 -90
rect 17410 -110 17420 -90
rect 17380 -140 17420 -110
rect 17380 -160 17390 -140
rect 17410 -160 17420 -140
rect 17380 -175 17420 -160
rect 17440 -90 17480 -75
rect 17440 -110 17450 -90
rect 17470 -110 17480 -90
rect 17440 -140 17480 -110
rect 17440 -160 17450 -140
rect 17470 -160 17480 -140
rect 17440 -175 17480 -160
rect 17500 -90 17540 -75
rect 17500 -110 17510 -90
rect 17530 -110 17540 -90
rect 17500 -140 17540 -110
rect 17500 -160 17510 -140
rect 17530 -160 17540 -140
rect 17500 -175 17540 -160
rect 17560 -90 17600 -75
rect 17560 -110 17570 -90
rect 17590 -110 17600 -90
rect 17560 -140 17600 -110
rect 17560 -160 17570 -140
rect 17590 -160 17600 -140
rect 17560 -175 17600 -160
rect 17620 -90 17660 -75
rect 17620 -110 17630 -90
rect 17650 -110 17660 -90
rect 17620 -140 17660 -110
rect 17620 -160 17630 -140
rect 17650 -160 17660 -140
rect 17620 -175 17660 -160
rect 17940 -90 17980 -75
rect 17940 -110 17950 -90
rect 17970 -110 17980 -90
rect 17940 -140 17980 -110
rect 17940 -160 17950 -140
rect 17970 -160 17980 -140
rect 17940 -175 17980 -160
rect 18000 -90 18040 -75
rect 18000 -110 18010 -90
rect 18030 -110 18040 -90
rect 18000 -140 18040 -110
rect 18000 -160 18010 -140
rect 18030 -160 18040 -140
rect 18000 -175 18040 -160
rect 18060 -90 18100 -75
rect 18060 -110 18070 -90
rect 18090 -110 18100 -90
rect 18060 -140 18100 -110
rect 18060 -160 18070 -140
rect 18090 -160 18100 -140
rect 18060 -175 18100 -160
rect 18120 -90 18160 -75
rect 18120 -110 18130 -90
rect 18150 -110 18160 -90
rect 18120 -140 18160 -110
rect 18120 -160 18130 -140
rect 18150 -160 18160 -140
rect 18120 -175 18160 -160
rect 18180 -90 18220 -75
rect 18180 -110 18190 -90
rect 18210 -110 18220 -90
rect 18180 -140 18220 -110
rect 18180 -160 18190 -140
rect 18210 -160 18220 -140
rect 18180 -175 18220 -160
rect 18240 -90 18280 -75
rect 18240 -110 18250 -90
rect 18270 -110 18280 -90
rect 18240 -140 18280 -110
rect 18240 -160 18250 -140
rect 18270 -160 18280 -140
rect 18240 -175 18280 -160
rect 18300 -90 18340 -75
rect 18300 -110 18310 -90
rect 18330 -110 18340 -90
rect 18300 -140 18340 -110
rect 18300 -160 18310 -140
rect 18330 -160 18340 -140
rect 18300 -175 18340 -160
rect 18360 -90 18400 -75
rect 18360 -110 18370 -90
rect 18390 -110 18400 -90
rect 18360 -140 18400 -110
rect 18360 -160 18370 -140
rect 18390 -160 18400 -140
rect 18360 -175 18400 -160
rect 18420 -90 18460 -75
rect 18420 -110 18430 -90
rect 18450 -110 18460 -90
rect 18420 -140 18460 -110
rect 18420 -160 18430 -140
rect 18450 -160 18460 -140
rect 18420 -175 18460 -160
rect 18480 -90 18520 -75
rect 18480 -110 18490 -90
rect 18510 -110 18520 -90
rect 18480 -140 18520 -110
rect 18480 -160 18490 -140
rect 18510 -160 18520 -140
rect 18480 -175 18520 -160
rect 18540 -90 18580 -75
rect 18540 -110 18550 -90
rect 18570 -110 18580 -90
rect 18540 -140 18580 -110
rect 18540 -160 18550 -140
rect 18570 -160 18580 -140
rect 18540 -175 18580 -160
rect 18600 -90 18640 -75
rect 18600 -110 18610 -90
rect 18630 -110 18640 -90
rect 18600 -140 18640 -110
rect 18600 -160 18610 -140
rect 18630 -160 18640 -140
rect 18600 -175 18640 -160
rect 18660 -90 18700 -75
rect 18660 -110 18670 -90
rect 18690 -110 18700 -90
rect 18660 -140 18700 -110
rect 18660 -160 18670 -140
rect 18690 -160 18700 -140
rect 18660 -175 18700 -160
rect 18720 -90 18760 -75
rect 18720 -110 18730 -90
rect 18750 -110 18760 -90
rect 18720 -140 18760 -110
rect 18720 -160 18730 -140
rect 18750 -160 18760 -140
rect 18720 -175 18760 -160
rect 18780 -90 18820 -75
rect 18780 -110 18790 -90
rect 18810 -110 18820 -90
rect 18780 -140 18820 -110
rect 18780 -160 18790 -140
rect 18810 -160 18820 -140
rect 18780 -175 18820 -160
rect 18840 -90 18880 -75
rect 18840 -110 18850 -90
rect 18870 -110 18880 -90
rect 18840 -140 18880 -110
rect 18840 -160 18850 -140
rect 18870 -160 18880 -140
rect 18840 -175 18880 -160
rect 18900 -90 18940 -75
rect 18900 -110 18910 -90
rect 18930 -110 18940 -90
rect 18900 -140 18940 -110
rect 18900 -160 18910 -140
rect 18930 -160 18940 -140
rect 18900 -175 18940 -160
rect 18960 -90 19000 -75
rect 18960 -110 18970 -90
rect 18990 -110 19000 -90
rect 18960 -140 19000 -110
rect 18960 -160 18970 -140
rect 18990 -160 19000 -140
rect 18960 -175 19000 -160
rect 19020 -90 19060 -75
rect 19020 -110 19030 -90
rect 19050 -110 19060 -90
rect 19020 -140 19060 -110
rect 19020 -160 19030 -140
rect 19050 -160 19060 -140
rect 19020 -175 19060 -160
rect 19080 -90 19120 -75
rect 19080 -110 19090 -90
rect 19110 -110 19120 -90
rect 19080 -140 19120 -110
rect 19080 -160 19090 -140
rect 19110 -160 19120 -140
rect 19080 -175 19120 -160
rect 19140 -90 19180 -75
rect 19140 -110 19150 -90
rect 19170 -110 19180 -90
rect 19140 -140 19180 -110
rect 19140 -160 19150 -140
rect 19170 -160 19180 -140
rect 19140 -175 19180 -160
<< ndiffc >>
rect 16970 -395 16990 -375
rect 16970 -445 16990 -425
rect 16970 -495 16990 -475
rect 16970 -545 16990 -525
rect 16970 -595 16990 -575
rect 17030 -395 17050 -375
rect 17030 -445 17050 -425
rect 17030 -495 17050 -475
rect 17030 -545 17050 -525
rect 17030 -595 17050 -575
rect 17090 -395 17110 -375
rect 18490 -395 18510 -375
rect 17090 -445 17110 -425
rect 17090 -495 17110 -475
rect 17090 -545 17110 -525
rect 17090 -595 17110 -575
rect 18490 -445 18510 -425
rect 18490 -495 18510 -475
rect 18490 -545 18510 -525
rect 18490 -595 18510 -575
rect 18550 -395 18570 -375
rect 18550 -445 18570 -425
rect 18550 -495 18570 -475
rect 18550 -545 18570 -525
rect 18550 -595 18570 -575
rect 18610 -395 18630 -375
rect 18610 -445 18630 -425
rect 18610 -495 18630 -475
rect 18610 -545 18630 -525
rect 18610 -595 18630 -575
rect 16540 -845 16560 -825
rect 16540 -895 16560 -875
rect 16540 -945 16560 -925
rect 16540 -995 16560 -975
rect 16540 -1045 16560 -1025
rect 17080 -845 17100 -825
rect 17160 -845 17180 -825
rect 17080 -895 17100 -875
rect 17160 -895 17180 -875
rect 17080 -945 17100 -925
rect 17160 -945 17180 -925
rect 17080 -995 17100 -975
rect 17160 -995 17180 -975
rect 17080 -1045 17100 -1025
rect 17160 -1045 17180 -1025
rect 17700 -845 17720 -825
rect 17700 -895 17720 -875
rect 17700 -945 17720 -925
rect 17700 -995 17720 -975
rect 17700 -1045 17720 -1025
rect 17880 -845 17900 -825
rect 17880 -895 17900 -875
rect 17880 -945 17900 -925
rect 17880 -995 17900 -975
rect 17880 -1045 17900 -1025
rect 18420 -845 18440 -825
rect 18500 -845 18520 -825
rect 18420 -895 18440 -875
rect 18500 -895 18520 -875
rect 18420 -945 18440 -925
rect 18500 -945 18520 -925
rect 18420 -995 18440 -975
rect 18500 -995 18520 -975
rect 18420 -1045 18440 -1025
rect 18500 -1045 18520 -1025
rect 19040 -845 19060 -825
rect 19040 -895 19060 -875
rect 19040 -945 19060 -925
rect 19040 -995 19060 -975
rect 19040 -1045 19060 -1025
rect 16750 -1225 16770 -1205
rect 16750 -1275 16770 -1255
rect 17790 -1225 17810 -1205
rect 17790 -1275 17810 -1255
rect 18830 -1225 18850 -1205
rect 18830 -1275 18850 -1255
rect 16550 -1575 16570 -1555
rect 16550 -1625 16570 -1605
rect 16605 -1575 16625 -1555
rect 16605 -1625 16625 -1605
rect 16660 -1575 16680 -1555
rect 16660 -1625 16680 -1605
rect 16715 -1575 16735 -1555
rect 16715 -1625 16735 -1605
rect 16770 -1575 16790 -1555
rect 16770 -1625 16790 -1605
rect 16825 -1575 16845 -1555
rect 16825 -1625 16845 -1605
rect 17035 -1575 17055 -1555
rect 17035 -1625 17055 -1605
rect 17090 -1575 17110 -1555
rect 17090 -1625 17110 -1605
rect 17145 -1575 17165 -1555
rect 17145 -1625 17165 -1605
rect 17200 -1575 17220 -1555
rect 17200 -1625 17220 -1605
rect 17255 -1575 17275 -1555
rect 17255 -1625 17275 -1605
rect 17310 -1575 17330 -1555
rect 17310 -1625 17330 -1605
rect 17365 -1575 17385 -1555
rect 17365 -1625 17385 -1605
rect 17420 -1575 17440 -1555
rect 17420 -1625 17440 -1605
rect 17475 -1575 17495 -1555
rect 17475 -1625 17495 -1605
rect 17625 -1575 17645 -1555
rect 17625 -1625 17645 -1605
rect 17680 -1575 17700 -1555
rect 17680 -1625 17700 -1605
rect 17735 -1575 17755 -1555
rect 17735 -1625 17755 -1605
rect 17790 -1575 17810 -1555
rect 17790 -1625 17810 -1605
rect 17845 -1575 17865 -1555
rect 17845 -1625 17865 -1605
rect 17900 -1575 17920 -1555
rect 17900 -1625 17920 -1605
rect 17955 -1575 17975 -1555
rect 17955 -1625 17975 -1605
rect 18105 -1575 18125 -1555
rect 18105 -1625 18125 -1605
rect 18160 -1575 18180 -1555
rect 18160 -1625 18180 -1605
rect 18215 -1575 18235 -1555
rect 18215 -1625 18235 -1605
rect 18270 -1575 18290 -1555
rect 18270 -1625 18290 -1605
rect 18325 -1575 18345 -1555
rect 18325 -1625 18345 -1605
rect 18380 -1575 18400 -1555
rect 18380 -1625 18400 -1605
rect 18435 -1575 18455 -1555
rect 18435 -1625 18455 -1605
rect 18490 -1575 18510 -1555
rect 18490 -1625 18510 -1605
rect 18545 -1575 18565 -1555
rect 18545 -1625 18565 -1605
<< pdiffc >>
rect 16385 1195 16405 1215
rect 16385 1145 16405 1165
rect 16440 1195 16460 1215
rect 16440 1145 16460 1165
rect 16495 1195 16515 1215
rect 16495 1145 16515 1165
rect 16550 1195 16570 1215
rect 16550 1145 16570 1165
rect 16605 1195 16625 1215
rect 16605 1145 16625 1165
rect 16895 1143 16915 1215
rect 16950 1143 16970 1215
rect 17005 1143 17025 1215
rect 17060 1143 17080 1215
rect 17115 1143 17135 1215
rect 17170 1143 17190 1215
rect 17225 1143 17245 1215
rect 17515 1195 17535 1215
rect 17515 1145 17535 1165
rect 17570 1195 17590 1215
rect 17570 1145 17590 1165
rect 17625 1195 17645 1215
rect 17625 1145 17645 1165
rect 17680 1195 17700 1215
rect 17680 1145 17700 1165
rect 17735 1195 17755 1215
rect 17735 1145 17755 1165
rect 17790 1195 17810 1215
rect 17790 1145 17810 1165
rect 17845 1195 17865 1215
rect 17845 1145 17865 1165
rect 17900 1195 17920 1215
rect 17900 1145 17920 1165
rect 17955 1195 17975 1215
rect 17955 1145 17975 1165
rect 18010 1195 18030 1215
rect 18010 1145 18030 1165
rect 18065 1195 18085 1215
rect 18065 1145 18085 1165
rect 18355 1145 18375 1215
rect 18410 1145 18430 1215
rect 18465 1145 18485 1215
rect 18520 1145 18540 1215
rect 18575 1145 18595 1215
rect 18630 1145 18650 1215
rect 18685 1145 18705 1215
rect 16980 730 17000 750
rect 16980 680 17000 700
rect 16445 630 16465 650
rect 16445 580 16465 600
rect 16500 630 16520 650
rect 16500 580 16520 600
rect 16555 630 16575 650
rect 16555 580 16575 600
rect 16610 630 16630 650
rect 16610 580 16630 600
rect 16665 630 16685 650
rect 16665 580 16685 600
rect 16980 630 17000 650
rect 16980 580 17000 600
rect 16980 530 17000 550
rect 16980 480 17000 500
rect 17070 730 17090 750
rect 17070 680 17090 700
rect 17070 630 17090 650
rect 17070 580 17090 600
rect 17070 530 17090 550
rect 17070 480 17090 500
rect 17160 730 17180 750
rect 17160 680 17180 700
rect 17160 630 17180 650
rect 17160 580 17180 600
rect 17160 530 17180 550
rect 17160 480 17180 500
rect 17250 730 17270 750
rect 17250 680 17270 700
rect 17250 630 17270 650
rect 17250 580 17270 600
rect 17250 530 17270 550
rect 17250 480 17270 500
rect 17340 730 17360 750
rect 17340 680 17360 700
rect 17340 630 17360 650
rect 17340 580 17360 600
rect 17340 530 17360 550
rect 17340 480 17360 500
rect 17430 730 17450 750
rect 17430 680 17450 700
rect 17430 630 17450 650
rect 17430 580 17450 600
rect 17430 530 17450 550
rect 17430 480 17450 500
rect 17520 730 17540 750
rect 17520 680 17540 700
rect 17520 630 17540 650
rect 17520 580 17540 600
rect 17520 530 17540 550
rect 17520 480 17540 500
rect 17610 730 17630 750
rect 17610 680 17630 700
rect 17610 630 17630 650
rect 17610 580 17630 600
rect 17610 530 17630 550
rect 17610 480 17630 500
rect 17700 730 17720 750
rect 17700 680 17720 700
rect 17700 630 17720 650
rect 17700 580 17720 600
rect 17700 530 17720 550
rect 17700 480 17720 500
rect 17790 730 17810 750
rect 17790 680 17810 700
rect 17790 630 17810 650
rect 17790 580 17810 600
rect 17790 530 17810 550
rect 17790 480 17810 500
rect 17880 730 17900 750
rect 17880 680 17900 700
rect 17880 630 17900 650
rect 17880 580 17900 600
rect 17880 530 17900 550
rect 17880 480 17900 500
rect 17970 730 17990 750
rect 17970 680 17990 700
rect 17970 630 17990 650
rect 17970 580 17990 600
rect 17970 530 17990 550
rect 17970 480 17990 500
rect 18060 730 18080 750
rect 18060 680 18080 700
rect 18060 630 18080 650
rect 18060 580 18080 600
rect 18060 530 18080 550
rect 18060 480 18080 500
rect 18150 730 18170 750
rect 18150 680 18170 700
rect 18150 630 18170 650
rect 18150 580 18170 600
rect 18150 530 18170 550
rect 18150 480 18170 500
rect 18240 730 18260 750
rect 18240 680 18260 700
rect 18240 630 18260 650
rect 18240 580 18260 600
rect 18240 530 18260 550
rect 18240 480 18260 500
rect 18330 730 18350 750
rect 18330 680 18350 700
rect 18330 630 18350 650
rect 18330 580 18350 600
rect 18330 530 18350 550
rect 18330 480 18350 500
rect 18420 730 18440 750
rect 18420 680 18440 700
rect 18420 630 18440 650
rect 18420 580 18440 600
rect 18420 530 18440 550
rect 18420 480 18440 500
rect 18510 730 18530 750
rect 18510 680 18530 700
rect 18510 630 18530 650
rect 18510 580 18530 600
rect 18510 530 18530 550
rect 18510 480 18530 500
rect 18600 730 18620 750
rect 18600 680 18620 700
rect 18600 630 18620 650
rect 18600 580 18620 600
rect 18915 730 18935 750
rect 18915 680 18935 700
rect 18915 630 18935 650
rect 18915 580 18935 600
rect 18970 730 18990 750
rect 18970 680 18990 700
rect 18970 630 18990 650
rect 18970 580 18990 600
rect 19025 730 19045 750
rect 19025 680 19045 700
rect 19025 630 19045 650
rect 19025 580 19045 600
rect 19080 730 19100 750
rect 19080 680 19100 700
rect 19080 630 19100 650
rect 19080 580 19100 600
rect 18600 530 18620 550
rect 18600 480 18620 500
rect 16430 -110 16450 -90
rect 16430 -160 16450 -140
rect 16490 -110 16510 -90
rect 16490 -160 16510 -140
rect 16550 -110 16570 -90
rect 16550 -160 16570 -140
rect 16610 -110 16630 -90
rect 16610 -160 16630 -140
rect 16670 -110 16690 -90
rect 16670 -160 16690 -140
rect 16730 -110 16750 -90
rect 16730 -160 16750 -140
rect 16790 -110 16810 -90
rect 16790 -160 16810 -140
rect 16850 -110 16870 -90
rect 16850 -160 16870 -140
rect 16910 -110 16930 -90
rect 16910 -160 16930 -140
rect 16970 -110 16990 -90
rect 16970 -160 16990 -140
rect 17030 -110 17050 -90
rect 17030 -160 17050 -140
rect 17090 -110 17110 -90
rect 17090 -160 17110 -140
rect 17150 -110 17170 -90
rect 17150 -160 17170 -140
rect 17210 -110 17230 -90
rect 17210 -160 17230 -140
rect 17270 -110 17290 -90
rect 17270 -160 17290 -140
rect 17330 -110 17350 -90
rect 17330 -160 17350 -140
rect 17390 -110 17410 -90
rect 17390 -160 17410 -140
rect 17450 -110 17470 -90
rect 17450 -160 17470 -140
rect 17510 -110 17530 -90
rect 17510 -160 17530 -140
rect 17570 -110 17590 -90
rect 17570 -160 17590 -140
rect 17630 -110 17650 -90
rect 17630 -160 17650 -140
rect 17950 -110 17970 -90
rect 17950 -160 17970 -140
rect 18010 -110 18030 -90
rect 18010 -160 18030 -140
rect 18070 -110 18090 -90
rect 18070 -160 18090 -140
rect 18130 -110 18150 -90
rect 18130 -160 18150 -140
rect 18190 -110 18210 -90
rect 18190 -160 18210 -140
rect 18250 -110 18270 -90
rect 18250 -160 18270 -140
rect 18310 -110 18330 -90
rect 18310 -160 18330 -140
rect 18370 -110 18390 -90
rect 18370 -160 18390 -140
rect 18430 -110 18450 -90
rect 18430 -160 18450 -140
rect 18490 -110 18510 -90
rect 18490 -160 18510 -140
rect 18550 -110 18570 -90
rect 18550 -160 18570 -140
rect 18610 -110 18630 -90
rect 18610 -160 18630 -140
rect 18670 -110 18690 -90
rect 18670 -160 18690 -140
rect 18730 -110 18750 -90
rect 18730 -160 18750 -140
rect 18790 -110 18810 -90
rect 18790 -160 18810 -140
rect 18850 -110 18870 -90
rect 18850 -160 18870 -140
rect 18910 -110 18930 -90
rect 18910 -160 18930 -140
rect 18970 -110 18990 -90
rect 18970 -160 18990 -140
rect 19030 -110 19050 -90
rect 19030 -160 19050 -140
rect 19090 -110 19110 -90
rect 19090 -160 19110 -140
rect 19150 -110 19170 -90
rect 19150 -160 19170 -140
<< psubdiff >>
rect 17560 -375 17600 -360
rect 17560 -395 17570 -375
rect 17590 -395 17600 -375
rect 17560 -410 17600 -395
rect 18000 -375 18040 -360
rect 18000 -395 18010 -375
rect 18030 -395 18040 -375
rect 18000 -410 18040 -395
rect 17110 -825 17150 -810
rect 17110 -845 17120 -825
rect 17140 -845 17150 -825
rect 17110 -875 17150 -845
rect 17110 -895 17120 -875
rect 17140 -895 17150 -875
rect 17110 -925 17150 -895
rect 17110 -945 17120 -925
rect 17140 -945 17150 -925
rect 17110 -975 17150 -945
rect 17110 -995 17120 -975
rect 17140 -995 17150 -975
rect 17110 -1025 17150 -995
rect 17110 -1045 17120 -1025
rect 17140 -1045 17150 -1025
rect 17110 -1055 17150 -1045
rect 18450 -825 18490 -810
rect 18450 -845 18460 -825
rect 18480 -845 18490 -825
rect 18450 -875 18490 -845
rect 18450 -895 18460 -875
rect 18480 -895 18490 -875
rect 18450 -925 18490 -895
rect 18450 -945 18460 -925
rect 18480 -945 18490 -925
rect 18450 -975 18490 -945
rect 18450 -995 18460 -975
rect 18480 -995 18490 -975
rect 18450 -1025 18490 -995
rect 18450 -1045 18460 -1025
rect 18480 -1045 18490 -1025
rect 18450 -1060 18490 -1045
rect 18860 -1205 18900 -1190
rect 18860 -1225 18870 -1205
rect 18890 -1225 18900 -1205
rect 18860 -1255 18900 -1225
rect 18860 -1275 18870 -1255
rect 18890 -1275 18900 -1255
rect 18860 -1290 18900 -1275
rect 16500 -1555 16540 -1540
rect 16500 -1575 16510 -1555
rect 16530 -1575 16540 -1555
rect 16500 -1605 16540 -1575
rect 16500 -1625 16510 -1605
rect 16530 -1625 16540 -1605
rect 16500 -1640 16540 -1625
rect 16855 -1555 16895 -1540
rect 16855 -1575 16865 -1555
rect 16885 -1575 16895 -1555
rect 16855 -1605 16895 -1575
rect 16855 -1625 16865 -1605
rect 16885 -1625 16895 -1605
rect 16855 -1640 16895 -1625
rect 16985 -1555 17025 -1540
rect 16985 -1575 16995 -1555
rect 17015 -1575 17025 -1555
rect 16985 -1605 17025 -1575
rect 16985 -1625 16995 -1605
rect 17015 -1625 17025 -1605
rect 16985 -1640 17025 -1625
rect 17505 -1555 17545 -1540
rect 17505 -1575 17515 -1555
rect 17535 -1575 17545 -1555
rect 17505 -1605 17545 -1575
rect 17505 -1625 17515 -1605
rect 17535 -1625 17545 -1605
rect 17505 -1640 17545 -1625
rect 17575 -1555 17615 -1540
rect 17575 -1575 17585 -1555
rect 17605 -1575 17615 -1555
rect 17575 -1605 17615 -1575
rect 17575 -1625 17585 -1605
rect 17605 -1625 17615 -1605
rect 17575 -1640 17615 -1625
rect 17985 -1555 18025 -1540
rect 17985 -1575 17995 -1555
rect 18015 -1575 18025 -1555
rect 17985 -1605 18025 -1575
rect 17985 -1625 17995 -1605
rect 18015 -1625 18025 -1605
rect 17985 -1640 18025 -1625
rect 18055 -1555 18095 -1540
rect 18055 -1575 18065 -1555
rect 18085 -1575 18095 -1555
rect 18055 -1605 18095 -1575
rect 18055 -1625 18065 -1605
rect 18085 -1625 18095 -1605
rect 18055 -1640 18095 -1625
rect 18575 -1555 18615 -1540
rect 18575 -1575 18585 -1555
rect 18605 -1575 18615 -1555
rect 18575 -1605 18615 -1575
rect 18575 -1625 18585 -1605
rect 18605 -1625 18615 -1605
rect 18575 -1640 18615 -1625
rect 17775 -4170 17825 -4155
rect 17775 -4190 17790 -4170
rect 17810 -4190 17825 -4170
rect 17775 -4220 17825 -4190
rect 17775 -4240 17790 -4220
rect 17810 -4240 17825 -4220
rect 17775 -4270 17825 -4240
rect 17775 -4290 17790 -4270
rect 17810 -4290 17825 -4270
rect 17775 -4305 17825 -4290
<< nsubdiff >>
rect 16335 1217 16375 1230
rect 16335 1195 16345 1217
rect 16365 1195 16375 1217
rect 16335 1165 16375 1195
rect 16335 1145 16345 1165
rect 16365 1145 16375 1165
rect 16335 1130 16375 1145
rect 16635 1217 16675 1230
rect 16635 1195 16645 1217
rect 16665 1195 16675 1217
rect 16635 1165 16675 1195
rect 16635 1145 16645 1165
rect 16665 1145 16675 1165
rect 16635 1130 16675 1145
rect 16845 1217 16885 1230
rect 16845 1145 16855 1217
rect 16875 1145 16885 1217
rect 16845 1130 16885 1145
rect 17255 1217 17295 1230
rect 17255 1145 17265 1217
rect 17285 1145 17295 1217
rect 17255 1130 17295 1145
rect 17465 1217 17505 1230
rect 17465 1195 17475 1217
rect 17495 1195 17505 1217
rect 17465 1165 17505 1195
rect 17465 1145 17475 1165
rect 17495 1145 17505 1165
rect 17465 1130 17505 1145
rect 18095 1217 18135 1230
rect 18095 1195 18105 1217
rect 18125 1195 18135 1217
rect 18095 1165 18135 1195
rect 18095 1145 18105 1165
rect 18125 1145 18135 1165
rect 18095 1130 18135 1145
rect 18305 1217 18345 1230
rect 18305 1145 18315 1217
rect 18335 1145 18345 1217
rect 18305 1130 18345 1145
rect 18715 1217 18755 1230
rect 18715 1145 18725 1217
rect 18745 1145 18755 1217
rect 18715 1130 18755 1145
rect 16930 750 16970 765
rect 16930 730 16940 750
rect 16960 730 16970 750
rect 16930 700 16970 730
rect 16930 680 16940 700
rect 16960 680 16970 700
rect 16395 650 16435 665
rect 16395 630 16405 650
rect 16425 630 16435 650
rect 16395 600 16435 630
rect 16395 580 16405 600
rect 16425 580 16435 600
rect 16395 565 16435 580
rect 16700 650 16740 665
rect 16700 630 16710 650
rect 16730 630 16740 650
rect 16700 600 16740 630
rect 16700 580 16710 600
rect 16730 580 16740 600
rect 16700 565 16740 580
rect 16930 650 16970 680
rect 16930 630 16940 650
rect 16960 630 16970 650
rect 16930 600 16970 630
rect 16930 580 16940 600
rect 16960 580 16970 600
rect 16930 550 16970 580
rect 16930 530 16940 550
rect 16960 530 16970 550
rect 16930 500 16970 530
rect 16930 480 16940 500
rect 16960 480 16970 500
rect 16930 465 16970 480
rect 18630 750 18670 765
rect 18630 730 18640 750
rect 18660 730 18670 750
rect 18630 700 18670 730
rect 18630 680 18640 700
rect 18660 680 18670 700
rect 18630 650 18670 680
rect 18630 630 18640 650
rect 18660 630 18670 650
rect 18630 600 18670 630
rect 18630 580 18640 600
rect 18660 580 18670 600
rect 18630 550 18670 580
rect 18865 750 18905 765
rect 18865 730 18875 750
rect 18895 730 18905 750
rect 18865 700 18905 730
rect 18865 680 18875 700
rect 18895 680 18905 700
rect 18865 650 18905 680
rect 18865 630 18875 650
rect 18895 630 18905 650
rect 18865 600 18905 630
rect 18865 580 18875 600
rect 18895 580 18905 600
rect 18865 565 18905 580
rect 19110 750 19150 765
rect 19110 730 19120 750
rect 19140 730 19150 750
rect 19110 700 19150 730
rect 19110 680 19120 700
rect 19140 680 19150 700
rect 19110 650 19150 680
rect 19110 630 19120 650
rect 19140 630 19150 650
rect 19110 600 19150 630
rect 19110 580 19120 600
rect 19140 580 19150 600
rect 19110 565 19150 580
rect 18630 530 18640 550
rect 18660 530 18670 550
rect 18630 500 18670 530
rect 18630 480 18640 500
rect 18660 480 18670 500
rect 18630 465 18670 480
rect 16380 -90 16420 -75
rect 16380 -110 16390 -90
rect 16410 -110 16420 -90
rect 16380 -140 16420 -110
rect 16380 -160 16390 -140
rect 16410 -160 16420 -140
rect 16380 -175 16420 -160
rect 17660 -90 17700 -75
rect 17660 -110 17670 -90
rect 17690 -110 17700 -90
rect 17660 -140 17700 -110
rect 17660 -160 17670 -140
rect 17690 -160 17700 -140
rect 17660 -175 17700 -160
rect 17900 -90 17940 -75
rect 17900 -110 17910 -90
rect 17930 -110 17940 -90
rect 17900 -140 17940 -110
rect 17900 -160 17910 -140
rect 17930 -160 17940 -140
rect 17900 -175 17940 -160
rect 19180 -90 19220 -75
rect 19180 -110 19190 -90
rect 19210 -110 19220 -90
rect 19180 -140 19220 -110
rect 19180 -160 19190 -140
rect 19210 -160 19220 -140
rect 19180 -175 19220 -160
<< psubdiffcont >>
rect 17570 -395 17590 -375
rect 18010 -395 18030 -375
rect 17120 -845 17140 -825
rect 17120 -895 17140 -875
rect 17120 -945 17140 -925
rect 17120 -995 17140 -975
rect 17120 -1045 17140 -1025
rect 18460 -845 18480 -825
rect 18460 -895 18480 -875
rect 18460 -945 18480 -925
rect 18460 -995 18480 -975
rect 18460 -1045 18480 -1025
rect 18870 -1225 18890 -1205
rect 18870 -1275 18890 -1255
rect 16510 -1575 16530 -1555
rect 16510 -1625 16530 -1605
rect 16865 -1575 16885 -1555
rect 16865 -1625 16885 -1605
rect 16995 -1575 17015 -1555
rect 16995 -1625 17015 -1605
rect 17515 -1575 17535 -1555
rect 17515 -1625 17535 -1605
rect 17585 -1575 17605 -1555
rect 17585 -1625 17605 -1605
rect 17995 -1575 18015 -1555
rect 17995 -1625 18015 -1605
rect 18065 -1575 18085 -1555
rect 18065 -1625 18085 -1605
rect 18585 -1575 18605 -1555
rect 18585 -1625 18605 -1605
rect 17790 -4190 17810 -4170
rect 17790 -4240 17810 -4220
rect 17790 -4290 17810 -4270
<< nsubdiffcont >>
rect 16345 1195 16365 1217
rect 16345 1145 16365 1165
rect 16645 1195 16665 1217
rect 16645 1145 16665 1165
rect 16855 1145 16875 1217
rect 17265 1145 17285 1217
rect 17475 1195 17495 1217
rect 17475 1145 17495 1165
rect 18105 1195 18125 1217
rect 18105 1145 18125 1165
rect 18315 1145 18335 1217
rect 18725 1145 18745 1217
rect 16940 730 16960 750
rect 16940 680 16960 700
rect 16405 630 16425 650
rect 16405 580 16425 600
rect 16710 630 16730 650
rect 16710 580 16730 600
rect 16940 630 16960 650
rect 16940 580 16960 600
rect 16940 530 16960 550
rect 16940 480 16960 500
rect 18640 730 18660 750
rect 18640 680 18660 700
rect 18640 630 18660 650
rect 18640 580 18660 600
rect 18875 730 18895 750
rect 18875 680 18895 700
rect 18875 630 18895 650
rect 18875 580 18895 600
rect 19120 730 19140 750
rect 19120 680 19140 700
rect 19120 630 19140 650
rect 19120 580 19140 600
rect 18640 530 18660 550
rect 18640 480 18660 500
rect 16390 -110 16410 -90
rect 16390 -160 16410 -140
rect 17670 -110 17690 -90
rect 17670 -160 17690 -140
rect 17910 -110 17930 -90
rect 17910 -160 17930 -140
rect 19190 -110 19210 -90
rect 19190 -160 19210 -140
<< poly >>
rect 16485 1455 16525 1465
rect 16485 1435 16495 1455
rect 16515 1435 16525 1455
rect 16485 1425 16525 1435
rect 17780 1455 17820 1465
rect 17780 1435 17790 1455
rect 17810 1435 17820 1455
rect 17780 1425 17820 1435
rect 16365 1275 16405 1285
rect 16365 1255 16375 1275
rect 16395 1260 16405 1275
rect 16395 1255 16430 1260
rect 16495 1255 16515 1425
rect 16605 1275 16645 1285
rect 16605 1260 16615 1275
rect 16580 1255 16615 1260
rect 16635 1255 16645 1275
rect 16365 1245 16430 1255
rect 16415 1230 16430 1245
rect 16470 1240 16540 1255
rect 16470 1230 16485 1240
rect 16525 1230 16540 1240
rect 16580 1245 16645 1255
rect 16885 1275 16925 1285
rect 16885 1255 16895 1275
rect 16915 1255 16925 1275
rect 17055 1275 17085 1285
rect 17055 1255 17060 1275
rect 17080 1255 17085 1275
rect 17215 1275 17255 1285
rect 17215 1255 17225 1275
rect 17245 1255 17255 1275
rect 16580 1230 16595 1245
rect 16885 1240 16940 1255
rect 16925 1230 16940 1240
rect 16980 1240 17160 1255
rect 16980 1230 16995 1240
rect 17035 1230 17050 1240
rect 17090 1230 17105 1240
rect 17145 1230 17160 1240
rect 17200 1240 17255 1255
rect 17495 1275 17535 1285
rect 17495 1255 17505 1275
rect 17525 1260 17535 1275
rect 17525 1255 17560 1260
rect 17790 1255 17810 1425
rect 18065 1275 18105 1285
rect 18065 1260 18075 1275
rect 18040 1255 18075 1260
rect 18095 1255 18105 1275
rect 17495 1245 17560 1255
rect 17200 1230 17215 1240
rect 17545 1230 17560 1245
rect 17600 1240 18000 1255
rect 17600 1230 17615 1240
rect 17655 1230 17670 1240
rect 17710 1230 17725 1240
rect 17765 1230 17780 1240
rect 17820 1230 17835 1240
rect 17875 1230 17890 1240
rect 17930 1230 17945 1240
rect 17985 1230 18000 1240
rect 18040 1245 18105 1255
rect 18345 1275 18385 1285
rect 18345 1255 18355 1275
rect 18375 1260 18385 1275
rect 18515 1275 18545 1285
rect 18375 1255 18400 1260
rect 18515 1255 18520 1275
rect 18540 1255 18545 1275
rect 18675 1275 18715 1285
rect 18675 1260 18685 1275
rect 18660 1255 18685 1260
rect 18705 1255 18715 1275
rect 18345 1245 18400 1255
rect 18040 1230 18055 1245
rect 18385 1230 18400 1245
rect 18440 1240 18620 1255
rect 18440 1230 18455 1240
rect 18495 1230 18510 1240
rect 18550 1230 18565 1240
rect 18605 1230 18620 1240
rect 18660 1245 18715 1255
rect 18660 1230 18675 1245
rect 16415 1115 16430 1130
rect 16470 1115 16485 1130
rect 16525 1115 16540 1130
rect 16580 1115 16595 1130
rect 16925 1115 16940 1130
rect 16980 1115 16995 1130
rect 17035 1115 17050 1130
rect 17090 1115 17105 1130
rect 17145 1115 17160 1130
rect 17200 1115 17215 1130
rect 17545 1115 17560 1130
rect 17600 1115 17615 1130
rect 17655 1115 17670 1130
rect 17710 1115 17725 1130
rect 17765 1115 17780 1130
rect 17820 1115 17835 1130
rect 17875 1115 17890 1130
rect 17930 1115 17945 1130
rect 17985 1115 18000 1130
rect 18040 1115 18055 1130
rect 18385 1115 18400 1130
rect 18440 1115 18455 1130
rect 18495 1115 18510 1130
rect 18550 1115 18565 1130
rect 18605 1115 18620 1130
rect 18660 1115 18675 1130
rect 16970 810 17010 820
rect 16970 790 16980 810
rect 17000 795 17010 810
rect 18590 810 18630 820
rect 18590 795 18600 810
rect 17000 790 17060 795
rect 16970 780 17060 790
rect 18540 790 18600 795
rect 18620 790 18630 810
rect 18540 780 18630 790
rect 18910 810 18940 820
rect 18910 790 18915 810
rect 18935 795 18940 810
rect 19080 810 19110 820
rect 19080 795 19085 810
rect 18935 790 18960 795
rect 18910 780 18960 790
rect 19055 790 19085 795
rect 19105 790 19110 810
rect 19055 780 19110 790
rect 17010 765 17060 780
rect 17100 765 17150 780
rect 17190 765 17240 780
rect 17280 765 17330 780
rect 17370 765 17420 780
rect 17460 765 17510 780
rect 17550 765 17600 780
rect 17640 765 17690 780
rect 17730 765 17780 780
rect 17820 765 17870 780
rect 17910 765 17960 780
rect 18000 765 18050 780
rect 18090 765 18140 780
rect 18180 765 18230 780
rect 18270 765 18320 780
rect 18360 765 18410 780
rect 18450 765 18500 780
rect 18540 765 18590 780
rect 18945 765 18960 780
rect 19000 765 19015 780
rect 19055 765 19070 780
rect 16440 710 16470 720
rect 16440 690 16445 710
rect 16465 690 16470 710
rect 16660 710 16690 720
rect 16660 690 16665 710
rect 16685 690 16690 710
rect 16440 675 16490 690
rect 16475 665 16490 675
rect 16530 665 16545 680
rect 16585 665 16600 680
rect 16640 675 16690 690
rect 16640 665 16655 675
rect 16475 550 16490 565
rect 16530 555 16545 565
rect 16585 555 16600 565
rect 16530 540 16600 555
rect 16640 550 16655 565
rect 16545 520 16555 540
rect 16575 520 16585 540
rect 16545 510 16585 520
rect 18945 550 18960 565
rect 19000 495 19015 565
rect 19055 550 19070 565
rect 19000 490 19040 495
rect 19000 470 19010 490
rect 19030 470 19040 490
rect 19000 465 19040 470
rect 17010 450 17060 465
rect 17100 455 17150 465
rect 17190 455 17240 465
rect 17280 455 17330 465
rect 17370 455 17420 465
rect 17460 455 17510 465
rect 17550 455 17600 465
rect 17640 455 17690 465
rect 17730 455 17780 465
rect 17820 455 17870 465
rect 17910 455 17960 465
rect 18000 455 18050 465
rect 18090 455 18140 465
rect 18180 455 18230 465
rect 18270 455 18320 465
rect 18360 455 18410 465
rect 18450 455 18500 465
rect 17100 440 18500 455
rect 18540 450 18590 465
rect 17690 420 17700 440
rect 17720 420 17730 440
rect 17690 410 17730 420
rect 18410 420 18420 440
rect 18440 420 18450 440
rect 18410 410 18450 420
rect 16425 -30 16455 -20
rect 16425 -50 16430 -30
rect 16450 -50 16455 -30
rect 17625 -30 17655 -20
rect 17625 -50 17630 -30
rect 17650 -50 17655 -30
rect 16425 -65 16480 -50
rect 16460 -75 16480 -65
rect 16520 -75 16540 -60
rect 16580 -75 16600 -60
rect 16640 -75 16660 -60
rect 16700 -75 16720 -60
rect 16760 -75 16780 -60
rect 16820 -75 16840 -60
rect 16880 -75 16900 -60
rect 16940 -75 16960 -60
rect 17000 -75 17020 -60
rect 17060 -75 17080 -60
rect 17120 -75 17140 -60
rect 17180 -75 17200 -60
rect 17240 -75 17260 -60
rect 17300 -75 17320 -60
rect 17360 -75 17380 -60
rect 17420 -75 17440 -60
rect 17480 -75 17500 -60
rect 17540 -75 17560 -60
rect 17600 -65 17655 -50
rect 17945 -30 17975 -20
rect 17945 -50 17950 -30
rect 17970 -50 17975 -30
rect 19145 -30 19175 -20
rect 19145 -50 19150 -30
rect 19170 -50 19175 -30
rect 17945 -65 18000 -50
rect 17600 -75 17620 -65
rect 17980 -75 18000 -65
rect 18040 -75 18060 -60
rect 18100 -75 18120 -60
rect 18160 -75 18180 -60
rect 18220 -75 18240 -60
rect 18280 -75 18300 -60
rect 18340 -75 18360 -60
rect 18400 -75 18420 -60
rect 18460 -75 18480 -60
rect 18520 -75 18540 -60
rect 18580 -75 18600 -60
rect 18640 -75 18660 -60
rect 18700 -75 18720 -60
rect 18760 -75 18780 -60
rect 18820 -75 18840 -60
rect 18880 -75 18900 -60
rect 18940 -75 18960 -60
rect 19000 -75 19020 -60
rect 19060 -75 19080 -60
rect 19120 -65 19175 -50
rect 19120 -75 19140 -65
rect 16460 -185 16480 -175
rect 16425 -200 16480 -185
rect 16520 -190 16540 -175
rect 16580 -185 16600 -175
rect 16640 -185 16660 -175
rect 16700 -185 16720 -175
rect 16760 -185 16780 -175
rect 16510 -200 16550 -190
rect 16580 -200 16780 -185
rect 16820 -185 16840 -175
rect 16880 -185 16900 -175
rect 16820 -200 16900 -185
rect 16940 -185 16960 -175
rect 17000 -185 17020 -175
rect 17060 -185 17080 -175
rect 17120 -185 17140 -175
rect 16940 -200 17140 -185
rect 17180 -185 17200 -175
rect 17240 -185 17260 -175
rect 17180 -200 17260 -185
rect 17300 -185 17320 -175
rect 17360 -185 17380 -175
rect 17420 -185 17440 -175
rect 17480 -185 17500 -175
rect 17300 -200 17500 -185
rect 17540 -190 17560 -175
rect 17600 -190 17620 -175
rect 17980 -185 18000 -175
rect 17535 -200 17565 -190
rect 16425 -220 16430 -200
rect 16450 -220 16455 -200
rect 16425 -230 16455 -220
rect 16510 -220 16520 -200
rect 16540 -220 16550 -200
rect 16510 -230 16550 -220
rect 16600 -220 16610 -200
rect 16630 -220 16640 -200
rect 16600 -230 16640 -220
rect 16840 -220 16850 -200
rect 16870 -220 16880 -200
rect 16840 -230 16880 -220
rect 16960 -220 16970 -200
rect 16990 -220 17000 -200
rect 16960 -230 17000 -220
rect 17200 -220 17210 -200
rect 17230 -220 17240 -200
rect 17200 -230 17240 -220
rect 17320 -220 17330 -200
rect 17350 -220 17360 -200
rect 17320 -230 17360 -220
rect 17535 -220 17540 -200
rect 17560 -220 17565 -200
rect 17535 -230 17565 -220
rect 17945 -200 18000 -185
rect 18040 -190 18060 -175
rect 18100 -185 18120 -175
rect 18160 -185 18180 -175
rect 18220 -185 18240 -175
rect 18280 -185 18300 -175
rect 18035 -200 18065 -190
rect 18100 -200 18300 -185
rect 18340 -185 18360 -175
rect 18400 -185 18420 -175
rect 18340 -200 18420 -185
rect 18460 -185 18480 -175
rect 18520 -185 18540 -175
rect 18580 -185 18600 -175
rect 18640 -185 18660 -175
rect 18460 -200 18660 -185
rect 18700 -185 18720 -175
rect 18760 -185 18780 -175
rect 18700 -200 18780 -185
rect 18820 -185 18840 -175
rect 18880 -185 18900 -175
rect 18940 -185 18960 -175
rect 19000 -185 19020 -175
rect 18820 -200 19020 -185
rect 19060 -190 19080 -175
rect 19120 -185 19140 -175
rect 19050 -200 19090 -190
rect 19120 -200 19175 -185
rect 17945 -220 17950 -200
rect 17970 -220 17975 -200
rect 17945 -230 17975 -220
rect 18035 -220 18040 -200
rect 18060 -220 18065 -200
rect 18035 -230 18065 -220
rect 18240 -220 18250 -200
rect 18270 -220 18280 -200
rect 18240 -230 18280 -220
rect 18360 -220 18370 -200
rect 18390 -220 18400 -200
rect 18360 -230 18400 -220
rect 18600 -220 18610 -200
rect 18630 -220 18640 -200
rect 18600 -230 18640 -220
rect 18720 -220 18730 -200
rect 18750 -220 18760 -200
rect 18720 -230 18760 -220
rect 18960 -220 18970 -200
rect 18990 -220 19000 -200
rect 18960 -230 19000 -220
rect 19050 -220 19060 -200
rect 19080 -220 19090 -200
rect 19050 -230 19090 -220
rect 19145 -220 19150 -200
rect 19170 -220 19175 -200
rect 19145 -230 19175 -220
rect 17007 -315 17037 -305
rect 17007 -330 17012 -315
rect 17000 -335 17012 -330
rect 17032 -335 17037 -315
rect 17000 -345 17037 -335
rect 18563 -315 18593 -305
rect 18563 -335 18568 -315
rect 18588 -330 18593 -315
rect 18588 -335 18600 -330
rect 18563 -345 18600 -335
rect 17000 -360 17020 -345
rect 17060 -360 17080 -345
rect 18520 -360 18540 -345
rect 18580 -360 18600 -345
rect 17000 -625 17020 -610
rect 17060 -625 17080 -610
rect 18520 -625 18540 -610
rect 18580 -625 18600 -610
rect 17060 -635 17105 -625
rect 17060 -655 17080 -635
rect 17100 -655 17105 -635
rect 17060 -665 17105 -655
rect 18495 -635 18540 -625
rect 18495 -655 18500 -635
rect 18520 -655 18540 -635
rect 18495 -665 18540 -655
rect 16620 -770 16660 -760
rect 16620 -790 16630 -770
rect 16650 -790 16660 -770
rect 16620 -795 16660 -790
rect 16740 -770 16780 -760
rect 16740 -790 16750 -770
rect 16770 -790 16780 -770
rect 16740 -795 16780 -790
rect 16860 -770 16900 -760
rect 16860 -790 16870 -770
rect 16890 -790 16900 -770
rect 16860 -795 16900 -790
rect 16980 -770 17020 -760
rect 16980 -790 16990 -770
rect 17010 -790 17020 -770
rect 16980 -795 17020 -790
rect 17300 -770 17340 -760
rect 17300 -790 17310 -770
rect 17330 -790 17340 -770
rect 17300 -795 17340 -790
rect 17420 -770 17460 -760
rect 17420 -790 17430 -770
rect 17450 -790 17460 -770
rect 17420 -795 17460 -790
rect 17540 -770 17580 -760
rect 17540 -790 17550 -770
rect 17570 -790 17580 -770
rect 17540 -795 17580 -790
rect 18020 -770 18060 -760
rect 18020 -790 18030 -770
rect 18050 -790 18060 -770
rect 18020 -795 18060 -790
rect 18140 -770 18180 -760
rect 18140 -790 18150 -770
rect 18170 -790 18180 -770
rect 18140 -795 18180 -790
rect 18260 -770 18300 -760
rect 18260 -790 18270 -770
rect 18290 -790 18300 -770
rect 18260 -795 18300 -790
rect 18580 -770 18620 -760
rect 18580 -790 18590 -770
rect 18610 -790 18620 -770
rect 18580 -795 18620 -790
rect 18700 -770 18740 -760
rect 18700 -790 18710 -770
rect 18730 -790 18740 -770
rect 18700 -795 18740 -790
rect 18820 -770 18860 -760
rect 18820 -790 18830 -770
rect 18850 -790 18860 -770
rect 18820 -795 18860 -790
rect 18940 -770 18980 -760
rect 18940 -790 18950 -770
rect 18970 -790 18980 -770
rect 18940 -795 18980 -790
rect 16570 -810 17070 -795
rect 17190 -810 17690 -795
rect 17910 -810 18410 -795
rect 18530 -810 19030 -795
rect 16570 -1075 17070 -1060
rect 17190 -1075 17690 -1060
rect 17910 -1075 18410 -1060
rect 18530 -1075 19030 -1060
rect 16820 -1145 16860 -1135
rect 16820 -1165 16830 -1145
rect 16850 -1165 16860 -1145
rect 16820 -1175 16860 -1165
rect 16900 -1145 16940 -1135
rect 16900 -1165 16910 -1145
rect 16930 -1165 16940 -1145
rect 16900 -1175 16940 -1165
rect 16980 -1145 17020 -1135
rect 16980 -1165 16990 -1145
rect 17010 -1165 17020 -1145
rect 16980 -1175 17020 -1165
rect 17060 -1145 17100 -1135
rect 17060 -1165 17070 -1145
rect 17090 -1165 17100 -1145
rect 17060 -1175 17100 -1165
rect 17140 -1145 17180 -1135
rect 17140 -1165 17150 -1145
rect 17170 -1165 17180 -1145
rect 17140 -1175 17180 -1165
rect 17220 -1145 17260 -1135
rect 17220 -1165 17230 -1145
rect 17250 -1165 17260 -1145
rect 17220 -1175 17260 -1165
rect 17300 -1145 17340 -1135
rect 17300 -1165 17310 -1145
rect 17330 -1165 17340 -1145
rect 17300 -1175 17340 -1165
rect 17380 -1145 17420 -1135
rect 17380 -1165 17390 -1145
rect 17410 -1165 17420 -1145
rect 17380 -1175 17420 -1165
rect 17460 -1145 17500 -1135
rect 17460 -1165 17470 -1145
rect 17490 -1165 17500 -1145
rect 17460 -1175 17500 -1165
rect 17540 -1145 17580 -1135
rect 17540 -1165 17550 -1145
rect 17570 -1165 17580 -1145
rect 17540 -1175 17580 -1165
rect 17620 -1145 17660 -1135
rect 17620 -1165 17630 -1145
rect 17650 -1165 17660 -1145
rect 17620 -1175 17660 -1165
rect 17700 -1145 17740 -1135
rect 17700 -1165 17710 -1145
rect 17730 -1165 17740 -1145
rect 17700 -1175 17740 -1165
rect 17860 -1145 17900 -1135
rect 17860 -1165 17870 -1145
rect 17890 -1165 17900 -1145
rect 17860 -1175 17900 -1165
rect 17940 -1145 17980 -1135
rect 17940 -1165 17950 -1145
rect 17970 -1165 17980 -1145
rect 17940 -1175 17980 -1165
rect 18020 -1145 18060 -1135
rect 18020 -1165 18030 -1145
rect 18050 -1165 18060 -1145
rect 18020 -1175 18060 -1165
rect 18100 -1145 18140 -1135
rect 18100 -1165 18110 -1145
rect 18130 -1165 18140 -1145
rect 18100 -1175 18140 -1165
rect 18180 -1145 18220 -1135
rect 18180 -1165 18190 -1145
rect 18210 -1165 18220 -1145
rect 18180 -1175 18220 -1165
rect 18260 -1145 18300 -1135
rect 18260 -1165 18270 -1145
rect 18290 -1165 18300 -1145
rect 18260 -1175 18300 -1165
rect 18340 -1145 18380 -1135
rect 18340 -1165 18350 -1145
rect 18370 -1165 18380 -1145
rect 18340 -1175 18380 -1165
rect 18420 -1145 18460 -1135
rect 18420 -1165 18430 -1145
rect 18450 -1165 18460 -1145
rect 18420 -1175 18460 -1165
rect 18500 -1145 18540 -1135
rect 18500 -1165 18510 -1145
rect 18530 -1165 18540 -1145
rect 18500 -1175 18540 -1165
rect 18580 -1145 18620 -1135
rect 18580 -1165 18590 -1145
rect 18610 -1165 18620 -1145
rect 18580 -1175 18620 -1165
rect 18660 -1145 18700 -1135
rect 18660 -1165 18670 -1145
rect 18690 -1165 18700 -1145
rect 18660 -1175 18700 -1165
rect 18740 -1145 18780 -1135
rect 18740 -1165 18750 -1145
rect 18770 -1165 18780 -1145
rect 18740 -1175 18780 -1165
rect 16780 -1190 17780 -1175
rect 17820 -1190 18820 -1175
rect 16780 -1305 17780 -1290
rect 17820 -1305 18820 -1290
rect 16540 -1495 16580 -1485
rect 16540 -1515 16550 -1495
rect 16570 -1510 16580 -1495
rect 16710 -1495 16740 -1485
rect 16570 -1515 16595 -1510
rect 16710 -1515 16715 -1495
rect 16735 -1515 16740 -1495
rect 16820 -1495 16860 -1485
rect 16820 -1510 16830 -1495
rect 16800 -1515 16830 -1510
rect 16850 -1515 16860 -1495
rect 16540 -1525 16595 -1515
rect 16580 -1540 16595 -1525
rect 16635 -1530 16760 -1515
rect 16635 -1540 16650 -1530
rect 16690 -1540 16705 -1530
rect 16745 -1540 16760 -1530
rect 16800 -1525 16860 -1515
rect 17025 -1495 17065 -1485
rect 17025 -1515 17035 -1495
rect 17055 -1510 17065 -1495
rect 17305 -1495 17335 -1485
rect 17055 -1515 17080 -1510
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17465 -1495 17505 -1485
rect 17465 -1510 17475 -1495
rect 17450 -1515 17475 -1510
rect 17495 -1515 17505 -1495
rect 17025 -1525 17080 -1515
rect 16800 -1540 16815 -1525
rect 17065 -1540 17080 -1525
rect 17120 -1530 17410 -1515
rect 17120 -1540 17135 -1530
rect 17175 -1540 17190 -1530
rect 17230 -1540 17245 -1530
rect 17285 -1540 17300 -1530
rect 17340 -1540 17355 -1530
rect 17395 -1540 17410 -1530
rect 17450 -1525 17505 -1515
rect 17615 -1495 17655 -1485
rect 17615 -1515 17625 -1495
rect 17645 -1510 17655 -1495
rect 17785 -1495 17815 -1485
rect 17645 -1515 17670 -1510
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17945 -1495 17985 -1485
rect 17945 -1510 17955 -1495
rect 17930 -1515 17955 -1510
rect 17975 -1515 17985 -1495
rect 17615 -1525 17670 -1515
rect 17450 -1540 17465 -1525
rect 17655 -1540 17670 -1525
rect 17710 -1530 17890 -1515
rect 17710 -1540 17725 -1530
rect 17765 -1540 17780 -1530
rect 17820 -1540 17835 -1530
rect 17875 -1540 17890 -1530
rect 17930 -1525 17985 -1515
rect 18095 -1495 18135 -1485
rect 18095 -1515 18105 -1495
rect 18125 -1510 18135 -1495
rect 18265 -1495 18295 -1485
rect 18125 -1515 18150 -1510
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18535 -1495 18575 -1485
rect 18535 -1510 18545 -1495
rect 18520 -1515 18545 -1510
rect 18565 -1515 18575 -1495
rect 18095 -1525 18150 -1515
rect 17930 -1540 17945 -1525
rect 18135 -1540 18150 -1525
rect 18190 -1530 18480 -1515
rect 18190 -1540 18205 -1530
rect 18245 -1540 18260 -1530
rect 18300 -1540 18315 -1530
rect 18355 -1540 18370 -1530
rect 18410 -1540 18425 -1530
rect 18465 -1540 18480 -1530
rect 18520 -1525 18575 -1515
rect 18520 -1540 18535 -1525
rect 16580 -1655 16595 -1640
rect 16635 -1655 16650 -1640
rect 16690 -1655 16705 -1640
rect 16745 -1655 16760 -1640
rect 16800 -1655 16815 -1640
rect 17065 -1655 17080 -1640
rect 17120 -1655 17135 -1640
rect 17175 -1655 17190 -1640
rect 17230 -1655 17245 -1640
rect 17285 -1655 17300 -1640
rect 17340 -1655 17355 -1640
rect 17395 -1655 17410 -1640
rect 17450 -1655 17465 -1640
rect 17655 -1655 17670 -1640
rect 17710 -1655 17725 -1640
rect 17765 -1655 17780 -1640
rect 17820 -1655 17835 -1640
rect 17875 -1655 17890 -1640
rect 17930 -1655 17945 -1640
rect 18135 -1655 18150 -1640
rect 18190 -1655 18205 -1640
rect 18245 -1655 18260 -1640
rect 18300 -1655 18315 -1640
rect 18355 -1655 18370 -1640
rect 18410 -1655 18425 -1640
rect 18465 -1655 18480 -1640
rect 18520 -1655 18535 -1640
<< polycont >>
rect 16495 1435 16515 1455
rect 17790 1435 17810 1455
rect 16375 1255 16395 1275
rect 16615 1255 16635 1275
rect 16895 1255 16915 1275
rect 17060 1255 17080 1275
rect 17225 1255 17245 1275
rect 17505 1255 17525 1275
rect 18075 1255 18095 1275
rect 18355 1255 18375 1275
rect 18520 1255 18540 1275
rect 18685 1255 18705 1275
rect 16980 790 17000 810
rect 18600 790 18620 810
rect 18915 790 18935 810
rect 19085 790 19105 810
rect 16445 690 16465 710
rect 16665 690 16685 710
rect 16555 520 16575 540
rect 19010 470 19030 490
rect 17700 420 17720 440
rect 18420 420 18440 440
rect 16430 -50 16450 -30
rect 17630 -50 17650 -30
rect 17950 -50 17970 -30
rect 19150 -50 19170 -30
rect 16430 -220 16450 -200
rect 16520 -220 16540 -200
rect 16610 -220 16630 -200
rect 16850 -220 16870 -200
rect 16970 -220 16990 -200
rect 17210 -220 17230 -200
rect 17330 -220 17350 -200
rect 17540 -220 17560 -200
rect 17950 -220 17970 -200
rect 18040 -220 18060 -200
rect 18250 -220 18270 -200
rect 18370 -220 18390 -200
rect 18610 -220 18630 -200
rect 18730 -220 18750 -200
rect 18970 -220 18990 -200
rect 19060 -220 19080 -200
rect 19150 -220 19170 -200
rect 17012 -335 17032 -315
rect 18568 -335 18588 -315
rect 17080 -655 17100 -635
rect 18500 -655 18520 -635
rect 16630 -790 16650 -770
rect 16750 -790 16770 -770
rect 16870 -790 16890 -770
rect 16990 -790 17010 -770
rect 17310 -790 17330 -770
rect 17430 -790 17450 -770
rect 17550 -790 17570 -770
rect 18030 -790 18050 -770
rect 18150 -790 18170 -770
rect 18270 -790 18290 -770
rect 18590 -790 18610 -770
rect 18710 -790 18730 -770
rect 18830 -790 18850 -770
rect 18950 -790 18970 -770
rect 16830 -1165 16850 -1145
rect 16910 -1165 16930 -1145
rect 16990 -1165 17010 -1145
rect 17070 -1165 17090 -1145
rect 17150 -1165 17170 -1145
rect 17230 -1165 17250 -1145
rect 17310 -1165 17330 -1145
rect 17390 -1165 17410 -1145
rect 17470 -1165 17490 -1145
rect 17550 -1165 17570 -1145
rect 17630 -1165 17650 -1145
rect 17710 -1165 17730 -1145
rect 17870 -1165 17890 -1145
rect 17950 -1165 17970 -1145
rect 18030 -1165 18050 -1145
rect 18110 -1165 18130 -1145
rect 18190 -1165 18210 -1145
rect 18270 -1165 18290 -1145
rect 18350 -1165 18370 -1145
rect 18430 -1165 18450 -1145
rect 18510 -1165 18530 -1145
rect 18590 -1165 18610 -1145
rect 18670 -1165 18690 -1145
rect 18750 -1165 18770 -1145
rect 16550 -1515 16570 -1495
rect 16715 -1515 16735 -1495
rect 16830 -1515 16850 -1495
rect 17035 -1515 17055 -1495
rect 17310 -1515 17330 -1495
rect 17475 -1515 17495 -1495
rect 17625 -1515 17645 -1495
rect 17790 -1515 17810 -1495
rect 17955 -1515 17975 -1495
rect 18105 -1515 18125 -1495
rect 18270 -1515 18290 -1495
rect 18545 -1515 18565 -1495
<< xpolycontact >>
rect 17470 -2035 17690 -2000
rect 17904 -2035 18124 -2000
rect 15950 -3376 15985 -3156
rect 15950 -3784 15985 -3565
rect 16160 -3285 16195 -3065
rect 16160 -3889 16195 -3669
rect 16220 -3285 16255 -3065
rect 16220 -3889 16255 -3669
rect 16280 -3285 16315 -3065
rect 16280 -3889 16315 -3669
rect 16485 -3160 16520 -2940
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19285 -3257 19320 -3037
rect 19285 -3889 19320 -3669
rect 19345 -3257 19380 -3037
rect 19345 -3889 19380 -3669
rect 19405 -3257 19440 -3037
rect 19405 -3889 19440 -3669
rect 19610 -3376 19645 -3156
rect 19610 -3784 19645 -3565
<< ppolyres >>
rect 15950 -3565 15985 -3376
rect 19610 -3565 19645 -3376
<< xpolyres >>
rect 17690 -2035 17904 -2000
rect 16160 -3669 16195 -3285
rect 16220 -3669 16255 -3285
rect 16280 -3669 16315 -3285
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19285 -3669 19320 -3257
rect 19345 -3669 19380 -3257
rect 19405 -3669 19440 -3257
<< locali >>
rect 16485 1455 16525 1465
rect 16485 1435 16495 1455
rect 16515 1435 16525 1455
rect 16485 1425 16525 1435
rect 17780 1455 17820 1465
rect 17780 1435 17790 1455
rect 17810 1435 17820 1455
rect 17780 1425 17820 1435
rect 16365 1275 16405 1285
rect 16365 1255 16375 1275
rect 16395 1255 16405 1275
rect 16365 1245 16405 1255
rect 16485 1275 16525 1285
rect 16485 1255 16495 1275
rect 16515 1255 16525 1275
rect 16485 1245 16525 1255
rect 16605 1275 16645 1285
rect 16605 1255 16615 1275
rect 16635 1255 16645 1275
rect 16605 1245 16645 1255
rect 16885 1275 16925 1285
rect 16885 1255 16895 1275
rect 16915 1255 16925 1275
rect 16885 1245 16925 1255
rect 16945 1275 16975 1285
rect 16945 1255 16950 1275
rect 16970 1255 16975 1275
rect 16945 1245 16975 1255
rect 16995 1275 17035 1285
rect 16995 1255 17005 1275
rect 17025 1255 17035 1275
rect 16995 1245 17035 1255
rect 17055 1275 17085 1285
rect 17055 1255 17060 1275
rect 17080 1255 17085 1275
rect 17055 1245 17085 1255
rect 17105 1275 17145 1285
rect 17105 1255 17115 1275
rect 17135 1255 17145 1275
rect 17105 1245 17145 1255
rect 17215 1275 17255 1285
rect 17215 1255 17225 1275
rect 17245 1255 17255 1275
rect 17215 1245 17255 1255
rect 17495 1275 17535 1285
rect 17495 1255 17505 1275
rect 17525 1255 17535 1275
rect 17495 1245 17535 1255
rect 17560 1275 17600 1285
rect 17560 1255 17570 1275
rect 17590 1255 17600 1275
rect 17560 1245 17600 1255
rect 17620 1275 17650 1285
rect 17620 1255 17625 1275
rect 17645 1255 17650 1275
rect 16385 1225 16405 1245
rect 16495 1225 16515 1245
rect 16605 1225 16625 1245
rect 16895 1225 16915 1245
rect 16950 1225 16970 1245
rect 17005 1225 17025 1245
rect 17115 1225 17135 1245
rect 17225 1225 17245 1245
rect 17515 1225 17535 1245
rect 17570 1225 17590 1245
rect 16340 1217 16410 1225
rect 16340 1195 16345 1217
rect 16365 1215 16410 1217
rect 16365 1195 16385 1215
rect 16405 1195 16410 1215
rect 16340 1165 16410 1195
rect 16340 1145 16345 1165
rect 16365 1145 16385 1165
rect 16405 1145 16410 1165
rect 16340 1135 16410 1145
rect 16435 1215 16465 1225
rect 16435 1195 16440 1215
rect 16460 1195 16465 1215
rect 16435 1165 16465 1195
rect 16435 1145 16440 1165
rect 16460 1145 16465 1165
rect 16435 1135 16465 1145
rect 16490 1215 16520 1225
rect 16490 1195 16495 1215
rect 16515 1195 16520 1215
rect 16490 1165 16520 1195
rect 16490 1145 16495 1165
rect 16515 1145 16520 1165
rect 16490 1135 16520 1145
rect 16545 1215 16575 1225
rect 16545 1195 16550 1215
rect 16570 1195 16575 1215
rect 16545 1165 16575 1195
rect 16545 1145 16550 1165
rect 16570 1145 16575 1165
rect 16545 1135 16575 1145
rect 16600 1217 16670 1225
rect 16600 1215 16645 1217
rect 16600 1195 16605 1215
rect 16625 1195 16645 1215
rect 16665 1195 16670 1217
rect 16600 1165 16670 1195
rect 16600 1145 16605 1165
rect 16625 1145 16645 1165
rect 16665 1145 16670 1165
rect 16600 1135 16670 1145
rect 16850 1217 16920 1225
rect 16850 1145 16855 1217
rect 16875 1215 16920 1217
rect 16875 1145 16895 1215
rect 16850 1143 16895 1145
rect 16915 1143 16920 1215
rect 16850 1135 16920 1143
rect 16945 1215 16975 1225
rect 16945 1143 16950 1215
rect 16970 1143 16975 1215
rect 16945 1135 16975 1143
rect 17000 1215 17030 1225
rect 17000 1143 17005 1215
rect 17025 1143 17030 1215
rect 17000 1135 17030 1143
rect 17055 1215 17085 1225
rect 17055 1143 17060 1215
rect 17080 1143 17085 1215
rect 17055 1135 17085 1143
rect 17110 1215 17140 1225
rect 17110 1143 17115 1215
rect 17135 1143 17140 1215
rect 17110 1135 17140 1143
rect 17165 1215 17195 1225
rect 17165 1143 17170 1215
rect 17190 1143 17195 1215
rect 17165 1135 17195 1143
rect 17220 1217 17290 1225
rect 17220 1215 17265 1217
rect 17220 1143 17225 1215
rect 17245 1145 17265 1215
rect 17285 1145 17290 1217
rect 17245 1143 17290 1145
rect 17220 1135 17290 1143
rect 17470 1217 17540 1225
rect 17470 1195 17475 1217
rect 17495 1215 17540 1217
rect 17495 1195 17515 1215
rect 17535 1195 17540 1215
rect 17470 1165 17540 1195
rect 17470 1145 17475 1165
rect 17495 1145 17515 1165
rect 17535 1145 17540 1165
rect 17470 1135 17540 1145
rect 17565 1215 17595 1225
rect 17565 1195 17570 1215
rect 17590 1195 17595 1215
rect 17565 1165 17595 1195
rect 17565 1145 17570 1165
rect 17590 1145 17595 1165
rect 17565 1135 17595 1145
rect 17620 1215 17650 1255
rect 17670 1275 17710 1285
rect 17670 1255 17680 1275
rect 17700 1255 17710 1275
rect 17670 1245 17710 1255
rect 17730 1275 17760 1285
rect 17730 1255 17735 1275
rect 17755 1255 17760 1275
rect 17680 1225 17700 1245
rect 17620 1195 17625 1215
rect 17645 1195 17650 1215
rect 17620 1165 17650 1195
rect 17620 1145 17625 1165
rect 17645 1145 17650 1165
rect 17620 1135 17650 1145
rect 17675 1215 17705 1225
rect 17675 1195 17680 1215
rect 17700 1195 17705 1215
rect 17675 1165 17705 1195
rect 17675 1145 17680 1165
rect 17700 1145 17705 1165
rect 17675 1135 17705 1145
rect 17730 1215 17760 1255
rect 17780 1275 17820 1285
rect 17780 1255 17790 1275
rect 17810 1255 17820 1275
rect 17780 1245 17820 1255
rect 17840 1275 17870 1285
rect 17840 1255 17845 1275
rect 17865 1255 17870 1275
rect 17790 1225 17810 1245
rect 17730 1195 17735 1215
rect 17755 1195 17760 1215
rect 17730 1165 17760 1195
rect 17730 1145 17735 1165
rect 17755 1145 17760 1165
rect 17730 1135 17760 1145
rect 17785 1215 17815 1225
rect 17785 1195 17790 1215
rect 17810 1195 17815 1215
rect 17785 1165 17815 1195
rect 17785 1145 17790 1165
rect 17810 1145 17815 1165
rect 17785 1135 17815 1145
rect 17840 1215 17870 1255
rect 17890 1275 17930 1285
rect 17890 1255 17900 1275
rect 17920 1255 17930 1275
rect 17890 1245 17930 1255
rect 17950 1275 17980 1285
rect 17950 1255 17955 1275
rect 17975 1255 17980 1275
rect 17900 1225 17920 1245
rect 17840 1195 17845 1215
rect 17865 1195 17870 1215
rect 17840 1165 17870 1195
rect 17840 1145 17845 1165
rect 17865 1145 17870 1165
rect 17840 1135 17870 1145
rect 17895 1215 17925 1225
rect 17895 1195 17900 1215
rect 17920 1195 17925 1215
rect 17895 1165 17925 1195
rect 17895 1145 17900 1165
rect 17920 1145 17925 1165
rect 17895 1135 17925 1145
rect 17950 1215 17980 1255
rect 18000 1275 18040 1285
rect 18000 1255 18010 1275
rect 18030 1255 18040 1275
rect 18000 1245 18040 1255
rect 18065 1275 18105 1285
rect 18065 1255 18075 1275
rect 18095 1255 18105 1275
rect 18065 1245 18105 1255
rect 18345 1275 18385 1285
rect 18345 1255 18355 1275
rect 18375 1255 18385 1275
rect 18345 1245 18385 1255
rect 18455 1275 18495 1285
rect 18455 1255 18465 1275
rect 18485 1255 18495 1275
rect 18455 1245 18495 1255
rect 18515 1275 18545 1285
rect 18515 1255 18520 1275
rect 18540 1255 18545 1275
rect 18515 1245 18545 1255
rect 18565 1275 18605 1285
rect 18565 1255 18575 1275
rect 18595 1255 18605 1275
rect 18565 1245 18605 1255
rect 18625 1275 18655 1285
rect 18625 1255 18630 1275
rect 18650 1255 18655 1275
rect 18625 1245 18655 1255
rect 18675 1275 18715 1285
rect 18675 1255 18685 1275
rect 18705 1255 18715 1275
rect 18675 1245 18715 1255
rect 18010 1225 18030 1245
rect 18065 1225 18085 1245
rect 18355 1225 18375 1245
rect 18465 1225 18485 1245
rect 18575 1225 18595 1245
rect 18630 1225 18650 1245
rect 18685 1225 18705 1245
rect 17950 1195 17955 1215
rect 17975 1195 17980 1215
rect 17950 1165 17980 1195
rect 17950 1145 17955 1165
rect 17975 1145 17980 1165
rect 17950 1135 17980 1145
rect 18005 1215 18035 1225
rect 18005 1195 18010 1215
rect 18030 1195 18035 1215
rect 18005 1165 18035 1195
rect 18005 1145 18010 1165
rect 18030 1145 18035 1165
rect 18005 1135 18035 1145
rect 18060 1217 18130 1225
rect 18060 1215 18105 1217
rect 18060 1195 18065 1215
rect 18085 1195 18105 1215
rect 18125 1195 18130 1217
rect 18060 1165 18130 1195
rect 18060 1145 18065 1165
rect 18085 1145 18105 1165
rect 18125 1145 18130 1165
rect 18060 1135 18130 1145
rect 18310 1217 18380 1225
rect 18310 1145 18315 1217
rect 18335 1215 18380 1217
rect 18335 1145 18355 1215
rect 18375 1145 18380 1215
rect 18310 1135 18380 1145
rect 18405 1215 18435 1225
rect 18405 1145 18410 1215
rect 18430 1145 18435 1215
rect 18405 1135 18435 1145
rect 18460 1215 18490 1225
rect 18460 1145 18465 1215
rect 18485 1145 18490 1215
rect 18460 1135 18490 1145
rect 18515 1215 18545 1225
rect 18515 1145 18520 1215
rect 18540 1145 18545 1215
rect 18515 1135 18545 1145
rect 18570 1215 18600 1225
rect 18570 1145 18575 1215
rect 18595 1145 18600 1215
rect 18570 1135 18600 1145
rect 18625 1215 18655 1225
rect 18625 1145 18630 1215
rect 18650 1145 18655 1215
rect 18625 1135 18655 1145
rect 18680 1217 18750 1225
rect 18680 1215 18725 1217
rect 18680 1145 18685 1215
rect 18705 1145 18725 1215
rect 18745 1145 18750 1217
rect 18680 1135 18750 1145
rect 16440 1115 16460 1135
rect 16550 1115 16570 1135
rect 16950 1115 16970 1135
rect 17060 1115 17080 1135
rect 17170 1115 17190 1135
rect 17625 1115 17645 1135
rect 17735 1115 17755 1135
rect 17845 1115 17865 1135
rect 17955 1115 17975 1135
rect 18410 1115 18430 1135
rect 18520 1115 18540 1135
rect 18630 1115 18650 1135
rect 16430 1105 16470 1115
rect 16430 1085 16440 1105
rect 16460 1085 16470 1105
rect 16430 1075 16470 1085
rect 16540 1105 16580 1115
rect 16540 1085 16550 1105
rect 16570 1085 16580 1105
rect 16540 1075 16580 1085
rect 16940 1105 16980 1115
rect 16940 1085 16950 1105
rect 16970 1085 16980 1105
rect 16940 1075 16980 1085
rect 17050 1105 17090 1115
rect 17050 1085 17060 1105
rect 17080 1085 17090 1105
rect 17050 1075 17090 1085
rect 17160 1105 17200 1115
rect 17160 1085 17170 1105
rect 17190 1085 17200 1105
rect 17160 1075 17200 1085
rect 17615 1105 17655 1115
rect 17615 1085 17625 1105
rect 17645 1085 17655 1105
rect 17615 1075 17655 1085
rect 17725 1105 17765 1115
rect 17725 1085 17735 1105
rect 17755 1085 17765 1105
rect 17725 1075 17765 1085
rect 17835 1105 17875 1115
rect 17835 1085 17845 1105
rect 17865 1085 17875 1105
rect 17835 1075 17875 1085
rect 17945 1105 17985 1115
rect 17945 1085 17955 1105
rect 17975 1085 17985 1105
rect 17945 1075 17985 1085
rect 18400 1105 18440 1115
rect 18400 1085 18410 1105
rect 18430 1085 18440 1105
rect 18400 1075 18440 1085
rect 18510 1105 18550 1115
rect 18510 1085 18520 1105
rect 18540 1085 18550 1105
rect 18510 1075 18550 1085
rect 18620 1105 18660 1115
rect 18620 1085 18630 1105
rect 18650 1085 18660 1105
rect 18620 1075 18660 1085
rect 16970 810 17010 820
rect 16970 790 16980 810
rect 17000 790 17010 810
rect 16970 780 17010 790
rect 17150 810 17190 820
rect 17150 790 17160 810
rect 17180 790 17190 810
rect 17150 780 17190 790
rect 17330 810 17370 820
rect 17330 790 17340 810
rect 17360 790 17370 810
rect 17330 780 17370 790
rect 17510 810 17550 820
rect 17510 790 17520 810
rect 17540 790 17550 810
rect 17510 780 17550 790
rect 17690 810 17730 820
rect 17690 790 17700 810
rect 17720 790 17730 810
rect 17690 780 17730 790
rect 17870 810 17910 820
rect 17870 790 17880 810
rect 17900 790 17910 810
rect 17870 780 17910 790
rect 18050 810 18090 820
rect 18050 790 18060 810
rect 18080 790 18090 810
rect 18050 780 18090 790
rect 18230 810 18270 820
rect 18230 790 18240 810
rect 18260 790 18270 810
rect 18230 780 18270 790
rect 18410 810 18450 820
rect 18410 790 18420 810
rect 18440 790 18450 810
rect 18410 780 18450 790
rect 18590 810 18630 820
rect 18590 790 18600 810
rect 18620 790 18630 810
rect 18590 780 18630 790
rect 18905 810 18945 820
rect 18905 790 18915 810
rect 18935 790 18945 810
rect 18905 780 18945 790
rect 19015 810 19055 820
rect 19015 790 19025 810
rect 19045 790 19055 810
rect 19015 780 19055 790
rect 19075 810 19115 820
rect 19075 790 19085 810
rect 19105 790 19115 810
rect 19075 780 19115 790
rect 16980 760 17000 780
rect 17160 760 17180 780
rect 17340 760 17360 780
rect 17520 760 17540 780
rect 17700 760 17720 780
rect 17880 760 17900 780
rect 18060 760 18080 780
rect 18240 760 18260 780
rect 18420 760 18440 780
rect 18600 760 18620 780
rect 18915 760 18935 780
rect 19025 760 19045 780
rect 19080 760 19100 780
rect 16935 750 17005 760
rect 16935 730 16940 750
rect 16960 730 16980 750
rect 17000 730 17005 750
rect 16440 710 16470 720
rect 16440 690 16445 710
rect 16465 690 16470 710
rect 16440 660 16470 690
rect 16545 710 16585 720
rect 16545 690 16555 710
rect 16575 690 16585 710
rect 16545 680 16585 690
rect 16655 710 16695 720
rect 16655 690 16665 710
rect 16685 690 16695 710
rect 16655 680 16695 690
rect 16935 700 17005 730
rect 16935 680 16940 700
rect 16960 680 16980 700
rect 17000 680 17005 700
rect 16555 660 16575 680
rect 16660 660 16690 680
rect 16400 650 16470 660
rect 16400 630 16405 650
rect 16425 630 16445 650
rect 16465 630 16470 650
rect 16400 600 16470 630
rect 16400 580 16405 600
rect 16425 580 16445 600
rect 16465 580 16470 600
rect 16400 570 16470 580
rect 16495 650 16525 660
rect 16495 630 16500 650
rect 16520 630 16525 650
rect 16495 600 16525 630
rect 16495 580 16500 600
rect 16520 580 16525 600
rect 16495 570 16525 580
rect 16550 650 16580 660
rect 16550 630 16555 650
rect 16575 630 16580 650
rect 16550 600 16580 630
rect 16550 580 16555 600
rect 16575 580 16580 600
rect 16550 570 16580 580
rect 16605 650 16635 660
rect 16605 630 16610 650
rect 16630 630 16635 650
rect 16605 600 16635 630
rect 16605 580 16610 600
rect 16630 580 16635 600
rect 16605 570 16635 580
rect 16660 650 16735 660
rect 16660 630 16665 650
rect 16685 630 16710 650
rect 16730 630 16735 650
rect 16660 600 16735 630
rect 16660 580 16665 600
rect 16685 580 16710 600
rect 16730 580 16735 600
rect 16660 570 16735 580
rect 16935 650 17005 680
rect 16935 630 16940 650
rect 16960 630 16980 650
rect 17000 630 17005 650
rect 16935 600 17005 630
rect 16935 580 16940 600
rect 16960 580 16980 600
rect 17000 580 17005 600
rect 16500 550 16520 570
rect 16610 550 16630 570
rect 16935 550 17005 580
rect 16480 540 16520 550
rect 16480 520 16490 540
rect 16510 520 16520 540
rect 16480 510 16520 520
rect 16545 540 16585 550
rect 16545 520 16555 540
rect 16575 520 16585 540
rect 16545 510 16585 520
rect 16610 540 16650 550
rect 16610 520 16620 540
rect 16640 520 16650 540
rect 16610 510 16650 520
rect 16935 530 16940 550
rect 16960 530 16980 550
rect 17000 530 17005 550
rect 16935 500 17005 530
rect 16935 480 16940 500
rect 16960 480 16980 500
rect 17000 480 17005 500
rect 16935 470 17005 480
rect 17065 750 17095 760
rect 17065 730 17070 750
rect 17090 730 17095 750
rect 17065 700 17095 730
rect 17065 680 17070 700
rect 17090 680 17095 700
rect 17065 650 17095 680
rect 17065 630 17070 650
rect 17090 630 17095 650
rect 17065 600 17095 630
rect 17065 580 17070 600
rect 17090 580 17095 600
rect 17065 550 17095 580
rect 17065 530 17070 550
rect 17090 530 17095 550
rect 17065 500 17095 530
rect 17065 480 17070 500
rect 17090 480 17095 500
rect 17065 470 17095 480
rect 17155 750 17185 760
rect 17155 730 17160 750
rect 17180 730 17185 750
rect 17155 700 17185 730
rect 17155 680 17160 700
rect 17180 680 17185 700
rect 17155 650 17185 680
rect 17155 630 17160 650
rect 17180 630 17185 650
rect 17155 600 17185 630
rect 17155 580 17160 600
rect 17180 580 17185 600
rect 17155 550 17185 580
rect 17155 530 17160 550
rect 17180 530 17185 550
rect 17155 500 17185 530
rect 17155 480 17160 500
rect 17180 480 17185 500
rect 17155 470 17185 480
rect 17245 750 17275 760
rect 17245 730 17250 750
rect 17270 730 17275 750
rect 17245 700 17275 730
rect 17245 680 17250 700
rect 17270 680 17275 700
rect 17245 650 17275 680
rect 17245 630 17250 650
rect 17270 630 17275 650
rect 17245 600 17275 630
rect 17245 580 17250 600
rect 17270 580 17275 600
rect 17245 550 17275 580
rect 17245 530 17250 550
rect 17270 530 17275 550
rect 17245 500 17275 530
rect 17245 480 17250 500
rect 17270 480 17275 500
rect 17245 470 17275 480
rect 17335 750 17365 760
rect 17335 730 17340 750
rect 17360 730 17365 750
rect 17335 700 17365 730
rect 17335 680 17340 700
rect 17360 680 17365 700
rect 17335 650 17365 680
rect 17335 630 17340 650
rect 17360 630 17365 650
rect 17335 600 17365 630
rect 17335 580 17340 600
rect 17360 580 17365 600
rect 17335 550 17365 580
rect 17335 530 17340 550
rect 17360 530 17365 550
rect 17335 500 17365 530
rect 17335 480 17340 500
rect 17360 480 17365 500
rect 17335 470 17365 480
rect 17425 750 17455 760
rect 17425 730 17430 750
rect 17450 730 17455 750
rect 17425 700 17455 730
rect 17425 680 17430 700
rect 17450 680 17455 700
rect 17425 650 17455 680
rect 17425 630 17430 650
rect 17450 630 17455 650
rect 17425 600 17455 630
rect 17425 580 17430 600
rect 17450 580 17455 600
rect 17425 550 17455 580
rect 17425 530 17430 550
rect 17450 530 17455 550
rect 17425 500 17455 530
rect 17425 480 17430 500
rect 17450 480 17455 500
rect 17425 470 17455 480
rect 17515 750 17545 760
rect 17515 730 17520 750
rect 17540 730 17545 750
rect 17515 700 17545 730
rect 17515 680 17520 700
rect 17540 680 17545 700
rect 17515 650 17545 680
rect 17515 630 17520 650
rect 17540 630 17545 650
rect 17515 600 17545 630
rect 17515 580 17520 600
rect 17540 580 17545 600
rect 17515 550 17545 580
rect 17515 530 17520 550
rect 17540 530 17545 550
rect 17515 500 17545 530
rect 17515 480 17520 500
rect 17540 480 17545 500
rect 17515 470 17545 480
rect 17605 750 17635 760
rect 17605 730 17610 750
rect 17630 730 17635 750
rect 17605 700 17635 730
rect 17605 680 17610 700
rect 17630 680 17635 700
rect 17605 650 17635 680
rect 17605 630 17610 650
rect 17630 630 17635 650
rect 17605 600 17635 630
rect 17605 580 17610 600
rect 17630 580 17635 600
rect 17605 550 17635 580
rect 17605 530 17610 550
rect 17630 530 17635 550
rect 17605 500 17635 530
rect 17605 480 17610 500
rect 17630 480 17635 500
rect 17605 470 17635 480
rect 17695 750 17725 760
rect 17695 730 17700 750
rect 17720 730 17725 750
rect 17695 700 17725 730
rect 17695 680 17700 700
rect 17720 680 17725 700
rect 17695 650 17725 680
rect 17695 630 17700 650
rect 17720 630 17725 650
rect 17695 600 17725 630
rect 17695 580 17700 600
rect 17720 580 17725 600
rect 17695 550 17725 580
rect 17695 530 17700 550
rect 17720 530 17725 550
rect 17695 500 17725 530
rect 17695 480 17700 500
rect 17720 480 17725 500
rect 17695 470 17725 480
rect 17785 750 17815 760
rect 17785 730 17790 750
rect 17810 730 17815 750
rect 17785 700 17815 730
rect 17785 680 17790 700
rect 17810 680 17815 700
rect 17785 650 17815 680
rect 17785 630 17790 650
rect 17810 630 17815 650
rect 17785 600 17815 630
rect 17785 580 17790 600
rect 17810 580 17815 600
rect 17785 550 17815 580
rect 17785 530 17790 550
rect 17810 530 17815 550
rect 17785 500 17815 530
rect 17785 480 17790 500
rect 17810 480 17815 500
rect 17785 470 17815 480
rect 17875 750 17905 760
rect 17875 730 17880 750
rect 17900 730 17905 750
rect 17875 700 17905 730
rect 17875 680 17880 700
rect 17900 680 17905 700
rect 17875 650 17905 680
rect 17875 630 17880 650
rect 17900 630 17905 650
rect 17875 600 17905 630
rect 17875 580 17880 600
rect 17900 580 17905 600
rect 17875 550 17905 580
rect 17875 530 17880 550
rect 17900 530 17905 550
rect 17875 500 17905 530
rect 17875 480 17880 500
rect 17900 480 17905 500
rect 17875 470 17905 480
rect 17965 750 17995 760
rect 17965 730 17970 750
rect 17990 730 17995 750
rect 17965 700 17995 730
rect 17965 680 17970 700
rect 17990 680 17995 700
rect 17965 650 17995 680
rect 17965 630 17970 650
rect 17990 630 17995 650
rect 17965 600 17995 630
rect 17965 580 17970 600
rect 17990 580 17995 600
rect 17965 550 17995 580
rect 17965 530 17970 550
rect 17990 530 17995 550
rect 17965 500 17995 530
rect 17965 480 17970 500
rect 17990 480 17995 500
rect 17965 470 17995 480
rect 18055 750 18085 760
rect 18055 730 18060 750
rect 18080 730 18085 750
rect 18055 700 18085 730
rect 18055 680 18060 700
rect 18080 680 18085 700
rect 18055 650 18085 680
rect 18055 630 18060 650
rect 18080 630 18085 650
rect 18055 600 18085 630
rect 18055 580 18060 600
rect 18080 580 18085 600
rect 18055 550 18085 580
rect 18055 530 18060 550
rect 18080 530 18085 550
rect 18055 500 18085 530
rect 18055 480 18060 500
rect 18080 480 18085 500
rect 18055 470 18085 480
rect 18145 750 18175 760
rect 18145 730 18150 750
rect 18170 730 18175 750
rect 18145 700 18175 730
rect 18145 680 18150 700
rect 18170 680 18175 700
rect 18145 650 18175 680
rect 18145 630 18150 650
rect 18170 630 18175 650
rect 18145 600 18175 630
rect 18145 580 18150 600
rect 18170 580 18175 600
rect 18145 550 18175 580
rect 18145 530 18150 550
rect 18170 530 18175 550
rect 18145 500 18175 530
rect 18145 480 18150 500
rect 18170 480 18175 500
rect 18145 470 18175 480
rect 18235 750 18265 760
rect 18235 730 18240 750
rect 18260 730 18265 750
rect 18235 700 18265 730
rect 18235 680 18240 700
rect 18260 680 18265 700
rect 18235 650 18265 680
rect 18235 630 18240 650
rect 18260 630 18265 650
rect 18235 600 18265 630
rect 18235 580 18240 600
rect 18260 580 18265 600
rect 18235 550 18265 580
rect 18235 530 18240 550
rect 18260 530 18265 550
rect 18235 500 18265 530
rect 18235 480 18240 500
rect 18260 480 18265 500
rect 18235 470 18265 480
rect 18325 750 18355 760
rect 18325 730 18330 750
rect 18350 730 18355 750
rect 18325 700 18355 730
rect 18325 680 18330 700
rect 18350 680 18355 700
rect 18325 650 18355 680
rect 18325 630 18330 650
rect 18350 630 18355 650
rect 18325 600 18355 630
rect 18325 580 18330 600
rect 18350 580 18355 600
rect 18325 550 18355 580
rect 18325 530 18330 550
rect 18350 530 18355 550
rect 18325 500 18355 530
rect 18325 480 18330 500
rect 18350 480 18355 500
rect 18325 470 18355 480
rect 18415 750 18445 760
rect 18415 730 18420 750
rect 18440 730 18445 750
rect 18415 700 18445 730
rect 18415 680 18420 700
rect 18440 680 18445 700
rect 18415 650 18445 680
rect 18415 630 18420 650
rect 18440 630 18445 650
rect 18415 600 18445 630
rect 18415 580 18420 600
rect 18440 580 18445 600
rect 18415 550 18445 580
rect 18415 530 18420 550
rect 18440 530 18445 550
rect 18415 500 18445 530
rect 18415 480 18420 500
rect 18440 480 18445 500
rect 18415 470 18445 480
rect 18505 750 18535 760
rect 18505 730 18510 750
rect 18530 730 18535 750
rect 18505 700 18535 730
rect 18505 680 18510 700
rect 18530 680 18535 700
rect 18505 650 18535 680
rect 18505 630 18510 650
rect 18530 630 18535 650
rect 18505 600 18535 630
rect 18505 580 18510 600
rect 18530 580 18535 600
rect 18505 550 18535 580
rect 18505 530 18510 550
rect 18530 530 18535 550
rect 18505 500 18535 530
rect 18505 480 18510 500
rect 18530 480 18535 500
rect 18505 470 18535 480
rect 18595 750 18665 760
rect 18595 730 18600 750
rect 18620 730 18640 750
rect 18660 730 18665 750
rect 18595 700 18665 730
rect 18595 680 18600 700
rect 18620 680 18640 700
rect 18660 680 18665 700
rect 18595 650 18665 680
rect 18595 630 18600 650
rect 18620 630 18640 650
rect 18660 630 18665 650
rect 18595 600 18665 630
rect 18595 580 18600 600
rect 18620 580 18640 600
rect 18660 580 18665 600
rect 18595 550 18665 580
rect 18870 750 18940 760
rect 18870 730 18875 750
rect 18895 730 18915 750
rect 18935 730 18940 750
rect 18870 700 18940 730
rect 18870 680 18875 700
rect 18895 680 18915 700
rect 18935 680 18940 700
rect 18870 650 18940 680
rect 18870 630 18875 650
rect 18895 630 18915 650
rect 18935 630 18940 650
rect 18870 600 18940 630
rect 18870 580 18875 600
rect 18895 580 18915 600
rect 18935 580 18940 600
rect 18870 570 18940 580
rect 18965 750 18995 760
rect 18965 730 18970 750
rect 18990 730 18995 750
rect 18965 700 18995 730
rect 18965 680 18970 700
rect 18990 680 18995 700
rect 18965 650 18995 680
rect 18965 630 18970 650
rect 18990 630 18995 650
rect 18965 600 18995 630
rect 18965 580 18970 600
rect 18990 580 18995 600
rect 18965 570 18995 580
rect 19020 750 19050 760
rect 19020 730 19025 750
rect 19045 730 19050 750
rect 19020 700 19050 730
rect 19020 680 19025 700
rect 19045 680 19050 700
rect 19020 650 19050 680
rect 19020 630 19025 650
rect 19045 630 19050 650
rect 19020 600 19050 630
rect 19020 580 19025 600
rect 19045 580 19050 600
rect 19020 570 19050 580
rect 19075 750 19145 760
rect 19075 730 19080 750
rect 19100 730 19120 750
rect 19140 730 19145 750
rect 19075 700 19145 730
rect 19075 680 19080 700
rect 19100 680 19120 700
rect 19140 680 19145 700
rect 19075 650 19145 680
rect 19075 630 19080 650
rect 19100 630 19120 650
rect 19140 630 19145 650
rect 19075 600 19145 630
rect 19075 580 19080 600
rect 19100 580 19120 600
rect 19140 580 19145 600
rect 19075 570 19145 580
rect 18970 550 18990 570
rect 18595 530 18600 550
rect 18620 530 18640 550
rect 18660 530 18665 550
rect 18595 500 18665 530
rect 18950 540 18990 550
rect 18950 520 18960 540
rect 18980 520 18990 540
rect 18950 510 18990 520
rect 18595 480 18600 500
rect 18620 480 18640 500
rect 18660 480 18665 500
rect 18595 470 18665 480
rect 19000 490 19040 495
rect 19000 470 19010 490
rect 19030 470 19040 490
rect 17070 450 17090 470
rect 17250 450 17270 470
rect 17430 450 17450 470
rect 17610 450 17630 470
rect 17790 450 17810 470
rect 17970 450 17990 470
rect 18150 450 18170 470
rect 18330 450 18350 470
rect 18510 450 18530 470
rect 19000 465 19040 470
rect 17060 440 17100 450
rect 17060 420 17070 440
rect 17090 420 17100 440
rect 17060 410 17100 420
rect 17240 440 17280 450
rect 17240 420 17250 440
rect 17270 420 17280 440
rect 17240 410 17280 420
rect 17420 440 17460 450
rect 17420 420 17430 440
rect 17450 420 17460 440
rect 17420 410 17460 420
rect 17600 440 17640 450
rect 17600 420 17610 440
rect 17630 420 17640 440
rect 17600 410 17640 420
rect 17690 440 17730 450
rect 17690 420 17700 440
rect 17720 420 17730 440
rect 17690 410 17730 420
rect 17780 440 17820 450
rect 17780 420 17790 440
rect 17810 420 17820 440
rect 17780 410 17820 420
rect 17960 440 18000 450
rect 17960 420 17970 440
rect 17990 420 18000 440
rect 17960 410 18000 420
rect 18140 440 18180 450
rect 18140 420 18150 440
rect 18170 420 18180 440
rect 18140 410 18180 420
rect 18320 440 18360 450
rect 18320 420 18330 440
rect 18350 420 18360 440
rect 18320 410 18360 420
rect 18410 440 18450 450
rect 18410 420 18420 440
rect 18440 420 18450 440
rect 18410 410 18450 420
rect 18500 440 18540 450
rect 18500 420 18510 440
rect 18530 420 18540 440
rect 18500 410 18540 420
rect 16425 -30 16455 -20
rect 16425 -50 16430 -30
rect 16450 -50 16455 -30
rect 16425 -80 16455 -50
rect 16480 -30 16520 -20
rect 16480 -50 16490 -30
rect 16510 -50 16520 -30
rect 16480 -60 16520 -50
rect 16545 -30 16575 -20
rect 16545 -50 16550 -30
rect 16570 -50 16575 -30
rect 16545 -60 16575 -50
rect 16665 -30 16695 -20
rect 16665 -50 16670 -30
rect 16690 -50 16695 -30
rect 16665 -60 16695 -50
rect 16785 -30 16815 -20
rect 16785 -50 16790 -30
rect 16810 -50 16815 -30
rect 16785 -60 16815 -50
rect 16840 -30 16880 -20
rect 16840 -50 16850 -30
rect 16870 -50 16880 -30
rect 16840 -60 16880 -50
rect 16905 -30 16935 -20
rect 16905 -50 16910 -30
rect 16930 -50 16935 -30
rect 16905 -60 16935 -50
rect 17025 -30 17055 -20
rect 17025 -50 17030 -30
rect 17050 -50 17055 -30
rect 17025 -60 17055 -50
rect 17145 -30 17175 -20
rect 17145 -50 17150 -30
rect 17170 -50 17175 -30
rect 17145 -60 17175 -50
rect 17200 -30 17240 -20
rect 17200 -50 17210 -30
rect 17230 -50 17240 -30
rect 17200 -60 17240 -50
rect 17265 -30 17295 -20
rect 17265 -50 17270 -30
rect 17290 -50 17295 -30
rect 17265 -60 17295 -50
rect 17385 -30 17415 -20
rect 17385 -50 17390 -30
rect 17410 -50 17415 -30
rect 17385 -60 17415 -50
rect 17505 -30 17535 -20
rect 17505 -50 17510 -30
rect 17530 -50 17535 -30
rect 17505 -60 17535 -50
rect 17560 -30 17600 -20
rect 17560 -50 17570 -30
rect 17590 -50 17600 -30
rect 17560 -60 17600 -50
rect 17625 -30 17655 -20
rect 17625 -50 17630 -30
rect 17650 -50 17655 -30
rect 16490 -80 16510 -60
rect 16550 -80 16570 -60
rect 16670 -80 16690 -60
rect 16790 -80 16810 -60
rect 16850 -80 16870 -60
rect 16910 -80 16930 -60
rect 17030 -80 17050 -60
rect 17150 -80 17170 -60
rect 17210 -80 17230 -60
rect 17270 -80 17290 -60
rect 17390 -80 17410 -60
rect 17510 -80 17530 -60
rect 17570 -80 17590 -60
rect 17625 -80 17655 -50
rect 17945 -30 17975 -20
rect 17945 -50 17950 -30
rect 17970 -50 17975 -30
rect 17945 -80 17975 -50
rect 18000 -30 18040 -20
rect 18000 -50 18010 -30
rect 18030 -50 18040 -30
rect 18000 -60 18040 -50
rect 18065 -30 18095 -20
rect 18065 -50 18070 -30
rect 18090 -50 18095 -30
rect 18065 -60 18095 -50
rect 18185 -30 18215 -20
rect 18185 -50 18190 -30
rect 18210 -50 18215 -30
rect 18185 -60 18215 -50
rect 18305 -30 18335 -20
rect 18305 -50 18310 -30
rect 18330 -50 18335 -30
rect 18305 -60 18335 -50
rect 18360 -30 18400 -20
rect 18360 -50 18370 -30
rect 18390 -50 18400 -30
rect 18360 -60 18400 -50
rect 18425 -30 18455 -20
rect 18425 -50 18430 -30
rect 18450 -50 18455 -30
rect 18425 -60 18455 -50
rect 18545 -30 18575 -20
rect 18545 -50 18550 -30
rect 18570 -50 18575 -30
rect 18545 -60 18575 -50
rect 18665 -30 18695 -20
rect 18665 -50 18670 -30
rect 18690 -50 18695 -30
rect 18665 -60 18695 -50
rect 18720 -30 18760 -20
rect 18720 -50 18730 -30
rect 18750 -50 18760 -30
rect 18720 -60 18760 -50
rect 18785 -30 18815 -20
rect 18785 -50 18790 -30
rect 18810 -50 18815 -30
rect 18785 -60 18815 -50
rect 18905 -30 18935 -20
rect 18905 -50 18910 -30
rect 18930 -50 18935 -30
rect 18905 -60 18935 -50
rect 19025 -30 19055 -20
rect 19025 -50 19030 -30
rect 19050 -50 19055 -30
rect 19025 -60 19055 -50
rect 19080 -30 19120 -20
rect 19080 -50 19090 -30
rect 19110 -50 19120 -30
rect 19080 -60 19120 -50
rect 19145 -30 19175 -20
rect 19145 -50 19150 -30
rect 19170 -50 19175 -30
rect 18010 -80 18030 -60
rect 18070 -80 18090 -60
rect 18190 -80 18210 -60
rect 18310 -80 18330 -60
rect 18370 -80 18390 -60
rect 18430 -80 18450 -60
rect 18550 -80 18570 -60
rect 18670 -80 18690 -60
rect 18730 -80 18750 -60
rect 18790 -80 18810 -60
rect 18910 -80 18930 -60
rect 19030 -80 19050 -60
rect 19090 -80 19110 -60
rect 19145 -80 19175 -50
rect 16385 -90 16455 -80
rect 16385 -110 16390 -90
rect 16410 -110 16430 -90
rect 16450 -110 16455 -90
rect 16385 -140 16455 -110
rect 16385 -160 16390 -140
rect 16410 -160 16430 -140
rect 16450 -160 16455 -140
rect 16385 -170 16455 -160
rect 16485 -90 16515 -80
rect 16485 -110 16490 -90
rect 16510 -110 16515 -90
rect 16485 -140 16515 -110
rect 16485 -160 16490 -140
rect 16510 -160 16515 -140
rect 16485 -170 16515 -160
rect 16545 -90 16575 -80
rect 16545 -110 16550 -90
rect 16570 -110 16575 -90
rect 16545 -140 16575 -110
rect 16545 -160 16550 -140
rect 16570 -160 16575 -140
rect 16545 -170 16575 -160
rect 16605 -90 16635 -80
rect 16605 -110 16610 -90
rect 16630 -110 16635 -90
rect 16605 -140 16635 -110
rect 16605 -160 16610 -140
rect 16630 -160 16635 -140
rect 16605 -170 16635 -160
rect 16665 -90 16695 -80
rect 16665 -110 16670 -90
rect 16690 -110 16695 -90
rect 16665 -140 16695 -110
rect 16665 -160 16670 -140
rect 16690 -160 16695 -140
rect 16665 -170 16695 -160
rect 16725 -90 16755 -80
rect 16725 -110 16730 -90
rect 16750 -110 16755 -90
rect 16725 -140 16755 -110
rect 16725 -160 16730 -140
rect 16750 -160 16755 -140
rect 16725 -170 16755 -160
rect 16785 -90 16815 -80
rect 16785 -110 16790 -90
rect 16810 -110 16815 -90
rect 16785 -140 16815 -110
rect 16785 -160 16790 -140
rect 16810 -160 16815 -140
rect 16785 -170 16815 -160
rect 16845 -90 16875 -80
rect 16845 -110 16850 -90
rect 16870 -110 16875 -90
rect 16845 -140 16875 -110
rect 16845 -160 16850 -140
rect 16870 -160 16875 -140
rect 16845 -170 16875 -160
rect 16905 -90 16935 -80
rect 16905 -110 16910 -90
rect 16930 -110 16935 -90
rect 16905 -140 16935 -110
rect 16905 -160 16910 -140
rect 16930 -160 16935 -140
rect 16905 -170 16935 -160
rect 16965 -90 16995 -80
rect 16965 -110 16970 -90
rect 16990 -110 16995 -90
rect 16965 -140 16995 -110
rect 16965 -160 16970 -140
rect 16990 -160 16995 -140
rect 16965 -170 16995 -160
rect 17025 -90 17055 -80
rect 17025 -110 17030 -90
rect 17050 -110 17055 -90
rect 17025 -140 17055 -110
rect 17025 -160 17030 -140
rect 17050 -160 17055 -140
rect 17025 -170 17055 -160
rect 17085 -90 17115 -80
rect 17085 -110 17090 -90
rect 17110 -110 17115 -90
rect 17085 -140 17115 -110
rect 17085 -160 17090 -140
rect 17110 -160 17115 -140
rect 17085 -170 17115 -160
rect 17145 -90 17175 -80
rect 17145 -110 17150 -90
rect 17170 -110 17175 -90
rect 17145 -140 17175 -110
rect 17145 -160 17150 -140
rect 17170 -160 17175 -140
rect 17145 -170 17175 -160
rect 17205 -90 17235 -80
rect 17205 -110 17210 -90
rect 17230 -110 17235 -90
rect 17205 -140 17235 -110
rect 17205 -160 17210 -140
rect 17230 -160 17235 -140
rect 17205 -170 17235 -160
rect 17265 -90 17295 -80
rect 17265 -110 17270 -90
rect 17290 -110 17295 -90
rect 17265 -140 17295 -110
rect 17265 -160 17270 -140
rect 17290 -160 17295 -140
rect 17265 -170 17295 -160
rect 17325 -90 17355 -80
rect 17325 -110 17330 -90
rect 17350 -110 17355 -90
rect 17325 -140 17355 -110
rect 17325 -160 17330 -140
rect 17350 -160 17355 -140
rect 17325 -170 17355 -160
rect 17385 -90 17415 -80
rect 17385 -110 17390 -90
rect 17410 -110 17415 -90
rect 17385 -140 17415 -110
rect 17385 -160 17390 -140
rect 17410 -160 17415 -140
rect 17385 -170 17415 -160
rect 17445 -90 17475 -80
rect 17445 -110 17450 -90
rect 17470 -110 17475 -90
rect 17445 -140 17475 -110
rect 17445 -160 17450 -140
rect 17470 -160 17475 -140
rect 17445 -170 17475 -160
rect 17505 -90 17535 -80
rect 17505 -110 17510 -90
rect 17530 -110 17535 -90
rect 17505 -140 17535 -110
rect 17505 -160 17510 -140
rect 17530 -160 17535 -140
rect 17505 -170 17535 -160
rect 17565 -90 17595 -80
rect 17565 -110 17570 -90
rect 17590 -110 17595 -90
rect 17565 -140 17595 -110
rect 17565 -160 17570 -140
rect 17590 -160 17595 -140
rect 17565 -170 17595 -160
rect 17625 -90 17695 -80
rect 17625 -110 17630 -90
rect 17650 -110 17670 -90
rect 17690 -110 17695 -90
rect 17625 -140 17695 -110
rect 17625 -160 17630 -140
rect 17650 -160 17670 -140
rect 17690 -160 17695 -140
rect 17625 -170 17695 -160
rect 17905 -90 17975 -80
rect 17905 -110 17910 -90
rect 17930 -110 17950 -90
rect 17970 -110 17975 -90
rect 17905 -140 17975 -110
rect 17905 -160 17910 -140
rect 17930 -160 17950 -140
rect 17970 -160 17975 -140
rect 17905 -170 17975 -160
rect 18005 -90 18035 -80
rect 18005 -110 18010 -90
rect 18030 -110 18035 -90
rect 18005 -140 18035 -110
rect 18005 -160 18010 -140
rect 18030 -160 18035 -140
rect 18005 -170 18035 -160
rect 18065 -90 18095 -80
rect 18065 -110 18070 -90
rect 18090 -110 18095 -90
rect 18065 -140 18095 -110
rect 18065 -160 18070 -140
rect 18090 -160 18095 -140
rect 18065 -170 18095 -160
rect 18125 -90 18155 -80
rect 18125 -110 18130 -90
rect 18150 -110 18155 -90
rect 18125 -140 18155 -110
rect 18125 -160 18130 -140
rect 18150 -160 18155 -140
rect 18125 -170 18155 -160
rect 18185 -90 18215 -80
rect 18185 -110 18190 -90
rect 18210 -110 18215 -90
rect 18185 -140 18215 -110
rect 18185 -160 18190 -140
rect 18210 -160 18215 -140
rect 18185 -170 18215 -160
rect 18245 -90 18275 -80
rect 18245 -110 18250 -90
rect 18270 -110 18275 -90
rect 18245 -140 18275 -110
rect 18245 -160 18250 -140
rect 18270 -160 18275 -140
rect 18245 -170 18275 -160
rect 18305 -90 18335 -80
rect 18305 -110 18310 -90
rect 18330 -110 18335 -90
rect 18305 -140 18335 -110
rect 18305 -160 18310 -140
rect 18330 -160 18335 -140
rect 18305 -170 18335 -160
rect 18365 -90 18395 -80
rect 18365 -110 18370 -90
rect 18390 -110 18395 -90
rect 18365 -140 18395 -110
rect 18365 -160 18370 -140
rect 18390 -160 18395 -140
rect 18365 -170 18395 -160
rect 18425 -90 18455 -80
rect 18425 -110 18430 -90
rect 18450 -110 18455 -90
rect 18425 -140 18455 -110
rect 18425 -160 18430 -140
rect 18450 -160 18455 -140
rect 18425 -170 18455 -160
rect 18485 -90 18515 -80
rect 18485 -110 18490 -90
rect 18510 -110 18515 -90
rect 18485 -140 18515 -110
rect 18485 -160 18490 -140
rect 18510 -160 18515 -140
rect 18485 -170 18515 -160
rect 18545 -90 18575 -80
rect 18545 -110 18550 -90
rect 18570 -110 18575 -90
rect 18545 -140 18575 -110
rect 18545 -160 18550 -140
rect 18570 -160 18575 -140
rect 18545 -170 18575 -160
rect 18605 -90 18635 -80
rect 18605 -110 18610 -90
rect 18630 -110 18635 -90
rect 18605 -140 18635 -110
rect 18605 -160 18610 -140
rect 18630 -160 18635 -140
rect 18605 -170 18635 -160
rect 18665 -90 18695 -80
rect 18665 -110 18670 -90
rect 18690 -110 18695 -90
rect 18665 -140 18695 -110
rect 18665 -160 18670 -140
rect 18690 -160 18695 -140
rect 18665 -170 18695 -160
rect 18725 -90 18755 -80
rect 18725 -110 18730 -90
rect 18750 -110 18755 -90
rect 18725 -140 18755 -110
rect 18725 -160 18730 -140
rect 18750 -160 18755 -140
rect 18725 -170 18755 -160
rect 18785 -90 18815 -80
rect 18785 -110 18790 -90
rect 18810 -110 18815 -90
rect 18785 -140 18815 -110
rect 18785 -160 18790 -140
rect 18810 -160 18815 -140
rect 18785 -170 18815 -160
rect 18845 -90 18875 -80
rect 18845 -110 18850 -90
rect 18870 -110 18875 -90
rect 18845 -140 18875 -110
rect 18845 -160 18850 -140
rect 18870 -160 18875 -140
rect 18845 -170 18875 -160
rect 18905 -90 18935 -80
rect 18905 -110 18910 -90
rect 18930 -110 18935 -90
rect 18905 -140 18935 -110
rect 18905 -160 18910 -140
rect 18930 -160 18935 -140
rect 18905 -170 18935 -160
rect 18965 -90 18995 -80
rect 18965 -110 18970 -90
rect 18990 -110 18995 -90
rect 18965 -140 18995 -110
rect 18965 -160 18970 -140
rect 18990 -160 18995 -140
rect 18965 -170 18995 -160
rect 19025 -90 19055 -80
rect 19025 -110 19030 -90
rect 19050 -110 19055 -90
rect 19025 -140 19055 -110
rect 19025 -160 19030 -140
rect 19050 -160 19055 -140
rect 19025 -170 19055 -160
rect 19085 -90 19115 -80
rect 19085 -110 19090 -90
rect 19110 -110 19115 -90
rect 19085 -140 19115 -110
rect 19085 -160 19090 -140
rect 19110 -160 19115 -140
rect 19085 -170 19115 -160
rect 19145 -90 19215 -80
rect 19145 -110 19150 -90
rect 19170 -110 19190 -90
rect 19210 -110 19215 -90
rect 19145 -140 19215 -110
rect 19145 -160 19150 -140
rect 19170 -160 19190 -140
rect 19210 -160 19215 -140
rect 19145 -170 19215 -160
rect 16425 -200 16455 -170
rect 16610 -190 16630 -170
rect 16730 -190 16750 -170
rect 16970 -190 16990 -170
rect 17090 -190 17110 -170
rect 17330 -190 17350 -170
rect 17450 -190 17470 -170
rect 16425 -220 16430 -200
rect 16450 -220 16455 -200
rect 16425 -230 16455 -220
rect 16510 -200 16550 -190
rect 16510 -220 16520 -200
rect 16540 -220 16550 -200
rect 16510 -230 16550 -220
rect 16600 -200 16640 -190
rect 16600 -220 16610 -200
rect 16630 -220 16640 -200
rect 16600 -230 16640 -220
rect 16720 -200 16760 -190
rect 16720 -220 16730 -200
rect 16750 -220 16760 -200
rect 16720 -230 16760 -220
rect 16840 -200 16880 -190
rect 16840 -220 16850 -200
rect 16870 -220 16880 -200
rect 16840 -230 16880 -220
rect 16960 -200 17000 -190
rect 16960 -220 16970 -200
rect 16990 -220 17000 -200
rect 16960 -230 17000 -220
rect 17080 -200 17120 -190
rect 17080 -220 17090 -200
rect 17110 -220 17120 -200
rect 17080 -230 17120 -220
rect 17200 -200 17240 -190
rect 17200 -220 17210 -200
rect 17230 -220 17240 -200
rect 17200 -230 17240 -220
rect 17320 -200 17360 -190
rect 17320 -220 17330 -200
rect 17350 -220 17360 -200
rect 17320 -230 17360 -220
rect 17440 -200 17480 -190
rect 17440 -220 17450 -200
rect 17470 -220 17480 -200
rect 17440 -230 17480 -220
rect 17535 -200 17565 -190
rect 17535 -220 17540 -200
rect 17560 -220 17565 -200
rect 17535 -230 17565 -220
rect 17945 -200 17975 -170
rect 18130 -190 18150 -170
rect 18250 -190 18270 -170
rect 18490 -190 18510 -170
rect 18610 -190 18630 -170
rect 18850 -190 18870 -170
rect 18970 -190 18990 -170
rect 19145 -175 19180 -170
rect 17945 -220 17950 -200
rect 17970 -220 17975 -200
rect 17945 -230 17975 -220
rect 18035 -200 18065 -190
rect 18035 -220 18040 -200
rect 18060 -220 18065 -200
rect 18035 -230 18065 -220
rect 18120 -200 18160 -190
rect 18120 -220 18130 -200
rect 18150 -220 18160 -200
rect 18120 -230 18160 -220
rect 18240 -200 18280 -190
rect 18240 -220 18250 -200
rect 18270 -220 18280 -200
rect 18240 -230 18280 -220
rect 18360 -200 18400 -190
rect 18360 -220 18370 -200
rect 18390 -220 18400 -200
rect 18360 -230 18400 -220
rect 18480 -200 18520 -190
rect 18480 -220 18490 -200
rect 18510 -220 18520 -200
rect 18480 -230 18520 -220
rect 18600 -200 18640 -190
rect 18600 -220 18610 -200
rect 18630 -220 18640 -200
rect 18600 -230 18640 -220
rect 18720 -200 18760 -190
rect 18720 -220 18730 -200
rect 18750 -220 18760 -200
rect 18720 -230 18760 -220
rect 18840 -200 18880 -190
rect 18840 -220 18850 -200
rect 18870 -220 18880 -200
rect 18840 -230 18880 -220
rect 18960 -200 19000 -190
rect 18960 -220 18970 -200
rect 18990 -220 19000 -200
rect 18960 -230 19000 -220
rect 19050 -200 19090 -190
rect 19050 -220 19060 -200
rect 19080 -220 19090 -200
rect 19050 -230 19090 -220
rect 19145 -200 19175 -175
rect 19145 -220 19150 -200
rect 19170 -220 19175 -200
rect 19145 -230 19175 -220
rect 16960 -315 16990 -305
rect 16960 -335 16965 -315
rect 16985 -335 16990 -315
rect 16960 -345 16990 -335
rect 17007 -315 17037 -305
rect 17007 -335 17012 -315
rect 17032 -335 17037 -315
rect 17007 -345 17037 -335
rect 17090 -315 17120 -305
rect 17090 -335 17095 -315
rect 17115 -335 17120 -315
rect 17090 -345 17120 -335
rect 18480 -315 18510 -305
rect 18480 -335 18485 -315
rect 18505 -335 18510 -315
rect 18480 -345 18510 -335
rect 18563 -315 18593 -305
rect 18563 -335 18568 -315
rect 18588 -335 18593 -315
rect 18563 -345 18593 -335
rect 18610 -315 18640 -305
rect 18610 -335 18615 -315
rect 18635 -335 18640 -315
rect 18610 -345 18640 -335
rect 16970 -365 16990 -345
rect 17090 -365 17110 -345
rect 18490 -365 18510 -345
rect 18610 -365 18630 -345
rect 16965 -375 16995 -365
rect 16965 -395 16970 -375
rect 16990 -395 16995 -375
rect 16965 -425 16995 -395
rect 16965 -445 16970 -425
rect 16990 -445 16995 -425
rect 16965 -475 16995 -445
rect 16965 -495 16970 -475
rect 16990 -495 16995 -475
rect 16965 -525 16995 -495
rect 16965 -545 16970 -525
rect 16990 -545 16995 -525
rect 16965 -575 16995 -545
rect 16965 -595 16970 -575
rect 16990 -595 16995 -575
rect 16965 -605 16995 -595
rect 17025 -375 17055 -365
rect 17025 -395 17030 -375
rect 17050 -395 17055 -375
rect 17025 -425 17055 -395
rect 17025 -445 17030 -425
rect 17050 -445 17055 -425
rect 17025 -475 17055 -445
rect 17025 -495 17030 -475
rect 17050 -495 17055 -475
rect 17025 -525 17055 -495
rect 17025 -545 17030 -525
rect 17050 -545 17055 -525
rect 17025 -575 17055 -545
rect 17025 -595 17030 -575
rect 17050 -595 17055 -575
rect 17025 -605 17055 -595
rect 17085 -375 17115 -365
rect 17085 -395 17090 -375
rect 17110 -395 17115 -375
rect 17085 -425 17115 -395
rect 17565 -375 17595 -365
rect 17565 -395 17570 -375
rect 17590 -395 17595 -375
rect 17565 -405 17595 -395
rect 18005 -375 18035 -365
rect 18005 -395 18010 -375
rect 18030 -395 18035 -375
rect 18005 -405 18035 -395
rect 18485 -375 18515 -365
rect 18485 -395 18490 -375
rect 18510 -395 18515 -375
rect 17085 -445 17090 -425
rect 17110 -445 17115 -425
rect 17085 -475 17115 -445
rect 17085 -495 17090 -475
rect 17110 -495 17115 -475
rect 17085 -525 17115 -495
rect 17085 -545 17090 -525
rect 17110 -545 17115 -525
rect 17085 -575 17115 -545
rect 17085 -595 17090 -575
rect 17110 -595 17115 -575
rect 17085 -605 17115 -595
rect 18485 -425 18515 -395
rect 18485 -445 18490 -425
rect 18510 -445 18515 -425
rect 18485 -475 18515 -445
rect 18485 -495 18490 -475
rect 18510 -495 18515 -475
rect 18485 -525 18515 -495
rect 18485 -545 18490 -525
rect 18510 -545 18515 -525
rect 18485 -575 18515 -545
rect 18485 -595 18490 -575
rect 18510 -595 18515 -575
rect 18485 -605 18515 -595
rect 18545 -375 18575 -365
rect 18545 -395 18550 -375
rect 18570 -395 18575 -375
rect 18545 -425 18575 -395
rect 18545 -445 18550 -425
rect 18570 -445 18575 -425
rect 18545 -475 18575 -445
rect 18545 -495 18550 -475
rect 18570 -495 18575 -475
rect 18545 -525 18575 -495
rect 18545 -545 18550 -525
rect 18570 -545 18575 -525
rect 18545 -575 18575 -545
rect 18545 -595 18550 -575
rect 18570 -595 18575 -575
rect 18545 -605 18575 -595
rect 18605 -375 18635 -365
rect 18605 -395 18610 -375
rect 18630 -395 18635 -375
rect 18605 -425 18635 -395
rect 18605 -445 18610 -425
rect 18630 -445 18635 -425
rect 18605 -475 18635 -445
rect 18605 -495 18610 -475
rect 18630 -495 18635 -475
rect 18605 -525 18635 -495
rect 18605 -545 18610 -525
rect 18630 -545 18635 -525
rect 18605 -575 18635 -545
rect 18605 -595 18610 -575
rect 18630 -595 18635 -575
rect 18605 -605 18635 -595
rect 18550 -625 18570 -605
rect 17075 -635 17105 -625
rect 17075 -655 17080 -635
rect 17100 -655 17105 -635
rect 17075 -665 17105 -655
rect 18495 -635 18525 -625
rect 18495 -655 18500 -635
rect 18520 -655 18525 -635
rect 18495 -665 18525 -655
rect 18545 -635 18575 -625
rect 18545 -655 18550 -635
rect 18570 -655 18575 -635
rect 18545 -665 18575 -655
rect 16620 -770 16660 -765
rect 16620 -790 16630 -770
rect 16650 -790 16660 -770
rect 16620 -800 16660 -790
rect 16740 -770 16780 -765
rect 16740 -790 16750 -770
rect 16770 -790 16780 -770
rect 16740 -800 16780 -790
rect 16860 -770 16900 -765
rect 16860 -790 16870 -770
rect 16890 -790 16900 -770
rect 16860 -800 16900 -790
rect 16980 -770 17020 -765
rect 16980 -790 16990 -770
rect 17010 -790 17020 -770
rect 16980 -800 17020 -790
rect 17300 -770 17340 -765
rect 17300 -790 17310 -770
rect 17330 -790 17340 -770
rect 17300 -800 17340 -790
rect 17420 -770 17460 -765
rect 17420 -790 17430 -770
rect 17450 -790 17460 -770
rect 17420 -800 17460 -790
rect 17540 -770 17580 -765
rect 17540 -790 17550 -770
rect 17570 -790 17580 -770
rect 18020 -770 18060 -760
rect 17540 -800 17580 -790
rect 17690 -785 17730 -775
rect 17690 -805 17700 -785
rect 17720 -805 17730 -785
rect 17690 -815 17730 -805
rect 17870 -785 17910 -775
rect 17870 -805 17880 -785
rect 17900 -805 17910 -785
rect 18020 -790 18030 -770
rect 18050 -790 18060 -770
rect 18020 -800 18060 -790
rect 18140 -770 18180 -760
rect 18140 -790 18150 -770
rect 18170 -790 18180 -770
rect 18140 -800 18180 -790
rect 18260 -770 18300 -760
rect 18260 -790 18270 -770
rect 18290 -790 18300 -770
rect 18260 -800 18300 -790
rect 18580 -770 18620 -760
rect 18580 -790 18590 -770
rect 18610 -790 18620 -770
rect 18580 -800 18620 -790
rect 18700 -770 18740 -760
rect 18700 -790 18710 -770
rect 18730 -790 18740 -770
rect 18700 -800 18740 -790
rect 18820 -770 18860 -760
rect 18820 -790 18830 -770
rect 18850 -790 18860 -770
rect 18820 -800 18860 -790
rect 18940 -770 18980 -760
rect 18940 -790 18950 -770
rect 18970 -790 18980 -770
rect 18940 -800 18980 -790
rect 19030 -785 19070 -775
rect 17870 -815 17910 -805
rect 19030 -805 19040 -785
rect 19060 -805 19070 -785
rect 19030 -815 19070 -805
rect 16535 -825 16565 -815
rect 16535 -845 16540 -825
rect 16560 -845 16565 -825
rect 16535 -875 16565 -845
rect 16535 -895 16540 -875
rect 16560 -895 16565 -875
rect 16535 -925 16565 -895
rect 16535 -945 16540 -925
rect 16560 -945 16565 -925
rect 16535 -975 16565 -945
rect 16535 -995 16540 -975
rect 16560 -995 16565 -975
rect 16535 -1025 16565 -995
rect 16535 -1045 16540 -1025
rect 16560 -1045 16565 -1025
rect 16535 -1055 16565 -1045
rect 17075 -825 17185 -815
rect 17075 -845 17080 -825
rect 17100 -845 17120 -825
rect 17140 -845 17160 -825
rect 17180 -845 17185 -825
rect 17075 -875 17185 -845
rect 17075 -895 17080 -875
rect 17100 -895 17120 -875
rect 17140 -895 17160 -875
rect 17180 -895 17185 -875
rect 17075 -925 17185 -895
rect 17075 -945 17080 -925
rect 17100 -945 17120 -925
rect 17140 -945 17160 -925
rect 17180 -945 17185 -925
rect 17075 -975 17185 -945
rect 17075 -995 17080 -975
rect 17100 -995 17120 -975
rect 17140 -995 17160 -975
rect 17180 -995 17185 -975
rect 17075 -1025 17185 -995
rect 17075 -1045 17080 -1025
rect 17100 -1045 17120 -1025
rect 17140 -1045 17160 -1025
rect 17180 -1045 17185 -1025
rect 17075 -1055 17185 -1045
rect 17695 -825 17725 -815
rect 17695 -845 17700 -825
rect 17720 -845 17725 -825
rect 17695 -875 17725 -845
rect 17695 -895 17700 -875
rect 17720 -895 17725 -875
rect 17695 -925 17725 -895
rect 17695 -945 17700 -925
rect 17720 -945 17725 -925
rect 17695 -975 17725 -945
rect 17695 -995 17700 -975
rect 17720 -995 17725 -975
rect 17695 -1025 17725 -995
rect 17695 -1045 17700 -1025
rect 17720 -1045 17725 -1025
rect 17695 -1055 17725 -1045
rect 17875 -825 17905 -815
rect 17875 -845 17880 -825
rect 17900 -845 17905 -825
rect 17875 -875 17905 -845
rect 17875 -895 17880 -875
rect 17900 -895 17905 -875
rect 17875 -925 17905 -895
rect 17875 -945 17880 -925
rect 17900 -945 17905 -925
rect 17875 -975 17905 -945
rect 17875 -995 17880 -975
rect 17900 -995 17905 -975
rect 17875 -1025 17905 -995
rect 17875 -1045 17880 -1025
rect 17900 -1045 17905 -1025
rect 17875 -1055 17905 -1045
rect 18415 -825 18525 -815
rect 18415 -845 18420 -825
rect 18440 -845 18460 -825
rect 18480 -845 18500 -825
rect 18520 -845 18525 -825
rect 18415 -875 18525 -845
rect 18415 -895 18420 -875
rect 18440 -895 18460 -875
rect 18480 -895 18500 -875
rect 18520 -895 18525 -875
rect 18415 -925 18525 -895
rect 18415 -945 18420 -925
rect 18440 -945 18460 -925
rect 18480 -945 18500 -925
rect 18520 -945 18525 -925
rect 18415 -975 18525 -945
rect 18415 -995 18420 -975
rect 18440 -995 18460 -975
rect 18480 -995 18500 -975
rect 18520 -995 18525 -975
rect 18415 -1025 18525 -995
rect 18415 -1045 18420 -1025
rect 18440 -1045 18460 -1025
rect 18480 -1045 18500 -1025
rect 18520 -1045 18525 -1025
rect 18415 -1055 18525 -1045
rect 19035 -825 19065 -815
rect 19035 -845 19040 -825
rect 19060 -845 19065 -825
rect 19035 -875 19065 -845
rect 19035 -895 19040 -875
rect 19060 -895 19065 -875
rect 19035 -925 19065 -895
rect 19035 -945 19040 -925
rect 19060 -945 19065 -925
rect 19035 -975 19065 -945
rect 19035 -995 19040 -975
rect 19060 -995 19065 -975
rect 19035 -1025 19065 -995
rect 19035 -1045 19040 -1025
rect 19060 -1045 19065 -1025
rect 19035 -1055 19065 -1045
rect 17120 -1075 17140 -1055
rect 18460 -1075 18480 -1055
rect 17110 -1085 17150 -1075
rect 17110 -1105 17120 -1085
rect 17140 -1105 17150 -1085
rect 17110 -1115 17150 -1105
rect 18450 -1085 18490 -1075
rect 18450 -1105 18460 -1085
rect 18480 -1105 18490 -1085
rect 18450 -1115 18490 -1105
rect 16740 -1145 16780 -1135
rect 16740 -1165 16750 -1145
rect 16770 -1165 16780 -1145
rect 16740 -1175 16780 -1165
rect 16820 -1145 16860 -1135
rect 16820 -1165 16830 -1145
rect 16850 -1165 16860 -1145
rect 16820 -1175 16860 -1165
rect 16900 -1145 16940 -1135
rect 16900 -1165 16910 -1145
rect 16930 -1165 16940 -1145
rect 16900 -1175 16940 -1165
rect 16980 -1145 17020 -1135
rect 16980 -1165 16990 -1145
rect 17010 -1165 17020 -1145
rect 16980 -1175 17020 -1165
rect 17060 -1145 17100 -1135
rect 17060 -1165 17070 -1145
rect 17090 -1165 17100 -1145
rect 17060 -1175 17100 -1165
rect 17140 -1145 17180 -1135
rect 17140 -1165 17150 -1145
rect 17170 -1165 17180 -1145
rect 17140 -1175 17180 -1165
rect 17220 -1145 17260 -1135
rect 17220 -1165 17230 -1145
rect 17250 -1165 17260 -1145
rect 17220 -1175 17260 -1165
rect 17300 -1145 17340 -1135
rect 17300 -1165 17310 -1145
rect 17330 -1165 17340 -1145
rect 17300 -1175 17340 -1165
rect 17380 -1145 17420 -1135
rect 17380 -1165 17390 -1145
rect 17410 -1165 17420 -1145
rect 17380 -1175 17420 -1165
rect 17460 -1145 17500 -1135
rect 17460 -1165 17470 -1145
rect 17490 -1165 17500 -1145
rect 17460 -1175 17500 -1165
rect 17540 -1145 17580 -1135
rect 17540 -1165 17550 -1145
rect 17570 -1165 17580 -1145
rect 17540 -1175 17580 -1165
rect 17620 -1145 17660 -1135
rect 17620 -1165 17630 -1145
rect 17650 -1165 17660 -1145
rect 17620 -1175 17660 -1165
rect 17700 -1145 17740 -1135
rect 17700 -1165 17710 -1145
rect 17730 -1165 17740 -1145
rect 17700 -1175 17740 -1165
rect 17780 -1145 17820 -1135
rect 17780 -1165 17790 -1145
rect 17810 -1165 17820 -1145
rect 17780 -1175 17820 -1165
rect 17860 -1145 17900 -1135
rect 17860 -1165 17870 -1145
rect 17890 -1165 17900 -1145
rect 17860 -1175 17900 -1165
rect 17940 -1145 17980 -1135
rect 17940 -1165 17950 -1145
rect 17970 -1165 17980 -1145
rect 17940 -1175 17980 -1165
rect 18020 -1145 18060 -1135
rect 18020 -1165 18030 -1145
rect 18050 -1165 18060 -1145
rect 18020 -1175 18060 -1165
rect 18100 -1145 18140 -1135
rect 18100 -1165 18110 -1145
rect 18130 -1165 18140 -1145
rect 18100 -1175 18140 -1165
rect 18180 -1145 18220 -1135
rect 18180 -1165 18190 -1145
rect 18210 -1165 18220 -1145
rect 18180 -1175 18220 -1165
rect 18260 -1145 18300 -1135
rect 18260 -1165 18270 -1145
rect 18290 -1165 18300 -1145
rect 18260 -1175 18300 -1165
rect 18340 -1145 18380 -1135
rect 18340 -1165 18350 -1145
rect 18370 -1165 18380 -1145
rect 18340 -1175 18380 -1165
rect 18420 -1145 18460 -1135
rect 18420 -1165 18430 -1145
rect 18450 -1165 18460 -1145
rect 18420 -1175 18460 -1165
rect 18500 -1145 18540 -1135
rect 18500 -1165 18510 -1145
rect 18530 -1165 18540 -1145
rect 18500 -1175 18540 -1165
rect 18580 -1145 18620 -1135
rect 18580 -1165 18590 -1145
rect 18610 -1165 18620 -1145
rect 18580 -1175 18620 -1165
rect 18660 -1145 18700 -1135
rect 18660 -1165 18670 -1145
rect 18690 -1165 18700 -1145
rect 18660 -1175 18700 -1165
rect 18740 -1145 18780 -1135
rect 18740 -1165 18750 -1145
rect 18770 -1165 18780 -1145
rect 18740 -1175 18780 -1165
rect 16750 -1195 16770 -1175
rect 17790 -1195 17810 -1175
rect 16745 -1205 16775 -1195
rect 16745 -1220 16750 -1205
rect 16700 -1225 16750 -1220
rect 16770 -1225 16775 -1205
rect 16700 -1230 16775 -1225
rect 16700 -1250 16710 -1230
rect 16730 -1250 16775 -1230
rect 16700 -1255 16775 -1250
rect 16700 -1260 16750 -1255
rect 16745 -1275 16750 -1260
rect 16770 -1275 16775 -1255
rect 16745 -1285 16775 -1275
rect 17785 -1205 17815 -1195
rect 17785 -1225 17790 -1205
rect 17810 -1225 17815 -1205
rect 17785 -1255 17815 -1225
rect 17785 -1275 17790 -1255
rect 17810 -1275 17815 -1255
rect 17785 -1285 17815 -1275
rect 18825 -1205 18895 -1195
rect 18825 -1225 18830 -1205
rect 18850 -1225 18870 -1205
rect 18890 -1220 18895 -1205
rect 18890 -1225 18935 -1220
rect 18825 -1230 18935 -1225
rect 18825 -1250 18905 -1230
rect 18925 -1250 18935 -1230
rect 18825 -1255 18935 -1250
rect 18825 -1275 18830 -1255
rect 18850 -1275 18870 -1255
rect 18890 -1260 18935 -1255
rect 18890 -1275 18895 -1260
rect 18825 -1285 18895 -1275
rect 16540 -1495 16580 -1485
rect 16540 -1515 16550 -1495
rect 16570 -1515 16580 -1495
rect 16540 -1525 16580 -1515
rect 16600 -1495 16630 -1485
rect 16600 -1515 16605 -1495
rect 16625 -1515 16630 -1495
rect 16600 -1525 16630 -1515
rect 16650 -1495 16690 -1485
rect 16650 -1515 16660 -1495
rect 16680 -1515 16690 -1495
rect 16650 -1525 16690 -1515
rect 16710 -1495 16740 -1485
rect 16710 -1515 16715 -1495
rect 16735 -1515 16740 -1495
rect 16710 -1525 16740 -1515
rect 16760 -1495 16800 -1485
rect 16760 -1515 16770 -1495
rect 16790 -1515 16800 -1495
rect 16760 -1525 16800 -1515
rect 16820 -1495 16860 -1485
rect 16820 -1515 16830 -1495
rect 16850 -1515 16860 -1495
rect 16820 -1525 16860 -1515
rect 17025 -1495 17065 -1485
rect 17025 -1515 17035 -1495
rect 17055 -1515 17065 -1495
rect 17025 -1525 17065 -1515
rect 17135 -1495 17175 -1485
rect 17135 -1515 17145 -1495
rect 17165 -1515 17175 -1495
rect 17135 -1525 17175 -1515
rect 17245 -1495 17285 -1485
rect 17245 -1515 17255 -1495
rect 17275 -1515 17285 -1495
rect 17245 -1525 17285 -1515
rect 17305 -1495 17335 -1485
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17305 -1525 17335 -1515
rect 17355 -1495 17395 -1485
rect 17355 -1515 17365 -1495
rect 17385 -1515 17395 -1495
rect 17355 -1525 17395 -1515
rect 17465 -1495 17505 -1485
rect 17465 -1515 17475 -1495
rect 17495 -1515 17505 -1495
rect 17465 -1525 17505 -1515
rect 17615 -1495 17655 -1485
rect 17615 -1515 17625 -1495
rect 17645 -1515 17655 -1495
rect 17615 -1525 17655 -1515
rect 17725 -1495 17765 -1485
rect 17725 -1515 17735 -1495
rect 17755 -1515 17765 -1495
rect 17725 -1525 17765 -1515
rect 17785 -1495 17815 -1485
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17785 -1525 17815 -1515
rect 17835 -1495 17875 -1485
rect 17835 -1515 17845 -1495
rect 17865 -1515 17875 -1495
rect 17835 -1525 17875 -1515
rect 17945 -1495 17985 -1485
rect 17945 -1515 17955 -1495
rect 17975 -1515 17985 -1495
rect 17945 -1525 17985 -1515
rect 18095 -1495 18135 -1485
rect 18095 -1515 18105 -1495
rect 18125 -1515 18135 -1495
rect 18095 -1525 18135 -1515
rect 18205 -1495 18245 -1485
rect 18205 -1515 18215 -1495
rect 18235 -1515 18245 -1495
rect 18205 -1525 18245 -1515
rect 18265 -1495 18295 -1485
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18265 -1525 18295 -1515
rect 18315 -1495 18355 -1485
rect 18315 -1515 18325 -1495
rect 18345 -1515 18355 -1495
rect 18315 -1525 18355 -1515
rect 18425 -1495 18465 -1485
rect 18425 -1515 18435 -1495
rect 18455 -1515 18465 -1495
rect 18425 -1525 18465 -1515
rect 18535 -1495 18575 -1485
rect 18535 -1515 18545 -1495
rect 18565 -1515 18575 -1495
rect 18535 -1525 18575 -1515
rect 16545 -1545 16575 -1525
rect 16605 -1545 16625 -1525
rect 16660 -1545 16680 -1525
rect 16770 -1545 16790 -1525
rect 16820 -1545 16850 -1525
rect 17030 -1545 17060 -1525
rect 17145 -1545 17165 -1525
rect 17255 -1545 17275 -1525
rect 17365 -1545 17385 -1525
rect 17470 -1545 17500 -1525
rect 17620 -1545 17650 -1525
rect 17735 -1545 17755 -1525
rect 17845 -1545 17865 -1525
rect 17950 -1545 17980 -1525
rect 18100 -1545 18130 -1525
rect 18215 -1545 18235 -1525
rect 18325 -1545 18345 -1525
rect 18435 -1545 18455 -1525
rect 18540 -1545 18570 -1525
rect 16505 -1555 16575 -1545
rect 16505 -1575 16510 -1555
rect 16530 -1575 16550 -1555
rect 16570 -1575 16575 -1555
rect 16505 -1605 16575 -1575
rect 16505 -1625 16510 -1605
rect 16530 -1625 16550 -1605
rect 16570 -1625 16575 -1605
rect 16505 -1635 16575 -1625
rect 16600 -1555 16630 -1545
rect 16600 -1575 16605 -1555
rect 16625 -1575 16630 -1555
rect 16600 -1605 16630 -1575
rect 16600 -1625 16605 -1605
rect 16625 -1625 16630 -1605
rect 16600 -1635 16630 -1625
rect 16655 -1555 16685 -1545
rect 16655 -1575 16660 -1555
rect 16680 -1575 16685 -1555
rect 16655 -1605 16685 -1575
rect 16655 -1625 16660 -1605
rect 16680 -1625 16685 -1605
rect 16655 -1635 16685 -1625
rect 16710 -1555 16740 -1545
rect 16710 -1575 16715 -1555
rect 16735 -1575 16740 -1555
rect 16710 -1605 16740 -1575
rect 16710 -1625 16715 -1605
rect 16735 -1625 16740 -1605
rect 16710 -1635 16740 -1625
rect 16765 -1555 16795 -1545
rect 16765 -1575 16770 -1555
rect 16790 -1575 16795 -1555
rect 16765 -1605 16795 -1575
rect 16765 -1625 16770 -1605
rect 16790 -1625 16795 -1605
rect 16765 -1635 16795 -1625
rect 16820 -1555 16890 -1545
rect 16820 -1575 16825 -1555
rect 16845 -1575 16865 -1555
rect 16885 -1575 16890 -1555
rect 16820 -1605 16890 -1575
rect 16820 -1625 16825 -1605
rect 16845 -1625 16865 -1605
rect 16885 -1625 16890 -1605
rect 16820 -1635 16890 -1625
rect 16990 -1555 17060 -1545
rect 16990 -1575 16995 -1555
rect 17015 -1575 17035 -1555
rect 17055 -1575 17060 -1555
rect 16990 -1605 17060 -1575
rect 16990 -1625 16995 -1605
rect 17015 -1625 17035 -1605
rect 17055 -1625 17060 -1605
rect 16990 -1635 17060 -1625
rect 17085 -1555 17115 -1545
rect 17085 -1575 17090 -1555
rect 17110 -1575 17115 -1555
rect 17085 -1605 17115 -1575
rect 17085 -1625 17090 -1605
rect 17110 -1625 17115 -1605
rect 17085 -1635 17115 -1625
rect 17140 -1555 17170 -1545
rect 17140 -1575 17145 -1555
rect 17165 -1575 17170 -1555
rect 17140 -1605 17170 -1575
rect 17140 -1625 17145 -1605
rect 17165 -1625 17170 -1605
rect 17140 -1635 17170 -1625
rect 17195 -1555 17225 -1545
rect 17195 -1575 17200 -1555
rect 17220 -1575 17225 -1555
rect 17195 -1605 17225 -1575
rect 17195 -1625 17200 -1605
rect 17220 -1625 17225 -1605
rect 17195 -1635 17225 -1625
rect 17250 -1555 17280 -1545
rect 17250 -1575 17255 -1555
rect 17275 -1575 17280 -1555
rect 17250 -1605 17280 -1575
rect 17250 -1625 17255 -1605
rect 17275 -1625 17280 -1605
rect 17250 -1635 17280 -1625
rect 17305 -1555 17335 -1545
rect 17305 -1575 17310 -1555
rect 17330 -1575 17335 -1555
rect 17305 -1605 17335 -1575
rect 17305 -1625 17310 -1605
rect 17330 -1625 17335 -1605
rect 17305 -1635 17335 -1625
rect 17360 -1555 17390 -1545
rect 17360 -1575 17365 -1555
rect 17385 -1575 17390 -1555
rect 17360 -1605 17390 -1575
rect 17360 -1625 17365 -1605
rect 17385 -1625 17390 -1605
rect 17360 -1635 17390 -1625
rect 17415 -1555 17445 -1545
rect 17415 -1575 17420 -1555
rect 17440 -1575 17445 -1555
rect 17415 -1605 17445 -1575
rect 17415 -1625 17420 -1605
rect 17440 -1625 17445 -1605
rect 17415 -1635 17445 -1625
rect 17470 -1555 17540 -1545
rect 17470 -1575 17475 -1555
rect 17495 -1575 17515 -1555
rect 17535 -1575 17540 -1555
rect 17470 -1605 17540 -1575
rect 17470 -1625 17475 -1605
rect 17495 -1625 17515 -1605
rect 17535 -1625 17540 -1605
rect 17470 -1635 17540 -1625
rect 17580 -1555 17650 -1545
rect 17580 -1575 17585 -1555
rect 17605 -1575 17625 -1555
rect 17645 -1575 17650 -1555
rect 17580 -1605 17650 -1575
rect 17580 -1625 17585 -1605
rect 17605 -1625 17625 -1605
rect 17645 -1625 17650 -1605
rect 17580 -1635 17650 -1625
rect 17675 -1555 17705 -1545
rect 17675 -1575 17680 -1555
rect 17700 -1575 17705 -1555
rect 17675 -1605 17705 -1575
rect 17675 -1625 17680 -1605
rect 17700 -1625 17705 -1605
rect 17675 -1635 17705 -1625
rect 17730 -1555 17760 -1545
rect 17730 -1575 17735 -1555
rect 17755 -1575 17760 -1555
rect 17730 -1605 17760 -1575
rect 17730 -1625 17735 -1605
rect 17755 -1625 17760 -1605
rect 17730 -1635 17760 -1625
rect 17785 -1555 17815 -1545
rect 17785 -1575 17790 -1555
rect 17810 -1575 17815 -1555
rect 17785 -1605 17815 -1575
rect 17785 -1625 17790 -1605
rect 17810 -1625 17815 -1605
rect 17785 -1635 17815 -1625
rect 17840 -1555 17870 -1545
rect 17840 -1575 17845 -1555
rect 17865 -1575 17870 -1555
rect 17840 -1605 17870 -1575
rect 17840 -1625 17845 -1605
rect 17865 -1625 17870 -1605
rect 17840 -1635 17870 -1625
rect 17895 -1555 17925 -1545
rect 17895 -1575 17900 -1555
rect 17920 -1575 17925 -1555
rect 17895 -1605 17925 -1575
rect 17895 -1625 17900 -1605
rect 17920 -1625 17925 -1605
rect 17895 -1635 17925 -1625
rect 17950 -1555 18020 -1545
rect 17950 -1575 17955 -1555
rect 17975 -1575 17995 -1555
rect 18015 -1575 18020 -1555
rect 17950 -1605 18020 -1575
rect 17950 -1625 17955 -1605
rect 17975 -1625 17995 -1605
rect 18015 -1625 18020 -1605
rect 17950 -1635 18020 -1625
rect 18060 -1555 18130 -1545
rect 18060 -1575 18065 -1555
rect 18085 -1575 18105 -1555
rect 18125 -1575 18130 -1555
rect 18060 -1605 18130 -1575
rect 18060 -1625 18065 -1605
rect 18085 -1625 18105 -1605
rect 18125 -1625 18130 -1605
rect 18060 -1635 18130 -1625
rect 18155 -1555 18185 -1545
rect 18155 -1575 18160 -1555
rect 18180 -1575 18185 -1555
rect 18155 -1605 18185 -1575
rect 18155 -1625 18160 -1605
rect 18180 -1625 18185 -1605
rect 18155 -1635 18185 -1625
rect 18210 -1555 18240 -1545
rect 18210 -1575 18215 -1555
rect 18235 -1575 18240 -1555
rect 18210 -1605 18240 -1575
rect 18210 -1625 18215 -1605
rect 18235 -1625 18240 -1605
rect 18210 -1635 18240 -1625
rect 18265 -1555 18295 -1545
rect 18265 -1575 18270 -1555
rect 18290 -1575 18295 -1555
rect 18265 -1605 18295 -1575
rect 18265 -1625 18270 -1605
rect 18290 -1625 18295 -1605
rect 18265 -1635 18295 -1625
rect 18320 -1555 18350 -1545
rect 18320 -1575 18325 -1555
rect 18345 -1575 18350 -1555
rect 18320 -1605 18350 -1575
rect 18320 -1625 18325 -1605
rect 18345 -1625 18350 -1605
rect 18320 -1635 18350 -1625
rect 18375 -1555 18405 -1545
rect 18375 -1575 18380 -1555
rect 18400 -1575 18405 -1555
rect 18375 -1605 18405 -1575
rect 18375 -1625 18380 -1605
rect 18400 -1625 18405 -1605
rect 18375 -1635 18405 -1625
rect 18430 -1555 18460 -1545
rect 18430 -1575 18435 -1555
rect 18455 -1575 18460 -1555
rect 18430 -1605 18460 -1575
rect 18430 -1625 18435 -1605
rect 18455 -1625 18460 -1605
rect 18430 -1635 18460 -1625
rect 18485 -1555 18515 -1545
rect 18485 -1575 18490 -1555
rect 18510 -1575 18515 -1555
rect 18485 -1605 18515 -1575
rect 18485 -1625 18490 -1605
rect 18510 -1625 18515 -1605
rect 18485 -1635 18515 -1625
rect 18540 -1555 18610 -1545
rect 18540 -1575 18545 -1555
rect 18565 -1575 18585 -1555
rect 18605 -1575 18610 -1555
rect 18540 -1605 18610 -1575
rect 18540 -1625 18545 -1605
rect 18565 -1625 18585 -1605
rect 18605 -1625 18610 -1605
rect 18540 -1635 18610 -1625
rect 16715 -1655 16735 -1635
rect 17090 -1655 17110 -1635
rect 17310 -1655 17330 -1635
rect 17680 -1655 17700 -1635
rect 17790 -1655 17810 -1635
rect 17900 -1655 17920 -1635
rect 18270 -1655 18290 -1635
rect 18490 -1655 18510 -1635
rect 16705 -1665 16745 -1655
rect 16705 -1685 16715 -1665
rect 16735 -1685 16745 -1665
rect 16705 -1695 16745 -1685
rect 17080 -1665 17120 -1655
rect 17080 -1685 17090 -1665
rect 17110 -1685 17120 -1665
rect 17080 -1695 17120 -1685
rect 17190 -1665 17230 -1655
rect 17190 -1685 17200 -1665
rect 17220 -1685 17230 -1665
rect 17190 -1695 17230 -1685
rect 17300 -1665 17340 -1655
rect 17300 -1685 17310 -1665
rect 17330 -1685 17340 -1665
rect 17300 -1695 17340 -1685
rect 17410 -1665 17450 -1655
rect 17410 -1685 17420 -1665
rect 17440 -1685 17450 -1665
rect 17410 -1695 17450 -1685
rect 17670 -1665 17710 -1655
rect 17670 -1685 17680 -1665
rect 17700 -1685 17710 -1665
rect 17670 -1695 17710 -1685
rect 17780 -1665 17820 -1655
rect 17780 -1685 17790 -1665
rect 17810 -1685 17820 -1665
rect 17780 -1695 17820 -1685
rect 17890 -1665 17930 -1655
rect 17890 -1685 17900 -1665
rect 17920 -1685 17930 -1665
rect 17890 -1695 17930 -1685
rect 18150 -1665 18190 -1655
rect 18150 -1685 18160 -1665
rect 18180 -1685 18190 -1665
rect 18150 -1695 18190 -1685
rect 18260 -1665 18300 -1655
rect 18260 -1685 18270 -1665
rect 18290 -1685 18300 -1665
rect 18260 -1695 18300 -1685
rect 18370 -1665 18410 -1655
rect 18370 -1685 18380 -1665
rect 18400 -1685 18410 -1665
rect 18370 -1695 18410 -1685
rect 18480 -1665 18520 -1655
rect 18480 -1685 18490 -1665
rect 18510 -1685 18520 -1665
rect 18480 -1695 18520 -1685
rect 17425 -2005 17470 -2000
rect 17425 -2030 17435 -2005
rect 17460 -2030 17470 -2005
rect 17425 -2035 17470 -2030
rect 18124 -2005 18169 -2000
rect 18124 -2030 18134 -2005
rect 18159 -2030 18169 -2005
rect 18124 -2035 18169 -2030
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16160 -3030 16195 -3020
rect 16160 -3055 16165 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3065 16195 -3055
rect 15950 -3121 15985 -3111
rect 15950 -3146 15955 -3121
rect 15980 -3146 15985 -3121
rect 15950 -3156 15985 -3146
rect 16255 -3100 16280 -3065
rect 16580 -2975 16605 -2940
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19405 -3002 19440 -2992
rect 19405 -3027 19410 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3037 19440 -3027
rect 19320 -3072 19345 -3037
rect 19610 -3121 19645 -3111
rect 19610 -3146 19615 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3156 19645 -3146
rect 16795 -3600 18805 -3475
rect 15950 -3794 15985 -3784
rect 15950 -3819 15955 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3829 15985 -3819
rect 16195 -3889 16220 -3854
rect 16280 -3899 16315 -3889
rect 16280 -3924 16285 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3934 16315 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4170 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19380 -3889 19405 -3854
rect 19610 -3794 19645 -3784
rect 19610 -3819 19615 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3829 19645 -3819
rect 19285 -3899 19320 -3889
rect 19285 -3924 19290 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3934 19320 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4190 17790 -4170
rect 17810 -4190 17820 -4170
rect 17780 -4220 17820 -4190
rect 17780 -4240 17790 -4220
rect 17810 -4240 17820 -4220
rect 17780 -4270 17820 -4240
rect 17780 -4290 17790 -4270
rect 17810 -4290 17820 -4270
rect 17780 -4300 17820 -4290
<< viali >>
rect 16495 1435 16515 1455
rect 17790 1435 17810 1455
rect 16375 1255 16395 1275
rect 16495 1255 16515 1275
rect 16615 1255 16635 1275
rect 16895 1255 16915 1275
rect 16950 1255 16970 1275
rect 17005 1255 17025 1275
rect 17060 1255 17080 1275
rect 17115 1255 17135 1275
rect 17225 1255 17245 1275
rect 17505 1255 17525 1275
rect 17570 1255 17590 1275
rect 17625 1255 17645 1275
rect 17680 1255 17700 1275
rect 17735 1255 17755 1275
rect 17790 1255 17810 1275
rect 17845 1255 17865 1275
rect 17900 1255 17920 1275
rect 17955 1255 17975 1275
rect 18010 1255 18030 1275
rect 18075 1255 18095 1275
rect 18355 1255 18375 1275
rect 18465 1255 18485 1275
rect 18520 1255 18540 1275
rect 18575 1255 18595 1275
rect 18630 1255 18650 1275
rect 18685 1255 18705 1275
rect 16440 1085 16460 1105
rect 16550 1085 16570 1105
rect 16950 1085 16970 1105
rect 17060 1085 17080 1105
rect 17170 1085 17190 1105
rect 17625 1085 17645 1105
rect 17735 1085 17755 1105
rect 17845 1085 17865 1105
rect 17955 1085 17975 1105
rect 18410 1085 18430 1105
rect 18520 1085 18540 1105
rect 18630 1085 18650 1105
rect 16980 790 17000 810
rect 17160 790 17180 810
rect 17340 790 17360 810
rect 17520 790 17540 810
rect 17700 790 17720 810
rect 17880 790 17900 810
rect 18060 790 18080 810
rect 18240 790 18260 810
rect 18420 790 18440 810
rect 18600 790 18620 810
rect 18915 790 18935 810
rect 19025 790 19045 810
rect 19085 790 19105 810
rect 16445 690 16465 710
rect 16555 690 16575 710
rect 16665 690 16685 710
rect 16490 520 16510 540
rect 16555 520 16575 540
rect 16620 520 16640 540
rect 18960 520 18980 540
rect 19010 470 19030 490
rect 17070 420 17090 440
rect 17250 420 17270 440
rect 17430 420 17450 440
rect 17610 420 17630 440
rect 17700 420 17720 440
rect 17790 420 17810 440
rect 17970 420 17990 440
rect 18150 420 18170 440
rect 18330 420 18350 440
rect 18420 420 18440 440
rect 18510 420 18530 440
rect 16430 -50 16450 -30
rect 16490 -50 16510 -30
rect 16550 -50 16570 -30
rect 16670 -50 16690 -30
rect 16790 -50 16810 -30
rect 16850 -50 16870 -30
rect 16910 -50 16930 -30
rect 17030 -50 17050 -30
rect 17150 -50 17170 -30
rect 17210 -50 17230 -30
rect 17270 -50 17290 -30
rect 17390 -50 17410 -30
rect 17510 -50 17530 -30
rect 17570 -50 17590 -30
rect 17630 -50 17650 -30
rect 17950 -50 17970 -30
rect 18010 -50 18030 -30
rect 18070 -50 18090 -30
rect 18190 -50 18210 -30
rect 18310 -50 18330 -30
rect 18370 -50 18390 -30
rect 18430 -50 18450 -30
rect 18550 -50 18570 -30
rect 18670 -50 18690 -30
rect 18730 -50 18750 -30
rect 18790 -50 18810 -30
rect 18910 -50 18930 -30
rect 19030 -50 19050 -30
rect 19090 -50 19110 -30
rect 19150 -50 19170 -30
rect 16520 -220 16540 -200
rect 16610 -220 16630 -200
rect 16730 -220 16750 -200
rect 16850 -220 16870 -200
rect 16970 -220 16990 -200
rect 17090 -220 17110 -200
rect 17210 -220 17230 -200
rect 17330 -220 17350 -200
rect 17450 -220 17470 -200
rect 17540 -220 17560 -200
rect 18040 -220 18060 -200
rect 18130 -220 18150 -200
rect 18250 -220 18270 -200
rect 18370 -220 18390 -200
rect 18490 -220 18510 -200
rect 18610 -220 18630 -200
rect 18730 -220 18750 -200
rect 18850 -220 18870 -200
rect 18970 -220 18990 -200
rect 19060 -220 19080 -200
rect 16965 -335 16985 -315
rect 17012 -335 17032 -315
rect 17095 -335 17115 -315
rect 18485 -335 18505 -315
rect 18568 -335 18588 -315
rect 18615 -335 18635 -315
rect 17030 -395 17050 -375
rect 17030 -445 17050 -425
rect 17030 -495 17050 -475
rect 17030 -545 17050 -525
rect 17030 -595 17050 -575
rect 17570 -395 17590 -375
rect 18010 -395 18030 -375
rect 17080 -655 17100 -635
rect 18500 -655 18520 -635
rect 18550 -655 18570 -635
rect 16630 -790 16650 -770
rect 16750 -790 16770 -770
rect 16870 -790 16890 -770
rect 16990 -790 17010 -770
rect 17310 -790 17330 -770
rect 17430 -790 17450 -770
rect 17550 -790 17570 -770
rect 17700 -805 17720 -785
rect 17880 -805 17900 -785
rect 18030 -790 18050 -770
rect 18150 -790 18170 -770
rect 18270 -790 18290 -770
rect 18590 -790 18610 -770
rect 18710 -790 18730 -770
rect 18830 -790 18850 -770
rect 18950 -790 18970 -770
rect 19040 -805 19060 -785
rect 16540 -845 16560 -825
rect 16540 -895 16560 -875
rect 16540 -945 16560 -925
rect 16540 -995 16560 -975
rect 16540 -1045 16560 -1025
rect 17120 -1105 17140 -1085
rect 18460 -1105 18480 -1085
rect 16750 -1165 16770 -1145
rect 16830 -1165 16850 -1145
rect 16910 -1165 16930 -1145
rect 16990 -1165 17010 -1145
rect 17070 -1165 17090 -1145
rect 17150 -1165 17170 -1145
rect 17230 -1165 17250 -1145
rect 17310 -1165 17330 -1145
rect 17390 -1165 17410 -1145
rect 17470 -1165 17490 -1145
rect 17550 -1165 17570 -1145
rect 17630 -1165 17650 -1145
rect 17710 -1165 17730 -1145
rect 17790 -1165 17810 -1145
rect 17870 -1165 17890 -1145
rect 17950 -1165 17970 -1145
rect 18030 -1165 18050 -1145
rect 18110 -1165 18130 -1145
rect 18190 -1165 18210 -1145
rect 18270 -1165 18290 -1145
rect 18350 -1165 18370 -1145
rect 18430 -1165 18450 -1145
rect 18510 -1165 18530 -1145
rect 18590 -1165 18610 -1145
rect 18670 -1165 18690 -1145
rect 18750 -1165 18770 -1145
rect 16710 -1250 16730 -1230
rect 18905 -1250 18925 -1230
rect 16550 -1515 16570 -1495
rect 16605 -1515 16625 -1495
rect 16660 -1515 16680 -1495
rect 16715 -1515 16735 -1495
rect 16770 -1515 16790 -1495
rect 16830 -1515 16850 -1495
rect 17035 -1515 17055 -1495
rect 17145 -1515 17165 -1495
rect 17255 -1515 17275 -1495
rect 17310 -1515 17330 -1495
rect 17365 -1515 17385 -1495
rect 17475 -1515 17495 -1495
rect 17625 -1515 17645 -1495
rect 17735 -1515 17755 -1495
rect 17790 -1515 17810 -1495
rect 17845 -1515 17865 -1495
rect 17955 -1515 17975 -1495
rect 18105 -1515 18125 -1495
rect 18215 -1515 18235 -1495
rect 18270 -1515 18290 -1495
rect 18325 -1515 18345 -1495
rect 18435 -1515 18455 -1495
rect 18545 -1515 18565 -1495
rect 17200 -1575 17220 -1555
rect 17200 -1625 17220 -1605
rect 17420 -1575 17440 -1555
rect 17420 -1625 17440 -1605
rect 18160 -1575 18180 -1555
rect 18160 -1625 18180 -1605
rect 18380 -1575 18400 -1555
rect 18380 -1625 18400 -1605
rect 16715 -1685 16735 -1665
rect 17090 -1685 17110 -1665
rect 17200 -1685 17220 -1665
rect 17310 -1685 17330 -1665
rect 17420 -1685 17440 -1665
rect 17680 -1685 17700 -1665
rect 17790 -1685 17810 -1665
rect 17900 -1685 17920 -1665
rect 18160 -1685 18180 -1665
rect 18270 -1685 18290 -1665
rect 18380 -1685 18400 -1665
rect 18490 -1685 18510 -1665
rect 17435 -2030 17460 -2005
rect 18134 -2030 18159 -2005
rect 16490 -2930 16515 -2905
rect 16165 -3055 16190 -3030
rect 15955 -3146 15980 -3121
rect 19085 -2930 19110 -2905
rect 19410 -3027 19435 -3002
rect 19615 -3146 19640 -3121
rect 15955 -3819 15980 -3794
rect 16285 -3924 16310 -3899
rect 16610 -3999 16635 -3974
rect 19615 -3819 19640 -3794
rect 19290 -3924 19315 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4290 17810 -4270
<< metal1 >>
rect 15725 -255 15765 -250
rect 15725 -285 15730 -255
rect 15760 -285 15765 -255
rect 15725 -290 15765 -285
rect 15735 -4310 15755 -290
rect 15785 -1770 15825 1595
rect 15950 -25 15990 -20
rect 15950 -55 15955 -25
rect 15985 -55 15990 -25
rect 15950 -60 15990 -55
rect 15785 -1800 15790 -1770
rect 15820 -1800 15825 -1770
rect 15785 -1810 15825 -1800
rect 15785 -1840 15790 -1810
rect 15820 -1840 15825 -1810
rect 15785 -1845 15825 -1840
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 -60
rect 16040 -1710 16060 1595
rect 16030 -1715 16070 -1710
rect 16030 -1745 16035 -1715
rect 16065 -1745 16070 -1715
rect 16030 -1750 16070 -1745
rect 16115 -1895 16135 1595
rect 16950 1510 16970 1595
rect 16940 1505 16980 1510
rect 16940 1475 16945 1505
rect 16975 1475 16980 1505
rect 16940 1470 16980 1475
rect 16485 1460 16525 1465
rect 16485 1430 16490 1460
rect 16520 1430 16525 1460
rect 16485 1425 16525 1430
rect 16365 1360 16405 1365
rect 16365 1330 16370 1360
rect 16400 1330 16405 1360
rect 16365 1320 16405 1330
rect 16365 1290 16370 1320
rect 16400 1290 16405 1320
rect 16365 1280 16405 1290
rect 16365 1250 16370 1280
rect 16400 1250 16405 1280
rect 16365 1245 16405 1250
rect 16485 1360 16525 1365
rect 16485 1330 16490 1360
rect 16520 1330 16525 1360
rect 16485 1320 16525 1330
rect 16485 1290 16490 1320
rect 16520 1290 16525 1320
rect 16485 1280 16525 1290
rect 16485 1250 16490 1280
rect 16520 1250 16525 1280
rect 16485 1245 16525 1250
rect 16605 1360 16645 1365
rect 16605 1330 16610 1360
rect 16640 1330 16645 1360
rect 16605 1320 16645 1330
rect 16605 1290 16610 1320
rect 16640 1290 16645 1320
rect 16605 1280 16645 1290
rect 16605 1250 16610 1280
rect 16640 1250 16645 1280
rect 16605 1245 16645 1250
rect 16885 1360 16925 1365
rect 16885 1330 16890 1360
rect 16920 1330 16925 1360
rect 16885 1320 16925 1330
rect 16885 1290 16890 1320
rect 16920 1290 16925 1320
rect 16885 1280 16925 1290
rect 16950 1285 16970 1470
rect 17050 1460 17090 1465
rect 17050 1430 17055 1460
rect 17085 1430 17090 1460
rect 17050 1425 17090 1430
rect 16995 1360 17035 1365
rect 16995 1330 17000 1360
rect 17030 1330 17035 1360
rect 16995 1320 17035 1330
rect 16995 1290 17000 1320
rect 17030 1290 17035 1320
rect 16885 1250 16890 1280
rect 16920 1250 16925 1280
rect 16885 1245 16925 1250
rect 16945 1275 16975 1285
rect 16945 1255 16950 1275
rect 16970 1255 16975 1275
rect 16945 1245 16975 1255
rect 16995 1280 17035 1290
rect 17060 1285 17080 1425
rect 17105 1360 17145 1365
rect 17105 1330 17110 1360
rect 17140 1330 17145 1360
rect 17105 1320 17145 1330
rect 17105 1290 17110 1320
rect 17140 1290 17145 1320
rect 16995 1250 17000 1280
rect 17030 1250 17035 1280
rect 16995 1245 17035 1250
rect 17055 1275 17085 1285
rect 17055 1255 17060 1275
rect 17080 1255 17085 1275
rect 17055 1245 17085 1255
rect 17105 1280 17145 1290
rect 17105 1250 17110 1280
rect 17140 1250 17145 1280
rect 17105 1245 17145 1250
rect 17215 1360 17255 1365
rect 17215 1330 17220 1360
rect 17250 1330 17255 1360
rect 17215 1320 17255 1330
rect 17215 1290 17220 1320
rect 17250 1290 17255 1320
rect 17215 1280 17255 1290
rect 17215 1250 17220 1280
rect 17250 1250 17255 1280
rect 17215 1245 17255 1250
rect 17495 1360 17535 1365
rect 17495 1330 17500 1360
rect 17530 1330 17535 1360
rect 17495 1320 17535 1330
rect 17495 1290 17500 1320
rect 17530 1290 17535 1320
rect 17495 1280 17535 1290
rect 17495 1250 17500 1280
rect 17530 1250 17535 1280
rect 17495 1245 17535 1250
rect 17560 1360 17600 1365
rect 17560 1330 17565 1360
rect 17595 1330 17600 1360
rect 17560 1320 17600 1330
rect 17560 1290 17565 1320
rect 17595 1290 17600 1320
rect 17560 1280 17600 1290
rect 17560 1250 17565 1280
rect 17595 1250 17600 1280
rect 17560 1245 17600 1250
rect 17620 1275 17650 1595
rect 17620 1255 17625 1275
rect 17645 1255 17650 1275
rect 17620 1245 17650 1255
rect 17670 1360 17710 1365
rect 17670 1330 17675 1360
rect 17705 1330 17710 1360
rect 17670 1320 17710 1330
rect 17670 1290 17675 1320
rect 17705 1290 17710 1320
rect 17670 1280 17710 1290
rect 17670 1250 17675 1280
rect 17705 1250 17710 1280
rect 17670 1245 17710 1250
rect 17730 1275 17760 1595
rect 17780 1460 17820 1465
rect 17780 1430 17785 1460
rect 17815 1430 17820 1460
rect 17780 1425 17820 1430
rect 17730 1255 17735 1275
rect 17755 1255 17760 1275
rect 17730 1245 17760 1255
rect 17780 1360 17820 1365
rect 17780 1330 17785 1360
rect 17815 1330 17820 1360
rect 17780 1320 17820 1330
rect 17780 1290 17785 1320
rect 17815 1290 17820 1320
rect 17780 1280 17820 1290
rect 17780 1250 17785 1280
rect 17815 1250 17820 1280
rect 17780 1245 17820 1250
rect 17840 1275 17870 1595
rect 17840 1255 17845 1275
rect 17865 1255 17870 1275
rect 17840 1245 17870 1255
rect 17890 1360 17930 1365
rect 17890 1330 17895 1360
rect 17925 1330 17930 1360
rect 17890 1320 17930 1330
rect 17890 1290 17895 1320
rect 17925 1290 17930 1320
rect 17890 1280 17930 1290
rect 17890 1250 17895 1280
rect 17925 1250 17930 1280
rect 17890 1245 17930 1250
rect 17950 1275 17980 1595
rect 18630 1510 18650 1595
rect 18620 1505 18660 1510
rect 18620 1475 18625 1505
rect 18655 1475 18660 1505
rect 18620 1470 18660 1475
rect 18200 1460 18240 1465
rect 18200 1430 18205 1460
rect 18235 1430 18240 1460
rect 18200 1425 18240 1430
rect 18510 1460 18550 1465
rect 18510 1430 18515 1460
rect 18545 1430 18550 1460
rect 18510 1425 18550 1430
rect 17950 1255 17955 1275
rect 17975 1255 17980 1275
rect 17950 1245 17980 1255
rect 18000 1360 18040 1365
rect 18000 1330 18005 1360
rect 18035 1330 18040 1360
rect 18000 1320 18040 1330
rect 18000 1290 18005 1320
rect 18035 1290 18040 1320
rect 18000 1280 18040 1290
rect 18000 1250 18005 1280
rect 18035 1250 18040 1280
rect 18000 1245 18040 1250
rect 18065 1360 18105 1365
rect 18065 1330 18070 1360
rect 18100 1330 18105 1360
rect 18065 1320 18105 1330
rect 18065 1290 18070 1320
rect 18100 1290 18105 1320
rect 18065 1280 18105 1290
rect 18065 1250 18070 1280
rect 18100 1250 18105 1280
rect 18065 1245 18105 1250
rect 16430 1110 16470 1115
rect 16430 1080 16435 1110
rect 16465 1080 16470 1110
rect 16430 1075 16470 1080
rect 16540 1110 16580 1115
rect 16540 1080 16545 1110
rect 16575 1080 16580 1110
rect 16540 1075 16580 1080
rect 16940 1110 16980 1115
rect 16940 1080 16945 1110
rect 16975 1080 16980 1110
rect 16940 1075 16980 1080
rect 17050 1110 17090 1115
rect 17050 1080 17055 1110
rect 17085 1080 17090 1110
rect 17050 1075 17090 1080
rect 17160 1110 17200 1115
rect 17160 1080 17165 1110
rect 17195 1080 17200 1110
rect 17160 1075 17200 1080
rect 17615 1110 17655 1115
rect 17615 1080 17620 1110
rect 17650 1080 17655 1110
rect 17615 1075 17655 1080
rect 17725 1110 17765 1115
rect 17725 1080 17730 1110
rect 17760 1080 17765 1110
rect 17725 1075 17765 1080
rect 17835 1110 17875 1115
rect 17835 1080 17840 1110
rect 17870 1080 17875 1110
rect 17835 1075 17875 1080
rect 17945 1110 17985 1115
rect 17945 1080 17950 1110
rect 17980 1080 17985 1110
rect 17945 1075 17985 1080
rect 16440 1015 16460 1075
rect 16550 1015 16570 1075
rect 18210 1060 18230 1425
rect 18345 1360 18385 1365
rect 18345 1330 18350 1360
rect 18380 1330 18385 1360
rect 18345 1320 18385 1330
rect 18345 1290 18350 1320
rect 18380 1290 18385 1320
rect 18345 1280 18385 1290
rect 18345 1250 18350 1280
rect 18380 1250 18385 1280
rect 18345 1245 18385 1250
rect 18455 1360 18495 1365
rect 18455 1330 18460 1360
rect 18490 1330 18495 1360
rect 18455 1320 18495 1330
rect 18455 1290 18460 1320
rect 18490 1290 18495 1320
rect 18455 1280 18495 1290
rect 18520 1285 18540 1425
rect 18565 1360 18605 1365
rect 18565 1330 18570 1360
rect 18600 1330 18605 1360
rect 18565 1320 18605 1330
rect 18565 1290 18570 1320
rect 18600 1290 18605 1320
rect 18455 1250 18460 1280
rect 18490 1250 18495 1280
rect 18455 1245 18495 1250
rect 18515 1275 18545 1285
rect 18515 1255 18520 1275
rect 18540 1255 18545 1275
rect 18515 1245 18545 1255
rect 18565 1280 18605 1290
rect 18630 1285 18650 1470
rect 18675 1360 18715 1365
rect 18675 1330 18680 1360
rect 18710 1330 18715 1360
rect 18675 1320 18715 1330
rect 18675 1290 18680 1320
rect 18710 1290 18715 1320
rect 18565 1250 18570 1280
rect 18600 1250 18605 1280
rect 18565 1245 18605 1250
rect 18625 1275 18655 1285
rect 18625 1255 18630 1275
rect 18650 1255 18655 1275
rect 18625 1245 18655 1255
rect 18675 1280 18715 1290
rect 18675 1250 18680 1280
rect 18710 1250 18715 1280
rect 18675 1245 18715 1250
rect 18400 1110 18440 1115
rect 18400 1080 18405 1110
rect 18435 1080 18440 1110
rect 18400 1075 18440 1080
rect 18510 1110 18550 1115
rect 18510 1080 18515 1110
rect 18545 1080 18550 1110
rect 18510 1075 18550 1080
rect 18620 1110 18660 1115
rect 18620 1080 18625 1110
rect 18655 1080 18660 1110
rect 18620 1075 18660 1080
rect 18200 1055 18240 1060
rect 18200 1025 18205 1055
rect 18235 1025 18240 1055
rect 18200 1020 18240 1025
rect 18720 1055 18760 1060
rect 18720 1025 18725 1055
rect 18755 1025 18760 1055
rect 18720 1020 18760 1025
rect 16160 1010 16200 1015
rect 16160 980 16165 1010
rect 16195 980 16200 1010
rect 16160 975 16200 980
rect 16430 1010 16470 1015
rect 16430 980 16435 1010
rect 16465 980 16470 1010
rect 16430 975 16470 980
rect 16540 1010 16580 1015
rect 16540 980 16545 1010
rect 16575 980 16580 1010
rect 16540 975 16580 980
rect 16170 -1320 16190 975
rect 16435 935 16475 940
rect 16435 905 16440 935
rect 16470 905 16475 935
rect 16435 895 16475 905
rect 16435 865 16440 895
rect 16470 865 16475 895
rect 16435 855 16475 865
rect 16435 825 16440 855
rect 16470 825 16475 855
rect 16435 815 16475 825
rect 16435 785 16440 815
rect 16470 785 16475 815
rect 16435 780 16475 785
rect 16655 935 16695 940
rect 16655 905 16660 935
rect 16690 905 16695 935
rect 16655 895 16695 905
rect 16655 865 16660 895
rect 16690 865 16695 895
rect 16655 855 16695 865
rect 16655 825 16660 855
rect 16690 825 16695 855
rect 16655 815 16695 825
rect 16655 785 16660 815
rect 16690 785 16695 815
rect 16655 780 16695 785
rect 16970 935 17010 940
rect 16970 905 16975 935
rect 17005 905 17010 935
rect 16970 895 17010 905
rect 16970 865 16975 895
rect 17005 865 17010 895
rect 16970 855 17010 865
rect 16970 825 16975 855
rect 17005 825 17010 855
rect 16970 815 17010 825
rect 16970 785 16975 815
rect 17005 785 17010 815
rect 16970 780 17010 785
rect 17150 935 17190 940
rect 17150 905 17155 935
rect 17185 905 17190 935
rect 17150 895 17190 905
rect 17150 865 17155 895
rect 17185 865 17190 895
rect 17150 855 17190 865
rect 17150 825 17155 855
rect 17185 825 17190 855
rect 17150 815 17190 825
rect 17150 785 17155 815
rect 17185 785 17190 815
rect 17150 780 17190 785
rect 17330 935 17370 940
rect 17330 905 17335 935
rect 17365 905 17370 935
rect 17330 895 17370 905
rect 17330 865 17335 895
rect 17365 865 17370 895
rect 17330 855 17370 865
rect 17330 825 17335 855
rect 17365 825 17370 855
rect 17330 815 17370 825
rect 17330 785 17335 815
rect 17365 785 17370 815
rect 17330 780 17370 785
rect 17510 935 17550 940
rect 17510 905 17515 935
rect 17545 905 17550 935
rect 17510 895 17550 905
rect 17510 865 17515 895
rect 17545 865 17550 895
rect 17510 855 17550 865
rect 17510 825 17515 855
rect 17545 825 17550 855
rect 17510 815 17550 825
rect 17510 785 17515 815
rect 17545 785 17550 815
rect 17510 780 17550 785
rect 17690 935 17730 940
rect 17690 905 17695 935
rect 17725 905 17730 935
rect 17690 895 17730 905
rect 17690 865 17695 895
rect 17725 865 17730 895
rect 17690 855 17730 865
rect 17690 825 17695 855
rect 17725 825 17730 855
rect 17690 815 17730 825
rect 17690 785 17695 815
rect 17725 785 17730 815
rect 17690 780 17730 785
rect 17870 935 17910 940
rect 17870 905 17875 935
rect 17905 905 17910 935
rect 17870 895 17910 905
rect 17870 865 17875 895
rect 17905 865 17910 895
rect 17870 855 17910 865
rect 17870 825 17875 855
rect 17905 825 17910 855
rect 17870 815 17910 825
rect 17870 785 17875 815
rect 17905 785 17910 815
rect 17870 780 17910 785
rect 18050 935 18090 940
rect 18050 905 18055 935
rect 18085 905 18090 935
rect 18050 895 18090 905
rect 18050 865 18055 895
rect 18085 865 18090 895
rect 18050 855 18090 865
rect 18050 825 18055 855
rect 18085 825 18090 855
rect 18050 815 18090 825
rect 18050 785 18055 815
rect 18085 785 18090 815
rect 18050 780 18090 785
rect 18230 935 18270 940
rect 18230 905 18235 935
rect 18265 905 18270 935
rect 18230 895 18270 905
rect 18230 865 18235 895
rect 18265 865 18270 895
rect 18230 855 18270 865
rect 18230 825 18235 855
rect 18265 825 18270 855
rect 18230 815 18270 825
rect 18230 785 18235 815
rect 18265 785 18270 815
rect 18230 780 18270 785
rect 18410 935 18450 940
rect 18410 905 18415 935
rect 18445 905 18450 935
rect 18410 895 18450 905
rect 18410 865 18415 895
rect 18445 865 18450 895
rect 18410 855 18450 865
rect 18410 825 18415 855
rect 18445 825 18450 855
rect 18410 815 18450 825
rect 18410 785 18415 815
rect 18445 785 18450 815
rect 18410 780 18450 785
rect 18590 935 18630 940
rect 18590 905 18595 935
rect 18625 905 18630 935
rect 18590 895 18630 905
rect 18590 865 18595 895
rect 18625 865 18630 895
rect 18590 855 18630 865
rect 18590 825 18595 855
rect 18625 825 18630 855
rect 18590 815 18630 825
rect 18590 785 18595 815
rect 18625 785 18630 815
rect 18590 780 18630 785
rect 16445 720 16465 780
rect 16665 720 16685 780
rect 16435 710 16475 720
rect 16435 690 16445 710
rect 16465 690 16475 710
rect 16435 680 16475 690
rect 16545 715 16585 720
rect 16545 685 16550 715
rect 16580 685 16585 715
rect 16545 680 16585 685
rect 16655 710 16695 720
rect 16655 690 16665 710
rect 16685 690 16695 710
rect 16655 680 16695 690
rect 16780 715 16820 720
rect 16780 685 16785 715
rect 16815 685 16820 715
rect 16780 680 16820 685
rect 16480 545 16520 550
rect 16480 515 16485 545
rect 16515 515 16520 545
rect 16480 510 16520 515
rect 16545 540 16585 550
rect 16545 520 16555 540
rect 16575 520 16585 540
rect 16545 510 16585 520
rect 16610 545 16650 550
rect 16610 515 16615 545
rect 16645 515 16650 545
rect 16610 510 16650 515
rect 16315 445 16355 450
rect 16315 415 16320 445
rect 16350 415 16355 445
rect 16260 390 16300 395
rect 16260 360 16265 390
rect 16295 360 16300 390
rect 16260 355 16300 360
rect 16205 345 16245 350
rect 16205 315 16210 345
rect 16240 315 16245 345
rect 16205 310 16245 315
rect 16215 -1220 16235 310
rect 16270 -305 16290 355
rect 16260 -310 16300 -305
rect 16260 -340 16265 -310
rect 16295 -340 16300 -310
rect 16260 -345 16300 -340
rect 16205 -1225 16245 -1220
rect 16205 -1255 16210 -1225
rect 16240 -1255 16245 -1225
rect 16205 -1260 16245 -1255
rect 16160 -1325 16200 -1320
rect 16160 -1355 16165 -1325
rect 16195 -1355 16200 -1325
rect 16160 -1360 16200 -1355
rect 16105 -1900 16145 -1895
rect 16105 -1930 16110 -1900
rect 16140 -1930 16145 -1900
rect 16105 -1935 16145 -1930
rect 16155 -1950 16195 -1945
rect 16155 -1980 16160 -1950
rect 16190 -1980 16195 -1950
rect 16155 -1985 16195 -1980
rect 16165 -3020 16185 -1985
rect 16270 -1995 16290 -345
rect 16315 -630 16355 415
rect 16555 350 16575 510
rect 16790 395 16810 680
rect 16840 545 16880 550
rect 16840 515 16845 545
rect 16875 515 16880 545
rect 16840 510 16880 515
rect 16780 390 16820 395
rect 16780 360 16785 390
rect 16815 360 16820 390
rect 16780 355 16820 360
rect 16545 345 16585 350
rect 16545 315 16550 345
rect 16580 315 16585 345
rect 16545 310 16585 315
rect 16420 110 16460 115
rect 16420 80 16425 110
rect 16455 80 16460 110
rect 16420 70 16460 80
rect 16420 40 16425 70
rect 16455 40 16460 70
rect 16420 30 16460 40
rect 16420 0 16425 30
rect 16455 0 16460 30
rect 16420 -5 16460 0
rect 16540 110 16580 115
rect 16540 80 16545 110
rect 16575 80 16580 110
rect 16540 70 16580 80
rect 16540 40 16545 70
rect 16575 40 16580 70
rect 16540 30 16580 40
rect 16540 0 16545 30
rect 16575 0 16580 30
rect 16540 -5 16580 0
rect 16660 110 16700 115
rect 16660 80 16665 110
rect 16695 80 16700 110
rect 16660 70 16700 80
rect 16660 40 16665 70
rect 16695 40 16700 70
rect 16660 30 16700 40
rect 16660 0 16665 30
rect 16695 0 16700 30
rect 16660 -5 16700 0
rect 16780 110 16820 115
rect 16780 80 16785 110
rect 16815 80 16820 110
rect 16780 70 16820 80
rect 16780 40 16785 70
rect 16815 40 16820 70
rect 16780 30 16820 40
rect 16780 0 16785 30
rect 16815 0 16820 30
rect 16780 -5 16820 0
rect 16430 -20 16450 -5
rect 16550 -20 16570 -5
rect 16670 -20 16690 -5
rect 16790 -20 16810 -5
rect 16850 -20 16870 510
rect 17060 440 17100 450
rect 17060 420 17070 440
rect 17090 420 17100 440
rect 17060 410 17100 420
rect 17240 440 17280 450
rect 17240 420 17250 440
rect 17270 420 17280 440
rect 17240 410 17280 420
rect 17420 440 17460 450
rect 17420 420 17430 440
rect 17450 420 17460 440
rect 17420 410 17460 420
rect 17600 445 17640 450
rect 17600 415 17605 445
rect 17635 415 17640 445
rect 17600 410 17640 415
rect 17690 440 17730 450
rect 17690 420 17700 440
rect 17720 420 17730 440
rect 17690 410 17730 420
rect 17780 440 17820 450
rect 17780 420 17790 440
rect 17810 420 17820 440
rect 17780 410 17820 420
rect 17960 445 18000 450
rect 17960 415 17965 445
rect 17995 415 18000 445
rect 17960 410 18000 415
rect 18140 440 18180 450
rect 18140 420 18150 440
rect 18170 420 18180 440
rect 18140 410 18180 420
rect 18320 440 18360 450
rect 18320 420 18330 440
rect 18350 420 18360 440
rect 18320 410 18360 420
rect 18410 440 18450 450
rect 18410 420 18420 440
rect 18440 420 18450 440
rect 18410 410 18450 420
rect 18500 440 18540 450
rect 18500 420 18510 440
rect 18530 420 18540 440
rect 18500 410 18540 420
rect 17070 305 17090 410
rect 17250 350 17270 410
rect 17430 395 17450 410
rect 17420 390 17460 395
rect 17420 360 17425 390
rect 17455 360 17460 390
rect 17420 355 17460 360
rect 17240 345 17280 350
rect 17240 315 17245 345
rect 17275 315 17280 345
rect 17240 310 17280 315
rect 17060 300 17100 305
rect 17060 270 17065 300
rect 17095 270 17100 300
rect 17060 265 17100 270
rect 16900 110 16940 115
rect 16900 80 16905 110
rect 16935 80 16940 110
rect 16900 70 16940 80
rect 16900 40 16905 70
rect 16935 40 16940 70
rect 16900 30 16940 40
rect 16900 0 16905 30
rect 16935 0 16940 30
rect 16900 -5 16940 0
rect 17020 110 17060 115
rect 17020 80 17025 110
rect 17055 80 17060 110
rect 17020 70 17060 80
rect 17020 40 17025 70
rect 17055 40 17060 70
rect 17020 30 17060 40
rect 17020 0 17025 30
rect 17055 0 17060 30
rect 17020 -5 17060 0
rect 17140 110 17180 115
rect 17140 80 17145 110
rect 17175 80 17180 110
rect 17140 70 17180 80
rect 17140 40 17145 70
rect 17175 40 17180 70
rect 17140 30 17180 40
rect 17140 0 17145 30
rect 17175 0 17180 30
rect 17140 -5 17180 0
rect 17260 110 17300 115
rect 17260 80 17265 110
rect 17295 80 17300 110
rect 17260 70 17300 80
rect 17260 40 17265 70
rect 17295 40 17300 70
rect 17260 30 17300 40
rect 17260 0 17265 30
rect 17295 0 17300 30
rect 17260 -5 17300 0
rect 17380 110 17420 115
rect 17380 80 17385 110
rect 17415 80 17420 110
rect 17380 70 17420 80
rect 17380 40 17385 70
rect 17415 40 17420 70
rect 17380 30 17420 40
rect 17380 0 17385 30
rect 17415 0 17420 30
rect 17380 -5 17420 0
rect 17500 110 17540 115
rect 17500 80 17505 110
rect 17535 80 17540 110
rect 17500 70 17540 80
rect 17500 40 17505 70
rect 17535 40 17540 70
rect 17500 30 17540 40
rect 17500 0 17505 30
rect 17535 0 17540 30
rect 17500 -5 17540 0
rect 17620 110 17660 115
rect 17620 80 17625 110
rect 17655 80 17660 110
rect 17620 70 17660 80
rect 17620 40 17625 70
rect 17655 40 17660 70
rect 17620 30 17660 40
rect 17620 0 17625 30
rect 17655 0 17660 30
rect 17620 -5 17660 0
rect 16910 -20 16930 -5
rect 17030 -20 17050 -5
rect 17150 -20 17170 -5
rect 17270 -20 17290 -5
rect 17390 -20 17410 -5
rect 17510 -20 17530 -5
rect 17630 -20 17650 -5
rect 17700 -20 17720 410
rect 17790 305 17810 410
rect 18150 395 18170 410
rect 18140 390 18180 395
rect 18140 360 18145 390
rect 18175 360 18180 390
rect 18140 355 18180 360
rect 18330 350 18350 410
rect 18420 405 18440 410
rect 18320 345 18360 350
rect 18320 315 18325 345
rect 18355 315 18360 345
rect 18320 310 18360 315
rect 18510 305 18530 410
rect 17780 300 17820 305
rect 17780 270 17785 300
rect 17815 270 17820 300
rect 17780 265 17820 270
rect 18500 300 18540 305
rect 18500 270 18505 300
rect 18535 270 18540 300
rect 18500 265 18540 270
rect 18730 255 18750 1020
rect 18905 935 18945 940
rect 18905 905 18910 935
rect 18940 905 18945 935
rect 18905 895 18945 905
rect 18905 865 18910 895
rect 18940 865 18945 895
rect 18905 855 18945 865
rect 18905 825 18910 855
rect 18940 825 18945 855
rect 18905 815 18945 825
rect 18905 785 18910 815
rect 18940 785 18945 815
rect 18905 780 18945 785
rect 19015 935 19055 940
rect 19015 905 19020 935
rect 19050 905 19055 935
rect 19015 895 19055 905
rect 19015 865 19020 895
rect 19050 865 19055 895
rect 19015 855 19055 865
rect 19015 825 19020 855
rect 19050 825 19055 855
rect 19015 815 19055 825
rect 19015 785 19020 815
rect 19050 785 19055 815
rect 19015 780 19055 785
rect 19075 935 19115 940
rect 19075 905 19080 935
rect 19110 905 19115 935
rect 19075 895 19115 905
rect 19075 865 19080 895
rect 19110 865 19115 895
rect 19075 855 19115 865
rect 19075 825 19080 855
rect 19110 825 19115 855
rect 19075 815 19115 825
rect 19075 785 19080 815
rect 19110 785 19115 815
rect 19075 780 19115 785
rect 19270 550 19290 1595
rect 19325 1010 19365 1015
rect 19325 980 19330 1010
rect 19360 980 19365 1010
rect 19325 975 19365 980
rect 18950 545 18990 550
rect 18950 515 18955 545
rect 18985 515 18990 545
rect 18950 510 18990 515
rect 19260 545 19300 550
rect 19260 515 19265 545
rect 19295 515 19300 545
rect 19260 510 19300 515
rect 19000 465 19005 495
rect 19035 465 19040 495
rect 19020 255 19040 465
rect 18000 250 18040 255
rect 18000 220 18005 250
rect 18035 220 18040 250
rect 18000 215 18040 220
rect 18720 250 18760 255
rect 18720 220 18725 250
rect 18755 220 18760 250
rect 18720 215 18760 220
rect 19010 250 19050 255
rect 19010 220 19015 250
rect 19045 220 19050 250
rect 19010 215 19050 220
rect 17940 110 17980 115
rect 17940 80 17945 110
rect 17975 80 17980 110
rect 17940 70 17980 80
rect 17940 40 17945 70
rect 17975 40 17980 70
rect 17940 30 17980 40
rect 17940 0 17945 30
rect 17975 0 17980 30
rect 17940 -5 17980 0
rect 17950 -20 17970 -5
rect 18010 -20 18030 215
rect 18060 110 18100 115
rect 18060 80 18065 110
rect 18095 80 18100 110
rect 18060 70 18100 80
rect 18060 40 18065 70
rect 18095 40 18100 70
rect 18060 30 18100 40
rect 18060 0 18065 30
rect 18095 0 18100 30
rect 18060 -5 18100 0
rect 18180 110 18220 115
rect 18180 80 18185 110
rect 18215 80 18220 110
rect 18180 70 18220 80
rect 18180 40 18185 70
rect 18215 40 18220 70
rect 18180 30 18220 40
rect 18180 0 18185 30
rect 18215 0 18220 30
rect 18180 -5 18220 0
rect 18300 110 18340 115
rect 18300 80 18305 110
rect 18335 80 18340 110
rect 18300 70 18340 80
rect 18300 40 18305 70
rect 18335 40 18340 70
rect 18300 30 18340 40
rect 18300 0 18305 30
rect 18335 0 18340 30
rect 18300 -5 18340 0
rect 18420 110 18460 115
rect 18420 80 18425 110
rect 18455 80 18460 110
rect 18420 70 18460 80
rect 18420 40 18425 70
rect 18455 40 18460 70
rect 18420 30 18460 40
rect 18420 0 18425 30
rect 18455 0 18460 30
rect 18420 -5 18460 0
rect 18540 110 18580 115
rect 18540 80 18545 110
rect 18575 80 18580 110
rect 18540 70 18580 80
rect 18540 40 18545 70
rect 18575 40 18580 70
rect 18540 30 18580 40
rect 18540 0 18545 30
rect 18575 0 18580 30
rect 18540 -5 18580 0
rect 18660 110 18700 115
rect 18660 80 18665 110
rect 18695 80 18700 110
rect 18660 70 18700 80
rect 18660 40 18665 70
rect 18695 40 18700 70
rect 18660 30 18700 40
rect 18660 0 18665 30
rect 18695 0 18700 30
rect 18660 -5 18700 0
rect 18780 110 18820 115
rect 18780 80 18785 110
rect 18815 80 18820 110
rect 18780 70 18820 80
rect 18780 40 18785 70
rect 18815 40 18820 70
rect 18780 30 18820 40
rect 18780 0 18785 30
rect 18815 0 18820 30
rect 18780 -5 18820 0
rect 18900 110 18940 115
rect 18900 80 18905 110
rect 18935 80 18940 110
rect 18900 70 18940 80
rect 18900 40 18905 70
rect 18935 40 18940 70
rect 18900 30 18940 40
rect 18900 0 18905 30
rect 18935 0 18940 30
rect 18900 -5 18940 0
rect 19020 110 19060 115
rect 19020 80 19025 110
rect 19055 80 19060 110
rect 19020 70 19060 80
rect 19020 40 19025 70
rect 19055 40 19060 70
rect 19020 30 19060 40
rect 19020 0 19025 30
rect 19055 0 19060 30
rect 19020 -5 19060 0
rect 19140 110 19180 115
rect 19140 80 19145 110
rect 19175 80 19180 110
rect 19140 70 19180 80
rect 19140 40 19145 70
rect 19175 40 19180 70
rect 19140 30 19180 40
rect 19140 0 19145 30
rect 19175 0 19180 30
rect 19140 -5 19180 0
rect 18070 -20 18090 -5
rect 18190 -20 18210 -5
rect 18310 -20 18330 -5
rect 18430 -20 18450 -5
rect 18550 -20 18570 -5
rect 18670 -20 18690 -5
rect 18790 -20 18810 -5
rect 18910 -20 18930 -5
rect 19030 -20 19050 -5
rect 19150 -20 19170 -5
rect 16425 -30 16455 -20
rect 16425 -50 16430 -30
rect 16450 -50 16455 -30
rect 16425 -65 16455 -50
rect 16480 -25 16520 -20
rect 16480 -55 16485 -25
rect 16515 -55 16520 -25
rect 16480 -60 16520 -55
rect 16545 -30 16575 -20
rect 16545 -50 16550 -30
rect 16570 -50 16575 -30
rect 16545 -60 16575 -50
rect 16665 -30 16695 -20
rect 16665 -50 16670 -30
rect 16690 -50 16695 -30
rect 16665 -60 16695 -50
rect 16785 -30 16815 -20
rect 16785 -50 16790 -30
rect 16810 -50 16815 -30
rect 16785 -60 16815 -50
rect 16840 -25 16880 -20
rect 16840 -55 16845 -25
rect 16875 -55 16880 -25
rect 16840 -60 16880 -55
rect 16905 -30 16935 -20
rect 16905 -50 16910 -30
rect 16930 -50 16935 -30
rect 16905 -60 16935 -50
rect 17025 -30 17055 -20
rect 17025 -50 17030 -30
rect 17050 -50 17055 -30
rect 17025 -60 17055 -50
rect 17145 -30 17175 -20
rect 17145 -50 17150 -30
rect 17170 -50 17175 -30
rect 17145 -60 17175 -50
rect 17200 -25 17240 -20
rect 17200 -55 17205 -25
rect 17235 -55 17240 -25
rect 17200 -60 17240 -55
rect 17265 -30 17295 -20
rect 17265 -50 17270 -30
rect 17290 -50 17295 -30
rect 17265 -60 17295 -50
rect 17385 -30 17415 -20
rect 17385 -50 17390 -30
rect 17410 -50 17415 -30
rect 17385 -60 17415 -50
rect 17505 -30 17535 -20
rect 17505 -50 17510 -30
rect 17530 -50 17535 -30
rect 17505 -60 17535 -50
rect 17560 -25 17600 -20
rect 17560 -55 17565 -25
rect 17595 -55 17600 -25
rect 17560 -60 17600 -55
rect 17625 -30 17655 -20
rect 17625 -50 17630 -30
rect 17650 -50 17655 -30
rect 17625 -65 17655 -50
rect 17690 -25 17730 -20
rect 17690 -55 17695 -25
rect 17725 -55 17730 -25
rect 17690 -60 17730 -55
rect 17870 -25 17910 -20
rect 17870 -55 17875 -25
rect 17905 -55 17910 -25
rect 17870 -60 17910 -55
rect 17945 -30 17975 -20
rect 17945 -50 17950 -30
rect 17970 -50 17975 -30
rect 16510 -200 16550 -190
rect 16510 -220 16520 -200
rect 16540 -220 16550 -200
rect 16510 -230 16550 -220
rect 16600 -195 16640 -190
rect 16600 -225 16605 -195
rect 16635 -225 16640 -195
rect 16600 -230 16640 -225
rect 16720 -200 16760 -190
rect 16720 -220 16730 -200
rect 16750 -220 16760 -200
rect 16720 -230 16760 -220
rect 16840 -200 16880 -190
rect 16840 -220 16850 -200
rect 16870 -220 16880 -200
rect 16840 -230 16880 -220
rect 16960 -195 17000 -190
rect 16960 -225 16965 -195
rect 16995 -225 17000 -195
rect 16960 -230 17000 -225
rect 17080 -200 17120 -190
rect 17080 -220 17090 -200
rect 17110 -220 17120 -200
rect 17080 -230 17120 -220
rect 17200 -200 17240 -190
rect 17200 -220 17210 -200
rect 17230 -220 17240 -200
rect 17200 -230 17240 -220
rect 17320 -195 17360 -190
rect 17320 -225 17325 -195
rect 17355 -225 17360 -195
rect 17320 -230 17360 -225
rect 17440 -200 17480 -190
rect 17440 -220 17450 -200
rect 17470 -220 17480 -200
rect 17440 -230 17480 -220
rect 17535 -200 17565 -190
rect 17535 -220 17540 -200
rect 17560 -220 17565 -200
rect 17535 -230 17565 -220
rect 16520 -250 16540 -230
rect 16730 -250 16750 -230
rect 16850 -250 16870 -230
rect 16510 -255 16550 -250
rect 16510 -285 16515 -255
rect 16545 -285 16550 -255
rect 16510 -290 16550 -285
rect 16720 -255 16760 -250
rect 16720 -285 16725 -255
rect 16755 -285 16760 -255
rect 16720 -290 16760 -285
rect 16840 -255 16880 -250
rect 16840 -285 16845 -255
rect 16875 -285 16880 -255
rect 16840 -290 16880 -285
rect 16970 -305 16990 -230
rect 17090 -250 17110 -230
rect 17210 -250 17230 -230
rect 17450 -250 17470 -230
rect 17540 -250 17560 -230
rect 17080 -255 17120 -250
rect 17080 -285 17085 -255
rect 17115 -285 17120 -255
rect 17080 -290 17120 -285
rect 17200 -255 17240 -250
rect 17200 -285 17205 -255
rect 17235 -285 17240 -255
rect 17200 -290 17240 -285
rect 17440 -255 17480 -250
rect 17440 -285 17445 -255
rect 17475 -285 17480 -255
rect 17440 -290 17480 -285
rect 17530 -255 17570 -250
rect 17530 -285 17535 -255
rect 17565 -285 17570 -255
rect 17530 -290 17570 -285
rect 17090 -305 17110 -290
rect 16960 -315 16990 -305
rect 16960 -335 16965 -315
rect 16985 -335 16990 -315
rect 16960 -345 16990 -335
rect 17007 -310 17037 -305
rect 17007 -345 17037 -340
rect 17090 -315 17120 -305
rect 17090 -335 17095 -315
rect 17115 -335 17120 -315
rect 17090 -345 17120 -335
rect 16315 -660 16320 -630
rect 16350 -660 16355 -630
rect 16315 -665 16355 -660
rect 17025 -375 17055 -365
rect 17025 -395 17030 -375
rect 17050 -395 17055 -375
rect 17025 -425 17055 -395
rect 17565 -370 17595 -365
rect 17565 -405 17595 -400
rect 17025 -445 17030 -425
rect 17050 -445 17055 -425
rect 17025 -475 17055 -445
rect 17025 -495 17030 -475
rect 17050 -495 17055 -475
rect 17025 -525 17055 -495
rect 17025 -545 17030 -525
rect 17050 -545 17055 -525
rect 17025 -575 17055 -545
rect 17025 -595 17030 -575
rect 17050 -595 17055 -575
rect 17025 -705 17055 -595
rect 17075 -630 17105 -625
rect 17075 -665 17105 -660
rect 16530 -710 16570 -705
rect 16530 -740 16535 -710
rect 16565 -740 16570 -710
rect 16530 -745 16570 -740
rect 17020 -710 17060 -705
rect 17020 -740 17025 -710
rect 17055 -740 17060 -710
rect 17020 -745 17060 -740
rect 16535 -825 16565 -745
rect 16620 -765 16660 -760
rect 16620 -795 16625 -765
rect 16655 -795 16660 -765
rect 16620 -800 16660 -795
rect 16740 -765 16780 -760
rect 16740 -795 16745 -765
rect 16775 -795 16780 -765
rect 16740 -800 16780 -795
rect 16860 -765 16900 -760
rect 16860 -795 16865 -765
rect 16895 -795 16900 -765
rect 16860 -800 16900 -795
rect 16980 -765 17020 -760
rect 16980 -795 16985 -765
rect 17015 -795 17020 -765
rect 16980 -800 17020 -795
rect 17300 -765 17340 -760
rect 17300 -795 17305 -765
rect 17335 -795 17340 -765
rect 17300 -800 17340 -795
rect 17420 -765 17460 -760
rect 17420 -795 17425 -765
rect 17455 -795 17460 -765
rect 17420 -800 17460 -795
rect 17540 -765 17580 -760
rect 17540 -795 17545 -765
rect 17575 -795 17580 -765
rect 17700 -775 17720 -60
rect 17780 -370 17820 -365
rect 17780 -400 17785 -370
rect 17815 -400 17820 -370
rect 17780 -405 17820 -400
rect 17540 -800 17580 -795
rect 17690 -785 17730 -775
rect 17690 -805 17700 -785
rect 17720 -805 17730 -785
rect 17690 -815 17730 -805
rect 16535 -845 16540 -825
rect 16560 -845 16565 -825
rect 16535 -875 16565 -845
rect 16535 -895 16540 -875
rect 16560 -895 16565 -875
rect 16535 -925 16565 -895
rect 16535 -945 16540 -925
rect 16560 -945 16565 -925
rect 16535 -975 16565 -945
rect 16535 -995 16540 -975
rect 16560 -995 16565 -975
rect 16535 -1025 16565 -995
rect 16535 -1045 16540 -1025
rect 16560 -1045 16565 -1025
rect 16535 -1055 16565 -1045
rect 17790 -1075 17810 -405
rect 17880 -775 17900 -60
rect 17945 -65 17975 -50
rect 18000 -25 18040 -20
rect 18000 -55 18005 -25
rect 18035 -55 18040 -25
rect 18000 -60 18040 -55
rect 18065 -30 18095 -20
rect 18065 -50 18070 -30
rect 18090 -50 18095 -30
rect 18065 -60 18095 -50
rect 18185 -30 18215 -20
rect 18185 -50 18190 -30
rect 18210 -50 18215 -30
rect 18185 -60 18215 -50
rect 18305 -30 18335 -20
rect 18305 -50 18310 -30
rect 18330 -50 18335 -30
rect 18305 -60 18335 -50
rect 18360 -25 18400 -20
rect 18360 -55 18365 -25
rect 18395 -55 18400 -25
rect 18360 -60 18400 -55
rect 18425 -30 18455 -20
rect 18425 -50 18430 -30
rect 18450 -50 18455 -30
rect 18425 -60 18455 -50
rect 18545 -30 18575 -20
rect 18545 -50 18550 -30
rect 18570 -50 18575 -30
rect 18545 -60 18575 -50
rect 18665 -30 18695 -20
rect 18665 -50 18670 -30
rect 18690 -50 18695 -30
rect 18665 -60 18695 -50
rect 18720 -25 18760 -20
rect 18720 -55 18725 -25
rect 18755 -55 18760 -25
rect 18720 -60 18760 -55
rect 18785 -30 18815 -20
rect 18785 -50 18790 -30
rect 18810 -50 18815 -30
rect 18785 -60 18815 -50
rect 18905 -30 18935 -20
rect 18905 -50 18910 -30
rect 18930 -50 18935 -30
rect 18905 -60 18935 -50
rect 19025 -30 19055 -20
rect 19025 -50 19030 -30
rect 19050 -50 19055 -30
rect 19025 -60 19055 -50
rect 19080 -25 19120 -20
rect 19080 -55 19085 -25
rect 19115 -55 19120 -25
rect 19080 -60 19120 -55
rect 19145 -30 19175 -20
rect 19145 -50 19150 -30
rect 19170 -50 19175 -30
rect 19145 -65 19175 -50
rect 18035 -200 18065 -190
rect 18035 -220 18040 -200
rect 18060 -220 18065 -200
rect 18035 -230 18065 -220
rect 18120 -200 18160 -190
rect 18120 -220 18130 -200
rect 18150 -220 18160 -200
rect 18120 -230 18160 -220
rect 18240 -195 18280 -190
rect 18240 -225 18245 -195
rect 18275 -225 18280 -195
rect 18240 -230 18280 -225
rect 18360 -200 18400 -190
rect 18360 -220 18370 -200
rect 18390 -220 18400 -200
rect 18360 -230 18400 -220
rect 18480 -200 18520 -190
rect 18480 -220 18490 -200
rect 18510 -220 18520 -200
rect 18480 -230 18520 -220
rect 18600 -195 18640 -190
rect 18600 -225 18605 -195
rect 18635 -225 18640 -195
rect 18600 -230 18640 -225
rect 18720 -200 18760 -190
rect 18720 -220 18730 -200
rect 18750 -220 18760 -200
rect 18720 -230 18760 -220
rect 18840 -200 18880 -190
rect 18840 -220 18850 -200
rect 18870 -220 18880 -200
rect 18840 -230 18880 -220
rect 18960 -195 19000 -190
rect 18960 -225 18965 -195
rect 18995 -225 19000 -195
rect 18960 -230 19000 -225
rect 19050 -200 19090 -190
rect 19050 -220 19060 -200
rect 19080 -220 19090 -200
rect 19050 -230 19090 -220
rect 18040 -250 18060 -230
rect 18130 -250 18150 -230
rect 18370 -250 18390 -230
rect 18490 -250 18510 -230
rect 18030 -255 18070 -250
rect 18030 -285 18035 -255
rect 18065 -285 18070 -255
rect 18030 -290 18070 -285
rect 18120 -255 18160 -250
rect 18120 -285 18125 -255
rect 18155 -285 18160 -255
rect 18120 -290 18160 -285
rect 18360 -255 18400 -250
rect 18360 -285 18365 -255
rect 18395 -285 18400 -255
rect 18360 -290 18400 -285
rect 18480 -255 18520 -250
rect 18480 -285 18485 -255
rect 18515 -285 18520 -255
rect 18480 -290 18520 -285
rect 18490 -305 18510 -290
rect 18610 -305 18630 -230
rect 18730 -250 18750 -230
rect 18850 -250 18870 -230
rect 19060 -250 19080 -230
rect 18720 -255 18760 -250
rect 18720 -285 18725 -255
rect 18755 -285 18760 -255
rect 18720 -290 18760 -285
rect 18840 -255 18880 -250
rect 18840 -285 18845 -255
rect 18875 -285 18880 -255
rect 18840 -290 18880 -285
rect 19050 -255 19090 -250
rect 19050 -285 19055 -255
rect 19085 -285 19090 -255
rect 19050 -290 19090 -285
rect 18480 -315 18510 -305
rect 18480 -335 18485 -315
rect 18505 -335 18510 -315
rect 18480 -345 18510 -335
rect 18563 -310 18593 -305
rect 18563 -345 18593 -340
rect 18610 -315 18640 -305
rect 18610 -335 18615 -315
rect 18635 -335 18640 -315
rect 18610 -345 18640 -335
rect 18005 -370 18035 -365
rect 18005 -405 18035 -400
rect 19335 -625 19355 975
rect 19415 305 19435 1595
rect 19460 445 19500 450
rect 19460 415 19465 445
rect 19495 415 19500 445
rect 19405 300 19445 305
rect 19405 270 19410 300
rect 19440 270 19445 300
rect 19405 265 19445 270
rect 19415 -305 19435 265
rect 19405 -310 19445 -305
rect 19405 -340 19410 -310
rect 19440 -340 19445 -310
rect 19405 -345 19445 -340
rect 18495 -630 18525 -625
rect 18495 -665 18525 -660
rect 18545 -635 18575 -625
rect 18545 -655 18550 -635
rect 18570 -655 18575 -635
rect 18545 -665 18575 -655
rect 19325 -630 19365 -625
rect 19325 -660 19330 -630
rect 19360 -660 19365 -630
rect 19325 -665 19365 -660
rect 18550 -705 18570 -665
rect 18540 -710 18580 -705
rect 18540 -740 18545 -710
rect 18575 -740 18580 -710
rect 18540 -745 18580 -740
rect 19030 -710 19070 -705
rect 19030 -740 19035 -710
rect 19065 -740 19070 -710
rect 19030 -745 19070 -740
rect 18020 -765 18060 -760
rect 17870 -785 17910 -775
rect 17870 -805 17880 -785
rect 17900 -805 17910 -785
rect 18020 -795 18025 -765
rect 18055 -795 18060 -765
rect 18020 -800 18060 -795
rect 18140 -765 18180 -760
rect 18140 -795 18145 -765
rect 18175 -795 18180 -765
rect 18140 -800 18180 -795
rect 18260 -765 18300 -760
rect 18260 -795 18265 -765
rect 18295 -795 18300 -765
rect 18260 -800 18300 -795
rect 18580 -765 18620 -760
rect 18580 -795 18585 -765
rect 18615 -795 18620 -765
rect 18580 -800 18620 -795
rect 18700 -765 18740 -760
rect 18700 -795 18705 -765
rect 18735 -795 18740 -765
rect 18700 -800 18740 -795
rect 18820 -765 18860 -760
rect 18820 -795 18825 -765
rect 18855 -795 18860 -765
rect 18820 -800 18860 -795
rect 18940 -765 18980 -760
rect 18940 -795 18945 -765
rect 18975 -795 18980 -765
rect 19040 -775 19060 -745
rect 18940 -800 18980 -795
rect 19030 -785 19070 -775
rect 17870 -815 17910 -805
rect 19030 -805 19040 -785
rect 19060 -805 19070 -785
rect 19030 -815 19070 -805
rect 17110 -1080 17150 -1075
rect 17110 -1110 17115 -1080
rect 17145 -1110 17150 -1080
rect 17110 -1115 17150 -1110
rect 17780 -1080 17820 -1075
rect 17780 -1110 17785 -1080
rect 17815 -1110 17820 -1080
rect 17780 -1115 17820 -1110
rect 18450 -1080 18490 -1075
rect 18450 -1110 18455 -1080
rect 18485 -1110 18490 -1080
rect 18450 -1115 18490 -1110
rect 16740 -1140 16780 -1135
rect 16740 -1170 16745 -1140
rect 16775 -1170 16780 -1140
rect 16740 -1175 16780 -1170
rect 16820 -1140 16860 -1135
rect 16820 -1170 16825 -1140
rect 16855 -1170 16860 -1140
rect 16820 -1175 16860 -1170
rect 16900 -1140 16940 -1135
rect 16900 -1170 16905 -1140
rect 16935 -1170 16940 -1140
rect 16900 -1175 16940 -1170
rect 16980 -1140 17020 -1135
rect 16980 -1170 16985 -1140
rect 17015 -1170 17020 -1140
rect 16980 -1175 17020 -1170
rect 17060 -1140 17100 -1135
rect 17060 -1170 17065 -1140
rect 17095 -1170 17100 -1140
rect 17060 -1175 17100 -1170
rect 17140 -1140 17180 -1135
rect 17140 -1170 17145 -1140
rect 17175 -1170 17180 -1140
rect 17140 -1175 17180 -1170
rect 17220 -1140 17260 -1135
rect 17220 -1170 17225 -1140
rect 17255 -1170 17260 -1140
rect 17220 -1175 17260 -1170
rect 17300 -1140 17340 -1135
rect 17300 -1170 17305 -1140
rect 17335 -1170 17340 -1140
rect 17300 -1175 17340 -1170
rect 17380 -1140 17420 -1135
rect 17380 -1170 17385 -1140
rect 17415 -1170 17420 -1140
rect 17380 -1175 17420 -1170
rect 17460 -1140 17500 -1135
rect 17460 -1170 17465 -1140
rect 17495 -1170 17500 -1140
rect 17460 -1175 17500 -1170
rect 17540 -1140 17580 -1135
rect 17540 -1170 17545 -1140
rect 17575 -1170 17580 -1140
rect 17540 -1175 17580 -1170
rect 17620 -1140 17660 -1135
rect 17620 -1170 17625 -1140
rect 17655 -1170 17660 -1140
rect 17620 -1175 17660 -1170
rect 17700 -1140 17740 -1135
rect 17700 -1170 17705 -1140
rect 17735 -1170 17740 -1140
rect 17700 -1175 17740 -1170
rect 17780 -1140 17820 -1135
rect 17780 -1170 17785 -1140
rect 17815 -1170 17820 -1140
rect 17780 -1175 17820 -1170
rect 17860 -1140 17900 -1135
rect 17860 -1170 17865 -1140
rect 17895 -1170 17900 -1140
rect 17860 -1175 17900 -1170
rect 17940 -1140 17980 -1135
rect 17940 -1170 17945 -1140
rect 17975 -1170 17980 -1140
rect 17940 -1175 17980 -1170
rect 18020 -1140 18060 -1135
rect 18020 -1170 18025 -1140
rect 18055 -1170 18060 -1140
rect 18020 -1175 18060 -1170
rect 18100 -1140 18140 -1135
rect 18100 -1170 18105 -1140
rect 18135 -1170 18140 -1140
rect 18100 -1175 18140 -1170
rect 18180 -1140 18220 -1135
rect 18180 -1170 18185 -1140
rect 18215 -1170 18220 -1140
rect 18180 -1175 18220 -1170
rect 18260 -1140 18300 -1135
rect 18260 -1170 18265 -1140
rect 18295 -1170 18300 -1140
rect 18260 -1175 18300 -1170
rect 18340 -1140 18380 -1135
rect 18340 -1170 18345 -1140
rect 18375 -1170 18380 -1140
rect 18340 -1175 18380 -1170
rect 18420 -1140 18460 -1135
rect 18420 -1170 18425 -1140
rect 18455 -1170 18460 -1140
rect 18420 -1175 18460 -1170
rect 18500 -1140 18540 -1135
rect 18500 -1170 18505 -1140
rect 18535 -1170 18540 -1140
rect 18500 -1175 18540 -1170
rect 18580 -1140 18620 -1135
rect 18580 -1170 18585 -1140
rect 18615 -1170 18620 -1140
rect 18580 -1175 18620 -1170
rect 18660 -1140 18700 -1135
rect 18660 -1170 18665 -1140
rect 18695 -1170 18700 -1140
rect 18660 -1175 18700 -1170
rect 18740 -1140 18780 -1135
rect 18740 -1170 18745 -1140
rect 18775 -1170 18780 -1140
rect 18740 -1175 18780 -1170
rect 16700 -1225 16740 -1220
rect 16700 -1255 16705 -1225
rect 16735 -1255 16740 -1225
rect 16700 -1260 16740 -1255
rect 18895 -1225 18935 -1220
rect 18895 -1255 18900 -1225
rect 18930 -1255 18935 -1225
rect 18895 -1260 18935 -1255
rect 16595 -1325 16635 -1320
rect 16595 -1355 16600 -1325
rect 16630 -1355 16635 -1325
rect 16595 -1360 16635 -1355
rect 16705 -1325 16745 -1320
rect 16705 -1355 16710 -1325
rect 16740 -1355 16745 -1325
rect 16705 -1360 16745 -1355
rect 17300 -1325 17340 -1320
rect 17300 -1355 17305 -1325
rect 17335 -1355 17340 -1325
rect 17300 -1360 17340 -1355
rect 17780 -1325 17820 -1320
rect 17780 -1355 17785 -1325
rect 17815 -1355 17820 -1325
rect 17780 -1360 17820 -1355
rect 18260 -1325 18300 -1320
rect 18260 -1355 18265 -1325
rect 18295 -1355 18300 -1325
rect 18260 -1360 18300 -1355
rect 16540 -1410 16580 -1405
rect 16540 -1440 16545 -1410
rect 16575 -1440 16580 -1410
rect 16540 -1450 16580 -1440
rect 16540 -1480 16545 -1450
rect 16575 -1480 16580 -1450
rect 16540 -1490 16580 -1480
rect 16605 -1485 16625 -1360
rect 16650 -1410 16690 -1405
rect 16650 -1440 16655 -1410
rect 16685 -1440 16690 -1410
rect 16650 -1450 16690 -1440
rect 16650 -1480 16655 -1450
rect 16685 -1480 16690 -1450
rect 16540 -1520 16545 -1490
rect 16575 -1520 16580 -1490
rect 16540 -1525 16580 -1520
rect 16600 -1495 16630 -1485
rect 16600 -1515 16605 -1495
rect 16625 -1515 16630 -1495
rect 16600 -1525 16630 -1515
rect 16650 -1490 16690 -1480
rect 16715 -1485 16735 -1360
rect 16760 -1410 16800 -1405
rect 16760 -1440 16765 -1410
rect 16795 -1440 16800 -1410
rect 16760 -1450 16800 -1440
rect 16760 -1480 16765 -1450
rect 16795 -1480 16800 -1450
rect 16650 -1520 16655 -1490
rect 16685 -1520 16690 -1490
rect 16650 -1525 16690 -1520
rect 16710 -1495 16740 -1485
rect 16710 -1515 16715 -1495
rect 16735 -1515 16740 -1495
rect 16710 -1525 16740 -1515
rect 16760 -1490 16800 -1480
rect 16760 -1520 16765 -1490
rect 16795 -1520 16800 -1490
rect 16760 -1525 16800 -1520
rect 16820 -1410 16860 -1405
rect 16820 -1440 16825 -1410
rect 16855 -1440 16860 -1410
rect 16820 -1450 16860 -1440
rect 16820 -1480 16825 -1450
rect 16855 -1480 16860 -1450
rect 16820 -1490 16860 -1480
rect 16820 -1520 16825 -1490
rect 16855 -1520 16860 -1490
rect 16820 -1525 16860 -1520
rect 17025 -1410 17065 -1405
rect 17025 -1440 17030 -1410
rect 17060 -1440 17065 -1410
rect 17025 -1450 17065 -1440
rect 17025 -1480 17030 -1450
rect 17060 -1480 17065 -1450
rect 17025 -1490 17065 -1480
rect 17025 -1520 17030 -1490
rect 17060 -1520 17065 -1490
rect 17025 -1525 17065 -1520
rect 17135 -1410 17175 -1405
rect 17135 -1440 17140 -1410
rect 17170 -1440 17175 -1410
rect 17135 -1450 17175 -1440
rect 17135 -1480 17140 -1450
rect 17170 -1480 17175 -1450
rect 17135 -1490 17175 -1480
rect 17135 -1520 17140 -1490
rect 17170 -1520 17175 -1490
rect 17135 -1525 17175 -1520
rect 17245 -1410 17285 -1405
rect 17245 -1440 17250 -1410
rect 17280 -1440 17285 -1410
rect 17245 -1450 17285 -1440
rect 17245 -1480 17250 -1450
rect 17280 -1480 17285 -1450
rect 17245 -1490 17285 -1480
rect 17310 -1485 17330 -1360
rect 17355 -1410 17395 -1405
rect 17355 -1440 17360 -1410
rect 17390 -1440 17395 -1410
rect 17355 -1450 17395 -1440
rect 17355 -1480 17360 -1450
rect 17390 -1480 17395 -1450
rect 17245 -1520 17250 -1490
rect 17280 -1520 17285 -1490
rect 17245 -1525 17285 -1520
rect 17305 -1495 17335 -1485
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17305 -1525 17335 -1515
rect 17355 -1490 17395 -1480
rect 17355 -1520 17360 -1490
rect 17390 -1520 17395 -1490
rect 17355 -1525 17395 -1520
rect 17465 -1410 17505 -1405
rect 17465 -1440 17470 -1410
rect 17500 -1440 17505 -1410
rect 17465 -1450 17505 -1440
rect 17465 -1480 17470 -1450
rect 17500 -1480 17505 -1450
rect 17465 -1490 17505 -1480
rect 17465 -1520 17470 -1490
rect 17500 -1520 17505 -1490
rect 17465 -1525 17505 -1520
rect 17615 -1410 17655 -1405
rect 17615 -1440 17620 -1410
rect 17650 -1440 17655 -1410
rect 17615 -1450 17655 -1440
rect 17615 -1480 17620 -1450
rect 17650 -1480 17655 -1450
rect 17615 -1490 17655 -1480
rect 17615 -1520 17620 -1490
rect 17650 -1520 17655 -1490
rect 17615 -1525 17655 -1520
rect 17725 -1410 17765 -1405
rect 17725 -1440 17730 -1410
rect 17760 -1440 17765 -1410
rect 17725 -1450 17765 -1440
rect 17725 -1480 17730 -1450
rect 17760 -1480 17765 -1450
rect 17725 -1490 17765 -1480
rect 17790 -1485 17810 -1360
rect 17835 -1410 17875 -1405
rect 17835 -1440 17840 -1410
rect 17870 -1440 17875 -1410
rect 17835 -1450 17875 -1440
rect 17835 -1480 17840 -1450
rect 17870 -1480 17875 -1450
rect 17725 -1520 17730 -1490
rect 17760 -1520 17765 -1490
rect 17725 -1525 17765 -1520
rect 17785 -1495 17815 -1485
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17785 -1525 17815 -1515
rect 17835 -1490 17875 -1480
rect 17835 -1520 17840 -1490
rect 17870 -1520 17875 -1490
rect 17835 -1525 17875 -1520
rect 17945 -1410 17985 -1405
rect 17945 -1440 17950 -1410
rect 17980 -1440 17985 -1410
rect 17945 -1450 17985 -1440
rect 17945 -1480 17950 -1450
rect 17980 -1480 17985 -1450
rect 17945 -1490 17985 -1480
rect 17945 -1520 17950 -1490
rect 17980 -1520 17985 -1490
rect 17945 -1525 17985 -1520
rect 18095 -1410 18135 -1405
rect 18095 -1440 18100 -1410
rect 18130 -1440 18135 -1410
rect 18095 -1450 18135 -1440
rect 18095 -1480 18100 -1450
rect 18130 -1480 18135 -1450
rect 18095 -1490 18135 -1480
rect 18095 -1520 18100 -1490
rect 18130 -1520 18135 -1490
rect 18095 -1525 18135 -1520
rect 18205 -1410 18245 -1405
rect 18205 -1440 18210 -1410
rect 18240 -1440 18245 -1410
rect 18205 -1450 18245 -1440
rect 18205 -1480 18210 -1450
rect 18240 -1480 18245 -1450
rect 18205 -1490 18245 -1480
rect 18270 -1485 18290 -1360
rect 18315 -1410 18355 -1405
rect 18315 -1440 18320 -1410
rect 18350 -1440 18355 -1410
rect 18315 -1450 18355 -1440
rect 18315 -1480 18320 -1450
rect 18350 -1480 18355 -1450
rect 18205 -1520 18210 -1490
rect 18240 -1520 18245 -1490
rect 18205 -1525 18245 -1520
rect 18265 -1495 18295 -1485
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18265 -1525 18295 -1515
rect 18315 -1490 18355 -1480
rect 18315 -1520 18320 -1490
rect 18350 -1520 18355 -1490
rect 18315 -1525 18355 -1520
rect 18425 -1410 18465 -1405
rect 18425 -1440 18430 -1410
rect 18460 -1440 18465 -1410
rect 18425 -1450 18465 -1440
rect 18425 -1480 18430 -1450
rect 18460 -1480 18465 -1450
rect 18425 -1490 18465 -1480
rect 18425 -1520 18430 -1490
rect 18460 -1520 18465 -1490
rect 18425 -1525 18465 -1520
rect 18535 -1410 18575 -1405
rect 18535 -1440 18540 -1410
rect 18570 -1440 18575 -1410
rect 18535 -1450 18575 -1440
rect 18535 -1480 18540 -1450
rect 18570 -1480 18575 -1450
rect 18535 -1490 18575 -1480
rect 18535 -1520 18540 -1490
rect 18570 -1520 18575 -1490
rect 18535 -1525 18575 -1520
rect 17195 -1555 17225 -1545
rect 17195 -1575 17200 -1555
rect 17220 -1575 17225 -1555
rect 17195 -1605 17225 -1575
rect 17195 -1625 17200 -1605
rect 17220 -1625 17225 -1605
rect 17195 -1655 17225 -1625
rect 17415 -1555 17445 -1545
rect 17415 -1575 17420 -1555
rect 17440 -1575 17445 -1555
rect 17415 -1605 17445 -1575
rect 17415 -1625 17420 -1605
rect 17440 -1625 17445 -1605
rect 17415 -1655 17445 -1625
rect 18155 -1555 18185 -1545
rect 18155 -1575 18160 -1555
rect 18180 -1575 18185 -1555
rect 18155 -1605 18185 -1575
rect 18155 -1625 18160 -1605
rect 18180 -1625 18185 -1605
rect 18155 -1655 18185 -1625
rect 18375 -1555 18405 -1545
rect 18375 -1575 18380 -1555
rect 18400 -1575 18405 -1555
rect 18375 -1605 18405 -1575
rect 18375 -1625 18380 -1605
rect 18400 -1625 18405 -1605
rect 18375 -1655 18405 -1625
rect 16705 -1665 16745 -1655
rect 16705 -1685 16715 -1665
rect 16735 -1685 16745 -1665
rect 16705 -1695 16745 -1685
rect 17080 -1665 17120 -1655
rect 17080 -1685 17090 -1665
rect 17110 -1685 17120 -1665
rect 17080 -1695 17120 -1685
rect 17190 -1660 17230 -1655
rect 17190 -1690 17195 -1660
rect 17225 -1690 17230 -1660
rect 16715 -1895 16735 -1695
rect 17090 -1710 17110 -1695
rect 17080 -1715 17120 -1710
rect 17080 -1745 17085 -1715
rect 17115 -1745 17120 -1715
rect 17080 -1750 17120 -1745
rect 17190 -1770 17230 -1690
rect 17300 -1665 17340 -1655
rect 17300 -1685 17310 -1665
rect 17330 -1685 17340 -1665
rect 17300 -1695 17340 -1685
rect 17410 -1660 17450 -1655
rect 17410 -1690 17415 -1660
rect 17445 -1690 17450 -1660
rect 17410 -1695 17450 -1690
rect 17670 -1660 17710 -1655
rect 17670 -1690 17675 -1660
rect 17705 -1690 17710 -1660
rect 17670 -1695 17710 -1690
rect 17780 -1660 17820 -1655
rect 17780 -1690 17785 -1660
rect 17815 -1690 17820 -1660
rect 17780 -1695 17820 -1690
rect 17890 -1660 17930 -1655
rect 17890 -1690 17895 -1660
rect 17925 -1690 17930 -1660
rect 17890 -1695 17930 -1690
rect 18150 -1660 18190 -1655
rect 18150 -1690 18155 -1660
rect 18185 -1690 18190 -1660
rect 18150 -1695 18190 -1690
rect 18260 -1665 18300 -1655
rect 18260 -1685 18270 -1665
rect 18290 -1685 18300 -1665
rect 18260 -1695 18300 -1685
rect 18370 -1660 18410 -1655
rect 18370 -1690 18375 -1660
rect 18405 -1690 18410 -1660
rect 17310 -1710 17330 -1695
rect 17300 -1715 17340 -1710
rect 17300 -1745 17305 -1715
rect 17335 -1745 17340 -1715
rect 17300 -1750 17340 -1745
rect 17190 -1800 17195 -1770
rect 17225 -1800 17230 -1770
rect 17190 -1810 17230 -1800
rect 17190 -1840 17195 -1810
rect 17225 -1840 17230 -1810
rect 17190 -1845 17230 -1840
rect 17790 -1895 17810 -1695
rect 18270 -1710 18290 -1695
rect 18260 -1715 18300 -1710
rect 18260 -1745 18265 -1715
rect 18295 -1745 18300 -1715
rect 18260 -1750 18300 -1745
rect 18370 -1770 18410 -1690
rect 18480 -1665 18520 -1655
rect 18480 -1685 18490 -1665
rect 18510 -1685 18520 -1665
rect 18480 -1695 18520 -1685
rect 18490 -1710 18510 -1695
rect 18480 -1715 18520 -1710
rect 18480 -1745 18485 -1715
rect 18515 -1745 18520 -1715
rect 18480 -1750 18520 -1745
rect 18370 -1800 18375 -1770
rect 18405 -1800 18410 -1770
rect 18370 -1810 18410 -1800
rect 18370 -1840 18375 -1810
rect 18405 -1840 18410 -1810
rect 18370 -1845 18410 -1840
rect 16705 -1900 16745 -1895
rect 16705 -1930 16710 -1900
rect 16740 -1930 16745 -1900
rect 16705 -1935 16745 -1930
rect 17780 -1900 17820 -1895
rect 17780 -1930 17785 -1900
rect 17815 -1930 17820 -1900
rect 17780 -1935 17820 -1930
rect 19335 -1945 19355 -665
rect 19325 -1950 19365 -1945
rect 19325 -1980 19330 -1950
rect 19360 -1980 19365 -1950
rect 19325 -1985 19365 -1980
rect 16260 -2000 16300 -1995
rect 16260 -2030 16265 -2000
rect 16295 -2030 16300 -2000
rect 16260 -2035 16300 -2030
rect 16480 -2000 16520 -1995
rect 16480 -2030 16485 -2000
rect 16515 -2030 16520 -2000
rect 16480 -2035 16520 -2030
rect 16730 -2000 16770 -1995
rect 16730 -2030 16735 -2000
rect 16765 -2030 16770 -2000
rect 16730 -2035 16770 -2030
rect 17195 -2000 17235 -1995
rect 17195 -2030 17200 -2000
rect 17230 -2030 17235 -2000
rect 16490 -2895 16510 -2035
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16160 -3025 16195 -3020
rect 16160 -3065 16195 -3060
rect 16740 -3100 16760 -2035
rect 17195 -2060 17235 -2030
rect 17425 -2035 17430 -2000
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2035 18169 -2000
rect 19080 -2005 19120 -2000
rect 19080 -2035 19085 -2005
rect 19115 -2035 19120 -2005
rect 17195 -2090 17200 -2060
rect 17230 -2090 17235 -2060
rect 17195 -2095 17235 -2090
rect 18830 -2060 18870 -2055
rect 18830 -2090 18835 -2060
rect 18865 -2090 18870 -2060
rect 18830 -2095 18870 -2090
rect 16945 -2615 18655 -2265
rect 16730 -3105 16770 -3100
rect 15820 -3145 15825 -3115
rect 15855 -3145 15860 -3115
rect 15820 -3150 15860 -3145
rect 15950 -3116 15985 -3111
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 15830 -4260 15850 -3150
rect 15950 -3156 15985 -3151
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18840 -3100 18860 -2095
rect 19080 -2895 19120 -2035
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19415 -2992 19435 -345
rect 19460 -2005 19500 415
rect 19545 -1895 19565 1595
rect 19610 250 19650 255
rect 19610 220 19615 250
rect 19645 220 19650 250
rect 19610 215 19650 220
rect 19535 -1900 19575 -1895
rect 19535 -1930 19540 -1900
rect 19570 -1930 19575 -1900
rect 19535 -1935 19575 -1930
rect 19460 -2035 19465 -2005
rect 19495 -2035 19500 -2005
rect 19460 -2040 19500 -2035
rect 19405 -2997 19440 -2992
rect 19405 -3037 19440 -3032
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -3100
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 19620 -3111 19640 215
rect 19720 -255 19760 -250
rect 19720 -285 19725 -255
rect 19755 -285 19760 -255
rect 19720 -290 19760 -285
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4295 15860 -4265
rect 15820 -4300 15860 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4345 15765 -4315
rect 15725 -4350 15765 -4345
rect 15960 -4355 15980 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 16290 -4185 16310 -3934
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 18960 -3969 18995 -3964
rect 16605 -4009 16640 -4004
rect 18960 -4009 18995 -4004
rect 16615 -4185 16635 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4220 16285 -4190
rect 16315 -4220 16320 -4190
rect 16280 -4225 16320 -4220
rect 16605 -4190 16645 -4185
rect 16605 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 17250 -4265 17300 -4255
rect 18965 -4260 18985 -4009
rect 19290 -4260 19310 -3934
rect 17250 -4295 17260 -4265
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4295 17820 -4265
rect 17780 -4300 17820 -4295
rect 18955 -4265 18995 -4260
rect 18955 -4295 18960 -4265
rect 18990 -4295 18995 -4265
rect 18955 -4300 18995 -4295
rect 19280 -4265 19320 -4260
rect 19280 -4295 19285 -4265
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 16900 -4315 16950 -4305
rect 16900 -4345 16910 -4315
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4345 18700 -4315
rect 18650 -4355 18700 -4345
rect 19620 -4355 19640 -3829
rect 19730 -4310 19750 -290
rect 19775 -1770 19815 1595
rect 19775 -1800 19780 -1770
rect 19810 -1800 19815 -1770
rect 19775 -1810 19815 -1800
rect 19775 -1840 19780 -1810
rect 19810 -1840 19815 -1810
rect 19775 -1845 19815 -1840
rect 19720 -4315 19760 -4310
rect 19720 -4345 19725 -4315
rect 19755 -4345 19760 -4315
rect 19720 -4350 19760 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4390 15990 -4360
rect 15950 -4395 15990 -4390
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 19355 -4395 19395 -4390
rect 19610 -4360 19650 -4355
rect 19610 -4390 19615 -4360
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4445 17995 -4440
<< via1 >>
rect 15730 -285 15760 -255
rect 15955 -55 15985 -25
rect 15790 -1800 15820 -1770
rect 15790 -1840 15820 -1810
rect 16035 -1745 16065 -1715
rect 16945 1475 16975 1505
rect 16490 1455 16520 1460
rect 16490 1435 16495 1455
rect 16495 1435 16515 1455
rect 16515 1435 16520 1455
rect 16490 1430 16520 1435
rect 16370 1330 16400 1360
rect 16370 1290 16400 1320
rect 16370 1275 16400 1280
rect 16370 1255 16375 1275
rect 16375 1255 16395 1275
rect 16395 1255 16400 1275
rect 16370 1250 16400 1255
rect 16490 1330 16520 1360
rect 16490 1290 16520 1320
rect 16490 1275 16520 1280
rect 16490 1255 16495 1275
rect 16495 1255 16515 1275
rect 16515 1255 16520 1275
rect 16490 1250 16520 1255
rect 16610 1330 16640 1360
rect 16610 1290 16640 1320
rect 16610 1275 16640 1280
rect 16610 1255 16615 1275
rect 16615 1255 16635 1275
rect 16635 1255 16640 1275
rect 16610 1250 16640 1255
rect 16890 1330 16920 1360
rect 16890 1290 16920 1320
rect 17055 1430 17085 1460
rect 17000 1330 17030 1360
rect 17000 1290 17030 1320
rect 16890 1275 16920 1280
rect 16890 1255 16895 1275
rect 16895 1255 16915 1275
rect 16915 1255 16920 1275
rect 16890 1250 16920 1255
rect 17110 1330 17140 1360
rect 17110 1290 17140 1320
rect 17000 1275 17030 1280
rect 17000 1255 17005 1275
rect 17005 1255 17025 1275
rect 17025 1255 17030 1275
rect 17000 1250 17030 1255
rect 17110 1275 17140 1280
rect 17110 1255 17115 1275
rect 17115 1255 17135 1275
rect 17135 1255 17140 1275
rect 17110 1250 17140 1255
rect 17220 1330 17250 1360
rect 17220 1290 17250 1320
rect 17220 1275 17250 1280
rect 17220 1255 17225 1275
rect 17225 1255 17245 1275
rect 17245 1255 17250 1275
rect 17220 1250 17250 1255
rect 17500 1330 17530 1360
rect 17500 1290 17530 1320
rect 17500 1275 17530 1280
rect 17500 1255 17505 1275
rect 17505 1255 17525 1275
rect 17525 1255 17530 1275
rect 17500 1250 17530 1255
rect 17565 1330 17595 1360
rect 17565 1290 17595 1320
rect 17565 1275 17595 1280
rect 17565 1255 17570 1275
rect 17570 1255 17590 1275
rect 17590 1255 17595 1275
rect 17565 1250 17595 1255
rect 17675 1330 17705 1360
rect 17675 1290 17705 1320
rect 17675 1275 17705 1280
rect 17675 1255 17680 1275
rect 17680 1255 17700 1275
rect 17700 1255 17705 1275
rect 17675 1250 17705 1255
rect 17785 1455 17815 1460
rect 17785 1435 17790 1455
rect 17790 1435 17810 1455
rect 17810 1435 17815 1455
rect 17785 1430 17815 1435
rect 17785 1330 17815 1360
rect 17785 1290 17815 1320
rect 17785 1275 17815 1280
rect 17785 1255 17790 1275
rect 17790 1255 17810 1275
rect 17810 1255 17815 1275
rect 17785 1250 17815 1255
rect 17895 1330 17925 1360
rect 17895 1290 17925 1320
rect 17895 1275 17925 1280
rect 17895 1255 17900 1275
rect 17900 1255 17920 1275
rect 17920 1255 17925 1275
rect 17895 1250 17925 1255
rect 18625 1475 18655 1505
rect 18205 1430 18235 1460
rect 18515 1430 18545 1460
rect 18005 1330 18035 1360
rect 18005 1290 18035 1320
rect 18005 1275 18035 1280
rect 18005 1255 18010 1275
rect 18010 1255 18030 1275
rect 18030 1255 18035 1275
rect 18005 1250 18035 1255
rect 18070 1330 18100 1360
rect 18070 1290 18100 1320
rect 18070 1275 18100 1280
rect 18070 1255 18075 1275
rect 18075 1255 18095 1275
rect 18095 1255 18100 1275
rect 18070 1250 18100 1255
rect 16435 1105 16465 1110
rect 16435 1085 16440 1105
rect 16440 1085 16460 1105
rect 16460 1085 16465 1105
rect 16435 1080 16465 1085
rect 16545 1105 16575 1110
rect 16545 1085 16550 1105
rect 16550 1085 16570 1105
rect 16570 1085 16575 1105
rect 16545 1080 16575 1085
rect 16945 1105 16975 1110
rect 16945 1085 16950 1105
rect 16950 1085 16970 1105
rect 16970 1085 16975 1105
rect 16945 1080 16975 1085
rect 17055 1105 17085 1110
rect 17055 1085 17060 1105
rect 17060 1085 17080 1105
rect 17080 1085 17085 1105
rect 17055 1080 17085 1085
rect 17165 1105 17195 1110
rect 17165 1085 17170 1105
rect 17170 1085 17190 1105
rect 17190 1085 17195 1105
rect 17165 1080 17195 1085
rect 17620 1105 17650 1110
rect 17620 1085 17625 1105
rect 17625 1085 17645 1105
rect 17645 1085 17650 1105
rect 17620 1080 17650 1085
rect 17730 1105 17760 1110
rect 17730 1085 17735 1105
rect 17735 1085 17755 1105
rect 17755 1085 17760 1105
rect 17730 1080 17760 1085
rect 17840 1105 17870 1110
rect 17840 1085 17845 1105
rect 17845 1085 17865 1105
rect 17865 1085 17870 1105
rect 17840 1080 17870 1085
rect 17950 1105 17980 1110
rect 17950 1085 17955 1105
rect 17955 1085 17975 1105
rect 17975 1085 17980 1105
rect 17950 1080 17980 1085
rect 18350 1330 18380 1360
rect 18350 1290 18380 1320
rect 18350 1275 18380 1280
rect 18350 1255 18355 1275
rect 18355 1255 18375 1275
rect 18375 1255 18380 1275
rect 18350 1250 18380 1255
rect 18460 1330 18490 1360
rect 18460 1290 18490 1320
rect 18570 1330 18600 1360
rect 18570 1290 18600 1320
rect 18460 1275 18490 1280
rect 18460 1255 18465 1275
rect 18465 1255 18485 1275
rect 18485 1255 18490 1275
rect 18460 1250 18490 1255
rect 18680 1330 18710 1360
rect 18680 1290 18710 1320
rect 18570 1275 18600 1280
rect 18570 1255 18575 1275
rect 18575 1255 18595 1275
rect 18595 1255 18600 1275
rect 18570 1250 18600 1255
rect 18680 1275 18710 1280
rect 18680 1255 18685 1275
rect 18685 1255 18705 1275
rect 18705 1255 18710 1275
rect 18680 1250 18710 1255
rect 18405 1105 18435 1110
rect 18405 1085 18410 1105
rect 18410 1085 18430 1105
rect 18430 1085 18435 1105
rect 18405 1080 18435 1085
rect 18515 1105 18545 1110
rect 18515 1085 18520 1105
rect 18520 1085 18540 1105
rect 18540 1085 18545 1105
rect 18515 1080 18545 1085
rect 18625 1105 18655 1110
rect 18625 1085 18630 1105
rect 18630 1085 18650 1105
rect 18650 1085 18655 1105
rect 18625 1080 18655 1085
rect 18205 1025 18235 1055
rect 18725 1025 18755 1055
rect 16165 980 16195 1010
rect 16435 980 16465 1010
rect 16545 980 16575 1010
rect 16440 905 16470 935
rect 16440 865 16470 895
rect 16440 825 16470 855
rect 16440 785 16470 815
rect 16660 905 16690 935
rect 16660 865 16690 895
rect 16660 825 16690 855
rect 16660 785 16690 815
rect 16975 905 17005 935
rect 16975 865 17005 895
rect 16975 825 17005 855
rect 16975 810 17005 815
rect 16975 790 16980 810
rect 16980 790 17000 810
rect 17000 790 17005 810
rect 16975 785 17005 790
rect 17155 905 17185 935
rect 17155 865 17185 895
rect 17155 825 17185 855
rect 17155 810 17185 815
rect 17155 790 17160 810
rect 17160 790 17180 810
rect 17180 790 17185 810
rect 17155 785 17185 790
rect 17335 905 17365 935
rect 17335 865 17365 895
rect 17335 825 17365 855
rect 17335 810 17365 815
rect 17335 790 17340 810
rect 17340 790 17360 810
rect 17360 790 17365 810
rect 17335 785 17365 790
rect 17515 905 17545 935
rect 17515 865 17545 895
rect 17515 825 17545 855
rect 17515 810 17545 815
rect 17515 790 17520 810
rect 17520 790 17540 810
rect 17540 790 17545 810
rect 17515 785 17545 790
rect 17695 905 17725 935
rect 17695 865 17725 895
rect 17695 825 17725 855
rect 17695 810 17725 815
rect 17695 790 17700 810
rect 17700 790 17720 810
rect 17720 790 17725 810
rect 17695 785 17725 790
rect 17875 905 17905 935
rect 17875 865 17905 895
rect 17875 825 17905 855
rect 17875 810 17905 815
rect 17875 790 17880 810
rect 17880 790 17900 810
rect 17900 790 17905 810
rect 17875 785 17905 790
rect 18055 905 18085 935
rect 18055 865 18085 895
rect 18055 825 18085 855
rect 18055 810 18085 815
rect 18055 790 18060 810
rect 18060 790 18080 810
rect 18080 790 18085 810
rect 18055 785 18085 790
rect 18235 905 18265 935
rect 18235 865 18265 895
rect 18235 825 18265 855
rect 18235 810 18265 815
rect 18235 790 18240 810
rect 18240 790 18260 810
rect 18260 790 18265 810
rect 18235 785 18265 790
rect 18415 905 18445 935
rect 18415 865 18445 895
rect 18415 825 18445 855
rect 18415 810 18445 815
rect 18415 790 18420 810
rect 18420 790 18440 810
rect 18440 790 18445 810
rect 18415 785 18445 790
rect 18595 905 18625 935
rect 18595 865 18625 895
rect 18595 825 18625 855
rect 18595 810 18625 815
rect 18595 790 18600 810
rect 18600 790 18620 810
rect 18620 790 18625 810
rect 18595 785 18625 790
rect 16550 710 16580 715
rect 16550 690 16555 710
rect 16555 690 16575 710
rect 16575 690 16580 710
rect 16550 685 16580 690
rect 16785 685 16815 715
rect 16485 540 16515 545
rect 16485 520 16490 540
rect 16490 520 16510 540
rect 16510 520 16515 540
rect 16485 515 16515 520
rect 16615 540 16645 545
rect 16615 520 16620 540
rect 16620 520 16640 540
rect 16640 520 16645 540
rect 16615 515 16645 520
rect 16320 415 16350 445
rect 16265 360 16295 390
rect 16210 315 16240 345
rect 16265 -340 16295 -310
rect 16210 -1255 16240 -1225
rect 16165 -1355 16195 -1325
rect 16110 -1930 16140 -1900
rect 16160 -1980 16190 -1950
rect 16845 515 16875 545
rect 16785 360 16815 390
rect 16550 315 16580 345
rect 16425 80 16455 110
rect 16425 40 16455 70
rect 16425 0 16455 30
rect 16545 80 16575 110
rect 16545 40 16575 70
rect 16545 0 16575 30
rect 16665 80 16695 110
rect 16665 40 16695 70
rect 16665 0 16695 30
rect 16785 80 16815 110
rect 16785 40 16815 70
rect 16785 0 16815 30
rect 17605 440 17635 445
rect 17605 420 17610 440
rect 17610 420 17630 440
rect 17630 420 17635 440
rect 17605 415 17635 420
rect 17965 440 17995 445
rect 17965 420 17970 440
rect 17970 420 17990 440
rect 17990 420 17995 440
rect 17965 415 17995 420
rect 17425 360 17455 390
rect 17245 315 17275 345
rect 17065 270 17095 300
rect 16905 80 16935 110
rect 16905 40 16935 70
rect 16905 0 16935 30
rect 17025 80 17055 110
rect 17025 40 17055 70
rect 17025 0 17055 30
rect 17145 80 17175 110
rect 17145 40 17175 70
rect 17145 0 17175 30
rect 17265 80 17295 110
rect 17265 40 17295 70
rect 17265 0 17295 30
rect 17385 80 17415 110
rect 17385 40 17415 70
rect 17385 0 17415 30
rect 17505 80 17535 110
rect 17505 40 17535 70
rect 17505 0 17535 30
rect 17625 80 17655 110
rect 17625 40 17655 70
rect 17625 0 17655 30
rect 18145 360 18175 390
rect 18325 315 18355 345
rect 17785 270 17815 300
rect 18505 270 18535 300
rect 18910 905 18940 935
rect 18910 865 18940 895
rect 18910 825 18940 855
rect 18910 810 18940 815
rect 18910 790 18915 810
rect 18915 790 18935 810
rect 18935 790 18940 810
rect 18910 785 18940 790
rect 19020 905 19050 935
rect 19020 865 19050 895
rect 19020 825 19050 855
rect 19020 810 19050 815
rect 19020 790 19025 810
rect 19025 790 19045 810
rect 19045 790 19050 810
rect 19020 785 19050 790
rect 19080 905 19110 935
rect 19080 865 19110 895
rect 19080 825 19110 855
rect 19080 810 19110 815
rect 19080 790 19085 810
rect 19085 790 19105 810
rect 19105 790 19110 810
rect 19080 785 19110 790
rect 19330 980 19360 1010
rect 18955 540 18985 545
rect 18955 520 18960 540
rect 18960 520 18980 540
rect 18980 520 18985 540
rect 18955 515 18985 520
rect 19265 515 19295 545
rect 19005 490 19035 495
rect 19005 470 19010 490
rect 19010 470 19030 490
rect 19030 470 19035 490
rect 19005 465 19035 470
rect 18005 220 18035 250
rect 18725 220 18755 250
rect 19015 220 19045 250
rect 17945 80 17975 110
rect 17945 40 17975 70
rect 17945 0 17975 30
rect 18065 80 18095 110
rect 18065 40 18095 70
rect 18065 0 18095 30
rect 18185 80 18215 110
rect 18185 40 18215 70
rect 18185 0 18215 30
rect 18305 80 18335 110
rect 18305 40 18335 70
rect 18305 0 18335 30
rect 18425 80 18455 110
rect 18425 40 18455 70
rect 18425 0 18455 30
rect 18545 80 18575 110
rect 18545 40 18575 70
rect 18545 0 18575 30
rect 18665 80 18695 110
rect 18665 40 18695 70
rect 18665 0 18695 30
rect 18785 80 18815 110
rect 18785 40 18815 70
rect 18785 0 18815 30
rect 18905 80 18935 110
rect 18905 40 18935 70
rect 18905 0 18935 30
rect 19025 80 19055 110
rect 19025 40 19055 70
rect 19025 0 19055 30
rect 19145 80 19175 110
rect 19145 40 19175 70
rect 19145 0 19175 30
rect 16485 -30 16515 -25
rect 16485 -50 16490 -30
rect 16490 -50 16510 -30
rect 16510 -50 16515 -30
rect 16485 -55 16515 -50
rect 16845 -30 16875 -25
rect 16845 -50 16850 -30
rect 16850 -50 16870 -30
rect 16870 -50 16875 -30
rect 16845 -55 16875 -50
rect 17205 -30 17235 -25
rect 17205 -50 17210 -30
rect 17210 -50 17230 -30
rect 17230 -50 17235 -30
rect 17205 -55 17235 -50
rect 17565 -30 17595 -25
rect 17565 -50 17570 -30
rect 17570 -50 17590 -30
rect 17590 -50 17595 -30
rect 17565 -55 17595 -50
rect 17695 -55 17725 -25
rect 17875 -55 17905 -25
rect 16605 -200 16635 -195
rect 16605 -220 16610 -200
rect 16610 -220 16630 -200
rect 16630 -220 16635 -200
rect 16605 -225 16635 -220
rect 16965 -200 16995 -195
rect 16965 -220 16970 -200
rect 16970 -220 16990 -200
rect 16990 -220 16995 -200
rect 16965 -225 16995 -220
rect 17325 -200 17355 -195
rect 17325 -220 17330 -200
rect 17330 -220 17350 -200
rect 17350 -220 17355 -200
rect 17325 -225 17355 -220
rect 16515 -285 16545 -255
rect 16725 -285 16755 -255
rect 16845 -285 16875 -255
rect 17085 -285 17115 -255
rect 17205 -285 17235 -255
rect 17445 -285 17475 -255
rect 17535 -285 17565 -255
rect 17007 -315 17037 -310
rect 17007 -335 17012 -315
rect 17012 -335 17032 -315
rect 17032 -335 17037 -315
rect 17007 -340 17037 -335
rect 16320 -660 16350 -630
rect 17565 -375 17595 -370
rect 17565 -395 17570 -375
rect 17570 -395 17590 -375
rect 17590 -395 17595 -375
rect 17565 -400 17595 -395
rect 17075 -635 17105 -630
rect 17075 -655 17080 -635
rect 17080 -655 17100 -635
rect 17100 -655 17105 -635
rect 17075 -660 17105 -655
rect 16535 -740 16565 -710
rect 17025 -740 17055 -710
rect 16625 -770 16655 -765
rect 16625 -790 16630 -770
rect 16630 -790 16650 -770
rect 16650 -790 16655 -770
rect 16625 -795 16655 -790
rect 16745 -770 16775 -765
rect 16745 -790 16750 -770
rect 16750 -790 16770 -770
rect 16770 -790 16775 -770
rect 16745 -795 16775 -790
rect 16865 -770 16895 -765
rect 16865 -790 16870 -770
rect 16870 -790 16890 -770
rect 16890 -790 16895 -770
rect 16865 -795 16895 -790
rect 16985 -770 17015 -765
rect 16985 -790 16990 -770
rect 16990 -790 17010 -770
rect 17010 -790 17015 -770
rect 16985 -795 17015 -790
rect 17305 -770 17335 -765
rect 17305 -790 17310 -770
rect 17310 -790 17330 -770
rect 17330 -790 17335 -770
rect 17305 -795 17335 -790
rect 17425 -770 17455 -765
rect 17425 -790 17430 -770
rect 17430 -790 17450 -770
rect 17450 -790 17455 -770
rect 17425 -795 17455 -790
rect 17545 -770 17575 -765
rect 17545 -790 17550 -770
rect 17550 -790 17570 -770
rect 17570 -790 17575 -770
rect 17545 -795 17575 -790
rect 17785 -400 17815 -370
rect 18005 -30 18035 -25
rect 18005 -50 18010 -30
rect 18010 -50 18030 -30
rect 18030 -50 18035 -30
rect 18005 -55 18035 -50
rect 18365 -30 18395 -25
rect 18365 -50 18370 -30
rect 18370 -50 18390 -30
rect 18390 -50 18395 -30
rect 18365 -55 18395 -50
rect 18725 -30 18755 -25
rect 18725 -50 18730 -30
rect 18730 -50 18750 -30
rect 18750 -50 18755 -30
rect 18725 -55 18755 -50
rect 19085 -30 19115 -25
rect 19085 -50 19090 -30
rect 19090 -50 19110 -30
rect 19110 -50 19115 -30
rect 19085 -55 19115 -50
rect 18245 -200 18275 -195
rect 18245 -220 18250 -200
rect 18250 -220 18270 -200
rect 18270 -220 18275 -200
rect 18245 -225 18275 -220
rect 18605 -200 18635 -195
rect 18605 -220 18610 -200
rect 18610 -220 18630 -200
rect 18630 -220 18635 -200
rect 18605 -225 18635 -220
rect 18965 -200 18995 -195
rect 18965 -220 18970 -200
rect 18970 -220 18990 -200
rect 18990 -220 18995 -200
rect 18965 -225 18995 -220
rect 18035 -285 18065 -255
rect 18125 -285 18155 -255
rect 18365 -285 18395 -255
rect 18485 -285 18515 -255
rect 18725 -285 18755 -255
rect 18845 -285 18875 -255
rect 19055 -285 19085 -255
rect 18563 -315 18593 -310
rect 18563 -335 18568 -315
rect 18568 -335 18588 -315
rect 18588 -335 18593 -315
rect 18563 -340 18593 -335
rect 18005 -375 18035 -370
rect 18005 -395 18010 -375
rect 18010 -395 18030 -375
rect 18030 -395 18035 -375
rect 18005 -400 18035 -395
rect 19465 415 19495 445
rect 19410 270 19440 300
rect 19410 -340 19440 -310
rect 18495 -635 18525 -630
rect 18495 -655 18500 -635
rect 18500 -655 18520 -635
rect 18520 -655 18525 -635
rect 18495 -660 18525 -655
rect 19330 -660 19360 -630
rect 18545 -740 18575 -710
rect 19035 -740 19065 -710
rect 18025 -770 18055 -765
rect 18025 -790 18030 -770
rect 18030 -790 18050 -770
rect 18050 -790 18055 -770
rect 18025 -795 18055 -790
rect 18145 -770 18175 -765
rect 18145 -790 18150 -770
rect 18150 -790 18170 -770
rect 18170 -790 18175 -770
rect 18145 -795 18175 -790
rect 18265 -770 18295 -765
rect 18265 -790 18270 -770
rect 18270 -790 18290 -770
rect 18290 -790 18295 -770
rect 18265 -795 18295 -790
rect 18585 -770 18615 -765
rect 18585 -790 18590 -770
rect 18590 -790 18610 -770
rect 18610 -790 18615 -770
rect 18585 -795 18615 -790
rect 18705 -770 18735 -765
rect 18705 -790 18710 -770
rect 18710 -790 18730 -770
rect 18730 -790 18735 -770
rect 18705 -795 18735 -790
rect 18825 -770 18855 -765
rect 18825 -790 18830 -770
rect 18830 -790 18850 -770
rect 18850 -790 18855 -770
rect 18825 -795 18855 -790
rect 18945 -770 18975 -765
rect 18945 -790 18950 -770
rect 18950 -790 18970 -770
rect 18970 -790 18975 -770
rect 18945 -795 18975 -790
rect 17115 -1085 17145 -1080
rect 17115 -1105 17120 -1085
rect 17120 -1105 17140 -1085
rect 17140 -1105 17145 -1085
rect 17115 -1110 17145 -1105
rect 17785 -1110 17815 -1080
rect 18455 -1085 18485 -1080
rect 18455 -1105 18460 -1085
rect 18460 -1105 18480 -1085
rect 18480 -1105 18485 -1085
rect 18455 -1110 18485 -1105
rect 16745 -1145 16775 -1140
rect 16745 -1165 16750 -1145
rect 16750 -1165 16770 -1145
rect 16770 -1165 16775 -1145
rect 16745 -1170 16775 -1165
rect 16825 -1145 16855 -1140
rect 16825 -1165 16830 -1145
rect 16830 -1165 16850 -1145
rect 16850 -1165 16855 -1145
rect 16825 -1170 16855 -1165
rect 16905 -1145 16935 -1140
rect 16905 -1165 16910 -1145
rect 16910 -1165 16930 -1145
rect 16930 -1165 16935 -1145
rect 16905 -1170 16935 -1165
rect 16985 -1145 17015 -1140
rect 16985 -1165 16990 -1145
rect 16990 -1165 17010 -1145
rect 17010 -1165 17015 -1145
rect 16985 -1170 17015 -1165
rect 17065 -1145 17095 -1140
rect 17065 -1165 17070 -1145
rect 17070 -1165 17090 -1145
rect 17090 -1165 17095 -1145
rect 17065 -1170 17095 -1165
rect 17145 -1145 17175 -1140
rect 17145 -1165 17150 -1145
rect 17150 -1165 17170 -1145
rect 17170 -1165 17175 -1145
rect 17145 -1170 17175 -1165
rect 17225 -1145 17255 -1140
rect 17225 -1165 17230 -1145
rect 17230 -1165 17250 -1145
rect 17250 -1165 17255 -1145
rect 17225 -1170 17255 -1165
rect 17305 -1145 17335 -1140
rect 17305 -1165 17310 -1145
rect 17310 -1165 17330 -1145
rect 17330 -1165 17335 -1145
rect 17305 -1170 17335 -1165
rect 17385 -1145 17415 -1140
rect 17385 -1165 17390 -1145
rect 17390 -1165 17410 -1145
rect 17410 -1165 17415 -1145
rect 17385 -1170 17415 -1165
rect 17465 -1145 17495 -1140
rect 17465 -1165 17470 -1145
rect 17470 -1165 17490 -1145
rect 17490 -1165 17495 -1145
rect 17465 -1170 17495 -1165
rect 17545 -1145 17575 -1140
rect 17545 -1165 17550 -1145
rect 17550 -1165 17570 -1145
rect 17570 -1165 17575 -1145
rect 17545 -1170 17575 -1165
rect 17625 -1145 17655 -1140
rect 17625 -1165 17630 -1145
rect 17630 -1165 17650 -1145
rect 17650 -1165 17655 -1145
rect 17625 -1170 17655 -1165
rect 17705 -1145 17735 -1140
rect 17705 -1165 17710 -1145
rect 17710 -1165 17730 -1145
rect 17730 -1165 17735 -1145
rect 17705 -1170 17735 -1165
rect 17785 -1145 17815 -1140
rect 17785 -1165 17790 -1145
rect 17790 -1165 17810 -1145
rect 17810 -1165 17815 -1145
rect 17785 -1170 17815 -1165
rect 17865 -1145 17895 -1140
rect 17865 -1165 17870 -1145
rect 17870 -1165 17890 -1145
rect 17890 -1165 17895 -1145
rect 17865 -1170 17895 -1165
rect 17945 -1145 17975 -1140
rect 17945 -1165 17950 -1145
rect 17950 -1165 17970 -1145
rect 17970 -1165 17975 -1145
rect 17945 -1170 17975 -1165
rect 18025 -1145 18055 -1140
rect 18025 -1165 18030 -1145
rect 18030 -1165 18050 -1145
rect 18050 -1165 18055 -1145
rect 18025 -1170 18055 -1165
rect 18105 -1145 18135 -1140
rect 18105 -1165 18110 -1145
rect 18110 -1165 18130 -1145
rect 18130 -1165 18135 -1145
rect 18105 -1170 18135 -1165
rect 18185 -1145 18215 -1140
rect 18185 -1165 18190 -1145
rect 18190 -1165 18210 -1145
rect 18210 -1165 18215 -1145
rect 18185 -1170 18215 -1165
rect 18265 -1145 18295 -1140
rect 18265 -1165 18270 -1145
rect 18270 -1165 18290 -1145
rect 18290 -1165 18295 -1145
rect 18265 -1170 18295 -1165
rect 18345 -1145 18375 -1140
rect 18345 -1165 18350 -1145
rect 18350 -1165 18370 -1145
rect 18370 -1165 18375 -1145
rect 18345 -1170 18375 -1165
rect 18425 -1145 18455 -1140
rect 18425 -1165 18430 -1145
rect 18430 -1165 18450 -1145
rect 18450 -1165 18455 -1145
rect 18425 -1170 18455 -1165
rect 18505 -1145 18535 -1140
rect 18505 -1165 18510 -1145
rect 18510 -1165 18530 -1145
rect 18530 -1165 18535 -1145
rect 18505 -1170 18535 -1165
rect 18585 -1145 18615 -1140
rect 18585 -1165 18590 -1145
rect 18590 -1165 18610 -1145
rect 18610 -1165 18615 -1145
rect 18585 -1170 18615 -1165
rect 18665 -1145 18695 -1140
rect 18665 -1165 18670 -1145
rect 18670 -1165 18690 -1145
rect 18690 -1165 18695 -1145
rect 18665 -1170 18695 -1165
rect 18745 -1145 18775 -1140
rect 18745 -1165 18750 -1145
rect 18750 -1165 18770 -1145
rect 18770 -1165 18775 -1145
rect 18745 -1170 18775 -1165
rect 16705 -1230 16735 -1225
rect 16705 -1250 16710 -1230
rect 16710 -1250 16730 -1230
rect 16730 -1250 16735 -1230
rect 16705 -1255 16735 -1250
rect 18900 -1230 18930 -1225
rect 18900 -1250 18905 -1230
rect 18905 -1250 18925 -1230
rect 18925 -1250 18930 -1230
rect 18900 -1255 18930 -1250
rect 16600 -1355 16630 -1325
rect 16710 -1355 16740 -1325
rect 17305 -1355 17335 -1325
rect 17785 -1355 17815 -1325
rect 18265 -1355 18295 -1325
rect 16545 -1440 16575 -1410
rect 16545 -1480 16575 -1450
rect 16655 -1440 16685 -1410
rect 16655 -1480 16685 -1450
rect 16545 -1495 16575 -1490
rect 16545 -1515 16550 -1495
rect 16550 -1515 16570 -1495
rect 16570 -1515 16575 -1495
rect 16545 -1520 16575 -1515
rect 16765 -1440 16795 -1410
rect 16765 -1480 16795 -1450
rect 16655 -1495 16685 -1490
rect 16655 -1515 16660 -1495
rect 16660 -1515 16680 -1495
rect 16680 -1515 16685 -1495
rect 16655 -1520 16685 -1515
rect 16765 -1495 16795 -1490
rect 16765 -1515 16770 -1495
rect 16770 -1515 16790 -1495
rect 16790 -1515 16795 -1495
rect 16765 -1520 16795 -1515
rect 16825 -1440 16855 -1410
rect 16825 -1480 16855 -1450
rect 16825 -1495 16855 -1490
rect 16825 -1515 16830 -1495
rect 16830 -1515 16850 -1495
rect 16850 -1515 16855 -1495
rect 16825 -1520 16855 -1515
rect 17030 -1440 17060 -1410
rect 17030 -1480 17060 -1450
rect 17030 -1495 17060 -1490
rect 17030 -1515 17035 -1495
rect 17035 -1515 17055 -1495
rect 17055 -1515 17060 -1495
rect 17030 -1520 17060 -1515
rect 17140 -1440 17170 -1410
rect 17140 -1480 17170 -1450
rect 17140 -1495 17170 -1490
rect 17140 -1515 17145 -1495
rect 17145 -1515 17165 -1495
rect 17165 -1515 17170 -1495
rect 17140 -1520 17170 -1515
rect 17250 -1440 17280 -1410
rect 17250 -1480 17280 -1450
rect 17360 -1440 17390 -1410
rect 17360 -1480 17390 -1450
rect 17250 -1495 17280 -1490
rect 17250 -1515 17255 -1495
rect 17255 -1515 17275 -1495
rect 17275 -1515 17280 -1495
rect 17250 -1520 17280 -1515
rect 17360 -1495 17390 -1490
rect 17360 -1515 17365 -1495
rect 17365 -1515 17385 -1495
rect 17385 -1515 17390 -1495
rect 17360 -1520 17390 -1515
rect 17470 -1440 17500 -1410
rect 17470 -1480 17500 -1450
rect 17470 -1495 17500 -1490
rect 17470 -1515 17475 -1495
rect 17475 -1515 17495 -1495
rect 17495 -1515 17500 -1495
rect 17470 -1520 17500 -1515
rect 17620 -1440 17650 -1410
rect 17620 -1480 17650 -1450
rect 17620 -1495 17650 -1490
rect 17620 -1515 17625 -1495
rect 17625 -1515 17645 -1495
rect 17645 -1515 17650 -1495
rect 17620 -1520 17650 -1515
rect 17730 -1440 17760 -1410
rect 17730 -1480 17760 -1450
rect 17840 -1440 17870 -1410
rect 17840 -1480 17870 -1450
rect 17730 -1495 17760 -1490
rect 17730 -1515 17735 -1495
rect 17735 -1515 17755 -1495
rect 17755 -1515 17760 -1495
rect 17730 -1520 17760 -1515
rect 17840 -1495 17870 -1490
rect 17840 -1515 17845 -1495
rect 17845 -1515 17865 -1495
rect 17865 -1515 17870 -1495
rect 17840 -1520 17870 -1515
rect 17950 -1440 17980 -1410
rect 17950 -1480 17980 -1450
rect 17950 -1495 17980 -1490
rect 17950 -1515 17955 -1495
rect 17955 -1515 17975 -1495
rect 17975 -1515 17980 -1495
rect 17950 -1520 17980 -1515
rect 18100 -1440 18130 -1410
rect 18100 -1480 18130 -1450
rect 18100 -1495 18130 -1490
rect 18100 -1515 18105 -1495
rect 18105 -1515 18125 -1495
rect 18125 -1515 18130 -1495
rect 18100 -1520 18130 -1515
rect 18210 -1440 18240 -1410
rect 18210 -1480 18240 -1450
rect 18320 -1440 18350 -1410
rect 18320 -1480 18350 -1450
rect 18210 -1495 18240 -1490
rect 18210 -1515 18215 -1495
rect 18215 -1515 18235 -1495
rect 18235 -1515 18240 -1495
rect 18210 -1520 18240 -1515
rect 18320 -1495 18350 -1490
rect 18320 -1515 18325 -1495
rect 18325 -1515 18345 -1495
rect 18345 -1515 18350 -1495
rect 18320 -1520 18350 -1515
rect 18430 -1440 18460 -1410
rect 18430 -1480 18460 -1450
rect 18430 -1495 18460 -1490
rect 18430 -1515 18435 -1495
rect 18435 -1515 18455 -1495
rect 18455 -1515 18460 -1495
rect 18430 -1520 18460 -1515
rect 18540 -1440 18570 -1410
rect 18540 -1480 18570 -1450
rect 18540 -1495 18570 -1490
rect 18540 -1515 18545 -1495
rect 18545 -1515 18565 -1495
rect 18565 -1515 18570 -1495
rect 18540 -1520 18570 -1515
rect 17195 -1665 17225 -1660
rect 17195 -1685 17200 -1665
rect 17200 -1685 17220 -1665
rect 17220 -1685 17225 -1665
rect 17195 -1690 17225 -1685
rect 17085 -1745 17115 -1715
rect 17415 -1665 17445 -1660
rect 17415 -1685 17420 -1665
rect 17420 -1685 17440 -1665
rect 17440 -1685 17445 -1665
rect 17415 -1690 17445 -1685
rect 17675 -1665 17705 -1660
rect 17675 -1685 17680 -1665
rect 17680 -1685 17700 -1665
rect 17700 -1685 17705 -1665
rect 17675 -1690 17705 -1685
rect 17785 -1665 17815 -1660
rect 17785 -1685 17790 -1665
rect 17790 -1685 17810 -1665
rect 17810 -1685 17815 -1665
rect 17785 -1690 17815 -1685
rect 17895 -1665 17925 -1660
rect 17895 -1685 17900 -1665
rect 17900 -1685 17920 -1665
rect 17920 -1685 17925 -1665
rect 17895 -1690 17925 -1685
rect 18155 -1665 18185 -1660
rect 18155 -1685 18160 -1665
rect 18160 -1685 18180 -1665
rect 18180 -1685 18185 -1665
rect 18155 -1690 18185 -1685
rect 18375 -1665 18405 -1660
rect 18375 -1685 18380 -1665
rect 18380 -1685 18400 -1665
rect 18400 -1685 18405 -1665
rect 18375 -1690 18405 -1685
rect 17305 -1745 17335 -1715
rect 17195 -1800 17225 -1770
rect 17195 -1840 17225 -1810
rect 18265 -1745 18295 -1715
rect 18485 -1745 18515 -1715
rect 18375 -1800 18405 -1770
rect 18375 -1840 18405 -1810
rect 16710 -1930 16740 -1900
rect 17785 -1930 17815 -1900
rect 19330 -1980 19360 -1950
rect 16265 -2030 16295 -2000
rect 16485 -2030 16515 -2000
rect 16735 -2030 16765 -2000
rect 17200 -2030 17230 -2000
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16160 -3030 16195 -3025
rect 16160 -3055 16165 -3030
rect 16165 -3055 16190 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3060 16195 -3055
rect 17430 -2005 17465 -2000
rect 17430 -2030 17435 -2005
rect 17435 -2030 17460 -2005
rect 17460 -2030 17465 -2005
rect 17430 -2035 17465 -2030
rect 18129 -2005 18164 -2000
rect 18129 -2030 18134 -2005
rect 18134 -2030 18159 -2005
rect 18159 -2030 18164 -2005
rect 18129 -2035 18164 -2030
rect 19085 -2035 19115 -2005
rect 17200 -2090 17230 -2060
rect 18835 -2090 18865 -2060
rect 15825 -3145 15855 -3115
rect 15950 -3121 15985 -3116
rect 15950 -3146 15955 -3121
rect 15955 -3146 15980 -3121
rect 15980 -3146 15985 -3121
rect 16735 -3135 16765 -3105
rect 15950 -3151 15985 -3146
rect 17785 -3135 17815 -3105
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19615 220 19645 250
rect 19540 -1930 19570 -1900
rect 19465 -2035 19495 -2005
rect 19405 -3002 19440 -2997
rect 19405 -3027 19410 -3002
rect 19410 -3027 19435 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3032 19440 -3027
rect 18620 -3135 18650 -3105
rect 18835 -3135 18865 -3105
rect 19725 -285 19755 -255
rect 19610 -3121 19645 -3116
rect 19610 -3146 19615 -3121
rect 19615 -3146 19640 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3151 19645 -3146
rect 15950 -3794 15985 -3789
rect 15950 -3819 15955 -3794
rect 15955 -3819 15980 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3824 15985 -3819
rect 15825 -4295 15855 -4265
rect 15730 -4345 15760 -4315
rect 16280 -3899 16315 -3894
rect 16280 -3924 16285 -3899
rect 16285 -3924 16310 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3929 16315 -3924
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 19610 -3794 19645 -3789
rect 19610 -3819 19615 -3794
rect 19615 -3819 19640 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3824 19645 -3819
rect 19285 -3899 19320 -3894
rect 19285 -3924 19290 -3899
rect 19290 -3924 19315 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3929 19320 -3924
rect 18960 -3974 18995 -3969
rect 16605 -4004 16640 -3999
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 16285 -4220 16315 -4190
rect 16610 -4220 16640 -4190
rect 17260 -4295 17290 -4265
rect 17785 -4270 17815 -4265
rect 17785 -4290 17790 -4270
rect 17790 -4290 17810 -4270
rect 17810 -4290 17815 -4270
rect 17785 -4295 17815 -4290
rect 18960 -4295 18990 -4265
rect 19285 -4295 19315 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 19780 -1800 19810 -1770
rect 19780 -1840 19810 -1810
rect 19725 -4345 19755 -4315
rect 15955 -4390 15985 -4360
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 19615 -4390 19645 -4360
rect 17960 -4440 17990 -4410
<< metal2 >>
rect 16940 1505 16980 1510
rect 16940 1475 16945 1505
rect 16975 1475 16980 1505
rect 16940 1470 16980 1475
rect 18620 1505 18660 1510
rect 18620 1475 18625 1505
rect 18655 1475 18660 1505
rect 18620 1470 18660 1475
rect 16485 1460 16525 1465
rect 16485 1430 16490 1460
rect 16520 1455 16525 1460
rect 17050 1460 17090 1465
rect 17050 1455 17055 1460
rect 16520 1435 17055 1455
rect 16520 1430 16525 1435
rect 16485 1425 16525 1430
rect 17050 1430 17055 1435
rect 17085 1455 17090 1460
rect 17780 1460 17820 1465
rect 17780 1455 17785 1460
rect 17085 1435 17785 1455
rect 17085 1430 17090 1435
rect 17050 1425 17090 1430
rect 17780 1430 17785 1435
rect 17815 1455 17820 1460
rect 18200 1460 18240 1465
rect 18200 1455 18205 1460
rect 17815 1435 18205 1455
rect 17815 1430 17820 1435
rect 17780 1425 17820 1430
rect 18200 1430 18205 1435
rect 18235 1455 18240 1460
rect 18510 1460 18550 1465
rect 18510 1455 18515 1460
rect 18235 1435 18515 1455
rect 18235 1430 18240 1435
rect 18200 1425 18240 1430
rect 18510 1430 18515 1435
rect 18545 1430 18550 1460
rect 18510 1425 18550 1430
rect 16365 1360 18715 1365
rect 16365 1330 16370 1360
rect 16400 1330 16490 1360
rect 16520 1330 16610 1360
rect 16640 1330 16890 1360
rect 16920 1330 17000 1360
rect 17030 1330 17110 1360
rect 17140 1330 17220 1360
rect 17250 1330 17500 1360
rect 17530 1330 17565 1360
rect 17595 1330 17675 1360
rect 17705 1330 17785 1360
rect 17815 1330 17895 1360
rect 17925 1330 18005 1360
rect 18035 1330 18070 1360
rect 18100 1330 18350 1360
rect 18380 1330 18460 1360
rect 18490 1330 18570 1360
rect 18600 1330 18680 1360
rect 18710 1330 18715 1360
rect 16365 1320 18715 1330
rect 16365 1290 16370 1320
rect 16400 1290 16490 1320
rect 16520 1290 16610 1320
rect 16640 1290 16890 1320
rect 16920 1290 17000 1320
rect 17030 1290 17110 1320
rect 17140 1290 17220 1320
rect 17250 1290 17500 1320
rect 17530 1290 17565 1320
rect 17595 1290 17675 1320
rect 17705 1290 17785 1320
rect 17815 1290 17895 1320
rect 17925 1290 18005 1320
rect 18035 1290 18070 1320
rect 18100 1290 18350 1320
rect 18380 1290 18460 1320
rect 18490 1290 18570 1320
rect 18600 1290 18680 1320
rect 18710 1290 18715 1320
rect 16365 1280 18715 1290
rect 16365 1250 16370 1280
rect 16400 1250 16490 1280
rect 16520 1250 16610 1280
rect 16640 1250 16890 1280
rect 16920 1250 17000 1280
rect 17030 1250 17110 1280
rect 17140 1250 17220 1280
rect 17250 1250 17500 1280
rect 17530 1250 17565 1280
rect 17595 1250 17675 1280
rect 17705 1250 17785 1280
rect 17815 1250 17895 1280
rect 17925 1250 18005 1280
rect 18035 1250 18070 1280
rect 18100 1250 18350 1280
rect 18380 1250 18460 1280
rect 18490 1250 18570 1280
rect 18600 1250 18680 1280
rect 18710 1250 18715 1280
rect 16365 1245 18715 1250
rect 16430 1110 16470 1115
rect 16430 1080 16435 1110
rect 16465 1080 16470 1110
rect 16430 1075 16470 1080
rect 16540 1110 16580 1115
rect 16540 1080 16545 1110
rect 16575 1080 16580 1110
rect 16540 1075 16580 1080
rect 16940 1110 16980 1115
rect 16940 1080 16945 1110
rect 16975 1105 16980 1110
rect 17050 1110 17090 1115
rect 17050 1105 17055 1110
rect 16975 1085 17055 1105
rect 16975 1080 16980 1085
rect 16940 1075 16980 1080
rect 17050 1080 17055 1085
rect 17085 1105 17090 1110
rect 17160 1110 17200 1115
rect 17160 1105 17165 1110
rect 17085 1085 17165 1105
rect 17085 1080 17090 1085
rect 17050 1075 17090 1080
rect 17160 1080 17165 1085
rect 17195 1080 17200 1110
rect 17160 1075 17200 1080
rect 17615 1110 17655 1115
rect 17615 1080 17620 1110
rect 17650 1105 17655 1110
rect 17725 1110 17765 1115
rect 17725 1105 17730 1110
rect 17650 1085 17730 1105
rect 17650 1080 17655 1085
rect 17615 1075 17655 1080
rect 17725 1080 17730 1085
rect 17760 1105 17765 1110
rect 17835 1110 17875 1115
rect 17835 1105 17840 1110
rect 17760 1085 17840 1105
rect 17760 1080 17765 1085
rect 17725 1075 17765 1080
rect 17835 1080 17840 1085
rect 17870 1105 17875 1110
rect 17945 1110 17985 1115
rect 17945 1105 17950 1110
rect 17870 1085 17950 1105
rect 17870 1080 17875 1085
rect 17835 1075 17875 1080
rect 17945 1080 17950 1085
rect 17980 1080 17985 1110
rect 17945 1075 17985 1080
rect 18400 1110 18440 1115
rect 18400 1080 18405 1110
rect 18435 1105 18440 1110
rect 18510 1110 18550 1115
rect 18510 1105 18515 1110
rect 18435 1085 18515 1105
rect 18435 1080 18440 1085
rect 18400 1075 18440 1080
rect 18510 1080 18515 1085
rect 18545 1105 18550 1110
rect 18620 1110 18660 1115
rect 18620 1105 18625 1110
rect 18545 1085 18625 1105
rect 18545 1080 18550 1085
rect 18510 1075 18550 1080
rect 18620 1080 18625 1085
rect 18655 1080 18660 1110
rect 18620 1075 18660 1080
rect 18200 1055 18240 1060
rect 18200 1025 18205 1055
rect 18235 1050 18240 1055
rect 18720 1055 18760 1060
rect 18720 1050 18725 1055
rect 18235 1030 18725 1050
rect 18235 1025 18240 1030
rect 18200 1020 18240 1025
rect 18720 1025 18725 1030
rect 18755 1025 18760 1055
rect 18720 1020 18760 1025
rect 16160 1010 16200 1015
rect 16160 980 16165 1010
rect 16195 1005 16200 1010
rect 16430 1010 16470 1015
rect 16430 1005 16435 1010
rect 16195 985 16435 1005
rect 16195 980 16200 985
rect 16160 975 16200 980
rect 16430 980 16435 985
rect 16465 980 16470 1010
rect 16430 975 16470 980
rect 16540 1010 16580 1015
rect 16540 980 16545 1010
rect 16575 1005 16580 1010
rect 19325 1010 19365 1015
rect 19325 1005 19330 1010
rect 16575 985 19330 1005
rect 16575 980 16580 985
rect 16540 975 16580 980
rect 19325 980 19330 985
rect 19360 980 19365 1010
rect 19325 975 19365 980
rect 16435 935 19115 940
rect 16435 905 16440 935
rect 16470 905 16660 935
rect 16690 905 16975 935
rect 17005 905 17155 935
rect 17185 905 17335 935
rect 17365 905 17515 935
rect 17545 905 17695 935
rect 17725 905 17875 935
rect 17905 905 18055 935
rect 18085 905 18235 935
rect 18265 905 18415 935
rect 18445 905 18595 935
rect 18625 905 18910 935
rect 18940 905 19020 935
rect 19050 905 19080 935
rect 19110 905 19115 935
rect 16435 895 19115 905
rect 16435 865 16440 895
rect 16470 865 16660 895
rect 16690 865 16975 895
rect 17005 865 17155 895
rect 17185 865 17335 895
rect 17365 865 17515 895
rect 17545 865 17695 895
rect 17725 865 17875 895
rect 17905 865 18055 895
rect 18085 865 18235 895
rect 18265 865 18415 895
rect 18445 865 18595 895
rect 18625 865 18910 895
rect 18940 865 19020 895
rect 19050 865 19080 895
rect 19110 865 19115 895
rect 16435 855 19115 865
rect 16435 825 16440 855
rect 16470 825 16660 855
rect 16690 825 16975 855
rect 17005 825 17155 855
rect 17185 825 17335 855
rect 17365 825 17515 855
rect 17545 825 17695 855
rect 17725 825 17875 855
rect 17905 825 18055 855
rect 18085 825 18235 855
rect 18265 825 18415 855
rect 18445 825 18595 855
rect 18625 825 18910 855
rect 18940 825 19020 855
rect 19050 825 19080 855
rect 19110 825 19115 855
rect 16435 815 19115 825
rect 16435 785 16440 815
rect 16470 785 16660 815
rect 16690 785 16975 815
rect 17005 785 17155 815
rect 17185 785 17335 815
rect 17365 785 17515 815
rect 17545 785 17695 815
rect 17725 785 17875 815
rect 17905 785 18055 815
rect 18085 785 18235 815
rect 18265 785 18415 815
rect 18445 785 18595 815
rect 18625 785 18910 815
rect 18940 785 19020 815
rect 19050 785 19080 815
rect 19110 785 19115 815
rect 16435 780 19115 785
rect 16545 715 16585 720
rect 16545 685 16550 715
rect 16580 710 16585 715
rect 16780 715 16820 720
rect 16780 710 16785 715
rect 16580 690 16785 710
rect 16580 685 16585 690
rect 16545 680 16585 685
rect 16780 685 16785 690
rect 16815 685 16820 715
rect 16780 680 16820 685
rect 16480 545 16520 550
rect 16480 515 16485 545
rect 16515 540 16520 545
rect 16610 545 16650 550
rect 16610 540 16615 545
rect 16515 520 16615 540
rect 16515 515 16520 520
rect 16480 510 16520 515
rect 16610 515 16615 520
rect 16645 540 16650 545
rect 16840 545 16880 550
rect 16840 540 16845 545
rect 16645 520 16845 540
rect 16645 515 16650 520
rect 16610 510 16650 515
rect 16840 515 16845 520
rect 16875 515 16880 545
rect 16840 510 16880 515
rect 18950 545 18990 550
rect 18950 515 18955 545
rect 18985 540 18990 545
rect 19260 545 19300 550
rect 19260 540 19265 545
rect 18985 520 19265 540
rect 18985 515 18990 520
rect 18950 510 18990 515
rect 19260 515 19265 520
rect 19295 515 19300 545
rect 19260 510 19300 515
rect 19000 465 19005 495
rect 19035 465 19040 495
rect 16315 445 19500 450
rect 16315 415 16320 445
rect 16350 415 17605 445
rect 17635 415 17965 445
rect 17995 415 19465 445
rect 19495 415 19500 445
rect 16315 410 19500 415
rect 16260 390 16300 395
rect 16260 360 16265 390
rect 16295 385 16300 390
rect 16780 390 16820 395
rect 16780 385 16785 390
rect 16295 365 16785 385
rect 16295 360 16300 365
rect 16260 355 16300 360
rect 16780 360 16785 365
rect 16815 385 16820 390
rect 17420 390 17460 395
rect 17420 385 17425 390
rect 16815 365 17425 385
rect 16815 360 16820 365
rect 16780 355 16820 360
rect 17420 360 17425 365
rect 17455 385 17460 390
rect 18140 390 18180 395
rect 18140 385 18145 390
rect 17455 365 18145 385
rect 17455 360 17460 365
rect 17420 355 17460 360
rect 18140 360 18145 365
rect 18175 360 18180 390
rect 18140 355 18180 360
rect 16205 345 16245 350
rect 16205 315 16210 345
rect 16240 340 16245 345
rect 16545 345 16585 350
rect 16545 340 16550 345
rect 16240 320 16550 340
rect 16240 315 16245 320
rect 16205 310 16245 315
rect 16545 315 16550 320
rect 16580 340 16585 345
rect 17240 345 17280 350
rect 17240 340 17245 345
rect 16580 320 17245 340
rect 16580 315 16585 320
rect 16545 310 16585 315
rect 17240 315 17245 320
rect 17275 340 17280 345
rect 18320 345 18360 350
rect 18320 340 18325 345
rect 17275 320 18325 340
rect 17275 315 17280 320
rect 17240 310 17280 315
rect 18320 315 18325 320
rect 18355 315 18360 345
rect 18320 310 18360 315
rect 17060 300 17100 305
rect 17060 270 17065 300
rect 17095 295 17100 300
rect 17780 300 17820 305
rect 17780 295 17785 300
rect 17095 275 17785 295
rect 17095 270 17100 275
rect 17060 265 17100 270
rect 17780 270 17785 275
rect 17815 295 17820 300
rect 18500 300 18540 305
rect 18500 295 18505 300
rect 17815 275 18505 295
rect 17815 270 17820 275
rect 17780 265 17820 270
rect 18500 270 18505 275
rect 18535 295 18540 300
rect 19405 300 19445 305
rect 19405 295 19410 300
rect 18535 275 19410 295
rect 18535 270 18540 275
rect 18500 265 18540 270
rect 19405 270 19410 275
rect 19440 270 19445 300
rect 19405 265 19445 270
rect 18000 250 18040 255
rect 18000 220 18005 250
rect 18035 245 18040 250
rect 18720 250 18760 255
rect 18720 245 18725 250
rect 18035 225 18725 245
rect 18035 220 18040 225
rect 18000 215 18040 220
rect 18720 220 18725 225
rect 18755 245 18760 250
rect 19010 250 19050 255
rect 19010 245 19015 250
rect 18755 225 19015 245
rect 18755 220 18760 225
rect 18720 215 18760 220
rect 19010 220 19015 225
rect 19045 245 19050 250
rect 19610 250 19650 255
rect 19610 245 19615 250
rect 19045 225 19615 245
rect 19045 220 19050 225
rect 19010 215 19050 220
rect 19610 220 19615 225
rect 19645 220 19650 250
rect 19610 215 19650 220
rect 16420 110 19180 115
rect 16420 80 16425 110
rect 16455 80 16545 110
rect 16575 80 16665 110
rect 16695 80 16785 110
rect 16815 80 16905 110
rect 16935 80 17025 110
rect 17055 80 17145 110
rect 17175 80 17265 110
rect 17295 80 17385 110
rect 17415 80 17505 110
rect 17535 80 17625 110
rect 17655 80 17945 110
rect 17975 80 18065 110
rect 18095 80 18185 110
rect 18215 80 18305 110
rect 18335 80 18425 110
rect 18455 80 18545 110
rect 18575 80 18665 110
rect 18695 80 18785 110
rect 18815 80 18905 110
rect 18935 80 19025 110
rect 19055 80 19145 110
rect 19175 80 19180 110
rect 16420 70 19180 80
rect 16420 40 16425 70
rect 16455 40 16545 70
rect 16575 40 16665 70
rect 16695 40 16785 70
rect 16815 40 16905 70
rect 16935 40 17025 70
rect 17055 40 17145 70
rect 17175 40 17265 70
rect 17295 40 17385 70
rect 17415 40 17505 70
rect 17535 40 17625 70
rect 17655 40 17945 70
rect 17975 40 18065 70
rect 18095 40 18185 70
rect 18215 40 18305 70
rect 18335 40 18425 70
rect 18455 40 18545 70
rect 18575 40 18665 70
rect 18695 40 18785 70
rect 18815 40 18905 70
rect 18935 40 19025 70
rect 19055 40 19145 70
rect 19175 40 19180 70
rect 16420 30 19180 40
rect 16420 0 16425 30
rect 16455 0 16545 30
rect 16575 0 16665 30
rect 16695 0 16785 30
rect 16815 0 16905 30
rect 16935 0 17025 30
rect 17055 0 17145 30
rect 17175 0 17265 30
rect 17295 0 17385 30
rect 17415 0 17505 30
rect 17535 0 17625 30
rect 17655 0 17945 30
rect 17975 0 18065 30
rect 18095 0 18185 30
rect 18215 0 18305 30
rect 18335 0 18425 30
rect 18455 0 18545 30
rect 18575 0 18665 30
rect 18695 0 18785 30
rect 18815 0 18905 30
rect 18935 0 19025 30
rect 19055 0 19145 30
rect 19175 0 19180 30
rect 16420 -5 19180 0
rect 15950 -25 15990 -20
rect 15950 -55 15955 -25
rect 15985 -30 15990 -25
rect 16480 -25 16520 -20
rect 16480 -30 16485 -25
rect 15985 -50 16485 -30
rect 15985 -55 15990 -50
rect 15950 -60 15990 -55
rect 16480 -55 16485 -50
rect 16515 -30 16520 -25
rect 16840 -25 16880 -20
rect 16840 -30 16845 -25
rect 16515 -50 16845 -30
rect 16515 -55 16520 -50
rect 16480 -60 16520 -55
rect 16840 -55 16845 -50
rect 16875 -30 16880 -25
rect 17200 -25 17240 -20
rect 17200 -30 17205 -25
rect 16875 -50 17205 -30
rect 16875 -55 16880 -50
rect 16840 -60 16880 -55
rect 17200 -55 17205 -50
rect 17235 -30 17240 -25
rect 17560 -25 17600 -20
rect 17560 -30 17565 -25
rect 17235 -50 17565 -30
rect 17235 -55 17240 -50
rect 17200 -60 17240 -55
rect 17560 -55 17565 -50
rect 17595 -30 17600 -25
rect 17690 -25 17730 -20
rect 17690 -30 17695 -25
rect 17595 -50 17695 -30
rect 17595 -55 17600 -50
rect 17560 -60 17600 -55
rect 17690 -55 17695 -50
rect 17725 -55 17730 -25
rect 17690 -60 17730 -55
rect 17870 -25 17910 -20
rect 17870 -55 17875 -25
rect 17905 -30 17910 -25
rect 18000 -25 18040 -20
rect 18000 -30 18005 -25
rect 17905 -50 18005 -30
rect 17905 -55 17910 -50
rect 17870 -60 17910 -55
rect 18000 -55 18005 -50
rect 18035 -30 18040 -25
rect 18360 -25 18400 -20
rect 18360 -30 18365 -25
rect 18035 -50 18365 -30
rect 18035 -55 18040 -50
rect 18000 -60 18040 -55
rect 18360 -55 18365 -50
rect 18395 -30 18400 -25
rect 18720 -25 18760 -20
rect 18720 -30 18725 -25
rect 18395 -50 18725 -30
rect 18395 -55 18400 -50
rect 18360 -60 18400 -55
rect 18720 -55 18725 -50
rect 18755 -30 18760 -25
rect 19080 -25 19120 -20
rect 19080 -30 19085 -25
rect 18755 -50 19085 -30
rect 18755 -55 18760 -50
rect 18720 -60 18760 -55
rect 19080 -55 19085 -50
rect 19115 -55 19120 -25
rect 19080 -60 19120 -55
rect 16600 -195 16640 -190
rect 16600 -225 16605 -195
rect 16635 -200 16640 -195
rect 16960 -195 17000 -190
rect 16960 -200 16965 -195
rect 16635 -220 16965 -200
rect 16635 -225 16640 -220
rect 16600 -230 16640 -225
rect 16960 -225 16965 -220
rect 16995 -200 17000 -195
rect 17320 -195 17360 -190
rect 17320 -200 17325 -195
rect 16995 -220 17325 -200
rect 16995 -225 17000 -220
rect 16960 -230 17000 -225
rect 17320 -225 17325 -220
rect 17355 -225 17360 -195
rect 17320 -230 17360 -225
rect 18240 -195 18280 -190
rect 18240 -225 18245 -195
rect 18275 -200 18280 -195
rect 18600 -195 18640 -190
rect 18600 -200 18605 -195
rect 18275 -220 18605 -200
rect 18275 -225 18280 -220
rect 18240 -230 18280 -225
rect 18600 -225 18605 -220
rect 18635 -200 18640 -195
rect 18960 -195 19000 -190
rect 18960 -200 18965 -195
rect 18635 -220 18965 -200
rect 18635 -225 18640 -220
rect 18600 -230 18640 -225
rect 18960 -225 18965 -220
rect 18995 -225 19000 -195
rect 18960 -230 19000 -225
rect 15725 -255 15765 -250
rect 15725 -285 15730 -255
rect 15760 -260 15765 -255
rect 16510 -255 16550 -250
rect 16510 -260 16515 -255
rect 15760 -280 16515 -260
rect 15760 -285 15765 -280
rect 15725 -290 15765 -285
rect 16510 -285 16515 -280
rect 16545 -260 16550 -255
rect 16720 -255 16760 -250
rect 16720 -260 16725 -255
rect 16545 -280 16725 -260
rect 16545 -285 16550 -280
rect 16510 -290 16550 -285
rect 16720 -285 16725 -280
rect 16755 -260 16760 -255
rect 16840 -255 16880 -250
rect 16840 -260 16845 -255
rect 16755 -280 16845 -260
rect 16755 -285 16760 -280
rect 16720 -290 16760 -285
rect 16840 -285 16845 -280
rect 16875 -260 16880 -255
rect 17080 -255 17120 -250
rect 17080 -260 17085 -255
rect 16875 -280 17085 -260
rect 16875 -285 16880 -280
rect 16840 -290 16880 -285
rect 17080 -285 17085 -280
rect 17115 -260 17120 -255
rect 17200 -255 17240 -250
rect 17200 -260 17205 -255
rect 17115 -280 17205 -260
rect 17115 -285 17120 -280
rect 17080 -290 17120 -285
rect 17200 -285 17205 -280
rect 17235 -260 17240 -255
rect 17440 -255 17480 -250
rect 17440 -260 17445 -255
rect 17235 -280 17445 -260
rect 17235 -285 17240 -280
rect 17200 -290 17240 -285
rect 17440 -285 17445 -280
rect 17475 -260 17480 -255
rect 17530 -255 17570 -250
rect 17530 -260 17535 -255
rect 17475 -280 17535 -260
rect 17475 -285 17480 -280
rect 17440 -290 17480 -285
rect 17530 -285 17535 -280
rect 17565 -285 17570 -255
rect 17530 -290 17570 -285
rect 18030 -255 18070 -250
rect 18030 -285 18035 -255
rect 18065 -260 18070 -255
rect 18120 -255 18160 -250
rect 18120 -260 18125 -255
rect 18065 -280 18125 -260
rect 18065 -285 18070 -280
rect 18030 -290 18070 -285
rect 18120 -285 18125 -280
rect 18155 -260 18160 -255
rect 18360 -255 18400 -250
rect 18360 -260 18365 -255
rect 18155 -280 18365 -260
rect 18155 -285 18160 -280
rect 18120 -290 18160 -285
rect 18360 -285 18365 -280
rect 18395 -260 18400 -255
rect 18480 -255 18520 -250
rect 18480 -260 18485 -255
rect 18395 -280 18485 -260
rect 18395 -285 18400 -280
rect 18360 -290 18400 -285
rect 18480 -285 18485 -280
rect 18515 -260 18520 -255
rect 18720 -255 18760 -250
rect 18720 -260 18725 -255
rect 18515 -280 18725 -260
rect 18515 -285 18520 -280
rect 18480 -290 18520 -285
rect 18720 -285 18725 -280
rect 18755 -260 18760 -255
rect 18840 -255 18880 -250
rect 18840 -260 18845 -255
rect 18755 -280 18845 -260
rect 18755 -285 18760 -280
rect 18720 -290 18760 -285
rect 18840 -285 18845 -280
rect 18875 -260 18880 -255
rect 19050 -255 19090 -250
rect 19050 -260 19055 -255
rect 18875 -280 19055 -260
rect 18875 -285 18880 -280
rect 18840 -290 18880 -285
rect 19050 -285 19055 -280
rect 19085 -260 19090 -255
rect 19720 -255 19760 -250
rect 19720 -260 19725 -255
rect 19085 -280 19725 -260
rect 19085 -285 19090 -280
rect 19050 -290 19090 -285
rect 19720 -285 19725 -280
rect 19755 -285 19760 -255
rect 19720 -290 19760 -285
rect 16260 -310 16300 -305
rect 16260 -340 16265 -310
rect 16295 -315 16300 -310
rect 17007 -310 17037 -305
rect 16295 -335 17007 -315
rect 16295 -340 16300 -335
rect 16260 -345 16300 -340
rect 18563 -310 18593 -305
rect 18562 -335 18563 -315
rect 17007 -345 17037 -340
rect 19405 -310 19445 -305
rect 19405 -315 19410 -310
rect 18593 -335 19410 -315
rect 18563 -345 18593 -340
rect 19405 -340 19410 -335
rect 19440 -340 19445 -310
rect 19405 -345 19445 -340
rect 17565 -370 17595 -365
rect 17780 -370 17820 -365
rect 17780 -375 17785 -370
rect 17595 -395 17785 -375
rect 17565 -405 17595 -400
rect 17780 -400 17785 -395
rect 17815 -375 17820 -370
rect 18005 -370 18035 -365
rect 17815 -395 18005 -375
rect 17815 -400 17820 -395
rect 17780 -405 17820 -400
rect 18005 -405 18035 -400
rect 16315 -630 17105 -625
rect 16315 -660 16320 -630
rect 16350 -660 17075 -630
rect 16315 -665 17105 -660
rect 18495 -630 18525 -625
rect 19325 -630 19365 -625
rect 19325 -635 19330 -630
rect 18525 -655 19330 -635
rect 18495 -665 18525 -660
rect 19325 -660 19330 -655
rect 19360 -660 19365 -630
rect 19325 -665 19365 -660
rect 16530 -710 17060 -705
rect 16530 -740 16535 -710
rect 16565 -740 17025 -710
rect 17055 -740 17060 -710
rect 16530 -745 17060 -740
rect 18540 -710 18580 -705
rect 18540 -740 18545 -710
rect 18575 -715 18580 -710
rect 19030 -710 19070 -705
rect 19030 -715 19035 -710
rect 18575 -735 19035 -715
rect 18575 -740 18580 -735
rect 18540 -745 18580 -740
rect 19030 -740 19035 -735
rect 19065 -740 19070 -710
rect 19030 -745 19070 -740
rect 16620 -765 18980 -760
rect 16620 -795 16625 -765
rect 16655 -795 16745 -765
rect 16775 -795 16865 -765
rect 16895 -795 16985 -765
rect 17015 -795 17305 -765
rect 17335 -795 17425 -765
rect 17455 -795 17545 -765
rect 17575 -795 18025 -765
rect 18055 -795 18145 -765
rect 18175 -795 18265 -765
rect 18295 -795 18585 -765
rect 18615 -795 18705 -765
rect 18735 -795 18825 -765
rect 18855 -795 18945 -765
rect 18975 -795 18980 -765
rect 16620 -800 18980 -795
rect 17110 -1080 17150 -1075
rect 17110 -1110 17115 -1080
rect 17145 -1085 17150 -1080
rect 17780 -1080 17820 -1075
rect 17780 -1085 17785 -1080
rect 17145 -1105 17785 -1085
rect 17145 -1110 17150 -1105
rect 17110 -1115 17150 -1110
rect 17780 -1110 17785 -1105
rect 17815 -1085 17820 -1080
rect 18450 -1080 18490 -1075
rect 18450 -1085 18455 -1080
rect 17815 -1105 18455 -1085
rect 17815 -1110 17820 -1105
rect 17780 -1115 17820 -1110
rect 18450 -1110 18455 -1105
rect 18485 -1110 18490 -1080
rect 18450 -1115 18490 -1110
rect 16740 -1140 16780 -1135
rect 16740 -1170 16745 -1140
rect 16775 -1145 16780 -1140
rect 16820 -1140 16860 -1135
rect 16820 -1145 16825 -1140
rect 16775 -1165 16825 -1145
rect 16775 -1170 16780 -1165
rect 16740 -1175 16780 -1170
rect 16820 -1170 16825 -1165
rect 16855 -1145 16860 -1140
rect 16900 -1140 16940 -1135
rect 16900 -1145 16905 -1140
rect 16855 -1165 16905 -1145
rect 16855 -1170 16860 -1165
rect 16820 -1175 16860 -1170
rect 16900 -1170 16905 -1165
rect 16935 -1145 16940 -1140
rect 16980 -1140 17020 -1135
rect 16980 -1145 16985 -1140
rect 16935 -1165 16985 -1145
rect 16935 -1170 16940 -1165
rect 16900 -1175 16940 -1170
rect 16980 -1170 16985 -1165
rect 17015 -1145 17020 -1140
rect 17060 -1140 17100 -1135
rect 17060 -1145 17065 -1140
rect 17015 -1165 17065 -1145
rect 17015 -1170 17020 -1165
rect 16980 -1175 17020 -1170
rect 17060 -1170 17065 -1165
rect 17095 -1145 17100 -1140
rect 17140 -1140 17180 -1135
rect 17140 -1145 17145 -1140
rect 17095 -1165 17145 -1145
rect 17095 -1170 17100 -1165
rect 17060 -1175 17100 -1170
rect 17140 -1170 17145 -1165
rect 17175 -1145 17180 -1140
rect 17220 -1140 17260 -1135
rect 17220 -1145 17225 -1140
rect 17175 -1165 17225 -1145
rect 17175 -1170 17180 -1165
rect 17140 -1175 17180 -1170
rect 17220 -1170 17225 -1165
rect 17255 -1145 17260 -1140
rect 17300 -1140 17340 -1135
rect 17300 -1145 17305 -1140
rect 17255 -1165 17305 -1145
rect 17255 -1170 17260 -1165
rect 17220 -1175 17260 -1170
rect 17300 -1170 17305 -1165
rect 17335 -1145 17340 -1140
rect 17380 -1140 17420 -1135
rect 17380 -1145 17385 -1140
rect 17335 -1165 17385 -1145
rect 17335 -1170 17340 -1165
rect 17300 -1175 17340 -1170
rect 17380 -1170 17385 -1165
rect 17415 -1145 17420 -1140
rect 17460 -1140 17500 -1135
rect 17460 -1145 17465 -1140
rect 17415 -1165 17465 -1145
rect 17415 -1170 17420 -1165
rect 17380 -1175 17420 -1170
rect 17460 -1170 17465 -1165
rect 17495 -1145 17500 -1140
rect 17540 -1140 17580 -1135
rect 17540 -1145 17545 -1140
rect 17495 -1165 17545 -1145
rect 17495 -1170 17500 -1165
rect 17460 -1175 17500 -1170
rect 17540 -1170 17545 -1165
rect 17575 -1145 17580 -1140
rect 17620 -1140 17660 -1135
rect 17620 -1145 17625 -1140
rect 17575 -1165 17625 -1145
rect 17575 -1170 17580 -1165
rect 17540 -1175 17580 -1170
rect 17620 -1170 17625 -1165
rect 17655 -1145 17660 -1140
rect 17700 -1140 17740 -1135
rect 17700 -1145 17705 -1140
rect 17655 -1165 17705 -1145
rect 17655 -1170 17660 -1165
rect 17620 -1175 17660 -1170
rect 17700 -1170 17705 -1165
rect 17735 -1170 17740 -1140
rect 17700 -1175 17740 -1170
rect 17780 -1140 17820 -1135
rect 17780 -1170 17785 -1140
rect 17815 -1145 17820 -1140
rect 17860 -1140 17900 -1135
rect 17860 -1145 17865 -1140
rect 17815 -1165 17865 -1145
rect 17815 -1170 17820 -1165
rect 17780 -1175 17820 -1170
rect 17860 -1170 17865 -1165
rect 17895 -1145 17900 -1140
rect 17940 -1140 17980 -1135
rect 17940 -1145 17945 -1140
rect 17895 -1165 17945 -1145
rect 17895 -1170 17900 -1165
rect 17860 -1175 17900 -1170
rect 17940 -1170 17945 -1165
rect 17975 -1145 17980 -1140
rect 18020 -1140 18060 -1135
rect 18020 -1145 18025 -1140
rect 17975 -1165 18025 -1145
rect 17975 -1170 17980 -1165
rect 17940 -1175 17980 -1170
rect 18020 -1170 18025 -1165
rect 18055 -1145 18060 -1140
rect 18100 -1140 18140 -1135
rect 18100 -1145 18105 -1140
rect 18055 -1165 18105 -1145
rect 18055 -1170 18060 -1165
rect 18020 -1175 18060 -1170
rect 18100 -1170 18105 -1165
rect 18135 -1145 18140 -1140
rect 18180 -1140 18220 -1135
rect 18180 -1145 18185 -1140
rect 18135 -1165 18185 -1145
rect 18135 -1170 18140 -1165
rect 18100 -1175 18140 -1170
rect 18180 -1170 18185 -1165
rect 18215 -1145 18220 -1140
rect 18260 -1140 18300 -1135
rect 18260 -1145 18265 -1140
rect 18215 -1165 18265 -1145
rect 18215 -1170 18220 -1165
rect 18180 -1175 18220 -1170
rect 18260 -1170 18265 -1165
rect 18295 -1145 18300 -1140
rect 18340 -1140 18380 -1135
rect 18340 -1145 18345 -1140
rect 18295 -1165 18345 -1145
rect 18295 -1170 18300 -1165
rect 18260 -1175 18300 -1170
rect 18340 -1170 18345 -1165
rect 18375 -1145 18380 -1140
rect 18420 -1140 18460 -1135
rect 18420 -1145 18425 -1140
rect 18375 -1165 18425 -1145
rect 18375 -1170 18380 -1165
rect 18340 -1175 18380 -1170
rect 18420 -1170 18425 -1165
rect 18455 -1145 18460 -1140
rect 18500 -1140 18540 -1135
rect 18500 -1145 18505 -1140
rect 18455 -1165 18505 -1145
rect 18455 -1170 18460 -1165
rect 18420 -1175 18460 -1170
rect 18500 -1170 18505 -1165
rect 18535 -1145 18540 -1140
rect 18580 -1140 18620 -1135
rect 18580 -1145 18585 -1140
rect 18535 -1165 18585 -1145
rect 18535 -1170 18540 -1165
rect 18500 -1175 18540 -1170
rect 18580 -1170 18585 -1165
rect 18615 -1145 18620 -1140
rect 18660 -1140 18700 -1135
rect 18660 -1145 18665 -1140
rect 18615 -1165 18665 -1145
rect 18615 -1170 18620 -1165
rect 18580 -1175 18620 -1170
rect 18660 -1170 18665 -1165
rect 18695 -1145 18700 -1140
rect 18740 -1140 18780 -1135
rect 18740 -1145 18745 -1140
rect 18695 -1165 18745 -1145
rect 18695 -1170 18700 -1165
rect 18660 -1175 18700 -1170
rect 18740 -1170 18745 -1165
rect 18775 -1170 18780 -1140
rect 18740 -1175 18780 -1170
rect 16205 -1225 16245 -1220
rect 16205 -1255 16210 -1225
rect 16240 -1230 16245 -1225
rect 16700 -1225 16740 -1220
rect 16700 -1230 16705 -1225
rect 16240 -1250 16705 -1230
rect 16240 -1255 16245 -1250
rect 16205 -1260 16245 -1255
rect 16700 -1255 16705 -1250
rect 16735 -1255 16740 -1225
rect 16700 -1260 16740 -1255
rect 18895 -1225 18935 -1220
rect 18895 -1255 18900 -1225
rect 18930 -1255 18935 -1225
rect 18895 -1260 18935 -1255
rect 16160 -1325 16200 -1320
rect 16160 -1355 16165 -1325
rect 16195 -1330 16200 -1325
rect 16595 -1325 16635 -1320
rect 16595 -1330 16600 -1325
rect 16195 -1350 16600 -1330
rect 16195 -1355 16200 -1350
rect 16160 -1360 16200 -1355
rect 16595 -1355 16600 -1350
rect 16630 -1330 16635 -1325
rect 16705 -1325 16745 -1320
rect 16705 -1330 16710 -1325
rect 16630 -1350 16710 -1330
rect 16630 -1355 16635 -1350
rect 16595 -1360 16635 -1355
rect 16705 -1355 16710 -1350
rect 16740 -1330 16745 -1325
rect 17300 -1325 17340 -1320
rect 17300 -1330 17305 -1325
rect 16740 -1350 17305 -1330
rect 16740 -1355 16745 -1350
rect 16705 -1360 16745 -1355
rect 17300 -1355 17305 -1350
rect 17335 -1330 17340 -1325
rect 17780 -1325 17820 -1320
rect 17780 -1330 17785 -1325
rect 17335 -1350 17785 -1330
rect 17335 -1355 17340 -1350
rect 17300 -1360 17340 -1355
rect 17780 -1355 17785 -1350
rect 17815 -1330 17820 -1325
rect 18260 -1325 18300 -1320
rect 18260 -1330 18265 -1325
rect 17815 -1350 18265 -1330
rect 17815 -1355 17820 -1350
rect 17780 -1360 17820 -1355
rect 18260 -1355 18265 -1350
rect 18295 -1355 18300 -1325
rect 18260 -1360 18300 -1355
rect 16540 -1410 18575 -1405
rect 16540 -1440 16545 -1410
rect 16575 -1440 16655 -1410
rect 16685 -1440 16765 -1410
rect 16795 -1440 16825 -1410
rect 16855 -1440 17030 -1410
rect 17060 -1440 17140 -1410
rect 17170 -1440 17250 -1410
rect 17280 -1440 17360 -1410
rect 17390 -1440 17470 -1410
rect 17500 -1440 17620 -1410
rect 17650 -1440 17730 -1410
rect 17760 -1440 17840 -1410
rect 17870 -1440 17950 -1410
rect 17980 -1440 18100 -1410
rect 18130 -1440 18210 -1410
rect 18240 -1440 18320 -1410
rect 18350 -1440 18430 -1410
rect 18460 -1440 18540 -1410
rect 18570 -1440 18575 -1410
rect 16540 -1450 18575 -1440
rect 16540 -1480 16545 -1450
rect 16575 -1480 16655 -1450
rect 16685 -1480 16765 -1450
rect 16795 -1480 16825 -1450
rect 16855 -1480 17030 -1450
rect 17060 -1480 17140 -1450
rect 17170 -1480 17250 -1450
rect 17280 -1480 17360 -1450
rect 17390 -1480 17470 -1450
rect 17500 -1480 17620 -1450
rect 17650 -1480 17730 -1450
rect 17760 -1480 17840 -1450
rect 17870 -1480 17950 -1450
rect 17980 -1480 18100 -1450
rect 18130 -1480 18210 -1450
rect 18240 -1480 18320 -1450
rect 18350 -1480 18430 -1450
rect 18460 -1480 18540 -1450
rect 18570 -1480 18575 -1450
rect 16540 -1490 18575 -1480
rect 16540 -1520 16545 -1490
rect 16575 -1520 16655 -1490
rect 16685 -1520 16765 -1490
rect 16795 -1520 16825 -1490
rect 16855 -1520 17030 -1490
rect 17060 -1520 17140 -1490
rect 17170 -1520 17250 -1490
rect 17280 -1520 17360 -1490
rect 17390 -1520 17470 -1490
rect 17500 -1520 17620 -1490
rect 17650 -1520 17730 -1490
rect 17760 -1520 17840 -1490
rect 17870 -1520 17950 -1490
rect 17980 -1520 18100 -1490
rect 18130 -1520 18210 -1490
rect 18240 -1520 18320 -1490
rect 18350 -1520 18430 -1490
rect 18460 -1520 18540 -1490
rect 18570 -1520 18575 -1490
rect 16540 -1525 18575 -1520
rect 17190 -1660 17450 -1655
rect 17190 -1690 17195 -1660
rect 17225 -1690 17415 -1660
rect 17445 -1690 17450 -1660
rect 17190 -1695 17450 -1690
rect 17670 -1660 17710 -1655
rect 17670 -1690 17675 -1660
rect 17705 -1665 17710 -1660
rect 17780 -1660 17820 -1655
rect 17780 -1665 17785 -1660
rect 17705 -1685 17785 -1665
rect 17705 -1690 17710 -1685
rect 17670 -1695 17710 -1690
rect 17780 -1690 17785 -1685
rect 17815 -1665 17820 -1660
rect 17890 -1660 17930 -1655
rect 17890 -1665 17895 -1660
rect 17815 -1685 17895 -1665
rect 17815 -1690 17820 -1685
rect 17780 -1695 17820 -1690
rect 17890 -1690 17895 -1685
rect 17925 -1690 17930 -1660
rect 17890 -1695 17930 -1690
rect 18150 -1660 18410 -1655
rect 18150 -1690 18155 -1660
rect 18185 -1690 18375 -1660
rect 18405 -1690 18410 -1660
rect 18150 -1695 18410 -1690
rect 16030 -1715 16070 -1710
rect 16030 -1745 16035 -1715
rect 16065 -1720 16070 -1715
rect 17080 -1715 17120 -1710
rect 17080 -1720 17085 -1715
rect 16065 -1740 17085 -1720
rect 16065 -1745 16070 -1740
rect 16030 -1750 16070 -1745
rect 17080 -1745 17085 -1740
rect 17115 -1720 17120 -1715
rect 17300 -1715 17340 -1710
rect 17300 -1720 17305 -1715
rect 17115 -1740 17305 -1720
rect 17115 -1745 17120 -1740
rect 17080 -1750 17120 -1745
rect 17300 -1745 17305 -1740
rect 17335 -1720 17340 -1715
rect 18260 -1715 18300 -1710
rect 18260 -1720 18265 -1715
rect 17335 -1740 18265 -1720
rect 17335 -1745 17340 -1740
rect 17300 -1750 17340 -1745
rect 18260 -1745 18265 -1740
rect 18295 -1720 18300 -1715
rect 18480 -1715 18520 -1710
rect 18480 -1720 18485 -1715
rect 18295 -1740 18485 -1720
rect 18295 -1745 18300 -1740
rect 18260 -1750 18300 -1745
rect 18480 -1745 18485 -1740
rect 18515 -1745 18520 -1715
rect 18480 -1750 18520 -1745
rect 15785 -1770 17230 -1765
rect 15785 -1800 15790 -1770
rect 15820 -1800 17195 -1770
rect 17225 -1800 17230 -1770
rect 15785 -1810 17230 -1800
rect 15785 -1840 15790 -1810
rect 15820 -1840 17195 -1810
rect 17225 -1840 17230 -1810
rect 15785 -1845 17230 -1840
rect 18370 -1770 19815 -1765
rect 18370 -1800 18375 -1770
rect 18405 -1800 19780 -1770
rect 19810 -1800 19815 -1770
rect 18370 -1810 19815 -1800
rect 18370 -1840 18375 -1810
rect 18405 -1840 19780 -1810
rect 19810 -1840 19815 -1810
rect 18370 -1845 19815 -1840
rect 16105 -1900 16145 -1895
rect 16105 -1930 16110 -1900
rect 16140 -1905 16145 -1900
rect 16705 -1900 16745 -1895
rect 16705 -1905 16710 -1900
rect 16140 -1925 16710 -1905
rect 16140 -1930 16145 -1925
rect 16105 -1935 16145 -1930
rect 16705 -1930 16710 -1925
rect 16740 -1930 16745 -1900
rect 16705 -1935 16745 -1930
rect 17780 -1900 17820 -1895
rect 17780 -1930 17785 -1900
rect 17815 -1905 17820 -1900
rect 19535 -1900 19575 -1895
rect 19535 -1905 19540 -1900
rect 17815 -1925 19540 -1905
rect 17815 -1930 17820 -1925
rect 17780 -1935 17820 -1930
rect 19535 -1930 19540 -1925
rect 19570 -1930 19575 -1900
rect 19535 -1935 19575 -1930
rect 16155 -1950 16195 -1945
rect 16155 -1980 16160 -1950
rect 16190 -1955 16195 -1950
rect 19325 -1950 19365 -1945
rect 19325 -1955 19330 -1950
rect 16190 -1975 19330 -1955
rect 16190 -1980 16195 -1975
rect 16155 -1985 16195 -1980
rect 19325 -1980 19330 -1975
rect 19360 -1980 19365 -1950
rect 19325 -1985 19365 -1980
rect 16260 -2000 16300 -1995
rect 16260 -2030 16265 -2000
rect 16295 -2005 16300 -2000
rect 16480 -2000 16520 -1995
rect 16480 -2005 16485 -2000
rect 16295 -2025 16485 -2005
rect 16295 -2030 16300 -2025
rect 16260 -2035 16300 -2030
rect 16480 -2030 16485 -2025
rect 16515 -2005 16520 -2000
rect 16730 -2000 16770 -1995
rect 16730 -2005 16735 -2000
rect 16515 -2025 16735 -2005
rect 16515 -2030 16520 -2025
rect 16480 -2035 16520 -2030
rect 16730 -2030 16735 -2025
rect 16765 -2030 16770 -2000
rect 16730 -2035 16770 -2030
rect 17195 -2000 17425 -1995
rect 17195 -2030 17200 -2000
rect 17230 -2030 17430 -2000
rect 17195 -2035 17430 -2030
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2005 19500 -2000
rect 18164 -2035 19085 -2005
rect 19115 -2035 19465 -2005
rect 19495 -2035 19500 -2005
rect 18165 -2040 19500 -2035
rect 17195 -2060 17235 -2055
rect 17195 -2090 17200 -2060
rect 17230 -2065 17235 -2060
rect 18830 -2060 18870 -2055
rect 18830 -2065 18835 -2060
rect 17230 -2085 18835 -2065
rect 17230 -2090 17235 -2085
rect 17195 -2095 17235 -2090
rect 18830 -2090 18835 -2085
rect 18865 -2090 18870 -2060
rect 18830 -2095 18870 -2090
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2997 19440 -2992
rect 16160 -3025 16195 -3020
rect 19405 -3037 19440 -3032
rect 16160 -3065 16195 -3060
rect 16730 -3105 16770 -3100
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3120 15860 -3115
rect 15950 -3116 15985 -3111
rect 15855 -3140 15950 -3120
rect 15855 -3145 15860 -3140
rect 15820 -3150 15860 -3145
rect 16730 -3135 16735 -3105
rect 16765 -3110 16770 -3105
rect 17780 -3105 17820 -3100
rect 17780 -3110 17785 -3105
rect 16765 -3130 17785 -3110
rect 16765 -3135 16770 -3130
rect 16730 -3140 16770 -3135
rect 17780 -3135 17785 -3130
rect 17815 -3135 17820 -3105
rect 17780 -3140 17820 -3135
rect 18615 -3105 18655 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3110 18655 -3105
rect 18830 -3105 18870 -3100
rect 18830 -3110 18835 -3105
rect 18650 -3130 18835 -3110
rect 18650 -3135 18655 -3130
rect 18615 -3140 18655 -3135
rect 18830 -3135 18835 -3130
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 15950 -3156 15985 -3151
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 15960 -3830 15980 -3829
rect 19620 -3830 19640 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 16290 -3935 16310 -3934
rect 19290 -3935 19310 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4195 16285 -4190
rect 15665 -4215 16285 -4195
rect 16280 -4220 16285 -4215
rect 16315 -4195 16320 -4190
rect 16605 -4190 16645 -4185
rect 16605 -4195 16610 -4190
rect 16315 -4215 16610 -4195
rect 16315 -4220 16320 -4215
rect 16280 -4225 16320 -4220
rect 16605 -4220 16610 -4215
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4270 15860 -4265
rect 17250 -4265 17300 -4255
rect 17250 -4270 17260 -4265
rect 15855 -4290 17260 -4270
rect 15855 -4295 15860 -4290
rect 15820 -4300 15860 -4295
rect 17250 -4295 17260 -4290
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4270 17820 -4265
rect 18955 -4265 18995 -4260
rect 18955 -4270 18960 -4265
rect 17815 -4290 18960 -4270
rect 17815 -4295 17820 -4290
rect 17780 -4300 17820 -4295
rect 18955 -4295 18960 -4290
rect 18990 -4270 18995 -4265
rect 19280 -4265 19320 -4260
rect 19280 -4270 19285 -4265
rect 18990 -4290 19285 -4270
rect 18990 -4295 18995 -4290
rect 18955 -4300 18995 -4295
rect 19280 -4295 19285 -4290
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4320 15765 -4315
rect 16900 -4315 16950 -4305
rect 16900 -4320 16910 -4315
rect 15760 -4340 16910 -4320
rect 15760 -4345 15765 -4340
rect 15725 -4350 15765 -4345
rect 16900 -4345 16910 -4340
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4320 18700 -4315
rect 19720 -4315 19760 -4310
rect 19720 -4320 19725 -4315
rect 18690 -4340 19725 -4320
rect 18690 -4345 18700 -4340
rect 18650 -4355 18700 -4345
rect 19720 -4345 19725 -4340
rect 19755 -4345 19760 -4315
rect 19720 -4350 19760 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4365 15990 -4360
rect 16205 -4360 16245 -4355
rect 16205 -4365 16210 -4360
rect 15985 -4385 16210 -4365
rect 15985 -4390 15990 -4385
rect 15950 -4395 15990 -4390
rect 16205 -4390 16210 -4385
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4365 19395 -4360
rect 19610 -4360 19650 -4355
rect 19610 -4365 19615 -4360
rect 19390 -4385 19615 -4365
rect 19390 -4390 19395 -4385
rect 19355 -4395 19395 -4390
rect 19610 -4390 19615 -4385
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4415 17995 -4410
rect 17990 -4435 19905 -4415
rect 17990 -4440 17995 -4435
rect 17955 -4445 17995 -4440
<< via2 >>
rect 17260 -4295 17290 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 17960 -4440 17990 -4410
<< metal3 >>
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 17250 -4305 17300 -4300
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4355 16950 -4350
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4355 18700 -4350
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4520 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4520 17995 -4440
rect 19355 -4520 19395 -4390
rect 15760 -4615 15990 -4520
rect 16110 -4615 16340 -4520
rect 16460 -4615 16690 -4520
rect 16810 -4615 17040 -4520
rect 15760 -4665 17040 -4615
rect 15760 -4750 15990 -4665
rect 16110 -4750 16340 -4665
rect 16460 -4750 16690 -4665
rect 16810 -4750 17040 -4665
rect 17160 -4615 17390 -4520
rect 17510 -4615 17740 -4520
rect 17860 -4615 18090 -4520
rect 18210 -4615 18440 -4520
rect 17160 -4665 18440 -4615
rect 17160 -4750 17390 -4665
rect 17510 -4750 17740 -4665
rect 17860 -4750 18090 -4665
rect 18210 -4750 18440 -4665
rect 18560 -4615 18790 -4520
rect 18910 -4615 19140 -4520
rect 19260 -4615 19490 -4520
rect 19610 -4615 19840 -4520
rect 18560 -4665 19840 -4615
rect 18560 -4750 18790 -4665
rect 18910 -4750 19140 -4665
rect 19260 -4750 19490 -4665
rect 19610 -4750 19840 -4665
rect 16200 -4870 16250 -4750
rect 17950 -4870 18000 -4750
rect 19350 -4870 19400 -4750
rect 15760 -4965 15990 -4870
rect 16110 -4965 16340 -4870
rect 16460 -4965 16690 -4870
rect 16810 -4965 17040 -4870
rect 15760 -5015 17040 -4965
rect 15760 -5100 15990 -5015
rect 16110 -5100 16340 -5015
rect 16460 -5100 16690 -5015
rect 16810 -5100 17040 -5015
rect 17160 -4965 17390 -4870
rect 17510 -4965 17740 -4870
rect 17860 -4965 18090 -4870
rect 18210 -4965 18440 -4870
rect 17160 -5015 18440 -4965
rect 17160 -5100 17390 -5015
rect 17510 -5100 17740 -5015
rect 17860 -5100 18090 -5015
rect 18210 -5100 18440 -5015
rect 18560 -4965 18790 -4870
rect 18910 -4965 19140 -4870
rect 19260 -4965 19490 -4870
rect 19610 -4965 19840 -4870
rect 18560 -5015 19840 -4965
rect 18560 -5100 18790 -5015
rect 18910 -5100 19140 -5015
rect 19260 -5100 19490 -5015
rect 19610 -5100 19840 -5015
rect 16200 -5220 16250 -5100
rect 17950 -5220 18000 -5100
rect 19350 -5220 19400 -5100
rect 15760 -5315 15990 -5220
rect 16110 -5315 16340 -5220
rect 16460 -5315 16690 -5220
rect 16810 -5315 17040 -5220
rect 15760 -5365 17040 -5315
rect 15760 -5450 15990 -5365
rect 16110 -5450 16340 -5365
rect 16460 -5450 16690 -5365
rect 16810 -5450 17040 -5365
rect 17160 -5315 17390 -5220
rect 17510 -5315 17740 -5220
rect 17860 -5315 18090 -5220
rect 18210 -5315 18440 -5220
rect 17160 -5365 18440 -5315
rect 17160 -5450 17390 -5365
rect 17510 -5450 17740 -5365
rect 17860 -5450 18090 -5365
rect 18210 -5450 18440 -5365
rect 18560 -5315 18790 -5220
rect 18910 -5315 19140 -5220
rect 19260 -5315 19490 -5220
rect 19610 -5315 19840 -5220
rect 18560 -5365 19840 -5315
rect 18560 -5450 18790 -5365
rect 18910 -5450 19140 -5365
rect 19260 -5450 19490 -5365
rect 19610 -5450 19840 -5365
rect 16200 -5570 16250 -5450
rect 17950 -5570 18000 -5450
rect 19350 -5570 19400 -5450
rect 15760 -5665 15990 -5570
rect 16110 -5665 16340 -5570
rect 16460 -5665 16690 -5570
rect 16810 -5665 17040 -5570
rect 15760 -5715 17040 -5665
rect 15760 -5800 15990 -5715
rect 16110 -5800 16340 -5715
rect 16460 -5800 16690 -5715
rect 16810 -5800 17040 -5715
rect 17160 -5665 17390 -5570
rect 17510 -5665 17740 -5570
rect 17860 -5665 18090 -5570
rect 18210 -5665 18440 -5570
rect 17160 -5715 18440 -5665
rect 17160 -5800 17390 -5715
rect 17510 -5800 17740 -5715
rect 17860 -5800 18090 -5715
rect 18210 -5800 18440 -5715
rect 18560 -5665 18790 -5570
rect 18910 -5665 19140 -5570
rect 19260 -5665 19490 -5570
rect 19610 -5665 19840 -5570
rect 18560 -5715 19840 -5665
rect 18560 -5800 18790 -5715
rect 18910 -5800 19140 -5715
rect 19260 -5800 19490 -5715
rect 19610 -5800 19840 -5715
rect 16200 -5920 16250 -5800
rect 17950 -5920 18000 -5800
rect 19350 -5920 19400 -5800
rect 15760 -6015 15990 -5920
rect 16110 -6015 16340 -5920
rect 16460 -6015 16690 -5920
rect 16810 -6015 17040 -5920
rect 15760 -6065 17040 -6015
rect 15760 -6150 15990 -6065
rect 16110 -6150 16340 -6065
rect 16460 -6150 16690 -6065
rect 16810 -6150 17040 -6065
rect 17160 -6015 17390 -5920
rect 17510 -6015 17740 -5920
rect 17860 -6015 18090 -5920
rect 18210 -6015 18440 -5920
rect 17160 -6065 18440 -6015
rect 17160 -6150 17390 -6065
rect 17510 -6150 17740 -6065
rect 17860 -6150 18090 -6065
rect 18210 -6150 18440 -6065
rect 18560 -6015 18790 -5920
rect 18910 -6015 19140 -5920
rect 19260 -6015 19490 -5920
rect 19610 -6015 19840 -5920
rect 18560 -6065 19840 -6015
rect 18560 -6150 18790 -6065
rect 18910 -6150 19140 -6065
rect 19260 -6150 19490 -6065
rect 19610 -6150 19840 -6065
<< via3 >>
rect 17255 -4265 17295 -4260
rect 17255 -4295 17260 -4265
rect 17260 -4295 17290 -4265
rect 17290 -4295 17295 -4265
rect 17255 -4300 17295 -4295
rect 16905 -4315 16945 -4310
rect 16905 -4345 16910 -4315
rect 16910 -4345 16940 -4315
rect 16940 -4345 16945 -4315
rect 16905 -4350 16945 -4345
rect 18655 -4315 18695 -4310
rect 18655 -4345 18660 -4315
rect 18660 -4345 18690 -4315
rect 18690 -4345 18695 -4315
rect 18655 -4350 18695 -4345
<< mimcap >>
rect 15775 -4620 15975 -4535
rect 15775 -4660 15855 -4620
rect 15895 -4660 15975 -4620
rect 15775 -4735 15975 -4660
rect 16125 -4620 16325 -4535
rect 16125 -4660 16205 -4620
rect 16245 -4660 16325 -4620
rect 16125 -4735 16325 -4660
rect 16475 -4620 16675 -4535
rect 16475 -4660 16555 -4620
rect 16595 -4660 16675 -4620
rect 16475 -4735 16675 -4660
rect 16825 -4620 17025 -4535
rect 16825 -4660 16905 -4620
rect 16945 -4660 17025 -4620
rect 16825 -4735 17025 -4660
rect 17175 -4620 17375 -4535
rect 17175 -4660 17255 -4620
rect 17295 -4660 17375 -4620
rect 17175 -4735 17375 -4660
rect 17525 -4620 17725 -4535
rect 17525 -4660 17605 -4620
rect 17645 -4660 17725 -4620
rect 17525 -4735 17725 -4660
rect 17875 -4620 18075 -4535
rect 17875 -4660 17955 -4620
rect 17995 -4660 18075 -4620
rect 17875 -4735 18075 -4660
rect 18225 -4620 18425 -4535
rect 18225 -4660 18305 -4620
rect 18345 -4660 18425 -4620
rect 18225 -4735 18425 -4660
rect 18575 -4620 18775 -4535
rect 18575 -4660 18655 -4620
rect 18695 -4660 18775 -4620
rect 18575 -4735 18775 -4660
rect 18925 -4620 19125 -4535
rect 18925 -4660 19005 -4620
rect 19045 -4660 19125 -4620
rect 18925 -4735 19125 -4660
rect 19275 -4620 19475 -4535
rect 19275 -4660 19355 -4620
rect 19395 -4660 19475 -4620
rect 19275 -4735 19475 -4660
rect 19625 -4620 19825 -4535
rect 19625 -4660 19705 -4620
rect 19745 -4660 19825 -4620
rect 19625 -4735 19825 -4660
rect 15775 -4970 15975 -4885
rect 15775 -5010 15855 -4970
rect 15895 -5010 15975 -4970
rect 15775 -5085 15975 -5010
rect 16125 -4970 16325 -4885
rect 16125 -5010 16205 -4970
rect 16245 -5010 16325 -4970
rect 16125 -5085 16325 -5010
rect 16475 -4970 16675 -4885
rect 16475 -5010 16555 -4970
rect 16595 -5010 16675 -4970
rect 16475 -5085 16675 -5010
rect 16825 -4970 17025 -4885
rect 16825 -5010 16905 -4970
rect 16945 -5010 17025 -4970
rect 16825 -5085 17025 -5010
rect 17175 -4970 17375 -4885
rect 17175 -5010 17255 -4970
rect 17295 -5010 17375 -4970
rect 17175 -5085 17375 -5010
rect 17525 -4970 17725 -4885
rect 17525 -5010 17605 -4970
rect 17645 -5010 17725 -4970
rect 17525 -5085 17725 -5010
rect 17875 -4970 18075 -4885
rect 17875 -5010 17955 -4970
rect 17995 -5010 18075 -4970
rect 17875 -5085 18075 -5010
rect 18225 -4970 18425 -4885
rect 18225 -5010 18305 -4970
rect 18345 -5010 18425 -4970
rect 18225 -5085 18425 -5010
rect 18575 -4970 18775 -4885
rect 18575 -5010 18655 -4970
rect 18695 -5010 18775 -4970
rect 18575 -5085 18775 -5010
rect 18925 -4970 19125 -4885
rect 18925 -5010 19005 -4970
rect 19045 -5010 19125 -4970
rect 18925 -5085 19125 -5010
rect 19275 -4970 19475 -4885
rect 19275 -5010 19355 -4970
rect 19395 -5010 19475 -4970
rect 19275 -5085 19475 -5010
rect 19625 -4970 19825 -4885
rect 19625 -5010 19705 -4970
rect 19745 -5010 19825 -4970
rect 19625 -5085 19825 -5010
rect 15775 -5320 15975 -5235
rect 15775 -5360 15855 -5320
rect 15895 -5360 15975 -5320
rect 15775 -5435 15975 -5360
rect 16125 -5320 16325 -5235
rect 16125 -5360 16205 -5320
rect 16245 -5360 16325 -5320
rect 16125 -5435 16325 -5360
rect 16475 -5320 16675 -5235
rect 16475 -5360 16555 -5320
rect 16595 -5360 16675 -5320
rect 16475 -5435 16675 -5360
rect 16825 -5320 17025 -5235
rect 16825 -5360 16905 -5320
rect 16945 -5360 17025 -5320
rect 16825 -5435 17025 -5360
rect 17175 -5320 17375 -5235
rect 17175 -5360 17255 -5320
rect 17295 -5360 17375 -5320
rect 17175 -5435 17375 -5360
rect 17525 -5320 17725 -5235
rect 17525 -5360 17605 -5320
rect 17645 -5360 17725 -5320
rect 17525 -5435 17725 -5360
rect 17875 -5320 18075 -5235
rect 17875 -5360 17955 -5320
rect 17995 -5360 18075 -5320
rect 17875 -5435 18075 -5360
rect 18225 -5320 18425 -5235
rect 18225 -5360 18305 -5320
rect 18345 -5360 18425 -5320
rect 18225 -5435 18425 -5360
rect 18575 -5320 18775 -5235
rect 18575 -5360 18655 -5320
rect 18695 -5360 18775 -5320
rect 18575 -5435 18775 -5360
rect 18925 -5320 19125 -5235
rect 18925 -5360 19005 -5320
rect 19045 -5360 19125 -5320
rect 18925 -5435 19125 -5360
rect 19275 -5320 19475 -5235
rect 19275 -5360 19355 -5320
rect 19395 -5360 19475 -5320
rect 19275 -5435 19475 -5360
rect 19625 -5320 19825 -5235
rect 19625 -5360 19705 -5320
rect 19745 -5360 19825 -5320
rect 19625 -5435 19825 -5360
rect 15775 -5670 15975 -5585
rect 15775 -5710 15855 -5670
rect 15895 -5710 15975 -5670
rect 15775 -5785 15975 -5710
rect 16125 -5670 16325 -5585
rect 16125 -5710 16205 -5670
rect 16245 -5710 16325 -5670
rect 16125 -5785 16325 -5710
rect 16475 -5670 16675 -5585
rect 16475 -5710 16555 -5670
rect 16595 -5710 16675 -5670
rect 16475 -5785 16675 -5710
rect 16825 -5670 17025 -5585
rect 16825 -5710 16905 -5670
rect 16945 -5710 17025 -5670
rect 16825 -5785 17025 -5710
rect 17175 -5670 17375 -5585
rect 17175 -5710 17255 -5670
rect 17295 -5710 17375 -5670
rect 17175 -5785 17375 -5710
rect 17525 -5670 17725 -5585
rect 17525 -5710 17605 -5670
rect 17645 -5710 17725 -5670
rect 17525 -5785 17725 -5710
rect 17875 -5670 18075 -5585
rect 17875 -5710 17955 -5670
rect 17995 -5710 18075 -5670
rect 17875 -5785 18075 -5710
rect 18225 -5670 18425 -5585
rect 18225 -5710 18305 -5670
rect 18345 -5710 18425 -5670
rect 18225 -5785 18425 -5710
rect 18575 -5670 18775 -5585
rect 18575 -5710 18655 -5670
rect 18695 -5710 18775 -5670
rect 18575 -5785 18775 -5710
rect 18925 -5670 19125 -5585
rect 18925 -5710 19005 -5670
rect 19045 -5710 19125 -5670
rect 18925 -5785 19125 -5710
rect 19275 -5670 19475 -5585
rect 19275 -5710 19355 -5670
rect 19395 -5710 19475 -5670
rect 19275 -5785 19475 -5710
rect 19625 -5670 19825 -5585
rect 19625 -5710 19705 -5670
rect 19745 -5710 19825 -5670
rect 19625 -5785 19825 -5710
rect 15775 -6020 15975 -5935
rect 15775 -6060 15855 -6020
rect 15895 -6060 15975 -6020
rect 15775 -6135 15975 -6060
rect 16125 -6020 16325 -5935
rect 16125 -6060 16205 -6020
rect 16245 -6060 16325 -6020
rect 16125 -6135 16325 -6060
rect 16475 -6020 16675 -5935
rect 16475 -6060 16555 -6020
rect 16595 -6060 16675 -6020
rect 16475 -6135 16675 -6060
rect 16825 -6020 17025 -5935
rect 16825 -6060 16905 -6020
rect 16945 -6060 17025 -6020
rect 16825 -6135 17025 -6060
rect 17175 -6020 17375 -5935
rect 17175 -6060 17255 -6020
rect 17295 -6060 17375 -6020
rect 17175 -6135 17375 -6060
rect 17525 -6020 17725 -5935
rect 17525 -6060 17605 -6020
rect 17645 -6060 17725 -6020
rect 17525 -6135 17725 -6060
rect 17875 -6020 18075 -5935
rect 17875 -6060 17955 -6020
rect 17995 -6060 18075 -6020
rect 17875 -6135 18075 -6060
rect 18225 -6020 18425 -5935
rect 18225 -6060 18305 -6020
rect 18345 -6060 18425 -6020
rect 18225 -6135 18425 -6060
rect 18575 -6020 18775 -5935
rect 18575 -6060 18655 -6020
rect 18695 -6060 18775 -6020
rect 18575 -6135 18775 -6060
rect 18925 -6020 19125 -5935
rect 18925 -6060 19005 -6020
rect 19045 -6060 19125 -6020
rect 18925 -6135 19125 -6060
rect 19275 -6020 19475 -5935
rect 19275 -6060 19355 -6020
rect 19395 -6060 19475 -6020
rect 19275 -6135 19475 -6060
rect 19625 -6020 19825 -5935
rect 19625 -6060 19705 -6020
rect 19745 -6060 19825 -6020
rect 19625 -6135 19825 -6060
<< mimcapcontact >>
rect 15855 -4660 15895 -4620
rect 16205 -4660 16245 -4620
rect 16555 -4660 16595 -4620
rect 16905 -4660 16945 -4620
rect 17255 -4660 17295 -4620
rect 17605 -4660 17645 -4620
rect 17955 -4660 17995 -4620
rect 18305 -4660 18345 -4620
rect 18655 -4660 18695 -4620
rect 19005 -4660 19045 -4620
rect 19355 -4660 19395 -4620
rect 19705 -4660 19745 -4620
rect 15855 -5010 15895 -4970
rect 16205 -5010 16245 -4970
rect 16555 -5010 16595 -4970
rect 16905 -5010 16945 -4970
rect 17255 -5010 17295 -4970
rect 17605 -5010 17645 -4970
rect 17955 -5010 17995 -4970
rect 18305 -5010 18345 -4970
rect 18655 -5010 18695 -4970
rect 19005 -5010 19045 -4970
rect 19355 -5010 19395 -4970
rect 19705 -5010 19745 -4970
rect 15855 -5360 15895 -5320
rect 16205 -5360 16245 -5320
rect 16555 -5360 16595 -5320
rect 16905 -5360 16945 -5320
rect 17255 -5360 17295 -5320
rect 17605 -5360 17645 -5320
rect 17955 -5360 17995 -5320
rect 18305 -5360 18345 -5320
rect 18655 -5360 18695 -5320
rect 19005 -5360 19045 -5320
rect 19355 -5360 19395 -5320
rect 19705 -5360 19745 -5320
rect 15855 -5710 15895 -5670
rect 16205 -5710 16245 -5670
rect 16555 -5710 16595 -5670
rect 16905 -5710 16945 -5670
rect 17255 -5710 17295 -5670
rect 17605 -5710 17645 -5670
rect 17955 -5710 17995 -5670
rect 18305 -5710 18345 -5670
rect 18655 -5710 18695 -5670
rect 19005 -5710 19045 -5670
rect 19355 -5710 19395 -5670
rect 19705 -5710 19745 -5670
rect 15855 -6060 15895 -6020
rect 16205 -6060 16245 -6020
rect 16555 -6060 16595 -6020
rect 16905 -6060 16945 -6020
rect 17255 -6060 17295 -6020
rect 17605 -6060 17645 -6020
rect 17955 -6060 17995 -6020
rect 18305 -6060 18345 -6020
rect 18655 -6060 18695 -6020
rect 19005 -6060 19045 -6020
rect 19355 -6060 19395 -6020
rect 19705 -6060 19745 -6020
<< metal4 >>
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4615 16950 -4350
rect 15850 -4620 16950 -4615
rect 15850 -4660 15855 -4620
rect 15895 -4660 16205 -4620
rect 16245 -4660 16555 -4620
rect 16595 -4660 16905 -4620
rect 16945 -4660 16950 -4620
rect 15850 -4665 16950 -4660
rect 17250 -4615 17300 -4300
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4615 18700 -4350
rect 17250 -4620 18350 -4615
rect 17250 -4660 17255 -4620
rect 17295 -4660 17605 -4620
rect 17645 -4660 17955 -4620
rect 17995 -4660 18305 -4620
rect 18345 -4660 18350 -4620
rect 17250 -4665 18350 -4660
rect 18650 -4620 19750 -4615
rect 18650 -4660 18655 -4620
rect 18695 -4660 19005 -4620
rect 19045 -4660 19355 -4620
rect 19395 -4660 19705 -4620
rect 19745 -4660 19750 -4620
rect 18650 -4665 19750 -4660
rect 16200 -4965 16250 -4665
rect 17950 -4965 18000 -4665
rect 19350 -4965 19400 -4665
rect 15850 -4970 16950 -4965
rect 15850 -5010 15855 -4970
rect 15895 -5010 16205 -4970
rect 16245 -5010 16555 -4970
rect 16595 -5010 16905 -4970
rect 16945 -5010 16950 -4970
rect 15850 -5015 16950 -5010
rect 17250 -4970 18350 -4965
rect 17250 -5010 17255 -4970
rect 17295 -5010 17605 -4970
rect 17645 -5010 17955 -4970
rect 17995 -5010 18305 -4970
rect 18345 -5010 18350 -4970
rect 17250 -5015 18350 -5010
rect 18650 -4970 19750 -4965
rect 18650 -5010 18655 -4970
rect 18695 -5010 19005 -4970
rect 19045 -5010 19355 -4970
rect 19395 -5010 19705 -4970
rect 19745 -5010 19750 -4970
rect 18650 -5015 19750 -5010
rect 16200 -5315 16250 -5015
rect 17950 -5315 18000 -5015
rect 19350 -5315 19400 -5015
rect 15850 -5320 16950 -5315
rect 15850 -5360 15855 -5320
rect 15895 -5360 16205 -5320
rect 16245 -5360 16555 -5320
rect 16595 -5360 16905 -5320
rect 16945 -5360 16950 -5320
rect 15850 -5365 16950 -5360
rect 17250 -5320 18350 -5315
rect 17250 -5360 17255 -5320
rect 17295 -5360 17605 -5320
rect 17645 -5360 17955 -5320
rect 17995 -5360 18305 -5320
rect 18345 -5360 18350 -5320
rect 17250 -5365 18350 -5360
rect 18650 -5320 19750 -5315
rect 18650 -5360 18655 -5320
rect 18695 -5360 19005 -5320
rect 19045 -5360 19355 -5320
rect 19395 -5360 19705 -5320
rect 19745 -5360 19750 -5320
rect 18650 -5365 19750 -5360
rect 16200 -5665 16250 -5365
rect 17950 -5665 18000 -5365
rect 19350 -5665 19400 -5365
rect 15850 -5670 16950 -5665
rect 15850 -5710 15855 -5670
rect 15895 -5710 16205 -5670
rect 16245 -5710 16555 -5670
rect 16595 -5710 16905 -5670
rect 16945 -5710 16950 -5670
rect 15850 -5715 16950 -5710
rect 17250 -5670 18350 -5665
rect 17250 -5710 17255 -5670
rect 17295 -5710 17605 -5670
rect 17645 -5710 17955 -5670
rect 17995 -5710 18305 -5670
rect 18345 -5710 18350 -5670
rect 17250 -5715 18350 -5710
rect 18650 -5670 19750 -5665
rect 18650 -5710 18655 -5670
rect 18695 -5710 19005 -5670
rect 19045 -5710 19355 -5670
rect 19395 -5710 19705 -5670
rect 19745 -5710 19750 -5670
rect 18650 -5715 19750 -5710
rect 16200 -6015 16250 -5715
rect 17950 -6015 18000 -5715
rect 19350 -6015 19400 -5715
rect 15850 -6020 16950 -6015
rect 15850 -6060 15855 -6020
rect 15895 -6060 16205 -6020
rect 16245 -6060 16555 -6020
rect 16595 -6060 16905 -6020
rect 16945 -6060 16950 -6020
rect 15850 -6065 16950 -6060
rect 17250 -6020 18350 -6015
rect 17250 -6060 17255 -6020
rect 17295 -6060 17605 -6020
rect 17645 -6060 17955 -6020
rect 17995 -6060 18305 -6020
rect 18345 -6060 18350 -6020
rect 17250 -6065 18350 -6060
rect 18650 -6020 19750 -6015
rect 18650 -6060 18655 -6020
rect 18695 -6060 19005 -6020
rect 19045 -6060 19355 -6020
rect 19395 -6060 19705 -6020
rect 19745 -6060 19750 -6020
rect 18650 -6065 19750 -6060
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel poly 18430 440 18430 440 5 FreeSans 400 0 0 -40 V_TOP
flabel metal2 15995 -4385 15995 -4385 5 FreeSans 400 0 0 -40 cap_res1
flabel metal3 19355 -4375 19355 -4375 7 FreeSans 400 180 -40 0 cap_res2
flabel metal1 16040 1585 16040 1585 7 FreeSans 240 0 -160 0 VB2_CUR_BIAS
port 11 w
flabel metal1 19415 1590 19415 1590 7 FreeSans 240 0 -160 0 ERR_AMP_REF
port 2 w
flabel metal1 19565 1590 19565 1590 3 FreeSans 240 0 160 0 VB3_CUR_BIAS
port 8 e
flabel via1 17800 1455 17800 1455 1 FreeSans 400 0 0 200 PFET_GATE_10uA
flabel metal1 16235 -1030 16235 -1030 3 FreeSans 400 0 200 0 START_UP
flabel metal1 18780 -1155 18780 -1155 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal1 16170 -1295 16170 -1295 7 FreeSans 400 0 -160 0 NFET_GATE_10uA
flabel metal2 18580 -745 18580 -745 3 FreeSans 400 180 200 0 V_p_2
flabel metal2 17060 -745 17060 -745 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 16670 -635 16670 -635 1 FreeSans 400 0 0 80 Vin+
flabel metal2 16665 -335 16665 -335 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 18930 -635 18930 -635 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 17570 -270 17570 -270 3 FreeSans 240 0 120 0 1st_Vout_1
flabel metal2 16620 -230 16620 -230 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 18030 -270 18030 -270 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 18980 -230 18980 -230 5 FreeSans 400 0 0 -40 V_mir2
flabel metal1 15805 1595 15805 1595 1 FreeSans 240 0 0 80 V_CMFB_S2
port 10 n
flabel metal1 17750 1595 17750 1595 1 FreeSans 240 0 0 80 TAIL_CUR_MIR_BIAS
port 5 n
flabel metal1 19795 1595 19795 1595 1 FreeSans 240 0 0 80 V_CMFB_S4
port 9 n
flabel metal1 16125 1595 16125 1595 1 FreeSans 240 0 0 80 ERR_AMP_CUR_BIAS
port 7 n
flabel metal1 19280 1590 19280 1590 1 FreeSans 240 0 0 80 VB1_CUR_BIAS
port 4 n
flabel metal1 18640 1595 18640 1595 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 16960 1595 16960 1595 1 FreeSans 240 0 0 80 V_CMFB_S1
port 6 n
<< end >>
