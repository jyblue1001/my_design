magic
tech sky130A
timestamp 1756311456
<< nwell >>
rect 2040 555 2220 575
rect 2060 540 2180 555
<< poly >>
rect -175 975 -135 985
rect -175 955 -165 975
rect -145 970 -135 975
rect -145 955 -90 970
rect -175 945 -135 955
rect 2180 940 2220 950
rect 2180 925 2190 940
rect 2090 920 2190 925
rect 2210 920 2220 940
rect 2090 910 2220 920
rect 3090 680 3130 690
rect 3090 660 3100 680
rect 3120 660 3130 680
rect 3090 650 3130 660
rect 3850 680 3890 690
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 3850 650 3890 660
rect 4070 490 4110 500
rect 4070 470 4080 490
rect 4100 470 4110 490
rect 4070 460 4110 470
rect -130 255 -90 265
rect -130 235 -120 255
rect -100 235 -90 255
rect -130 225 -90 235
rect 2075 80 2115 90
rect 2075 60 2085 80
rect 2105 60 2115 80
rect 2075 50 2115 60
rect 6010 -355 6050 -345
rect 6010 -375 6020 -355
rect 6040 -375 6050 -355
rect 6010 -385 6050 -375
rect 4965 -645 4985 -630
<< polycont >>
rect -165 955 -145 975
rect 2190 920 2210 940
rect 3100 660 3120 680
rect 3860 660 3880 680
rect 4080 470 4100 490
rect -120 235 -100 255
rect 2085 60 2105 80
rect 6020 -375 6040 -355
<< locali >>
rect 2775 2815 2825 2830
rect 2775 2795 2790 2815
rect 2810 2795 2825 2815
rect 2775 2780 2825 2795
rect 4820 2540 4860 2550
rect 4820 2520 4830 2540
rect 4850 2520 4860 2540
rect 4820 2510 4860 2520
rect 2775 2220 2825 2235
rect 2775 2200 2790 2220
rect 2810 2200 2825 2220
rect 2775 2185 2825 2200
rect 2380 1210 2430 1220
rect 2380 1205 2390 1210
rect 2355 1185 2390 1205
rect 2380 1180 2390 1185
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2030 1150 2070 1160
rect 2030 1130 2040 1150
rect 2060 1130 2070 1150
rect 2030 1120 2070 1130
rect 2040 1100 2060 1120
rect 2735 1015 2785 1030
rect 2735 995 2750 1015
rect 2770 995 2785 1015
rect -175 975 -135 985
rect 2735 980 2785 995
rect -175 955 -165 975
rect -145 955 -135 975
rect -175 945 -135 955
rect 2180 940 2220 950
rect 2180 920 2190 940
rect 2210 920 2220 940
rect 2180 910 2220 920
rect 2300 940 2340 950
rect 2300 920 2310 940
rect 2330 920 2340 940
rect 2300 910 2340 920
rect 3090 680 3130 690
rect 3090 660 3100 680
rect 3120 660 3130 680
rect 3850 680 3890 690
rect 3090 650 3130 660
rect 3155 635 3195 665
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 3850 650 3890 660
rect -190 620 -140 630
rect -190 590 -180 620
rect -150 615 -140 620
rect 2460 620 2510 635
rect 2460 615 2475 620
rect -150 595 -130 615
rect 2370 595 2400 615
rect 2420 600 2475 615
rect 2495 600 2510 620
rect 3155 615 3165 635
rect 3185 615 3195 635
rect 3155 605 3195 615
rect 2420 595 2510 600
rect -150 590 -140 595
rect -190 580 -140 590
rect 2460 585 2510 595
rect 4450 595 4490 605
rect 4450 575 4460 595
rect 4480 575 4490 595
rect 2040 555 2220 575
rect 4450 565 4490 575
rect 2040 505 2060 555
rect 2180 545 2220 555
rect 2180 525 2190 545
rect 2210 525 2220 545
rect 2180 515 2220 525
rect 4070 490 4110 500
rect 4070 470 4080 490
rect 4100 470 4110 490
rect 4070 460 4110 470
rect 2305 275 2345 285
rect -130 255 -90 265
rect -130 235 -120 255
rect -100 235 -90 255
rect 2305 255 2315 275
rect 2335 255 2345 275
rect 2305 245 2345 255
rect -130 225 -90 235
rect 2735 165 2785 180
rect 2735 145 2750 165
rect 2770 145 2785 165
rect 2735 130 2785 145
rect 2075 80 2115 90
rect 2075 60 2085 80
rect 2105 60 2115 80
rect 2075 50 2115 60
rect 2380 30 2430 40
rect 2380 25 2390 30
rect 2355 5 2390 25
rect 2380 0 2390 5
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 2380 -170 2430 -160
rect 2380 -200 2390 -170
rect 2420 -180 2430 -170
rect 7550 -180 7570 30
rect 2420 -200 2460 -180
rect 2480 -200 2510 -180
rect 2530 -200 2560 -180
rect 2580 -200 2610 -180
rect 2630 -200 2660 -180
rect 2680 -200 2710 -180
rect 2730 -200 2760 -180
rect 2780 -200 2810 -180
rect 2830 -200 2860 -180
rect 2880 -200 2910 -180
rect 2930 -200 2960 -180
rect 2980 -200 3010 -180
rect 3030 -200 3060 -180
rect 3080 -200 3110 -180
rect 3130 -200 3160 -180
rect 3180 -200 3210 -180
rect 3230 -200 3260 -180
rect 3280 -200 3310 -180
rect 3330 -200 3360 -180
rect 3380 -200 3410 -180
rect 3430 -200 3460 -180
rect 3480 -200 3510 -180
rect 3530 -200 3560 -180
rect 3580 -200 3610 -180
rect 3630 -200 3660 -180
rect 3680 -200 3710 -180
rect 3730 -200 3760 -180
rect 3780 -200 3810 -180
rect 3830 -200 3860 -180
rect 3880 -200 3910 -180
rect 3930 -200 3960 -180
rect 3980 -200 4010 -180
rect 4030 -200 4060 -180
rect 4080 -200 4110 -180
rect 4130 -200 4160 -180
rect 4180 -200 4210 -180
rect 4230 -200 4260 -180
rect 4280 -200 4310 -180
rect 4330 -200 4360 -180
rect 4380 -200 4410 -180
rect 4430 -200 4460 -180
rect 4480 -200 4510 -180
rect 4530 -200 4560 -180
rect 4580 -200 4610 -180
rect 4630 -200 4660 -180
rect 4680 -200 4710 -180
rect 4730 -200 4760 -180
rect 4780 -200 4810 -180
rect 4830 -200 4860 -180
rect 4880 -200 4910 -180
rect 4930 -200 4945 -180
rect 6180 -200 6210 -180
rect 6230 -200 6260 -180
rect 6280 -200 6310 -180
rect 6330 -200 6360 -180
rect 6380 -200 6410 -180
rect 6430 -200 6460 -180
rect 6480 -200 6510 -180
rect 6530 -200 6560 -180
rect 6580 -200 6610 -180
rect 6630 -200 6660 -180
rect 6680 -200 6710 -180
rect 6730 -200 6760 -180
rect 6780 -200 6810 -180
rect 6830 -200 6860 -180
rect 6880 -200 6910 -180
rect 6930 -200 6960 -180
rect 6980 -200 7010 -180
rect 7030 -200 7060 -180
rect 7080 -200 7110 -180
rect 7130 -200 7160 -180
rect 7180 -200 7210 -180
rect 7230 -200 7260 -180
rect 7280 -200 7310 -180
rect 7330 -200 7360 -180
rect 7380 -200 7410 -180
rect 7430 -200 7460 -180
rect 7480 -200 7510 -180
rect 7530 -200 7570 -180
rect 2380 -210 2430 -200
rect 6010 -355 6050 -345
rect 6010 -375 6020 -355
rect 6040 -375 6050 -355
rect 6010 -385 6050 -375
rect -335 -630 -295 -620
rect -335 -650 -325 -630
rect -305 -640 -295 -630
rect -305 -650 -280 -640
rect -335 -660 -280 -650
rect -330 -820 -280 -810
rect -330 -850 -320 -820
rect -290 -850 -280 -820
rect -330 -860 -280 -850
<< viali >>
rect 2790 2795 2810 2815
rect 4830 2520 4850 2540
rect 2790 2200 2810 2220
rect 2390 1180 2420 1210
rect 2040 1130 2060 1150
rect 2750 995 2770 1015
rect -165 955 -145 975
rect 2190 920 2210 940
rect 2310 920 2330 940
rect 3100 660 3120 680
rect 3860 660 3880 680
rect -180 590 -150 620
rect 2350 595 2370 615
rect 2400 595 2420 615
rect 2475 600 2495 620
rect 3165 615 3185 635
rect 4460 575 4480 595
rect 2190 525 2210 545
rect 3065 525 3085 545
rect 4080 470 4100 490
rect -120 235 -100 255
rect 2315 255 2335 275
rect 2750 145 2770 165
rect 2085 60 2105 80
rect 2390 0 2420 30
rect 2390 -200 2420 -170
rect 2460 -200 2480 -180
rect 2510 -200 2530 -180
rect 2560 -200 2580 -180
rect 2610 -200 2630 -180
rect 2660 -200 2680 -180
rect 2710 -200 2730 -180
rect 2760 -200 2780 -180
rect 2810 -200 2830 -180
rect 2860 -200 2880 -180
rect 2910 -200 2930 -180
rect 2960 -200 2980 -180
rect 3010 -200 3030 -180
rect 3060 -200 3080 -180
rect 3110 -200 3130 -180
rect 3160 -200 3180 -180
rect 3210 -200 3230 -180
rect 3260 -200 3280 -180
rect 3310 -200 3330 -180
rect 3360 -200 3380 -180
rect 3410 -200 3430 -180
rect 3460 -200 3480 -180
rect 3510 -200 3530 -180
rect 3560 -200 3580 -180
rect 3610 -200 3630 -180
rect 3660 -200 3680 -180
rect 3710 -200 3730 -180
rect 3760 -200 3780 -180
rect 3810 -200 3830 -180
rect 3860 -200 3880 -180
rect 3910 -200 3930 -180
rect 3960 -200 3980 -180
rect 4010 -200 4030 -180
rect 4060 -200 4080 -180
rect 4110 -200 4130 -180
rect 4160 -200 4180 -180
rect 4210 -200 4230 -180
rect 4260 -200 4280 -180
rect 4310 -200 4330 -180
rect 4360 -200 4380 -180
rect 4410 -200 4430 -180
rect 4460 -200 4480 -180
rect 4510 -200 4530 -180
rect 4560 -200 4580 -180
rect 4610 -200 4630 -180
rect 4660 -200 4680 -180
rect 4710 -200 4730 -180
rect 4760 -200 4780 -180
rect 4810 -200 4830 -180
rect 4860 -200 4880 -180
rect 4910 -200 4930 -180
rect 6160 -200 6180 -180
rect 6210 -200 6230 -180
rect 6260 -200 6280 -180
rect 6310 -200 6330 -180
rect 6360 -200 6380 -180
rect 6410 -200 6430 -180
rect 6460 -200 6480 -180
rect 6510 -200 6530 -180
rect 6560 -200 6580 -180
rect 6610 -200 6630 -180
rect 6660 -200 6680 -180
rect 6710 -200 6730 -180
rect 6760 -200 6780 -180
rect 6810 -200 6830 -180
rect 6860 -200 6880 -180
rect 6910 -200 6930 -180
rect 6960 -200 6980 -180
rect 7010 -200 7030 -180
rect 7060 -200 7080 -180
rect 7110 -200 7130 -180
rect 7160 -200 7180 -180
rect 7210 -200 7230 -180
rect 7260 -200 7280 -180
rect 7310 -200 7330 -180
rect 7360 -200 7380 -180
rect 7410 -200 7430 -180
rect 7460 -200 7480 -180
rect 7510 -200 7530 -180
rect 6020 -375 6040 -355
rect -325 -650 -305 -630
rect -320 -850 -290 -820
<< metal1 >>
rect 1825 6285 1905 6290
rect 1825 6255 1830 6285
rect 1860 6255 1870 6285
rect 1900 6255 1905 6285
rect 1825 6245 1905 6255
rect 1825 6215 1830 6245
rect 1860 6215 1870 6245
rect 1900 6215 1905 6245
rect 1825 6205 1905 6215
rect 1825 6175 1830 6205
rect 1860 6175 1870 6205
rect 1900 6175 1905 6205
rect 1825 3870 1905 6175
rect 1825 3840 1830 3870
rect 1860 3840 1870 3870
rect 1900 3840 1905 3870
rect 1825 3830 1905 3840
rect 1825 3800 1830 3830
rect 1860 3800 1870 3830
rect 1900 3800 1905 3830
rect 1825 3795 1905 3800
rect 2465 3315 2505 5475
rect 2460 3295 2510 3315
rect 2460 3265 2470 3295
rect 2500 3265 2510 3295
rect 2460 3245 2510 3265
rect 2460 3215 2470 3245
rect 2500 3215 2510 3245
rect 2460 3195 2510 3215
rect 2775 2820 2825 2830
rect 2775 2790 2785 2820
rect 2815 2790 2825 2820
rect 2775 2780 2825 2790
rect 2635 2595 2675 2600
rect 2635 2565 2640 2595
rect 2670 2565 2675 2595
rect 2635 2560 2675 2565
rect 2895 2590 2935 2595
rect 2895 2560 2900 2590
rect 2930 2560 2935 2590
rect 2580 2510 2620 2515
rect 2580 2480 2585 2510
rect 2615 2480 2620 2510
rect 2580 2475 2620 2480
rect -565 1345 -445 1350
rect -565 1315 -560 1345
rect -530 1315 -520 1345
rect -490 1315 -480 1345
rect -450 1315 -445 1345
rect -565 1305 -445 1315
rect -565 1275 -560 1305
rect -530 1275 -520 1305
rect -490 1275 -480 1305
rect -450 1275 -445 1305
rect -565 1265 -445 1275
rect -565 1235 -560 1265
rect -530 1235 -520 1265
rect -490 1235 -480 1265
rect -450 1235 -445 1265
rect -565 -30 -445 1235
rect 675 1345 715 1365
rect 675 1315 680 1345
rect 710 1315 715 1345
rect 675 1305 715 1315
rect 675 1275 680 1305
rect 710 1275 715 1305
rect 675 1265 715 1275
rect 675 1235 680 1265
rect 710 1235 715 1265
rect 675 1230 715 1235
rect 785 1345 825 1365
rect 785 1315 790 1345
rect 820 1315 825 1345
rect 785 1305 825 1315
rect 785 1275 790 1305
rect 820 1275 825 1305
rect 785 1265 825 1275
rect 785 1235 790 1265
rect 820 1235 825 1265
rect 785 1230 825 1235
rect 895 1345 935 1365
rect 895 1315 900 1345
rect 930 1315 935 1345
rect 895 1305 935 1315
rect 895 1275 900 1305
rect 930 1275 935 1305
rect 895 1265 935 1275
rect 895 1235 900 1265
rect 930 1235 935 1265
rect 895 1230 935 1235
rect 1005 1345 1045 1365
rect 1005 1315 1010 1345
rect 1040 1315 1045 1345
rect 1005 1305 1045 1315
rect 1005 1275 1010 1305
rect 1040 1275 1045 1305
rect 1005 1265 1045 1275
rect 1005 1235 1010 1265
rect 1040 1235 1045 1265
rect 1005 1230 1045 1235
rect 1115 1345 1155 1365
rect 1115 1315 1120 1345
rect 1150 1315 1155 1345
rect 1115 1305 1155 1315
rect 1115 1275 1120 1305
rect 1150 1275 1155 1305
rect 1115 1265 1155 1275
rect 1115 1235 1120 1265
rect 1150 1235 1155 1265
rect 1115 1230 1155 1235
rect 1225 1345 1265 1365
rect 1225 1315 1230 1345
rect 1260 1315 1265 1345
rect 2590 1340 2610 2475
rect 1225 1305 1265 1315
rect 1225 1275 1230 1305
rect 1260 1275 1265 1305
rect 2580 1335 2620 1340
rect 2580 1305 2585 1335
rect 2615 1305 2620 1335
rect 2580 1300 2620 1305
rect 1225 1265 1265 1275
rect 1225 1235 1230 1265
rect 1260 1235 1265 1265
rect 2535 1280 2575 1285
rect 2535 1250 2540 1280
rect 2570 1250 2575 1280
rect 2535 1245 2575 1250
rect 1225 1230 1265 1235
rect 2380 1215 2430 1220
rect 2355 1210 2430 1215
rect 2355 1180 2390 1210
rect 2420 1180 2430 1210
rect 2355 1175 2430 1180
rect 2380 1170 2430 1175
rect 2030 1155 2070 1160
rect 2030 1125 2035 1155
rect 2065 1125 2070 1155
rect 2030 1120 2070 1125
rect 2545 1095 2565 1245
rect 2580 1155 2620 1160
rect 2580 1125 2585 1155
rect 2615 1125 2620 1155
rect 2580 1120 2620 1125
rect 2180 1090 2220 1095
rect 2180 1060 2185 1090
rect 2215 1060 2220 1090
rect 2180 1055 2220 1060
rect 2535 1090 2575 1095
rect 2535 1060 2540 1090
rect 2570 1060 2575 1090
rect 2535 1055 2575 1060
rect -175 980 -135 985
rect -175 950 -170 980
rect -140 950 -135 980
rect 2190 950 2210 1055
rect -175 945 -135 950
rect 2180 945 2220 950
rect 2180 915 2185 945
rect 2215 915 2220 945
rect 2180 910 2220 915
rect 2300 945 2340 950
rect 2300 915 2305 945
rect 2335 915 2340 945
rect 2300 910 2340 915
rect 2535 945 2575 950
rect 2535 915 2540 945
rect 2570 915 2575 945
rect 2535 910 2575 915
rect -190 625 -140 630
rect 2460 625 2510 635
rect -190 620 -115 625
rect -190 590 -180 620
rect -150 590 -115 620
rect 2355 615 2470 625
rect 2370 595 2400 615
rect 2420 595 2470 615
rect 2500 595 2510 625
rect 2545 610 2565 910
rect 2590 690 2610 1120
rect 2580 685 2620 690
rect 2580 655 2585 685
rect 2615 655 2620 685
rect 2580 650 2620 655
rect 2645 645 2665 2560
rect 2895 2555 2935 2560
rect 4820 2540 4860 2550
rect 5975 2545 6015 2550
rect 5975 2540 5980 2545
rect 4820 2520 4830 2540
rect 4850 2525 5980 2540
rect 4850 2520 4860 2525
rect 2895 2510 2935 2515
rect 4820 2510 4860 2520
rect 5975 2515 5980 2525
rect 6010 2515 6015 2545
rect 5975 2510 6015 2515
rect 2895 2480 2900 2510
rect 2930 2480 2935 2510
rect 2895 2475 2935 2480
rect 2775 2225 2825 2235
rect 2775 2195 2785 2225
rect 2815 2195 2825 2225
rect 2775 2185 2825 2195
rect 2690 1390 2730 1395
rect 2690 1360 2695 1390
rect 2725 1360 2730 1390
rect 2690 1355 2730 1360
rect 5975 1385 6015 1390
rect 5975 1355 5980 1385
rect 6010 1355 6015 1385
rect 2700 690 2720 1355
rect 5975 1350 6015 1355
rect 5450 1335 5490 1340
rect 5450 1305 5455 1335
rect 5485 1305 5490 1335
rect 5450 1300 5490 1305
rect 2735 1020 2785 1030
rect 2735 990 2745 1020
rect 2775 990 2785 1020
rect 2735 980 2785 990
rect 2690 685 2730 690
rect 2690 655 2695 685
rect 2725 655 2730 685
rect 2690 650 2730 655
rect 3090 685 3130 690
rect 3090 655 3095 685
rect 3125 655 3130 685
rect 3090 650 3130 655
rect 3850 680 3890 690
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 2635 640 2675 645
rect 2635 610 2640 640
rect 2670 610 2675 640
rect -190 585 -115 590
rect 2355 585 2510 595
rect 2535 605 2575 610
rect 2635 605 2675 610
rect 3155 640 3195 645
rect 3155 610 3160 640
rect 3190 610 3195 640
rect 3155 605 3195 610
rect -190 580 -140 585
rect 2535 575 2540 605
rect 2570 575 2575 605
rect 2535 570 2575 575
rect 3850 595 3890 660
rect 5460 605 5480 1300
rect 3850 565 3855 595
rect 3885 565 3890 595
rect 4450 600 4490 605
rect 4450 570 4455 600
rect 4485 570 4490 600
rect 4450 565 4490 570
rect 5450 600 5490 605
rect 5450 570 5455 600
rect 5485 570 5490 600
rect 5450 565 5490 570
rect 3850 560 3890 565
rect 2180 550 2220 555
rect 2180 520 2185 550
rect 2215 520 2220 550
rect 2180 515 2220 520
rect 2495 550 2615 555
rect 2495 520 2500 550
rect 2530 520 2540 550
rect 2570 520 2580 550
rect 2610 520 2615 550
rect 2305 280 2345 285
rect -335 260 -295 265
rect -335 230 -330 260
rect -300 255 -295 260
rect -130 255 -90 265
rect -300 240 -120 255
rect -300 230 -295 240
rect -335 225 -295 230
rect -130 235 -120 240
rect -100 235 -90 255
rect 2305 250 2310 280
rect 2340 250 2345 280
rect 2305 245 2345 250
rect -130 225 -90 235
rect -565 -60 -560 -30
rect -530 -60 -520 -30
rect -490 -60 -480 -30
rect -450 -60 -445 -30
rect -565 -70 -445 -60
rect -565 -100 -560 -70
rect -530 -100 -520 -70
rect -490 -100 -480 -70
rect -450 -100 -445 -70
rect -565 -110 -445 -100
rect -565 -140 -560 -110
rect -530 -140 -520 -110
rect -490 -140 -480 -110
rect -450 -140 -445 -110
rect -565 -145 -445 -140
rect -325 -620 -305 225
rect 2075 85 2115 90
rect 2075 55 2080 85
rect 2110 55 2115 85
rect 2075 50 2115 55
rect 2380 35 2430 40
rect 2355 30 2430 35
rect 2355 0 2390 30
rect 2420 0 2430 30
rect 2355 -5 2430 0
rect 2380 -10 2430 -5
rect 2495 -30 2615 520
rect 3055 550 3095 555
rect 3055 520 3060 550
rect 3090 520 3095 550
rect 3055 515 3095 520
rect 4070 495 4110 500
rect 2735 490 2775 495
rect 2735 460 2740 490
rect 2770 460 2775 490
rect 4070 465 4075 495
rect 4105 465 4110 495
rect 4070 460 4110 465
rect 2735 455 2775 460
rect 2745 285 2765 455
rect 2735 280 2775 285
rect 2735 250 2740 280
rect 2770 250 2775 280
rect 2735 245 2775 250
rect 2735 170 2785 180
rect 2735 140 2745 170
rect 2775 140 2785 170
rect 2735 130 2785 140
rect 5460 0 5480 565
rect 2495 -60 2500 -30
rect 2530 -60 2540 -30
rect 2570 -60 2580 -30
rect 2610 -60 2615 -30
rect 5450 -5 5490 0
rect 5450 -35 5455 -5
rect 5485 -35 5490 -5
rect 5450 -40 5490 -35
rect 6010 -5 6065 0
rect 6010 -35 6015 -5
rect 6045 -15 6065 -5
rect 6045 -30 6115 -15
rect 6045 -35 6065 -30
rect 6010 -40 6065 -35
rect 2495 -70 2615 -60
rect 2495 -100 2500 -70
rect 2530 -100 2540 -70
rect 2570 -100 2580 -70
rect 2610 -100 2615 -70
rect 2495 -110 2615 -100
rect 2495 -140 2500 -110
rect 2530 -140 2540 -110
rect 2570 -140 2580 -110
rect 2610 -140 2615 -110
rect 2495 -145 2615 -140
rect 2380 -170 2430 -160
rect 2380 -200 2390 -170
rect 2420 -180 4945 -170
rect 6180 -180 7570 -170
rect 2420 -200 2460 -180
rect 2480 -200 2510 -180
rect 2530 -200 2560 -180
rect 2580 -200 2610 -180
rect 2630 -200 2660 -180
rect 2680 -200 2710 -180
rect 2730 -200 2760 -180
rect 2780 -200 2810 -180
rect 2830 -200 2860 -180
rect 2880 -200 2910 -180
rect 2930 -200 2960 -180
rect 2980 -200 3010 -180
rect 3030 -200 3060 -180
rect 3080 -200 3110 -180
rect 3130 -200 3160 -180
rect 3180 -200 3210 -180
rect 3230 -200 3260 -180
rect 3280 -200 3310 -180
rect 3330 -200 3360 -180
rect 3380 -200 3410 -180
rect 3430 -200 3460 -180
rect 3480 -200 3510 -180
rect 3530 -200 3560 -180
rect 3580 -200 3610 -180
rect 3630 -200 3660 -180
rect 3680 -200 3710 -180
rect 3730 -200 3760 -180
rect 3780 -200 3810 -180
rect 3830 -200 3860 -180
rect 3880 -200 3910 -180
rect 3930 -200 3960 -180
rect 3980 -200 4010 -180
rect 4030 -200 4060 -180
rect 4080 -200 4110 -180
rect 4130 -200 4160 -180
rect 4180 -200 4210 -180
rect 4230 -200 4260 -180
rect 4280 -200 4310 -180
rect 4330 -200 4360 -180
rect 4380 -200 4410 -180
rect 4430 -200 4460 -180
rect 4480 -200 4510 -180
rect 4530 -200 4560 -180
rect 4580 -200 4610 -180
rect 4630 -200 4660 -180
rect 4680 -200 4710 -180
rect 4730 -200 4760 -180
rect 4780 -200 4810 -180
rect 4830 -200 4860 -180
rect 4880 -200 4910 -180
rect 4930 -200 4945 -180
rect 6180 -200 6210 -180
rect 6230 -200 6260 -180
rect 6280 -200 6310 -180
rect 6330 -200 6360 -180
rect 6380 -200 6410 -180
rect 6430 -200 6460 -180
rect 6480 -200 6510 -180
rect 6530 -200 6560 -180
rect 6580 -200 6610 -180
rect 6630 -200 6660 -180
rect 6680 -200 6710 -180
rect 6730 -200 6760 -180
rect 6780 -200 6810 -180
rect 6830 -200 6860 -180
rect 6880 -200 6910 -180
rect 6930 -200 6960 -180
rect 6980 -200 7010 -180
rect 7030 -200 7060 -180
rect 7080 -200 7110 -180
rect 7130 -200 7160 -180
rect 7180 -200 7210 -180
rect 7230 -200 7260 -180
rect 7280 -200 7310 -180
rect 7330 -200 7360 -180
rect 7380 -200 7410 -180
rect 7430 -200 7460 -180
rect 7480 -200 7510 -180
rect 7530 -200 7570 -180
rect 2380 -210 4945 -200
rect 6180 -210 7570 -200
rect 6010 -350 6050 -345
rect 6010 -380 6015 -350
rect 6045 -380 6050 -350
rect 6010 -385 6050 -380
rect -335 -625 -295 -620
rect -335 -655 -330 -625
rect -300 -655 -295 -625
rect -335 -660 -295 -655
rect -330 -820 -280 -810
rect -330 -850 -320 -820
rect -290 -850 -280 -820
rect -330 -860 -280 -850
<< via1 >>
rect 1830 6255 1860 6285
rect 1870 6255 1900 6285
rect 1830 6215 1860 6245
rect 1870 6215 1900 6245
rect 1830 6175 1860 6205
rect 1870 6175 1900 6205
rect 1830 3840 1860 3870
rect 1870 3840 1900 3870
rect 1830 3800 1860 3830
rect 1870 3800 1900 3830
rect 2470 3265 2500 3295
rect 2470 3215 2500 3245
rect 2785 2815 2815 2820
rect 2785 2795 2790 2815
rect 2790 2795 2810 2815
rect 2810 2795 2815 2815
rect 2785 2790 2815 2795
rect 2640 2565 2670 2595
rect 2900 2560 2930 2590
rect 2585 2480 2615 2510
rect -560 1315 -530 1345
rect -520 1315 -490 1345
rect -480 1315 -450 1345
rect -560 1275 -530 1305
rect -520 1275 -490 1305
rect -480 1275 -450 1305
rect -560 1235 -530 1265
rect -520 1235 -490 1265
rect -480 1235 -450 1265
rect 680 1315 710 1345
rect 680 1275 710 1305
rect 680 1235 710 1265
rect 790 1315 820 1345
rect 790 1275 820 1305
rect 790 1235 820 1265
rect 900 1315 930 1345
rect 900 1275 930 1305
rect 900 1235 930 1265
rect 1010 1315 1040 1345
rect 1010 1275 1040 1305
rect 1010 1235 1040 1265
rect 1120 1315 1150 1345
rect 1120 1275 1150 1305
rect 1120 1235 1150 1265
rect 1230 1315 1260 1345
rect 1230 1275 1260 1305
rect 2585 1305 2615 1335
rect 1230 1235 1260 1265
rect 2540 1250 2570 1280
rect 2390 1180 2420 1210
rect 2035 1150 2065 1155
rect 2035 1130 2040 1150
rect 2040 1130 2060 1150
rect 2060 1130 2065 1150
rect 2035 1125 2065 1130
rect 2585 1125 2615 1155
rect 2185 1060 2215 1090
rect 2540 1060 2570 1090
rect -170 975 -140 980
rect -170 955 -165 975
rect -165 955 -145 975
rect -145 955 -140 975
rect -170 950 -140 955
rect 2185 940 2215 945
rect 2185 920 2190 940
rect 2190 920 2210 940
rect 2210 920 2215 940
rect 2185 915 2215 920
rect 2305 940 2335 945
rect 2305 920 2310 940
rect 2310 920 2330 940
rect 2330 920 2335 940
rect 2305 915 2335 920
rect 2540 915 2570 945
rect -180 590 -150 620
rect 2470 620 2500 625
rect 2470 600 2475 620
rect 2475 600 2495 620
rect 2495 600 2500 620
rect 2470 595 2500 600
rect 2585 655 2615 685
rect 5980 2515 6010 2545
rect 2900 2480 2930 2510
rect 2785 2220 2815 2225
rect 2785 2200 2790 2220
rect 2790 2200 2810 2220
rect 2810 2200 2815 2220
rect 2785 2195 2815 2200
rect 2695 1360 2725 1390
rect 5980 1355 6010 1385
rect 5455 1305 5485 1335
rect 2745 1015 2775 1020
rect 2745 995 2750 1015
rect 2750 995 2770 1015
rect 2770 995 2775 1015
rect 2745 990 2775 995
rect 2695 655 2725 685
rect 3095 680 3125 685
rect 3095 660 3100 680
rect 3100 660 3120 680
rect 3120 660 3125 680
rect 3095 655 3125 660
rect 2640 610 2670 640
rect 3160 635 3190 640
rect 3160 615 3165 635
rect 3165 615 3185 635
rect 3185 615 3190 635
rect 3160 610 3190 615
rect 2540 575 2570 605
rect 3855 565 3885 595
rect 4455 595 4485 600
rect 4455 575 4460 595
rect 4460 575 4480 595
rect 4480 575 4485 595
rect 4455 570 4485 575
rect 5455 570 5485 600
rect 2185 545 2215 550
rect 2185 525 2190 545
rect 2190 525 2210 545
rect 2210 525 2215 545
rect 2185 520 2215 525
rect 2500 520 2530 550
rect 2540 520 2570 550
rect 2580 520 2610 550
rect -330 230 -300 260
rect 2310 275 2340 280
rect 2310 255 2315 275
rect 2315 255 2335 275
rect 2335 255 2340 275
rect 2310 250 2340 255
rect -560 -60 -530 -30
rect -520 -60 -490 -30
rect -480 -60 -450 -30
rect -560 -100 -530 -70
rect -520 -100 -490 -70
rect -480 -100 -450 -70
rect -560 -140 -530 -110
rect -520 -140 -490 -110
rect -480 -140 -450 -110
rect 2080 80 2110 85
rect 2080 60 2085 80
rect 2085 60 2105 80
rect 2105 60 2110 80
rect 2080 55 2110 60
rect 2390 0 2420 30
rect 3060 545 3090 550
rect 3060 525 3065 545
rect 3065 525 3085 545
rect 3085 525 3090 545
rect 3060 520 3090 525
rect 2740 460 2770 490
rect 4075 490 4105 495
rect 4075 470 4080 490
rect 4080 470 4100 490
rect 4100 470 4105 490
rect 4075 465 4105 470
rect 2740 250 2770 280
rect 2745 165 2775 170
rect 2745 145 2750 165
rect 2750 145 2770 165
rect 2770 145 2775 165
rect 2745 140 2775 145
rect 2500 -60 2530 -30
rect 2540 -60 2570 -30
rect 2580 -60 2610 -30
rect 5455 -35 5485 -5
rect 6015 -35 6045 -5
rect 2500 -100 2530 -70
rect 2540 -100 2570 -70
rect 2580 -100 2610 -70
rect 2500 -140 2530 -110
rect 2540 -140 2570 -110
rect 2580 -140 2610 -110
rect 2390 -200 2420 -170
rect 6015 -355 6045 -350
rect 6015 -375 6020 -355
rect 6020 -375 6040 -355
rect 6040 -375 6045 -355
rect 6015 -380 6045 -375
rect -330 -630 -300 -625
rect -330 -650 -325 -630
rect -325 -650 -305 -630
rect -305 -650 -300 -630
rect -330 -655 -300 -650
rect -320 -850 -290 -820
<< metal2 >>
rect 1795 6285 1905 6290
rect 1795 6255 1830 6285
rect 1860 6255 1870 6285
rect 1900 6255 1905 6285
rect 1795 6245 1905 6255
rect 1795 6215 1830 6245
rect 1860 6215 1870 6245
rect 1900 6215 1905 6245
rect 1795 6205 1905 6215
rect 1795 6175 1830 6205
rect 1860 6175 1870 6205
rect 1900 6175 1905 6205
rect 1795 6170 1905 6175
rect 1630 3870 2430 3875
rect 1630 3840 1830 3870
rect 1860 3840 1870 3870
rect 1900 3850 2430 3870
rect 1900 3840 2390 3850
rect 1630 3830 2390 3840
rect 1630 3800 1830 3830
rect 1860 3800 1870 3830
rect 1900 3820 2390 3830
rect 2420 3820 2430 3850
rect 1900 3800 2430 3820
rect 1630 3795 2430 3800
rect 1185 3695 2430 3715
rect 1185 3665 2390 3695
rect 2420 3665 2430 3695
rect 1185 3645 2430 3665
rect 1185 3615 2390 3645
rect 2420 3615 2430 3645
rect 1185 3595 2430 3615
rect 1675 3295 2510 3315
rect 1675 3265 2470 3295
rect 2500 3265 2510 3295
rect 1675 3245 2510 3265
rect 1675 3215 2470 3245
rect 2500 3215 2510 3245
rect 1675 3195 2510 3215
rect 2775 2820 2825 2830
rect 2775 2790 2785 2820
rect 2815 2790 2825 2820
rect 2775 2780 2825 2790
rect 2635 2595 2675 2600
rect 2635 2565 2640 2595
rect 2670 2580 2675 2595
rect 2895 2590 2935 2595
rect 2895 2580 2900 2590
rect 2670 2565 2900 2580
rect 2635 2560 2675 2565
rect 2895 2560 2900 2565
rect 2930 2560 2935 2590
rect 2895 2555 2935 2560
rect 5975 2545 6015 2550
rect 5975 2515 5980 2545
rect 6010 2515 6015 2545
rect 2580 2510 2620 2515
rect 1875 2465 2510 2485
rect 2580 2480 2585 2510
rect 2615 2500 2620 2510
rect 2895 2510 2935 2515
rect 5975 2510 6015 2515
rect 2895 2500 2900 2510
rect 2615 2485 2900 2500
rect 2615 2480 2620 2485
rect 2580 2475 2620 2480
rect 2895 2480 2900 2485
rect 2930 2480 2935 2510
rect 2895 2475 2935 2480
rect 1875 2435 2470 2465
rect 2500 2435 2510 2465
rect 1875 2415 2510 2435
rect 1875 2385 2470 2415
rect 2500 2385 2510 2415
rect 1875 2365 2510 2385
rect 2775 2225 2825 2235
rect 2775 2195 2785 2225
rect 2815 2195 2825 2225
rect 2775 2185 2825 2195
rect 1860 1740 2510 1760
rect 1860 1710 2470 1740
rect 2500 1710 2510 1740
rect 1860 1690 2510 1710
rect 1860 1660 2470 1690
rect 2500 1660 2510 1690
rect 1860 1640 2510 1660
rect 2460 1460 2510 1465
rect 1860 1455 2510 1460
rect 1860 1425 2470 1455
rect 2500 1425 2510 1455
rect 1860 1420 2510 1425
rect 2460 1415 2510 1420
rect 2690 1390 2730 1395
rect 5985 1390 6000 2510
rect 2690 1360 2695 1390
rect 2725 1380 2730 1390
rect 5975 1385 6015 1390
rect 5975 1380 5980 1385
rect 2725 1365 5980 1380
rect 2725 1360 2730 1365
rect 2690 1355 2730 1360
rect 5975 1355 5980 1365
rect 6010 1355 6015 1385
rect 5975 1350 6015 1355
rect -565 1345 1265 1350
rect -565 1315 -560 1345
rect -530 1315 -520 1345
rect -490 1315 -480 1345
rect -450 1315 680 1345
rect 710 1315 790 1345
rect 820 1315 900 1345
rect 930 1315 1010 1345
rect 1040 1315 1120 1345
rect 1150 1315 1230 1345
rect 1260 1315 1265 1345
rect -565 1305 1265 1315
rect -565 1275 -560 1305
rect -530 1275 -520 1305
rect -490 1275 -480 1305
rect -450 1275 680 1305
rect 710 1275 790 1305
rect 820 1275 900 1305
rect 930 1275 1010 1305
rect 1040 1275 1120 1305
rect 1150 1275 1230 1305
rect 1260 1275 1265 1305
rect 2580 1335 2620 1340
rect 2580 1305 2585 1335
rect 2615 1330 2620 1335
rect 5450 1335 5490 1340
rect 5450 1330 5455 1335
rect 2615 1310 5455 1330
rect 2615 1305 2620 1310
rect 2580 1300 2620 1305
rect 5450 1305 5455 1310
rect 5485 1305 5490 1335
rect 5450 1300 5490 1305
rect -565 1265 1265 1275
rect -565 1235 -560 1265
rect -530 1235 -520 1265
rect -490 1235 -480 1265
rect -450 1235 680 1265
rect 710 1235 790 1265
rect 820 1235 900 1265
rect 930 1235 1010 1265
rect 1040 1235 1120 1265
rect 1150 1235 1230 1265
rect 1260 1235 1265 1265
rect 2535 1280 2575 1285
rect 2535 1250 2540 1280
rect 2570 1275 2575 1280
rect 2570 1260 2735 1275
rect 2570 1250 2575 1260
rect 2535 1245 2575 1250
rect -565 1230 1265 1235
rect 2380 1210 2430 1220
rect 2380 1180 2390 1210
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2030 1155 2070 1160
rect 2030 1125 2035 1155
rect 2065 1150 2070 1155
rect 2580 1155 2620 1160
rect 2580 1150 2585 1155
rect 2065 1130 2585 1150
rect 2065 1125 2070 1130
rect 2030 1120 2070 1125
rect 2580 1125 2585 1130
rect 2615 1125 2620 1155
rect 2580 1120 2620 1125
rect 2180 1090 2220 1095
rect 2180 1060 2185 1090
rect 2215 1085 2220 1090
rect 2535 1090 2575 1095
rect 2535 1085 2540 1090
rect 2215 1065 2540 1085
rect 2215 1060 2220 1065
rect 2180 1055 2220 1060
rect 2535 1060 2540 1065
rect 2570 1060 2575 1090
rect 2535 1055 2575 1060
rect 2735 1020 2785 1030
rect 2735 990 2745 1020
rect 2775 990 2785 1020
rect -1140 980 -135 985
rect 2735 980 2785 990
rect -1140 950 -170 980
rect -140 950 -135 980
rect -1140 945 -135 950
rect 2180 945 2220 950
rect 2180 915 2185 945
rect 2215 915 2220 945
rect 2180 910 2220 915
rect 2300 945 2340 950
rect 2300 915 2305 945
rect 2335 940 2340 945
rect 2535 945 2575 950
rect 2535 940 2540 945
rect 2335 920 2540 940
rect 2335 915 2340 920
rect 2300 910 2340 915
rect 2535 915 2540 920
rect 2570 915 2575 945
rect 2535 910 2575 915
rect 2580 685 2620 690
rect 2580 655 2585 685
rect 2615 680 2620 685
rect 2690 685 2730 690
rect 2690 680 2695 685
rect 2615 660 2695 680
rect 2615 655 2620 660
rect 2580 650 2620 655
rect 2690 655 2695 660
rect 2725 680 2730 685
rect 3090 685 3130 690
rect 3090 680 3095 685
rect 2725 660 3095 680
rect 2725 655 2730 660
rect 2690 650 2730 655
rect 3090 655 3095 660
rect 3125 655 3130 685
rect 3090 650 3130 655
rect 2635 640 2675 645
rect -190 620 -140 630
rect -190 590 -180 620
rect -150 590 -140 620
rect -190 580 -140 590
rect 2460 625 2510 635
rect 2460 595 2470 625
rect 2500 595 2510 625
rect 2635 610 2640 640
rect 2670 635 2675 640
rect 3155 640 3195 645
rect 3155 635 3160 640
rect 2670 615 3160 635
rect 2670 610 2675 615
rect 2460 585 2510 595
rect 2535 605 2575 610
rect 2635 605 2675 610
rect 3155 610 3160 615
rect 3190 610 3195 640
rect 3155 605 3195 610
rect 2535 575 2540 605
rect 2570 590 2575 605
rect 4450 600 4490 605
rect 3850 595 3890 600
rect 3850 590 3855 595
rect 2570 575 3855 590
rect 2535 570 3855 575
rect 3850 565 3855 570
rect 3885 565 3890 595
rect 4450 570 4455 600
rect 4485 595 4490 600
rect 5450 600 5490 605
rect 5450 595 5455 600
rect 4485 575 5455 595
rect 4485 570 4490 575
rect 4450 565 4490 570
rect 5450 570 5455 575
rect 5485 570 5490 600
rect 5450 565 5490 570
rect 3850 560 3890 565
rect 2180 550 3095 555
rect 2180 520 2185 550
rect 2215 520 2500 550
rect 2530 520 2540 550
rect 2570 520 2580 550
rect 2610 520 3060 550
rect 3090 520 3095 550
rect 2180 515 3095 520
rect 4070 495 4110 500
rect 2735 490 2775 495
rect 4070 490 4075 495
rect 2735 460 2740 490
rect 2770 470 4075 490
rect 2770 460 2775 470
rect 4070 465 4075 470
rect 4105 465 4110 495
rect 4070 460 4110 465
rect 2735 455 2775 460
rect 2305 280 2345 285
rect -335 260 -295 265
rect -335 230 -330 260
rect -300 230 -295 260
rect 2305 250 2310 280
rect 2340 275 2345 280
rect 2735 280 2775 285
rect 2735 275 2740 280
rect 2340 255 2740 275
rect 2340 250 2345 255
rect 2305 245 2345 250
rect 2735 250 2740 255
rect 2770 250 2775 280
rect 2735 245 2775 250
rect -335 225 -295 230
rect 2735 170 2785 180
rect 2735 140 2745 170
rect 2775 140 2785 170
rect 2735 130 2785 140
rect 2075 85 2115 90
rect 2075 55 2080 85
rect 2110 70 2740 85
rect 2110 55 2115 70
rect 2075 50 2115 55
rect 2380 30 2430 40
rect 2380 0 2390 30
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 5450 -5 5490 0
rect -565 -30 2615 -25
rect -565 -60 -560 -30
rect -530 -60 -520 -30
rect -490 -60 -480 -30
rect -450 -60 2500 -30
rect 2530 -60 2540 -30
rect 2570 -60 2580 -30
rect 2610 -60 2615 -30
rect 5450 -35 5455 -5
rect 5485 -10 5490 -5
rect 6010 -5 6065 0
rect 6010 -10 6015 -5
rect 5485 -30 6015 -10
rect 5485 -35 5490 -30
rect 5450 -40 5490 -35
rect 6010 -35 6015 -30
rect 6045 -35 6065 -5
rect 6010 -40 6065 -35
rect -565 -70 2615 -60
rect -565 -100 -560 -70
rect -530 -100 -520 -70
rect -490 -100 -480 -70
rect -450 -100 2500 -70
rect 2530 -100 2540 -70
rect 2570 -100 2580 -70
rect 2610 -100 2615 -70
rect -565 -110 2615 -100
rect -565 -140 -560 -110
rect -530 -140 -520 -110
rect -490 -140 -480 -110
rect -450 -140 2500 -110
rect 2530 -140 2540 -110
rect 2570 -140 2580 -110
rect 2610 -140 2615 -110
rect -565 -145 2615 -140
rect 2380 -170 2430 -160
rect 2380 -200 2390 -170
rect 2420 -200 2430 -170
rect 2380 -210 2430 -200
rect 6020 -345 6035 -40
rect 6010 -350 6050 -345
rect 6010 -380 6015 -350
rect 6045 -380 6050 -350
rect 6010 -385 6050 -380
rect -335 -625 -295 -620
rect -335 -655 -330 -625
rect -300 -655 -295 -625
rect -335 -660 -295 -655
rect -330 -820 -280 -810
rect -330 -850 -320 -820
rect -290 -850 -280 -820
rect -330 -860 -280 -850
<< via2 >>
rect 2390 3820 2420 3850
rect 2390 3665 2420 3695
rect 2390 3615 2420 3645
rect 2470 3265 2500 3295
rect 2470 3215 2500 3245
rect 2785 2790 2815 2820
rect 2470 2435 2500 2465
rect 2470 2385 2500 2415
rect 2785 2195 2815 2225
rect 2470 1710 2500 1740
rect 2470 1660 2500 1690
rect 2470 1425 2500 1455
rect 2390 1180 2420 1210
rect 2745 990 2775 1020
rect -180 590 -150 620
rect 2470 595 2500 625
rect 2745 140 2775 170
rect 2390 0 2420 30
rect 2390 -200 2420 -170
rect -320 -850 -290 -820
<< metal3 >>
rect 2380 3855 2430 3860
rect 2380 3815 2385 3855
rect 2425 3815 2430 3855
rect 2380 3810 2430 3815
rect 2380 3700 2430 3705
rect 2380 3660 2385 3700
rect 2425 3660 2430 3700
rect 2380 3650 2430 3660
rect 2380 3610 2385 3650
rect 2425 3610 2430 3650
rect 2380 3605 2430 3610
rect 2460 3300 2510 3305
rect 2460 3260 2465 3300
rect 2505 3260 2510 3300
rect 2460 3250 2510 3260
rect 2460 3210 2465 3250
rect 2505 3210 2510 3250
rect 2460 3205 2510 3210
rect 2380 2825 2825 2830
rect 2380 2785 2385 2825
rect 2425 2820 2825 2825
rect 2425 2790 2785 2820
rect 2815 2790 2825 2820
rect 2425 2785 2825 2790
rect 2380 2780 2825 2785
rect 2460 2470 2510 2475
rect 2460 2430 2465 2470
rect 2505 2430 2510 2470
rect 2460 2420 2510 2430
rect 2460 2380 2465 2420
rect 2505 2380 2510 2420
rect 2460 2375 2510 2380
rect 2460 2230 2825 2235
rect 2460 2190 2465 2230
rect 2505 2225 2825 2230
rect 2505 2195 2785 2225
rect 2815 2195 2825 2225
rect 2505 2190 2825 2195
rect 2460 2185 2825 2190
rect 2460 1745 2510 1750
rect 2460 1705 2465 1745
rect 2505 1705 2510 1745
rect 2460 1695 2510 1705
rect 2460 1655 2465 1695
rect 2505 1655 2510 1695
rect 2460 1650 2510 1655
rect 2460 1460 2510 1465
rect 2460 1420 2465 1460
rect 2505 1420 2510 1460
rect 2460 1415 2510 1420
rect 2380 1215 2430 1220
rect 2380 1175 2385 1215
rect 2425 1175 2430 1215
rect 2380 1170 2430 1175
rect 2460 1025 2785 1030
rect 2460 985 2465 1025
rect 2505 1020 2785 1025
rect 2505 990 2745 1020
rect 2775 990 2785 1020
rect 2505 985 2785 990
rect 2460 980 2785 985
rect 2460 630 2510 635
rect -430 625 -140 630
rect -430 585 -425 625
rect -385 620 -140 625
rect -385 590 -180 620
rect -150 590 -140 620
rect -385 585 -140 590
rect 2460 590 2465 630
rect 2505 590 2510 630
rect 2460 585 2510 590
rect -430 580 -140 585
rect 2380 175 2785 180
rect 2380 135 2385 175
rect 2425 170 2785 175
rect 2425 140 2745 170
rect 2775 140 2785 170
rect 2425 135 2785 140
rect 2380 130 2785 135
rect 2380 35 2430 40
rect 2380 -5 2385 35
rect 2425 -5 2430 35
rect 2380 -10 2430 -5
rect 2380 -165 2430 -160
rect 2380 -205 2385 -165
rect 2425 -205 2430 -165
rect 2380 -210 2430 -205
rect -430 -815 -280 -810
rect -430 -855 -425 -815
rect -385 -820 -280 -815
rect -385 -850 -320 -820
rect -290 -850 -280 -820
rect -385 -855 -280 -850
rect -430 -860 -280 -855
<< via3 >>
rect 2385 3850 2425 3855
rect 2385 3820 2390 3850
rect 2390 3820 2420 3850
rect 2420 3820 2425 3850
rect 2385 3815 2425 3820
rect 2385 3695 2425 3700
rect 2385 3665 2390 3695
rect 2390 3665 2420 3695
rect 2420 3665 2425 3695
rect 2385 3660 2425 3665
rect 2385 3645 2425 3650
rect 2385 3615 2390 3645
rect 2390 3615 2420 3645
rect 2420 3615 2425 3645
rect 2385 3610 2425 3615
rect 2465 3295 2505 3300
rect 2465 3265 2470 3295
rect 2470 3265 2500 3295
rect 2500 3265 2505 3295
rect 2465 3260 2505 3265
rect 2465 3245 2505 3250
rect 2465 3215 2470 3245
rect 2470 3215 2500 3245
rect 2500 3215 2505 3245
rect 2465 3210 2505 3215
rect 2385 2785 2425 2825
rect 2465 2465 2505 2470
rect 2465 2435 2470 2465
rect 2470 2435 2500 2465
rect 2500 2435 2505 2465
rect 2465 2430 2505 2435
rect 2465 2415 2505 2420
rect 2465 2385 2470 2415
rect 2470 2385 2500 2415
rect 2500 2385 2505 2415
rect 2465 2380 2505 2385
rect 2465 2190 2505 2230
rect 2465 1740 2505 1745
rect 2465 1710 2470 1740
rect 2470 1710 2500 1740
rect 2500 1710 2505 1740
rect 2465 1705 2505 1710
rect 2465 1690 2505 1695
rect 2465 1660 2470 1690
rect 2470 1660 2500 1690
rect 2500 1660 2505 1690
rect 2465 1655 2505 1660
rect 2465 1455 2505 1460
rect 2465 1425 2470 1455
rect 2470 1425 2500 1455
rect 2500 1425 2505 1455
rect 2465 1420 2505 1425
rect 2385 1210 2425 1215
rect 2385 1180 2390 1210
rect 2390 1180 2420 1210
rect 2420 1180 2425 1210
rect 2385 1175 2425 1180
rect 2465 985 2505 1025
rect -425 585 -385 625
rect 2465 625 2505 630
rect 2465 595 2470 625
rect 2470 595 2500 625
rect 2500 595 2505 625
rect 2465 590 2505 595
rect 2385 135 2425 175
rect 2385 30 2425 35
rect 2385 0 2390 30
rect 2390 0 2420 30
rect 2420 0 2425 30
rect 2385 -5 2425 0
rect 2385 -170 2425 -165
rect 2385 -200 2390 -170
rect 2390 -200 2420 -170
rect 2420 -200 2425 -170
rect 2385 -205 2425 -200
rect -425 -855 -385 -815
<< metal4 >>
rect 2380 3855 2430 3875
rect 2380 3815 2385 3855
rect 2425 3815 2430 3855
rect 2380 3700 2430 3815
rect 2380 3660 2385 3700
rect 2425 3660 2430 3700
rect 2380 3650 2430 3660
rect 2380 3610 2385 3650
rect 2425 3610 2430 3650
rect 2380 2825 2430 3610
rect 2380 2785 2385 2825
rect 2425 2785 2430 2825
rect 2380 1215 2430 2785
rect 2380 1175 2385 1215
rect 2425 1175 2430 1215
rect -430 625 -380 630
rect -430 585 -425 625
rect -385 585 -380 625
rect -430 -815 -380 585
rect 2380 175 2430 1175
rect 2460 3300 2510 3315
rect 2460 3260 2465 3300
rect 2505 3260 2510 3300
rect 2460 3250 2510 3260
rect 2460 3210 2465 3250
rect 2505 3210 2510 3250
rect 2460 2470 2510 3210
rect 2460 2430 2465 2470
rect 2505 2430 2510 2470
rect 2460 2420 2510 2430
rect 2460 2380 2465 2420
rect 2505 2380 2510 2420
rect 2460 2230 2510 2380
rect 2460 2190 2465 2230
rect 2505 2190 2510 2230
rect 2460 1745 2510 2190
rect 2460 1705 2465 1745
rect 2505 1705 2510 1745
rect 2460 1695 2510 1705
rect 2460 1655 2465 1695
rect 2505 1655 2510 1695
rect 2460 1460 2510 1655
rect 2460 1420 2465 1460
rect 2505 1420 2510 1460
rect 2460 1025 2510 1420
rect 2460 985 2465 1025
rect 2505 985 2510 1025
rect 2460 630 2510 985
rect 2460 590 2465 630
rect 2505 590 2510 630
rect 2460 585 2510 590
rect -280 100 -230 150
rect 2380 135 2385 175
rect 2425 135 2430 175
rect 2380 35 2430 135
rect 2380 -5 2385 35
rect 2425 -5 2430 35
rect 2380 -165 2430 -5
rect 2380 -205 2385 -165
rect 2425 -205 2430 -165
rect 2380 -210 2430 -205
rect -430 -855 -425 -815
rect -385 -855 -380 -815
rect -430 -860 -380 -855
use bgr  bgr_0
timestamp 1756256667
transform -1 0 18295 0 -1 2015
box 12350 -4330 19435 650
use charge_pump_cell_6  charge_pump_cell_6_0
timestamp 1756257297
transform 1 0 -6370 0 1 -1565
box 9105 1615 11630 2860
use loop_filter_2  loop_filter_2_0
timestamp 1740116583
transform 1 0 4930 0 -1 290
box 1135 -5975 9720 330
use opamp_cell_4  opamp_cell_4_0
timestamp 1740145811
transform 1 0 -425 0 -1 4625
box 3110 897 6365 3205
use pfd_8  pfd_8_0
timestamp 1739770731
transform 1 0 -930 0 1 4650
box 650 -4655 3290 -3435
use VCO_FD_magic  VCO_FD_magic_0
timestamp 1740284885
transform -1 0 6180 0 -1 -110
box 0 60 6470 1150
<< labels >>
flabel metal1 5480 985 5480 985 3 FreeSans 400 0 200 0 V_CONT
flabel poly 4975 -630 4975 -630 1 FreeSans 400 0 0 200 V_OSC
port 1 n
flabel poly -130 245 -130 245 7 FreeSans 400 0 -200 0 F_VCO
flabel metal1 -140 605 -140 605 7 FreeSans 400 0 -200 0 VDDA
port 2 w
flabel metal4 -280 125 -280 125 7 FreeSans 400 0 -200 0 GNDA
port 3 w
flabel poly -130 960 -130 960 7 FreeSans 400 0 -200 0 F_REF
port 4 w
flabel metal1 2615 -85 2615 -85 3 FreeSans 800 0 400 0 BGR_CURRENT_OUT
<< end >>
