* NGSPICE file created from loop_filter.ext - technology: sky130A

**.subckt loop_filter
X0 GNDA V_OUT sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X1 GNDA a_7952_500# sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X2 V_OUT a_7952_500# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=7.52
.ends

