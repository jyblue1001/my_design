* PEX produced on Thu Aug  7 12:54:54 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_18.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_18 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VOUT-.t19 two_stage_opamp_dummy_magic_25_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 VDDA.t241 two_stage_opamp_dummy_magic_25_0.Vb3.t8 two_stage_opamp_dummy_magic_25_0.VD4.t25 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X2 VDDA.t239 two_stage_opamp_dummy_magic_25_0.Vb3.t9 two_stage_opamp_dummy_magic_25_0.VD3.t31 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X3 VOUT+.t19 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_25_0.VD3.t37 two_stage_opamp_dummy_magic_25_0.Vb2.t11 two_stage_opamp_dummy_magic_25_0.X.t15 two_stage_opamp_dummy_magic_25_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X5 GNDA.t248 GNDA.t246 two_stage_opamp_dummy_magic_25_0.Vb2.t6 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 VOUT-.t20 two_stage_opamp_dummy_magic_25_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 two_stage_opamp_dummy_magic_25_0.VD2.t16 VIN+.t0 two_stage_opamp_dummy_magic_25_0.V_source.t13 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X8 VOUT-.t21 two_stage_opamp_dummy_magic_25_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 bgr_11_0.V_mir2.t11 bgr_11_0.V_mir2.t10 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X10 two_stage_opamp_dummy_magic_25_0.V_source.t11 two_stage_opamp_dummy_magic_25_0.Vb1.t12 two_stage_opamp_dummy_magic_25_0.Vb1_2.t4 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X11 VOUT+.t17 two_stage_opamp_dummy_magic_25_0.Y.t25 VDDA.t387 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X12 bgr_11_0.V_TOP.t14 VDDA.t147 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 GNDA.t285 VDDA.t356 VDDA.t358 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X14 GNDA.t3 a_6470_28110.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X15 GNDA.t331 two_stage_opamp_dummy_magic_25_0.Y.t26 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t10 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X16 VOUT-.t22 two_stage_opamp_dummy_magic_25_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 GNDA.t294 bgr_11_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t2 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X18 VDDA.t121 two_stage_opamp_dummy_magic_25_0.Y.t27 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t12 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X19 VOUT+.t20 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 two_stage_opamp_dummy_magic_25_0.Vb2.t5 GNDA.t243 GNDA.t245 GNDA.t244 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X21 VOUT-.t23 two_stage_opamp_dummy_magic_25_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t408 bgr_11_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t16 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X23 bgr_11_0.V_TOP.t15 VDDA.t148 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t15 VDDA.t353 VDDA.t355 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X25 VOUT-.t24 two_stage_opamp_dummy_magic_25_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 bgr_11_0.1st_Vout_1.t6 bgr_11_0.V_mir1.t13 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X27 VDDA.t237 two_stage_opamp_dummy_magic_25_0.Vb3.t10 two_stage_opamp_dummy_magic_25_0.VD4.t28 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X28 two_stage_opamp_dummy_magic_25_0.V_err_gate.t4 VDDA.t350 VDDA.t352 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X29 two_stage_opamp_dummy_magic_25_0.V_err_p.t2 two_stage_opamp_dummy_magic_25_0.V_tot.t4 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t0 VDDA.t364 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X30 two_stage_opamp_dummy_magic_25_0.VD1.t9 two_stage_opamp_dummy_magic_25_0.Vb1.t13 two_stage_opamp_dummy_magic_25_0.X.t18 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X31 VOUT-.t25 two_stage_opamp_dummy_magic_25_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 a_12070_29568.t0 bgr_11_0.V_CUR_REF_REG.t0 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=4
X33 two_stage_opamp_dummy_magic_25_0.VD3.t33 VDDA.t347 VDDA.t349 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X34 two_stage_opamp_dummy_magic_25_0.VD2.t3 two_stage_opamp_dummy_magic_25_0.Vb1.t14 two_stage_opamp_dummy_magic_25_0.Y.t9 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X35 bgr_11_0.1st_Vout_2.t7 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VOUT-.t1 two_stage_opamp_dummy_magic_25_0.X.t25 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X37 two_stage_opamp_dummy_magic_25_0.VD1.t8 two_stage_opamp_dummy_magic_25_0.Vb1.t15 two_stage_opamp_dummy_magic_25_0.X.t19 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X38 VOUT+.t21 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT-.t2 two_stage_opamp_dummy_magic_25_0.X.t26 VDDA.t49 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X40 GNDA.t122 two_stage_opamp_dummy_magic_25_0.X.t27 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t10 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X41 two_stage_opamp_dummy_magic_25_0.V_err_gate.t1 bgr_11_0.NFET_GATE_10uA.t6 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X42 bgr_11_0.V_TOP.t6 bgr_11_0.1st_Vout_1.t7 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X43 VDDA.t235 two_stage_opamp_dummy_magic_25_0.Vb3.t11 two_stage_opamp_dummy_magic_25_0.VD4.t27 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X44 GNDA.t242 GNDA.t240 VDDA.t50 GNDA.t241 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X45 VOUT+.t22 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 VOUT-.t26 two_stage_opamp_dummy_magic_25_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VOUT-.t27 two_stage_opamp_dummy_magic_25_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT-.t28 two_stage_opamp_dummy_magic_25_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VOUT-.t29 two_stage_opamp_dummy_magic_25_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VDDA.t367 two_stage_opamp_dummy_magic_25_0.X.t28 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t12 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X51 VOUT-.t30 two_stage_opamp_dummy_magic_25_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VOUT+.t23 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 bgr_11_0.START_UP.t3 bgr_11_0.V_TOP.t16 VDDA.t419 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X54 VDDA.t346 VDDA.t344 two_stage_opamp_dummy_magic_25_0.V_err_gate.t3 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X55 VOUT+.t24 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 VDDA.t343 VDDA.t341 VDDA.t343 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X57 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t1 GNDA.t237 GNDA.t239 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X58 two_stage_opamp_dummy_magic_25_0.VD1.t16 VIN-.t0 two_stage_opamp_dummy_magic_25_0.V_source.t26 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X59 VDDA.t156 bgr_11_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t10 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X60 VOUT+.t25 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 bgr_11_0.V_TOP.t12 bgr_11_0.1st_Vout_1.t8 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X62 VOUT+.t26 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 two_stage_opamp_dummy_magic_25_0.VD3.t17 two_stage_opamp_dummy_magic_25_0.Vb2.t12 two_stage_opamp_dummy_magic_25_0.X.t14 two_stage_opamp_dummy_magic_25_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X64 bgr_11_0.1st_Vout_2.t8 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 two_stage_opamp_dummy_magic_25_0.VD2.t18 GNDA.t234 GNDA.t236 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X66 two_stage_opamp_dummy_magic_25_0.Vb1.t5 two_stage_opamp_dummy_magic_25_0.Vb1.t4 two_stage_opamp_dummy_magic_25_0.Vb1_2.t3 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X67 a_5700_29568.t0 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t0 GNDA.t46 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X68 VOUT+.t27 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 bgr_11_0.V_TOP.t17 VDDA.t420 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 GNDA.t292 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_25_0.V_source.t33 GNDA.t291 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X71 two_stage_opamp_dummy_magic_25_0.X.t13 two_stage_opamp_dummy_magic_25_0.Vb2.t13 two_stage_opamp_dummy_magic_25_0.VD3.t35 two_stage_opamp_dummy_magic_25_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X72 VOUT+.t15 VDDA.t338 VDDA.t340 VDDA.t339 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X73 GNDA.t233 GNDA.t231 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t2 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X74 two_stage_opamp_dummy_magic_25_0.VD1.t12 VIN-.t1 two_stage_opamp_dummy_magic_25_0.V_source.t2 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X75 VOUT-.t31 two_stage_opamp_dummy_magic_25_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t14 bgr_11_0.PFET_GATE_10uA.t12 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X77 VOUT+.t6 two_stage_opamp_dummy_magic_25_0.Y.t28 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X78 bgr_11_0.1st_Vout_1.t9 bgr_11_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 GNDA.t8 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t2 VOUT+.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X80 two_stage_opamp_dummy_magic_25_0.VD4.t12 two_stage_opamp_dummy_magic_25_0.Vb2.t14 two_stage_opamp_dummy_magic_25_0.Y.t19 two_stage_opamp_dummy_magic_25_0.VD4.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X81 GNDA.t74 two_stage_opamp_dummy_magic_25_0.Y.t29 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t9 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X82 VOUT-.t32 two_stage_opamp_dummy_magic_25_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VDDA.t233 two_stage_opamp_dummy_magic_25_0.Vb3.t12 two_stage_opamp_dummy_magic_25_0.VD4.t26 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X84 VOUT-.t33 two_stage_opamp_dummy_magic_25_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT-.t34 two_stage_opamp_dummy_magic_25_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 two_stage_opamp_dummy_magic_25_0.V_source.t6 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t13 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X87 VOUT+.t28 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 bgr_11_0.V_TOP.t13 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t7 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X89 GNDA.t284 VDDA.t421 bgr_11_0.V_p_2.t2 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X90 VOUT+.t29 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VOUT+.t30 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 VDDA.t337 VDDA.t335 bgr_11_0.V_TOP.t11 VDDA.t336 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X93 VOUT+.t31 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 bgr_11_0.V_mir1.t12 bgr_11_0.V_mir1.t11 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X95 two_stage_opamp_dummy_magic_25_0.Vb2_2.t8 two_stage_opamp_dummy_magic_25_0.Vb2_2.t6 two_stage_opamp_dummy_magic_25_0.Vb2_2.t8 two_stage_opamp_dummy_magic_25_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X96 two_stage_opamp_dummy_magic_25_0.V_p_mir.t1 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t14 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X97 two_stage_opamp_dummy_magic_25_0.VD3.t30 two_stage_opamp_dummy_magic_25_0.Vb3.t13 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X98 bgr_11_0.V_TOP.t10 VDDA.t332 VDDA.t334 VDDA.t333 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X99 two_stage_opamp_dummy_magic_25_0.VD1.t7 two_stage_opamp_dummy_magic_25_0.Vb1.t16 two_stage_opamp_dummy_magic_25_0.X.t22 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X100 VOUT-.t35 two_stage_opamp_dummy_magic_25_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 GNDA.t230 GNDA.t228 VOUT+.t4 GNDA.t229 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X102 VOUT+.t32 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 bgr_11_0.V_TOP.t18 VDDA.t391 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VOUT-.t36 two_stage_opamp_dummy_magic_25_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 GNDA.t296 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_25_0.V_source.t34 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X106 VOUT-.t37 two_stage_opamp_dummy_magic_25_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT-.t38 two_stage_opamp_dummy_magic_25_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VOUT+.t33 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VDDA.t331 VDDA.t329 GNDA.t278 VDDA.t330 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X110 two_stage_opamp_dummy_magic_25_0.VD2.t0 two_stage_opamp_dummy_magic_25_0.Vb1.t17 two_stage_opamp_dummy_magic_25_0.Y.t8 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X111 VOUT-.t39 two_stage_opamp_dummy_magic_25_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT-.t40 two_stage_opamp_dummy_magic_25_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT-.t7 two_stage_opamp_dummy_magic_25_0.X.t29 VDDA.t100 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X114 VDDA.t393 bgr_11_0.V_TOP.t19 bgr_11_0.Vin+.t5 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X115 two_stage_opamp_dummy_magic_25_0.VD1.t6 two_stage_opamp_dummy_magic_25_0.Vb1.t18 two_stage_opamp_dummy_magic_25_0.X.t20 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X116 VOUT-.t41 two_stage_opamp_dummy_magic_25_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 GNDA.t116 two_stage_opamp_dummy_magic_25_0.X.t30 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t9 VDDA.t403 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X118 VDDA.t16 bgr_11_0.V_mir2.t13 bgr_11_0.1st_Vout_2.t5 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X119 VOUT+.t34 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT+.t35 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 VOUT+.t36 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT+.t37 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 bgr_11_0.1st_Vout_2.t9 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 bgr_11_0.V_mir1.t10 bgr_11_0.V_mir1.t9 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X125 two_stage_opamp_dummy_magic_25_0.Y.t24 two_stage_opamp_dummy_magic_25_0.VD4.t32 two_stage_opamp_dummy_magic_25_0.VD4.t34 two_stage_opamp_dummy_magic_25_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X126 VDDA.t30 GNDA.t225 GNDA.t227 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X127 two_stage_opamp_dummy_magic_25_0.VD4.t19 two_stage_opamp_dummy_magic_25_0.Vb3.t14 VDDA.t229 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X128 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_25_0.V_err_gate.t6 VDDA.t398 VDDA.t397 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X129 VOUT+.t38 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 two_stage_opamp_dummy_magic_25_0.X.t12 two_stage_opamp_dummy_magic_25_0.Vb2.t15 two_stage_opamp_dummy_magic_25_0.VD3.t21 two_stage_opamp_dummy_magic_25_0.VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X131 two_stage_opamp_dummy_magic_25_0.VD3.t29 two_stage_opamp_dummy_magic_25_0.Vb3.t15 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X132 two_stage_opamp_dummy_magic_25_0.VD1.t17 VIN-.t2 two_stage_opamp_dummy_magic_25_0.V_source.t27 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X133 bgr_11_0.PFET_GATE_10uA.t8 VDDA.t326 VDDA.t328 VDDA.t327 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X134 VOUT-.t42 two_stage_opamp_dummy_magic_25_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 VOUT+.t39 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 VOUT-.t43 two_stage_opamp_dummy_magic_25_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 VOUT+.t40 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VOUT+.t41 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 a_6350_29718.t1 bgr_11_0.Vin+.t1 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X140 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t6 bgr_11_0.V_TOP.t20 VDDA.t415 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X141 VOUT-.t44 two_stage_opamp_dummy_magic_25_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 VOUT-.t45 two_stage_opamp_dummy_magic_25_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 two_stage_opamp_dummy_magic_25_0.Vb1.t1 two_stage_opamp_dummy_magic_25_0.Vb1.t0 two_stage_opamp_dummy_magic_25_0.Vb1_2.t2 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 two_stage_opamp_dummy_magic_25_0.VD1.t13 VIN-.t3 two_stage_opamp_dummy_magic_25_0.V_source.t9 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X145 VOUT+.t2 two_stage_opamp_dummy_magic_25_0.Y.t30 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X146 VOUT+.t42 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT+.t43 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT-.t46 two_stage_opamp_dummy_magic_25_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t44 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 bgr_11_0.1st_Vout_2.t10 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 VDDA.t301 VDDA.t299 two_stage_opamp_dummy_magic_25_0.Vb1.t11 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X152 VDDA.t44 bgr_11_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t9 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X153 GNDA.t287 bgr_11_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_25_0.Vb3.t5 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X154 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t8 bgr_11_0.PFET_GATE_10uA.t14 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X155 a_13840_3288.t0 two_stage_opamp_dummy_magic_25_0.V_tot.t2 GNDA.t70 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X156 VDDA.t123 bgr_11_0.V_mir2.t8 bgr_11_0.V_mir2.t9 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X157 VOUT+.t45 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 GNDA.t224 GNDA.t222 two_stage_opamp_dummy_magic_25_0.VD1.t15 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X159 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 GNDA.t221 GNDA.t219 two_stage_opamp_dummy_magic_25_0.V_source.t24 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X161 GNDA.t134 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_25_0.V_source.t22 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X162 VOUT-.t47 two_stage_opamp_dummy_magic_25_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VOUT-.t48 two_stage_opamp_dummy_magic_25_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VOUT-.t49 two_stage_opamp_dummy_magic_25_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT+.t46 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VDDA.t417 bgr_11_0.V_TOP.t21 bgr_11_0.START_UP.t2 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X167 VOUT+.t47 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 bgr_11_0.Vin-.t4 bgr_11_0.V_TOP.t22 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X169 VOUT+.t48 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VDDA.t225 two_stage_opamp_dummy_magic_25_0.Vb3.t16 two_stage_opamp_dummy_magic_25_0.VD3.t28 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X171 bgr_11_0.1st_Vout_1.t10 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 GNDA.t218 GNDA.t216 two_stage_opamp_dummy_magic_25_0.VD2.t17 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X173 VOUT+.t49 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 two_stage_opamp_dummy_magic_25_0.V_source.t30 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t17 GNDA.t270 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X175 VOUT-.t50 two_stage_opamp_dummy_magic_25_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VDDA.t325 VDDA.t323 VOUT+.t14 VDDA.t324 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X177 VOUT+.t50 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VOUT+.t9 GNDA.t213 GNDA.t215 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X179 two_stage_opamp_dummy_magic_25_0.Y.t18 two_stage_opamp_dummy_magic_25_0.Vb2.t16 two_stage_opamp_dummy_magic_25_0.VD4.t14 two_stage_opamp_dummy_magic_25_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X180 VOUT+.t51 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT+.t52 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 bgr_11_0.1st_Vout_2.t6 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t0 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X184 two_stage_opamp_dummy_magic_25_0.VD4.t22 two_stage_opamp_dummy_magic_25_0.Vb3.t17 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X185 VOUT+.t53 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VOUT+.t54 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 VOUT+.t55 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X189 VOUT-.t5 two_stage_opamp_dummy_magic_25_0.X.t31 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X190 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X191 two_stage_opamp_dummy_magic_25_0.VD1.t5 two_stage_opamp_dummy_magic_25_0.Vb1.t19 two_stage_opamp_dummy_magic_25_0.X.t24 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X192 VDDA.t187 bgr_11_0.1st_Vout_2.t12 bgr_11_0.PFET_GATE_10uA.t5 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X193 GNDA.t277 VDDA.t320 VDDA.t322 VDDA.t321 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X194 VOUT-.t51 two_stage_opamp_dummy_magic_25_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT+.t56 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT-.t52 two_stage_opamp_dummy_magic_25_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VOUT-.t53 two_stage_opamp_dummy_magic_25_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 VOUT-.t54 two_stage_opamp_dummy_magic_25_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 GNDA.t31 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_25_0.Vb2.t1 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X200 two_stage_opamp_dummy_magic_25_0.X.t11 two_stage_opamp_dummy_magic_25_0.Vb2.t17 two_stage_opamp_dummy_magic_25_0.VD3.t7 two_stage_opamp_dummy_magic_25_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X201 VOUT+.t57 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 two_stage_opamp_dummy_magic_25_0.X.t21 two_stage_opamp_dummy_magic_25_0.Vb1.t20 two_stage_opamp_dummy_magic_25_0.VD1.t4 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X203 VOUT-.t55 two_stage_opamp_dummy_magic_25_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VOUT+.t10 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t3 GNDA.t100 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X205 VOUT+.t58 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT-.t56 two_stage_opamp_dummy_magic_25_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT+.t59 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 bgr_11_0.V_TOP.t23 VDDA.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 two_stage_opamp_dummy_magic_25_0.Vb2.t9 bgr_11_0.NFET_GATE_10uA.t9 GNDA.t314 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X210 VOUT-.t57 two_stage_opamp_dummy_magic_25_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 bgr_11_0.NFET_GATE_10uA.t3 bgr_11_0.PFET_GATE_10uA.t15 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X213 two_stage_opamp_dummy_magic_25_0.Vb1.t10 GNDA.t210 GNDA.t212 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X214 two_stage_opamp_dummy_magic_25_0.Y.t17 two_stage_opamp_dummy_magic_25_0.Vb2.t18 two_stage_opamp_dummy_magic_25_0.VD4.t2 two_stage_opamp_dummy_magic_25_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X215 two_stage_opamp_dummy_magic_25_0.Y.t7 two_stage_opamp_dummy_magic_25_0.Vb1.t21 two_stage_opamp_dummy_magic_25_0.VD2.t19 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X216 VOUT+.t60 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 two_stage_opamp_dummy_magic_25_0.VD4.t21 two_stage_opamp_dummy_magic_25_0.Vb3.t18 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X218 two_stage_opamp_dummy_magic_25_0.VD1.t14 GNDA.t207 GNDA.t209 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X219 bgr_11_0.V_TOP.t24 VDDA.t145 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 bgr_11_0.1st_Vout_1.t5 bgr_11_0.V_mir1.t14 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X221 VOUT-.t58 two_stage_opamp_dummy_magic_25_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT-.t59 two_stage_opamp_dummy_magic_25_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT-.t60 two_stage_opamp_dummy_magic_25_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 GNDA.t206 GNDA.t204 VDDA.t129 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X225 VDDA.t219 two_stage_opamp_dummy_magic_25_0.Vb3.t19 two_stage_opamp_dummy_magic_25_0.VD3.t27 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X226 bgr_11_0.NFET_GATE_10uA.t1 bgr_11_0.NFET_GATE_10uA.t0 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X227 VOUT-.t61 two_stage_opamp_dummy_magic_25_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VOUT-.t62 two_stage_opamp_dummy_magic_25_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 a_3690_3288.t1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t13 GNDA.t124 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X230 VOUT+.t61 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 bgr_11_0.V_TOP.t25 VDDA.t146 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_11_0.Vin+.t0 GNDA.t97 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X233 VOUT-.t63 two_stage_opamp_dummy_magic_25_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 a_13960_3288.t1 two_stage_opamp_dummy_magic_25_0.V_tot.t3 GNDA.t86 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X235 VOUT+.t62 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VOUT-.t64 two_stage_opamp_dummy_magic_25_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 two_stage_opamp_dummy_magic_25_0.V_source.t12 VIN+.t1 two_stage_opamp_dummy_magic_25_0.VD2.t15 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X238 bgr_11_0.V_TOP.t26 VDDA.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDDA.t134 bgr_11_0.V_mir2.t6 bgr_11_0.V_mir2.t7 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X240 VDDA.t8 bgr_11_0.V_mir1.t7 bgr_11_0.V_mir1.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X241 VOUT-.t12 VDDA.t317 VDDA.t319 VDDA.t318 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X242 two_stage_opamp_dummy_magic_25_0.X.t10 two_stage_opamp_dummy_magic_25_0.Vb2.t19 two_stage_opamp_dummy_magic_25_0.VD3.t19 two_stage_opamp_dummy_magic_25_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X243 VOUT+.t63 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_25_0.Y.t31 VDDA.t385 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X245 two_stage_opamp_dummy_magic_25_0.VD4.t8 two_stage_opamp_dummy_magic_25_0.Vb2.t20 two_stage_opamp_dummy_magic_25_0.Y.t16 two_stage_opamp_dummy_magic_25_0.VD4.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X246 bgr_11_0.V_TOP.t27 VDDA.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 a_11420_29718.t1 bgr_11_0.Vin-.t5 GNDA.t325 sky130_fd_pr__res_xhigh_po_0p35 l=6
X248 VOUT-.t65 two_stage_opamp_dummy_magic_25_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 GNDA.t307 a_11950_28360.t1 GNDA.t306 sky130_fd_pr__res_xhigh_po_0p35 l=4
X250 VDDA.t217 two_stage_opamp_dummy_magic_25_0.Vb3.t20 two_stage_opamp_dummy_magic_25_0.VD3.t26 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X251 VOUT-.t66 two_stage_opamp_dummy_magic_25_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 VOUT-.t67 two_stage_opamp_dummy_magic_25_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VOUT+.t64 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 two_stage_opamp_dummy_magic_25_0.VD3.t15 two_stage_opamp_dummy_magic_25_0.VD3.t13 two_stage_opamp_dummy_magic_25_0.X.t4 two_stage_opamp_dummy_magic_25_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X255 VOUT+.t65 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VOUT+.t66 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 VOUT+.t67 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 two_stage_opamp_dummy_magic_25_0.err_amp_out.t3 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t5 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X260 VOUT+.t68 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 VOUT+.t69 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 bgr_11_0.1st_Vout_1.t13 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 two_stage_opamp_dummy_magic_25_0.Vb2.t2 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t53 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X264 bgr_11_0.1st_Vout_2.t14 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 GNDA.t203 GNDA.t201 VOUT-.t8 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X266 two_stage_opamp_dummy_magic_25_0.Y.t6 two_stage_opamp_dummy_magic_25_0.Vb1.t22 two_stage_opamp_dummy_magic_25_0.VD2.t21 GNDA.t333 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X267 two_stage_opamp_dummy_magic_25_0.Y.t5 two_stage_opamp_dummy_magic_25_0.Vb1.t23 two_stage_opamp_dummy_magic_25_0.VD2.t6 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X268 VDDA.t164 bgr_11_0.1st_Vout_2.t15 bgr_11_0.PFET_GATE_10uA.t4 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X269 VOUT-.t68 two_stage_opamp_dummy_magic_25_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VOUT+.t70 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 VOUT-.t69 two_stage_opamp_dummy_magic_25_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 VDDA.t316 VDDA.t314 GNDA.t276 VDDA.t315 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X273 VOUT-.t70 two_stage_opamp_dummy_magic_25_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 VOUT+.t71 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t1 bgr_11_0.NFET_GATE_10uA.t11 GNDA.t261 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X276 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t11 two_stage_opamp_dummy_magic_25_0.X.t32 VDDA.t196 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X277 VOUT+.t72 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 bgr_11_0.1st_Vout_2.t16 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VDDA.t313 VDDA.t311 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t14 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X280 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_25_0.X.t33 VDDA.t85 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X281 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t0 bgr_11_0.PFET_GATE_10uA.t16 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X282 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VOUT-.t71 two_stage_opamp_dummy_magic_25_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 bgr_11_0.V_TOP.t28 VDDA.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 bgr_11_0.V_mir1.t0 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t1 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X287 VDDA.t105 bgr_11_0.V_TOP.t29 bgr_11_0.START_UP.t1 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X288 two_stage_opamp_dummy_magic_25_0.V_source.t19 VIN+.t2 two_stage_opamp_dummy_magic_25_0.VD2.t14 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X289 VDDA.t142 bgr_11_0.V_mir2.t14 bgr_11_0.1st_Vout_2.t4 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X290 two_stage_opamp_dummy_magic_25_0.VD4.t6 two_stage_opamp_dummy_magic_25_0.Vb2.t21 two_stage_opamp_dummy_magic_25_0.Y.t15 two_stage_opamp_dummy_magic_25_0.VD4.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X291 VOUT-.t72 two_stage_opamp_dummy_magic_25_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t1 GNDA.t198 GNDA.t200 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X293 two_stage_opamp_dummy_magic_25_0.Vb3.t6 two_stage_opamp_dummy_magic_25_0.Vb2.t22 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X294 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_25_0.Y.t32 GNDA.t18 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X295 VOUT-.t73 two_stage_opamp_dummy_magic_25_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 two_stage_opamp_dummy_magic_25_0.cap_res_X.t138 two_stage_opamp_dummy_magic_25_0.X.t23 GNDA.t332 sky130_fd_pr__res_high_po_1p41 l=1.41
X297 VOUT+.t73 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VOUT-.t74 two_stage_opamp_dummy_magic_25_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 VOUT+.t74 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT-.t75 two_stage_opamp_dummy_magic_25_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 GNDA.t197 GNDA.t194 GNDA.t196 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X302 VOUT+.t75 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_25_0.Y.t33 VDDA.t120 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X304 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_25_0.Y.t34 VDDA.t169 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X305 VOUT+.t76 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 VOUT+.t77 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 two_stage_opamp_dummy_magic_25_0.VD3.t1 two_stage_opamp_dummy_magic_25_0.Vb2.t23 two_stage_opamp_dummy_magic_25_0.X.t9 two_stage_opamp_dummy_magic_25_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X308 VDDA.t160 bgr_11_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t7 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X309 VOUT+.t78 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 GNDA.t145 GNDA.t193 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X311 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t6 bgr_11_0.PFET_GATE_10uA.t18 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X312 two_stage_opamp_dummy_magic_25_0.err_amp_out.t1 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_25_0.V_err_p.t3 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X313 bgr_11_0.V_TOP.t30 VDDA.t388 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VOUT+.t79 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 GNDA.t145 GNDA.t192 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X316 VOUT-.t76 two_stage_opamp_dummy_magic_25_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_25_0.VD4.t10 two_stage_opamp_dummy_magic_25_0.Vb2.t24 two_stage_opamp_dummy_magic_25_0.Y.t14 two_stage_opamp_dummy_magic_25_0.VD4.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X318 VDDA.t310 VDDA.t308 two_stage_opamp_dummy_magic_25_0.VD4.t37 VDDA.t309 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X319 VOUT-.t77 two_stage_opamp_dummy_magic_25_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 two_stage_opamp_dummy_magic_25_0.Y.t4 two_stage_opamp_dummy_magic_25_0.Vb1.t24 two_stage_opamp_dummy_magic_25_0.VD2.t2 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X321 two_stage_opamp_dummy_magic_25_0.V_source.t36 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t18 GNDA.t302 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X322 bgr_11_0.cap_res1.t0 bgr_11_0.V_TOP.t1 GNDA.t67 sky130_fd_pr__res_high_po_0p35 l=2.05
X323 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t13 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 VDDA.t58 bgr_11_0.V_mir2.t4 bgr_11_0.V_mir2.t5 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X325 VDDA.t40 bgr_11_0.PFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t12 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 VOUT+.t80 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VOUT-.t78 two_stage_opamp_dummy_magic_25_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT-.t18 GNDA.t189 GNDA.t191 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X329 VDDA.t307 VDDA.t305 VOUT-.t0 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X330 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_25_0.X.t34 GNDA.t117 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X331 VDDA.t304 VDDA.t302 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t16 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X332 VOUT+.t81 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 two_stage_opamp_dummy_magic_25_0.VD3.t25 two_stage_opamp_dummy_magic_25_0.Vb3.t21 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X334 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_25_0.X.t35 GNDA.t118 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X335 GNDA.t272 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_25_0.V_source.t31 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X336 bgr_11_0.Vin-.t6 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t3 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X337 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_25_0.X.t36 VDDA.t47 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X338 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t5 bgr_11_0.V_TOP.t31 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X339 VOUT+.t82 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VOUT-.t79 two_stage_opamp_dummy_magic_25_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VOUT-.t80 two_stage_opamp_dummy_magic_25_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 GNDA.t145 GNDA.t146 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X343 VOUT-.t81 two_stage_opamp_dummy_magic_25_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 VOUT-.t82 two_stage_opamp_dummy_magic_25_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VOUT+.t83 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VDDA.t5 bgr_11_0.V_mir1.t15 bgr_11_0.1st_Vout_1.t4 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X347 VOUT+.t84 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 bgr_11_0.V_p_2.t1 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t8 bgr_11_0.V_mir2.t12 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X349 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t10 VDDA.t296 VDDA.t298 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X350 VOUT-.t83 two_stage_opamp_dummy_magic_25_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VOUT-.t14 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t4 GNDA.t269 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X352 bgr_11_0.START_UP.t5 bgr_11_0.START_UP.t4 bgr_11_0.START_UP_NFET1.t0 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X353 two_stage_opamp_dummy_magic_25_0.V_source.t21 VIN+.t3 two_stage_opamp_dummy_magic_25_0.VD2.t13 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X354 VOUT-.t84 two_stage_opamp_dummy_magic_25_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VOUT-.t85 two_stage_opamp_dummy_magic_25_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 two_stage_opamp_dummy_magic_25_0.VD3.t9 two_stage_opamp_dummy_magic_25_0.Vb2.t25 two_stage_opamp_dummy_magic_25_0.X.t8 two_stage_opamp_dummy_magic_25_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X357 VDDA.t152 two_stage_opamp_dummy_magic_25_0.Y.t35 VOUT+.t11 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X358 VOUT+.t85 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT+.t86 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 GNDA.t20 a_11300_28110.t1 GNDA.t19 sky130_fd_pr__res_xhigh_po_0p35 l=6
X361 VOUT+.t87 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 VOUT+.t88 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_25_0.Y.t36 GNDA.t319 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X365 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t0 a_13940_n584.t1 GNDA.t310 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X366 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_25_0.Y.t37 GNDA.t330 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X367 VDDA.t295 VDDA.t293 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t2 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X368 two_stage_opamp_dummy_magic_25_0.VD3.t24 two_stage_opamp_dummy_magic_25_0.Vb3.t22 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X369 VOUT+.t89 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_25_0.Y.t38 VDDA.t119 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X371 VOUT+.t90 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VDDA.t292 VDDA.t290 bgr_11_0.V_TOP.t9 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X373 VOUT-.t86 two_stage_opamp_dummy_magic_25_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 VOUT-.t87 two_stage_opamp_dummy_magic_25_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_25_0.V_err_gate.t2 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X377 VOUT+.t91 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VOUT-.t88 two_stage_opamp_dummy_magic_25_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 VDDA.t42 two_stage_opamp_dummy_magic_25_0.V_err_gate.t7 two_stage_opamp_dummy_magic_25_0.V_err_p.t1 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X380 VOUT+.t92 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 VOUT+.t93 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VOUT-.t89 two_stage_opamp_dummy_magic_25_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VOUT-.t90 two_stage_opamp_dummy_magic_25_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VDDA.t78 bgr_11_0.1st_Vout_1.t17 bgr_11_0.V_TOP.t2 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X386 VOUT+.t94 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VOUT+.t95 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 two_stage_opamp_dummy_magic_25_0.Y.t3 two_stage_opamp_dummy_magic_25_0.Vb1.t25 two_stage_opamp_dummy_magic_25_0.VD2.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X389 VDDA.t98 two_stage_opamp_dummy_magic_25_0.X.t37 VOUT-.t6 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X390 a_5700_29568.t1 a_5820_28304.t0 GNDA.t46 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X391 VDDA.t405 bgr_11_0.V_TOP.t32 bgr_11_0.Vin-.t3 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X392 VOUT+.t96 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 VDDA.t150 two_stage_opamp_dummy_magic_25_0.X.t38 VOUT-.t10 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X394 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_25_0.X.t39 GNDA.t104 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X395 VOUT-.t91 two_stage_opamp_dummy_magic_25_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 two_stage_opamp_dummy_magic_25_0.Vb1.t8 bgr_11_0.PFET_GATE_10uA.t21 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X397 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t5 bgr_11_0.PFET_GATE_10uA.t22 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X398 VOUT-.t92 two_stage_opamp_dummy_magic_25_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 GNDA.t188 GNDA.t186 two_stage_opamp_dummy_magic_25_0.Vb3.t7 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X400 VOUT-.t93 two_stage_opamp_dummy_magic_25_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_25_0.X.t40 VDDA.t29 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X402 VOUT-.t94 two_stage_opamp_dummy_magic_25_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 GNDA.t300 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t3 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t4 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X405 VOUT+.t97 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 two_stage_opamp_dummy_magic_25_0.V_source.t1 VIN-.t4 two_stage_opamp_dummy_magic_25_0.VD1.t11 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X407 VOUT+.t98 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 bgr_11_0.V_TOP.t33 VDDA.t406 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 two_stage_opamp_dummy_magic_25_0.V_source.t23 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t20 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X410 VDDA.t195 bgr_11_0.V_mir1.t5 bgr_11_0.V_mir1.t6 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X411 two_stage_opamp_dummy_magic_25_0.Y.t13 two_stage_opamp_dummy_magic_25_0.Vb2.t26 two_stage_opamp_dummy_magic_25_0.VD4.t4 two_stage_opamp_dummy_magic_25_0.VD4.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X412 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_25_0.Vb3.t0 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X413 bgr_11_0.1st_Vout_1.t19 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VDDA.t52 bgr_11_0.1st_Vout_1.t20 bgr_11_0.V_TOP.t0 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X415 VOUT+.t99 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT-.t95 two_stage_opamp_dummy_magic_25_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 two_stage_opamp_dummy_magic_25_0.V_source.t14 VIN+.t4 two_stage_opamp_dummy_magic_25_0.VD2.t12 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X418 GNDA.t185 GNDA.t183 two_stage_opamp_dummy_magic_25_0.Vb1.t9 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X419 GNDA.t72 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t21 two_stage_opamp_dummy_magic_25_0.V_source.t8 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X420 VOUT+.t100 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VDDA.t74 two_stage_opamp_dummy_magic_25_0.Y.t39 VOUT+.t5 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X422 two_stage_opamp_dummy_magic_25_0.V_source.t28 VIN-.t5 two_stage_opamp_dummy_magic_25_0.VD1.t18 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X423 VDDA.t82 two_stage_opamp_dummy_magic_25_0.Y.t40 VOUT+.t7 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X424 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_25_0.Y.t41 GNDA.t318 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X425 VOUT+.t101 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT-.t96 two_stage_opamp_dummy_magic_25_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VOUT-.t97 two_stage_opamp_dummy_magic_25_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 GNDA.t132 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_25_0.V_p_mir.t0 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X429 VOUT-.t98 two_stage_opamp_dummy_magic_25_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 bgr_11_0.PFET_GATE_10uA.t3 bgr_11_0.1st_Vout_2.t19 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X431 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_25_0.Y.t42 VDDA.t13 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X432 VOUT+.t102 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VOUT-.t99 two_stage_opamp_dummy_magic_25_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+.t103 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT-.t100 two_stage_opamp_dummy_magic_25_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 bgr_11_0.Vin-.t2 bgr_11_0.V_TOP.t34 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X437 VOUT+.t104 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 bgr_11_0.V_TOP.t35 VDDA.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VOUT+.t105 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT+.t106 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_25_0.V_source.t25 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t23 GNDA.t253 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X442 GNDA.t180 GNDA.t178 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t14 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X443 GNDA.t145 GNDA.t181 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X444 VDDA.t158 bgr_11_0.V_mir1.t3 bgr_11_0.V_mir1.t4 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X445 two_stage_opamp_dummy_magic_25_0.Y.t12 two_stage_opamp_dummy_magic_25_0.Vb2.t27 two_stage_opamp_dummy_magic_25_0.VD4.t18 two_stage_opamp_dummy_magic_25_0.VD4.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X446 two_stage_opamp_dummy_magic_25_0.X.t0 two_stage_opamp_dummy_magic_25_0.Vb1.t26 two_stage_opamp_dummy_magic_25_0.VD1.t3 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X447 VOUT-.t101 two_stage_opamp_dummy_magic_25_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t2 VDDA.t287 VDDA.t289 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X449 VOUT+.t107 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 bgr_11_0.V_TOP.t36 VDDA.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 GNDA.t145 GNDA.t182 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X452 GNDA.t14 bgr_11_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t2 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X453 VDDA.t10 bgr_11_0.1st_Vout_2.t20 bgr_11_0.PFET_GATE_10uA.t0 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X454 GNDA.t66 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_25_0.V_source.t7 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X455 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t284 VDDA.t286 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X456 VOUT+.t108 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 a_6350_29718.t0 a_6470_28110.t1 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X458 VDDA.t113 bgr_11_0.PFET_GATE_10uA.t23 bgr_11_0.V_CUR_REF_REG.t1 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X459 VOUT+.t109 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 bgr_11_0.1st_Vout_2.t21 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VDDA.t211 two_stage_opamp_dummy_magic_25_0.Vb3.t23 two_stage_opamp_dummy_magic_25_0.VD3.t23 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X462 two_stage_opamp_dummy_magic_25_0.Y.t22 GNDA.t175 GNDA.t177 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X463 VDDA.t72 two_stage_opamp_dummy_magic_25_0.X.t41 VOUT-.t4 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X464 two_stage_opamp_dummy_magic_25_0.X.t17 two_stage_opamp_dummy_magic_25_0.Vb1.t27 two_stage_opamp_dummy_magic_25_0.VD1.t2 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X465 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_25_0.X.t42 GNDA.t113 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X466 VOUT-.t102 two_stage_opamp_dummy_magic_25_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 VOUT-.t103 two_stage_opamp_dummy_magic_25_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 VDDA.t118 two_stage_opamp_dummy_magic_25_0.Y.t43 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t6 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X469 VOUT+.t110 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT-.t104 two_stage_opamp_dummy_magic_25_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT+.t111 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t7 two_stage_opamp_dummy_magic_25_0.X.t43 VDDA.t95 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X475 VOUT+.t3 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t5 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X476 GNDA.t24 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_25_0.V_err_gate.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X477 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t1 a_3830_n584.t1 GNDA.t324 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X478 VDDA.t366 bgr_11_0.V_mir2.t15 bgr_11_0.1st_Vout_2.t3 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X479 VDDA.t209 two_stage_opamp_dummy_magic_25_0.Vb3.t24 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t9 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X480 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_25_0.Y.t20 GNDA.t126 sky130_fd_pr__res_high_po_1p41 l=1.41
X481 two_stage_opamp_dummy_magic_25_0.V_err_gate.t5 two_stage_opamp_dummy_magic_25_0.V_tot.t5 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t2 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X482 two_stage_opamp_dummy_magic_25_0.V_source.t0 VIN-.t6 two_stage_opamp_dummy_magic_25_0.VD1.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X483 VOUT-.t105 two_stage_opamp_dummy_magic_25_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 GNDA.t145 GNDA.t167 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X485 VOUT+.t112 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT-.t106 two_stage_opamp_dummy_magic_25_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VOUT+.t113 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 a_12070_29568.t1 a_11950_28360.t0 GNDA.t68 sky130_fd_pr__res_xhigh_po_0p35 l=4
X490 a_3810_3288.t0 two_stage_opamp_dummy_magic_25_0.V_tot.t1 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X491 VOUT+.t114 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 a_13840_3288.t1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t14 GNDA.t323 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X494 two_stage_opamp_dummy_magic_25_0.Vb1_2.t1 two_stage_opamp_dummy_magic_25_0.Vb1.t2 two_stage_opamp_dummy_magic_25_0.Vb1.t3 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X495 VDDA.t283 VDDA.t281 two_stage_opamp_dummy_magic_25_0.VD3.t32 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X496 two_stage_opamp_dummy_magic_25_0.V_source.t18 VIN+.t5 two_stage_opamp_dummy_magic_25_0.VD2.t11 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X497 VOUT-.t107 two_stage_opamp_dummy_magic_25_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t11 VIN-.t7 two_stage_opamp_dummy_magic_25_0.V_p_mir.t3 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X499 two_stage_opamp_dummy_magic_25_0.V_source.t38 VIN-.t8 two_stage_opamp_dummy_magic_25_0.VD1.t21 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X500 VDDA.t93 bgr_11_0.V_TOP.t37 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t4 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X501 VDDA.t168 two_stage_opamp_dummy_magic_25_0.Y.t44 VOUT+.t13 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X502 VOUT-.t108 two_stage_opamp_dummy_magic_25_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 two_stage_opamp_dummy_magic_25_0.Vb3.t1 bgr_11_0.NFET_GATE_10uA.t14 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X504 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_25_0.Y.t45 GNDA.t35 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X505 VOUT+.t115 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 VOUT-.t109 two_stage_opamp_dummy_magic_25_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT-.t110 two_stage_opamp_dummy_magic_25_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT+.t116 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 bgr_11_0.1st_Vout_2.t24 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 two_stage_opamp_dummy_magic_25_0.V_source.t40 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t25 GNDA.t338 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X512 VOUT+.t117 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 bgr_11_0.V_mir2.t3 bgr_11_0.V_mir2.t2 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X514 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 bgr_11_0.1st_Vout_2.t25 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 GNDA.t41 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_25_0.V_source.t4 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X517 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t1 bgr_11_0.NFET_GATE_10uA.t15 GNDA.t252 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X518 two_stage_opamp_dummy_magic_25_0.X.t16 two_stage_opamp_dummy_magic_25_0.Vb1.t28 two_stage_opamp_dummy_magic_25_0.VD1.t1 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X519 GNDA.t335 bgr_11_0.NFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t0 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X520 GNDA.t174 GNDA.t171 GNDA.t173 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X521 VOUT-.t111 two_stage_opamp_dummy_magic_25_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VOUT+.t118 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 GNDA.t6 two_stage_opamp_dummy_magic_25_0.Y.t46 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t3 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X524 VOUT+.t119 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VDDA.t376 two_stage_opamp_dummy_magic_25_0.X.t44 VOUT-.t16 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X526 two_stage_opamp_dummy_magic_25_0.X.t5 two_stage_opamp_dummy_magic_25_0.Vb1.t29 two_stage_opamp_dummy_magic_25_0.VD1.t0 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X527 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_25_0.X.t45 GNDA.t105 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X528 two_stage_opamp_dummy_magic_25_0.Vb2.t0 bgr_11_0.NFET_GATE_10uA.t17 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X529 VDDA.t80 bgr_11_0.V_mir1.t16 bgr_11_0.1st_Vout_1.t3 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X530 GNDA.t136 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_25_0.Vb2.t8 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X531 VOUT-.t112 two_stage_opamp_dummy_magic_25_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t12 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X533 VOUT+.t120 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VDDA.t179 bgr_11_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t13 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X535 two_stage_opamp_dummy_magic_25_0.VD4.t16 two_stage_opamp_dummy_magic_25_0.Vb2.t28 two_stage_opamp_dummy_magic_25_0.Y.t11 two_stage_opamp_dummy_magic_25_0.VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X536 bgr_11_0.V_TOP.t38 VDDA.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VDDA.t181 two_stage_opamp_dummy_magic_25_0.V_err_gate.t8 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t0 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X538 GNDA.t170 GNDA.t168 two_stage_opamp_dummy_magic_25_0.X.t2 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X539 VOUT-.t113 two_stage_opamp_dummy_magic_25_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VOUT+.t121 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 bgr_11_0.V_TOP.t39 VDDA.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VOUT-.t114 two_stage_opamp_dummy_magic_25_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VOUT-.t115 two_stage_opamp_dummy_magic_25_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VOUT-.t116 two_stage_opamp_dummy_magic_25_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 two_stage_opamp_dummy_magic_25_0.Vb1_2.t0 two_stage_opamp_dummy_magic_25_0.Vb1.t6 two_stage_opamp_dummy_magic_25_0.Vb1.t7 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X546 GNDA.t166 GNDA.t164 two_stage_opamp_dummy_magic_25_0.Y.t21 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X547 VOUT-.t117 two_stage_opamp_dummy_magic_25_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 VDDA.t207 two_stage_opamp_dummy_magic_25_0.Vb3.t25 two_stage_opamp_dummy_magic_25_0.VD4.t23 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X549 a_3690_3288.t0 two_stage_opamp_dummy_magic_25_0.V_tot.t0 GNDA.t34 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X550 VOUT+.t122 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VOUT+.t123 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 bgr_11_0.1st_Vout_2.t2 bgr_11_0.V_mir2.t16 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X553 VDDA.t185 bgr_11_0.1st_Vout_1.t25 bgr_11_0.V_TOP.t4 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X554 VDDA.t382 two_stage_opamp_dummy_magic_25_0.Y.t47 VOUT+.t16 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X555 two_stage_opamp_dummy_magic_25_0.V_source.t32 VIN-.t9 two_stage_opamp_dummy_magic_25_0.VD1.t20 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X556 VOUT+.t124 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 VDDA.t360 bgr_11_0.V_mir1.t17 bgr_11_0.1st_Vout_1.t2 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X558 VOUT-.t118 two_stage_opamp_dummy_magic_25_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 GNDA.t128 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t6 VOUT+.t12 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X560 VOUT+.t125 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 two_stage_opamp_dummy_magic_25_0.VD4.t31 two_stage_opamp_dummy_magic_25_0.VD4.t29 two_stage_opamp_dummy_magic_25_0.Y.t23 two_stage_opamp_dummy_magic_25_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X562 VOUT-.t119 two_stage_opamp_dummy_magic_25_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 VOUT-.t120 two_stage_opamp_dummy_magic_25_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 two_stage_opamp_dummy_magic_25_0.VD1.t19 VIN-.t10 two_stage_opamp_dummy_magic_25_0.V_source.t29 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X565 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t4 bgr_11_0.PFET_GATE_10uA.t26 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X566 VOUT-.t121 two_stage_opamp_dummy_magic_25_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 VOUT-.t122 two_stage_opamp_dummy_magic_25_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 bgr_11_0.V_TOP.t40 VDDA.t372 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT-.t123 two_stage_opamp_dummy_magic_25_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 two_stage_opamp_dummy_magic_25_0.VD3.t22 two_stage_opamp_dummy_magic_25_0.Vb3.t26 VDDA.t205 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X571 two_stage_opamp_dummy_magic_25_0.V_source.t5 two_stage_opamp_dummy_magic_25_0.err_amp_out.t4 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X572 VDDA.t280 VDDA.t277 VDDA.t279 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X573 two_stage_opamp_dummy_magic_25_0.VD2.t10 VIN+.t6 two_stage_opamp_dummy_magic_25_0.V_source.t17 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X574 two_stage_opamp_dummy_magic_25_0.V_source.t39 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t27 GNDA.t312 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X575 VOUT+.t18 two_stage_opamp_dummy_magic_25_0.Y.t48 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X576 VDDA.t175 bgr_11_0.PFET_GATE_10uA.t27 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t11 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X577 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t15 VDDA.t274 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X578 VDDA.t401 two_stage_opamp_dummy_magic_25_0.X.t46 VOUT-.t17 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X579 two_stage_opamp_dummy_magic_25_0.X.t1 GNDA.t161 GNDA.t163 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X580 VDDA.t374 bgr_11_0.V_TOP.t41 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t3 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X581 GNDA.t79 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_25_0.V_source.t10 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X582 VDDA.t117 two_stage_opamp_dummy_magic_25_0.Y.t49 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t5 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X583 VOUT+.t126 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 bgr_11_0.V_mir2.t1 bgr_11_0.V_mir2.t0 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X585 VOUT+.t1 a_3830_n584.t0 GNDA.t43 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X586 bgr_11_0.V_TOP.t8 VDDA.t271 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X587 VOUT-.t124 two_stage_opamp_dummy_magic_25_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 VDDA.t270 VDDA.t268 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X589 two_stage_opamp_dummy_magic_25_0.X.t7 two_stage_opamp_dummy_magic_25_0.Vb2.t29 two_stage_opamp_dummy_magic_25_0.VD3.t3 two_stage_opamp_dummy_magic_25_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X590 VOUT-.t125 two_stage_opamp_dummy_magic_25_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 VOUT-.t126 two_stage_opamp_dummy_magic_25_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 a_3810_3288.t1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t11 GNDA.t73 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X594 GNDA.t160 GNDA.t158 two_stage_opamp_dummy_magic_25_0.err_amp_out.t0 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X595 VOUT+.t127 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 a_13960_3288.t0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t0 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X597 VOUT-.t127 two_stage_opamp_dummy_magic_25_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 VOUT+.t128 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 VOUT+.t129 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 VOUT+.t130 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 VOUT-.t128 two_stage_opamp_dummy_magic_25_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 GNDA.t282 VDDA.t422 bgr_11_0.V_TOP.t7 GNDA.t281 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X603 two_stage_opamp_dummy_magic_25_0.Vb2.t7 two_stage_opamp_dummy_magic_25_0.Vb2_2.t3 two_stage_opamp_dummy_magic_25_0.Vb2_2.t5 two_stage_opamp_dummy_magic_25_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X604 two_stage_opamp_dummy_magic_25_0.VD2.t5 two_stage_opamp_dummy_magic_25_0.Vb1.t30 two_stage_opamp_dummy_magic_25_0.Y.t2 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X605 bgr_11_0.PFET_GATE_10uA.t1 bgr_11_0.1st_Vout_2.t26 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X606 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t1 VDDA.t265 VDDA.t267 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X607 VOUT+.t131 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 VOUT+.t132 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 bgr_11_0.cap_res2.t20 bgr_11_0.PFET_GATE_10uA.t9 GNDA.t322 sky130_fd_pr__res_high_po_0p35 l=2.05
X610 VOUT-.t129 two_stage_opamp_dummy_magic_25_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VOUT-.t130 two_stage_opamp_dummy_magic_25_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VOUT-.t131 two_stage_opamp_dummy_magic_25_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 VOUT-.t132 two_stage_opamp_dummy_magic_25_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 VOUT-.t133 two_stage_opamp_dummy_magic_25_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 bgr_11_0.V_p_1.t2 VDDA.t423 GNDA.t280 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X617 bgr_11_0.START_UP.t0 bgr_11_0.V_TOP.t42 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X618 VDDA.t22 two_stage_opamp_dummy_magic_25_0.X.t47 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t6 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X619 VOUT+.t133 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VDDA.t264 VDDA.t262 two_stage_opamp_dummy_magic_25_0.Vb2_2.t9 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X621 GNDA.t145 GNDA.t157 bgr_11_0.Vin-.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X622 VOUT+.t134 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 VOUT-.t15 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t7 GNDA.t289 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X624 VOUT+.t135 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 bgr_11_0.1st_Vout_1.t28 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 GNDA.t145 GNDA.t147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X627 two_stage_opamp_dummy_magic_25_0.VD2.t9 VIN+.t7 two_stage_opamp_dummy_magic_25_0.V_source.t20 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X628 VOUT+.t136 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 bgr_11_0.Vin+.t4 bgr_11_0.V_TOP.t43 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X630 two_stage_opamp_dummy_magic_25_0.VD4.t0 VDDA.t259 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X631 two_stage_opamp_dummy_magic_25_0.V_p_mir.t2 VIN+.t8 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t0 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X632 two_stage_opamp_dummy_magic_25_0.VD2.t8 VIN+.t9 two_stage_opamp_dummy_magic_25_0.V_source.t16 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X633 VOUT+.t137 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 GNDA.t317 two_stage_opamp_dummy_magic_25_0.Y.t50 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t2 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X635 VOUT-.t134 two_stage_opamp_dummy_magic_25_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 VOUT-.t135 two_stage_opamp_dummy_magic_25_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 VOUT-.t136 two_stage_opamp_dummy_magic_25_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VOUT-.t137 two_stage_opamp_dummy_magic_25_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 VOUT+.t138 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 VOUT-.t138 two_stage_opamp_dummy_magic_25_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 bgr_11_0.1st_Vout_2.t1 bgr_11_0.V_mir2.t17 VDDA.t132 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X642 VDDA.t258 VDDA.t255 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X643 VDDA.t254 VDDA.t251 VDDA.t253 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X644 two_stage_opamp_dummy_magic_25_0.Y.t10 two_stage_opamp_dummy_magic_25_0.Vb2.t30 two_stage_opamp_dummy_magic_25_0.VD4.t36 two_stage_opamp_dummy_magic_25_0.VD4.t35 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X645 VDDA.t409 two_stage_opamp_dummy_magic_25_0.Y.t51 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t4 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X646 bgr_11_0.V_TOP.t44 VDDA.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 VOUT+.t139 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 two_stage_opamp_dummy_magic_25_0.Vb3.t4 bgr_11_0.NFET_GATE_10uA.t19 GNDA.t258 GNDA.t257 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X649 VDDA.t395 bgr_11_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t3 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X650 VOUT+.t140 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 VOUT-.t139 two_stage_opamp_dummy_magic_25_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 bgr_11_0.1st_Vout_2.t27 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 GNDA.t145 GNDA.t144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X654 VDDA.t250 VDDA.t248 two_stage_opamp_dummy_magic_25_0.err_amp_out.t2 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X655 VDDA.t61 bgr_11_0.V_TOP.t45 bgr_11_0.Vin-.t1 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X656 VOUT+.t141 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VOUT-.t140 two_stage_opamp_dummy_magic_25_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 VOUT-.t141 two_stage_opamp_dummy_magic_25_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 bgr_11_0.V_mir1.t2 bgr_11_0.V_mir1.t1 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X660 two_stage_opamp_dummy_magic_25_0.VD4.t20 two_stage_opamp_dummy_magic_25_0.Vb3.t27 VDDA.t203 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X661 VOUT+.t142 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 VOUT+.t143 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 VOUT-.t142 two_stage_opamp_dummy_magic_25_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 two_stage_opamp_dummy_magic_25_0.V_source.t35 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t29 GNDA.t298 GNDA.t297 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X666 two_stage_opamp_dummy_magic_25_0.VD2.t4 two_stage_opamp_dummy_magic_25_0.Vb1.t31 two_stage_opamp_dummy_magic_25_0.Y.t1 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X667 VOUT+.t144 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 VOUT-.t143 two_stage_opamp_dummy_magic_25_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 VOUT-.t144 two_stage_opamp_dummy_magic_25_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 VOUT-.t145 two_stage_opamp_dummy_magic_25_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 bgr_11_0.1st_Vout_1.t29 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 a_11420_29718.t0 a_11300_28110.t0 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6
X673 VOUT-.t146 two_stage_opamp_dummy_magic_25_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VOUT+.t145 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 GNDA.t110 two_stage_opamp_dummy_magic_25_0.X.t48 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t3 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X676 VOUT+.t146 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 VDDA.t107 two_stage_opamp_dummy_magic_25_0.X.t49 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t5 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X678 VOUT+.t147 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VOUT-.t147 two_stage_opamp_dummy_magic_25_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 VDDA.t96 two_stage_opamp_dummy_magic_25_0.X.t50 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t4 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X682 VOUT-.t148 two_stage_opamp_dummy_magic_25_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VDDA.t136 bgr_11_0.V_TOP.t46 bgr_11_0.Vin+.t3 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X684 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t0 bgr_11_0.NFET_GATE_10uA.t20 GNDA.t81 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X685 VOUT+.t148 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 VOUT-.t149 two_stage_opamp_dummy_magic_25_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 two_stage_opamp_dummy_magic_25_0.Vb2_2.t2 two_stage_opamp_dummy_magic_25_0.Vb2.t31 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X688 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 GNDA.t328 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_25_0.Vb2.t10 GNDA.t327 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X690 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t13 GNDA.t154 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X691 two_stage_opamp_dummy_magic_25_0.VD2.t7 VIN+.t10 two_stage_opamp_dummy_magic_25_0.V_source.t15 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X692 VDDA.t247 VDDA.t245 bgr_11_0.NFET_GATE_10uA.t4 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X693 VOUT+.t8 two_stage_opamp_dummy_magic_25_0.Y.t52 VDDA.t116 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X694 bgr_11_0.PFET_GATE_10uA.t2 bgr_11_0.1st_Vout_2.t31 VDDA.t140 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X695 two_stage_opamp_dummy_magic_25_0.X.t3 two_stage_opamp_dummy_magic_25_0.VD3.t10 two_stage_opamp_dummy_magic_25_0.VD3.t12 two_stage_opamp_dummy_magic_25_0.VD3.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X696 bgr_11_0.1st_Vout_1.t30 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 VOUT+.t149 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 bgr_11_0.1st_Vout_2.t32 bgr_11_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 GNDA.t85 two_stage_opamp_dummy_magic_25_0.Y.t53 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t1 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X700 bgr_11_0.PFET_GATE_10uA.t6 VDDA.t424 GNDA.t275 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X701 two_stage_opamp_dummy_magic_25_0.VD3.t5 two_stage_opamp_dummy_magic_25_0.Vb2.t32 two_stage_opamp_dummy_magic_25_0.X.t6 two_stage_opamp_dummy_magic_25_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X702 GNDA.t315 a_5820_28304.t1 GNDA.t46 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X703 VDDA.t114 GNDA.t151 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X704 VDDA.t379 two_stage_opamp_dummy_magic_25_0.Y.t54 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t3 GNDA.t316 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X705 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 bgr_11_0.Vin+.t2 bgr_11_0.V_TOP.t47 VDDA.t138 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X707 two_stage_opamp_dummy_magic_25_0.VD4.t24 two_stage_opamp_dummy_magic_25_0.Vb3.t28 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X708 GNDA.t63 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t8 VOUT-.t3 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X709 GNDA.t150 GNDA.t148 bgr_11_0.NFET_GATE_10uA.t2 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X710 VOUT+.t150 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 VOUT-.t150 two_stage_opamp_dummy_magic_25_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 VOUT+.t151 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 bgr_11_0.V_p_1.t0 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t0 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X714 two_stage_opamp_dummy_magic_25_0.V_err_p.t0 two_stage_opamp_dummy_magic_25_0.V_err_gate.t9 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X715 bgr_11_0.1st_Vout_2.t0 bgr_11_0.V_mir2.t18 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X716 two_stage_opamp_dummy_magic_25_0.Vb2_2.t1 two_stage_opamp_dummy_magic_25_0.Vb2.t3 two_stage_opamp_dummy_magic_25_0.Vb2.t4 two_stage_opamp_dummy_magic_25_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X717 bgr_11_0.V_TOP.t5 bgr_11_0.1st_Vout_1.t32 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X718 VOUT-.t151 two_stage_opamp_dummy_magic_25_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 VOUT+.t152 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT-.t152 two_stage_opamp_dummy_magic_25_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VOUT-.t153 two_stage_opamp_dummy_magic_25_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 VOUT+.t153 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 two_stage_opamp_dummy_magic_25_0.Vb3.t2 GNDA.t141 GNDA.t143 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X724 two_stage_opamp_dummy_magic_25_0.VD2.t20 two_stage_opamp_dummy_magic_25_0.Vb1.t32 two_stage_opamp_dummy_magic_25_0.Y.t0 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X725 bgr_11_0.1st_Vout_1.t1 bgr_11_0.V_mir1.t18 VDDA.t362 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X726 VOUT+.t154 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 VOUT+.t155 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 GNDA.t250 bgr_11_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_25_0.Vb3.t3 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X729 VOUT-.t11 two_stage_opamp_dummy_magic_25_0.X.t51 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X730 VOUT+.t156 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VOUT-.t9 a_13940_n584.t0 GNDA.t102 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X732 GNDA.t265 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t9 VOUT-.t13 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X733 GNDA.t107 two_stage_opamp_dummy_magic_25_0.X.t52 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t2 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X734 VOUT-.t154 two_stage_opamp_dummy_magic_25_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 bgr_11_0.V_TOP.t48 VDDA.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 GNDA.t106 two_stage_opamp_dummy_magic_25_0.X.t53 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t1 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X737 GNDA.t38 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_25_0.V_source.t3 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X738 VDDA.t197 two_stage_opamp_dummy_magic_25_0.X.t54 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t3 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X739 VOUT-.t155 two_stage_opamp_dummy_magic_25_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 VDDA.t244 VDDA.t242 bgr_11_0.PFET_GATE_10uA.t7 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X741 bgr_11_0.V_TOP.t49 VDDA.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 VOUT-.t156 two_stage_opamp_dummy_magic_25_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 two_stage_opamp_dummy_magic_25_0.V_source.t37 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t31 GNDA.t305 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
R0 VOUT-.n178 VOUT-.t9 110.191
R1 VOUT-.n39 VOUT-.n38 34.9935
R2 VOUT-.n28 VOUT-.n27 34.9935
R3 VOUT-.n30 VOUT-.n29 34.9935
R4 VOUT-.n33 VOUT-.n32 34.9935
R5 VOUT-.n36 VOUT-.n35 34.9935
R6 VOUT-.n42 VOUT-.n41 34.9935
R7 VOUT-.n185 VOUT-.n184 9.73997
R8 VOUT-.n181 VOUT-.n180 9.73997
R9 VOUT-.n188 VOUT-.n187 9.73997
R10 VOUT-.n186 VOUT-.n181 6.64633
R11 VOUT-.n186 VOUT-.n185 6.64633
R12 VOUT-.n38 VOUT-.t17 6.56717
R13 VOUT-.n38 VOUT-.t12 6.56717
R14 VOUT-.n27 VOUT-.t0 6.56717
R15 VOUT-.n27 VOUT-.t11 6.56717
R16 VOUT-.n29 VOUT-.t10 6.56717
R17 VOUT-.n29 VOUT-.t2 6.56717
R18 VOUT-.n32 VOUT-.t6 6.56717
R19 VOUT-.n32 VOUT-.t1 6.56717
R20 VOUT-.n35 VOUT-.t4 6.56717
R21 VOUT-.n35 VOUT-.t7 6.56717
R22 VOUT-.n41 VOUT-.t16 6.56717
R23 VOUT-.n41 VOUT-.t5 6.56717
R24 VOUT-.n31 VOUT-.n28 6.3755
R25 VOUT-.n40 VOUT-.n39 6.3755
R26 VOUT-.n188 VOUT-.n186 6.02133
R27 VOUT-.n31 VOUT-.n30 5.813
R28 VOUT-.n34 VOUT-.n33 5.813
R29 VOUT-.n37 VOUT-.n36 5.813
R30 VOUT-.n42 VOUT-.n40 5.813
R31 VOUT-.n46 VOUT-.n26 5.063
R32 VOUT-.n43 VOUT-.n19 5.063
R33 VOUT-.n109 VOUT-.t35 4.8295
R34 VOUT-.n108 VOUT-.t71 4.8295
R35 VOUT-.n107 VOUT-.t106 4.8295
R36 VOUT-.n106 VOUT-.t141 4.8295
R37 VOUT-.n105 VOUT-.t54 4.8295
R38 VOUT-.n104 VOUT-.t100 4.8295
R39 VOUT-.n110 VOUT-.t147 4.8295
R40 VOUT-.n121 VOUT-.t132 4.8295
R41 VOUT-.n122 VOUT-.t42 4.8295
R42 VOUT-.n124 VOUT-.t103 4.8295
R43 VOUT-.n125 VOUT-.t86 4.8295
R44 VOUT-.n127 VOUT-.t67 4.8295
R45 VOUT-.n128 VOUT-.t48 4.8295
R46 VOUT-.n130 VOUT-.t98 4.8295
R47 VOUT-.n131 VOUT-.t80 4.8295
R48 VOUT-.n133 VOUT-.t61 4.8295
R49 VOUT-.n134 VOUT-.t43 4.8295
R50 VOUT-.n136 VOUT-.t19 4.8295
R51 VOUT-.n137 VOUT-.t142 4.8295
R52 VOUT-.n139 VOUT-.t55 4.8295
R53 VOUT-.n140 VOUT-.t36 4.8295
R54 VOUT-.n142 VOUT-.t151 4.8295
R55 VOUT-.n143 VOUT-.t134 4.8295
R56 VOUT-.n145 VOUT-.t111 4.8295
R57 VOUT-.n146 VOUT-.t97 4.8295
R58 VOUT-.n148 VOUT-.t74 4.8295
R59 VOUT-.n149 VOUT-.t59 4.8295
R60 VOUT-.n71 VOUT-.t96 4.8295
R61 VOUT-.n73 VOUT-.t58 4.8295
R62 VOUT-.n86 VOUT-.t117 4.8295
R63 VOUT-.n87 VOUT-.t102 4.8295
R64 VOUT-.n89 VOUT-.t153 4.8295
R65 VOUT-.n90 VOUT-.t136 4.8295
R66 VOUT-.n92 VOUT-.t62 4.8295
R67 VOUT-.n93 VOUT-.t30 4.8295
R68 VOUT-.n95 VOUT-.t66 4.8295
R69 VOUT-.n96 VOUT-.t47 4.8295
R70 VOUT-.n98 VOUT-.t29 4.8295
R71 VOUT-.n99 VOUT-.t150 4.8295
R72 VOUT-.n101 VOUT-.t70 4.8295
R73 VOUT-.n102 VOUT-.t53 4.8295
R74 VOUT-.n151 VOUT-.t108 4.8295
R75 VOUT-.n112 VOUT-.t75 4.8154
R76 VOUT-.n74 VOUT-.t146 4.806
R77 VOUT-.n75 VOUT-.t119 4.806
R78 VOUT-.n76 VOUT-.t139 4.806
R79 VOUT-.n77 VOUT-.t38 4.806
R80 VOUT-.n78 VOUT-.t154 4.806
R81 VOUT-.n79 VOUT-.t56 4.806
R82 VOUT-.n80 VOUT-.t91 4.806
R83 VOUT-.n81 VOUT-.t127 4.806
R84 VOUT-.n82 VOUT-.t107 4.806
R85 VOUT-.n83 VOUT-.t148 4.806
R86 VOUT-.n84 VOUT-.t45 4.806
R87 VOUT-.n109 VOUT-.t52 4.5005
R88 VOUT-.n108 VOUT-.t90 4.5005
R89 VOUT-.n107 VOUT-.t125 4.5005
R90 VOUT-.n106 VOUT-.t25 4.5005
R91 VOUT-.n105 VOUT-.t145 4.5005
R92 VOUT-.n104 VOUT-.t64 4.5005
R93 VOUT-.n120 VOUT-.t23 4.5005
R94 VOUT-.n119 VOUT-.t46 4.5005
R95 VOUT-.n118 VOUT-.t149 4.5005
R96 VOUT-.n117 VOUT-.t109 4.5005
R97 VOUT-.n116 VOUT-.t128 4.5005
R98 VOUT-.n115 VOUT-.t94 4.5005
R99 VOUT-.n114 VOUT-.t57 4.5005
R100 VOUT-.n113 VOUT-.t155 4.5005
R101 VOUT-.n112 VOUT-.t41 4.5005
R102 VOUT-.n111 VOUT-.t140 4.5005
R103 VOUT-.n110 VOUT-.t122 4.5005
R104 VOUT-.n121 VOUT-.t95 4.5005
R105 VOUT-.n123 VOUT-.t60 4.5005
R106 VOUT-.n122 VOUT-.t78 4.5005
R107 VOUT-.n124 VOUT-.t69 4.5005
R108 VOUT-.n126 VOUT-.t32 4.5005
R109 VOUT-.n125 VOUT-.t120 4.5005
R110 VOUT-.n127 VOUT-.t27 4.5005
R111 VOUT-.n129 VOUT-.t131 4.5005
R112 VOUT-.n128 VOUT-.t82 4.5005
R113 VOUT-.n130 VOUT-.t65 4.5005
R114 VOUT-.n132 VOUT-.t26 4.5005
R115 VOUT-.n131 VOUT-.t113 4.5005
R116 VOUT-.n133 VOUT-.t24 4.5005
R117 VOUT-.n135 VOUT-.t126 4.5005
R118 VOUT-.n134 VOUT-.t76 4.5005
R119 VOUT-.n136 VOUT-.t123 4.5005
R120 VOUT-.n138 VOUT-.t88 4.5005
R121 VOUT-.n137 VOUT-.t37 4.5005
R122 VOUT-.n139 VOUT-.t156 4.5005
R123 VOUT-.n141 VOUT-.t121 4.5005
R124 VOUT-.n140 VOUT-.t72 4.5005
R125 VOUT-.n142 VOUT-.t115 4.5005
R126 VOUT-.n144 VOUT-.t83 4.5005
R127 VOUT-.n143 VOUT-.t31 4.5005
R128 VOUT-.n145 VOUT-.t77 4.5005
R129 VOUT-.n147 VOUT-.t44 4.5005
R130 VOUT-.n146 VOUT-.t129 4.5005
R131 VOUT-.n148 VOUT-.t40 4.5005
R132 VOUT-.n150 VOUT-.t143 4.5005
R133 VOUT-.n149 VOUT-.t93 4.5005
R134 VOUT-.n71 VOUT-.t63 4.5005
R135 VOUT-.n72 VOUT-.t22 4.5005
R136 VOUT-.n73 VOUT-.t20 4.5005
R137 VOUT-.n85 VOUT-.t118 4.5005
R138 VOUT-.n84 VOUT-.t144 4.5005
R139 VOUT-.n83 VOUT-.t105 4.5005
R140 VOUT-.n82 VOUT-.t68 4.5005
R141 VOUT-.n81 VOUT-.t89 4.5005
R142 VOUT-.n80 VOUT-.t51 4.5005
R143 VOUT-.n79 VOUT-.t152 4.5005
R144 VOUT-.n78 VOUT-.t112 4.5005
R145 VOUT-.n77 VOUT-.t135 4.5005
R146 VOUT-.n76 VOUT-.t101 4.5005
R147 VOUT-.n75 VOUT-.t79 4.5005
R148 VOUT-.n74 VOUT-.t104 4.5005
R149 VOUT-.n86 VOUT-.t85 4.5005
R150 VOUT-.n88 VOUT-.t50 4.5005
R151 VOUT-.n87 VOUT-.t137 4.5005
R152 VOUT-.n89 VOUT-.t116 4.5005
R153 VOUT-.n91 VOUT-.t84 4.5005
R154 VOUT-.n90 VOUT-.t33 4.5005
R155 VOUT-.n92 VOUT-.t110 4.5005
R156 VOUT-.n94 VOUT-.t21 4.5005
R157 VOUT-.n93 VOUT-.t114 4.5005
R158 VOUT-.n95 VOUT-.t28 4.5005
R159 VOUT-.n97 VOUT-.t130 4.5005
R160 VOUT-.n96 VOUT-.t81 4.5005
R161 VOUT-.n98 VOUT-.t133 4.5005
R162 VOUT-.n100 VOUT-.t99 4.5005
R163 VOUT-.n99 VOUT-.t49 4.5005
R164 VOUT-.n101 VOUT-.t34 4.5005
R165 VOUT-.n103 VOUT-.t138 4.5005
R166 VOUT-.n102 VOUT-.t87 4.5005
R167 VOUT-.n151 VOUT-.t73 4.5005
R168 VOUT-.n152 VOUT-.t39 4.5005
R169 VOUT-.n153 VOUT-.t124 4.5005
R170 VOUT-.n154 VOUT-.t92 4.5005
R171 VOUT-.n47 VOUT-.n46 4.5005
R172 VOUT-.n45 VOUT-.n24 4.5005
R173 VOUT-.n44 VOUT-.n23 4.5005
R174 VOUT-.n43 VOUT-.n20 4.5005
R175 VOUT-.n65 VOUT-.n64 4.5005
R176 VOUT-.n16 VOUT-.n13 4.5005
R177 VOUT-.n65 VOUT-.n13 4.5005
R178 VOUT-.n66 VOUT-.n9 4.5005
R179 VOUT-.n66 VOUT-.n11 4.5005
R180 VOUT-.n66 VOUT-.n65 4.5005
R181 VOUT-.n163 VOUT-.n69 4.5005
R182 VOUT-.n164 VOUT-.n163 4.5005
R183 VOUT-.n164 VOUT-.n5 4.5005
R184 VOUT-.n165 VOUT-.n4 4.5005
R185 VOUT-.n165 VOUT-.n164 4.5005
R186 VOUT-.n177 VOUT-.n176 4.5005
R187 VOUT-.n177 VOUT-.n1 4.5005
R188 VOUT-.n173 VOUT-.n1 4.5005
R189 VOUT-.n170 VOUT-.n1 4.5005
R190 VOUT-.n171 VOUT-.n1 4.5005
R191 VOUT-.n173 VOUT-.n172 4.5005
R192 VOUT-.n172 VOUT-.n170 4.5005
R193 VOUT-.n172 VOUT-.n171 4.5005
R194 VOUT-.n184 VOUT-.t3 3.42907
R195 VOUT-.n184 VOUT-.t18 3.42907
R196 VOUT-.n180 VOUT-.t8 3.42907
R197 VOUT-.n180 VOUT-.t15 3.42907
R198 VOUT-.n187 VOUT-.t13 3.42907
R199 VOUT-.n187 VOUT-.t14 3.42907
R200 VOUT-.n63 VOUT-.n62 2.24601
R201 VOUT-.n14 VOUT-.n8 2.24601
R202 VOUT-.n175 VOUT-.n174 2.24601
R203 VOUT-.n169 VOUT-.n168 2.24601
R204 VOUT-.n162 VOUT-.n161 2.24477
R205 VOUT-.n7 VOUT-.n2 2.24477
R206 VOUT-.n66 VOUT-.n10 2.24063
R207 VOUT-.n165 VOUT-.n3 2.24063
R208 VOUT-.n172 VOUT-.n0 2.24063
R209 VOUT-.n13 VOUT-.n12 2.24063
R210 VOUT-.n163 VOUT-.n67 2.24063
R211 VOUT-.n68 VOUT-.n5 2.24063
R212 VOUT-.n176 VOUT-.n167 2.24063
R213 VOUT-.n176 VOUT-.n166 2.24063
R214 VOUT-.n64 VOUT-.n17 2.23934
R215 VOUT-.n64 VOUT-.n15 2.23934
R216 VOUT-.n185 VOUT-.n183 1.62886
R217 VOUT-.n196 VOUT-.n181 1.52133
R218 VOUT-.n189 VOUT-.n188 1.52133
R219 VOUT-.n50 VOUT-.n25 1.5005
R220 VOUT-.n52 VOUT-.n51 1.5005
R221 VOUT-.n53 VOUT-.n22 1.5005
R222 VOUT-.n55 VOUT-.n54 1.5005
R223 VOUT-.n56 VOUT-.n21 1.5005
R224 VOUT-.n58 VOUT-.n57 1.5005
R225 VOUT-.n59 VOUT-.n18 1.5005
R226 VOUT-.n61 VOUT-.n60 1.5005
R227 VOUT-.n191 VOUT-.n190 1.5005
R228 VOUT-.n192 VOUT-.n182 1.5005
R229 VOUT-.n194 VOUT-.n193 1.5005
R230 VOUT-.n195 VOUT-.n179 1.5005
R231 VOUT-.n197 VOUT-.n196 1.5005
R232 VOUT-.n30 VOUT-.n20 1.313
R233 VOUT-.n33 VOUT-.n23 1.313
R234 VOUT-.n36 VOUT-.n24 1.313
R235 VOUT-.n47 VOUT-.n42 1.313
R236 VOUT-.n28 VOUT-.n19 1.313
R237 VOUT-.n39 VOUT-.n26 1.313
R238 VOUT-.n161 VOUT-.n160 1.1455
R239 VOUT-.n155 VOUT-.n6 1.13717
R240 VOUT-.n157 VOUT-.n156 1.13717
R241 VOUT-.n159 VOUT-.n158 1.13717
R242 VOUT-.n164 VOUT-.n6 1.13717
R243 VOUT-.n157 VOUT-.n7 1.13717
R244 VOUT-.n158 VOUT-.n4 1.13717
R245 VOUT-.n70 VOUT-.n69 1.13717
R246 VOUT-.n49 VOUT-.n26 0.715216
R247 VOUT-.n58 VOUT-.n20 0.65675
R248 VOUT-.n54 VOUT-.n23 0.65675
R249 VOUT-.n52 VOUT-.n24 0.65675
R250 VOUT-.n48 VOUT-.n47 0.65675
R251 VOUT-.n60 VOUT-.n19 0.65675
R252 VOUT-.n160 VOUT-.n159 0.585
R253 VOUT-.n176 VOUT-.n165 0.5705
R254 VOUT-.n50 VOUT-.n49 0.564601
R255 VOUT-.n46 VOUT-.n45 0.563
R256 VOUT-.n45 VOUT-.n44 0.563
R257 VOUT-.n44 VOUT-.n43 0.563
R258 VOUT-.n34 VOUT-.n31 0.563
R259 VOUT-.n37 VOUT-.n34 0.563
R260 VOUT-.n40 VOUT-.n37 0.563
R261 VOUT-.n62 VOUT-.n61 0.495292
R262 VOUT-.n120 VOUT-.n104 0.3295
R263 VOUT-.n120 VOUT-.n119 0.3295
R264 VOUT-.n119 VOUT-.n118 0.3295
R265 VOUT-.n118 VOUT-.n117 0.3295
R266 VOUT-.n117 VOUT-.n116 0.3295
R267 VOUT-.n116 VOUT-.n115 0.3295
R268 VOUT-.n115 VOUT-.n114 0.3295
R269 VOUT-.n114 VOUT-.n113 0.3295
R270 VOUT-.n113 VOUT-.n112 0.3295
R271 VOUT-.n112 VOUT-.n111 0.3295
R272 VOUT-.n111 VOUT-.n110 0.3295
R273 VOUT-.n123 VOUT-.n121 0.3295
R274 VOUT-.n123 VOUT-.n122 0.3295
R275 VOUT-.n126 VOUT-.n124 0.3295
R276 VOUT-.n126 VOUT-.n125 0.3295
R277 VOUT-.n129 VOUT-.n127 0.3295
R278 VOUT-.n129 VOUT-.n128 0.3295
R279 VOUT-.n132 VOUT-.n130 0.3295
R280 VOUT-.n132 VOUT-.n131 0.3295
R281 VOUT-.n135 VOUT-.n133 0.3295
R282 VOUT-.n135 VOUT-.n134 0.3295
R283 VOUT-.n138 VOUT-.n136 0.3295
R284 VOUT-.n138 VOUT-.n137 0.3295
R285 VOUT-.n141 VOUT-.n139 0.3295
R286 VOUT-.n141 VOUT-.n140 0.3295
R287 VOUT-.n144 VOUT-.n142 0.3295
R288 VOUT-.n144 VOUT-.n143 0.3295
R289 VOUT-.n147 VOUT-.n145 0.3295
R290 VOUT-.n147 VOUT-.n146 0.3295
R291 VOUT-.n150 VOUT-.n148 0.3295
R292 VOUT-.n150 VOUT-.n149 0.3295
R293 VOUT-.n72 VOUT-.n71 0.3295
R294 VOUT-.n85 VOUT-.n73 0.3295
R295 VOUT-.n85 VOUT-.n84 0.3295
R296 VOUT-.n84 VOUT-.n83 0.3295
R297 VOUT-.n83 VOUT-.n82 0.3295
R298 VOUT-.n82 VOUT-.n81 0.3295
R299 VOUT-.n81 VOUT-.n80 0.3295
R300 VOUT-.n80 VOUT-.n79 0.3295
R301 VOUT-.n79 VOUT-.n78 0.3295
R302 VOUT-.n78 VOUT-.n77 0.3295
R303 VOUT-.n77 VOUT-.n76 0.3295
R304 VOUT-.n76 VOUT-.n75 0.3295
R305 VOUT-.n75 VOUT-.n74 0.3295
R306 VOUT-.n88 VOUT-.n86 0.3295
R307 VOUT-.n88 VOUT-.n87 0.3295
R308 VOUT-.n91 VOUT-.n89 0.3295
R309 VOUT-.n91 VOUT-.n90 0.3295
R310 VOUT-.n94 VOUT-.n92 0.3295
R311 VOUT-.n94 VOUT-.n93 0.3295
R312 VOUT-.n97 VOUT-.n95 0.3295
R313 VOUT-.n97 VOUT-.n96 0.3295
R314 VOUT-.n100 VOUT-.n98 0.3295
R315 VOUT-.n100 VOUT-.n99 0.3295
R316 VOUT-.n103 VOUT-.n101 0.3295
R317 VOUT-.n103 VOUT-.n102 0.3295
R318 VOUT-.n152 VOUT-.n151 0.3295
R319 VOUT-.n153 VOUT-.n152 0.3295
R320 VOUT-.n113 VOUT-.n109 0.3154
R321 VOUT-.n191 VOUT-.n183 0.314966
R322 VOUT-.n154 VOUT-.n153 0.3107
R323 VOUT-.n114 VOUT-.n108 0.306
R324 VOUT-.n115 VOUT-.n107 0.306
R325 VOUT-.n116 VOUT-.n106 0.306
R326 VOUT-.n117 VOUT-.n105 0.306
R327 VOUT-.n123 VOUT-.n120 0.2825
R328 VOUT-.n126 VOUT-.n123 0.2825
R329 VOUT-.n129 VOUT-.n126 0.2825
R330 VOUT-.n132 VOUT-.n129 0.2825
R331 VOUT-.n135 VOUT-.n132 0.2825
R332 VOUT-.n138 VOUT-.n135 0.2825
R333 VOUT-.n141 VOUT-.n138 0.2825
R334 VOUT-.n144 VOUT-.n141 0.2825
R335 VOUT-.n147 VOUT-.n144 0.2825
R336 VOUT-.n150 VOUT-.n147 0.2825
R337 VOUT-.n85 VOUT-.n72 0.2825
R338 VOUT-.n88 VOUT-.n85 0.2825
R339 VOUT-.n91 VOUT-.n88 0.2825
R340 VOUT-.n94 VOUT-.n91 0.2825
R341 VOUT-.n97 VOUT-.n94 0.2825
R342 VOUT-.n100 VOUT-.n97 0.2825
R343 VOUT-.n103 VOUT-.n100 0.2825
R344 VOUT-.n152 VOUT-.n103 0.2825
R345 VOUT-.n152 VOUT-.n150 0.2825
R346 VOUT-.n163 VOUT-.n66 0.2655
R347 VOUT- VOUT-.n178 0.198417
R348 VOUT-.n178 VOUT-.n177 0.193208
R349 VOUT- VOUT-.n197 0.182792
R350 VOUT-.n155 VOUT-.n154 0.138367
R351 VOUT-.n189 VOUT-.n183 0.0891864
R352 VOUT-.n60 VOUT-.n59 0.0577917
R353 VOUT-.n59 VOUT-.n58 0.0577917
R354 VOUT-.n58 VOUT-.n21 0.0577917
R355 VOUT-.n54 VOUT-.n21 0.0577917
R356 VOUT-.n54 VOUT-.n53 0.0577917
R357 VOUT-.n53 VOUT-.n52 0.0577917
R358 VOUT-.n52 VOUT-.n25 0.0577917
R359 VOUT-.n48 VOUT-.n25 0.0577917
R360 VOUT-.n61 VOUT-.n18 0.0577917
R361 VOUT-.n57 VOUT-.n18 0.0577917
R362 VOUT-.n57 VOUT-.n56 0.0577917
R363 VOUT-.n56 VOUT-.n55 0.0577917
R364 VOUT-.n55 VOUT-.n22 0.0577917
R365 VOUT-.n51 VOUT-.n22 0.0577917
R366 VOUT-.n51 VOUT-.n50 0.0577917
R367 VOUT-.n49 VOUT-.n48 0.054517
R368 VOUT-.n170 VOUT-.n169 0.047375
R369 VOUT-.n174 VOUT-.n173 0.047375
R370 VOUT-.n164 VOUT-.n7 0.0421667
R371 VOUT-.n65 VOUT-.n14 0.0421667
R372 VOUT-.n196 VOUT-.n195 0.0421667
R373 VOUT-.n195 VOUT-.n194 0.0421667
R374 VOUT-.n194 VOUT-.n182 0.0421667
R375 VOUT-.n190 VOUT-.n182 0.0421667
R376 VOUT-.n190 VOUT-.n189 0.0421667
R377 VOUT-.n197 VOUT-.n179 0.0421667
R378 VOUT-.n193 VOUT-.n179 0.0421667
R379 VOUT-.n193 VOUT-.n192 0.0421667
R380 VOUT-.n192 VOUT-.n191 0.0421667
R381 VOUT-.n15 VOUT-.n14 0.0243161
R382 VOUT-.n17 VOUT-.n9 0.0243161
R383 VOUT-.n17 VOUT-.n16 0.0243161
R384 VOUT-.n15 VOUT-.n11 0.0243161
R385 VOUT-.n161 VOUT-.n3 0.0217373
R386 VOUT-.n62 VOUT-.n10 0.0217373
R387 VOUT-.n16 VOUT-.n10 0.0217373
R388 VOUT-.n69 VOUT-.n3 0.0217373
R389 VOUT-.n177 VOUT-.n0 0.0217373
R390 VOUT-.n174 VOUT-.n0 0.0217373
R391 VOUT-.n67 VOUT-.n7 0.0217373
R392 VOUT-.n69 VOUT-.n68 0.0217373
R393 VOUT-.n12 VOUT-.n9 0.0217373
R394 VOUT-.n12 VOUT-.n11 0.0217373
R395 VOUT-.n67 VOUT-.n4 0.0217373
R396 VOUT-.n68 VOUT-.n4 0.0217373
R397 VOUT-.n171 VOUT-.n166 0.0217373
R398 VOUT-.n170 VOUT-.n167 0.0217373
R399 VOUT-.n173 VOUT-.n167 0.0217373
R400 VOUT-.n169 VOUT-.n166 0.0217373
R401 VOUT-.n156 VOUT-.n155 0.0161667
R402 VOUT-.n159 VOUT-.n156 0.0161667
R403 VOUT-.n157 VOUT-.n6 0.0161667
R404 VOUT-.n158 VOUT-.n157 0.0161667
R405 VOUT-.n158 VOUT-.n70 0.0161667
R406 VOUT-.n162 VOUT-.n5 0.0134654
R407 VOUT-.n165 VOUT-.n2 0.0134654
R408 VOUT-.n163 VOUT-.n162 0.0134654
R409 VOUT-.n5 VOUT-.n2 0.0134654
R410 VOUT-.n63 VOUT-.n13 0.0109778
R411 VOUT-.n66 VOUT-.n8 0.0109778
R412 VOUT-.n175 VOUT-.n1 0.0109778
R413 VOUT-.n172 VOUT-.n168 0.0109778
R414 VOUT-.n64 VOUT-.n63 0.0109778
R415 VOUT-.n13 VOUT-.n8 0.0109778
R416 VOUT-.n176 VOUT-.n175 0.0109778
R417 VOUT-.n168 VOUT-.n1 0.0109778
R418 VOUT-.n160 VOUT-.n70 0.00872683
R419 two_stage_opamp_dummy_magic_25_0.cap_res_X two_stage_opamp_dummy_magic_25_0.cap_res_X.t138 49.4254
R420 two_stage_opamp_dummy_magic_25_0.cap_res_X two_stage_opamp_dummy_magic_25_0.cap_res_X.t15 1.481
R421 two_stage_opamp_dummy_magic_25_0.cap_res_X.t34 two_stage_opamp_dummy_magic_25_0.cap_res_X.t9 0.1603
R422 two_stage_opamp_dummy_magic_25_0.cap_res_X.t16 two_stage_opamp_dummy_magic_25_0.cap_res_X.t34 0.1603
R423 two_stage_opamp_dummy_magic_25_0.cap_res_X.t115 two_stage_opamp_dummy_magic_25_0.cap_res_X.t81 0.1603
R424 two_stage_opamp_dummy_magic_25_0.cap_res_X.t104 two_stage_opamp_dummy_magic_25_0.cap_res_X.t121 0.1603
R425 two_stage_opamp_dummy_magic_25_0.cap_res_X.t1 two_stage_opamp_dummy_magic_25_0.cap_res_X.t104 0.1603
R426 two_stage_opamp_dummy_magic_25_0.cap_res_X.t66 two_stage_opamp_dummy_magic_25_0.cap_res_X.t85 0.1603
R427 two_stage_opamp_dummy_magic_25_0.cap_res_X.t99 two_stage_opamp_dummy_magic_25_0.cap_res_X.t66 0.1603
R428 two_stage_opamp_dummy_magic_25_0.cap_res_X.t31 two_stage_opamp_dummy_magic_25_0.cap_res_X.t50 0.1603
R429 two_stage_opamp_dummy_magic_25_0.cap_res_X.t62 two_stage_opamp_dummy_magic_25_0.cap_res_X.t31 0.1603
R430 two_stage_opamp_dummy_magic_25_0.cap_res_X.t92 two_stage_opamp_dummy_magic_25_0.cap_res_X.t56 0.1603
R431 two_stage_opamp_dummy_magic_25_0.cap_res_X.t78 two_stage_opamp_dummy_magic_25_0.cap_res_X.t114 0.1603
R432 two_stage_opamp_dummy_magic_25_0.cap_res_X.t61 two_stage_opamp_dummy_magic_25_0.cap_res_X.t24 0.1603
R433 two_stage_opamp_dummy_magic_25_0.cap_res_X.t36 two_stage_opamp_dummy_magic_25_0.cap_res_X.t70 0.1603
R434 two_stage_opamp_dummy_magic_25_0.cap_res_X.t87 two_stage_opamp_dummy_magic_25_0.cap_res_X.t53 0.1603
R435 two_stage_opamp_dummy_magic_25_0.cap_res_X.t74 two_stage_opamp_dummy_magic_25_0.cap_res_X.t108 0.1603
R436 two_stage_opamp_dummy_magic_25_0.cap_res_X.t129 two_stage_opamp_dummy_magic_25_0.cap_res_X.t89 0.1603
R437 two_stage_opamp_dummy_magic_25_0.cap_res_X.t43 two_stage_opamp_dummy_magic_25_0.cap_res_X.t76 0.1603
R438 two_stage_opamp_dummy_magic_25_0.cap_res_X.t91 two_stage_opamp_dummy_magic_25_0.cap_res_X.t58 0.1603
R439 two_stage_opamp_dummy_magic_25_0.cap_res_X.t80 two_stage_opamp_dummy_magic_25_0.cap_res_X.t113 0.1603
R440 two_stage_opamp_dummy_magic_25_0.cap_res_X.t132 two_stage_opamp_dummy_magic_25_0.cap_res_X.t95 0.1603
R441 two_stage_opamp_dummy_magic_25_0.cap_res_X.t119 two_stage_opamp_dummy_magic_25_0.cap_res_X.t14 0.1603
R442 two_stage_opamp_dummy_magic_25_0.cap_res_X.t33 two_stage_opamp_dummy_magic_25_0.cap_res_X.t137 0.1603
R443 two_stage_opamp_dummy_magic_25_0.cap_res_X.t84 two_stage_opamp_dummy_magic_25_0.cap_res_X.t120 0.1603
R444 two_stage_opamp_dummy_magic_25_0.cap_res_X.t0 two_stage_opamp_dummy_magic_25_0.cap_res_X.t101 0.1603
R445 two_stage_opamp_dummy_magic_25_0.cap_res_X.t125 two_stage_opamp_dummy_magic_25_0.cap_res_X.t22 0.1603
R446 two_stage_opamp_dummy_magic_25_0.cap_res_X.t41 two_stage_opamp_dummy_magic_25_0.cap_res_X.t5 0.1603
R447 two_stage_opamp_dummy_magic_25_0.cap_res_X.t27 two_stage_opamp_dummy_magic_25_0.cap_res_X.t59 0.1603
R448 two_stage_opamp_dummy_magic_25_0.cap_res_X.t79 two_stage_opamp_dummy_magic_25_0.cap_res_X.t45 0.1603
R449 two_stage_opamp_dummy_magic_25_0.cap_res_X.t63 two_stage_opamp_dummy_magic_25_0.cap_res_X.t97 0.1603
R450 two_stage_opamp_dummy_magic_25_0.cap_res_X.t116 two_stage_opamp_dummy_magic_25_0.cap_res_X.t82 0.1603
R451 two_stage_opamp_dummy_magic_25_0.cap_res_X.t32 two_stage_opamp_dummy_magic_25_0.cap_res_X.t64 0.1603
R452 two_stage_opamp_dummy_magic_25_0.cap_res_X.t83 two_stage_opamp_dummy_magic_25_0.cap_res_X.t48 0.1603
R453 two_stage_opamp_dummy_magic_25_0.cap_res_X.t69 two_stage_opamp_dummy_magic_25_0.cap_res_X.t103 0.1603
R454 two_stage_opamp_dummy_magic_25_0.cap_res_X.t122 two_stage_opamp_dummy_magic_25_0.cap_res_X.t86 0.1603
R455 two_stage_opamp_dummy_magic_25_0.cap_res_X.t107 two_stage_opamp_dummy_magic_25_0.cap_res_X.t6 0.1603
R456 two_stage_opamp_dummy_magic_25_0.cap_res_X.t23 two_stage_opamp_dummy_magic_25_0.cap_res_X.t127 0.1603
R457 two_stage_opamp_dummy_magic_25_0.cap_res_X.t75 two_stage_opamp_dummy_magic_25_0.cap_res_X.t109 0.1603
R458 two_stage_opamp_dummy_magic_25_0.cap_res_X.t128 two_stage_opamp_dummy_magic_25_0.cap_res_X.t90 0.1603
R459 two_stage_opamp_dummy_magic_25_0.cap_res_X.t42 two_stage_opamp_dummy_magic_25_0.cap_res_X.t126 0.1603
R460 two_stage_opamp_dummy_magic_25_0.cap_res_X.t46 two_stage_opamp_dummy_magic_25_0.cap_res_X.t94 0.1603
R461 two_stage_opamp_dummy_magic_25_0.cap_res_X.t123 two_stage_opamp_dummy_magic_25_0.cap_res_X.t20 0.1603
R462 two_stage_opamp_dummy_magic_25_0.cap_res_X.t40 two_stage_opamp_dummy_magic_25_0.cap_res_X.t3 0.1603
R463 two_stage_opamp_dummy_magic_25_0.cap_res_X.t19 two_stage_opamp_dummy_magic_25_0.cap_res_X.t54 0.1603
R464 two_stage_opamp_dummy_magic_25_0.cap_res_X.t71 two_stage_opamp_dummy_magic_25_0.cap_res_X.t39 0.1603
R465 two_stage_opamp_dummy_magic_25_0.cap_res_X.t52 two_stage_opamp_dummy_magic_25_0.cap_res_X.t10 0.1603
R466 two_stage_opamp_dummy_magic_25_0.cap_res_X.t77 two_stage_opamp_dummy_magic_25_0.cap_res_X.t37 0.1603
R467 two_stage_opamp_dummy_magic_25_0.cap_res_X.t55 two_stage_opamp_dummy_magic_25_0.cap_res_X.t17 0.1603
R468 two_stage_opamp_dummy_magic_25_0.cap_res_X.t21 two_stage_opamp_dummy_magic_25_0.cap_res_X.t118 0.1603
R469 two_stage_opamp_dummy_magic_25_0.cap_res_X.t44 two_stage_opamp_dummy_magic_25_0.cap_res_X.t2 0.1603
R470 two_stage_opamp_dummy_magic_25_0.cap_res_X.t4 two_stage_opamp_dummy_magic_25_0.cap_res_X.t100 0.1603
R471 two_stage_opamp_dummy_magic_25_0.cap_res_X.t105 two_stage_opamp_dummy_magic_25_0.cap_res_X.t65 0.1603
R472 two_stage_opamp_dummy_magic_25_0.cap_res_X.t67 two_stage_opamp_dummy_magic_25_0.cap_res_X.t29 0.1603
R473 two_stage_opamp_dummy_magic_25_0.cap_res_X.t88 two_stage_opamp_dummy_magic_25_0.cap_res_X.t49 0.1603
R474 two_stage_opamp_dummy_magic_25_0.cap_res_X.t51 two_stage_opamp_dummy_magic_25_0.cap_res_X.t8 0.1603
R475 two_stage_opamp_dummy_magic_25_0.cap_res_X.t12 two_stage_opamp_dummy_magic_25_0.cap_res_X.t111 0.1603
R476 two_stage_opamp_dummy_magic_25_0.cap_res_X.t136 two_stage_opamp_dummy_magic_25_0.cap_res_X.t98 0.1603
R477 two_stage_opamp_dummy_magic_25_0.cap_res_X.t93 two_stage_opamp_dummy_magic_25_0.cap_res_X.t60 0.1603
R478 two_stage_opamp_dummy_magic_25_0.cap_res_X.t7 two_stage_opamp_dummy_magic_25_0.cap_res_X.t110 0.1603
R479 two_stage_opamp_dummy_magic_25_0.cap_res_X.t11 two_stage_opamp_dummy_magic_25_0.cap_res_X.t102 0.1603
R480 two_stage_opamp_dummy_magic_25_0.cap_res_X.t47 two_stage_opamp_dummy_magic_25_0.cap_res_X.t11 0.1603
R481 two_stage_opamp_dummy_magic_25_0.cap_res_X.t131 two_stage_opamp_dummy_magic_25_0.cap_res_X.t28 0.1603
R482 two_stage_opamp_dummy_magic_25_0.cap_res_X.t15 two_stage_opamp_dummy_magic_25_0.cap_res_X.t131 0.1603
R483 two_stage_opamp_dummy_magic_25_0.cap_res_X.t38 two_stage_opamp_dummy_magic_25_0.cap_res_X.n10 0.159278
R484 two_stage_opamp_dummy_magic_25_0.cap_res_X.t106 two_stage_opamp_dummy_magic_25_0.cap_res_X.n11 0.159278
R485 two_stage_opamp_dummy_magic_25_0.cap_res_X.t72 two_stage_opamp_dummy_magic_25_0.cap_res_X.n12 0.159278
R486 two_stage_opamp_dummy_magic_25_0.cap_res_X.t135 two_stage_opamp_dummy_magic_25_0.cap_res_X.n13 0.159278
R487 two_stage_opamp_dummy_magic_25_0.cap_res_X.t26 two_stage_opamp_dummy_magic_25_0.cap_res_X.n14 0.159278
R488 two_stage_opamp_dummy_magic_25_0.cap_res_X.t57 two_stage_opamp_dummy_magic_25_0.cap_res_X.n15 0.159278
R489 two_stage_opamp_dummy_magic_25_0.cap_res_X.t18 two_stage_opamp_dummy_magic_25_0.cap_res_X.n16 0.159278
R490 two_stage_opamp_dummy_magic_25_0.cap_res_X.t117 two_stage_opamp_dummy_magic_25_0.cap_res_X.n17 0.159278
R491 two_stage_opamp_dummy_magic_25_0.cap_res_X.t13 two_stage_opamp_dummy_magic_25_0.cap_res_X.n18 0.159278
R492 two_stage_opamp_dummy_magic_25_0.cap_res_X.t112 two_stage_opamp_dummy_magic_25_0.cap_res_X.n19 0.159278
R493 two_stage_opamp_dummy_magic_25_0.cap_res_X.t73 two_stage_opamp_dummy_magic_25_0.cap_res_X.n20 0.159278
R494 two_stage_opamp_dummy_magic_25_0.cap_res_X.t35 two_stage_opamp_dummy_magic_25_0.cap_res_X.n21 0.159278
R495 two_stage_opamp_dummy_magic_25_0.cap_res_X.t68 two_stage_opamp_dummy_magic_25_0.cap_res_X.n22 0.159278
R496 two_stage_opamp_dummy_magic_25_0.cap_res_X.t30 two_stage_opamp_dummy_magic_25_0.cap_res_X.n23 0.159278
R497 two_stage_opamp_dummy_magic_25_0.cap_res_X.t130 two_stage_opamp_dummy_magic_25_0.cap_res_X.n24 0.159278
R498 two_stage_opamp_dummy_magic_25_0.cap_res_X.t25 two_stage_opamp_dummy_magic_25_0.cap_res_X.n25 0.159278
R499 two_stage_opamp_dummy_magic_25_0.cap_res_X.t124 two_stage_opamp_dummy_magic_25_0.cap_res_X.n26 0.159278
R500 two_stage_opamp_dummy_magic_25_0.cap_res_X.t96 two_stage_opamp_dummy_magic_25_0.cap_res_X.n27 0.159278
R501 two_stage_opamp_dummy_magic_25_0.cap_res_X.t133 two_stage_opamp_dummy_magic_25_0.cap_res_X.n28 0.159278
R502 two_stage_opamp_dummy_magic_25_0.cap_res_X.n31 two_stage_opamp_dummy_magic_25_0.cap_res_X.t16 0.1368
R503 two_stage_opamp_dummy_magic_25_0.cap_res_X.n29 two_stage_opamp_dummy_magic_25_0.cap_res_X.t92 0.1368
R504 two_stage_opamp_dummy_magic_25_0.cap_res_X.n28 two_stage_opamp_dummy_magic_25_0.cap_res_X.t78 0.1368
R505 two_stage_opamp_dummy_magic_25_0.cap_res_X.n28 two_stage_opamp_dummy_magic_25_0.cap_res_X.t61 0.1368
R506 two_stage_opamp_dummy_magic_25_0.cap_res_X.n27 two_stage_opamp_dummy_magic_25_0.cap_res_X.t36 0.1368
R507 two_stage_opamp_dummy_magic_25_0.cap_res_X.n27 two_stage_opamp_dummy_magic_25_0.cap_res_X.t87 0.1368
R508 two_stage_opamp_dummy_magic_25_0.cap_res_X.n26 two_stage_opamp_dummy_magic_25_0.cap_res_X.t74 0.1368
R509 two_stage_opamp_dummy_magic_25_0.cap_res_X.n26 two_stage_opamp_dummy_magic_25_0.cap_res_X.t129 0.1368
R510 two_stage_opamp_dummy_magic_25_0.cap_res_X.n25 two_stage_opamp_dummy_magic_25_0.cap_res_X.t43 0.1368
R511 two_stage_opamp_dummy_magic_25_0.cap_res_X.n25 two_stage_opamp_dummy_magic_25_0.cap_res_X.t91 0.1368
R512 two_stage_opamp_dummy_magic_25_0.cap_res_X.n24 two_stage_opamp_dummy_magic_25_0.cap_res_X.t80 0.1368
R513 two_stage_opamp_dummy_magic_25_0.cap_res_X.n24 two_stage_opamp_dummy_magic_25_0.cap_res_X.t132 0.1368
R514 two_stage_opamp_dummy_magic_25_0.cap_res_X.n23 two_stage_opamp_dummy_magic_25_0.cap_res_X.t119 0.1368
R515 two_stage_opamp_dummy_magic_25_0.cap_res_X.n23 two_stage_opamp_dummy_magic_25_0.cap_res_X.t33 0.1368
R516 two_stage_opamp_dummy_magic_25_0.cap_res_X.n22 two_stage_opamp_dummy_magic_25_0.cap_res_X.t84 0.1368
R517 two_stage_opamp_dummy_magic_25_0.cap_res_X.n22 two_stage_opamp_dummy_magic_25_0.cap_res_X.t0 0.1368
R518 two_stage_opamp_dummy_magic_25_0.cap_res_X.n21 two_stage_opamp_dummy_magic_25_0.cap_res_X.t125 0.1368
R519 two_stage_opamp_dummy_magic_25_0.cap_res_X.n21 two_stage_opamp_dummy_magic_25_0.cap_res_X.t41 0.1368
R520 two_stage_opamp_dummy_magic_25_0.cap_res_X.n20 two_stage_opamp_dummy_magic_25_0.cap_res_X.t27 0.1368
R521 two_stage_opamp_dummy_magic_25_0.cap_res_X.n20 two_stage_opamp_dummy_magic_25_0.cap_res_X.t79 0.1368
R522 two_stage_opamp_dummy_magic_25_0.cap_res_X.n19 two_stage_opamp_dummy_magic_25_0.cap_res_X.t63 0.1368
R523 two_stage_opamp_dummy_magic_25_0.cap_res_X.n19 two_stage_opamp_dummy_magic_25_0.cap_res_X.t116 0.1368
R524 two_stage_opamp_dummy_magic_25_0.cap_res_X.n18 two_stage_opamp_dummy_magic_25_0.cap_res_X.t32 0.1368
R525 two_stage_opamp_dummy_magic_25_0.cap_res_X.n18 two_stage_opamp_dummy_magic_25_0.cap_res_X.t83 0.1368
R526 two_stage_opamp_dummy_magic_25_0.cap_res_X.n17 two_stage_opamp_dummy_magic_25_0.cap_res_X.t69 0.1368
R527 two_stage_opamp_dummy_magic_25_0.cap_res_X.n17 two_stage_opamp_dummy_magic_25_0.cap_res_X.t122 0.1368
R528 two_stage_opamp_dummy_magic_25_0.cap_res_X.n16 two_stage_opamp_dummy_magic_25_0.cap_res_X.t107 0.1368
R529 two_stage_opamp_dummy_magic_25_0.cap_res_X.n16 two_stage_opamp_dummy_magic_25_0.cap_res_X.t23 0.1368
R530 two_stage_opamp_dummy_magic_25_0.cap_res_X.n15 two_stage_opamp_dummy_magic_25_0.cap_res_X.t75 0.1368
R531 two_stage_opamp_dummy_magic_25_0.cap_res_X.n15 two_stage_opamp_dummy_magic_25_0.cap_res_X.t128 0.1368
R532 two_stage_opamp_dummy_magic_25_0.cap_res_X.n14 two_stage_opamp_dummy_magic_25_0.cap_res_X.t42 0.1368
R533 two_stage_opamp_dummy_magic_25_0.cap_res_X.n14 two_stage_opamp_dummy_magic_25_0.cap_res_X.t46 0.1368
R534 two_stage_opamp_dummy_magic_25_0.cap_res_X.n13 two_stage_opamp_dummy_magic_25_0.cap_res_X.t123 0.1368
R535 two_stage_opamp_dummy_magic_25_0.cap_res_X.n13 two_stage_opamp_dummy_magic_25_0.cap_res_X.t40 0.1368
R536 two_stage_opamp_dummy_magic_25_0.cap_res_X.n12 two_stage_opamp_dummy_magic_25_0.cap_res_X.t19 0.1368
R537 two_stage_opamp_dummy_magic_25_0.cap_res_X.n12 two_stage_opamp_dummy_magic_25_0.cap_res_X.t71 0.1368
R538 two_stage_opamp_dummy_magic_25_0.cap_res_X.n11 two_stage_opamp_dummy_magic_25_0.cap_res_X.t136 0.1368
R539 two_stage_opamp_dummy_magic_25_0.cap_res_X.n10 two_stage_opamp_dummy_magic_25_0.cap_res_X.t93 0.1368
R540 two_stage_opamp_dummy_magic_25_0.cap_res_X.t110 two_stage_opamp_dummy_magic_25_0.cap_res_X.n29 0.1368
R541 two_stage_opamp_dummy_magic_25_0.cap_res_X.n30 two_stage_opamp_dummy_magic_25_0.cap_res_X.t7 0.1368
R542 two_stage_opamp_dummy_magic_25_0.cap_res_X.n0 two_stage_opamp_dummy_magic_25_0.cap_res_X.t52 0.114322
R543 two_stage_opamp_dummy_magic_25_0.cap_res_X.n32 two_stage_opamp_dummy_magic_25_0.cap_res_X.n31 0.1133
R544 two_stage_opamp_dummy_magic_25_0.cap_res_X.n33 two_stage_opamp_dummy_magic_25_0.cap_res_X.n32 0.1133
R545 two_stage_opamp_dummy_magic_25_0.cap_res_X.n34 two_stage_opamp_dummy_magic_25_0.cap_res_X.n33 0.1133
R546 two_stage_opamp_dummy_magic_25_0.cap_res_X.n1 two_stage_opamp_dummy_magic_25_0.cap_res_X.n0 0.1133
R547 two_stage_opamp_dummy_magic_25_0.cap_res_X.n2 two_stage_opamp_dummy_magic_25_0.cap_res_X.n1 0.1133
R548 two_stage_opamp_dummy_magic_25_0.cap_res_X.n3 two_stage_opamp_dummy_magic_25_0.cap_res_X.n2 0.1133
R549 two_stage_opamp_dummy_magic_25_0.cap_res_X.n4 two_stage_opamp_dummy_magic_25_0.cap_res_X.n3 0.1133
R550 two_stage_opamp_dummy_magic_25_0.cap_res_X.n5 two_stage_opamp_dummy_magic_25_0.cap_res_X.n4 0.1133
R551 two_stage_opamp_dummy_magic_25_0.cap_res_X.n6 two_stage_opamp_dummy_magic_25_0.cap_res_X.n5 0.1133
R552 two_stage_opamp_dummy_magic_25_0.cap_res_X.n7 two_stage_opamp_dummy_magic_25_0.cap_res_X.n6 0.1133
R553 two_stage_opamp_dummy_magic_25_0.cap_res_X.n8 two_stage_opamp_dummy_magic_25_0.cap_res_X.n7 0.1133
R554 two_stage_opamp_dummy_magic_25_0.cap_res_X.n9 two_stage_opamp_dummy_magic_25_0.cap_res_X.n8 0.1133
R555 two_stage_opamp_dummy_magic_25_0.cap_res_X.n11 two_stage_opamp_dummy_magic_25_0.cap_res_X.n9 0.1133
R556 two_stage_opamp_dummy_magic_25_0.cap_res_X.n35 two_stage_opamp_dummy_magic_25_0.cap_res_X.n30 0.1133
R557 two_stage_opamp_dummy_magic_25_0.cap_res_X.n35 two_stage_opamp_dummy_magic_25_0.cap_res_X.n34 0.1133
R558 two_stage_opamp_dummy_magic_25_0.cap_res_X.n31 two_stage_opamp_dummy_magic_25_0.cap_res_X.t115 0.00152174
R559 two_stage_opamp_dummy_magic_25_0.cap_res_X.n32 two_stage_opamp_dummy_magic_25_0.cap_res_X.t1 0.00152174
R560 two_stage_opamp_dummy_magic_25_0.cap_res_X.n33 two_stage_opamp_dummy_magic_25_0.cap_res_X.t99 0.00152174
R561 two_stage_opamp_dummy_magic_25_0.cap_res_X.n34 two_stage_opamp_dummy_magic_25_0.cap_res_X.t62 0.00152174
R562 two_stage_opamp_dummy_magic_25_0.cap_res_X.n0 two_stage_opamp_dummy_magic_25_0.cap_res_X.t77 0.00152174
R563 two_stage_opamp_dummy_magic_25_0.cap_res_X.n1 two_stage_opamp_dummy_magic_25_0.cap_res_X.t55 0.00152174
R564 two_stage_opamp_dummy_magic_25_0.cap_res_X.n2 two_stage_opamp_dummy_magic_25_0.cap_res_X.t21 0.00152174
R565 two_stage_opamp_dummy_magic_25_0.cap_res_X.n3 two_stage_opamp_dummy_magic_25_0.cap_res_X.t44 0.00152174
R566 two_stage_opamp_dummy_magic_25_0.cap_res_X.n4 two_stage_opamp_dummy_magic_25_0.cap_res_X.t4 0.00152174
R567 two_stage_opamp_dummy_magic_25_0.cap_res_X.n5 two_stage_opamp_dummy_magic_25_0.cap_res_X.t105 0.00152174
R568 two_stage_opamp_dummy_magic_25_0.cap_res_X.n6 two_stage_opamp_dummy_magic_25_0.cap_res_X.t67 0.00152174
R569 two_stage_opamp_dummy_magic_25_0.cap_res_X.n7 two_stage_opamp_dummy_magic_25_0.cap_res_X.t88 0.00152174
R570 two_stage_opamp_dummy_magic_25_0.cap_res_X.n8 two_stage_opamp_dummy_magic_25_0.cap_res_X.t51 0.00152174
R571 two_stage_opamp_dummy_magic_25_0.cap_res_X.n9 two_stage_opamp_dummy_magic_25_0.cap_res_X.t12 0.00152174
R572 two_stage_opamp_dummy_magic_25_0.cap_res_X.n10 two_stage_opamp_dummy_magic_25_0.cap_res_X.t134 0.00152174
R573 two_stage_opamp_dummy_magic_25_0.cap_res_X.n11 two_stage_opamp_dummy_magic_25_0.cap_res_X.t38 0.00152174
R574 two_stage_opamp_dummy_magic_25_0.cap_res_X.n12 two_stage_opamp_dummy_magic_25_0.cap_res_X.t106 0.00152174
R575 two_stage_opamp_dummy_magic_25_0.cap_res_X.n13 two_stage_opamp_dummy_magic_25_0.cap_res_X.t72 0.00152174
R576 two_stage_opamp_dummy_magic_25_0.cap_res_X.n14 two_stage_opamp_dummy_magic_25_0.cap_res_X.t135 0.00152174
R577 two_stage_opamp_dummy_magic_25_0.cap_res_X.n15 two_stage_opamp_dummy_magic_25_0.cap_res_X.t26 0.00152174
R578 two_stage_opamp_dummy_magic_25_0.cap_res_X.n16 two_stage_opamp_dummy_magic_25_0.cap_res_X.t57 0.00152174
R579 two_stage_opamp_dummy_magic_25_0.cap_res_X.n17 two_stage_opamp_dummy_magic_25_0.cap_res_X.t18 0.00152174
R580 two_stage_opamp_dummy_magic_25_0.cap_res_X.n18 two_stage_opamp_dummy_magic_25_0.cap_res_X.t117 0.00152174
R581 two_stage_opamp_dummy_magic_25_0.cap_res_X.n19 two_stage_opamp_dummy_magic_25_0.cap_res_X.t13 0.00152174
R582 two_stage_opamp_dummy_magic_25_0.cap_res_X.n20 two_stage_opamp_dummy_magic_25_0.cap_res_X.t112 0.00152174
R583 two_stage_opamp_dummy_magic_25_0.cap_res_X.n21 two_stage_opamp_dummy_magic_25_0.cap_res_X.t73 0.00152174
R584 two_stage_opamp_dummy_magic_25_0.cap_res_X.n22 two_stage_opamp_dummy_magic_25_0.cap_res_X.t35 0.00152174
R585 two_stage_opamp_dummy_magic_25_0.cap_res_X.n23 two_stage_opamp_dummy_magic_25_0.cap_res_X.t68 0.00152174
R586 two_stage_opamp_dummy_magic_25_0.cap_res_X.n24 two_stage_opamp_dummy_magic_25_0.cap_res_X.t30 0.00152174
R587 two_stage_opamp_dummy_magic_25_0.cap_res_X.n25 two_stage_opamp_dummy_magic_25_0.cap_res_X.t130 0.00152174
R588 two_stage_opamp_dummy_magic_25_0.cap_res_X.n26 two_stage_opamp_dummy_magic_25_0.cap_res_X.t25 0.00152174
R589 two_stage_opamp_dummy_magic_25_0.cap_res_X.n27 two_stage_opamp_dummy_magic_25_0.cap_res_X.t124 0.00152174
R590 two_stage_opamp_dummy_magic_25_0.cap_res_X.n28 two_stage_opamp_dummy_magic_25_0.cap_res_X.t96 0.00152174
R591 two_stage_opamp_dummy_magic_25_0.cap_res_X.n29 two_stage_opamp_dummy_magic_25_0.cap_res_X.t133 0.00152174
R592 two_stage_opamp_dummy_magic_25_0.cap_res_X.n30 two_stage_opamp_dummy_magic_25_0.cap_res_X.t47 0.00152174
R593 two_stage_opamp_dummy_magic_25_0.cap_res_X.t28 two_stage_opamp_dummy_magic_25_0.cap_res_X.n35 0.00152174
R594 two_stage_opamp_dummy_magic_25_0.Vb3.n25 two_stage_opamp_dummy_magic_25_0.Vb3.t24 768.551
R595 two_stage_opamp_dummy_magic_25_0.Vb3.n19 two_stage_opamp_dummy_magic_25_0.Vb3.t18 611.739
R596 two_stage_opamp_dummy_magic_25_0.Vb3.n15 two_stage_opamp_dummy_magic_25_0.Vb3.t8 611.739
R597 two_stage_opamp_dummy_magic_25_0.Vb3.n10 two_stage_opamp_dummy_magic_25_0.Vb3.t22 611.739
R598 two_stage_opamp_dummy_magic_25_0.Vb3.n6 two_stage_opamp_dummy_magic_25_0.Vb3.t16 611.739
R599 two_stage_opamp_dummy_magic_25_0.Vb3.n24 two_stage_opamp_dummy_magic_25_0.Vb3.n23 431.07
R600 two_stage_opamp_dummy_magic_25_0.Vb3.n24 two_stage_opamp_dummy_magic_25_0.Vb3.n14 430.507
R601 two_stage_opamp_dummy_magic_25_0.Vb3.n19 two_stage_opamp_dummy_magic_25_0.Vb3.t12 421.75
R602 two_stage_opamp_dummy_magic_25_0.Vb3.n20 two_stage_opamp_dummy_magic_25_0.Vb3.t28 421.75
R603 two_stage_opamp_dummy_magic_25_0.Vb3.n21 two_stage_opamp_dummy_magic_25_0.Vb3.t10 421.75
R604 two_stage_opamp_dummy_magic_25_0.Vb3.n22 two_stage_opamp_dummy_magic_25_0.Vb3.t27 421.75
R605 two_stage_opamp_dummy_magic_25_0.Vb3.n15 two_stage_opamp_dummy_magic_25_0.Vb3.t14 421.75
R606 two_stage_opamp_dummy_magic_25_0.Vb3.n16 two_stage_opamp_dummy_magic_25_0.Vb3.t11 421.75
R607 two_stage_opamp_dummy_magic_25_0.Vb3.n17 two_stage_opamp_dummy_magic_25_0.Vb3.t17 421.75
R608 two_stage_opamp_dummy_magic_25_0.Vb3.n18 two_stage_opamp_dummy_magic_25_0.Vb3.t25 421.75
R609 two_stage_opamp_dummy_magic_25_0.Vb3.n10 two_stage_opamp_dummy_magic_25_0.Vb3.t20 421.75
R610 two_stage_opamp_dummy_magic_25_0.Vb3.n11 two_stage_opamp_dummy_magic_25_0.Vb3.t15 421.75
R611 two_stage_opamp_dummy_magic_25_0.Vb3.n12 two_stage_opamp_dummy_magic_25_0.Vb3.t9 421.75
R612 two_stage_opamp_dummy_magic_25_0.Vb3.n13 two_stage_opamp_dummy_magic_25_0.Vb3.t26 421.75
R613 two_stage_opamp_dummy_magic_25_0.Vb3.n6 two_stage_opamp_dummy_magic_25_0.Vb3.t13 421.75
R614 two_stage_opamp_dummy_magic_25_0.Vb3.n7 two_stage_opamp_dummy_magic_25_0.Vb3.t19 421.75
R615 two_stage_opamp_dummy_magic_25_0.Vb3.n8 two_stage_opamp_dummy_magic_25_0.Vb3.t21 421.75
R616 two_stage_opamp_dummy_magic_25_0.Vb3.n9 two_stage_opamp_dummy_magic_25_0.Vb3.t23 421.75
R617 two_stage_opamp_dummy_magic_25_0.Vb3.n20 two_stage_opamp_dummy_magic_25_0.Vb3.n19 167.094
R618 two_stage_opamp_dummy_magic_25_0.Vb3.n21 two_stage_opamp_dummy_magic_25_0.Vb3.n20 167.094
R619 two_stage_opamp_dummy_magic_25_0.Vb3.n22 two_stage_opamp_dummy_magic_25_0.Vb3.n21 167.094
R620 two_stage_opamp_dummy_magic_25_0.Vb3.n16 two_stage_opamp_dummy_magic_25_0.Vb3.n15 167.094
R621 two_stage_opamp_dummy_magic_25_0.Vb3.n17 two_stage_opamp_dummy_magic_25_0.Vb3.n16 167.094
R622 two_stage_opamp_dummy_magic_25_0.Vb3.n18 two_stage_opamp_dummy_magic_25_0.Vb3.n17 167.094
R623 two_stage_opamp_dummy_magic_25_0.Vb3.n11 two_stage_opamp_dummy_magic_25_0.Vb3.n10 167.094
R624 two_stage_opamp_dummy_magic_25_0.Vb3.n12 two_stage_opamp_dummy_magic_25_0.Vb3.n11 167.094
R625 two_stage_opamp_dummy_magic_25_0.Vb3.n13 two_stage_opamp_dummy_magic_25_0.Vb3.n12 167.094
R626 two_stage_opamp_dummy_magic_25_0.Vb3.n7 two_stage_opamp_dummy_magic_25_0.Vb3.n6 167.094
R627 two_stage_opamp_dummy_magic_25_0.Vb3.n8 two_stage_opamp_dummy_magic_25_0.Vb3.n7 167.094
R628 two_stage_opamp_dummy_magic_25_0.Vb3.n9 two_stage_opamp_dummy_magic_25_0.Vb3.n8 167.094
R629 two_stage_opamp_dummy_magic_25_0.Vb3.n2 two_stage_opamp_dummy_magic_25_0.Vb3.n0 139.639
R630 two_stage_opamp_dummy_magic_25_0.Vb3.n2 two_stage_opamp_dummy_magic_25_0.Vb3.n1 139.638
R631 two_stage_opamp_dummy_magic_25_0.Vb3.n4 two_stage_opamp_dummy_magic_25_0.Vb3.n3 134.577
R632 two_stage_opamp_dummy_magic_25_0.Vb3.n26 two_stage_opamp_dummy_magic_25_0.Vb3.n5 73.3081
R633 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_25_0.Vb3.n26 68.0005
R634 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_25_0.Vb3.n4 42.1255
R635 two_stage_opamp_dummy_magic_25_0.Vb3.n23 two_stage_opamp_dummy_magic_25_0.Vb3.n22 35.3472
R636 two_stage_opamp_dummy_magic_25_0.Vb3.n23 two_stage_opamp_dummy_magic_25_0.Vb3.n18 35.3472
R637 two_stage_opamp_dummy_magic_25_0.Vb3.n14 two_stage_opamp_dummy_magic_25_0.Vb3.n13 35.3472
R638 two_stage_opamp_dummy_magic_25_0.Vb3.n14 two_stage_opamp_dummy_magic_25_0.Vb3.n9 35.3472
R639 two_stage_opamp_dummy_magic_25_0.Vb3.n3 two_stage_opamp_dummy_magic_25_0.Vb3.t5 24.0005
R640 two_stage_opamp_dummy_magic_25_0.Vb3.n3 two_stage_opamp_dummy_magic_25_0.Vb3.t1 24.0005
R641 two_stage_opamp_dummy_magic_25_0.Vb3.n1 two_stage_opamp_dummy_magic_25_0.Vb3.t3 24.0005
R642 two_stage_opamp_dummy_magic_25_0.Vb3.n1 two_stage_opamp_dummy_magic_25_0.Vb3.t2 24.0005
R643 two_stage_opamp_dummy_magic_25_0.Vb3.n0 two_stage_opamp_dummy_magic_25_0.Vb3.t7 24.0005
R644 two_stage_opamp_dummy_magic_25_0.Vb3.n0 two_stage_opamp_dummy_magic_25_0.Vb3.t4 24.0005
R645 two_stage_opamp_dummy_magic_25_0.Vb3.n25 two_stage_opamp_dummy_magic_25_0.Vb3.n24 15.563
R646 two_stage_opamp_dummy_magic_25_0.Vb3.n5 two_stage_opamp_dummy_magic_25_0.Vb3.t0 11.2576
R647 two_stage_opamp_dummy_magic_25_0.Vb3.n5 two_stage_opamp_dummy_magic_25_0.Vb3.t6 11.2576
R648 two_stage_opamp_dummy_magic_25_0.Vb3.n4 two_stage_opamp_dummy_magic_25_0.Vb3.n2 4.5005
R649 two_stage_opamp_dummy_magic_25_0.Vb3.n26 two_stage_opamp_dummy_magic_25_0.Vb3.n25 1.21231
R650 two_stage_opamp_dummy_magic_25_0.VD4.n35 two_stage_opamp_dummy_magic_25_0.VD4.t32 672.293
R651 two_stage_opamp_dummy_magic_25_0.VD4.n32 two_stage_opamp_dummy_magic_25_0.VD4.t29 672.293
R652 two_stage_opamp_dummy_magic_25_0.VD4.t30 two_stage_opamp_dummy_magic_25_0.VD4.n33 213.131
R653 two_stage_opamp_dummy_magic_25_0.VD4.n34 two_stage_opamp_dummy_magic_25_0.VD4.t33 213.131
R654 two_stage_opamp_dummy_magic_25_0.VD4.t17 two_stage_opamp_dummy_magic_25_0.VD4.t30 146.155
R655 two_stage_opamp_dummy_magic_25_0.VD4.t9 two_stage_opamp_dummy_magic_25_0.VD4.t17 146.155
R656 two_stage_opamp_dummy_magic_25_0.VD4.t1 two_stage_opamp_dummy_magic_25_0.VD4.t9 146.155
R657 two_stage_opamp_dummy_magic_25_0.VD4.t11 two_stage_opamp_dummy_magic_25_0.VD4.t1 146.155
R658 two_stage_opamp_dummy_magic_25_0.VD4.t35 two_stage_opamp_dummy_magic_25_0.VD4.t11 146.155
R659 two_stage_opamp_dummy_magic_25_0.VD4.t15 two_stage_opamp_dummy_magic_25_0.VD4.t35 146.155
R660 two_stage_opamp_dummy_magic_25_0.VD4.t3 two_stage_opamp_dummy_magic_25_0.VD4.t15 146.155
R661 two_stage_opamp_dummy_magic_25_0.VD4.t5 two_stage_opamp_dummy_magic_25_0.VD4.t3 146.155
R662 two_stage_opamp_dummy_magic_25_0.VD4.t13 two_stage_opamp_dummy_magic_25_0.VD4.t5 146.155
R663 two_stage_opamp_dummy_magic_25_0.VD4.t7 two_stage_opamp_dummy_magic_25_0.VD4.t13 146.155
R664 two_stage_opamp_dummy_magic_25_0.VD4.t33 two_stage_opamp_dummy_magic_25_0.VD4.t7 146.155
R665 two_stage_opamp_dummy_magic_25_0.VD4.n33 two_stage_opamp_dummy_magic_25_0.VD4.t31 76.2576
R666 two_stage_opamp_dummy_magic_25_0.VD4.n34 two_stage_opamp_dummy_magic_25_0.VD4.t34 76.2576
R667 two_stage_opamp_dummy_magic_25_0.VD4.n2 two_stage_opamp_dummy_magic_25_0.VD4.n31 66.9922
R668 two_stage_opamp_dummy_magic_25_0.VD4.n2 two_stage_opamp_dummy_magic_25_0.VD4.n9 66.9922
R669 two_stage_opamp_dummy_magic_25_0.VD4.n2 two_stage_opamp_dummy_magic_25_0.VD4.n10 66.9922
R670 two_stage_opamp_dummy_magic_25_0.VD4.n4 two_stage_opamp_dummy_magic_25_0.VD4.n11 66.9922
R671 two_stage_opamp_dummy_magic_25_0.VD4.n36 two_stage_opamp_dummy_magic_25_0.VD4.n2 66.9922
R672 two_stage_opamp_dummy_magic_25_0.VD4.n16 two_stage_opamp_dummy_magic_25_0.VD4.n15 66.0338
R673 two_stage_opamp_dummy_magic_25_0.VD4.n18 two_stage_opamp_dummy_magic_25_0.VD4.n17 66.0338
R674 two_stage_opamp_dummy_magic_25_0.VD4.n26 two_stage_opamp_dummy_magic_25_0.VD4.n25 66.0338
R675 two_stage_opamp_dummy_magic_25_0.VD4.n29 two_stage_opamp_dummy_magic_25_0.VD4.n28 66.0338
R676 two_stage_opamp_dummy_magic_25_0.VD4.n21 two_stage_opamp_dummy_magic_25_0.VD4.n20 66.0338
R677 two_stage_opamp_dummy_magic_25_0.VD4.n13 two_stage_opamp_dummy_magic_25_0.VD4.n12 66.0338
R678 two_stage_opamp_dummy_magic_25_0.VD4.n31 two_stage_opamp_dummy_magic_25_0.VD4.t18 11.2576
R679 two_stage_opamp_dummy_magic_25_0.VD4.n31 two_stage_opamp_dummy_magic_25_0.VD4.t10 11.2576
R680 two_stage_opamp_dummy_magic_25_0.VD4.n9 two_stage_opamp_dummy_magic_25_0.VD4.t36 11.2576
R681 two_stage_opamp_dummy_magic_25_0.VD4.n9 two_stage_opamp_dummy_magic_25_0.VD4.t16 11.2576
R682 two_stage_opamp_dummy_magic_25_0.VD4.n10 two_stage_opamp_dummy_magic_25_0.VD4.t4 11.2576
R683 two_stage_opamp_dummy_magic_25_0.VD4.n10 two_stage_opamp_dummy_magic_25_0.VD4.t6 11.2576
R684 two_stage_opamp_dummy_magic_25_0.VD4.n11 two_stage_opamp_dummy_magic_25_0.VD4.t14 11.2576
R685 two_stage_opamp_dummy_magic_25_0.VD4.n11 two_stage_opamp_dummy_magic_25_0.VD4.t8 11.2576
R686 two_stage_opamp_dummy_magic_25_0.VD4.n15 two_stage_opamp_dummy_magic_25_0.VD4.t28 11.2576
R687 two_stage_opamp_dummy_magic_25_0.VD4.n15 two_stage_opamp_dummy_magic_25_0.VD4.t20 11.2576
R688 two_stage_opamp_dummy_magic_25_0.VD4.n17 two_stage_opamp_dummy_magic_25_0.VD4.t23 11.2576
R689 two_stage_opamp_dummy_magic_25_0.VD4.n17 two_stage_opamp_dummy_magic_25_0.VD4.t22 11.2576
R690 two_stage_opamp_dummy_magic_25_0.VD4.n25 two_stage_opamp_dummy_magic_25_0.VD4.t27 11.2576
R691 two_stage_opamp_dummy_magic_25_0.VD4.n25 two_stage_opamp_dummy_magic_25_0.VD4.t19 11.2576
R692 two_stage_opamp_dummy_magic_25_0.VD4.n28 two_stage_opamp_dummy_magic_25_0.VD4.t25 11.2576
R693 two_stage_opamp_dummy_magic_25_0.VD4.n28 two_stage_opamp_dummy_magic_25_0.VD4.t0 11.2576
R694 two_stage_opamp_dummy_magic_25_0.VD4.n20 two_stage_opamp_dummy_magic_25_0.VD4.t26 11.2576
R695 two_stage_opamp_dummy_magic_25_0.VD4.n20 two_stage_opamp_dummy_magic_25_0.VD4.t24 11.2576
R696 two_stage_opamp_dummy_magic_25_0.VD4.n12 two_stage_opamp_dummy_magic_25_0.VD4.t37 11.2576
R697 two_stage_opamp_dummy_magic_25_0.VD4.n12 two_stage_opamp_dummy_magic_25_0.VD4.t21 11.2576
R698 two_stage_opamp_dummy_magic_25_0.VD4.t2 two_stage_opamp_dummy_magic_25_0.VD4.n36 11.2576
R699 two_stage_opamp_dummy_magic_25_0.VD4.n36 two_stage_opamp_dummy_magic_25_0.VD4.t12 11.2576
R700 two_stage_opamp_dummy_magic_25_0.VD4.n29 two_stage_opamp_dummy_magic_25_0.VD4.n27 5.91717
R701 two_stage_opamp_dummy_magic_25_0.VD4.n22 two_stage_opamp_dummy_magic_25_0.VD4.n13 5.91717
R702 two_stage_opamp_dummy_magic_25_0.VD4.n24 two_stage_opamp_dummy_magic_25_0.VD4.n18 5.29217
R703 two_stage_opamp_dummy_magic_25_0.VD4.n27 two_stage_opamp_dummy_magic_25_0.VD4.n26 5.29217
R704 two_stage_opamp_dummy_magic_25_0.VD4.n22 two_stage_opamp_dummy_magic_25_0.VD4.n21 5.29217
R705 two_stage_opamp_dummy_magic_25_0.VD4.n23 two_stage_opamp_dummy_magic_25_0.VD4.n16 5.29217
R706 two_stage_opamp_dummy_magic_25_0.VD4.n1 two_stage_opamp_dummy_magic_25_0.VD4.n7 0.351294
R707 two_stage_opamp_dummy_magic_25_0.VD4.n1 two_stage_opamp_dummy_magic_25_0.VD4.n8 0.48314
R708 two_stage_opamp_dummy_magic_25_0.VD4.n6 two_stage_opamp_dummy_magic_25_0.VD4.n0 0.48314
R709 two_stage_opamp_dummy_magic_25_0.VD4.n4 two_stage_opamp_dummy_magic_25_0.VD4.n5 0.214731
R710 two_stage_opamp_dummy_magic_25_0.VD4.n2 two_stage_opamp_dummy_magic_25_0.VD4.n3 0.0894566
R711 two_stage_opamp_dummy_magic_25_0.VD4.n33 two_stage_opamp_dummy_magic_25_0.VD4.n32 1.03383
R712 two_stage_opamp_dummy_magic_25_0.VD4.n35 two_stage_opamp_dummy_magic_25_0.VD4.n34 1.03383
R713 two_stage_opamp_dummy_magic_25_0.VD4.n30 two_stage_opamp_dummy_magic_25_0.VD4.n29 1.02322
R714 two_stage_opamp_dummy_magic_25_0.VD4.n4 two_stage_opamp_dummy_magic_25_0.VD4.n35 0.958833
R715 two_stage_opamp_dummy_magic_25_0.VD4.n6 two_stage_opamp_dummy_magic_25_0.VD4.n18 1.00018
R716 two_stage_opamp_dummy_magic_25_0.VD4.n26 two_stage_opamp_dummy_magic_25_0.VD4.n19 0.958833
R717 two_stage_opamp_dummy_magic_25_0.VD4.n21 two_stage_opamp_dummy_magic_25_0.VD4.n14 0.958833
R718 two_stage_opamp_dummy_magic_25_0.VD4.n8 two_stage_opamp_dummy_magic_25_0.VD4.n13 1.00018
R719 two_stage_opamp_dummy_magic_25_0.VD4.n7 two_stage_opamp_dummy_magic_25_0.VD4.n16 1.02002
R720 two_stage_opamp_dummy_magic_25_0.VD4.n27 two_stage_opamp_dummy_magic_25_0.VD4.n24 0.6255
R721 two_stage_opamp_dummy_magic_25_0.VD4.n24 two_stage_opamp_dummy_magic_25_0.VD4.n23 0.6255
R722 two_stage_opamp_dummy_magic_25_0.VD4.n23 two_stage_opamp_dummy_magic_25_0.VD4.n22 0.6255
R723 two_stage_opamp_dummy_magic_25_0.VD4.n0 two_stage_opamp_dummy_magic_25_0.VD4.n30 0.427973
R724 two_stage_opamp_dummy_magic_25_0.VD4.n30 two_stage_opamp_dummy_magic_25_0.VD4.n19 0.0587394
R725 two_stage_opamp_dummy_magic_25_0.VD4.n6 two_stage_opamp_dummy_magic_25_0.VD4.n19 0.0838727
R726 two_stage_opamp_dummy_magic_25_0.VD4.n8 two_stage_opamp_dummy_magic_25_0.VD4.n14 0.0838727
R727 two_stage_opamp_dummy_magic_25_0.VD4.n7 two_stage_opamp_dummy_magic_25_0.VD4.n14 0.0616865
R728 two_stage_opamp_dummy_magic_25_0.VD4.n32 two_stage_opamp_dummy_magic_25_0.VD4.n3 1.19908
R729 two_stage_opamp_dummy_magic_25_0.VD4.n3 two_stage_opamp_dummy_magic_25_0.VD4.n5 0.32698
R730 two_stage_opamp_dummy_magic_25_0.VD4.n5 two_stage_opamp_dummy_magic_25_0.VD4.n1 0.883997
R731 two_stage_opamp_dummy_magic_25_0.VD4.n1 two_stage_opamp_dummy_magic_25_0.VD4.n0 0.458833
R732 two_stage_opamp_dummy_magic_25_0.VD4.n4 two_stage_opamp_dummy_magic_25_0.VD4.n2 0.333833
R733 VDDA.n402 VDDA.t323 1231.74
R734 VDDA.n399 VDDA.t338 1231.74
R735 VDDA.n2298 VDDA.t305 1231.74
R736 VDDA.n2301 VDDA.t317 1231.74
R737 VDDA.n2357 VDDA.t248 826.801
R738 VDDA.n2389 VDDA.t350 826.801
R739 VDDA.n2363 VDDA.t344 826.801
R740 VDDA.n446 VDDA.t287 826.801
R741 VDDA.n1993 VDDA.t244 708.125
R742 VDDA.t244 VDDA.n1970 708.125
R743 VDDA.n2000 VDDA.t292 708.125
R744 VDDA.t292 VDDA.n1951 708.125
R745 VDDA.t272 VDDA.n2076 676.966
R746 VDDA.n2404 VDDA.t308 672.293
R747 VDDA.n365 VDDA.t259 672.293
R748 VDDA.n2266 VDDA.t281 672.293
R749 VDDA.n452 VDDA.t347 672.293
R750 VDDA.n378 VDDA.t268 661.375
R751 VDDA.n381 VDDA.t296 661.375
R752 VDDA.t333 VDDA.n1998 660.001
R753 VDDA.n1992 VDDA.t243 657.76
R754 VDDA.n1999 VDDA.t291 657.76
R755 VDDA.n2077 VDDA.t336 643.038
R756 VDDA.t312 VDDA.n2110 643.037
R757 VDDA.n2111 VDDA.t354 643.037
R758 VDDA.t303 VDDA.n2095 643.037
R759 VDDA.n2096 VDDA.t275 643.037
R760 VDDA.n2105 VDDA.t252 642.992
R761 VDDA.t342 VDDA.n2104 642.992
R762 VDDA.n2090 VDDA.t285 642.992
R763 VDDA.t246 VDDA.n2089 642.992
R764 VDDA.n1766 VDDA.t255 605.143
R765 VDDA.n1787 VDDA.t299 589.076
R766 VDDA.n2325 VDDA.t314 589.076
R767 VDDA.n2328 VDDA.t320 589.076
R768 VDDA.n433 VDDA.t329 589.076
R769 VDDA.n430 VDDA.t356 589.076
R770 VDDA.n2028 VDDA.n2026 587.407
R771 VDDA.n2032 VDDA.n2029 587.407
R772 VDDA.n2058 VDDA.n2057 587.407
R773 VDDA.n2053 VDDA.n2019 587.407
R774 VDDA.n2057 VDDA.n2056 585
R775 VDDA.n2055 VDDA.n2053 585
R776 VDDA.n2039 VDDA.n2028 585
R777 VDDA.n2036 VDDA.n2029 585
R778 VDDA.n2388 VDDA.n440 585
R779 VDDA.n2376 VDDA.n2375 585
R780 VDDA.n2373 VDDA.n2372 585
R781 VDDA.n2356 VDDA.n2355 585
R782 VDDA.t327 VDDA.n1991 540.818
R783 VDDA.n1777 VDDA.t301 464.281
R784 VDDA.t301 VDDA.n1393 464.281
R785 VDDA.n1772 VDDA.t258 464.281
R786 VDDA.t258 VDDA.n1771 464.281
R787 VDDA.n374 VDDA.t262 456.526
R788 VDDA.n371 VDDA.t277 456.526
R789 VDDA.n2098 VDDA.t341 441.2
R790 VDDA.n2106 VDDA.t251 441.2
R791 VDDA.n2087 VDDA.t245 441.2
R792 VDDA.n2091 VDDA.t284 441.2
R793 VDDA.n2078 VDDA.t335 413.084
R794 VDDA.n2075 VDDA.t271 413.084
R795 VDDA.n2107 VDDA.t311 409.067
R796 VDDA.n2112 VDDA.t353 409.067
R797 VDDA.t243 VDDA.t161 407.144
R798 VDDA.t161 VDDA.t15 407.144
R799 VDDA.t15 VDDA.t55 407.144
R800 VDDA.t55 VDDA.t133 407.144
R801 VDDA.t133 VDDA.t143 407.144
R802 VDDA.t143 VDDA.t186 407.144
R803 VDDA.t186 VDDA.t37 407.144
R804 VDDA.t37 VDDA.t141 407.144
R805 VDDA.t141 VDDA.t170 407.144
R806 VDDA.t170 VDDA.t122 407.144
R807 VDDA.t122 VDDA.t11 407.144
R808 VDDA.t11 VDDA.t163 407.144
R809 VDDA.t163 VDDA.t139 407.144
R810 VDDA.t139 VDDA.t365 407.144
R811 VDDA.t365 VDDA.t131 407.144
R812 VDDA.t131 VDDA.t57 407.144
R813 VDDA.t57 VDDA.t172 407.144
R814 VDDA.t172 VDDA.t9 407.144
R815 VDDA.t9 VDDA.t327 407.144
R816 VDDA.t291 VDDA.t198 407.144
R817 VDDA.t198 VDDA.t7 407.144
R818 VDDA.t7 VDDA.t192 407.144
R819 VDDA.t192 VDDA.t4 407.144
R820 VDDA.t4 VDDA.t188 407.144
R821 VDDA.t188 VDDA.t184 407.144
R822 VDDA.t184 VDDA.t190 407.144
R823 VDDA.t190 VDDA.t194 407.144
R824 VDDA.t194 VDDA.t64 407.144
R825 VDDA.t64 VDDA.t79 407.144
R826 VDDA.t79 VDDA.t69 407.144
R827 VDDA.t69 VDDA.t77 407.144
R828 VDDA.t77 VDDA.t368 407.144
R829 VDDA.t368 VDDA.t157 407.144
R830 VDDA.t157 VDDA.t0 407.144
R831 VDDA.t0 VDDA.t359 407.144
R832 VDDA.t359 VDDA.t361 407.144
R833 VDDA.t361 VDDA.t51 407.144
R834 VDDA.t51 VDDA.t333 407.144
R835 VDDA.n373 VDDA.t263 397.784
R836 VDDA.t278 VDDA.n372 397.784
R837 VDDA.n2092 VDDA.t302 390.322
R838 VDDA.n2097 VDDA.t274 390.322
R839 VDDA.t242 VDDA.n1993 379.582
R840 VDDA.t290 VDDA.n2000 379.582
R841 VDDA.n1990 VDDA.t326 379.277
R842 VDDA.t108 VDDA.t312 373.214
R843 VDDA.t407 VDDA.t108 373.214
R844 VDDA.t2 VDDA.t407 373.214
R845 VDDA.t178 VDDA.t2 373.214
R846 VDDA.t354 VDDA.t178 373.214
R847 VDDA.t159 VDDA.t342 373.214
R848 VDDA.t176 VDDA.t159 373.214
R849 VDDA.t155 VDDA.t176 373.214
R850 VDDA.t377 VDDA.t155 373.214
R851 VDDA.t394 VDDA.t377 373.214
R852 VDDA.t370 VDDA.t394 373.214
R853 VDDA.t43 VDDA.t370 373.214
R854 VDDA.t110 VDDA.t43 373.214
R855 VDDA.t252 VDDA.t110 373.214
R856 VDDA.t33 VDDA.t303 373.214
R857 VDDA.t174 VDDA.t33 373.214
R858 VDDA.t45 VDDA.t174 373.214
R859 VDDA.t39 VDDA.t45 373.214
R860 VDDA.t275 VDDA.t39 373.214
R861 VDDA.t182 VDDA.t246 373.214
R862 VDDA.t112 VDDA.t182 373.214
R863 VDDA.t285 VDDA.t112 373.214
R864 VDDA.t336 VDDA.t396 373.214
R865 VDDA.t396 VDDA.t84 373.214
R866 VDDA.t84 VDDA.t272 373.214
R867 VDDA.n2010 VDDA.t293 360.868
R868 VDDA.n2064 VDDA.t265 360.868
R869 VDDA.t326 VDDA.n1988 358.858
R870 VDDA.n1994 VDDA.t242 358.858
R871 VDDA.n1997 VDDA.t332 358.858
R872 VDDA.n2001 VDDA.t290 358.858
R873 VDDA.n2105 VDDA.t254 354.154
R874 VDDA.n2104 VDDA.t343 354.154
R875 VDDA.n2090 VDDA.t286 354.154
R876 VDDA.n2089 VDDA.t247 354.154
R877 VDDA.n1998 VDDA.t334 354.065
R878 VDDA.n2077 VDDA.t337 354.063
R879 VDDA.n1989 VDDA.t328 351.793
R880 VDDA.n2076 VDDA.t273 347.224
R881 VDDA.t315 VDDA.n2326 343.882
R882 VDDA.n2327 VDDA.t321 343.882
R883 VDDA.n432 VDDA.t330 343.882
R884 VDDA.t357 VDDA.n431 343.882
R885 VDDA.n2124 VDDA.n2094 342.197
R886 VDDA.n2125 VDDA.n2093 342.197
R887 VDDA.n2113 VDDA.n2109 341.769
R888 VDDA.n2114 VDDA.n2108 341.769
R889 VDDA.n1987 VDDA.n1986 338.714
R890 VDDA.n1985 VDDA.n1984 338.714
R891 VDDA.n1983 VDDA.n1982 338.714
R892 VDDA.n1981 VDDA.n1980 338.714
R893 VDDA.n1979 VDDA.n1978 338.714
R894 VDDA.n1977 VDDA.n1976 338.714
R895 VDDA.n1975 VDDA.n1974 338.714
R896 VDDA.n1973 VDDA.n1972 338.714
R897 VDDA.n1969 VDDA.n1968 338.714
R898 VDDA.n1967 VDDA.n1966 338.714
R899 VDDA.n1965 VDDA.n1964 338.714
R900 VDDA.n1963 VDDA.n1962 338.714
R901 VDDA.n1961 VDDA.n1960 338.714
R902 VDDA.n1959 VDDA.n1958 338.714
R903 VDDA.n1957 VDDA.n1956 338.714
R904 VDDA.n1955 VDDA.n1954 338.714
R905 VDDA.n1953 VDDA.n1952 338.714
R906 VDDA.n1950 VDDA.n1949 338.714
R907 VDDA.n2117 VDDA.n2103 336.341
R908 VDDA.n2118 VDDA.n2102 336.341
R909 VDDA.n2119 VDDA.n2101 336.341
R910 VDDA.n2120 VDDA.n2100 336.341
R911 VDDA.n2121 VDDA.n2099 336.341
R912 VDDA.n2128 VDDA.n2088 336.341
R913 VDDA.n2095 VDDA.t304 332.267
R914 VDDA.n2096 VDDA.t276 332.267
R915 VDDA.n2110 VDDA.t313 332.084
R916 VDDA.n2111 VDDA.t355 332.084
R917 VDDA.n2375 VDDA.n2367 291.053
R918 VDDA.n2375 VDDA.n2374 291.053
R919 VDDA.n2372 VDDA.n2365 291.053
R920 VDDA.n2372 VDDA.n2371 291.053
R921 VDDA.n2381 VDDA.n440 290.233
R922 VDDA.n2382 VDDA.n440 290.233
R923 VDDA.n2355 VDDA.n2345 290.233
R924 VDDA.n2355 VDDA.n2354 290.233
R925 VDDA.n1783 VDDA.t300 267.188
R926 VDDA.t256 VDDA.n1775 267.188
R927 VDDA.t263 VDDA.t25 259.091
R928 VDDA.t25 VDDA.t278 259.091
R929 VDDA.t414 VDDA.t294 251.471
R930 VDDA.t416 VDDA.t414 251.471
R931 VDDA.t17 VDDA.t416 251.471
R932 VDDA.t404 VDDA.t17 251.471
R933 VDDA.t126 VDDA.t404 251.471
R934 VDDA.t135 VDDA.t126 251.471
R935 VDDA.t137 VDDA.t135 251.471
R936 VDDA.t92 VDDA.t137 251.471
R937 VDDA.t389 VDDA.t92 251.471
R938 VDDA.t392 VDDA.t389 251.471
R939 VDDA.t19 VDDA.t392 251.471
R940 VDDA.t60 VDDA.t19 251.471
R941 VDDA.t88 VDDA.t60 251.471
R942 VDDA.t104 VDDA.t88 251.471
R943 VDDA.t418 VDDA.t104 251.471
R944 VDDA.t373 VDDA.t418 251.471
R945 VDDA.t266 VDDA.t373 251.471
R946 VDDA.n2382 VDDA.n2379 242.903
R947 VDDA.n2354 VDDA.n2353 242.903
R948 VDDA.n1774 VDDA.n1773 238.367
R949 VDDA.n1400 VDDA.n1396 238.367
R950 VDDA.n2060 VDDA.n2059 238.367
R951 VDDA.n1991 VDDA.n1990 238.367
R952 VDDA.n1991 VDDA.n1971 238.367
R953 VDDA.n2388 VDDA.n2387 238.367
R954 VDDA.n2377 VDDA.n2376 238.367
R955 VDDA.n2373 VDDA.n443 238.367
R956 VDDA.t294 VDDA.n2044 237.5
R957 VDDA.n2061 VDDA.t266 237.5
R958 VDDA.n2352 VDDA.t249 221.121
R959 VDDA.n2378 VDDA.t288 221.121
R960 VDDA.t345 VDDA.n2378 221.121
R961 VDDA.n2386 VDDA.t351 221.121
R962 VDDA.t300 VDDA.t31 217.708
R963 VDDA.t31 VDDA.t256 217.708
R964 VDDA.t165 VDDA.t315 217.708
R965 VDDA.t130 VDDA.t165 217.708
R966 VDDA.t23 VDDA.t130 217.708
R967 VDDA.t54 VDDA.t23 217.708
R968 VDDA.t106 VDDA.t54 217.708
R969 VDDA.t166 VDDA.t106 217.708
R970 VDDA.t53 VDDA.t166 217.708
R971 VDDA.t402 VDDA.t53 217.708
R972 VDDA.t403 VDDA.t402 217.708
R973 VDDA.t399 VDDA.t403 217.708
R974 VDDA.t321 VDDA.t399 217.708
R975 VDDA.t330 VDDA.t6 217.708
R976 VDDA.t6 VDDA.t412 217.708
R977 VDDA.t412 VDDA.t413 217.708
R978 VDDA.t413 VDDA.t383 217.708
R979 VDDA.t383 VDDA.t83 217.708
R980 VDDA.t83 VDDA.t21 217.708
R981 VDDA.t21 VDDA.t380 217.708
R982 VDDA.t380 VDDA.t14 217.708
R983 VDDA.t14 VDDA.t94 217.708
R984 VDDA.t94 VDDA.t384 217.708
R985 VDDA.t384 VDDA.t357 217.708
R986 VDDA.n439 VDDA.n438 216.677
R987 VDDA.n2360 VDDA.n2359 216.677
R988 VDDA.t269 VDDA.n379 213.131
R989 VDDA.n380 VDDA.t297 213.131
R990 VDDA.n2403 VDDA.t309 213.131
R991 VDDA.t260 VDDA.n2402 213.131
R992 VDDA.n2265 VDDA.t282 213.131
R993 VDDA.t348 VDDA.n2264 213.131
R994 VDDA.n1399 VDDA.n1397 185
R995 VDDA.n1770 VDDA.n1769 185
R996 VDDA.n1782 VDDA.n1781 185
R997 VDDA.n1783 VDDA.n1782 185
R998 VDDA.n1779 VDDA.n1776 185
R999 VDDA.n1778 VDDA.n1394 185
R1000 VDDA.n1785 VDDA.n1784 185
R1001 VDDA.n1784 VDDA.n1783 185
R1002 VDDA.n2049 VDDA.n2047 185
R1003 VDDA.n2056 VDDA.n2046 185
R1004 VDDA.n2061 VDDA.n2046 185
R1005 VDDA.n2055 VDDA.n2054 185
R1006 VDDA.n2052 VDDA.n2021 185
R1007 VDDA.n2063 VDDA.n2062 185
R1008 VDDA.n2062 VDDA.n2061 185
R1009 VDDA.n2043 VDDA.n2042 185
R1010 VDDA.n2044 VDDA.n2043 185
R1011 VDDA.n2040 VDDA.n2025 185
R1012 VDDA.n2039 VDDA.n2038 185
R1013 VDDA.n2037 VDDA.n2036 185
R1014 VDDA.n2031 VDDA.n2030 185
R1015 VDDA.n2033 VDDA.n2024 185
R1016 VDDA.n2044 VDDA.n2024 185
R1017 VDDA.n2366 VDDA.n445 185
R1018 VDDA.n2370 VDDA.n444 185
R1019 VDDA.n2378 VDDA.n444 185
R1020 VDDA.n2369 VDDA.n2368 185
R1021 VDDA.n442 VDDA.n441 185
R1022 VDDA.n2385 VDDA.n2384 185
R1023 VDDA.n2386 VDDA.n2385 185
R1024 VDDA.n2383 VDDA.n2380 185
R1025 VDDA.n2356 VDDA.n2343 185
R1026 VDDA.n2352 VDDA.n2343 185
R1027 VDDA.n2348 VDDA.n2344 185
R1028 VDDA.n2350 VDDA.n2349 185
R1029 VDDA.n2347 VDDA.n2346 185
R1030 VDDA.t249 VDDA.t68 180.173
R1031 VDDA.t68 VDDA.t66 180.173
R1032 VDDA.t66 VDDA.t41 180.173
R1033 VDDA.t41 VDDA.t364 180.173
R1034 VDDA.t364 VDDA.t288 180.173
R1035 VDDA.t363 VDDA.t345 180.173
R1036 VDDA.t397 VDDA.t363 180.173
R1037 VDDA.t180 VDDA.t397 180.173
R1038 VDDA.t24 VDDA.t180 180.173
R1039 VDDA.t351 VDDA.t24 180.173
R1040 VDDA.n373 VDDA.t264 168.139
R1041 VDDA.n372 VDDA.t280 168.139
R1042 VDDA.n370 VDDA.n369 150.643
R1043 VDDA.n1769 VDDA.n1397 150
R1044 VDDA.n1782 VDDA.n1776 150
R1045 VDDA.n1784 VDDA.n1394 150
R1046 VDDA.n2047 VDDA.n2046 150
R1047 VDDA.n2054 VDDA.n2046 150
R1048 VDDA.n2062 VDDA.n2021 150
R1049 VDDA.n2043 VDDA.n2025 150
R1050 VDDA.n2038 VDDA.n2037 150
R1051 VDDA.n2030 VDDA.n2024 150
R1052 VDDA.n2385 VDDA.n442 150
R1053 VDDA.n2385 VDDA.n2380 150
R1054 VDDA.n445 VDDA.n444 150
R1055 VDDA.n2368 VDDA.n444 150
R1056 VDDA.n2348 VDDA.n2343 150
R1057 VDDA.n2350 VDDA.n2347 150
R1058 VDDA.n1402 VDDA.n1401 149.112
R1059 VDDA.t208 VDDA.t269 146.155
R1060 VDDA.t297 VDDA.t208 146.155
R1061 VDDA.t309 VDDA.t220 146.155
R1062 VDDA.t220 VDDA.t232 146.155
R1063 VDDA.t232 VDDA.t200 146.155
R1064 VDDA.t200 VDDA.t236 146.155
R1065 VDDA.t236 VDDA.t202 146.155
R1066 VDDA.t202 VDDA.t206 146.155
R1067 VDDA.t206 VDDA.t222 146.155
R1068 VDDA.t222 VDDA.t234 146.155
R1069 VDDA.t234 VDDA.t228 146.155
R1070 VDDA.t228 VDDA.t240 146.155
R1071 VDDA.t240 VDDA.t260 146.155
R1072 VDDA.t282 VDDA.t212 146.155
R1073 VDDA.t212 VDDA.t216 146.155
R1074 VDDA.t216 VDDA.t226 146.155
R1075 VDDA.t226 VDDA.t238 146.155
R1076 VDDA.t238 VDDA.t204 146.155
R1077 VDDA.t204 VDDA.t210 146.155
R1078 VDDA.t210 VDDA.t214 146.155
R1079 VDDA.t214 VDDA.t218 146.155
R1080 VDDA.t218 VDDA.t230 146.155
R1081 VDDA.t230 VDDA.t224 146.155
R1082 VDDA.t224 VDDA.t348 146.155
R1083 VDDA.n2065 VDDA.n2018 141.712
R1084 VDDA.n2066 VDDA.n2017 141.712
R1085 VDDA.n2067 VDDA.n2016 141.712
R1086 VDDA.n2068 VDDA.n2015 141.712
R1087 VDDA.n2069 VDDA.n2014 141.712
R1088 VDDA.n2070 VDDA.n2013 141.712
R1089 VDDA.n2071 VDDA.n2012 141.712
R1090 VDDA.n2072 VDDA.n2011 141.712
R1091 VDDA.n2326 VDDA.t316 136.701
R1092 VDDA.n2327 VDDA.t322 136.701
R1093 VDDA.n432 VDDA.t331 136.701
R1094 VDDA.n431 VDDA.t358 136.701
R1095 VDDA.t295 VDDA.n2028 123.126
R1096 VDDA.n2029 VDDA.t295 123.126
R1097 VDDA.n2057 VDDA.t267 123.126
R1098 VDDA.n2053 VDDA.t267 123.126
R1099 VDDA.n401 VDDA.t324 122.829
R1100 VDDA.t339 VDDA.n400 122.829
R1101 VDDA.t306 VDDA.n2299 122.829
R1102 VDDA.n2300 VDDA.t318 122.829
R1103 VDDA.t324 VDDA.t410 81.6411
R1104 VDDA.t410 VDDA.t81 81.6411
R1105 VDDA.t81 VDDA.t75 81.6411
R1106 VDDA.t75 VDDA.t167 81.6411
R1107 VDDA.t167 VDDA.t35 81.6411
R1108 VDDA.t35 VDDA.t381 81.6411
R1109 VDDA.t381 VDDA.t115 81.6411
R1110 VDDA.t115 VDDA.t151 81.6411
R1111 VDDA.t151 VDDA.t386 81.6411
R1112 VDDA.t386 VDDA.t73 81.6411
R1113 VDDA.t73 VDDA.t339 81.6411
R1114 VDDA.t153 VDDA.t306 81.6411
R1115 VDDA.t149 VDDA.t153 81.6411
R1116 VDDA.t48 VDDA.t149 81.6411
R1117 VDDA.t97 VDDA.t48 81.6411
R1118 VDDA.t27 VDDA.t97 81.6411
R1119 VDDA.t71 VDDA.t27 81.6411
R1120 VDDA.t99 VDDA.t71 81.6411
R1121 VDDA.t375 VDDA.t99 81.6411
R1122 VDDA.t86 VDDA.t375 81.6411
R1123 VDDA.t400 VDDA.t86 81.6411
R1124 VDDA.t318 VDDA.t400 81.6411
R1125 VDDA.n379 VDDA.t270 76.2576
R1126 VDDA.n380 VDDA.t298 76.2576
R1127 VDDA.n2403 VDDA.t310 76.2576
R1128 VDDA.n2402 VDDA.t261 76.2576
R1129 VDDA.n2265 VDDA.t283 76.2576
R1130 VDDA.n2264 VDDA.t349 76.2576
R1131 VDDA.n2416 VDDA.n2415 71.3255
R1132 VDDA.n2414 VDDA.n2413 71.3255
R1133 VDDA.n2409 VDDA.n2408 71.3255
R1134 VDDA.n2407 VDDA.n2406 71.3255
R1135 VDDA.n2278 VDDA.n2277 71.3255
R1136 VDDA.n2276 VDDA.n2275 71.3255
R1137 VDDA.n2271 VDDA.n2270 71.3255
R1138 VDDA.n2269 VDDA.n2268 71.3255
R1139 VDDA.n377 VDDA.n376 68.4557
R1140 VDDA.n2411 VDDA.n2410 66.8255
R1141 VDDA.n2273 VDDA.n2272 66.8255
R1142 VDDA.n1775 VDDA.n1774 65.8183
R1143 VDDA.n1775 VDDA.n1396 65.8183
R1144 VDDA.n1783 VDDA.n1395 65.8183
R1145 VDDA.n2061 VDDA.n2060 65.8183
R1146 VDDA.n2061 VDDA.n2045 65.8183
R1147 VDDA.n2044 VDDA.n2022 65.8183
R1148 VDDA.n2044 VDDA.n2023 65.8183
R1149 VDDA.n2378 VDDA.n2377 65.8183
R1150 VDDA.n2378 VDDA.n443 65.8183
R1151 VDDA.n2387 VDDA.n2386 65.8183
R1152 VDDA.n2386 VDDA.n2379 65.8183
R1153 VDDA.n2352 VDDA.n2351 65.8183
R1154 VDDA.n2353 VDDA.n2352 65.8183
R1155 VDDA.n1940 VDDA.t422 58.8005
R1156 VDDA.n1939 VDDA.t424 58.8005
R1157 VDDA.n2389 VDDA.n2388 58.0576
R1158 VDDA.n2357 VDDA.n2356 58.0576
R1159 VDDA.n2364 VDDA.n2363 54.4005
R1160 VDDA.n2364 VDDA.n446 54.4005
R1161 VDDA.n1774 VDDA.n1397 53.3664
R1162 VDDA.n1769 VDDA.n1396 53.3664
R1163 VDDA.n1776 VDDA.n1395 53.3664
R1164 VDDA.n1395 VDDA.n1394 53.3664
R1165 VDDA.n2054 VDDA.n2045 53.3664
R1166 VDDA.n2060 VDDA.n2047 53.3664
R1167 VDDA.n2045 VDDA.n2021 53.3664
R1168 VDDA.n2025 VDDA.n2022 53.3664
R1169 VDDA.n2037 VDDA.n2023 53.3664
R1170 VDDA.n2038 VDDA.n2022 53.3664
R1171 VDDA.n2030 VDDA.n2023 53.3664
R1172 VDDA.n2380 VDDA.n2379 53.3664
R1173 VDDA.n2368 VDDA.n443 53.3664
R1174 VDDA.n2377 VDDA.n445 53.3664
R1175 VDDA.n2387 VDDA.n442 53.3664
R1176 VDDA.n2351 VDDA.n2348 53.3664
R1177 VDDA.n2353 VDDA.n2347 53.3664
R1178 VDDA.n2351 VDDA.n2350 53.3664
R1179 VDDA.n1939 VDDA.t421 49.1638
R1180 VDDA.n1941 VDDA.t423 48.5162
R1181 VDDA.n401 VDDA.t325 40.9789
R1182 VDDA.n400 VDDA.t340 40.9789
R1183 VDDA.n2299 VDDA.t307 40.9789
R1184 VDDA.n2300 VDDA.t319 40.9789
R1185 VDDA.n2109 VDDA.t3 39.4005
R1186 VDDA.n2109 VDDA.t179 39.4005
R1187 VDDA.n2108 VDDA.t109 39.4005
R1188 VDDA.n2108 VDDA.t408 39.4005
R1189 VDDA.n2103 VDDA.t111 39.4005
R1190 VDDA.n2103 VDDA.t253 39.4005
R1191 VDDA.n2102 VDDA.t371 39.4005
R1192 VDDA.n2102 VDDA.t44 39.4005
R1193 VDDA.n2101 VDDA.t378 39.4005
R1194 VDDA.n2101 VDDA.t395 39.4005
R1195 VDDA.n2100 VDDA.t177 39.4005
R1196 VDDA.n2100 VDDA.t156 39.4005
R1197 VDDA.t343 VDDA.n2099 39.4005
R1198 VDDA.n2099 VDDA.t160 39.4005
R1199 VDDA.n2094 VDDA.t46 39.4005
R1200 VDDA.n2094 VDDA.t40 39.4005
R1201 VDDA.n2093 VDDA.t34 39.4005
R1202 VDDA.n2093 VDDA.t175 39.4005
R1203 VDDA.n2088 VDDA.t183 39.4005
R1204 VDDA.n2088 VDDA.t113 39.4005
R1205 VDDA.n1986 VDDA.t173 39.4005
R1206 VDDA.n1986 VDDA.t10 39.4005
R1207 VDDA.n1984 VDDA.t132 39.4005
R1208 VDDA.n1984 VDDA.t58 39.4005
R1209 VDDA.n1982 VDDA.t140 39.4005
R1210 VDDA.n1982 VDDA.t366 39.4005
R1211 VDDA.n1980 VDDA.t12 39.4005
R1212 VDDA.n1980 VDDA.t164 39.4005
R1213 VDDA.n1978 VDDA.t171 39.4005
R1214 VDDA.n1978 VDDA.t123 39.4005
R1215 VDDA.n1976 VDDA.t38 39.4005
R1216 VDDA.n1976 VDDA.t142 39.4005
R1217 VDDA.n1974 VDDA.t144 39.4005
R1218 VDDA.n1974 VDDA.t187 39.4005
R1219 VDDA.n1972 VDDA.t56 39.4005
R1220 VDDA.n1972 VDDA.t134 39.4005
R1221 VDDA.n1968 VDDA.t162 39.4005
R1222 VDDA.n1968 VDDA.t16 39.4005
R1223 VDDA.n1966 VDDA.t362 39.4005
R1224 VDDA.n1966 VDDA.t52 39.4005
R1225 VDDA.n1964 VDDA.t1 39.4005
R1226 VDDA.n1964 VDDA.t360 39.4005
R1227 VDDA.n1962 VDDA.t369 39.4005
R1228 VDDA.n1962 VDDA.t158 39.4005
R1229 VDDA.n1960 VDDA.t70 39.4005
R1230 VDDA.n1960 VDDA.t78 39.4005
R1231 VDDA.n1958 VDDA.t65 39.4005
R1232 VDDA.n1958 VDDA.t80 39.4005
R1233 VDDA.n1956 VDDA.t191 39.4005
R1234 VDDA.n1956 VDDA.t195 39.4005
R1235 VDDA.n1954 VDDA.t189 39.4005
R1236 VDDA.n1954 VDDA.t185 39.4005
R1237 VDDA.n1952 VDDA.t193 39.4005
R1238 VDDA.n1952 VDDA.t5 39.4005
R1239 VDDA.n1949 VDDA.t199 39.4005
R1240 VDDA.n1949 VDDA.t8 39.4005
R1241 VDDA.n398 VDDA.n397 38.2279
R1242 VDDA.n396 VDDA.n395 38.2279
R1243 VDDA.n394 VDDA.n393 38.2279
R1244 VDDA.n392 VDDA.n391 38.2279
R1245 VDDA.n390 VDDA.n389 38.2279
R1246 VDDA.n2289 VDDA.n2288 38.2279
R1247 VDDA.n2291 VDDA.n2290 38.2279
R1248 VDDA.n2293 VDDA.n2292 38.2279
R1249 VDDA.n2295 VDDA.n2294 38.2279
R1250 VDDA.n2297 VDDA.n2296 38.2279
R1251 VDDA.n2112 VDDA.n2111 27.2462
R1252 VDDA.n2110 VDDA.n2107 27.2462
R1253 VDDA.n2097 VDDA.n2096 27.2462
R1254 VDDA.n2095 VDDA.n2092 27.2462
R1255 VDDA.n415 VDDA.n413 26.9096
R1256 VDDA.n2311 VDDA.n2309 26.8887
R1257 VDDA.n415 VDDA.n414 26.795
R1258 VDDA.n417 VDDA.n416 26.795
R1259 VDDA.n419 VDDA.n418 26.795
R1260 VDDA.n421 VDDA.n420 26.795
R1261 VDDA.n423 VDDA.n422 26.795
R1262 VDDA.n2319 VDDA.n2318 26.7741
R1263 VDDA.n2317 VDDA.n2316 26.7741
R1264 VDDA.n2315 VDDA.n2314 26.7741
R1265 VDDA.n2313 VDDA.n2312 26.7741
R1266 VDDA.n2311 VDDA.n2310 26.7741
R1267 VDDA.n2106 VDDA.n2105 24.9931
R1268 VDDA.n2104 VDDA.n2098 24.9931
R1269 VDDA.n2091 VDDA.n2090 24.9931
R1270 VDDA.n2089 VDDA.n2087 24.9931
R1271 VDDA.n1461 VDDA.t124 23.2175
R1272 VDDA.n2078 VDDA.n2077 22.9536
R1273 VDDA.n1998 VDDA.n1997 22.9536
R1274 VDDA.n2064 VDDA.n2063 22.8576
R1275 VDDA.n2033 VDDA.n2010 22.8576
R1276 VDDA.n369 VDDA.t26 21.8894
R1277 VDDA.n369 VDDA.t279 21.8894
R1278 VDDA.n1988 VDDA.n1971 20.7243
R1279 VDDA.n1994 VDDA.n1970 20.7243
R1280 VDDA.n2001 VDDA.n1951 20.7243
R1281 VDDA.n2076 VDDA.n2075 20.4312
R1282 VDDA.n1401 VDDA.t32 19.7005
R1283 VDDA.n1401 VDDA.t257 19.7005
R1284 VDDA.n2355 VDDA.t250 15.7605
R1285 VDDA.n440 VDDA.t352 15.7605
R1286 VDDA.n2372 VDDA.t346 15.7605
R1287 VDDA.n2375 VDDA.t289 15.7605
R1288 VDDA.n438 VDDA.t398 15.7605
R1289 VDDA.n438 VDDA.t181 15.7605
R1290 VDDA.n2359 VDDA.t67 15.7605
R1291 VDDA.n2359 VDDA.t42 15.7605
R1292 VDDA.n2018 VDDA.t419 13.1338
R1293 VDDA.n2018 VDDA.t374 13.1338
R1294 VDDA.n2017 VDDA.t89 13.1338
R1295 VDDA.n2017 VDDA.t105 13.1338
R1296 VDDA.n2016 VDDA.t20 13.1338
R1297 VDDA.n2016 VDDA.t61 13.1338
R1298 VDDA.n2015 VDDA.t390 13.1338
R1299 VDDA.n2015 VDDA.t393 13.1338
R1300 VDDA.n2014 VDDA.t138 13.1338
R1301 VDDA.n2014 VDDA.t93 13.1338
R1302 VDDA.n2013 VDDA.t127 13.1338
R1303 VDDA.n2013 VDDA.t136 13.1338
R1304 VDDA.n2012 VDDA.t18 13.1338
R1305 VDDA.n2012 VDDA.t405 13.1338
R1306 VDDA.n2011 VDDA.t415 13.1338
R1307 VDDA.n2011 VDDA.t417 13.1338
R1308 VDDA.n2075 VDDA.n2074 11.37
R1309 VDDA.n2079 VDDA.n2078 11.37
R1310 VDDA.t270 VDDA.n377 11.2576
R1311 VDDA.n377 VDDA.t209 11.2576
R1312 VDDA.n2415 VDDA.t229 11.2576
R1313 VDDA.n2415 VDDA.t241 11.2576
R1314 VDDA.n2413 VDDA.t223 11.2576
R1315 VDDA.n2413 VDDA.t235 11.2576
R1316 VDDA.n2410 VDDA.t203 11.2576
R1317 VDDA.n2410 VDDA.t207 11.2576
R1318 VDDA.n2408 VDDA.t201 11.2576
R1319 VDDA.n2408 VDDA.t237 11.2576
R1320 VDDA.n2406 VDDA.t221 11.2576
R1321 VDDA.n2406 VDDA.t233 11.2576
R1322 VDDA.n2277 VDDA.t231 11.2576
R1323 VDDA.n2277 VDDA.t225 11.2576
R1324 VDDA.n2275 VDDA.t215 11.2576
R1325 VDDA.n2275 VDDA.t219 11.2576
R1326 VDDA.n2272 VDDA.t205 11.2576
R1327 VDDA.n2272 VDDA.t211 11.2576
R1328 VDDA.n2270 VDDA.t227 11.2576
R1329 VDDA.n2270 VDDA.t239 11.2576
R1330 VDDA.n2268 VDDA.t213 11.2576
R1331 VDDA.n2268 VDDA.t217 11.2576
R1332 VDDA.n1988 VDDA.n1987 11.2346
R1333 VDDA.n1995 VDDA.n1994 11.1096
R1334 VDDA.n2002 VDDA.n2001 11.1096
R1335 VDDA.n1997 VDDA.n1996 11.1096
R1336 VDDA.n2065 VDDA.n2064 11.0575
R1337 VDDA.n2113 VDDA.n2112 10.9846
R1338 VDDA.n2115 VDDA.n2107 10.87
R1339 VDDA.n2122 VDDA.n2098 10.87
R1340 VDDA.n2126 VDDA.n2092 10.87
R1341 VDDA.n2129 VDDA.n2087 10.87
R1342 VDDA.n2127 VDDA.n2091 10.87
R1343 VDDA.n2123 VDDA.n2097 10.87
R1344 VDDA.n2116 VDDA.n2106 10.87
R1345 VDDA.n2073 VDDA.n2010 10.87
R1346 VDDA.n2358 VDDA.n2357 10.8696
R1347 VDDA.n2361 VDDA.n446 10.869
R1348 VDDA.n2363 VDDA.n2362 10.869
R1349 VDDA.n2390 VDDA.n2389 10.869
R1350 VDDA.n1773 VDDA.n1398 9.50883
R1351 VDDA.n1781 VDDA.n1780 9.50883
R1352 VDDA.n2042 VDDA.n2041 9.50883
R1353 VDDA.n2034 VDDA.n2033 9.50883
R1354 VDDA.n2059 VDDA.n2048 9.50883
R1355 VDDA.n2063 VDDA.n2020 9.50883
R1356 VDDA.n1770 VDDA.n1768 9.3005
R1357 VDDA.n1399 VDDA.n1398 9.3005
R1358 VDDA.n1767 VDDA.n1400 9.3005
R1359 VDDA.n1778 VDDA.n1392 9.3005
R1360 VDDA.n1780 VDDA.n1779 9.3005
R1361 VDDA.n1786 VDDA.n1785 9.3005
R1362 VDDA.n2052 VDDA.n2020 9.3005
R1363 VDDA.n2055 VDDA.n2051 9.3005
R1364 VDDA.n2056 VDDA.n2050 9.3005
R1365 VDDA.n2049 VDDA.n2048 9.3005
R1366 VDDA.n2034 VDDA.n2031 9.3005
R1367 VDDA.n2036 VDDA.n2035 9.3005
R1368 VDDA.n2039 VDDA.n2027 9.3005
R1369 VDDA.n2041 VDDA.n2040 9.3005
R1370 VDDA.n1770 VDDA.n1399 9.14336
R1371 VDDA.n1779 VDDA.n1778 9.14336
R1372 VDDA.n2056 VDDA.n2049 9.14336
R1373 VDDA.n2056 VDDA.n2055 9.14336
R1374 VDDA.n2055 VDDA.n2052 9.14336
R1375 VDDA.n2040 VDDA.n2039 9.14336
R1376 VDDA.n2039 VDDA.n2036 9.14336
R1377 VDDA.n2036 VDDA.n2031 9.14336
R1378 VDDA.n2388 VDDA.n441 9.14336
R1379 VDDA.n2384 VDDA.n2383 9.14336
R1380 VDDA.n2356 VDDA.n2344 9.14336
R1381 VDDA.n2349 VDDA.n2346 9.14336
R1382 VDDA.n2318 VDDA.t95 8.0005
R1383 VDDA.n2318 VDDA.t30 8.0005
R1384 VDDA.n2316 VDDA.t29 8.0005
R1385 VDDA.n2316 VDDA.t367 8.0005
R1386 VDDA.n2314 VDDA.t47 8.0005
R1387 VDDA.n2314 VDDA.t197 8.0005
R1388 VDDA.n2312 VDDA.t196 8.0005
R1389 VDDA.n2312 VDDA.t107 8.0005
R1390 VDDA.n2310 VDDA.t85 8.0005
R1391 VDDA.n2310 VDDA.t96 8.0005
R1392 VDDA.n2309 VDDA.t129 8.0005
R1393 VDDA.n2309 VDDA.t22 8.0005
R1394 VDDA.n413 VDDA.t120 8.0005
R1395 VDDA.n413 VDDA.t114 8.0005
R1396 VDDA.n414 VDDA.t385 8.0005
R1397 VDDA.n414 VDDA.t409 8.0005
R1398 VDDA.n416 VDDA.t13 8.0005
R1399 VDDA.n416 VDDA.t117 8.0005
R1400 VDDA.n418 VDDA.t119 8.0005
R1401 VDDA.n418 VDDA.t121 8.0005
R1402 VDDA.n420 VDDA.t169 8.0005
R1403 VDDA.n420 VDDA.t379 8.0005
R1404 VDDA.n422 VDDA.t50 8.0005
R1405 VDDA.n422 VDDA.t118 8.0005
R1406 VDDA.n397 VDDA.t387 6.56717
R1407 VDDA.n397 VDDA.t74 6.56717
R1408 VDDA.n395 VDDA.t116 6.56717
R1409 VDDA.n395 VDDA.t152 6.56717
R1410 VDDA.n393 VDDA.t36 6.56717
R1411 VDDA.n393 VDDA.t382 6.56717
R1412 VDDA.n391 VDDA.t76 6.56717
R1413 VDDA.n391 VDDA.t168 6.56717
R1414 VDDA.n389 VDDA.t411 6.56717
R1415 VDDA.n389 VDDA.t82 6.56717
R1416 VDDA.n2288 VDDA.t87 6.56717
R1417 VDDA.n2288 VDDA.t401 6.56717
R1418 VDDA.n2290 VDDA.t100 6.56717
R1419 VDDA.n2290 VDDA.t376 6.56717
R1420 VDDA.n2292 VDDA.t28 6.56717
R1421 VDDA.n2292 VDDA.t72 6.56717
R1422 VDDA.n2294 VDDA.t49 6.56717
R1423 VDDA.n2294 VDDA.t98 6.56717
R1424 VDDA.n2296 VDDA.t154 6.56717
R1425 VDDA.n2296 VDDA.t150 6.56717
R1426 VDDA.n1773 VDDA.n1772 5.33286
R1427 VDDA.n1771 VDDA.n1400 5.33286
R1428 VDDA.n1781 VDDA.n1777 5.33286
R1429 VDDA.n1785 VDDA.n1393 5.33286
R1430 VDDA.n2059 VDDA.n2058 5.33286
R1431 VDDA.n2063 VDDA.n2019 5.33286
R1432 VDDA.n2042 VDDA.n2026 5.33286
R1433 VDDA.n2033 VDDA.n2032 5.33286
R1434 VDDA.n2407 VDDA.n2405 5.1255
R1435 VDDA.n2417 VDDA.n2416 5.1255
R1436 VDDA.n2269 VDDA.n2267 5.1255
R1437 VDDA.n2279 VDDA.n2278 5.1255
R1438 VDDA.n1989 VDDA.n1971 4.54311
R1439 VDDA.n1990 VDDA.n1989 4.54311
R1440 VDDA.n2381 VDDA.n441 4.53698
R1441 VDDA.n2383 VDDA.n2382 4.53698
R1442 VDDA.n2384 VDDA.n2381 4.53698
R1443 VDDA.n2345 VDDA.n2344 4.53698
R1444 VDDA.n2354 VDDA.n2346 4.53698
R1445 VDDA.n2349 VDDA.n2345 4.53698
R1446 VDDA.n1790 VDDA.n1789 4.5005
R1447 VDDA.n1793 VDDA.n1792 4.5005
R1448 VDDA.n1794 VDDA.n1390 4.5005
R1449 VDDA.n1798 VDDA.n1795 4.5005
R1450 VDDA.n1799 VDDA.n1389 4.5005
R1451 VDDA.n1803 VDDA.n1802 4.5005
R1452 VDDA.n1804 VDDA.n1388 4.5005
R1453 VDDA.n1808 VDDA.n1805 4.5005
R1454 VDDA.n1809 VDDA.n1387 4.5005
R1455 VDDA.n1813 VDDA.n1812 4.5005
R1456 VDDA.n1814 VDDA.n1386 4.5005
R1457 VDDA.n1818 VDDA.n1815 4.5005
R1458 VDDA.n1819 VDDA.n1385 4.5005
R1459 VDDA.n1823 VDDA.n1822 4.5005
R1460 VDDA.n1824 VDDA.n1384 4.5005
R1461 VDDA.n1828 VDDA.n1825 4.5005
R1462 VDDA.n1829 VDDA.n1383 4.5005
R1463 VDDA.n1833 VDDA.n1832 4.5005
R1464 VDDA.n1834 VDDA.n1382 4.5005
R1465 VDDA.n1838 VDDA.n1835 4.5005
R1466 VDDA.n1839 VDDA.n1381 4.5005
R1467 VDDA.n1843 VDDA.n1842 4.5005
R1468 VDDA.n1844 VDDA.n1380 4.5005
R1469 VDDA.n1848 VDDA.n1845 4.5005
R1470 VDDA.n1849 VDDA.n1379 4.5005
R1471 VDDA.n1853 VDDA.n1852 4.5005
R1472 VDDA.n1854 VDDA.n1378 4.5005
R1473 VDDA.n1858 VDDA.n1855 4.5005
R1474 VDDA.n1859 VDDA.n1377 4.5005
R1475 VDDA.n1863 VDDA.n1862 4.5005
R1476 VDDA.n1864 VDDA.n1376 4.5005
R1477 VDDA.n1868 VDDA.n1865 4.5005
R1478 VDDA.n1869 VDDA.n1375 4.5005
R1479 VDDA.n1873 VDDA.n1872 4.5005
R1480 VDDA.n1874 VDDA.n1374 4.5005
R1481 VDDA.n1878 VDDA.n1875 4.5005
R1482 VDDA.n1879 VDDA.n1373 4.5005
R1483 VDDA.n1883 VDDA.n1882 4.5005
R1484 VDDA.n1884 VDDA.n1372 4.5005
R1485 VDDA.n1888 VDDA.n1885 4.5005
R1486 VDDA.n1889 VDDA.n1371 4.5005
R1487 VDDA.n1893 VDDA.n1892 4.5005
R1488 VDDA.n1894 VDDA.n1370 4.5005
R1489 VDDA.n1898 VDDA.n1895 4.5005
R1490 VDDA.n1899 VDDA.n1369 4.5005
R1491 VDDA.n1903 VDDA.n1902 4.5005
R1492 VDDA.n1462 VDDA.n1461 4.5005
R1493 VDDA.n1465 VDDA.n1464 4.5005
R1494 VDDA.n1466 VDDA.n1455 4.5005
R1495 VDDA.n1470 VDDA.n1467 4.5005
R1496 VDDA.n1471 VDDA.n1454 4.5005
R1497 VDDA.n1475 VDDA.n1474 4.5005
R1498 VDDA.n1476 VDDA.n1453 4.5005
R1499 VDDA.n1480 VDDA.n1477 4.5005
R1500 VDDA.n1481 VDDA.n1452 4.5005
R1501 VDDA.n1485 VDDA.n1484 4.5005
R1502 VDDA.n1486 VDDA.n1451 4.5005
R1503 VDDA.n1490 VDDA.n1487 4.5005
R1504 VDDA.n1491 VDDA.n1450 4.5005
R1505 VDDA.n1495 VDDA.n1494 4.5005
R1506 VDDA.n1496 VDDA.n1449 4.5005
R1507 VDDA.n1500 VDDA.n1497 4.5005
R1508 VDDA.n1501 VDDA.n1448 4.5005
R1509 VDDA.n1505 VDDA.n1504 4.5005
R1510 VDDA.n1506 VDDA.n1447 4.5005
R1511 VDDA.n1510 VDDA.n1507 4.5005
R1512 VDDA.n1511 VDDA.n1446 4.5005
R1513 VDDA.n1515 VDDA.n1514 4.5005
R1514 VDDA.n1516 VDDA.n1445 4.5005
R1515 VDDA.n1520 VDDA.n1517 4.5005
R1516 VDDA.n1521 VDDA.n1444 4.5005
R1517 VDDA.n1525 VDDA.n1524 4.5005
R1518 VDDA.n1526 VDDA.n1443 4.5005
R1519 VDDA.n1530 VDDA.n1527 4.5005
R1520 VDDA.n1531 VDDA.n1442 4.5005
R1521 VDDA.n1535 VDDA.n1534 4.5005
R1522 VDDA.n1536 VDDA.n1441 4.5005
R1523 VDDA.n1540 VDDA.n1537 4.5005
R1524 VDDA.n1541 VDDA.n1440 4.5005
R1525 VDDA.n1545 VDDA.n1544 4.5005
R1526 VDDA.n1546 VDDA.n1439 4.5005
R1527 VDDA.n1550 VDDA.n1547 4.5005
R1528 VDDA.n1551 VDDA.n1438 4.5005
R1529 VDDA.n1555 VDDA.n1554 4.5005
R1530 VDDA.n1556 VDDA.n1437 4.5005
R1531 VDDA.n1560 VDDA.n1557 4.5005
R1532 VDDA.n1561 VDDA.n1436 4.5005
R1533 VDDA.n1565 VDDA.n1564 4.5005
R1534 VDDA.n1566 VDDA.n1435 4.5005
R1535 VDDA.n1570 VDDA.n1567 4.5005
R1536 VDDA.n1571 VDDA.n1434 4.5005
R1537 VDDA.n1575 VDDA.n1574 4.5005
R1538 VDDA.n1945 VDDA.n1944 4.5005
R1539 VDDA.n2006 VDDA.n2005 4.5005
R1540 VDDA.n2083 VDDA.n2082 4.5005
R1541 VDDA.n2133 VDDA.n2132 4.5005
R1542 VDDA.n2137 VDDA.n2136 4.5005
R1543 VDDA.n2140 VDDA.n2139 4.5005
R1544 VDDA.n2141 VDDA.n1930 4.5005
R1545 VDDA.n2145 VDDA.n2142 4.5005
R1546 VDDA.n2146 VDDA.n1929 4.5005
R1547 VDDA.n2150 VDDA.n2149 4.5005
R1548 VDDA.n2151 VDDA.n1928 4.5005
R1549 VDDA.n2155 VDDA.n2152 4.5005
R1550 VDDA.n2156 VDDA.n1927 4.5005
R1551 VDDA.n2160 VDDA.n2159 4.5005
R1552 VDDA.n2161 VDDA.n1926 4.5005
R1553 VDDA.n2165 VDDA.n2162 4.5005
R1554 VDDA.n2166 VDDA.n1925 4.5005
R1555 VDDA.n2170 VDDA.n2169 4.5005
R1556 VDDA.n2171 VDDA.n1924 4.5005
R1557 VDDA.n2175 VDDA.n2172 4.5005
R1558 VDDA.n2176 VDDA.n1923 4.5005
R1559 VDDA.n2180 VDDA.n2179 4.5005
R1560 VDDA.n2181 VDDA.n1922 4.5005
R1561 VDDA.n2185 VDDA.n2182 4.5005
R1562 VDDA.n2186 VDDA.n1921 4.5005
R1563 VDDA.n2190 VDDA.n2189 4.5005
R1564 VDDA.n2191 VDDA.n1920 4.5005
R1565 VDDA.n2195 VDDA.n2192 4.5005
R1566 VDDA.n2196 VDDA.n1919 4.5005
R1567 VDDA.n2200 VDDA.n2199 4.5005
R1568 VDDA.n2201 VDDA.n1918 4.5005
R1569 VDDA.n2205 VDDA.n2202 4.5005
R1570 VDDA.n2206 VDDA.n1917 4.5005
R1571 VDDA.n2210 VDDA.n2209 4.5005
R1572 VDDA.n2211 VDDA.n1916 4.5005
R1573 VDDA.n2215 VDDA.n2212 4.5005
R1574 VDDA.n2216 VDDA.n1915 4.5005
R1575 VDDA.n2220 VDDA.n2219 4.5005
R1576 VDDA.n2221 VDDA.n1914 4.5005
R1577 VDDA.n2225 VDDA.n2222 4.5005
R1578 VDDA.n2226 VDDA.n1913 4.5005
R1579 VDDA.n2230 VDDA.n2229 4.5005
R1580 VDDA.n2231 VDDA.n1912 4.5005
R1581 VDDA.n2235 VDDA.n2232 4.5005
R1582 VDDA.n2236 VDDA.n1911 4.5005
R1583 VDDA.n2240 VDDA.n2239 4.5005
R1584 VDDA.n2241 VDDA.n1910 4.5005
R1585 VDDA.n2245 VDDA.n2242 4.5005
R1586 VDDA.n2246 VDDA.n1909 4.5005
R1587 VDDA.n2250 VDDA.n2249 4.5005
R1588 VDDA.n91 VDDA.n85 4.5005
R1589 VDDA.n93 VDDA.n92 4.5005
R1590 VDDA.n94 VDDA.n84 4.5005
R1591 VDDA.n98 VDDA.n97 4.5005
R1592 VDDA.n99 VDDA.n81 4.5005
R1593 VDDA.n101 VDDA.n100 4.5005
R1594 VDDA.n102 VDDA.n80 4.5005
R1595 VDDA.n106 VDDA.n105 4.5005
R1596 VDDA.n107 VDDA.n77 4.5005
R1597 VDDA.n109 VDDA.n108 4.5005
R1598 VDDA.n110 VDDA.n76 4.5005
R1599 VDDA.n114 VDDA.n113 4.5005
R1600 VDDA.n115 VDDA.n73 4.5005
R1601 VDDA.n117 VDDA.n116 4.5005
R1602 VDDA.n118 VDDA.n72 4.5005
R1603 VDDA.n122 VDDA.n121 4.5005
R1604 VDDA.n123 VDDA.n69 4.5005
R1605 VDDA.n125 VDDA.n124 4.5005
R1606 VDDA.n126 VDDA.n68 4.5005
R1607 VDDA.n130 VDDA.n129 4.5005
R1608 VDDA.n131 VDDA.n65 4.5005
R1609 VDDA.n133 VDDA.n132 4.5005
R1610 VDDA.n134 VDDA.n64 4.5005
R1611 VDDA.n138 VDDA.n137 4.5005
R1612 VDDA.n139 VDDA.n61 4.5005
R1613 VDDA.n141 VDDA.n140 4.5005
R1614 VDDA.n142 VDDA.n60 4.5005
R1615 VDDA.n146 VDDA.n145 4.5005
R1616 VDDA.n147 VDDA.n57 4.5005
R1617 VDDA.n149 VDDA.n148 4.5005
R1618 VDDA.n150 VDDA.n56 4.5005
R1619 VDDA.n154 VDDA.n153 4.5005
R1620 VDDA.n155 VDDA.n53 4.5005
R1621 VDDA.n157 VDDA.n156 4.5005
R1622 VDDA.n158 VDDA.n52 4.5005
R1623 VDDA.n162 VDDA.n161 4.5005
R1624 VDDA.n163 VDDA.n49 4.5005
R1625 VDDA.n165 VDDA.n164 4.5005
R1626 VDDA.n166 VDDA.n48 4.5005
R1627 VDDA.n170 VDDA.n169 4.5005
R1628 VDDA.n171 VDDA.n45 4.5005
R1629 VDDA.n173 VDDA.n172 4.5005
R1630 VDDA.n174 VDDA.n44 4.5005
R1631 VDDA.n178 VDDA.n177 4.5005
R1632 VDDA.n179 VDDA.n43 4.5005
R1633 VDDA.n2944 VDDA.n2943 4.5005
R1634 VDDA.n2813 VDDA.n2812 4.5005
R1635 VDDA.n2823 VDDA.n2822 4.5005
R1636 VDDA.n2824 VDDA.n2811 4.5005
R1637 VDDA.n2826 VDDA.n2825 4.5005
R1638 VDDA.n2809 VDDA.n2808 4.5005
R1639 VDDA.n2833 VDDA.n2832 4.5005
R1640 VDDA.n2834 VDDA.n2807 4.5005
R1641 VDDA.n2836 VDDA.n2835 4.5005
R1642 VDDA.n2805 VDDA.n2804 4.5005
R1643 VDDA.n2843 VDDA.n2842 4.5005
R1644 VDDA.n2844 VDDA.n2803 4.5005
R1645 VDDA.n2846 VDDA.n2845 4.5005
R1646 VDDA.n2801 VDDA.n2800 4.5005
R1647 VDDA.n2853 VDDA.n2852 4.5005
R1648 VDDA.n2854 VDDA.n2799 4.5005
R1649 VDDA.n2856 VDDA.n2855 4.5005
R1650 VDDA.n2797 VDDA.n2796 4.5005
R1651 VDDA.n2863 VDDA.n2862 4.5005
R1652 VDDA.n2864 VDDA.n2795 4.5005
R1653 VDDA.n2866 VDDA.n2865 4.5005
R1654 VDDA.n2793 VDDA.n2792 4.5005
R1655 VDDA.n2873 VDDA.n2872 4.5005
R1656 VDDA.n2874 VDDA.n2791 4.5005
R1657 VDDA.n2876 VDDA.n2875 4.5005
R1658 VDDA.n2789 VDDA.n2788 4.5005
R1659 VDDA.n2883 VDDA.n2882 4.5005
R1660 VDDA.n2884 VDDA.n2787 4.5005
R1661 VDDA.n2886 VDDA.n2885 4.5005
R1662 VDDA.n2785 VDDA.n2784 4.5005
R1663 VDDA.n2893 VDDA.n2892 4.5005
R1664 VDDA.n2894 VDDA.n2783 4.5005
R1665 VDDA.n2896 VDDA.n2895 4.5005
R1666 VDDA.n2781 VDDA.n2780 4.5005
R1667 VDDA.n2903 VDDA.n2902 4.5005
R1668 VDDA.n2904 VDDA.n2779 4.5005
R1669 VDDA.n2906 VDDA.n2905 4.5005
R1670 VDDA.n2777 VDDA.n2776 4.5005
R1671 VDDA.n2913 VDDA.n2912 4.5005
R1672 VDDA.n2914 VDDA.n2775 4.5005
R1673 VDDA.n2916 VDDA.n2915 4.5005
R1674 VDDA.n2773 VDDA.n2772 4.5005
R1675 VDDA.n2923 VDDA.n2922 4.5005
R1676 VDDA.n2924 VDDA.n2771 4.5005
R1677 VDDA.n2926 VDDA.n2925 4.5005
R1678 VDDA.n2769 VDDA.n2768 4.5005
R1679 VDDA.n2932 VDDA.n2931 4.5005
R1680 VDDA.n2668 VDDA.n2664 4.5005
R1681 VDDA.n2672 VDDA.n2671 4.5005
R1682 VDDA.n2673 VDDA.n2661 4.5005
R1683 VDDA.n2675 VDDA.n2674 4.5005
R1684 VDDA.n2676 VDDA.n2660 4.5005
R1685 VDDA.n2680 VDDA.n2679 4.5005
R1686 VDDA.n2681 VDDA.n2657 4.5005
R1687 VDDA.n2683 VDDA.n2682 4.5005
R1688 VDDA.n2684 VDDA.n2656 4.5005
R1689 VDDA.n2688 VDDA.n2687 4.5005
R1690 VDDA.n2689 VDDA.n2653 4.5005
R1691 VDDA.n2691 VDDA.n2690 4.5005
R1692 VDDA.n2692 VDDA.n2652 4.5005
R1693 VDDA.n2696 VDDA.n2695 4.5005
R1694 VDDA.n2697 VDDA.n2649 4.5005
R1695 VDDA.n2699 VDDA.n2698 4.5005
R1696 VDDA.n2700 VDDA.n2648 4.5005
R1697 VDDA.n2704 VDDA.n2703 4.5005
R1698 VDDA.n2705 VDDA.n2645 4.5005
R1699 VDDA.n2707 VDDA.n2706 4.5005
R1700 VDDA.n2708 VDDA.n2644 4.5005
R1701 VDDA.n2712 VDDA.n2711 4.5005
R1702 VDDA.n2713 VDDA.n2641 4.5005
R1703 VDDA.n2715 VDDA.n2714 4.5005
R1704 VDDA.n2716 VDDA.n2640 4.5005
R1705 VDDA.n2720 VDDA.n2719 4.5005
R1706 VDDA.n2721 VDDA.n2637 4.5005
R1707 VDDA.n2723 VDDA.n2722 4.5005
R1708 VDDA.n2724 VDDA.n2636 4.5005
R1709 VDDA.n2728 VDDA.n2727 4.5005
R1710 VDDA.n2729 VDDA.n2633 4.5005
R1711 VDDA.n2731 VDDA.n2730 4.5005
R1712 VDDA.n2732 VDDA.n2632 4.5005
R1713 VDDA.n2736 VDDA.n2735 4.5005
R1714 VDDA.n2737 VDDA.n2629 4.5005
R1715 VDDA.n2739 VDDA.n2738 4.5005
R1716 VDDA.n2740 VDDA.n2628 4.5005
R1717 VDDA.n2744 VDDA.n2743 4.5005
R1718 VDDA.n2745 VDDA.n2625 4.5005
R1719 VDDA.n2747 VDDA.n2746 4.5005
R1720 VDDA.n2748 VDDA.n2624 4.5005
R1721 VDDA.n2752 VDDA.n2751 4.5005
R1722 VDDA.n2753 VDDA.n2623 4.5005
R1723 VDDA.n2755 VDDA.n2754 4.5005
R1724 VDDA.n193 VDDA.n192 4.5005
R1725 VDDA.n2761 VDDA.n2760 4.5005
R1726 VDDA.n269 VDDA.n263 4.5005
R1727 VDDA.n271 VDDA.n270 4.5005
R1728 VDDA.n272 VDDA.n262 4.5005
R1729 VDDA.n276 VDDA.n275 4.5005
R1730 VDDA.n277 VDDA.n259 4.5005
R1731 VDDA.n279 VDDA.n278 4.5005
R1732 VDDA.n280 VDDA.n258 4.5005
R1733 VDDA.n284 VDDA.n283 4.5005
R1734 VDDA.n285 VDDA.n255 4.5005
R1735 VDDA.n287 VDDA.n286 4.5005
R1736 VDDA.n288 VDDA.n254 4.5005
R1737 VDDA.n292 VDDA.n291 4.5005
R1738 VDDA.n293 VDDA.n251 4.5005
R1739 VDDA.n295 VDDA.n294 4.5005
R1740 VDDA.n296 VDDA.n250 4.5005
R1741 VDDA.n300 VDDA.n299 4.5005
R1742 VDDA.n301 VDDA.n247 4.5005
R1743 VDDA.n303 VDDA.n302 4.5005
R1744 VDDA.n304 VDDA.n246 4.5005
R1745 VDDA.n308 VDDA.n307 4.5005
R1746 VDDA.n309 VDDA.n243 4.5005
R1747 VDDA.n311 VDDA.n310 4.5005
R1748 VDDA.n312 VDDA.n242 4.5005
R1749 VDDA.n316 VDDA.n315 4.5005
R1750 VDDA.n317 VDDA.n239 4.5005
R1751 VDDA.n319 VDDA.n318 4.5005
R1752 VDDA.n320 VDDA.n238 4.5005
R1753 VDDA.n324 VDDA.n323 4.5005
R1754 VDDA.n325 VDDA.n235 4.5005
R1755 VDDA.n327 VDDA.n326 4.5005
R1756 VDDA.n328 VDDA.n234 4.5005
R1757 VDDA.n332 VDDA.n331 4.5005
R1758 VDDA.n333 VDDA.n231 4.5005
R1759 VDDA.n335 VDDA.n334 4.5005
R1760 VDDA.n336 VDDA.n230 4.5005
R1761 VDDA.n340 VDDA.n339 4.5005
R1762 VDDA.n341 VDDA.n227 4.5005
R1763 VDDA.n343 VDDA.n342 4.5005
R1764 VDDA.n344 VDDA.n226 4.5005
R1765 VDDA.n348 VDDA.n347 4.5005
R1766 VDDA.n349 VDDA.n223 4.5005
R1767 VDDA.n351 VDDA.n350 4.5005
R1768 VDDA.n352 VDDA.n222 4.5005
R1769 VDDA.n356 VDDA.n355 4.5005
R1770 VDDA.n357 VDDA.n221 4.5005
R1771 VDDA.n2596 VDDA.n2595 4.5005
R1772 VDDA.n2465 VDDA.n2464 4.5005
R1773 VDDA.n2475 VDDA.n2474 4.5005
R1774 VDDA.n2476 VDDA.n2463 4.5005
R1775 VDDA.n2478 VDDA.n2477 4.5005
R1776 VDDA.n2461 VDDA.n2460 4.5005
R1777 VDDA.n2485 VDDA.n2484 4.5005
R1778 VDDA.n2486 VDDA.n2459 4.5005
R1779 VDDA.n2488 VDDA.n2487 4.5005
R1780 VDDA.n2457 VDDA.n2456 4.5005
R1781 VDDA.n2495 VDDA.n2494 4.5005
R1782 VDDA.n2496 VDDA.n2455 4.5005
R1783 VDDA.n2498 VDDA.n2497 4.5005
R1784 VDDA.n2453 VDDA.n2452 4.5005
R1785 VDDA.n2505 VDDA.n2504 4.5005
R1786 VDDA.n2506 VDDA.n2451 4.5005
R1787 VDDA.n2508 VDDA.n2507 4.5005
R1788 VDDA.n2449 VDDA.n2448 4.5005
R1789 VDDA.n2515 VDDA.n2514 4.5005
R1790 VDDA.n2516 VDDA.n2447 4.5005
R1791 VDDA.n2518 VDDA.n2517 4.5005
R1792 VDDA.n2445 VDDA.n2444 4.5005
R1793 VDDA.n2525 VDDA.n2524 4.5005
R1794 VDDA.n2526 VDDA.n2443 4.5005
R1795 VDDA.n2528 VDDA.n2527 4.5005
R1796 VDDA.n2441 VDDA.n2440 4.5005
R1797 VDDA.n2535 VDDA.n2534 4.5005
R1798 VDDA.n2536 VDDA.n2439 4.5005
R1799 VDDA.n2538 VDDA.n2537 4.5005
R1800 VDDA.n2437 VDDA.n2436 4.5005
R1801 VDDA.n2545 VDDA.n2544 4.5005
R1802 VDDA.n2546 VDDA.n2435 4.5005
R1803 VDDA.n2548 VDDA.n2547 4.5005
R1804 VDDA.n2433 VDDA.n2432 4.5005
R1805 VDDA.n2555 VDDA.n2554 4.5005
R1806 VDDA.n2556 VDDA.n2431 4.5005
R1807 VDDA.n2558 VDDA.n2557 4.5005
R1808 VDDA.n2429 VDDA.n2428 4.5005
R1809 VDDA.n2565 VDDA.n2564 4.5005
R1810 VDDA.n2566 VDDA.n2427 4.5005
R1811 VDDA.n2568 VDDA.n2567 4.5005
R1812 VDDA.n2425 VDDA.n2424 4.5005
R1813 VDDA.n2575 VDDA.n2574 4.5005
R1814 VDDA.n2576 VDDA.n2423 4.5005
R1815 VDDA.n2578 VDDA.n2577 4.5005
R1816 VDDA.n2421 VDDA.n2420 4.5005
R1817 VDDA.n2584 VDDA.n2583 4.5005
R1818 VDDA.n1228 VDDA.n1224 4.5005
R1819 VDDA.n1232 VDDA.n1231 4.5005
R1820 VDDA.n1233 VDDA.n1221 4.5005
R1821 VDDA.n1235 VDDA.n1234 4.5005
R1822 VDDA.n1236 VDDA.n1220 4.5005
R1823 VDDA.n1240 VDDA.n1239 4.5005
R1824 VDDA.n1241 VDDA.n1217 4.5005
R1825 VDDA.n1243 VDDA.n1242 4.5005
R1826 VDDA.n1244 VDDA.n1216 4.5005
R1827 VDDA.n1248 VDDA.n1247 4.5005
R1828 VDDA.n1249 VDDA.n1213 4.5005
R1829 VDDA.n1251 VDDA.n1250 4.5005
R1830 VDDA.n1252 VDDA.n1212 4.5005
R1831 VDDA.n1256 VDDA.n1255 4.5005
R1832 VDDA.n1257 VDDA.n1209 4.5005
R1833 VDDA.n1259 VDDA.n1258 4.5005
R1834 VDDA.n1260 VDDA.n1208 4.5005
R1835 VDDA.n1264 VDDA.n1263 4.5005
R1836 VDDA.n1265 VDDA.n1205 4.5005
R1837 VDDA.n1267 VDDA.n1266 4.5005
R1838 VDDA.n1268 VDDA.n1204 4.5005
R1839 VDDA.n1272 VDDA.n1271 4.5005
R1840 VDDA.n1273 VDDA.n1201 4.5005
R1841 VDDA.n1275 VDDA.n1274 4.5005
R1842 VDDA.n1276 VDDA.n1200 4.5005
R1843 VDDA.n1280 VDDA.n1279 4.5005
R1844 VDDA.n1281 VDDA.n1197 4.5005
R1845 VDDA.n1283 VDDA.n1282 4.5005
R1846 VDDA.n1284 VDDA.n1196 4.5005
R1847 VDDA.n1288 VDDA.n1287 4.5005
R1848 VDDA.n1289 VDDA.n1193 4.5005
R1849 VDDA.n1291 VDDA.n1290 4.5005
R1850 VDDA.n1292 VDDA.n1192 4.5005
R1851 VDDA.n1296 VDDA.n1295 4.5005
R1852 VDDA.n1297 VDDA.n1189 4.5005
R1853 VDDA.n1299 VDDA.n1298 4.5005
R1854 VDDA.n1300 VDDA.n1188 4.5005
R1855 VDDA.n1304 VDDA.n1303 4.5005
R1856 VDDA.n1305 VDDA.n1185 4.5005
R1857 VDDA.n1307 VDDA.n1306 4.5005
R1858 VDDA.n1308 VDDA.n1184 4.5005
R1859 VDDA.n1312 VDDA.n1311 4.5005
R1860 VDDA.n1313 VDDA.n1183 4.5005
R1861 VDDA.n1315 VDDA.n1314 4.5005
R1862 VDDA.n459 VDDA.n458 4.5005
R1863 VDDA.n2257 VDDA.n2256 4.5005
R1864 VDDA.n2412 VDDA.n2411 4.5005
R1865 VDDA.n407 VDDA.n406 4.5005
R1866 VDDA.n410 VDDA.n409 4.5005
R1867 VDDA.n2391 VDDA.n387 4.5005
R1868 VDDA.n2393 VDDA.n2392 4.5005
R1869 VDDA.n2392 VDDA.n2391 4.5005
R1870 VDDA.n2287 VDDA.n448 4.5005
R1871 VDDA.n2305 VDDA.n2304 4.5005
R1872 VDDA.n2308 VDDA.n2307 4.5005
R1873 VDDA.n2274 VDDA.n2273 4.5005
R1874 VDDA.n535 VDDA.n529 4.5005
R1875 VDDA.n537 VDDA.n536 4.5005
R1876 VDDA.n538 VDDA.n528 4.5005
R1877 VDDA.n542 VDDA.n541 4.5005
R1878 VDDA.n543 VDDA.n525 4.5005
R1879 VDDA.n545 VDDA.n544 4.5005
R1880 VDDA.n546 VDDA.n524 4.5005
R1881 VDDA.n550 VDDA.n549 4.5005
R1882 VDDA.n551 VDDA.n521 4.5005
R1883 VDDA.n553 VDDA.n552 4.5005
R1884 VDDA.n554 VDDA.n520 4.5005
R1885 VDDA.n558 VDDA.n557 4.5005
R1886 VDDA.n559 VDDA.n517 4.5005
R1887 VDDA.n561 VDDA.n560 4.5005
R1888 VDDA.n562 VDDA.n516 4.5005
R1889 VDDA.n566 VDDA.n565 4.5005
R1890 VDDA.n567 VDDA.n513 4.5005
R1891 VDDA.n569 VDDA.n568 4.5005
R1892 VDDA.n570 VDDA.n512 4.5005
R1893 VDDA.n574 VDDA.n573 4.5005
R1894 VDDA.n575 VDDA.n509 4.5005
R1895 VDDA.n577 VDDA.n576 4.5005
R1896 VDDA.n578 VDDA.n508 4.5005
R1897 VDDA.n582 VDDA.n581 4.5005
R1898 VDDA.n583 VDDA.n505 4.5005
R1899 VDDA.n585 VDDA.n584 4.5005
R1900 VDDA.n586 VDDA.n504 4.5005
R1901 VDDA.n590 VDDA.n589 4.5005
R1902 VDDA.n591 VDDA.n501 4.5005
R1903 VDDA.n593 VDDA.n592 4.5005
R1904 VDDA.n594 VDDA.n500 4.5005
R1905 VDDA.n598 VDDA.n597 4.5005
R1906 VDDA.n599 VDDA.n497 4.5005
R1907 VDDA.n601 VDDA.n600 4.5005
R1908 VDDA.n602 VDDA.n496 4.5005
R1909 VDDA.n606 VDDA.n605 4.5005
R1910 VDDA.n607 VDDA.n493 4.5005
R1911 VDDA.n609 VDDA.n608 4.5005
R1912 VDDA.n610 VDDA.n492 4.5005
R1913 VDDA.n614 VDDA.n613 4.5005
R1914 VDDA.n615 VDDA.n489 4.5005
R1915 VDDA.n617 VDDA.n616 4.5005
R1916 VDDA.n618 VDDA.n488 4.5005
R1917 VDDA.n622 VDDA.n621 4.5005
R1918 VDDA.n623 VDDA.n487 4.5005
R1919 VDDA.n1156 VDDA.n1155 4.5005
R1920 VDDA.n1025 VDDA.n1024 4.5005
R1921 VDDA.n1035 VDDA.n1034 4.5005
R1922 VDDA.n1036 VDDA.n1023 4.5005
R1923 VDDA.n1038 VDDA.n1037 4.5005
R1924 VDDA.n1021 VDDA.n1020 4.5005
R1925 VDDA.n1045 VDDA.n1044 4.5005
R1926 VDDA.n1046 VDDA.n1019 4.5005
R1927 VDDA.n1048 VDDA.n1047 4.5005
R1928 VDDA.n1017 VDDA.n1016 4.5005
R1929 VDDA.n1055 VDDA.n1054 4.5005
R1930 VDDA.n1056 VDDA.n1015 4.5005
R1931 VDDA.n1058 VDDA.n1057 4.5005
R1932 VDDA.n1013 VDDA.n1012 4.5005
R1933 VDDA.n1065 VDDA.n1064 4.5005
R1934 VDDA.n1066 VDDA.n1011 4.5005
R1935 VDDA.n1068 VDDA.n1067 4.5005
R1936 VDDA.n1009 VDDA.n1008 4.5005
R1937 VDDA.n1075 VDDA.n1074 4.5005
R1938 VDDA.n1076 VDDA.n1007 4.5005
R1939 VDDA.n1078 VDDA.n1077 4.5005
R1940 VDDA.n1005 VDDA.n1004 4.5005
R1941 VDDA.n1085 VDDA.n1084 4.5005
R1942 VDDA.n1086 VDDA.n1003 4.5005
R1943 VDDA.n1088 VDDA.n1087 4.5005
R1944 VDDA.n1001 VDDA.n1000 4.5005
R1945 VDDA.n1095 VDDA.n1094 4.5005
R1946 VDDA.n1096 VDDA.n999 4.5005
R1947 VDDA.n1098 VDDA.n1097 4.5005
R1948 VDDA.n997 VDDA.n996 4.5005
R1949 VDDA.n1105 VDDA.n1104 4.5005
R1950 VDDA.n1106 VDDA.n995 4.5005
R1951 VDDA.n1108 VDDA.n1107 4.5005
R1952 VDDA.n993 VDDA.n992 4.5005
R1953 VDDA.n1115 VDDA.n1114 4.5005
R1954 VDDA.n1116 VDDA.n991 4.5005
R1955 VDDA.n1118 VDDA.n1117 4.5005
R1956 VDDA.n989 VDDA.n988 4.5005
R1957 VDDA.n1125 VDDA.n1124 4.5005
R1958 VDDA.n1126 VDDA.n987 4.5005
R1959 VDDA.n1128 VDDA.n1127 4.5005
R1960 VDDA.n985 VDDA.n984 4.5005
R1961 VDDA.n1135 VDDA.n1134 4.5005
R1962 VDDA.n1136 VDDA.n983 4.5005
R1963 VDDA.n1138 VDDA.n1137 4.5005
R1964 VDDA.n981 VDDA.n980 4.5005
R1965 VDDA.n1144 VDDA.n1143 4.5005
R1966 VDDA.n880 VDDA.n876 4.5005
R1967 VDDA.n884 VDDA.n883 4.5005
R1968 VDDA.n885 VDDA.n873 4.5005
R1969 VDDA.n887 VDDA.n886 4.5005
R1970 VDDA.n888 VDDA.n872 4.5005
R1971 VDDA.n892 VDDA.n891 4.5005
R1972 VDDA.n893 VDDA.n869 4.5005
R1973 VDDA.n895 VDDA.n894 4.5005
R1974 VDDA.n896 VDDA.n868 4.5005
R1975 VDDA.n900 VDDA.n899 4.5005
R1976 VDDA.n901 VDDA.n865 4.5005
R1977 VDDA.n903 VDDA.n902 4.5005
R1978 VDDA.n904 VDDA.n864 4.5005
R1979 VDDA.n908 VDDA.n907 4.5005
R1980 VDDA.n909 VDDA.n861 4.5005
R1981 VDDA.n911 VDDA.n910 4.5005
R1982 VDDA.n912 VDDA.n860 4.5005
R1983 VDDA.n916 VDDA.n915 4.5005
R1984 VDDA.n917 VDDA.n857 4.5005
R1985 VDDA.n919 VDDA.n918 4.5005
R1986 VDDA.n920 VDDA.n856 4.5005
R1987 VDDA.n924 VDDA.n923 4.5005
R1988 VDDA.n925 VDDA.n853 4.5005
R1989 VDDA.n927 VDDA.n926 4.5005
R1990 VDDA.n928 VDDA.n852 4.5005
R1991 VDDA.n932 VDDA.n931 4.5005
R1992 VDDA.n933 VDDA.n849 4.5005
R1993 VDDA.n935 VDDA.n934 4.5005
R1994 VDDA.n936 VDDA.n848 4.5005
R1995 VDDA.n940 VDDA.n939 4.5005
R1996 VDDA.n941 VDDA.n845 4.5005
R1997 VDDA.n943 VDDA.n942 4.5005
R1998 VDDA.n944 VDDA.n844 4.5005
R1999 VDDA.n948 VDDA.n947 4.5005
R2000 VDDA.n949 VDDA.n841 4.5005
R2001 VDDA.n951 VDDA.n950 4.5005
R2002 VDDA.n952 VDDA.n840 4.5005
R2003 VDDA.n956 VDDA.n955 4.5005
R2004 VDDA.n957 VDDA.n837 4.5005
R2005 VDDA.n959 VDDA.n958 4.5005
R2006 VDDA.n960 VDDA.n836 4.5005
R2007 VDDA.n964 VDDA.n963 4.5005
R2008 VDDA.n965 VDDA.n835 4.5005
R2009 VDDA.n967 VDDA.n966 4.5005
R2010 VDDA.n636 VDDA.n635 4.5005
R2011 VDDA.n973 VDDA.n972 4.5005
R2012 VDDA.n976 VDDA.n634 4.5005
R2013 VDDA.n978 VDDA.n977 4.5005
R2014 VDDA.n977 VDDA.n976 4.5005
R2015 VDDA.n1147 VDDA.n979 4.5005
R2016 VDDA.n1149 VDDA.n1148 4.5005
R2017 VDDA.n1148 VDDA.n1147 4.5005
R2018 VDDA.n1152 VDDA.n1151 4.5005
R2019 VDDA.n1150 VDDA.n456 4.5005
R2020 VDDA.n1151 VDDA.n1150 4.5005
R2021 VDDA.n2285 VDDA.n2281 4.5005
R2022 VDDA.n2286 VDDA.n450 4.5005
R2023 VDDA.n2286 VDDA.n2285 4.5005
R2024 VDDA.n2400 VDDA.n2399 4.5005
R2025 VDDA.n2399 VDDA.n2398 4.5005
R2026 VDDA.n2398 VDDA.n385 4.5005
R2027 VDDA.n2260 VDDA.n457 4.5005
R2028 VDDA.n2262 VDDA.n2261 4.5005
R2029 VDDA.n2261 VDDA.n2260 4.5005
R2030 VDDA.n2587 VDDA.n2419 4.5005
R2031 VDDA.n2589 VDDA.n2588 4.5005
R2032 VDDA.n2588 VDDA.n2587 4.5005
R2033 VDDA.n2592 VDDA.n2591 4.5005
R2034 VDDA.n2590 VDDA.n190 4.5005
R2035 VDDA.n2591 VDDA.n2590 4.5005
R2036 VDDA.n2764 VDDA.n191 4.5005
R2037 VDDA.n2766 VDDA.n2765 4.5005
R2038 VDDA.n2765 VDDA.n2764 4.5005
R2039 VDDA.n2935 VDDA.n2767 4.5005
R2040 VDDA.n2937 VDDA.n2936 4.5005
R2041 VDDA.n2936 VDDA.n2935 4.5005
R2042 VDDA.n2938 VDDA.n181 4.5005
R2043 VDDA.n2940 VDDA.n2939 4.5005
R2044 VDDA.n2939 VDDA.n2938 4.5005
R2045 VDDA.n804 VDDA.n801 4.5005
R2046 VDDA.n689 VDDA.n685 4.5005
R2047 VDDA.n693 VDDA.n690 4.5005
R2048 VDDA.n694 VDDA.n684 4.5005
R2049 VDDA.n698 VDDA.n697 4.5005
R2050 VDDA.n699 VDDA.n683 4.5005
R2051 VDDA.n703 VDDA.n700 4.5005
R2052 VDDA.n704 VDDA.n682 4.5005
R2053 VDDA.n708 VDDA.n707 4.5005
R2054 VDDA.n709 VDDA.n681 4.5005
R2055 VDDA.n713 VDDA.n710 4.5005
R2056 VDDA.n714 VDDA.n680 4.5005
R2057 VDDA.n718 VDDA.n717 4.5005
R2058 VDDA.n719 VDDA.n679 4.5005
R2059 VDDA.n723 VDDA.n720 4.5005
R2060 VDDA.n724 VDDA.n678 4.5005
R2061 VDDA.n728 VDDA.n727 4.5005
R2062 VDDA.n729 VDDA.n677 4.5005
R2063 VDDA.n733 VDDA.n730 4.5005
R2064 VDDA.n734 VDDA.n676 4.5005
R2065 VDDA.n738 VDDA.n737 4.5005
R2066 VDDA.n739 VDDA.n675 4.5005
R2067 VDDA.n743 VDDA.n740 4.5005
R2068 VDDA.n744 VDDA.n674 4.5005
R2069 VDDA.n748 VDDA.n747 4.5005
R2070 VDDA.n749 VDDA.n673 4.5005
R2071 VDDA.n753 VDDA.n750 4.5005
R2072 VDDA.n754 VDDA.n672 4.5005
R2073 VDDA.n758 VDDA.n757 4.5005
R2074 VDDA.n759 VDDA.n671 4.5005
R2075 VDDA.n763 VDDA.n760 4.5005
R2076 VDDA.n764 VDDA.n670 4.5005
R2077 VDDA.n768 VDDA.n767 4.5005
R2078 VDDA.n769 VDDA.n669 4.5005
R2079 VDDA.n773 VDDA.n770 4.5005
R2080 VDDA.n774 VDDA.n668 4.5005
R2081 VDDA.n778 VDDA.n777 4.5005
R2082 VDDA.n779 VDDA.n667 4.5005
R2083 VDDA.n783 VDDA.n780 4.5005
R2084 VDDA.n784 VDDA.n666 4.5005
R2085 VDDA.n788 VDDA.n787 4.5005
R2086 VDDA.n789 VDDA.n665 4.5005
R2087 VDDA.n793 VDDA.n790 4.5005
R2088 VDDA.n794 VDDA.n664 4.5005
R2089 VDDA.n798 VDDA.n797 4.5005
R2090 VDDA.n799 VDDA.n663 4.5005
R2091 VDDA.n808 VDDA.n807 4.5005
R2092 VDDA.n1992 VDDA.n1970 4.48641
R2093 VDDA.n1993 VDDA.n1992 4.48641
R2094 VDDA.n1999 VDDA.n1951 4.48641
R2095 VDDA.n2000 VDDA.n1999 4.48641
R2096 VDDA.n1772 VDDA.n1399 3.75335
R2097 VDDA.n1771 VDDA.n1770 3.75335
R2098 VDDA.n1779 VDDA.n1777 3.75335
R2099 VDDA.n1778 VDDA.n1393 3.75335
R2100 VDDA.n2058 VDDA.n2049 3.75335
R2101 VDDA.n2052 VDDA.n2019 3.75335
R2102 VDDA.n2040 VDDA.n2026 3.75335
R2103 VDDA.n2032 VDDA.n2031 3.75335
R2104 VDDA.n1905 VDDA.n1904 3.4877
R2105 VDDA.n1577 VDDA.n1576 3.47821
R2106 VDDA.n2252 VDDA.n2251 3.47821
R2107 VDDA.n90 VDDA.n18 3.47821
R2108 VDDA.n2815 VDDA.n2814 3.47821
R2109 VDDA.n2665 VDDA.n2599 3.47821
R2110 VDDA.n268 VDDA.n196 3.47821
R2111 VDDA.n2467 VDDA.n2466 3.47821
R2112 VDDA.n1225 VDDA.n1159 3.47821
R2113 VDDA.n534 VDDA.n462 3.47821
R2114 VDDA.n1027 VDDA.n1026 3.47821
R2115 VDDA.n877 VDDA.n811 3.47821
R2116 VDDA.n688 VDDA.n638 3.47821
R2117 VDDA.n1368 VDDA.n1367 3.4105
R2118 VDDA.n1902 VDDA.n1901 3.4105
R2119 VDDA.n1900 VDDA.n1899 3.4105
R2120 VDDA.n1898 VDDA.n1897 3.4105
R2121 VDDA.n1896 VDDA.n1370 3.4105
R2122 VDDA.n1892 VDDA.n1891 3.4105
R2123 VDDA.n1890 VDDA.n1889 3.4105
R2124 VDDA.n1888 VDDA.n1887 3.4105
R2125 VDDA.n1886 VDDA.n1372 3.4105
R2126 VDDA.n1882 VDDA.n1881 3.4105
R2127 VDDA.n1880 VDDA.n1879 3.4105
R2128 VDDA.n1878 VDDA.n1877 3.4105
R2129 VDDA.n1876 VDDA.n1374 3.4105
R2130 VDDA.n1872 VDDA.n1871 3.4105
R2131 VDDA.n1870 VDDA.n1869 3.4105
R2132 VDDA.n1868 VDDA.n1867 3.4105
R2133 VDDA.n1866 VDDA.n1376 3.4105
R2134 VDDA.n1862 VDDA.n1861 3.4105
R2135 VDDA.n1860 VDDA.n1859 3.4105
R2136 VDDA.n1858 VDDA.n1857 3.4105
R2137 VDDA.n1856 VDDA.n1378 3.4105
R2138 VDDA.n1852 VDDA.n1851 3.4105
R2139 VDDA.n1850 VDDA.n1849 3.4105
R2140 VDDA.n1848 VDDA.n1847 3.4105
R2141 VDDA.n1846 VDDA.n1380 3.4105
R2142 VDDA.n1842 VDDA.n1841 3.4105
R2143 VDDA.n1840 VDDA.n1839 3.4105
R2144 VDDA.n1838 VDDA.n1837 3.4105
R2145 VDDA.n1836 VDDA.n1382 3.4105
R2146 VDDA.n1832 VDDA.n1831 3.4105
R2147 VDDA.n1830 VDDA.n1829 3.4105
R2148 VDDA.n1828 VDDA.n1827 3.4105
R2149 VDDA.n1826 VDDA.n1384 3.4105
R2150 VDDA.n1822 VDDA.n1821 3.4105
R2151 VDDA.n1820 VDDA.n1819 3.4105
R2152 VDDA.n1818 VDDA.n1817 3.4105
R2153 VDDA.n1816 VDDA.n1386 3.4105
R2154 VDDA.n1812 VDDA.n1811 3.4105
R2155 VDDA.n1810 VDDA.n1809 3.4105
R2156 VDDA.n1808 VDDA.n1807 3.4105
R2157 VDDA.n1806 VDDA.n1388 3.4105
R2158 VDDA.n1802 VDDA.n1801 3.4105
R2159 VDDA.n1800 VDDA.n1799 3.4105
R2160 VDDA.n1798 VDDA.n1797 3.4105
R2161 VDDA.n1796 VDDA.n1390 3.4105
R2162 VDDA.n1792 VDDA.n1791 3.4105
R2163 VDDA.n1790 VDDA.n1342 3.4105
R2164 VDDA.n1433 VDDA.n1432 3.4105
R2165 VDDA.n1574 VDDA.n1573 3.4105
R2166 VDDA.n1572 VDDA.n1571 3.4105
R2167 VDDA.n1570 VDDA.n1569 3.4105
R2168 VDDA.n1568 VDDA.n1435 3.4105
R2169 VDDA.n1564 VDDA.n1563 3.4105
R2170 VDDA.n1562 VDDA.n1561 3.4105
R2171 VDDA.n1560 VDDA.n1559 3.4105
R2172 VDDA.n1558 VDDA.n1437 3.4105
R2173 VDDA.n1554 VDDA.n1553 3.4105
R2174 VDDA.n1552 VDDA.n1551 3.4105
R2175 VDDA.n1550 VDDA.n1549 3.4105
R2176 VDDA.n1548 VDDA.n1439 3.4105
R2177 VDDA.n1544 VDDA.n1543 3.4105
R2178 VDDA.n1542 VDDA.n1541 3.4105
R2179 VDDA.n1540 VDDA.n1539 3.4105
R2180 VDDA.n1538 VDDA.n1441 3.4105
R2181 VDDA.n1534 VDDA.n1533 3.4105
R2182 VDDA.n1532 VDDA.n1531 3.4105
R2183 VDDA.n1530 VDDA.n1529 3.4105
R2184 VDDA.n1528 VDDA.n1443 3.4105
R2185 VDDA.n1524 VDDA.n1523 3.4105
R2186 VDDA.n1522 VDDA.n1521 3.4105
R2187 VDDA.n1520 VDDA.n1519 3.4105
R2188 VDDA.n1518 VDDA.n1445 3.4105
R2189 VDDA.n1514 VDDA.n1513 3.4105
R2190 VDDA.n1512 VDDA.n1511 3.4105
R2191 VDDA.n1510 VDDA.n1509 3.4105
R2192 VDDA.n1508 VDDA.n1447 3.4105
R2193 VDDA.n1504 VDDA.n1503 3.4105
R2194 VDDA.n1502 VDDA.n1501 3.4105
R2195 VDDA.n1500 VDDA.n1499 3.4105
R2196 VDDA.n1498 VDDA.n1449 3.4105
R2197 VDDA.n1494 VDDA.n1493 3.4105
R2198 VDDA.n1492 VDDA.n1491 3.4105
R2199 VDDA.n1490 VDDA.n1489 3.4105
R2200 VDDA.n1488 VDDA.n1451 3.4105
R2201 VDDA.n1484 VDDA.n1483 3.4105
R2202 VDDA.n1482 VDDA.n1481 3.4105
R2203 VDDA.n1480 VDDA.n1479 3.4105
R2204 VDDA.n1478 VDDA.n1453 3.4105
R2205 VDDA.n1474 VDDA.n1473 3.4105
R2206 VDDA.n1472 VDDA.n1471 3.4105
R2207 VDDA.n1470 VDDA.n1469 3.4105
R2208 VDDA.n1468 VDDA.n1455 3.4105
R2209 VDDA.n1464 VDDA.n1463 3.4105
R2210 VDDA.n1462 VDDA.n1408 3.4105
R2211 VDDA.n1908 VDDA.n1907 3.4105
R2212 VDDA.n2249 VDDA.n2248 3.4105
R2213 VDDA.n2247 VDDA.n2246 3.4105
R2214 VDDA.n2245 VDDA.n2244 3.4105
R2215 VDDA.n2243 VDDA.n1910 3.4105
R2216 VDDA.n2239 VDDA.n2238 3.4105
R2217 VDDA.n2237 VDDA.n2236 3.4105
R2218 VDDA.n2235 VDDA.n2234 3.4105
R2219 VDDA.n2233 VDDA.n1912 3.4105
R2220 VDDA.n2229 VDDA.n2228 3.4105
R2221 VDDA.n2227 VDDA.n2226 3.4105
R2222 VDDA.n2225 VDDA.n2224 3.4105
R2223 VDDA.n2223 VDDA.n1914 3.4105
R2224 VDDA.n2219 VDDA.n2218 3.4105
R2225 VDDA.n2217 VDDA.n2216 3.4105
R2226 VDDA.n2215 VDDA.n2214 3.4105
R2227 VDDA.n2213 VDDA.n1916 3.4105
R2228 VDDA.n2209 VDDA.n2208 3.4105
R2229 VDDA.n2207 VDDA.n2206 3.4105
R2230 VDDA.n2205 VDDA.n2204 3.4105
R2231 VDDA.n2203 VDDA.n1918 3.4105
R2232 VDDA.n2199 VDDA.n2198 3.4105
R2233 VDDA.n2197 VDDA.n2196 3.4105
R2234 VDDA.n2195 VDDA.n2194 3.4105
R2235 VDDA.n2193 VDDA.n1920 3.4105
R2236 VDDA.n2189 VDDA.n2188 3.4105
R2237 VDDA.n2187 VDDA.n2186 3.4105
R2238 VDDA.n2185 VDDA.n2184 3.4105
R2239 VDDA.n2183 VDDA.n1922 3.4105
R2240 VDDA.n2179 VDDA.n2178 3.4105
R2241 VDDA.n2177 VDDA.n2176 3.4105
R2242 VDDA.n2175 VDDA.n2174 3.4105
R2243 VDDA.n2173 VDDA.n1924 3.4105
R2244 VDDA.n2169 VDDA.n2168 3.4105
R2245 VDDA.n2167 VDDA.n2166 3.4105
R2246 VDDA.n2165 VDDA.n2164 3.4105
R2247 VDDA.n2163 VDDA.n1926 3.4105
R2248 VDDA.n2159 VDDA.n2158 3.4105
R2249 VDDA.n2157 VDDA.n2156 3.4105
R2250 VDDA.n2155 VDDA.n2154 3.4105
R2251 VDDA.n2153 VDDA.n1928 3.4105
R2252 VDDA.n2149 VDDA.n2148 3.4105
R2253 VDDA.n2147 VDDA.n2146 3.4105
R2254 VDDA.n2145 VDDA.n2144 3.4105
R2255 VDDA.n2143 VDDA.n1930 3.4105
R2256 VDDA.n2139 VDDA.n2138 3.4105
R2257 VDDA.n2137 VDDA.n1318 3.4105
R2258 VDDA.n43 VDDA.n42 3.4105
R2259 VDDA.n177 VDDA.n176 3.4105
R2260 VDDA.n175 VDDA.n174 3.4105
R2261 VDDA.n173 VDDA.n47 3.4105
R2262 VDDA.n46 VDDA.n45 3.4105
R2263 VDDA.n169 VDDA.n168 3.4105
R2264 VDDA.n167 VDDA.n166 3.4105
R2265 VDDA.n165 VDDA.n51 3.4105
R2266 VDDA.n50 VDDA.n49 3.4105
R2267 VDDA.n161 VDDA.n160 3.4105
R2268 VDDA.n159 VDDA.n158 3.4105
R2269 VDDA.n157 VDDA.n55 3.4105
R2270 VDDA.n54 VDDA.n53 3.4105
R2271 VDDA.n153 VDDA.n152 3.4105
R2272 VDDA.n151 VDDA.n150 3.4105
R2273 VDDA.n149 VDDA.n59 3.4105
R2274 VDDA.n58 VDDA.n57 3.4105
R2275 VDDA.n145 VDDA.n144 3.4105
R2276 VDDA.n143 VDDA.n142 3.4105
R2277 VDDA.n141 VDDA.n63 3.4105
R2278 VDDA.n62 VDDA.n61 3.4105
R2279 VDDA.n137 VDDA.n136 3.4105
R2280 VDDA.n135 VDDA.n134 3.4105
R2281 VDDA.n133 VDDA.n67 3.4105
R2282 VDDA.n66 VDDA.n65 3.4105
R2283 VDDA.n129 VDDA.n128 3.4105
R2284 VDDA.n127 VDDA.n126 3.4105
R2285 VDDA.n125 VDDA.n71 3.4105
R2286 VDDA.n70 VDDA.n69 3.4105
R2287 VDDA.n121 VDDA.n120 3.4105
R2288 VDDA.n119 VDDA.n118 3.4105
R2289 VDDA.n117 VDDA.n75 3.4105
R2290 VDDA.n74 VDDA.n73 3.4105
R2291 VDDA.n113 VDDA.n112 3.4105
R2292 VDDA.n111 VDDA.n110 3.4105
R2293 VDDA.n109 VDDA.n79 3.4105
R2294 VDDA.n78 VDDA.n77 3.4105
R2295 VDDA.n105 VDDA.n104 3.4105
R2296 VDDA.n103 VDDA.n102 3.4105
R2297 VDDA.n101 VDDA.n83 3.4105
R2298 VDDA.n82 VDDA.n81 3.4105
R2299 VDDA.n97 VDDA.n96 3.4105
R2300 VDDA.n95 VDDA.n94 3.4105
R2301 VDDA.n93 VDDA.n87 3.4105
R2302 VDDA.n86 VDDA.n85 3.4105
R2303 VDDA.n89 VDDA.n88 3.4105
R2304 VDDA.n2945 VDDA.n2944 3.4105
R2305 VDDA.n2929 VDDA.n2769 3.4105
R2306 VDDA.n2927 VDDA.n2926 3.4105
R2307 VDDA.n2771 VDDA.n2770 3.4105
R2308 VDDA.n2922 VDDA.n2921 3.4105
R2309 VDDA.n2919 VDDA.n2773 3.4105
R2310 VDDA.n2917 VDDA.n2916 3.4105
R2311 VDDA.n2775 VDDA.n2774 3.4105
R2312 VDDA.n2912 VDDA.n2911 3.4105
R2313 VDDA.n2909 VDDA.n2777 3.4105
R2314 VDDA.n2907 VDDA.n2906 3.4105
R2315 VDDA.n2779 VDDA.n2778 3.4105
R2316 VDDA.n2902 VDDA.n2901 3.4105
R2317 VDDA.n2899 VDDA.n2781 3.4105
R2318 VDDA.n2897 VDDA.n2896 3.4105
R2319 VDDA.n2783 VDDA.n2782 3.4105
R2320 VDDA.n2892 VDDA.n2891 3.4105
R2321 VDDA.n2889 VDDA.n2785 3.4105
R2322 VDDA.n2887 VDDA.n2886 3.4105
R2323 VDDA.n2787 VDDA.n2786 3.4105
R2324 VDDA.n2882 VDDA.n2881 3.4105
R2325 VDDA.n2879 VDDA.n2789 3.4105
R2326 VDDA.n2877 VDDA.n2876 3.4105
R2327 VDDA.n2791 VDDA.n2790 3.4105
R2328 VDDA.n2872 VDDA.n2871 3.4105
R2329 VDDA.n2869 VDDA.n2793 3.4105
R2330 VDDA.n2867 VDDA.n2866 3.4105
R2331 VDDA.n2795 VDDA.n2794 3.4105
R2332 VDDA.n2862 VDDA.n2861 3.4105
R2333 VDDA.n2859 VDDA.n2797 3.4105
R2334 VDDA.n2857 VDDA.n2856 3.4105
R2335 VDDA.n2799 VDDA.n2798 3.4105
R2336 VDDA.n2852 VDDA.n2851 3.4105
R2337 VDDA.n2849 VDDA.n2801 3.4105
R2338 VDDA.n2847 VDDA.n2846 3.4105
R2339 VDDA.n2803 VDDA.n2802 3.4105
R2340 VDDA.n2842 VDDA.n2841 3.4105
R2341 VDDA.n2839 VDDA.n2805 3.4105
R2342 VDDA.n2837 VDDA.n2836 3.4105
R2343 VDDA.n2807 VDDA.n2806 3.4105
R2344 VDDA.n2832 VDDA.n2831 3.4105
R2345 VDDA.n2829 VDDA.n2809 3.4105
R2346 VDDA.n2827 VDDA.n2826 3.4105
R2347 VDDA.n2811 VDDA.n2810 3.4105
R2348 VDDA.n2822 VDDA.n2821 3.4105
R2349 VDDA.n2819 VDDA.n2813 3.4105
R2350 VDDA.n2817 VDDA.n2816 3.4105
R2351 VDDA.n2931 VDDA.n2930 3.4105
R2352 VDDA.n194 VDDA.n193 3.4105
R2353 VDDA.n2756 VDDA.n2755 3.4105
R2354 VDDA.n2623 VDDA.n2622 3.4105
R2355 VDDA.n2751 VDDA.n2750 3.4105
R2356 VDDA.n2749 VDDA.n2748 3.4105
R2357 VDDA.n2747 VDDA.n2627 3.4105
R2358 VDDA.n2626 VDDA.n2625 3.4105
R2359 VDDA.n2743 VDDA.n2742 3.4105
R2360 VDDA.n2741 VDDA.n2740 3.4105
R2361 VDDA.n2739 VDDA.n2631 3.4105
R2362 VDDA.n2630 VDDA.n2629 3.4105
R2363 VDDA.n2735 VDDA.n2734 3.4105
R2364 VDDA.n2733 VDDA.n2732 3.4105
R2365 VDDA.n2731 VDDA.n2635 3.4105
R2366 VDDA.n2634 VDDA.n2633 3.4105
R2367 VDDA.n2727 VDDA.n2726 3.4105
R2368 VDDA.n2725 VDDA.n2724 3.4105
R2369 VDDA.n2723 VDDA.n2639 3.4105
R2370 VDDA.n2638 VDDA.n2637 3.4105
R2371 VDDA.n2719 VDDA.n2718 3.4105
R2372 VDDA.n2717 VDDA.n2716 3.4105
R2373 VDDA.n2715 VDDA.n2643 3.4105
R2374 VDDA.n2642 VDDA.n2641 3.4105
R2375 VDDA.n2711 VDDA.n2710 3.4105
R2376 VDDA.n2709 VDDA.n2708 3.4105
R2377 VDDA.n2707 VDDA.n2647 3.4105
R2378 VDDA.n2646 VDDA.n2645 3.4105
R2379 VDDA.n2703 VDDA.n2702 3.4105
R2380 VDDA.n2701 VDDA.n2700 3.4105
R2381 VDDA.n2699 VDDA.n2651 3.4105
R2382 VDDA.n2650 VDDA.n2649 3.4105
R2383 VDDA.n2695 VDDA.n2694 3.4105
R2384 VDDA.n2693 VDDA.n2692 3.4105
R2385 VDDA.n2691 VDDA.n2655 3.4105
R2386 VDDA.n2654 VDDA.n2653 3.4105
R2387 VDDA.n2687 VDDA.n2686 3.4105
R2388 VDDA.n2685 VDDA.n2684 3.4105
R2389 VDDA.n2683 VDDA.n2659 3.4105
R2390 VDDA.n2658 VDDA.n2657 3.4105
R2391 VDDA.n2679 VDDA.n2678 3.4105
R2392 VDDA.n2677 VDDA.n2676 3.4105
R2393 VDDA.n2675 VDDA.n2663 3.4105
R2394 VDDA.n2662 VDDA.n2661 3.4105
R2395 VDDA.n2671 VDDA.n2670 3.4105
R2396 VDDA.n2669 VDDA.n2668 3.4105
R2397 VDDA.n2667 VDDA.n2666 3.4105
R2398 VDDA.n2760 VDDA.n2759 3.4105
R2399 VDDA.n221 VDDA.n220 3.4105
R2400 VDDA.n355 VDDA.n354 3.4105
R2401 VDDA.n353 VDDA.n352 3.4105
R2402 VDDA.n351 VDDA.n225 3.4105
R2403 VDDA.n224 VDDA.n223 3.4105
R2404 VDDA.n347 VDDA.n346 3.4105
R2405 VDDA.n345 VDDA.n344 3.4105
R2406 VDDA.n343 VDDA.n229 3.4105
R2407 VDDA.n228 VDDA.n227 3.4105
R2408 VDDA.n339 VDDA.n338 3.4105
R2409 VDDA.n337 VDDA.n336 3.4105
R2410 VDDA.n335 VDDA.n233 3.4105
R2411 VDDA.n232 VDDA.n231 3.4105
R2412 VDDA.n331 VDDA.n330 3.4105
R2413 VDDA.n329 VDDA.n328 3.4105
R2414 VDDA.n327 VDDA.n237 3.4105
R2415 VDDA.n236 VDDA.n235 3.4105
R2416 VDDA.n323 VDDA.n322 3.4105
R2417 VDDA.n321 VDDA.n320 3.4105
R2418 VDDA.n319 VDDA.n241 3.4105
R2419 VDDA.n240 VDDA.n239 3.4105
R2420 VDDA.n315 VDDA.n314 3.4105
R2421 VDDA.n313 VDDA.n312 3.4105
R2422 VDDA.n311 VDDA.n245 3.4105
R2423 VDDA.n244 VDDA.n243 3.4105
R2424 VDDA.n307 VDDA.n306 3.4105
R2425 VDDA.n305 VDDA.n304 3.4105
R2426 VDDA.n303 VDDA.n249 3.4105
R2427 VDDA.n248 VDDA.n247 3.4105
R2428 VDDA.n299 VDDA.n298 3.4105
R2429 VDDA.n297 VDDA.n296 3.4105
R2430 VDDA.n295 VDDA.n253 3.4105
R2431 VDDA.n252 VDDA.n251 3.4105
R2432 VDDA.n291 VDDA.n290 3.4105
R2433 VDDA.n289 VDDA.n288 3.4105
R2434 VDDA.n287 VDDA.n257 3.4105
R2435 VDDA.n256 VDDA.n255 3.4105
R2436 VDDA.n283 VDDA.n282 3.4105
R2437 VDDA.n281 VDDA.n280 3.4105
R2438 VDDA.n279 VDDA.n261 3.4105
R2439 VDDA.n260 VDDA.n259 3.4105
R2440 VDDA.n275 VDDA.n274 3.4105
R2441 VDDA.n273 VDDA.n272 3.4105
R2442 VDDA.n271 VDDA.n265 3.4105
R2443 VDDA.n264 VDDA.n263 3.4105
R2444 VDDA.n267 VDDA.n266 3.4105
R2445 VDDA.n2597 VDDA.n2596 3.4105
R2446 VDDA.n2581 VDDA.n2421 3.4105
R2447 VDDA.n2579 VDDA.n2578 3.4105
R2448 VDDA.n2423 VDDA.n2422 3.4105
R2449 VDDA.n2574 VDDA.n2573 3.4105
R2450 VDDA.n2571 VDDA.n2425 3.4105
R2451 VDDA.n2569 VDDA.n2568 3.4105
R2452 VDDA.n2427 VDDA.n2426 3.4105
R2453 VDDA.n2564 VDDA.n2563 3.4105
R2454 VDDA.n2561 VDDA.n2429 3.4105
R2455 VDDA.n2559 VDDA.n2558 3.4105
R2456 VDDA.n2431 VDDA.n2430 3.4105
R2457 VDDA.n2554 VDDA.n2553 3.4105
R2458 VDDA.n2551 VDDA.n2433 3.4105
R2459 VDDA.n2549 VDDA.n2548 3.4105
R2460 VDDA.n2435 VDDA.n2434 3.4105
R2461 VDDA.n2544 VDDA.n2543 3.4105
R2462 VDDA.n2541 VDDA.n2437 3.4105
R2463 VDDA.n2539 VDDA.n2538 3.4105
R2464 VDDA.n2439 VDDA.n2438 3.4105
R2465 VDDA.n2534 VDDA.n2533 3.4105
R2466 VDDA.n2531 VDDA.n2441 3.4105
R2467 VDDA.n2529 VDDA.n2528 3.4105
R2468 VDDA.n2443 VDDA.n2442 3.4105
R2469 VDDA.n2524 VDDA.n2523 3.4105
R2470 VDDA.n2521 VDDA.n2445 3.4105
R2471 VDDA.n2519 VDDA.n2518 3.4105
R2472 VDDA.n2447 VDDA.n2446 3.4105
R2473 VDDA.n2514 VDDA.n2513 3.4105
R2474 VDDA.n2511 VDDA.n2449 3.4105
R2475 VDDA.n2509 VDDA.n2508 3.4105
R2476 VDDA.n2451 VDDA.n2450 3.4105
R2477 VDDA.n2504 VDDA.n2503 3.4105
R2478 VDDA.n2501 VDDA.n2453 3.4105
R2479 VDDA.n2499 VDDA.n2498 3.4105
R2480 VDDA.n2455 VDDA.n2454 3.4105
R2481 VDDA.n2494 VDDA.n2493 3.4105
R2482 VDDA.n2491 VDDA.n2457 3.4105
R2483 VDDA.n2489 VDDA.n2488 3.4105
R2484 VDDA.n2459 VDDA.n2458 3.4105
R2485 VDDA.n2484 VDDA.n2483 3.4105
R2486 VDDA.n2481 VDDA.n2461 3.4105
R2487 VDDA.n2479 VDDA.n2478 3.4105
R2488 VDDA.n2463 VDDA.n2462 3.4105
R2489 VDDA.n2474 VDDA.n2473 3.4105
R2490 VDDA.n2471 VDDA.n2465 3.4105
R2491 VDDA.n2469 VDDA.n2468 3.4105
R2492 VDDA.n2583 VDDA.n2582 3.4105
R2493 VDDA.n460 VDDA.n459 3.4105
R2494 VDDA.n1316 VDDA.n1315 3.4105
R2495 VDDA.n1183 VDDA.n1182 3.4105
R2496 VDDA.n1311 VDDA.n1310 3.4105
R2497 VDDA.n1309 VDDA.n1308 3.4105
R2498 VDDA.n1307 VDDA.n1187 3.4105
R2499 VDDA.n1186 VDDA.n1185 3.4105
R2500 VDDA.n1303 VDDA.n1302 3.4105
R2501 VDDA.n1301 VDDA.n1300 3.4105
R2502 VDDA.n1299 VDDA.n1191 3.4105
R2503 VDDA.n1190 VDDA.n1189 3.4105
R2504 VDDA.n1295 VDDA.n1294 3.4105
R2505 VDDA.n1293 VDDA.n1292 3.4105
R2506 VDDA.n1291 VDDA.n1195 3.4105
R2507 VDDA.n1194 VDDA.n1193 3.4105
R2508 VDDA.n1287 VDDA.n1286 3.4105
R2509 VDDA.n1285 VDDA.n1284 3.4105
R2510 VDDA.n1283 VDDA.n1199 3.4105
R2511 VDDA.n1198 VDDA.n1197 3.4105
R2512 VDDA.n1279 VDDA.n1278 3.4105
R2513 VDDA.n1277 VDDA.n1276 3.4105
R2514 VDDA.n1275 VDDA.n1203 3.4105
R2515 VDDA.n1202 VDDA.n1201 3.4105
R2516 VDDA.n1271 VDDA.n1270 3.4105
R2517 VDDA.n1269 VDDA.n1268 3.4105
R2518 VDDA.n1267 VDDA.n1207 3.4105
R2519 VDDA.n1206 VDDA.n1205 3.4105
R2520 VDDA.n1263 VDDA.n1262 3.4105
R2521 VDDA.n1261 VDDA.n1260 3.4105
R2522 VDDA.n1259 VDDA.n1211 3.4105
R2523 VDDA.n1210 VDDA.n1209 3.4105
R2524 VDDA.n1255 VDDA.n1254 3.4105
R2525 VDDA.n1253 VDDA.n1252 3.4105
R2526 VDDA.n1251 VDDA.n1215 3.4105
R2527 VDDA.n1214 VDDA.n1213 3.4105
R2528 VDDA.n1247 VDDA.n1246 3.4105
R2529 VDDA.n1245 VDDA.n1244 3.4105
R2530 VDDA.n1243 VDDA.n1219 3.4105
R2531 VDDA.n1218 VDDA.n1217 3.4105
R2532 VDDA.n1239 VDDA.n1238 3.4105
R2533 VDDA.n1237 VDDA.n1236 3.4105
R2534 VDDA.n1235 VDDA.n1223 3.4105
R2535 VDDA.n1222 VDDA.n1221 3.4105
R2536 VDDA.n1231 VDDA.n1230 3.4105
R2537 VDDA.n1229 VDDA.n1228 3.4105
R2538 VDDA.n1227 VDDA.n1226 3.4105
R2539 VDDA.n2256 VDDA.n2255 3.4105
R2540 VDDA.n487 VDDA.n486 3.4105
R2541 VDDA.n621 VDDA.n620 3.4105
R2542 VDDA.n619 VDDA.n618 3.4105
R2543 VDDA.n617 VDDA.n491 3.4105
R2544 VDDA.n490 VDDA.n489 3.4105
R2545 VDDA.n613 VDDA.n612 3.4105
R2546 VDDA.n611 VDDA.n610 3.4105
R2547 VDDA.n609 VDDA.n495 3.4105
R2548 VDDA.n494 VDDA.n493 3.4105
R2549 VDDA.n605 VDDA.n604 3.4105
R2550 VDDA.n603 VDDA.n602 3.4105
R2551 VDDA.n601 VDDA.n499 3.4105
R2552 VDDA.n498 VDDA.n497 3.4105
R2553 VDDA.n597 VDDA.n596 3.4105
R2554 VDDA.n595 VDDA.n594 3.4105
R2555 VDDA.n593 VDDA.n503 3.4105
R2556 VDDA.n502 VDDA.n501 3.4105
R2557 VDDA.n589 VDDA.n588 3.4105
R2558 VDDA.n587 VDDA.n586 3.4105
R2559 VDDA.n585 VDDA.n507 3.4105
R2560 VDDA.n506 VDDA.n505 3.4105
R2561 VDDA.n581 VDDA.n580 3.4105
R2562 VDDA.n579 VDDA.n578 3.4105
R2563 VDDA.n577 VDDA.n511 3.4105
R2564 VDDA.n510 VDDA.n509 3.4105
R2565 VDDA.n573 VDDA.n572 3.4105
R2566 VDDA.n571 VDDA.n570 3.4105
R2567 VDDA.n569 VDDA.n515 3.4105
R2568 VDDA.n514 VDDA.n513 3.4105
R2569 VDDA.n565 VDDA.n564 3.4105
R2570 VDDA.n563 VDDA.n562 3.4105
R2571 VDDA.n561 VDDA.n519 3.4105
R2572 VDDA.n518 VDDA.n517 3.4105
R2573 VDDA.n557 VDDA.n556 3.4105
R2574 VDDA.n555 VDDA.n554 3.4105
R2575 VDDA.n553 VDDA.n523 3.4105
R2576 VDDA.n522 VDDA.n521 3.4105
R2577 VDDA.n549 VDDA.n548 3.4105
R2578 VDDA.n547 VDDA.n546 3.4105
R2579 VDDA.n545 VDDA.n527 3.4105
R2580 VDDA.n526 VDDA.n525 3.4105
R2581 VDDA.n541 VDDA.n540 3.4105
R2582 VDDA.n539 VDDA.n538 3.4105
R2583 VDDA.n537 VDDA.n531 3.4105
R2584 VDDA.n530 VDDA.n529 3.4105
R2585 VDDA.n533 VDDA.n532 3.4105
R2586 VDDA.n1157 VDDA.n1156 3.4105
R2587 VDDA.n1141 VDDA.n981 3.4105
R2588 VDDA.n1139 VDDA.n1138 3.4105
R2589 VDDA.n983 VDDA.n982 3.4105
R2590 VDDA.n1134 VDDA.n1133 3.4105
R2591 VDDA.n1131 VDDA.n985 3.4105
R2592 VDDA.n1129 VDDA.n1128 3.4105
R2593 VDDA.n987 VDDA.n986 3.4105
R2594 VDDA.n1124 VDDA.n1123 3.4105
R2595 VDDA.n1121 VDDA.n989 3.4105
R2596 VDDA.n1119 VDDA.n1118 3.4105
R2597 VDDA.n991 VDDA.n990 3.4105
R2598 VDDA.n1114 VDDA.n1113 3.4105
R2599 VDDA.n1111 VDDA.n993 3.4105
R2600 VDDA.n1109 VDDA.n1108 3.4105
R2601 VDDA.n995 VDDA.n994 3.4105
R2602 VDDA.n1104 VDDA.n1103 3.4105
R2603 VDDA.n1101 VDDA.n997 3.4105
R2604 VDDA.n1099 VDDA.n1098 3.4105
R2605 VDDA.n999 VDDA.n998 3.4105
R2606 VDDA.n1094 VDDA.n1093 3.4105
R2607 VDDA.n1091 VDDA.n1001 3.4105
R2608 VDDA.n1089 VDDA.n1088 3.4105
R2609 VDDA.n1003 VDDA.n1002 3.4105
R2610 VDDA.n1084 VDDA.n1083 3.4105
R2611 VDDA.n1081 VDDA.n1005 3.4105
R2612 VDDA.n1079 VDDA.n1078 3.4105
R2613 VDDA.n1007 VDDA.n1006 3.4105
R2614 VDDA.n1074 VDDA.n1073 3.4105
R2615 VDDA.n1071 VDDA.n1009 3.4105
R2616 VDDA.n1069 VDDA.n1068 3.4105
R2617 VDDA.n1011 VDDA.n1010 3.4105
R2618 VDDA.n1064 VDDA.n1063 3.4105
R2619 VDDA.n1061 VDDA.n1013 3.4105
R2620 VDDA.n1059 VDDA.n1058 3.4105
R2621 VDDA.n1015 VDDA.n1014 3.4105
R2622 VDDA.n1054 VDDA.n1053 3.4105
R2623 VDDA.n1051 VDDA.n1017 3.4105
R2624 VDDA.n1049 VDDA.n1048 3.4105
R2625 VDDA.n1019 VDDA.n1018 3.4105
R2626 VDDA.n1044 VDDA.n1043 3.4105
R2627 VDDA.n1041 VDDA.n1021 3.4105
R2628 VDDA.n1039 VDDA.n1038 3.4105
R2629 VDDA.n1023 VDDA.n1022 3.4105
R2630 VDDA.n1034 VDDA.n1033 3.4105
R2631 VDDA.n1031 VDDA.n1025 3.4105
R2632 VDDA.n1029 VDDA.n1028 3.4105
R2633 VDDA.n1143 VDDA.n1142 3.4105
R2634 VDDA.n637 VDDA.n636 3.4105
R2635 VDDA.n968 VDDA.n967 3.4105
R2636 VDDA.n835 VDDA.n834 3.4105
R2637 VDDA.n963 VDDA.n962 3.4105
R2638 VDDA.n961 VDDA.n960 3.4105
R2639 VDDA.n959 VDDA.n839 3.4105
R2640 VDDA.n838 VDDA.n837 3.4105
R2641 VDDA.n955 VDDA.n954 3.4105
R2642 VDDA.n953 VDDA.n952 3.4105
R2643 VDDA.n951 VDDA.n843 3.4105
R2644 VDDA.n842 VDDA.n841 3.4105
R2645 VDDA.n947 VDDA.n946 3.4105
R2646 VDDA.n945 VDDA.n944 3.4105
R2647 VDDA.n943 VDDA.n847 3.4105
R2648 VDDA.n846 VDDA.n845 3.4105
R2649 VDDA.n939 VDDA.n938 3.4105
R2650 VDDA.n937 VDDA.n936 3.4105
R2651 VDDA.n935 VDDA.n851 3.4105
R2652 VDDA.n850 VDDA.n849 3.4105
R2653 VDDA.n931 VDDA.n930 3.4105
R2654 VDDA.n929 VDDA.n928 3.4105
R2655 VDDA.n927 VDDA.n855 3.4105
R2656 VDDA.n854 VDDA.n853 3.4105
R2657 VDDA.n923 VDDA.n922 3.4105
R2658 VDDA.n921 VDDA.n920 3.4105
R2659 VDDA.n919 VDDA.n859 3.4105
R2660 VDDA.n858 VDDA.n857 3.4105
R2661 VDDA.n915 VDDA.n914 3.4105
R2662 VDDA.n913 VDDA.n912 3.4105
R2663 VDDA.n911 VDDA.n863 3.4105
R2664 VDDA.n862 VDDA.n861 3.4105
R2665 VDDA.n907 VDDA.n906 3.4105
R2666 VDDA.n905 VDDA.n904 3.4105
R2667 VDDA.n903 VDDA.n867 3.4105
R2668 VDDA.n866 VDDA.n865 3.4105
R2669 VDDA.n899 VDDA.n898 3.4105
R2670 VDDA.n897 VDDA.n896 3.4105
R2671 VDDA.n895 VDDA.n871 3.4105
R2672 VDDA.n870 VDDA.n869 3.4105
R2673 VDDA.n891 VDDA.n890 3.4105
R2674 VDDA.n889 VDDA.n888 3.4105
R2675 VDDA.n887 VDDA.n875 3.4105
R2676 VDDA.n874 VDDA.n873 3.4105
R2677 VDDA.n883 VDDA.n882 3.4105
R2678 VDDA.n881 VDDA.n880 3.4105
R2679 VDDA.n879 VDDA.n878 3.4105
R2680 VDDA.n972 VDDA.n971 3.4105
R2681 VDDA.n663 VDDA.n662 3.4105
R2682 VDDA.n797 VDDA.n796 3.4105
R2683 VDDA.n795 VDDA.n794 3.4105
R2684 VDDA.n793 VDDA.n792 3.4105
R2685 VDDA.n791 VDDA.n665 3.4105
R2686 VDDA.n787 VDDA.n786 3.4105
R2687 VDDA.n785 VDDA.n784 3.4105
R2688 VDDA.n783 VDDA.n782 3.4105
R2689 VDDA.n781 VDDA.n667 3.4105
R2690 VDDA.n777 VDDA.n776 3.4105
R2691 VDDA.n775 VDDA.n774 3.4105
R2692 VDDA.n773 VDDA.n772 3.4105
R2693 VDDA.n771 VDDA.n669 3.4105
R2694 VDDA.n767 VDDA.n766 3.4105
R2695 VDDA.n765 VDDA.n764 3.4105
R2696 VDDA.n763 VDDA.n762 3.4105
R2697 VDDA.n761 VDDA.n671 3.4105
R2698 VDDA.n757 VDDA.n756 3.4105
R2699 VDDA.n755 VDDA.n754 3.4105
R2700 VDDA.n753 VDDA.n752 3.4105
R2701 VDDA.n751 VDDA.n673 3.4105
R2702 VDDA.n747 VDDA.n746 3.4105
R2703 VDDA.n745 VDDA.n744 3.4105
R2704 VDDA.n743 VDDA.n742 3.4105
R2705 VDDA.n741 VDDA.n675 3.4105
R2706 VDDA.n737 VDDA.n736 3.4105
R2707 VDDA.n735 VDDA.n734 3.4105
R2708 VDDA.n733 VDDA.n732 3.4105
R2709 VDDA.n731 VDDA.n677 3.4105
R2710 VDDA.n727 VDDA.n726 3.4105
R2711 VDDA.n725 VDDA.n724 3.4105
R2712 VDDA.n723 VDDA.n722 3.4105
R2713 VDDA.n721 VDDA.n679 3.4105
R2714 VDDA.n717 VDDA.n716 3.4105
R2715 VDDA.n715 VDDA.n714 3.4105
R2716 VDDA.n713 VDDA.n712 3.4105
R2717 VDDA.n711 VDDA.n681 3.4105
R2718 VDDA.n707 VDDA.n706 3.4105
R2719 VDDA.n705 VDDA.n704 3.4105
R2720 VDDA.n703 VDDA.n702 3.4105
R2721 VDDA.n701 VDDA.n683 3.4105
R2722 VDDA.n697 VDDA.n696 3.4105
R2723 VDDA.n695 VDDA.n694 3.4105
R2724 VDDA.n693 VDDA.n692 3.4105
R2725 VDDA.n691 VDDA.n685 3.4105
R2726 VDDA.n687 VDDA.n686 3.4105
R2727 VDDA.n809 VDDA.n808 3.4105
R2728 VDDA.n810 VDDA.n638 3.4105
R2729 VDDA.n810 VDDA.n809 3.4105
R2730 VDDA.n970 VDDA.n811 3.4105
R2731 VDDA.n971 VDDA.n970 3.4105
R2732 VDDA.n1026 VDDA.n461 3.4105
R2733 VDDA.n1142 VDDA.n461 3.4105
R2734 VDDA.n1158 VDDA.n462 3.4105
R2735 VDDA.n1158 VDDA.n1157 3.4105
R2736 VDDA.n2254 VDDA.n1159 3.4105
R2737 VDDA.n2255 VDDA.n2254 3.4105
R2738 VDDA.n2253 VDDA.n1318 3.4105
R2739 VDDA.n2253 VDDA.n2252 3.4105
R2740 VDDA.n2466 VDDA.n195 3.4105
R2741 VDDA.n2582 VDDA.n195 3.4105
R2742 VDDA.n2598 VDDA.n196 3.4105
R2743 VDDA.n2598 VDDA.n2597 3.4105
R2744 VDDA.n2758 VDDA.n2599 3.4105
R2745 VDDA.n2759 VDDA.n2758 3.4105
R2746 VDDA.n2814 VDDA.n17 3.4105
R2747 VDDA.n2930 VDDA.n17 3.4105
R2748 VDDA.n2946 VDDA.n18 3.4105
R2749 VDDA.n2946 VDDA.n2945 3.4105
R2750 VDDA.n1578 VDDA.n1408 3.4105
R2751 VDDA.n1578 VDDA.n1577 3.4105
R2752 VDDA.n1906 VDDA.n1342 3.4105
R2753 VDDA.n1906 VDDA.n1905 3.4105
R2754 VDDA.n1579 VDDA.n1407 3.4105
R2755 VDDA.n1644 VDDA.n1579 3.4105
R2756 VDDA.n3053 VDDA.n15 3.4105
R2757 VDDA.n3053 VDDA.n16 3.4105
R2758 VDDA.n3053 VDDA.n3052 3.4105
R2759 VDDA.n3023 VDDA.n2964 3.4105
R2760 VDDA.n3052 VDDA.n2964 3.4105
R2761 VDDA.n3023 VDDA.n2961 3.4105
R2762 VDDA.n3022 VDDA.n2961 3.4105
R2763 VDDA.n3026 VDDA.n2961 3.4105
R2764 VDDA.n3021 VDDA.n2961 3.4105
R2765 VDDA.n3028 VDDA.n2961 3.4105
R2766 VDDA.n3020 VDDA.n2961 3.4105
R2767 VDDA.n3030 VDDA.n2961 3.4105
R2768 VDDA.n3019 VDDA.n2961 3.4105
R2769 VDDA.n3032 VDDA.n2961 3.4105
R2770 VDDA.n3018 VDDA.n2961 3.4105
R2771 VDDA.n3034 VDDA.n2961 3.4105
R2772 VDDA.n3017 VDDA.n2961 3.4105
R2773 VDDA.n3036 VDDA.n2961 3.4105
R2774 VDDA.n3016 VDDA.n2961 3.4105
R2775 VDDA.n3038 VDDA.n2961 3.4105
R2776 VDDA.n3015 VDDA.n2961 3.4105
R2777 VDDA.n3040 VDDA.n2961 3.4105
R2778 VDDA.n3014 VDDA.n2961 3.4105
R2779 VDDA.n3042 VDDA.n2961 3.4105
R2780 VDDA.n3013 VDDA.n2961 3.4105
R2781 VDDA.n3044 VDDA.n2961 3.4105
R2782 VDDA.n3012 VDDA.n2961 3.4105
R2783 VDDA.n3046 VDDA.n2961 3.4105
R2784 VDDA.n3011 VDDA.n2961 3.4105
R2785 VDDA.n3048 VDDA.n2961 3.4105
R2786 VDDA.n3010 VDDA.n2961 3.4105
R2787 VDDA.n3050 VDDA.n2961 3.4105
R2788 VDDA.n3009 VDDA.n2961 3.4105
R2789 VDDA.n2961 VDDA.n16 3.4105
R2790 VDDA.n3052 VDDA.n2961 3.4105
R2791 VDDA.n3023 VDDA.n2967 3.4105
R2792 VDDA.n3022 VDDA.n2967 3.4105
R2793 VDDA.n3026 VDDA.n2967 3.4105
R2794 VDDA.n3021 VDDA.n2967 3.4105
R2795 VDDA.n3028 VDDA.n2967 3.4105
R2796 VDDA.n3020 VDDA.n2967 3.4105
R2797 VDDA.n3030 VDDA.n2967 3.4105
R2798 VDDA.n3019 VDDA.n2967 3.4105
R2799 VDDA.n3032 VDDA.n2967 3.4105
R2800 VDDA.n3018 VDDA.n2967 3.4105
R2801 VDDA.n3034 VDDA.n2967 3.4105
R2802 VDDA.n3017 VDDA.n2967 3.4105
R2803 VDDA.n3036 VDDA.n2967 3.4105
R2804 VDDA.n3016 VDDA.n2967 3.4105
R2805 VDDA.n3038 VDDA.n2967 3.4105
R2806 VDDA.n3015 VDDA.n2967 3.4105
R2807 VDDA.n3040 VDDA.n2967 3.4105
R2808 VDDA.n3014 VDDA.n2967 3.4105
R2809 VDDA.n3042 VDDA.n2967 3.4105
R2810 VDDA.n3013 VDDA.n2967 3.4105
R2811 VDDA.n3044 VDDA.n2967 3.4105
R2812 VDDA.n3012 VDDA.n2967 3.4105
R2813 VDDA.n3046 VDDA.n2967 3.4105
R2814 VDDA.n3011 VDDA.n2967 3.4105
R2815 VDDA.n3048 VDDA.n2967 3.4105
R2816 VDDA.n3010 VDDA.n2967 3.4105
R2817 VDDA.n3050 VDDA.n2967 3.4105
R2818 VDDA.n3009 VDDA.n2967 3.4105
R2819 VDDA.n2967 VDDA.n16 3.4105
R2820 VDDA.n3052 VDDA.n2967 3.4105
R2821 VDDA.n3023 VDDA.n2960 3.4105
R2822 VDDA.n3022 VDDA.n2960 3.4105
R2823 VDDA.n3026 VDDA.n2960 3.4105
R2824 VDDA.n3021 VDDA.n2960 3.4105
R2825 VDDA.n3028 VDDA.n2960 3.4105
R2826 VDDA.n3020 VDDA.n2960 3.4105
R2827 VDDA.n3030 VDDA.n2960 3.4105
R2828 VDDA.n3019 VDDA.n2960 3.4105
R2829 VDDA.n3032 VDDA.n2960 3.4105
R2830 VDDA.n3018 VDDA.n2960 3.4105
R2831 VDDA.n3034 VDDA.n2960 3.4105
R2832 VDDA.n3017 VDDA.n2960 3.4105
R2833 VDDA.n3036 VDDA.n2960 3.4105
R2834 VDDA.n3016 VDDA.n2960 3.4105
R2835 VDDA.n3038 VDDA.n2960 3.4105
R2836 VDDA.n3015 VDDA.n2960 3.4105
R2837 VDDA.n3040 VDDA.n2960 3.4105
R2838 VDDA.n3014 VDDA.n2960 3.4105
R2839 VDDA.n3042 VDDA.n2960 3.4105
R2840 VDDA.n3013 VDDA.n2960 3.4105
R2841 VDDA.n3044 VDDA.n2960 3.4105
R2842 VDDA.n3012 VDDA.n2960 3.4105
R2843 VDDA.n3046 VDDA.n2960 3.4105
R2844 VDDA.n3011 VDDA.n2960 3.4105
R2845 VDDA.n3048 VDDA.n2960 3.4105
R2846 VDDA.n3010 VDDA.n2960 3.4105
R2847 VDDA.n3050 VDDA.n2960 3.4105
R2848 VDDA.n3009 VDDA.n2960 3.4105
R2849 VDDA.n2960 VDDA.n16 3.4105
R2850 VDDA.n3052 VDDA.n2960 3.4105
R2851 VDDA.n3023 VDDA.n2970 3.4105
R2852 VDDA.n3022 VDDA.n2970 3.4105
R2853 VDDA.n3026 VDDA.n2970 3.4105
R2854 VDDA.n3021 VDDA.n2970 3.4105
R2855 VDDA.n3028 VDDA.n2970 3.4105
R2856 VDDA.n3020 VDDA.n2970 3.4105
R2857 VDDA.n3030 VDDA.n2970 3.4105
R2858 VDDA.n3019 VDDA.n2970 3.4105
R2859 VDDA.n3032 VDDA.n2970 3.4105
R2860 VDDA.n3018 VDDA.n2970 3.4105
R2861 VDDA.n3034 VDDA.n2970 3.4105
R2862 VDDA.n3017 VDDA.n2970 3.4105
R2863 VDDA.n3036 VDDA.n2970 3.4105
R2864 VDDA.n3016 VDDA.n2970 3.4105
R2865 VDDA.n3038 VDDA.n2970 3.4105
R2866 VDDA.n3015 VDDA.n2970 3.4105
R2867 VDDA.n3040 VDDA.n2970 3.4105
R2868 VDDA.n3014 VDDA.n2970 3.4105
R2869 VDDA.n3042 VDDA.n2970 3.4105
R2870 VDDA.n3013 VDDA.n2970 3.4105
R2871 VDDA.n3044 VDDA.n2970 3.4105
R2872 VDDA.n3012 VDDA.n2970 3.4105
R2873 VDDA.n3046 VDDA.n2970 3.4105
R2874 VDDA.n3011 VDDA.n2970 3.4105
R2875 VDDA.n3048 VDDA.n2970 3.4105
R2876 VDDA.n3010 VDDA.n2970 3.4105
R2877 VDDA.n3050 VDDA.n2970 3.4105
R2878 VDDA.n3009 VDDA.n2970 3.4105
R2879 VDDA.n2970 VDDA.n16 3.4105
R2880 VDDA.n3052 VDDA.n2970 3.4105
R2881 VDDA.n3023 VDDA.n2959 3.4105
R2882 VDDA.n3022 VDDA.n2959 3.4105
R2883 VDDA.n3026 VDDA.n2959 3.4105
R2884 VDDA.n3021 VDDA.n2959 3.4105
R2885 VDDA.n3028 VDDA.n2959 3.4105
R2886 VDDA.n3020 VDDA.n2959 3.4105
R2887 VDDA.n3030 VDDA.n2959 3.4105
R2888 VDDA.n3019 VDDA.n2959 3.4105
R2889 VDDA.n3032 VDDA.n2959 3.4105
R2890 VDDA.n3018 VDDA.n2959 3.4105
R2891 VDDA.n3034 VDDA.n2959 3.4105
R2892 VDDA.n3017 VDDA.n2959 3.4105
R2893 VDDA.n3036 VDDA.n2959 3.4105
R2894 VDDA.n3016 VDDA.n2959 3.4105
R2895 VDDA.n3038 VDDA.n2959 3.4105
R2896 VDDA.n3015 VDDA.n2959 3.4105
R2897 VDDA.n3040 VDDA.n2959 3.4105
R2898 VDDA.n3014 VDDA.n2959 3.4105
R2899 VDDA.n3042 VDDA.n2959 3.4105
R2900 VDDA.n3013 VDDA.n2959 3.4105
R2901 VDDA.n3044 VDDA.n2959 3.4105
R2902 VDDA.n3012 VDDA.n2959 3.4105
R2903 VDDA.n3046 VDDA.n2959 3.4105
R2904 VDDA.n3011 VDDA.n2959 3.4105
R2905 VDDA.n3048 VDDA.n2959 3.4105
R2906 VDDA.n3010 VDDA.n2959 3.4105
R2907 VDDA.n3050 VDDA.n2959 3.4105
R2908 VDDA.n3009 VDDA.n2959 3.4105
R2909 VDDA.n2959 VDDA.n16 3.4105
R2910 VDDA.n3052 VDDA.n2959 3.4105
R2911 VDDA.n3023 VDDA.n2973 3.4105
R2912 VDDA.n3022 VDDA.n2973 3.4105
R2913 VDDA.n3026 VDDA.n2973 3.4105
R2914 VDDA.n3021 VDDA.n2973 3.4105
R2915 VDDA.n3028 VDDA.n2973 3.4105
R2916 VDDA.n3020 VDDA.n2973 3.4105
R2917 VDDA.n3030 VDDA.n2973 3.4105
R2918 VDDA.n3019 VDDA.n2973 3.4105
R2919 VDDA.n3032 VDDA.n2973 3.4105
R2920 VDDA.n3018 VDDA.n2973 3.4105
R2921 VDDA.n3034 VDDA.n2973 3.4105
R2922 VDDA.n3017 VDDA.n2973 3.4105
R2923 VDDA.n3036 VDDA.n2973 3.4105
R2924 VDDA.n3016 VDDA.n2973 3.4105
R2925 VDDA.n3038 VDDA.n2973 3.4105
R2926 VDDA.n3015 VDDA.n2973 3.4105
R2927 VDDA.n3040 VDDA.n2973 3.4105
R2928 VDDA.n3014 VDDA.n2973 3.4105
R2929 VDDA.n3042 VDDA.n2973 3.4105
R2930 VDDA.n3013 VDDA.n2973 3.4105
R2931 VDDA.n3044 VDDA.n2973 3.4105
R2932 VDDA.n3012 VDDA.n2973 3.4105
R2933 VDDA.n3046 VDDA.n2973 3.4105
R2934 VDDA.n3011 VDDA.n2973 3.4105
R2935 VDDA.n3048 VDDA.n2973 3.4105
R2936 VDDA.n3010 VDDA.n2973 3.4105
R2937 VDDA.n3050 VDDA.n2973 3.4105
R2938 VDDA.n3009 VDDA.n2973 3.4105
R2939 VDDA.n2973 VDDA.n16 3.4105
R2940 VDDA.n3052 VDDA.n2973 3.4105
R2941 VDDA.n3023 VDDA.n2958 3.4105
R2942 VDDA.n3022 VDDA.n2958 3.4105
R2943 VDDA.n3026 VDDA.n2958 3.4105
R2944 VDDA.n3021 VDDA.n2958 3.4105
R2945 VDDA.n3028 VDDA.n2958 3.4105
R2946 VDDA.n3020 VDDA.n2958 3.4105
R2947 VDDA.n3030 VDDA.n2958 3.4105
R2948 VDDA.n3019 VDDA.n2958 3.4105
R2949 VDDA.n3032 VDDA.n2958 3.4105
R2950 VDDA.n3018 VDDA.n2958 3.4105
R2951 VDDA.n3034 VDDA.n2958 3.4105
R2952 VDDA.n3017 VDDA.n2958 3.4105
R2953 VDDA.n3036 VDDA.n2958 3.4105
R2954 VDDA.n3016 VDDA.n2958 3.4105
R2955 VDDA.n3038 VDDA.n2958 3.4105
R2956 VDDA.n3015 VDDA.n2958 3.4105
R2957 VDDA.n3040 VDDA.n2958 3.4105
R2958 VDDA.n3014 VDDA.n2958 3.4105
R2959 VDDA.n3042 VDDA.n2958 3.4105
R2960 VDDA.n3013 VDDA.n2958 3.4105
R2961 VDDA.n3044 VDDA.n2958 3.4105
R2962 VDDA.n3012 VDDA.n2958 3.4105
R2963 VDDA.n3046 VDDA.n2958 3.4105
R2964 VDDA.n3011 VDDA.n2958 3.4105
R2965 VDDA.n3048 VDDA.n2958 3.4105
R2966 VDDA.n3010 VDDA.n2958 3.4105
R2967 VDDA.n3050 VDDA.n2958 3.4105
R2968 VDDA.n3009 VDDA.n2958 3.4105
R2969 VDDA.n2958 VDDA.n16 3.4105
R2970 VDDA.n3052 VDDA.n2958 3.4105
R2971 VDDA.n3023 VDDA.n2976 3.4105
R2972 VDDA.n3022 VDDA.n2976 3.4105
R2973 VDDA.n3026 VDDA.n2976 3.4105
R2974 VDDA.n3021 VDDA.n2976 3.4105
R2975 VDDA.n3028 VDDA.n2976 3.4105
R2976 VDDA.n3020 VDDA.n2976 3.4105
R2977 VDDA.n3030 VDDA.n2976 3.4105
R2978 VDDA.n3019 VDDA.n2976 3.4105
R2979 VDDA.n3032 VDDA.n2976 3.4105
R2980 VDDA.n3018 VDDA.n2976 3.4105
R2981 VDDA.n3034 VDDA.n2976 3.4105
R2982 VDDA.n3017 VDDA.n2976 3.4105
R2983 VDDA.n3036 VDDA.n2976 3.4105
R2984 VDDA.n3016 VDDA.n2976 3.4105
R2985 VDDA.n3038 VDDA.n2976 3.4105
R2986 VDDA.n3015 VDDA.n2976 3.4105
R2987 VDDA.n3040 VDDA.n2976 3.4105
R2988 VDDA.n3014 VDDA.n2976 3.4105
R2989 VDDA.n3042 VDDA.n2976 3.4105
R2990 VDDA.n3013 VDDA.n2976 3.4105
R2991 VDDA.n3044 VDDA.n2976 3.4105
R2992 VDDA.n3012 VDDA.n2976 3.4105
R2993 VDDA.n3046 VDDA.n2976 3.4105
R2994 VDDA.n3011 VDDA.n2976 3.4105
R2995 VDDA.n3048 VDDA.n2976 3.4105
R2996 VDDA.n3010 VDDA.n2976 3.4105
R2997 VDDA.n3050 VDDA.n2976 3.4105
R2998 VDDA.n3009 VDDA.n2976 3.4105
R2999 VDDA.n2976 VDDA.n16 3.4105
R3000 VDDA.n3052 VDDA.n2976 3.4105
R3001 VDDA.n3023 VDDA.n2957 3.4105
R3002 VDDA.n3022 VDDA.n2957 3.4105
R3003 VDDA.n3026 VDDA.n2957 3.4105
R3004 VDDA.n3021 VDDA.n2957 3.4105
R3005 VDDA.n3028 VDDA.n2957 3.4105
R3006 VDDA.n3020 VDDA.n2957 3.4105
R3007 VDDA.n3030 VDDA.n2957 3.4105
R3008 VDDA.n3019 VDDA.n2957 3.4105
R3009 VDDA.n3032 VDDA.n2957 3.4105
R3010 VDDA.n3018 VDDA.n2957 3.4105
R3011 VDDA.n3034 VDDA.n2957 3.4105
R3012 VDDA.n3017 VDDA.n2957 3.4105
R3013 VDDA.n3036 VDDA.n2957 3.4105
R3014 VDDA.n3016 VDDA.n2957 3.4105
R3015 VDDA.n3038 VDDA.n2957 3.4105
R3016 VDDA.n3015 VDDA.n2957 3.4105
R3017 VDDA.n3040 VDDA.n2957 3.4105
R3018 VDDA.n3014 VDDA.n2957 3.4105
R3019 VDDA.n3042 VDDA.n2957 3.4105
R3020 VDDA.n3013 VDDA.n2957 3.4105
R3021 VDDA.n3044 VDDA.n2957 3.4105
R3022 VDDA.n3012 VDDA.n2957 3.4105
R3023 VDDA.n3046 VDDA.n2957 3.4105
R3024 VDDA.n3011 VDDA.n2957 3.4105
R3025 VDDA.n3048 VDDA.n2957 3.4105
R3026 VDDA.n3010 VDDA.n2957 3.4105
R3027 VDDA.n3050 VDDA.n2957 3.4105
R3028 VDDA.n3009 VDDA.n2957 3.4105
R3029 VDDA.n2957 VDDA.n16 3.4105
R3030 VDDA.n3052 VDDA.n2957 3.4105
R3031 VDDA.n3023 VDDA.n2979 3.4105
R3032 VDDA.n3022 VDDA.n2979 3.4105
R3033 VDDA.n3026 VDDA.n2979 3.4105
R3034 VDDA.n3021 VDDA.n2979 3.4105
R3035 VDDA.n3028 VDDA.n2979 3.4105
R3036 VDDA.n3020 VDDA.n2979 3.4105
R3037 VDDA.n3030 VDDA.n2979 3.4105
R3038 VDDA.n3019 VDDA.n2979 3.4105
R3039 VDDA.n3032 VDDA.n2979 3.4105
R3040 VDDA.n3018 VDDA.n2979 3.4105
R3041 VDDA.n3034 VDDA.n2979 3.4105
R3042 VDDA.n3017 VDDA.n2979 3.4105
R3043 VDDA.n3036 VDDA.n2979 3.4105
R3044 VDDA.n3016 VDDA.n2979 3.4105
R3045 VDDA.n3038 VDDA.n2979 3.4105
R3046 VDDA.n3015 VDDA.n2979 3.4105
R3047 VDDA.n3040 VDDA.n2979 3.4105
R3048 VDDA.n3014 VDDA.n2979 3.4105
R3049 VDDA.n3042 VDDA.n2979 3.4105
R3050 VDDA.n3013 VDDA.n2979 3.4105
R3051 VDDA.n3044 VDDA.n2979 3.4105
R3052 VDDA.n3012 VDDA.n2979 3.4105
R3053 VDDA.n3046 VDDA.n2979 3.4105
R3054 VDDA.n3011 VDDA.n2979 3.4105
R3055 VDDA.n3048 VDDA.n2979 3.4105
R3056 VDDA.n3010 VDDA.n2979 3.4105
R3057 VDDA.n3050 VDDA.n2979 3.4105
R3058 VDDA.n3009 VDDA.n2979 3.4105
R3059 VDDA.n2979 VDDA.n16 3.4105
R3060 VDDA.n3052 VDDA.n2979 3.4105
R3061 VDDA.n3023 VDDA.n2956 3.4105
R3062 VDDA.n3022 VDDA.n2956 3.4105
R3063 VDDA.n3026 VDDA.n2956 3.4105
R3064 VDDA.n3021 VDDA.n2956 3.4105
R3065 VDDA.n3028 VDDA.n2956 3.4105
R3066 VDDA.n3020 VDDA.n2956 3.4105
R3067 VDDA.n3030 VDDA.n2956 3.4105
R3068 VDDA.n3019 VDDA.n2956 3.4105
R3069 VDDA.n3032 VDDA.n2956 3.4105
R3070 VDDA.n3018 VDDA.n2956 3.4105
R3071 VDDA.n3034 VDDA.n2956 3.4105
R3072 VDDA.n3017 VDDA.n2956 3.4105
R3073 VDDA.n3036 VDDA.n2956 3.4105
R3074 VDDA.n3016 VDDA.n2956 3.4105
R3075 VDDA.n3038 VDDA.n2956 3.4105
R3076 VDDA.n3015 VDDA.n2956 3.4105
R3077 VDDA.n3040 VDDA.n2956 3.4105
R3078 VDDA.n3014 VDDA.n2956 3.4105
R3079 VDDA.n3042 VDDA.n2956 3.4105
R3080 VDDA.n3013 VDDA.n2956 3.4105
R3081 VDDA.n3044 VDDA.n2956 3.4105
R3082 VDDA.n3012 VDDA.n2956 3.4105
R3083 VDDA.n3046 VDDA.n2956 3.4105
R3084 VDDA.n3011 VDDA.n2956 3.4105
R3085 VDDA.n3048 VDDA.n2956 3.4105
R3086 VDDA.n3010 VDDA.n2956 3.4105
R3087 VDDA.n3050 VDDA.n2956 3.4105
R3088 VDDA.n3009 VDDA.n2956 3.4105
R3089 VDDA.n2956 VDDA.n16 3.4105
R3090 VDDA.n3052 VDDA.n2956 3.4105
R3091 VDDA.n3023 VDDA.n2982 3.4105
R3092 VDDA.n3022 VDDA.n2982 3.4105
R3093 VDDA.n3026 VDDA.n2982 3.4105
R3094 VDDA.n3021 VDDA.n2982 3.4105
R3095 VDDA.n3028 VDDA.n2982 3.4105
R3096 VDDA.n3020 VDDA.n2982 3.4105
R3097 VDDA.n3030 VDDA.n2982 3.4105
R3098 VDDA.n3019 VDDA.n2982 3.4105
R3099 VDDA.n3032 VDDA.n2982 3.4105
R3100 VDDA.n3018 VDDA.n2982 3.4105
R3101 VDDA.n3034 VDDA.n2982 3.4105
R3102 VDDA.n3017 VDDA.n2982 3.4105
R3103 VDDA.n3036 VDDA.n2982 3.4105
R3104 VDDA.n3016 VDDA.n2982 3.4105
R3105 VDDA.n3038 VDDA.n2982 3.4105
R3106 VDDA.n3015 VDDA.n2982 3.4105
R3107 VDDA.n3040 VDDA.n2982 3.4105
R3108 VDDA.n3014 VDDA.n2982 3.4105
R3109 VDDA.n3042 VDDA.n2982 3.4105
R3110 VDDA.n3013 VDDA.n2982 3.4105
R3111 VDDA.n3044 VDDA.n2982 3.4105
R3112 VDDA.n3012 VDDA.n2982 3.4105
R3113 VDDA.n3046 VDDA.n2982 3.4105
R3114 VDDA.n3011 VDDA.n2982 3.4105
R3115 VDDA.n3048 VDDA.n2982 3.4105
R3116 VDDA.n3010 VDDA.n2982 3.4105
R3117 VDDA.n3050 VDDA.n2982 3.4105
R3118 VDDA.n3009 VDDA.n2982 3.4105
R3119 VDDA.n2982 VDDA.n16 3.4105
R3120 VDDA.n3052 VDDA.n2982 3.4105
R3121 VDDA.n3023 VDDA.n2955 3.4105
R3122 VDDA.n3022 VDDA.n2955 3.4105
R3123 VDDA.n3026 VDDA.n2955 3.4105
R3124 VDDA.n3021 VDDA.n2955 3.4105
R3125 VDDA.n3028 VDDA.n2955 3.4105
R3126 VDDA.n3020 VDDA.n2955 3.4105
R3127 VDDA.n3030 VDDA.n2955 3.4105
R3128 VDDA.n3019 VDDA.n2955 3.4105
R3129 VDDA.n3032 VDDA.n2955 3.4105
R3130 VDDA.n3018 VDDA.n2955 3.4105
R3131 VDDA.n3034 VDDA.n2955 3.4105
R3132 VDDA.n3017 VDDA.n2955 3.4105
R3133 VDDA.n3036 VDDA.n2955 3.4105
R3134 VDDA.n3016 VDDA.n2955 3.4105
R3135 VDDA.n3038 VDDA.n2955 3.4105
R3136 VDDA.n3015 VDDA.n2955 3.4105
R3137 VDDA.n3040 VDDA.n2955 3.4105
R3138 VDDA.n3014 VDDA.n2955 3.4105
R3139 VDDA.n3042 VDDA.n2955 3.4105
R3140 VDDA.n3013 VDDA.n2955 3.4105
R3141 VDDA.n3044 VDDA.n2955 3.4105
R3142 VDDA.n3012 VDDA.n2955 3.4105
R3143 VDDA.n3046 VDDA.n2955 3.4105
R3144 VDDA.n3011 VDDA.n2955 3.4105
R3145 VDDA.n3048 VDDA.n2955 3.4105
R3146 VDDA.n3010 VDDA.n2955 3.4105
R3147 VDDA.n3050 VDDA.n2955 3.4105
R3148 VDDA.n3009 VDDA.n2955 3.4105
R3149 VDDA.n2955 VDDA.n16 3.4105
R3150 VDDA.n3052 VDDA.n2955 3.4105
R3151 VDDA.n3023 VDDA.n2985 3.4105
R3152 VDDA.n3022 VDDA.n2985 3.4105
R3153 VDDA.n3026 VDDA.n2985 3.4105
R3154 VDDA.n3021 VDDA.n2985 3.4105
R3155 VDDA.n3028 VDDA.n2985 3.4105
R3156 VDDA.n3020 VDDA.n2985 3.4105
R3157 VDDA.n3030 VDDA.n2985 3.4105
R3158 VDDA.n3019 VDDA.n2985 3.4105
R3159 VDDA.n3032 VDDA.n2985 3.4105
R3160 VDDA.n3018 VDDA.n2985 3.4105
R3161 VDDA.n3034 VDDA.n2985 3.4105
R3162 VDDA.n3017 VDDA.n2985 3.4105
R3163 VDDA.n3036 VDDA.n2985 3.4105
R3164 VDDA.n3016 VDDA.n2985 3.4105
R3165 VDDA.n3038 VDDA.n2985 3.4105
R3166 VDDA.n3015 VDDA.n2985 3.4105
R3167 VDDA.n3040 VDDA.n2985 3.4105
R3168 VDDA.n3014 VDDA.n2985 3.4105
R3169 VDDA.n3042 VDDA.n2985 3.4105
R3170 VDDA.n3013 VDDA.n2985 3.4105
R3171 VDDA.n3044 VDDA.n2985 3.4105
R3172 VDDA.n3012 VDDA.n2985 3.4105
R3173 VDDA.n3046 VDDA.n2985 3.4105
R3174 VDDA.n3011 VDDA.n2985 3.4105
R3175 VDDA.n3048 VDDA.n2985 3.4105
R3176 VDDA.n3010 VDDA.n2985 3.4105
R3177 VDDA.n3050 VDDA.n2985 3.4105
R3178 VDDA.n3009 VDDA.n2985 3.4105
R3179 VDDA.n2985 VDDA.n16 3.4105
R3180 VDDA.n3052 VDDA.n2985 3.4105
R3181 VDDA.n3023 VDDA.n2954 3.4105
R3182 VDDA.n3022 VDDA.n2954 3.4105
R3183 VDDA.n3026 VDDA.n2954 3.4105
R3184 VDDA.n3021 VDDA.n2954 3.4105
R3185 VDDA.n3028 VDDA.n2954 3.4105
R3186 VDDA.n3020 VDDA.n2954 3.4105
R3187 VDDA.n3030 VDDA.n2954 3.4105
R3188 VDDA.n3019 VDDA.n2954 3.4105
R3189 VDDA.n3032 VDDA.n2954 3.4105
R3190 VDDA.n3018 VDDA.n2954 3.4105
R3191 VDDA.n3034 VDDA.n2954 3.4105
R3192 VDDA.n3017 VDDA.n2954 3.4105
R3193 VDDA.n3036 VDDA.n2954 3.4105
R3194 VDDA.n3016 VDDA.n2954 3.4105
R3195 VDDA.n3038 VDDA.n2954 3.4105
R3196 VDDA.n3015 VDDA.n2954 3.4105
R3197 VDDA.n3040 VDDA.n2954 3.4105
R3198 VDDA.n3014 VDDA.n2954 3.4105
R3199 VDDA.n3042 VDDA.n2954 3.4105
R3200 VDDA.n3013 VDDA.n2954 3.4105
R3201 VDDA.n3044 VDDA.n2954 3.4105
R3202 VDDA.n3012 VDDA.n2954 3.4105
R3203 VDDA.n3046 VDDA.n2954 3.4105
R3204 VDDA.n3011 VDDA.n2954 3.4105
R3205 VDDA.n3048 VDDA.n2954 3.4105
R3206 VDDA.n3010 VDDA.n2954 3.4105
R3207 VDDA.n3050 VDDA.n2954 3.4105
R3208 VDDA.n3009 VDDA.n2954 3.4105
R3209 VDDA.n2954 VDDA.n16 3.4105
R3210 VDDA.n3052 VDDA.n2954 3.4105
R3211 VDDA.n3023 VDDA.n2988 3.4105
R3212 VDDA.n3022 VDDA.n2988 3.4105
R3213 VDDA.n3026 VDDA.n2988 3.4105
R3214 VDDA.n3021 VDDA.n2988 3.4105
R3215 VDDA.n3028 VDDA.n2988 3.4105
R3216 VDDA.n3020 VDDA.n2988 3.4105
R3217 VDDA.n3030 VDDA.n2988 3.4105
R3218 VDDA.n3019 VDDA.n2988 3.4105
R3219 VDDA.n3032 VDDA.n2988 3.4105
R3220 VDDA.n3018 VDDA.n2988 3.4105
R3221 VDDA.n3034 VDDA.n2988 3.4105
R3222 VDDA.n3017 VDDA.n2988 3.4105
R3223 VDDA.n3036 VDDA.n2988 3.4105
R3224 VDDA.n3016 VDDA.n2988 3.4105
R3225 VDDA.n3038 VDDA.n2988 3.4105
R3226 VDDA.n3015 VDDA.n2988 3.4105
R3227 VDDA.n3040 VDDA.n2988 3.4105
R3228 VDDA.n3014 VDDA.n2988 3.4105
R3229 VDDA.n3042 VDDA.n2988 3.4105
R3230 VDDA.n3013 VDDA.n2988 3.4105
R3231 VDDA.n3044 VDDA.n2988 3.4105
R3232 VDDA.n3012 VDDA.n2988 3.4105
R3233 VDDA.n3046 VDDA.n2988 3.4105
R3234 VDDA.n3011 VDDA.n2988 3.4105
R3235 VDDA.n3048 VDDA.n2988 3.4105
R3236 VDDA.n3010 VDDA.n2988 3.4105
R3237 VDDA.n3050 VDDA.n2988 3.4105
R3238 VDDA.n3009 VDDA.n2988 3.4105
R3239 VDDA.n2988 VDDA.n16 3.4105
R3240 VDDA.n3052 VDDA.n2988 3.4105
R3241 VDDA.n3023 VDDA.n2953 3.4105
R3242 VDDA.n3022 VDDA.n2953 3.4105
R3243 VDDA.n3026 VDDA.n2953 3.4105
R3244 VDDA.n3021 VDDA.n2953 3.4105
R3245 VDDA.n3028 VDDA.n2953 3.4105
R3246 VDDA.n3020 VDDA.n2953 3.4105
R3247 VDDA.n3030 VDDA.n2953 3.4105
R3248 VDDA.n3019 VDDA.n2953 3.4105
R3249 VDDA.n3032 VDDA.n2953 3.4105
R3250 VDDA.n3018 VDDA.n2953 3.4105
R3251 VDDA.n3034 VDDA.n2953 3.4105
R3252 VDDA.n3017 VDDA.n2953 3.4105
R3253 VDDA.n3036 VDDA.n2953 3.4105
R3254 VDDA.n3016 VDDA.n2953 3.4105
R3255 VDDA.n3038 VDDA.n2953 3.4105
R3256 VDDA.n3015 VDDA.n2953 3.4105
R3257 VDDA.n3040 VDDA.n2953 3.4105
R3258 VDDA.n3014 VDDA.n2953 3.4105
R3259 VDDA.n3042 VDDA.n2953 3.4105
R3260 VDDA.n3013 VDDA.n2953 3.4105
R3261 VDDA.n3044 VDDA.n2953 3.4105
R3262 VDDA.n3012 VDDA.n2953 3.4105
R3263 VDDA.n3046 VDDA.n2953 3.4105
R3264 VDDA.n3011 VDDA.n2953 3.4105
R3265 VDDA.n3048 VDDA.n2953 3.4105
R3266 VDDA.n3010 VDDA.n2953 3.4105
R3267 VDDA.n3050 VDDA.n2953 3.4105
R3268 VDDA.n3009 VDDA.n2953 3.4105
R3269 VDDA.n2953 VDDA.n16 3.4105
R3270 VDDA.n3052 VDDA.n2953 3.4105
R3271 VDDA.n3023 VDDA.n2991 3.4105
R3272 VDDA.n3022 VDDA.n2991 3.4105
R3273 VDDA.n3026 VDDA.n2991 3.4105
R3274 VDDA.n3021 VDDA.n2991 3.4105
R3275 VDDA.n3028 VDDA.n2991 3.4105
R3276 VDDA.n3020 VDDA.n2991 3.4105
R3277 VDDA.n3030 VDDA.n2991 3.4105
R3278 VDDA.n3019 VDDA.n2991 3.4105
R3279 VDDA.n3032 VDDA.n2991 3.4105
R3280 VDDA.n3018 VDDA.n2991 3.4105
R3281 VDDA.n3034 VDDA.n2991 3.4105
R3282 VDDA.n3017 VDDA.n2991 3.4105
R3283 VDDA.n3036 VDDA.n2991 3.4105
R3284 VDDA.n3016 VDDA.n2991 3.4105
R3285 VDDA.n3038 VDDA.n2991 3.4105
R3286 VDDA.n3015 VDDA.n2991 3.4105
R3287 VDDA.n3040 VDDA.n2991 3.4105
R3288 VDDA.n3014 VDDA.n2991 3.4105
R3289 VDDA.n3042 VDDA.n2991 3.4105
R3290 VDDA.n3013 VDDA.n2991 3.4105
R3291 VDDA.n3044 VDDA.n2991 3.4105
R3292 VDDA.n3012 VDDA.n2991 3.4105
R3293 VDDA.n3046 VDDA.n2991 3.4105
R3294 VDDA.n3011 VDDA.n2991 3.4105
R3295 VDDA.n3048 VDDA.n2991 3.4105
R3296 VDDA.n3010 VDDA.n2991 3.4105
R3297 VDDA.n3050 VDDA.n2991 3.4105
R3298 VDDA.n3009 VDDA.n2991 3.4105
R3299 VDDA.n2991 VDDA.n16 3.4105
R3300 VDDA.n3052 VDDA.n2991 3.4105
R3301 VDDA.n3023 VDDA.n2952 3.4105
R3302 VDDA.n3022 VDDA.n2952 3.4105
R3303 VDDA.n3026 VDDA.n2952 3.4105
R3304 VDDA.n3021 VDDA.n2952 3.4105
R3305 VDDA.n3028 VDDA.n2952 3.4105
R3306 VDDA.n3020 VDDA.n2952 3.4105
R3307 VDDA.n3030 VDDA.n2952 3.4105
R3308 VDDA.n3019 VDDA.n2952 3.4105
R3309 VDDA.n3032 VDDA.n2952 3.4105
R3310 VDDA.n3018 VDDA.n2952 3.4105
R3311 VDDA.n3034 VDDA.n2952 3.4105
R3312 VDDA.n3017 VDDA.n2952 3.4105
R3313 VDDA.n3036 VDDA.n2952 3.4105
R3314 VDDA.n3016 VDDA.n2952 3.4105
R3315 VDDA.n3038 VDDA.n2952 3.4105
R3316 VDDA.n3015 VDDA.n2952 3.4105
R3317 VDDA.n3040 VDDA.n2952 3.4105
R3318 VDDA.n3014 VDDA.n2952 3.4105
R3319 VDDA.n3042 VDDA.n2952 3.4105
R3320 VDDA.n3013 VDDA.n2952 3.4105
R3321 VDDA.n3044 VDDA.n2952 3.4105
R3322 VDDA.n3012 VDDA.n2952 3.4105
R3323 VDDA.n3046 VDDA.n2952 3.4105
R3324 VDDA.n3011 VDDA.n2952 3.4105
R3325 VDDA.n3048 VDDA.n2952 3.4105
R3326 VDDA.n3010 VDDA.n2952 3.4105
R3327 VDDA.n3050 VDDA.n2952 3.4105
R3328 VDDA.n3009 VDDA.n2952 3.4105
R3329 VDDA.n2952 VDDA.n16 3.4105
R3330 VDDA.n3052 VDDA.n2952 3.4105
R3331 VDDA.n3023 VDDA.n2994 3.4105
R3332 VDDA.n3022 VDDA.n2994 3.4105
R3333 VDDA.n3026 VDDA.n2994 3.4105
R3334 VDDA.n3021 VDDA.n2994 3.4105
R3335 VDDA.n3028 VDDA.n2994 3.4105
R3336 VDDA.n3020 VDDA.n2994 3.4105
R3337 VDDA.n3030 VDDA.n2994 3.4105
R3338 VDDA.n3019 VDDA.n2994 3.4105
R3339 VDDA.n3032 VDDA.n2994 3.4105
R3340 VDDA.n3018 VDDA.n2994 3.4105
R3341 VDDA.n3034 VDDA.n2994 3.4105
R3342 VDDA.n3017 VDDA.n2994 3.4105
R3343 VDDA.n3036 VDDA.n2994 3.4105
R3344 VDDA.n3016 VDDA.n2994 3.4105
R3345 VDDA.n3038 VDDA.n2994 3.4105
R3346 VDDA.n3015 VDDA.n2994 3.4105
R3347 VDDA.n3040 VDDA.n2994 3.4105
R3348 VDDA.n3014 VDDA.n2994 3.4105
R3349 VDDA.n3042 VDDA.n2994 3.4105
R3350 VDDA.n3013 VDDA.n2994 3.4105
R3351 VDDA.n3044 VDDA.n2994 3.4105
R3352 VDDA.n3012 VDDA.n2994 3.4105
R3353 VDDA.n3046 VDDA.n2994 3.4105
R3354 VDDA.n3011 VDDA.n2994 3.4105
R3355 VDDA.n3048 VDDA.n2994 3.4105
R3356 VDDA.n3010 VDDA.n2994 3.4105
R3357 VDDA.n3050 VDDA.n2994 3.4105
R3358 VDDA.n3009 VDDA.n2994 3.4105
R3359 VDDA.n2994 VDDA.n16 3.4105
R3360 VDDA.n3052 VDDA.n2994 3.4105
R3361 VDDA.n3023 VDDA.n2951 3.4105
R3362 VDDA.n3022 VDDA.n2951 3.4105
R3363 VDDA.n3026 VDDA.n2951 3.4105
R3364 VDDA.n3021 VDDA.n2951 3.4105
R3365 VDDA.n3028 VDDA.n2951 3.4105
R3366 VDDA.n3020 VDDA.n2951 3.4105
R3367 VDDA.n3030 VDDA.n2951 3.4105
R3368 VDDA.n3019 VDDA.n2951 3.4105
R3369 VDDA.n3032 VDDA.n2951 3.4105
R3370 VDDA.n3018 VDDA.n2951 3.4105
R3371 VDDA.n3034 VDDA.n2951 3.4105
R3372 VDDA.n3017 VDDA.n2951 3.4105
R3373 VDDA.n3036 VDDA.n2951 3.4105
R3374 VDDA.n3016 VDDA.n2951 3.4105
R3375 VDDA.n3038 VDDA.n2951 3.4105
R3376 VDDA.n3015 VDDA.n2951 3.4105
R3377 VDDA.n3040 VDDA.n2951 3.4105
R3378 VDDA.n3014 VDDA.n2951 3.4105
R3379 VDDA.n3042 VDDA.n2951 3.4105
R3380 VDDA.n3013 VDDA.n2951 3.4105
R3381 VDDA.n3044 VDDA.n2951 3.4105
R3382 VDDA.n3012 VDDA.n2951 3.4105
R3383 VDDA.n3046 VDDA.n2951 3.4105
R3384 VDDA.n3011 VDDA.n2951 3.4105
R3385 VDDA.n3048 VDDA.n2951 3.4105
R3386 VDDA.n3010 VDDA.n2951 3.4105
R3387 VDDA.n3050 VDDA.n2951 3.4105
R3388 VDDA.n3009 VDDA.n2951 3.4105
R3389 VDDA.n2951 VDDA.n16 3.4105
R3390 VDDA.n3052 VDDA.n2951 3.4105
R3391 VDDA.n3023 VDDA.n2997 3.4105
R3392 VDDA.n3022 VDDA.n2997 3.4105
R3393 VDDA.n3026 VDDA.n2997 3.4105
R3394 VDDA.n3021 VDDA.n2997 3.4105
R3395 VDDA.n3028 VDDA.n2997 3.4105
R3396 VDDA.n3020 VDDA.n2997 3.4105
R3397 VDDA.n3030 VDDA.n2997 3.4105
R3398 VDDA.n3019 VDDA.n2997 3.4105
R3399 VDDA.n3032 VDDA.n2997 3.4105
R3400 VDDA.n3018 VDDA.n2997 3.4105
R3401 VDDA.n3034 VDDA.n2997 3.4105
R3402 VDDA.n3017 VDDA.n2997 3.4105
R3403 VDDA.n3036 VDDA.n2997 3.4105
R3404 VDDA.n3016 VDDA.n2997 3.4105
R3405 VDDA.n3038 VDDA.n2997 3.4105
R3406 VDDA.n3015 VDDA.n2997 3.4105
R3407 VDDA.n3040 VDDA.n2997 3.4105
R3408 VDDA.n3014 VDDA.n2997 3.4105
R3409 VDDA.n3042 VDDA.n2997 3.4105
R3410 VDDA.n3013 VDDA.n2997 3.4105
R3411 VDDA.n3044 VDDA.n2997 3.4105
R3412 VDDA.n3012 VDDA.n2997 3.4105
R3413 VDDA.n3046 VDDA.n2997 3.4105
R3414 VDDA.n3011 VDDA.n2997 3.4105
R3415 VDDA.n3048 VDDA.n2997 3.4105
R3416 VDDA.n3010 VDDA.n2997 3.4105
R3417 VDDA.n3050 VDDA.n2997 3.4105
R3418 VDDA.n3009 VDDA.n2997 3.4105
R3419 VDDA.n2997 VDDA.n16 3.4105
R3420 VDDA.n3052 VDDA.n2997 3.4105
R3421 VDDA.n3023 VDDA.n2950 3.4105
R3422 VDDA.n3022 VDDA.n2950 3.4105
R3423 VDDA.n3026 VDDA.n2950 3.4105
R3424 VDDA.n3021 VDDA.n2950 3.4105
R3425 VDDA.n3028 VDDA.n2950 3.4105
R3426 VDDA.n3020 VDDA.n2950 3.4105
R3427 VDDA.n3030 VDDA.n2950 3.4105
R3428 VDDA.n3019 VDDA.n2950 3.4105
R3429 VDDA.n3032 VDDA.n2950 3.4105
R3430 VDDA.n3018 VDDA.n2950 3.4105
R3431 VDDA.n3034 VDDA.n2950 3.4105
R3432 VDDA.n3017 VDDA.n2950 3.4105
R3433 VDDA.n3036 VDDA.n2950 3.4105
R3434 VDDA.n3016 VDDA.n2950 3.4105
R3435 VDDA.n3038 VDDA.n2950 3.4105
R3436 VDDA.n3015 VDDA.n2950 3.4105
R3437 VDDA.n3040 VDDA.n2950 3.4105
R3438 VDDA.n3014 VDDA.n2950 3.4105
R3439 VDDA.n3042 VDDA.n2950 3.4105
R3440 VDDA.n3013 VDDA.n2950 3.4105
R3441 VDDA.n3044 VDDA.n2950 3.4105
R3442 VDDA.n3012 VDDA.n2950 3.4105
R3443 VDDA.n3046 VDDA.n2950 3.4105
R3444 VDDA.n3011 VDDA.n2950 3.4105
R3445 VDDA.n3048 VDDA.n2950 3.4105
R3446 VDDA.n3010 VDDA.n2950 3.4105
R3447 VDDA.n3050 VDDA.n2950 3.4105
R3448 VDDA.n3009 VDDA.n2950 3.4105
R3449 VDDA.n2950 VDDA.n16 3.4105
R3450 VDDA.n3052 VDDA.n2950 3.4105
R3451 VDDA.n3023 VDDA.n3000 3.4105
R3452 VDDA.n3022 VDDA.n3000 3.4105
R3453 VDDA.n3026 VDDA.n3000 3.4105
R3454 VDDA.n3021 VDDA.n3000 3.4105
R3455 VDDA.n3028 VDDA.n3000 3.4105
R3456 VDDA.n3020 VDDA.n3000 3.4105
R3457 VDDA.n3030 VDDA.n3000 3.4105
R3458 VDDA.n3019 VDDA.n3000 3.4105
R3459 VDDA.n3032 VDDA.n3000 3.4105
R3460 VDDA.n3018 VDDA.n3000 3.4105
R3461 VDDA.n3034 VDDA.n3000 3.4105
R3462 VDDA.n3017 VDDA.n3000 3.4105
R3463 VDDA.n3036 VDDA.n3000 3.4105
R3464 VDDA.n3016 VDDA.n3000 3.4105
R3465 VDDA.n3038 VDDA.n3000 3.4105
R3466 VDDA.n3015 VDDA.n3000 3.4105
R3467 VDDA.n3040 VDDA.n3000 3.4105
R3468 VDDA.n3014 VDDA.n3000 3.4105
R3469 VDDA.n3042 VDDA.n3000 3.4105
R3470 VDDA.n3013 VDDA.n3000 3.4105
R3471 VDDA.n3044 VDDA.n3000 3.4105
R3472 VDDA.n3012 VDDA.n3000 3.4105
R3473 VDDA.n3046 VDDA.n3000 3.4105
R3474 VDDA.n3011 VDDA.n3000 3.4105
R3475 VDDA.n3048 VDDA.n3000 3.4105
R3476 VDDA.n3010 VDDA.n3000 3.4105
R3477 VDDA.n3050 VDDA.n3000 3.4105
R3478 VDDA.n3009 VDDA.n3000 3.4105
R3479 VDDA.n3000 VDDA.n16 3.4105
R3480 VDDA.n3052 VDDA.n3000 3.4105
R3481 VDDA.n3023 VDDA.n2949 3.4105
R3482 VDDA.n3022 VDDA.n2949 3.4105
R3483 VDDA.n3026 VDDA.n2949 3.4105
R3484 VDDA.n3021 VDDA.n2949 3.4105
R3485 VDDA.n3028 VDDA.n2949 3.4105
R3486 VDDA.n3020 VDDA.n2949 3.4105
R3487 VDDA.n3030 VDDA.n2949 3.4105
R3488 VDDA.n3019 VDDA.n2949 3.4105
R3489 VDDA.n3032 VDDA.n2949 3.4105
R3490 VDDA.n3018 VDDA.n2949 3.4105
R3491 VDDA.n3034 VDDA.n2949 3.4105
R3492 VDDA.n3017 VDDA.n2949 3.4105
R3493 VDDA.n3036 VDDA.n2949 3.4105
R3494 VDDA.n3016 VDDA.n2949 3.4105
R3495 VDDA.n3038 VDDA.n2949 3.4105
R3496 VDDA.n3015 VDDA.n2949 3.4105
R3497 VDDA.n3040 VDDA.n2949 3.4105
R3498 VDDA.n3014 VDDA.n2949 3.4105
R3499 VDDA.n3042 VDDA.n2949 3.4105
R3500 VDDA.n3013 VDDA.n2949 3.4105
R3501 VDDA.n3044 VDDA.n2949 3.4105
R3502 VDDA.n3012 VDDA.n2949 3.4105
R3503 VDDA.n3046 VDDA.n2949 3.4105
R3504 VDDA.n3011 VDDA.n2949 3.4105
R3505 VDDA.n3048 VDDA.n2949 3.4105
R3506 VDDA.n3010 VDDA.n2949 3.4105
R3507 VDDA.n3050 VDDA.n2949 3.4105
R3508 VDDA.n3009 VDDA.n2949 3.4105
R3509 VDDA.n2949 VDDA.n16 3.4105
R3510 VDDA.n3052 VDDA.n2949 3.4105
R3511 VDDA.n3023 VDDA.n3003 3.4105
R3512 VDDA.n3022 VDDA.n3003 3.4105
R3513 VDDA.n3026 VDDA.n3003 3.4105
R3514 VDDA.n3021 VDDA.n3003 3.4105
R3515 VDDA.n3028 VDDA.n3003 3.4105
R3516 VDDA.n3020 VDDA.n3003 3.4105
R3517 VDDA.n3030 VDDA.n3003 3.4105
R3518 VDDA.n3019 VDDA.n3003 3.4105
R3519 VDDA.n3032 VDDA.n3003 3.4105
R3520 VDDA.n3018 VDDA.n3003 3.4105
R3521 VDDA.n3034 VDDA.n3003 3.4105
R3522 VDDA.n3017 VDDA.n3003 3.4105
R3523 VDDA.n3036 VDDA.n3003 3.4105
R3524 VDDA.n3016 VDDA.n3003 3.4105
R3525 VDDA.n3038 VDDA.n3003 3.4105
R3526 VDDA.n3015 VDDA.n3003 3.4105
R3527 VDDA.n3040 VDDA.n3003 3.4105
R3528 VDDA.n3014 VDDA.n3003 3.4105
R3529 VDDA.n3042 VDDA.n3003 3.4105
R3530 VDDA.n3013 VDDA.n3003 3.4105
R3531 VDDA.n3044 VDDA.n3003 3.4105
R3532 VDDA.n3012 VDDA.n3003 3.4105
R3533 VDDA.n3046 VDDA.n3003 3.4105
R3534 VDDA.n3011 VDDA.n3003 3.4105
R3535 VDDA.n3048 VDDA.n3003 3.4105
R3536 VDDA.n3010 VDDA.n3003 3.4105
R3537 VDDA.n3050 VDDA.n3003 3.4105
R3538 VDDA.n3009 VDDA.n3003 3.4105
R3539 VDDA.n3003 VDDA.n16 3.4105
R3540 VDDA.n3052 VDDA.n3003 3.4105
R3541 VDDA.n3023 VDDA.n2948 3.4105
R3542 VDDA.n3022 VDDA.n2948 3.4105
R3543 VDDA.n3026 VDDA.n2948 3.4105
R3544 VDDA.n3021 VDDA.n2948 3.4105
R3545 VDDA.n3028 VDDA.n2948 3.4105
R3546 VDDA.n3020 VDDA.n2948 3.4105
R3547 VDDA.n3030 VDDA.n2948 3.4105
R3548 VDDA.n3019 VDDA.n2948 3.4105
R3549 VDDA.n3032 VDDA.n2948 3.4105
R3550 VDDA.n3018 VDDA.n2948 3.4105
R3551 VDDA.n3034 VDDA.n2948 3.4105
R3552 VDDA.n3017 VDDA.n2948 3.4105
R3553 VDDA.n3036 VDDA.n2948 3.4105
R3554 VDDA.n3016 VDDA.n2948 3.4105
R3555 VDDA.n3038 VDDA.n2948 3.4105
R3556 VDDA.n3015 VDDA.n2948 3.4105
R3557 VDDA.n3040 VDDA.n2948 3.4105
R3558 VDDA.n3014 VDDA.n2948 3.4105
R3559 VDDA.n3042 VDDA.n2948 3.4105
R3560 VDDA.n3013 VDDA.n2948 3.4105
R3561 VDDA.n3044 VDDA.n2948 3.4105
R3562 VDDA.n3012 VDDA.n2948 3.4105
R3563 VDDA.n3046 VDDA.n2948 3.4105
R3564 VDDA.n3011 VDDA.n2948 3.4105
R3565 VDDA.n3048 VDDA.n2948 3.4105
R3566 VDDA.n3010 VDDA.n2948 3.4105
R3567 VDDA.n3050 VDDA.n2948 3.4105
R3568 VDDA.n3009 VDDA.n2948 3.4105
R3569 VDDA.n2948 VDDA.n16 3.4105
R3570 VDDA.n3052 VDDA.n2948 3.4105
R3571 VDDA.n3023 VDDA.n3006 3.4105
R3572 VDDA.n3022 VDDA.n3006 3.4105
R3573 VDDA.n3026 VDDA.n3006 3.4105
R3574 VDDA.n3021 VDDA.n3006 3.4105
R3575 VDDA.n3028 VDDA.n3006 3.4105
R3576 VDDA.n3020 VDDA.n3006 3.4105
R3577 VDDA.n3030 VDDA.n3006 3.4105
R3578 VDDA.n3019 VDDA.n3006 3.4105
R3579 VDDA.n3032 VDDA.n3006 3.4105
R3580 VDDA.n3018 VDDA.n3006 3.4105
R3581 VDDA.n3034 VDDA.n3006 3.4105
R3582 VDDA.n3017 VDDA.n3006 3.4105
R3583 VDDA.n3036 VDDA.n3006 3.4105
R3584 VDDA.n3016 VDDA.n3006 3.4105
R3585 VDDA.n3038 VDDA.n3006 3.4105
R3586 VDDA.n3015 VDDA.n3006 3.4105
R3587 VDDA.n3040 VDDA.n3006 3.4105
R3588 VDDA.n3014 VDDA.n3006 3.4105
R3589 VDDA.n3042 VDDA.n3006 3.4105
R3590 VDDA.n3013 VDDA.n3006 3.4105
R3591 VDDA.n3044 VDDA.n3006 3.4105
R3592 VDDA.n3012 VDDA.n3006 3.4105
R3593 VDDA.n3046 VDDA.n3006 3.4105
R3594 VDDA.n3011 VDDA.n3006 3.4105
R3595 VDDA.n3048 VDDA.n3006 3.4105
R3596 VDDA.n3010 VDDA.n3006 3.4105
R3597 VDDA.n3050 VDDA.n3006 3.4105
R3598 VDDA.n3009 VDDA.n3006 3.4105
R3599 VDDA.n3006 VDDA.n16 3.4105
R3600 VDDA.n3052 VDDA.n3006 3.4105
R3601 VDDA.n3023 VDDA.n2947 3.4105
R3602 VDDA.n3022 VDDA.n2947 3.4105
R3603 VDDA.n3026 VDDA.n2947 3.4105
R3604 VDDA.n3021 VDDA.n2947 3.4105
R3605 VDDA.n3028 VDDA.n2947 3.4105
R3606 VDDA.n3020 VDDA.n2947 3.4105
R3607 VDDA.n3030 VDDA.n2947 3.4105
R3608 VDDA.n3019 VDDA.n2947 3.4105
R3609 VDDA.n3032 VDDA.n2947 3.4105
R3610 VDDA.n3018 VDDA.n2947 3.4105
R3611 VDDA.n3034 VDDA.n2947 3.4105
R3612 VDDA.n3017 VDDA.n2947 3.4105
R3613 VDDA.n3036 VDDA.n2947 3.4105
R3614 VDDA.n3016 VDDA.n2947 3.4105
R3615 VDDA.n3038 VDDA.n2947 3.4105
R3616 VDDA.n3015 VDDA.n2947 3.4105
R3617 VDDA.n3040 VDDA.n2947 3.4105
R3618 VDDA.n3014 VDDA.n2947 3.4105
R3619 VDDA.n3042 VDDA.n2947 3.4105
R3620 VDDA.n3013 VDDA.n2947 3.4105
R3621 VDDA.n3044 VDDA.n2947 3.4105
R3622 VDDA.n3012 VDDA.n2947 3.4105
R3623 VDDA.n3046 VDDA.n2947 3.4105
R3624 VDDA.n3011 VDDA.n2947 3.4105
R3625 VDDA.n3048 VDDA.n2947 3.4105
R3626 VDDA.n3010 VDDA.n2947 3.4105
R3627 VDDA.n3050 VDDA.n2947 3.4105
R3628 VDDA.n3009 VDDA.n2947 3.4105
R3629 VDDA.n2947 VDDA.n16 3.4105
R3630 VDDA.n3052 VDDA.n2947 3.4105
R3631 VDDA.n3051 VDDA.n3022 3.4105
R3632 VDDA.n3051 VDDA.n3026 3.4105
R3633 VDDA.n3051 VDDA.n3021 3.4105
R3634 VDDA.n3051 VDDA.n3028 3.4105
R3635 VDDA.n3051 VDDA.n3020 3.4105
R3636 VDDA.n3051 VDDA.n3030 3.4105
R3637 VDDA.n3051 VDDA.n3019 3.4105
R3638 VDDA.n3051 VDDA.n3032 3.4105
R3639 VDDA.n3051 VDDA.n3018 3.4105
R3640 VDDA.n3051 VDDA.n3034 3.4105
R3641 VDDA.n3051 VDDA.n3017 3.4105
R3642 VDDA.n3051 VDDA.n3036 3.4105
R3643 VDDA.n3051 VDDA.n3016 3.4105
R3644 VDDA.n3051 VDDA.n3038 3.4105
R3645 VDDA.n3051 VDDA.n3015 3.4105
R3646 VDDA.n3051 VDDA.n3040 3.4105
R3647 VDDA.n3051 VDDA.n3014 3.4105
R3648 VDDA.n3051 VDDA.n3042 3.4105
R3649 VDDA.n3051 VDDA.n3013 3.4105
R3650 VDDA.n3051 VDDA.n3044 3.4105
R3651 VDDA.n3051 VDDA.n3012 3.4105
R3652 VDDA.n3051 VDDA.n3046 3.4105
R3653 VDDA.n3051 VDDA.n3011 3.4105
R3654 VDDA.n3051 VDDA.n3048 3.4105
R3655 VDDA.n3051 VDDA.n3010 3.4105
R3656 VDDA.n3051 VDDA.n3050 3.4105
R3657 VDDA.n3051 VDDA.n3009 3.4105
R3658 VDDA.n3051 VDDA.n16 3.4105
R3659 VDDA.n3052 VDDA.n3051 3.4105
R3660 VDDA.n384 VDDA.n383 3.06776
R3661 VDDA.n2329 VDDA.n2325 2.96402
R3662 VDDA.n434 VDDA.n430 2.96402
R3663 VDDA.n2366 VDDA.n2365 2.8957
R3664 VDDA.n2367 VDDA.n2366 2.8957
R3665 VDDA.n2371 VDDA.n2369 2.8957
R3666 VDDA.n2374 VDDA.n2369 2.8957
R3667 VDDA.n2370 VDDA.n2367 2.8957
R3668 VDDA.n2374 VDDA.n2373 2.8957
R3669 VDDA.n2376 VDDA.n2365 2.8957
R3670 VDDA.n2371 VDDA.n2370 2.8957
R3671 VDDA.n372 VDDA.n371 2.8255
R3672 VDDA.n374 VDDA.n373 2.8255
R3673 VDDA.n2328 VDDA.n2327 2.423
R3674 VDDA.n2326 VDDA.n2325 2.423
R3675 VDDA.n431 VDDA.n430 2.423
R3676 VDDA.n433 VDDA.n432 2.423
R3677 VDDA.n1904 VDDA.n1903 2.41009
R3678 VDDA.n2376 VDDA.n2364 2.32777
R3679 VDDA.n91 VDDA.n90 2.30736
R3680 VDDA.n2815 VDDA.n2812 2.30736
R3681 VDDA.n2665 VDDA.n2664 2.30736
R3682 VDDA.n269 VDDA.n268 2.30736
R3683 VDDA.n2467 VDDA.n2464 2.30736
R3684 VDDA.n1225 VDDA.n1224 2.30736
R3685 VDDA.n535 VDDA.n534 2.30736
R3686 VDDA.n1027 VDDA.n1024 2.30736
R3687 VDDA.n877 VDDA.n876 2.30736
R3688 VDDA.n1576 VDDA.n1575 2.30736
R3689 VDDA.n2251 VDDA.n2250 2.30736
R3690 VDDA.n689 VDDA.n688 2.30736
R3691 VDDA.n2329 VDDA.n2328 2.27652
R3692 VDDA.n434 VDDA.n433 2.27652
R3693 VDDA.n1946 VDDA.n1938 2.26187
R3694 VDDA.n2007 VDDA.n1936 2.26187
R3695 VDDA.n2084 VDDA.n1934 2.26187
R3696 VDDA.n2134 VDDA.n1932 2.26187
R3697 VDDA.n427 VDDA.n405 2.26187
R3698 VDDA.n411 VDDA.n408 2.26187
R3699 VDDA.n412 VDDA.n411 2.26187
R3700 VDDA.n2322 VDDA.n2321 2.26187
R3701 VDDA.n803 VDDA.n800 2.26187
R3702 VDDA.n803 VDDA.n802 2.26187
R3703 VDDA.n1943 VDDA.n1938 2.26187
R3704 VDDA.n2323 VDDA.n2322 2.26187
R3705 VDDA.n2334 VDDA.n2333 2.26187
R3706 VDDA.n2284 VDDA.n2283 2.26187
R3707 VDDA.n1763 VDDA.n1403 2.2505
R3708 VDDA.n1762 VDDA.n1761 2.2505
R3709 VDDA.n1405 VDDA.n1404 2.2505
R3710 VDDA.n1583 VDDA.n1580 2.2505
R3711 VDDA.n1753 VDDA.n1752 2.2505
R3712 VDDA.n1751 VDDA.n1582 2.2505
R3713 VDDA.n1750 VDDA.n1749 2.2505
R3714 VDDA.n1585 VDDA.n1584 2.2505
R3715 VDDA.n1743 VDDA.n1742 2.2505
R3716 VDDA.n1741 VDDA.n1589 2.2505
R3717 VDDA.n1740 VDDA.n1739 2.2505
R3718 VDDA.n1591 VDDA.n1590 2.2505
R3719 VDDA.n1733 VDDA.n1732 2.2505
R3720 VDDA.n1731 VDDA.n1595 2.2505
R3721 VDDA.n1730 VDDA.n1729 2.2505
R3722 VDDA.n1597 VDDA.n1596 2.2505
R3723 VDDA.n1723 VDDA.n1722 2.2505
R3724 VDDA.n1721 VDDA.n1601 2.2505
R3725 VDDA.n1720 VDDA.n1719 2.2505
R3726 VDDA.n1603 VDDA.n1602 2.2505
R3727 VDDA.n1713 VDDA.n1712 2.2505
R3728 VDDA.n1711 VDDA.n1607 2.2505
R3729 VDDA.n1710 VDDA.n1709 2.2505
R3730 VDDA.n1609 VDDA.n1608 2.2505
R3731 VDDA.n1703 VDDA.n1702 2.2505
R3732 VDDA.n1701 VDDA.n1613 2.2505
R3733 VDDA.n1700 VDDA.n1699 2.2505
R3734 VDDA.n1615 VDDA.n1614 2.2505
R3735 VDDA.n1693 VDDA.n1692 2.2505
R3736 VDDA.n1691 VDDA.n1619 2.2505
R3737 VDDA.n1690 VDDA.n1689 2.2505
R3738 VDDA.n1621 VDDA.n1620 2.2505
R3739 VDDA.n1683 VDDA.n1682 2.2505
R3740 VDDA.n1681 VDDA.n1625 2.2505
R3741 VDDA.n1680 VDDA.n1679 2.2505
R3742 VDDA.n1627 VDDA.n1626 2.2505
R3743 VDDA.n1673 VDDA.n1672 2.2505
R3744 VDDA.n1671 VDDA.n1631 2.2505
R3745 VDDA.n1670 VDDA.n1669 2.2505
R3746 VDDA.n1633 VDDA.n1632 2.2505
R3747 VDDA.n1663 VDDA.n1662 2.2505
R3748 VDDA.n1661 VDDA.n1637 2.2505
R3749 VDDA.n1660 VDDA.n1659 2.2505
R3750 VDDA.n1639 VDDA.n1638 2.2505
R3751 VDDA.n1653 VDDA.n1652 2.2505
R3752 VDDA.n1651 VDDA.n1643 2.2505
R3753 VDDA.n1947 VDDA.n1937 2.24063
R3754 VDDA.n2008 VDDA.n1935 2.24063
R3755 VDDA.n2085 VDDA.n1933 2.24063
R3756 VDDA.n2135 VDDA.n1931 2.24063
R3757 VDDA.n429 VDDA.n428 2.24063
R3758 VDDA.n2394 VDDA.n2393 2.24063
R3759 VDDA.n404 VDDA.n388 2.24063
R3760 VDDA.n2338 VDDA.n2337 2.24063
R3761 VDDA.n2336 VDDA.n447 2.24063
R3762 VDDA.n2331 VDDA.n2330 2.24063
R3763 VDDA.n2333 VDDA.n2332 2.24063
R3764 VDDA.n2321 VDDA.n2320 2.24063
R3765 VDDA.n978 VDDA.n631 2.24063
R3766 VDDA.n632 VDDA.n630 2.24063
R3767 VDDA.n1149 VDDA.n628 2.24063
R3768 VDDA.n629 VDDA.n627 2.24063
R3769 VDDA.n1153 VDDA.n456 2.24063
R3770 VDDA.n626 VDDA.n625 2.24063
R3771 VDDA.n2283 VDDA.n450 2.24063
R3772 VDDA.n2282 VDDA.n449 2.24063
R3773 VDDA.n2400 VDDA.n367 2.24063
R3774 VDDA.n368 VDDA.n366 2.24063
R3775 VDDA.n2397 VDDA.n2396 2.24063
R3776 VDDA.n2262 VDDA.n454 2.24063
R3777 VDDA.n455 VDDA.n453 2.24063
R3778 VDDA.n2589 VDDA.n362 2.24063
R3779 VDDA.n363 VDDA.n361 2.24063
R3780 VDDA.n2593 VDDA.n190 2.24063
R3781 VDDA.n360 VDDA.n359 2.24063
R3782 VDDA.n2766 VDDA.n188 2.24063
R3783 VDDA.n189 VDDA.n187 2.24063
R3784 VDDA.n2937 VDDA.n185 2.24063
R3785 VDDA.n186 VDDA.n184 2.24063
R3786 VDDA.n2941 VDDA.n2940 2.24063
R3787 VDDA.n183 VDDA.n182 2.24063
R3788 VDDA.n1943 VDDA.n1942 2.24063
R3789 VDDA.n1948 VDDA.n1936 2.24063
R3790 VDDA.n2004 VDDA.n2003 2.24063
R3791 VDDA.n2009 VDDA.n1934 2.24063
R3792 VDDA.n2081 VDDA.n2080 2.24063
R3793 VDDA.n2086 VDDA.n1932 2.24063
R3794 VDDA.n2131 VDDA.n2130 2.24063
R3795 VDDA.n437 VDDA.n405 2.24063
R3796 VDDA.n436 VDDA.n435 2.24063
R3797 VDDA.n426 VDDA.n408 2.24063
R3798 VDDA.n425 VDDA.n424 2.24063
R3799 VDDA.n2395 VDDA.n386 2.24063
R3800 VDDA.n2340 VDDA.n2339 2.24063
R3801 VDDA.n2342 VDDA.n2341 2.24063
R3802 VDDA.n2335 VDDA.n2303 2.24063
R3803 VDDA.n2324 VDDA.n2306 2.24063
R3804 VDDA.n975 VDDA.n974 2.24063
R3805 VDDA.n1146 VDDA.n1145 2.24063
R3806 VDDA.n1154 VDDA.n624 2.24063
R3807 VDDA.n2259 VDDA.n2258 2.24063
R3808 VDDA.n2586 VDDA.n2585 2.24063
R3809 VDDA.n2594 VDDA.n358 2.24063
R3810 VDDA.n2763 VDDA.n2762 2.24063
R3811 VDDA.n2934 VDDA.n2933 2.24063
R3812 VDDA.n2942 VDDA.n180 2.24063
R3813 VDDA.n806 VDDA.n800 2.24063
R3814 VDDA.n805 VDDA.n633 2.24063
R3815 VDDA.n2943 VDDA.n2942 2.16196
R3816 VDDA.n2933 VDDA.n2932 2.16196
R3817 VDDA.n2762 VDDA.n2761 2.16196
R3818 VDDA.n2595 VDDA.n2594 2.16196
R3819 VDDA.n2585 VDDA.n2584 2.16196
R3820 VDDA.n2258 VDDA.n2257 2.16196
R3821 VDDA.n1155 VDDA.n1154 2.16196
R3822 VDDA.n1145 VDDA.n1144 2.16196
R3823 VDDA.n974 VDDA.n973 2.16196
R3824 VDDA.n807 VDDA.n806 2.16196
R3825 VDDA.n2411 VDDA.n364 2.16194
R3826 VDDA.n2418 VDDA.n2417 2.16194
R3827 VDDA.n2405 VDDA.n2401 2.16194
R3828 VDDA.n2273 VDDA.n451 2.16194
R3829 VDDA.n2280 VDDA.n2279 2.16194
R3830 VDDA.n2267 VDDA.n2263 2.16194
R3831 VDDA.n383 VDDA.n382 2.12369
R3832 VDDA.n1789 VDDA.n1788 2.05049
R3833 VDDA.n1764 VDDA.n1402 1.9823
R3834 VDDA.n1765 VDDA.n1764 1.9823
R3835 VDDA.n400 VDDA.n399 1.97758
R3836 VDDA.n402 VDDA.n401 1.97758
R3837 VDDA.n2301 VDDA.n2300 1.97758
R3838 VDDA.n2299 VDDA.n2298 1.97758
R3839 VDDA.n399 VDDA.n398 1.95361
R3840 VDDA.n2298 VDDA.n2297 1.95361
R3841 VDDA.n381 VDDA.n380 1.888
R3842 VDDA.n379 VDDA.n378 1.888
R3843 VDDA.n403 VDDA.n402 1.83902
R3844 VDDA.n2302 VDDA.n2301 1.83902
R3845 VDDA.n1650 VDDA.n1644 1.74133
R3846 VDDA.n2962 VDDA.n0 1.70567
R3847 VDDA.n2965 VDDA.n2962 1.70567
R3848 VDDA.n2968 VDDA.n2962 1.70567
R3849 VDDA.n2971 VDDA.n2962 1.70567
R3850 VDDA.n2974 VDDA.n2962 1.70567
R3851 VDDA.n2977 VDDA.n2962 1.70567
R3852 VDDA.n2980 VDDA.n2962 1.70567
R3853 VDDA.n2983 VDDA.n2962 1.70567
R3854 VDDA.n2986 VDDA.n2962 1.70567
R3855 VDDA.n2989 VDDA.n2962 1.70567
R3856 VDDA.n2992 VDDA.n2962 1.70567
R3857 VDDA.n2995 VDDA.n2962 1.70567
R3858 VDDA.n2998 VDDA.n2962 1.70567
R3859 VDDA.n3001 VDDA.n2962 1.70567
R3860 VDDA.n3004 VDDA.n2962 1.70567
R3861 VDDA.n3007 VDDA.n2962 1.70567
R3862 VDDA.n3053 VDDA.n14 1.70565
R3863 VDDA.n3053 VDDA.n12 1.70565
R3864 VDDA.n3053 VDDA.n10 1.70565
R3865 VDDA.n3053 VDDA.n8 1.70565
R3866 VDDA.n3053 VDDA.n6 1.70565
R3867 VDDA.n3053 VDDA.n4 1.70565
R3868 VDDA.n3053 VDDA.n2 1.70565
R3869 VDDA.n3029 VDDA.n2964 1.70565
R3870 VDDA.n3031 VDDA.n2964 1.70565
R3871 VDDA.n3037 VDDA.n2964 1.70565
R3872 VDDA.n3039 VDDA.n2964 1.70565
R3873 VDDA.n3045 VDDA.n2964 1.70565
R3874 VDDA.n3047 VDDA.n2964 1.70565
R3875 VDDA.n3051 VDDA.n3024 1.70565
R3876 VDDA.n3053 VDDA.n13 1.70563
R3877 VDDA.n3053 VDDA.n9 1.70563
R3878 VDDA.n3053 VDDA.n5 1.70563
R3879 VDDA.n3053 VDDA.n1 1.70563
R3880 VDDA.n3025 VDDA.n2964 1.70563
R3881 VDDA.n3027 VDDA.n2964 1.70563
R3882 VDDA.n3033 VDDA.n2964 1.70563
R3883 VDDA.n3035 VDDA.n2964 1.70563
R3884 VDDA.n3041 VDDA.n2964 1.70563
R3885 VDDA.n3043 VDDA.n2964 1.70563
R3886 VDDA.n3049 VDDA.n2964 1.70563
R3887 VDDA.n3008 VDDA.n2964 1.70563
R3888 VDDA.n2963 VDDA.n15 1.70563
R3889 VDDA.n2969 VDDA.n15 1.70563
R3890 VDDA.n2975 VDDA.n15 1.70563
R3891 VDDA.n2981 VDDA.n15 1.70563
R3892 VDDA.n2987 VDDA.n15 1.70563
R3893 VDDA.n2993 VDDA.n15 1.70563
R3894 VDDA.n2999 VDDA.n15 1.70563
R3895 VDDA.n3005 VDDA.n15 1.70563
R3896 VDDA.n3053 VDDA.n11 1.70556
R3897 VDDA.n3053 VDDA.n7 1.70556
R3898 VDDA.n3053 VDDA.n3 1.70556
R3899 VDDA.n2966 VDDA.n15 1.70556
R3900 VDDA.n2972 VDDA.n15 1.70556
R3901 VDDA.n2978 VDDA.n15 1.70556
R3902 VDDA.n2984 VDDA.n15 1.70556
R3903 VDDA.n2990 VDDA.n15 1.70556
R3904 VDDA.n2996 VDDA.n15 1.70556
R3905 VDDA.n3002 VDDA.n15 1.70556
R3906 VDDA.n1649 VDDA.n1648 1.7055
R3907 VDDA.n1645 VDDA.n1643 1.7055
R3908 VDDA.n1654 VDDA.n1653 1.7055
R3909 VDDA.n1656 VDDA.n1639 1.7055
R3910 VDDA.n1659 VDDA.n1658 1.7055
R3911 VDDA.n1640 VDDA.n1637 1.7055
R3912 VDDA.n1664 VDDA.n1663 1.7055
R3913 VDDA.n1666 VDDA.n1633 1.7055
R3914 VDDA.n1669 VDDA.n1668 1.7055
R3915 VDDA.n1634 VDDA.n1631 1.7055
R3916 VDDA.n1674 VDDA.n1673 1.7055
R3917 VDDA.n1676 VDDA.n1627 1.7055
R3918 VDDA.n1679 VDDA.n1678 1.7055
R3919 VDDA.n1628 VDDA.n1625 1.7055
R3920 VDDA.n1684 VDDA.n1683 1.7055
R3921 VDDA.n1686 VDDA.n1621 1.7055
R3922 VDDA.n1689 VDDA.n1688 1.7055
R3923 VDDA.n1622 VDDA.n1619 1.7055
R3924 VDDA.n1694 VDDA.n1693 1.7055
R3925 VDDA.n1696 VDDA.n1615 1.7055
R3926 VDDA.n1699 VDDA.n1698 1.7055
R3927 VDDA.n1616 VDDA.n1613 1.7055
R3928 VDDA.n1704 VDDA.n1703 1.7055
R3929 VDDA.n1706 VDDA.n1609 1.7055
R3930 VDDA.n1709 VDDA.n1708 1.7055
R3931 VDDA.n1610 VDDA.n1607 1.7055
R3932 VDDA.n1714 VDDA.n1713 1.7055
R3933 VDDA.n1716 VDDA.n1603 1.7055
R3934 VDDA.n1719 VDDA.n1718 1.7055
R3935 VDDA.n1604 VDDA.n1601 1.7055
R3936 VDDA.n1724 VDDA.n1723 1.7055
R3937 VDDA.n1726 VDDA.n1597 1.7055
R3938 VDDA.n1729 VDDA.n1728 1.7055
R3939 VDDA.n1598 VDDA.n1595 1.7055
R3940 VDDA.n1734 VDDA.n1733 1.7055
R3941 VDDA.n1736 VDDA.n1591 1.7055
R3942 VDDA.n1739 VDDA.n1738 1.7055
R3943 VDDA.n1592 VDDA.n1589 1.7055
R3944 VDDA.n1744 VDDA.n1743 1.7055
R3945 VDDA.n1746 VDDA.n1585 1.7055
R3946 VDDA.n1749 VDDA.n1748 1.7055
R3947 VDDA.n1586 VDDA.n1582 1.7055
R3948 VDDA.n1754 VDDA.n1753 1.7055
R3949 VDDA.n1756 VDDA.n1580 1.7055
R3950 VDDA.n1758 VDDA.n1405 1.7055
R3951 VDDA.n1761 VDDA.n1760 1.7055
R3952 VDDA.n1407 VDDA.n1403 1.7055
R3953 VDDA.n1641 VDDA.n1579 1.69989
R3954 VDDA.n1675 VDDA.n1579 1.69989
R3955 VDDA.n1623 VDDA.n1579 1.69989
R3956 VDDA.n1705 VDDA.n1579 1.69989
R3957 VDDA.n1605 VDDA.n1579 1.69989
R3958 VDDA.n1735 VDDA.n1579 1.69989
R3959 VDDA.n1587 VDDA.n1579 1.69989
R3960 VDDA.n1657 VDDA.n1366 1.69938
R3961 VDDA.n1636 VDDA.n1366 1.69938
R3962 VDDA.n1630 VDDA.n1366 1.69938
R3963 VDDA.n1677 VDDA.n1366 1.69938
R3964 VDDA.n1687 VDDA.n1366 1.69938
R3965 VDDA.n1618 VDDA.n1366 1.69938
R3966 VDDA.n1612 VDDA.n1366 1.69938
R3967 VDDA.n1707 VDDA.n1366 1.69938
R3968 VDDA.n1717 VDDA.n1366 1.69938
R3969 VDDA.n1600 VDDA.n1366 1.69938
R3970 VDDA.n1594 VDDA.n1366 1.69938
R3971 VDDA.n1737 VDDA.n1366 1.69938
R3972 VDDA.n1747 VDDA.n1366 1.69938
R3973 VDDA.n1581 VDDA.n1366 1.69938
R3974 VDDA.n1406 VDDA.n1366 1.69938
R3975 VDDA.n1647 VDDA.n1366 1.69938
R3976 VDDA.n1646 VDDA.n1579 1.69888
R3977 VDDA.n1642 VDDA.n1366 1.69888
R3978 VDDA.n1655 VDDA.n1579 1.69888
R3979 VDDA.n1665 VDDA.n1579 1.69888
R3980 VDDA.n1667 VDDA.n1366 1.69888
R3981 VDDA.n1635 VDDA.n1579 1.69888
R3982 VDDA.n1629 VDDA.n1579 1.69888
R3983 VDDA.n1624 VDDA.n1366 1.69888
R3984 VDDA.n1685 VDDA.n1579 1.69888
R3985 VDDA.n1695 VDDA.n1579 1.69888
R3986 VDDA.n1697 VDDA.n1366 1.69888
R3987 VDDA.n1617 VDDA.n1579 1.69888
R3988 VDDA.n1611 VDDA.n1579 1.69888
R3989 VDDA.n1606 VDDA.n1366 1.69888
R3990 VDDA.n1715 VDDA.n1579 1.69888
R3991 VDDA.n1725 VDDA.n1579 1.69888
R3992 VDDA.n1727 VDDA.n1366 1.69888
R3993 VDDA.n1599 VDDA.n1579 1.69888
R3994 VDDA.n1593 VDDA.n1579 1.69888
R3995 VDDA.n1588 VDDA.n1366 1.69888
R3996 VDDA.n1745 VDDA.n1579 1.69888
R3997 VDDA.n1755 VDDA.n1579 1.69888
R3998 VDDA.n1757 VDDA.n1366 1.69888
R3999 VDDA.n1759 VDDA.n1579 1.69888
R4000 VDDA.n810 VDDA.n659 1.69433
R4001 VDDA.n810 VDDA.n656 1.69433
R4002 VDDA.n810 VDDA.n653 1.69433
R4003 VDDA.n810 VDDA.n650 1.69433
R4004 VDDA.n810 VDDA.n647 1.69433
R4005 VDDA.n810 VDDA.n644 1.69433
R4006 VDDA.n810 VDDA.n641 1.69433
R4007 VDDA.n970 VDDA.n832 1.69433
R4008 VDDA.n970 VDDA.n829 1.69433
R4009 VDDA.n970 VDDA.n826 1.69433
R4010 VDDA.n970 VDDA.n823 1.69433
R4011 VDDA.n970 VDDA.n820 1.69433
R4012 VDDA.n970 VDDA.n817 1.69433
R4013 VDDA.n970 VDDA.n814 1.69433
R4014 VDDA.n1130 VDDA.n461 1.69433
R4015 VDDA.n1112 VDDA.n461 1.69433
R4016 VDDA.n1100 VDDA.n461 1.69433
R4017 VDDA.n1082 VDDA.n461 1.69433
R4018 VDDA.n1070 VDDA.n461 1.69433
R4019 VDDA.n1052 VDDA.n461 1.69433
R4020 VDDA.n1040 VDDA.n461 1.69433
R4021 VDDA.n1158 VDDA.n483 1.69433
R4022 VDDA.n1158 VDDA.n480 1.69433
R4023 VDDA.n1158 VDDA.n477 1.69433
R4024 VDDA.n1158 VDDA.n474 1.69433
R4025 VDDA.n1158 VDDA.n471 1.69433
R4026 VDDA.n1158 VDDA.n468 1.69433
R4027 VDDA.n1158 VDDA.n465 1.69433
R4028 VDDA.n2254 VDDA.n1180 1.69433
R4029 VDDA.n2254 VDDA.n1177 1.69433
R4030 VDDA.n2254 VDDA.n1174 1.69433
R4031 VDDA.n2254 VDDA.n1171 1.69433
R4032 VDDA.n2254 VDDA.n1168 1.69433
R4033 VDDA.n2254 VDDA.n1165 1.69433
R4034 VDDA.n2254 VDDA.n1162 1.69433
R4035 VDDA.n2253 VDDA.n1339 1.69433
R4036 VDDA.n2253 VDDA.n1336 1.69433
R4037 VDDA.n2253 VDDA.n1333 1.69433
R4038 VDDA.n2253 VDDA.n1330 1.69433
R4039 VDDA.n2253 VDDA.n1327 1.69433
R4040 VDDA.n2253 VDDA.n1324 1.69433
R4041 VDDA.n2253 VDDA.n1321 1.69433
R4042 VDDA.n2570 VDDA.n195 1.69433
R4043 VDDA.n2552 VDDA.n195 1.69433
R4044 VDDA.n2540 VDDA.n195 1.69433
R4045 VDDA.n2522 VDDA.n195 1.69433
R4046 VDDA.n2510 VDDA.n195 1.69433
R4047 VDDA.n2492 VDDA.n195 1.69433
R4048 VDDA.n2480 VDDA.n195 1.69433
R4049 VDDA.n2598 VDDA.n217 1.69433
R4050 VDDA.n2598 VDDA.n214 1.69433
R4051 VDDA.n2598 VDDA.n211 1.69433
R4052 VDDA.n2598 VDDA.n208 1.69433
R4053 VDDA.n2598 VDDA.n205 1.69433
R4054 VDDA.n2598 VDDA.n202 1.69433
R4055 VDDA.n2598 VDDA.n199 1.69433
R4056 VDDA.n2758 VDDA.n2620 1.69433
R4057 VDDA.n2758 VDDA.n2617 1.69433
R4058 VDDA.n2758 VDDA.n2614 1.69433
R4059 VDDA.n2758 VDDA.n2611 1.69433
R4060 VDDA.n2758 VDDA.n2608 1.69433
R4061 VDDA.n2758 VDDA.n2605 1.69433
R4062 VDDA.n2758 VDDA.n2602 1.69433
R4063 VDDA.n2918 VDDA.n17 1.69433
R4064 VDDA.n2900 VDDA.n17 1.69433
R4065 VDDA.n2888 VDDA.n17 1.69433
R4066 VDDA.n2870 VDDA.n17 1.69433
R4067 VDDA.n2858 VDDA.n17 1.69433
R4068 VDDA.n2840 VDDA.n17 1.69433
R4069 VDDA.n2828 VDDA.n17 1.69433
R4070 VDDA.n2946 VDDA.n39 1.69433
R4071 VDDA.n2946 VDDA.n36 1.69433
R4072 VDDA.n2946 VDDA.n33 1.69433
R4073 VDDA.n2946 VDDA.n30 1.69433
R4074 VDDA.n2946 VDDA.n27 1.69433
R4075 VDDA.n2946 VDDA.n24 1.69433
R4076 VDDA.n2946 VDDA.n21 1.69433
R4077 VDDA.n1578 VDDA.n1429 1.69433
R4078 VDDA.n1578 VDDA.n1426 1.69433
R4079 VDDA.n1578 VDDA.n1423 1.69433
R4080 VDDA.n1578 VDDA.n1420 1.69433
R4081 VDDA.n1578 VDDA.n1417 1.69433
R4082 VDDA.n1578 VDDA.n1414 1.69433
R4083 VDDA.n1578 VDDA.n1411 1.69433
R4084 VDDA.n1906 VDDA.n1363 1.69328
R4085 VDDA.n1906 VDDA.n1360 1.69328
R4086 VDDA.n1906 VDDA.n1357 1.69328
R4087 VDDA.n1906 VDDA.n1354 1.69328
R4088 VDDA.n1906 VDDA.n1351 1.69328
R4089 VDDA.n1906 VDDA.n1348 1.69328
R4090 VDDA.n1906 VDDA.n1345 1.69328
R4091 VDDA.n810 VDDA.n661 1.6924
R4092 VDDA.n810 VDDA.n660 1.6924
R4093 VDDA.n810 VDDA.n658 1.6924
R4094 VDDA.n810 VDDA.n657 1.6924
R4095 VDDA.n810 VDDA.n655 1.6924
R4096 VDDA.n810 VDDA.n654 1.6924
R4097 VDDA.n810 VDDA.n652 1.6924
R4098 VDDA.n810 VDDA.n651 1.6924
R4099 VDDA.n810 VDDA.n649 1.6924
R4100 VDDA.n810 VDDA.n648 1.6924
R4101 VDDA.n810 VDDA.n646 1.6924
R4102 VDDA.n810 VDDA.n645 1.6924
R4103 VDDA.n810 VDDA.n643 1.6924
R4104 VDDA.n810 VDDA.n642 1.6924
R4105 VDDA.n810 VDDA.n640 1.6924
R4106 VDDA.n810 VDDA.n639 1.6924
R4107 VDDA.n970 VDDA.n969 1.6924
R4108 VDDA.n970 VDDA.n833 1.6924
R4109 VDDA.n970 VDDA.n831 1.6924
R4110 VDDA.n970 VDDA.n830 1.6924
R4111 VDDA.n970 VDDA.n828 1.6924
R4112 VDDA.n970 VDDA.n827 1.6924
R4113 VDDA.n970 VDDA.n825 1.6924
R4114 VDDA.n970 VDDA.n824 1.6924
R4115 VDDA.n970 VDDA.n822 1.6924
R4116 VDDA.n970 VDDA.n821 1.6924
R4117 VDDA.n970 VDDA.n819 1.6924
R4118 VDDA.n970 VDDA.n818 1.6924
R4119 VDDA.n970 VDDA.n816 1.6924
R4120 VDDA.n970 VDDA.n815 1.6924
R4121 VDDA.n970 VDDA.n813 1.6924
R4122 VDDA.n970 VDDA.n812 1.6924
R4123 VDDA.n1140 VDDA.n461 1.6924
R4124 VDDA.n1132 VDDA.n461 1.6924
R4125 VDDA.n1122 VDDA.n461 1.6924
R4126 VDDA.n1120 VDDA.n461 1.6924
R4127 VDDA.n1110 VDDA.n461 1.6924
R4128 VDDA.n1102 VDDA.n461 1.6924
R4129 VDDA.n1092 VDDA.n461 1.6924
R4130 VDDA.n1090 VDDA.n461 1.6924
R4131 VDDA.n1080 VDDA.n461 1.6924
R4132 VDDA.n1072 VDDA.n461 1.6924
R4133 VDDA.n1062 VDDA.n461 1.6924
R4134 VDDA.n1060 VDDA.n461 1.6924
R4135 VDDA.n1050 VDDA.n461 1.6924
R4136 VDDA.n1042 VDDA.n461 1.6924
R4137 VDDA.n1032 VDDA.n461 1.6924
R4138 VDDA.n1030 VDDA.n461 1.6924
R4139 VDDA.n1158 VDDA.n485 1.6924
R4140 VDDA.n1158 VDDA.n484 1.6924
R4141 VDDA.n1158 VDDA.n482 1.6924
R4142 VDDA.n1158 VDDA.n481 1.6924
R4143 VDDA.n1158 VDDA.n479 1.6924
R4144 VDDA.n1158 VDDA.n478 1.6924
R4145 VDDA.n1158 VDDA.n476 1.6924
R4146 VDDA.n1158 VDDA.n475 1.6924
R4147 VDDA.n1158 VDDA.n473 1.6924
R4148 VDDA.n1158 VDDA.n472 1.6924
R4149 VDDA.n1158 VDDA.n470 1.6924
R4150 VDDA.n1158 VDDA.n469 1.6924
R4151 VDDA.n1158 VDDA.n467 1.6924
R4152 VDDA.n1158 VDDA.n466 1.6924
R4153 VDDA.n1158 VDDA.n464 1.6924
R4154 VDDA.n1158 VDDA.n463 1.6924
R4155 VDDA.n2254 VDDA.n1317 1.6924
R4156 VDDA.n2254 VDDA.n1181 1.6924
R4157 VDDA.n2254 VDDA.n1179 1.6924
R4158 VDDA.n2254 VDDA.n1178 1.6924
R4159 VDDA.n2254 VDDA.n1176 1.6924
R4160 VDDA.n2254 VDDA.n1175 1.6924
R4161 VDDA.n2254 VDDA.n1173 1.6924
R4162 VDDA.n2254 VDDA.n1172 1.6924
R4163 VDDA.n2254 VDDA.n1170 1.6924
R4164 VDDA.n2254 VDDA.n1169 1.6924
R4165 VDDA.n2254 VDDA.n1167 1.6924
R4166 VDDA.n2254 VDDA.n1166 1.6924
R4167 VDDA.n2254 VDDA.n1164 1.6924
R4168 VDDA.n2254 VDDA.n1163 1.6924
R4169 VDDA.n2254 VDDA.n1161 1.6924
R4170 VDDA.n2254 VDDA.n1160 1.6924
R4171 VDDA.n2253 VDDA.n1341 1.6924
R4172 VDDA.n2253 VDDA.n1340 1.6924
R4173 VDDA.n2253 VDDA.n1338 1.6924
R4174 VDDA.n2253 VDDA.n1337 1.6924
R4175 VDDA.n2253 VDDA.n1335 1.6924
R4176 VDDA.n2253 VDDA.n1334 1.6924
R4177 VDDA.n2253 VDDA.n1332 1.6924
R4178 VDDA.n2253 VDDA.n1331 1.6924
R4179 VDDA.n2253 VDDA.n1329 1.6924
R4180 VDDA.n2253 VDDA.n1328 1.6924
R4181 VDDA.n2253 VDDA.n1326 1.6924
R4182 VDDA.n2253 VDDA.n1325 1.6924
R4183 VDDA.n2253 VDDA.n1323 1.6924
R4184 VDDA.n2253 VDDA.n1322 1.6924
R4185 VDDA.n2253 VDDA.n1320 1.6924
R4186 VDDA.n2253 VDDA.n1319 1.6924
R4187 VDDA.n2580 VDDA.n195 1.6924
R4188 VDDA.n2572 VDDA.n195 1.6924
R4189 VDDA.n2562 VDDA.n195 1.6924
R4190 VDDA.n2560 VDDA.n195 1.6924
R4191 VDDA.n2550 VDDA.n195 1.6924
R4192 VDDA.n2542 VDDA.n195 1.6924
R4193 VDDA.n2532 VDDA.n195 1.6924
R4194 VDDA.n2530 VDDA.n195 1.6924
R4195 VDDA.n2520 VDDA.n195 1.6924
R4196 VDDA.n2512 VDDA.n195 1.6924
R4197 VDDA.n2502 VDDA.n195 1.6924
R4198 VDDA.n2500 VDDA.n195 1.6924
R4199 VDDA.n2490 VDDA.n195 1.6924
R4200 VDDA.n2482 VDDA.n195 1.6924
R4201 VDDA.n2472 VDDA.n195 1.6924
R4202 VDDA.n2470 VDDA.n195 1.6924
R4203 VDDA.n2598 VDDA.n219 1.6924
R4204 VDDA.n2598 VDDA.n218 1.6924
R4205 VDDA.n2598 VDDA.n216 1.6924
R4206 VDDA.n2598 VDDA.n215 1.6924
R4207 VDDA.n2598 VDDA.n213 1.6924
R4208 VDDA.n2598 VDDA.n212 1.6924
R4209 VDDA.n2598 VDDA.n210 1.6924
R4210 VDDA.n2598 VDDA.n209 1.6924
R4211 VDDA.n2598 VDDA.n207 1.6924
R4212 VDDA.n2598 VDDA.n206 1.6924
R4213 VDDA.n2598 VDDA.n204 1.6924
R4214 VDDA.n2598 VDDA.n203 1.6924
R4215 VDDA.n2598 VDDA.n201 1.6924
R4216 VDDA.n2598 VDDA.n200 1.6924
R4217 VDDA.n2598 VDDA.n198 1.6924
R4218 VDDA.n2598 VDDA.n197 1.6924
R4219 VDDA.n2758 VDDA.n2757 1.6924
R4220 VDDA.n2758 VDDA.n2621 1.6924
R4221 VDDA.n2758 VDDA.n2619 1.6924
R4222 VDDA.n2758 VDDA.n2618 1.6924
R4223 VDDA.n2758 VDDA.n2616 1.6924
R4224 VDDA.n2758 VDDA.n2615 1.6924
R4225 VDDA.n2758 VDDA.n2613 1.6924
R4226 VDDA.n2758 VDDA.n2612 1.6924
R4227 VDDA.n2758 VDDA.n2610 1.6924
R4228 VDDA.n2758 VDDA.n2609 1.6924
R4229 VDDA.n2758 VDDA.n2607 1.6924
R4230 VDDA.n2758 VDDA.n2606 1.6924
R4231 VDDA.n2758 VDDA.n2604 1.6924
R4232 VDDA.n2758 VDDA.n2603 1.6924
R4233 VDDA.n2758 VDDA.n2601 1.6924
R4234 VDDA.n2758 VDDA.n2600 1.6924
R4235 VDDA.n2928 VDDA.n17 1.6924
R4236 VDDA.n2920 VDDA.n17 1.6924
R4237 VDDA.n2910 VDDA.n17 1.6924
R4238 VDDA.n2908 VDDA.n17 1.6924
R4239 VDDA.n2898 VDDA.n17 1.6924
R4240 VDDA.n2890 VDDA.n17 1.6924
R4241 VDDA.n2880 VDDA.n17 1.6924
R4242 VDDA.n2878 VDDA.n17 1.6924
R4243 VDDA.n2868 VDDA.n17 1.6924
R4244 VDDA.n2860 VDDA.n17 1.6924
R4245 VDDA.n2850 VDDA.n17 1.6924
R4246 VDDA.n2848 VDDA.n17 1.6924
R4247 VDDA.n2838 VDDA.n17 1.6924
R4248 VDDA.n2830 VDDA.n17 1.6924
R4249 VDDA.n2820 VDDA.n17 1.6924
R4250 VDDA.n2818 VDDA.n17 1.6924
R4251 VDDA.n2946 VDDA.n41 1.6924
R4252 VDDA.n2946 VDDA.n40 1.6924
R4253 VDDA.n2946 VDDA.n38 1.6924
R4254 VDDA.n2946 VDDA.n37 1.6924
R4255 VDDA.n2946 VDDA.n35 1.6924
R4256 VDDA.n2946 VDDA.n34 1.6924
R4257 VDDA.n2946 VDDA.n32 1.6924
R4258 VDDA.n2946 VDDA.n31 1.6924
R4259 VDDA.n2946 VDDA.n29 1.6924
R4260 VDDA.n2946 VDDA.n28 1.6924
R4261 VDDA.n2946 VDDA.n26 1.6924
R4262 VDDA.n2946 VDDA.n25 1.6924
R4263 VDDA.n2946 VDDA.n23 1.6924
R4264 VDDA.n2946 VDDA.n22 1.6924
R4265 VDDA.n2946 VDDA.n20 1.6924
R4266 VDDA.n2946 VDDA.n19 1.6924
R4267 VDDA.n1578 VDDA.n1431 1.6924
R4268 VDDA.n1578 VDDA.n1430 1.6924
R4269 VDDA.n1578 VDDA.n1428 1.6924
R4270 VDDA.n1578 VDDA.n1427 1.6924
R4271 VDDA.n1578 VDDA.n1425 1.6924
R4272 VDDA.n1578 VDDA.n1424 1.6924
R4273 VDDA.n1578 VDDA.n1422 1.6924
R4274 VDDA.n1578 VDDA.n1421 1.6924
R4275 VDDA.n1578 VDDA.n1419 1.6924
R4276 VDDA.n1578 VDDA.n1418 1.6924
R4277 VDDA.n1578 VDDA.n1416 1.6924
R4278 VDDA.n1578 VDDA.n1415 1.6924
R4279 VDDA.n1578 VDDA.n1413 1.6924
R4280 VDDA.n1578 VDDA.n1412 1.6924
R4281 VDDA.n1578 VDDA.n1410 1.6924
R4282 VDDA.n1578 VDDA.n1409 1.6924
R4283 VDDA.n1906 VDDA.n1365 1.69118
R4284 VDDA.n1906 VDDA.n1364 1.69118
R4285 VDDA.n1906 VDDA.n1362 1.69118
R4286 VDDA.n1906 VDDA.n1361 1.69118
R4287 VDDA.n1906 VDDA.n1359 1.69118
R4288 VDDA.n1906 VDDA.n1358 1.69118
R4289 VDDA.n1906 VDDA.n1356 1.69118
R4290 VDDA.n1906 VDDA.n1355 1.69118
R4291 VDDA.n1906 VDDA.n1353 1.69118
R4292 VDDA.n1906 VDDA.n1352 1.69118
R4293 VDDA.n1906 VDDA.n1350 1.69118
R4294 VDDA.n1906 VDDA.n1349 1.69118
R4295 VDDA.n1906 VDDA.n1347 1.69118
R4296 VDDA.n1906 VDDA.n1346 1.69118
R4297 VDDA.n1906 VDDA.n1344 1.69118
R4298 VDDA.n1906 VDDA.n1343 1.69118
R4299 VDDA.n371 VDDA.n370 1.63212
R4300 VDDA.n378 VDDA.n376 1.63212
R4301 VDDA.n383 VDDA.n375 1.59823
R4302 VDDA.n375 VDDA.n374 1.56962
R4303 VDDA.n382 VDDA.n381 1.56962
R4304 VDDA.n1788 VDDA.n1391 1.56177
R4305 VDDA.n1765 VDDA.n1391 1.50969
R4306 VDDA.n1402 VDDA.n1391 1.44719
R4307 VDDA.n450 VDDA.n384 1.31821
R4308 VDDA.n2398 VDDA.n384 1.31821
R4309 VDDA.n1651 VDDA.n1650 1.20209
R4310 VDDA.n1942 VDDA.n1941 1.1893
R4311 VDDA.n2392 VDDA.n437 1.13592
R4312 VDDA.n2336 VDDA.n2335 1.13592
R4313 VDDA.n428 VDDA.n426 1.07342
R4314 VDDA.n2332 VDDA.n2324 1.06821
R4315 VDDA.n2402 VDDA.n365 1.03383
R4316 VDDA.n2404 VDDA.n2403 1.03383
R4317 VDDA.n2264 VDDA.n452 1.03383
R4318 VDDA.n2266 VDDA.n2265 1.03383
R4319 VDDA.n2358 VDDA.n2342 0.932792
R4320 VDDA.n2391 VDDA.n2390 0.932792
R4321 VDDA.n2396 VDDA.n2395 0.922375
R4322 VDDA.n2340 VDDA.n2286 0.922375
R4323 VDDA.n2080 VDDA.n2079 0.807792
R4324 VDDA.n1948 VDDA.n1947 0.802583
R4325 VDDA.n2003 VDDA.n2002 0.792167
R4326 VDDA.n2417 VDDA.n365 0.792167
R4327 VDDA.n2405 VDDA.n2404 0.792167
R4328 VDDA.n2279 VDDA.n452 0.792167
R4329 VDDA.n2267 VDDA.n2266 0.792167
R4330 VDDA.n1940 VDDA.n1939 0.75233
R4331 VDDA.n2130 VDDA.n2129 0.734875
R4332 VDDA.n2009 VDDA.n2008 0.661958
R4333 VDDA.n1941 VDDA.n1940 0.648711
R4334 VDDA.n2260 VDDA.n456 0.646333
R4335 VDDA.n2591 VDDA.n2589 0.646333
R4336 VDDA.n2409 VDDA.n2407 0.6255
R4337 VDDA.n2412 VDDA.n2409 0.6255
R4338 VDDA.n2414 VDDA.n2412 0.6255
R4339 VDDA.n2416 VDDA.n2414 0.6255
R4340 VDDA.n2271 VDDA.n2269 0.6255
R4341 VDDA.n2274 VDDA.n2271 0.6255
R4342 VDDA.n2276 VDDA.n2274 0.6255
R4343 VDDA.n2278 VDDA.n2276 0.6255
R4344 VDDA.n2263 VDDA.n2262 0.490083
R4345 VDDA.n2587 VDDA.n2418 0.490083
R4346 VDDA.n2263 VDDA.n451 0.3755
R4347 VDDA.n2280 VDDA.n451 0.3755
R4348 VDDA.n2401 VDDA.n364 0.3755
R4349 VDDA.n2418 VDDA.n364 0.3755
R4350 VDDA.n1996 VDDA.n1995 0.333833
R4351 VDDA.n2074 VDDA.n2073 0.328625
R4352 VDDA.n2320 VDDA.n2319 0.323417
R4353 VDDA.n424 VDDA.n423 0.323417
R4354 VDDA.n2127 VDDA.n2126 0.292167
R4355 VDDA.n2123 VDDA.n2122 0.292167
R4356 VDDA.n2116 VDDA.n2115 0.292167
R4357 VDDA.n2086 VDDA.n2085 0.292167
R4358 VDDA.n976 VDDA.n633 0.28175
R4359 VDDA.n1147 VDDA.n978 0.28175
R4360 VDDA.n1151 VDDA.n1149 0.28175
R4361 VDDA.n2764 VDDA.n190 0.28175
R4362 VDDA.n2935 VDDA.n2766 0.28175
R4363 VDDA.n2938 VDDA.n2937 0.28175
R4364 VDDA.n2136 VDDA.n2135 0.276542
R4365 VDDA.n2330 VDDA.n2329 0.266125
R4366 VDDA.n435 VDDA.n434 0.266125
R4367 VDDA.n2338 VDDA.n2302 0.266125
R4368 VDDA.n2393 VDDA.n403 0.266125
R4369 VDDA.n2285 VDDA.n2280 0.234875
R4370 VDDA.n2401 VDDA.n2400 0.234875
R4371 VDDA.n1767 VDDA.n1766 0.229667
R4372 VDDA.n1787 VDDA.n1786 0.229667
R4373 VDDA.n2079 VDDA.n2074 0.229667
R4374 VDDA.n1768 VDDA.n1398 0.208833
R4375 VDDA.n1768 VDDA.n1767 0.208833
R4376 VDDA.n1780 VDDA.n1392 0.208833
R4377 VDDA.n1786 VDDA.n1392 0.208833
R4378 VDDA.n2041 VDDA.n2027 0.208833
R4379 VDDA.n2035 VDDA.n2027 0.208833
R4380 VDDA.n2035 VDDA.n2034 0.208833
R4381 VDDA.n2050 VDDA.n2048 0.208833
R4382 VDDA.n2051 VDDA.n2050 0.208833
R4383 VDDA.n2051 VDDA.n2020 0.208833
R4384 VDDA.n2073 VDDA.n2072 0.188
R4385 VDDA.n2072 VDDA.n2071 0.188
R4386 VDDA.n2071 VDDA.n2070 0.188
R4387 VDDA.n2070 VDDA.n2069 0.188
R4388 VDDA.n2069 VDDA.n2068 0.188
R4389 VDDA.n2068 VDDA.n2067 0.188
R4390 VDDA.n2067 VDDA.n2066 0.188
R4391 VDDA.n2066 VDDA.n2065 0.188
R4392 VDDA.n2360 VDDA.n2358 0.172375
R4393 VDDA.n2361 VDDA.n2360 0.172375
R4394 VDDA.n2362 VDDA.n439 0.172375
R4395 VDDA.n2390 VDDA.n439 0.172375
R4396 VDDA.t128 VDDA.t420 0.1603
R4397 VDDA.t406 VDDA.t103 0.1603
R4398 VDDA.t146 VDDA.t391 0.1603
R4399 VDDA.t90 VDDA.t388 0.1603
R4400 VDDA.t59 VDDA.t101 0.1603
R4401 VDDA.n1794 VDDA.n1793 0.159591
R4402 VDDA.n1795 VDDA.n1794 0.159591
R4403 VDDA.n1795 VDDA.n1389 0.159591
R4404 VDDA.n1805 VDDA.n1387 0.159591
R4405 VDDA.n1813 VDDA.n1387 0.159591
R4406 VDDA.n1814 VDDA.n1813 0.159591
R4407 VDDA.n1824 VDDA.n1823 0.159591
R4408 VDDA.n1825 VDDA.n1824 0.159591
R4409 VDDA.n1825 VDDA.n1383 0.159591
R4410 VDDA.n1835 VDDA.n1381 0.159591
R4411 VDDA.n1843 VDDA.n1381 0.159591
R4412 VDDA.n1844 VDDA.n1843 0.159591
R4413 VDDA.n1854 VDDA.n1853 0.159591
R4414 VDDA.n1855 VDDA.n1854 0.159591
R4415 VDDA.n1855 VDDA.n1377 0.159591
R4416 VDDA.n1865 VDDA.n1375 0.159591
R4417 VDDA.n1873 VDDA.n1375 0.159591
R4418 VDDA.n1874 VDDA.n1873 0.159591
R4419 VDDA.n1884 VDDA.n1883 0.159591
R4420 VDDA.n1885 VDDA.n1884 0.159591
R4421 VDDA.n1885 VDDA.n1371 0.159591
R4422 VDDA.n1895 VDDA.n1369 0.159591
R4423 VDDA.n1903 VDDA.n1369 0.159591
R4424 VDDA.n1792 VDDA.n1390 0.159591
R4425 VDDA.n1798 VDDA.n1390 0.159591
R4426 VDDA.n1799 VDDA.n1798 0.159591
R4427 VDDA.n1809 VDDA.n1808 0.159591
R4428 VDDA.n1812 VDDA.n1809 0.159591
R4429 VDDA.n1812 VDDA.n1386 0.159591
R4430 VDDA.n1822 VDDA.n1384 0.159591
R4431 VDDA.n1828 VDDA.n1384 0.159591
R4432 VDDA.n1829 VDDA.n1828 0.159591
R4433 VDDA.n1839 VDDA.n1838 0.159591
R4434 VDDA.n1842 VDDA.n1839 0.159591
R4435 VDDA.n1842 VDDA.n1380 0.159591
R4436 VDDA.n1852 VDDA.n1378 0.159591
R4437 VDDA.n1858 VDDA.n1378 0.159591
R4438 VDDA.n1859 VDDA.n1858 0.159591
R4439 VDDA.n1869 VDDA.n1868 0.159591
R4440 VDDA.n1872 VDDA.n1869 0.159591
R4441 VDDA.n1872 VDDA.n1374 0.159591
R4442 VDDA.n1882 VDDA.n1372 0.159591
R4443 VDDA.n1888 VDDA.n1372 0.159591
R4444 VDDA.n1889 VDDA.n1888 0.159591
R4445 VDDA.n1899 VDDA.n1898 0.159591
R4446 VDDA.n1902 VDDA.n1899 0.159591
R4447 VDDA.n1902 VDDA.n1368 0.159591
R4448 VDDA.n1457 VDDA.t91 0.159278
R4449 VDDA.n1458 VDDA.t62 0.159278
R4450 VDDA.n1459 VDDA.t147 0.159278
R4451 VDDA.n1460 VDDA.t145 0.159278
R4452 VDDA.n1793 VDDA.n1789 0.148227
R4453 VDDA.n1803 VDDA.n1389 0.148227
R4454 VDDA.n1805 VDDA.n1804 0.148227
R4455 VDDA.n1815 VDDA.n1814 0.148227
R4456 VDDA.n1823 VDDA.n1385 0.148227
R4457 VDDA.n1833 VDDA.n1383 0.148227
R4458 VDDA.n1835 VDDA.n1834 0.148227
R4459 VDDA.n1845 VDDA.n1844 0.148227
R4460 VDDA.n1853 VDDA.n1379 0.148227
R4461 VDDA.n1863 VDDA.n1377 0.148227
R4462 VDDA.n1865 VDDA.n1864 0.148227
R4463 VDDA.n1875 VDDA.n1874 0.148227
R4464 VDDA.n1883 VDDA.n1373 0.148227
R4465 VDDA.n1893 VDDA.n1371 0.148227
R4466 VDDA.n1895 VDDA.n1894 0.148227
R4467 VDDA.n1792 VDDA.n1790 0.148227
R4468 VDDA.n1802 VDDA.n1799 0.148227
R4469 VDDA.n1808 VDDA.n1388 0.148227
R4470 VDDA.n1818 VDDA.n1386 0.148227
R4471 VDDA.n1822 VDDA.n1819 0.148227
R4472 VDDA.n1832 VDDA.n1829 0.148227
R4473 VDDA.n1838 VDDA.n1382 0.148227
R4474 VDDA.n1848 VDDA.n1380 0.148227
R4475 VDDA.n1852 VDDA.n1849 0.148227
R4476 VDDA.n1862 VDDA.n1859 0.148227
R4477 VDDA.n1868 VDDA.n1376 0.148227
R4478 VDDA.n1878 VDDA.n1374 0.148227
R4479 VDDA.n1882 VDDA.n1879 0.148227
R4480 VDDA.n1892 VDDA.n1889 0.148227
R4481 VDDA.n1898 VDDA.n1370 0.148227
R4482 VDDA.n1464 VDDA.n1455 0.146333
R4483 VDDA.n1470 VDDA.n1455 0.146333
R4484 VDDA.n1471 VDDA.n1470 0.146333
R4485 VDDA.n1481 VDDA.n1480 0.146333
R4486 VDDA.n1484 VDDA.n1481 0.146333
R4487 VDDA.n1484 VDDA.n1451 0.146333
R4488 VDDA.n1494 VDDA.n1449 0.146333
R4489 VDDA.n1500 VDDA.n1449 0.146333
R4490 VDDA.n1501 VDDA.n1500 0.146333
R4491 VDDA.n1511 VDDA.n1510 0.146333
R4492 VDDA.n1514 VDDA.n1511 0.146333
R4493 VDDA.n1514 VDDA.n1445 0.146333
R4494 VDDA.n1524 VDDA.n1443 0.146333
R4495 VDDA.n1530 VDDA.n1443 0.146333
R4496 VDDA.n1531 VDDA.n1530 0.146333
R4497 VDDA.n1541 VDDA.n1540 0.146333
R4498 VDDA.n1544 VDDA.n1541 0.146333
R4499 VDDA.n1544 VDDA.n1439 0.146333
R4500 VDDA.n1554 VDDA.n1437 0.146333
R4501 VDDA.n1560 VDDA.n1437 0.146333
R4502 VDDA.n1561 VDDA.n1560 0.146333
R4503 VDDA.n1571 VDDA.n1570 0.146333
R4504 VDDA.n1574 VDDA.n1571 0.146333
R4505 VDDA.n1574 VDDA.n1433 0.146333
R4506 VDDA.n2139 VDDA.n1930 0.146333
R4507 VDDA.n2145 VDDA.n1930 0.146333
R4508 VDDA.n2146 VDDA.n2145 0.146333
R4509 VDDA.n2156 VDDA.n2155 0.146333
R4510 VDDA.n2159 VDDA.n2156 0.146333
R4511 VDDA.n2159 VDDA.n1926 0.146333
R4512 VDDA.n2169 VDDA.n1924 0.146333
R4513 VDDA.n2175 VDDA.n1924 0.146333
R4514 VDDA.n2176 VDDA.n2175 0.146333
R4515 VDDA.n2186 VDDA.n2185 0.146333
R4516 VDDA.n2189 VDDA.n2186 0.146333
R4517 VDDA.n2189 VDDA.n1920 0.146333
R4518 VDDA.n2199 VDDA.n1918 0.146333
R4519 VDDA.n2205 VDDA.n1918 0.146333
R4520 VDDA.n2206 VDDA.n2205 0.146333
R4521 VDDA.n2216 VDDA.n2215 0.146333
R4522 VDDA.n2219 VDDA.n2216 0.146333
R4523 VDDA.n2219 VDDA.n1914 0.146333
R4524 VDDA.n2229 VDDA.n1912 0.146333
R4525 VDDA.n2235 VDDA.n1912 0.146333
R4526 VDDA.n2236 VDDA.n2235 0.146333
R4527 VDDA.n2246 VDDA.n2245 0.146333
R4528 VDDA.n2249 VDDA.n2246 0.146333
R4529 VDDA.n2249 VDDA.n1908 0.146333
R4530 VDDA.n89 VDDA.n85 0.146333
R4531 VDDA.n93 VDDA.n85 0.146333
R4532 VDDA.n94 VDDA.n93 0.146333
R4533 VDDA.n102 VDDA.n101 0.146333
R4534 VDDA.n105 VDDA.n102 0.146333
R4535 VDDA.n105 VDDA.n77 0.146333
R4536 VDDA.n113 VDDA.n73 0.146333
R4537 VDDA.n117 VDDA.n73 0.146333
R4538 VDDA.n118 VDDA.n117 0.146333
R4539 VDDA.n126 VDDA.n125 0.146333
R4540 VDDA.n129 VDDA.n126 0.146333
R4541 VDDA.n129 VDDA.n65 0.146333
R4542 VDDA.n137 VDDA.n61 0.146333
R4543 VDDA.n141 VDDA.n61 0.146333
R4544 VDDA.n142 VDDA.n141 0.146333
R4545 VDDA.n150 VDDA.n149 0.146333
R4546 VDDA.n153 VDDA.n150 0.146333
R4547 VDDA.n153 VDDA.n53 0.146333
R4548 VDDA.n161 VDDA.n49 0.146333
R4549 VDDA.n165 VDDA.n49 0.146333
R4550 VDDA.n166 VDDA.n165 0.146333
R4551 VDDA.n174 VDDA.n173 0.146333
R4552 VDDA.n177 VDDA.n174 0.146333
R4553 VDDA.n177 VDDA.n43 0.146333
R4554 VDDA.n2816 VDDA.n2813 0.146333
R4555 VDDA.n2822 VDDA.n2813 0.146333
R4556 VDDA.n2822 VDDA.n2811 0.146333
R4557 VDDA.n2832 VDDA.n2807 0.146333
R4558 VDDA.n2836 VDDA.n2807 0.146333
R4559 VDDA.n2836 VDDA.n2805 0.146333
R4560 VDDA.n2846 VDDA.n2801 0.146333
R4561 VDDA.n2852 VDDA.n2801 0.146333
R4562 VDDA.n2852 VDDA.n2799 0.146333
R4563 VDDA.n2862 VDDA.n2795 0.146333
R4564 VDDA.n2866 VDDA.n2795 0.146333
R4565 VDDA.n2866 VDDA.n2793 0.146333
R4566 VDDA.n2876 VDDA.n2789 0.146333
R4567 VDDA.n2882 VDDA.n2789 0.146333
R4568 VDDA.n2882 VDDA.n2787 0.146333
R4569 VDDA.n2892 VDDA.n2783 0.146333
R4570 VDDA.n2896 VDDA.n2783 0.146333
R4571 VDDA.n2896 VDDA.n2781 0.146333
R4572 VDDA.n2906 VDDA.n2777 0.146333
R4573 VDDA.n2912 VDDA.n2777 0.146333
R4574 VDDA.n2912 VDDA.n2775 0.146333
R4575 VDDA.n2922 VDDA.n2771 0.146333
R4576 VDDA.n2926 VDDA.n2771 0.146333
R4577 VDDA.n2926 VDDA.n2769 0.146333
R4578 VDDA.n2668 VDDA.n2667 0.146333
R4579 VDDA.n2671 VDDA.n2668 0.146333
R4580 VDDA.n2671 VDDA.n2661 0.146333
R4581 VDDA.n2679 VDDA.n2657 0.146333
R4582 VDDA.n2683 VDDA.n2657 0.146333
R4583 VDDA.n2684 VDDA.n2683 0.146333
R4584 VDDA.n2692 VDDA.n2691 0.146333
R4585 VDDA.n2695 VDDA.n2692 0.146333
R4586 VDDA.n2695 VDDA.n2649 0.146333
R4587 VDDA.n2703 VDDA.n2645 0.146333
R4588 VDDA.n2707 VDDA.n2645 0.146333
R4589 VDDA.n2708 VDDA.n2707 0.146333
R4590 VDDA.n2716 VDDA.n2715 0.146333
R4591 VDDA.n2719 VDDA.n2716 0.146333
R4592 VDDA.n2719 VDDA.n2637 0.146333
R4593 VDDA.n2727 VDDA.n2633 0.146333
R4594 VDDA.n2731 VDDA.n2633 0.146333
R4595 VDDA.n2732 VDDA.n2731 0.146333
R4596 VDDA.n2740 VDDA.n2739 0.146333
R4597 VDDA.n2743 VDDA.n2740 0.146333
R4598 VDDA.n2743 VDDA.n2625 0.146333
R4599 VDDA.n2751 VDDA.n2623 0.146333
R4600 VDDA.n2755 VDDA.n2623 0.146333
R4601 VDDA.n2755 VDDA.n193 0.146333
R4602 VDDA.n267 VDDA.n263 0.146333
R4603 VDDA.n271 VDDA.n263 0.146333
R4604 VDDA.n272 VDDA.n271 0.146333
R4605 VDDA.n280 VDDA.n279 0.146333
R4606 VDDA.n283 VDDA.n280 0.146333
R4607 VDDA.n283 VDDA.n255 0.146333
R4608 VDDA.n291 VDDA.n251 0.146333
R4609 VDDA.n295 VDDA.n251 0.146333
R4610 VDDA.n296 VDDA.n295 0.146333
R4611 VDDA.n304 VDDA.n303 0.146333
R4612 VDDA.n307 VDDA.n304 0.146333
R4613 VDDA.n307 VDDA.n243 0.146333
R4614 VDDA.n315 VDDA.n239 0.146333
R4615 VDDA.n319 VDDA.n239 0.146333
R4616 VDDA.n320 VDDA.n319 0.146333
R4617 VDDA.n328 VDDA.n327 0.146333
R4618 VDDA.n331 VDDA.n328 0.146333
R4619 VDDA.n331 VDDA.n231 0.146333
R4620 VDDA.n339 VDDA.n227 0.146333
R4621 VDDA.n343 VDDA.n227 0.146333
R4622 VDDA.n344 VDDA.n343 0.146333
R4623 VDDA.n352 VDDA.n351 0.146333
R4624 VDDA.n355 VDDA.n352 0.146333
R4625 VDDA.n355 VDDA.n221 0.146333
R4626 VDDA.n2468 VDDA.n2465 0.146333
R4627 VDDA.n2474 VDDA.n2465 0.146333
R4628 VDDA.n2474 VDDA.n2463 0.146333
R4629 VDDA.n2484 VDDA.n2459 0.146333
R4630 VDDA.n2488 VDDA.n2459 0.146333
R4631 VDDA.n2488 VDDA.n2457 0.146333
R4632 VDDA.n2498 VDDA.n2453 0.146333
R4633 VDDA.n2504 VDDA.n2453 0.146333
R4634 VDDA.n2504 VDDA.n2451 0.146333
R4635 VDDA.n2514 VDDA.n2447 0.146333
R4636 VDDA.n2518 VDDA.n2447 0.146333
R4637 VDDA.n2518 VDDA.n2445 0.146333
R4638 VDDA.n2528 VDDA.n2441 0.146333
R4639 VDDA.n2534 VDDA.n2441 0.146333
R4640 VDDA.n2534 VDDA.n2439 0.146333
R4641 VDDA.n2544 VDDA.n2435 0.146333
R4642 VDDA.n2548 VDDA.n2435 0.146333
R4643 VDDA.n2548 VDDA.n2433 0.146333
R4644 VDDA.n2558 VDDA.n2429 0.146333
R4645 VDDA.n2564 VDDA.n2429 0.146333
R4646 VDDA.n2564 VDDA.n2427 0.146333
R4647 VDDA.n2574 VDDA.n2423 0.146333
R4648 VDDA.n2578 VDDA.n2423 0.146333
R4649 VDDA.n2578 VDDA.n2421 0.146333
R4650 VDDA.n1228 VDDA.n1227 0.146333
R4651 VDDA.n1231 VDDA.n1228 0.146333
R4652 VDDA.n1231 VDDA.n1221 0.146333
R4653 VDDA.n1239 VDDA.n1217 0.146333
R4654 VDDA.n1243 VDDA.n1217 0.146333
R4655 VDDA.n1244 VDDA.n1243 0.146333
R4656 VDDA.n1252 VDDA.n1251 0.146333
R4657 VDDA.n1255 VDDA.n1252 0.146333
R4658 VDDA.n1255 VDDA.n1209 0.146333
R4659 VDDA.n1263 VDDA.n1205 0.146333
R4660 VDDA.n1267 VDDA.n1205 0.146333
R4661 VDDA.n1268 VDDA.n1267 0.146333
R4662 VDDA.n1276 VDDA.n1275 0.146333
R4663 VDDA.n1279 VDDA.n1276 0.146333
R4664 VDDA.n1279 VDDA.n1197 0.146333
R4665 VDDA.n1287 VDDA.n1193 0.146333
R4666 VDDA.n1291 VDDA.n1193 0.146333
R4667 VDDA.n1292 VDDA.n1291 0.146333
R4668 VDDA.n1300 VDDA.n1299 0.146333
R4669 VDDA.n1303 VDDA.n1300 0.146333
R4670 VDDA.n1303 VDDA.n1185 0.146333
R4671 VDDA.n1311 VDDA.n1183 0.146333
R4672 VDDA.n1315 VDDA.n1183 0.146333
R4673 VDDA.n1315 VDDA.n459 0.146333
R4674 VDDA.n533 VDDA.n529 0.146333
R4675 VDDA.n537 VDDA.n529 0.146333
R4676 VDDA.n538 VDDA.n537 0.146333
R4677 VDDA.n546 VDDA.n545 0.146333
R4678 VDDA.n549 VDDA.n546 0.146333
R4679 VDDA.n549 VDDA.n521 0.146333
R4680 VDDA.n557 VDDA.n517 0.146333
R4681 VDDA.n561 VDDA.n517 0.146333
R4682 VDDA.n562 VDDA.n561 0.146333
R4683 VDDA.n570 VDDA.n569 0.146333
R4684 VDDA.n573 VDDA.n570 0.146333
R4685 VDDA.n573 VDDA.n509 0.146333
R4686 VDDA.n581 VDDA.n505 0.146333
R4687 VDDA.n585 VDDA.n505 0.146333
R4688 VDDA.n586 VDDA.n585 0.146333
R4689 VDDA.n594 VDDA.n593 0.146333
R4690 VDDA.n597 VDDA.n594 0.146333
R4691 VDDA.n597 VDDA.n497 0.146333
R4692 VDDA.n605 VDDA.n493 0.146333
R4693 VDDA.n609 VDDA.n493 0.146333
R4694 VDDA.n610 VDDA.n609 0.146333
R4695 VDDA.n618 VDDA.n617 0.146333
R4696 VDDA.n621 VDDA.n618 0.146333
R4697 VDDA.n621 VDDA.n487 0.146333
R4698 VDDA.n1028 VDDA.n1025 0.146333
R4699 VDDA.n1034 VDDA.n1025 0.146333
R4700 VDDA.n1034 VDDA.n1023 0.146333
R4701 VDDA.n1044 VDDA.n1019 0.146333
R4702 VDDA.n1048 VDDA.n1019 0.146333
R4703 VDDA.n1048 VDDA.n1017 0.146333
R4704 VDDA.n1058 VDDA.n1013 0.146333
R4705 VDDA.n1064 VDDA.n1013 0.146333
R4706 VDDA.n1064 VDDA.n1011 0.146333
R4707 VDDA.n1074 VDDA.n1007 0.146333
R4708 VDDA.n1078 VDDA.n1007 0.146333
R4709 VDDA.n1078 VDDA.n1005 0.146333
R4710 VDDA.n1088 VDDA.n1001 0.146333
R4711 VDDA.n1094 VDDA.n1001 0.146333
R4712 VDDA.n1094 VDDA.n999 0.146333
R4713 VDDA.n1104 VDDA.n995 0.146333
R4714 VDDA.n1108 VDDA.n995 0.146333
R4715 VDDA.n1108 VDDA.n993 0.146333
R4716 VDDA.n1118 VDDA.n989 0.146333
R4717 VDDA.n1124 VDDA.n989 0.146333
R4718 VDDA.n1124 VDDA.n987 0.146333
R4719 VDDA.n1134 VDDA.n983 0.146333
R4720 VDDA.n1138 VDDA.n983 0.146333
R4721 VDDA.n1138 VDDA.n981 0.146333
R4722 VDDA.n880 VDDA.n879 0.146333
R4723 VDDA.n883 VDDA.n880 0.146333
R4724 VDDA.n883 VDDA.n873 0.146333
R4725 VDDA.n891 VDDA.n869 0.146333
R4726 VDDA.n895 VDDA.n869 0.146333
R4727 VDDA.n896 VDDA.n895 0.146333
R4728 VDDA.n904 VDDA.n903 0.146333
R4729 VDDA.n907 VDDA.n904 0.146333
R4730 VDDA.n907 VDDA.n861 0.146333
R4731 VDDA.n915 VDDA.n857 0.146333
R4732 VDDA.n919 VDDA.n857 0.146333
R4733 VDDA.n920 VDDA.n919 0.146333
R4734 VDDA.n928 VDDA.n927 0.146333
R4735 VDDA.n931 VDDA.n928 0.146333
R4736 VDDA.n931 VDDA.n849 0.146333
R4737 VDDA.n939 VDDA.n845 0.146333
R4738 VDDA.n943 VDDA.n845 0.146333
R4739 VDDA.n944 VDDA.n943 0.146333
R4740 VDDA.n952 VDDA.n951 0.146333
R4741 VDDA.n955 VDDA.n952 0.146333
R4742 VDDA.n955 VDDA.n837 0.146333
R4743 VDDA.n963 VDDA.n835 0.146333
R4744 VDDA.n967 VDDA.n835 0.146333
R4745 VDDA.n967 VDDA.n636 0.146333
R4746 VDDA.n687 VDDA.n685 0.146333
R4747 VDDA.n693 VDDA.n685 0.146333
R4748 VDDA.n694 VDDA.n693 0.146333
R4749 VDDA.n704 VDDA.n703 0.146333
R4750 VDDA.n707 VDDA.n704 0.146333
R4751 VDDA.n707 VDDA.n681 0.146333
R4752 VDDA.n717 VDDA.n679 0.146333
R4753 VDDA.n723 VDDA.n679 0.146333
R4754 VDDA.n724 VDDA.n723 0.146333
R4755 VDDA.n734 VDDA.n733 0.146333
R4756 VDDA.n737 VDDA.n734 0.146333
R4757 VDDA.n737 VDDA.n675 0.146333
R4758 VDDA.n747 VDDA.n673 0.146333
R4759 VDDA.n753 VDDA.n673 0.146333
R4760 VDDA.n754 VDDA.n753 0.146333
R4761 VDDA.n764 VDDA.n763 0.146333
R4762 VDDA.n767 VDDA.n764 0.146333
R4763 VDDA.n767 VDDA.n669 0.146333
R4764 VDDA.n777 VDDA.n667 0.146333
R4765 VDDA.n783 VDDA.n667 0.146333
R4766 VDDA.n784 VDDA.n783 0.146333
R4767 VDDA.n794 VDDA.n793 0.146333
R4768 VDDA.n797 VDDA.n794 0.146333
R4769 VDDA.n797 VDDA.n663 0.146333
R4770 VDDA.n1804 VDDA.n1803 0.136864
R4771 VDDA.n1815 VDDA.n1385 0.136864
R4772 VDDA.n1834 VDDA.n1833 0.136864
R4773 VDDA.n1845 VDDA.n1379 0.136864
R4774 VDDA.n1864 VDDA.n1863 0.136864
R4775 VDDA.n1875 VDDA.n1373 0.136864
R4776 VDDA.n1894 VDDA.n1893 0.136864
R4777 VDDA.n1802 VDDA.n1388 0.136864
R4778 VDDA.n1819 VDDA.n1818 0.136864
R4779 VDDA.n1832 VDDA.n1382 0.136864
R4780 VDDA.n1849 VDDA.n1848 0.136864
R4781 VDDA.n1862 VDDA.n1376 0.136864
R4782 VDDA.n1879 VDDA.n1878 0.136864
R4783 VDDA.n1892 VDDA.n1370 0.136864
R4784 VDDA.n1460 VDDA.t102 0.1368
R4785 VDDA.n1460 VDDA.t128 0.1368
R4786 VDDA.n1459 VDDA.t125 0.1368
R4787 VDDA.n1459 VDDA.t406 0.1368
R4788 VDDA.n1458 VDDA.t372 0.1368
R4789 VDDA.n1458 VDDA.t146 0.1368
R4790 VDDA.n1457 VDDA.t148 0.1368
R4791 VDDA.n1457 VDDA.t90 0.1368
R4792 VDDA.n1456 VDDA.t63 0.1368
R4793 VDDA.n1456 VDDA.t59 0.1368
R4794 VDDA.n1464 VDDA.n1462 0.135917
R4795 VDDA.n1474 VDDA.n1471 0.135917
R4796 VDDA.n1480 VDDA.n1453 0.135917
R4797 VDDA.n1490 VDDA.n1451 0.135917
R4798 VDDA.n1494 VDDA.n1491 0.135917
R4799 VDDA.n1504 VDDA.n1501 0.135917
R4800 VDDA.n1510 VDDA.n1447 0.135917
R4801 VDDA.n1520 VDDA.n1445 0.135917
R4802 VDDA.n1524 VDDA.n1521 0.135917
R4803 VDDA.n1534 VDDA.n1531 0.135917
R4804 VDDA.n1540 VDDA.n1441 0.135917
R4805 VDDA.n1550 VDDA.n1439 0.135917
R4806 VDDA.n1554 VDDA.n1551 0.135917
R4807 VDDA.n1564 VDDA.n1561 0.135917
R4808 VDDA.n1570 VDDA.n1435 0.135917
R4809 VDDA.n2139 VDDA.n2137 0.135917
R4810 VDDA.n2149 VDDA.n2146 0.135917
R4811 VDDA.n2155 VDDA.n1928 0.135917
R4812 VDDA.n2165 VDDA.n1926 0.135917
R4813 VDDA.n2169 VDDA.n2166 0.135917
R4814 VDDA.n2179 VDDA.n2176 0.135917
R4815 VDDA.n2185 VDDA.n1922 0.135917
R4816 VDDA.n2195 VDDA.n1920 0.135917
R4817 VDDA.n2199 VDDA.n2196 0.135917
R4818 VDDA.n2209 VDDA.n2206 0.135917
R4819 VDDA.n2215 VDDA.n1916 0.135917
R4820 VDDA.n2225 VDDA.n1914 0.135917
R4821 VDDA.n2229 VDDA.n2226 0.135917
R4822 VDDA.n2239 VDDA.n2236 0.135917
R4823 VDDA.n2245 VDDA.n1910 0.135917
R4824 VDDA.n97 VDDA.n94 0.135917
R4825 VDDA.n101 VDDA.n81 0.135917
R4826 VDDA.n109 VDDA.n77 0.135917
R4827 VDDA.n113 VDDA.n110 0.135917
R4828 VDDA.n121 VDDA.n118 0.135917
R4829 VDDA.n125 VDDA.n69 0.135917
R4830 VDDA.n133 VDDA.n65 0.135917
R4831 VDDA.n137 VDDA.n134 0.135917
R4832 VDDA.n145 VDDA.n142 0.135917
R4833 VDDA.n149 VDDA.n57 0.135917
R4834 VDDA.n157 VDDA.n53 0.135917
R4835 VDDA.n161 VDDA.n158 0.135917
R4836 VDDA.n169 VDDA.n166 0.135917
R4837 VDDA.n173 VDDA.n45 0.135917
R4838 VDDA.n2944 VDDA.n43 0.135917
R4839 VDDA.n2826 VDDA.n2811 0.135917
R4840 VDDA.n2832 VDDA.n2809 0.135917
R4841 VDDA.n2842 VDDA.n2805 0.135917
R4842 VDDA.n2846 VDDA.n2803 0.135917
R4843 VDDA.n2856 VDDA.n2799 0.135917
R4844 VDDA.n2862 VDDA.n2797 0.135917
R4845 VDDA.n2872 VDDA.n2793 0.135917
R4846 VDDA.n2876 VDDA.n2791 0.135917
R4847 VDDA.n2886 VDDA.n2787 0.135917
R4848 VDDA.n2892 VDDA.n2785 0.135917
R4849 VDDA.n2902 VDDA.n2781 0.135917
R4850 VDDA.n2906 VDDA.n2779 0.135917
R4851 VDDA.n2916 VDDA.n2775 0.135917
R4852 VDDA.n2922 VDDA.n2773 0.135917
R4853 VDDA.n2931 VDDA.n2769 0.135917
R4854 VDDA.n2675 VDDA.n2661 0.135917
R4855 VDDA.n2679 VDDA.n2676 0.135917
R4856 VDDA.n2687 VDDA.n2684 0.135917
R4857 VDDA.n2691 VDDA.n2653 0.135917
R4858 VDDA.n2699 VDDA.n2649 0.135917
R4859 VDDA.n2703 VDDA.n2700 0.135917
R4860 VDDA.n2711 VDDA.n2708 0.135917
R4861 VDDA.n2715 VDDA.n2641 0.135917
R4862 VDDA.n2723 VDDA.n2637 0.135917
R4863 VDDA.n2727 VDDA.n2724 0.135917
R4864 VDDA.n2735 VDDA.n2732 0.135917
R4865 VDDA.n2739 VDDA.n2629 0.135917
R4866 VDDA.n2747 VDDA.n2625 0.135917
R4867 VDDA.n2751 VDDA.n2748 0.135917
R4868 VDDA.n2760 VDDA.n193 0.135917
R4869 VDDA.n275 VDDA.n272 0.135917
R4870 VDDA.n279 VDDA.n259 0.135917
R4871 VDDA.n287 VDDA.n255 0.135917
R4872 VDDA.n291 VDDA.n288 0.135917
R4873 VDDA.n299 VDDA.n296 0.135917
R4874 VDDA.n303 VDDA.n247 0.135917
R4875 VDDA.n311 VDDA.n243 0.135917
R4876 VDDA.n315 VDDA.n312 0.135917
R4877 VDDA.n323 VDDA.n320 0.135917
R4878 VDDA.n327 VDDA.n235 0.135917
R4879 VDDA.n335 VDDA.n231 0.135917
R4880 VDDA.n339 VDDA.n336 0.135917
R4881 VDDA.n347 VDDA.n344 0.135917
R4882 VDDA.n351 VDDA.n223 0.135917
R4883 VDDA.n2596 VDDA.n221 0.135917
R4884 VDDA.n2478 VDDA.n2463 0.135917
R4885 VDDA.n2484 VDDA.n2461 0.135917
R4886 VDDA.n2494 VDDA.n2457 0.135917
R4887 VDDA.n2498 VDDA.n2455 0.135917
R4888 VDDA.n2508 VDDA.n2451 0.135917
R4889 VDDA.n2514 VDDA.n2449 0.135917
R4890 VDDA.n2524 VDDA.n2445 0.135917
R4891 VDDA.n2528 VDDA.n2443 0.135917
R4892 VDDA.n2538 VDDA.n2439 0.135917
R4893 VDDA.n2544 VDDA.n2437 0.135917
R4894 VDDA.n2554 VDDA.n2433 0.135917
R4895 VDDA.n2558 VDDA.n2431 0.135917
R4896 VDDA.n2568 VDDA.n2427 0.135917
R4897 VDDA.n2574 VDDA.n2425 0.135917
R4898 VDDA.n2583 VDDA.n2421 0.135917
R4899 VDDA.n1235 VDDA.n1221 0.135917
R4900 VDDA.n1239 VDDA.n1236 0.135917
R4901 VDDA.n1247 VDDA.n1244 0.135917
R4902 VDDA.n1251 VDDA.n1213 0.135917
R4903 VDDA.n1259 VDDA.n1209 0.135917
R4904 VDDA.n1263 VDDA.n1260 0.135917
R4905 VDDA.n1271 VDDA.n1268 0.135917
R4906 VDDA.n1275 VDDA.n1201 0.135917
R4907 VDDA.n1283 VDDA.n1197 0.135917
R4908 VDDA.n1287 VDDA.n1284 0.135917
R4909 VDDA.n1295 VDDA.n1292 0.135917
R4910 VDDA.n1299 VDDA.n1189 0.135917
R4911 VDDA.n1307 VDDA.n1185 0.135917
R4912 VDDA.n1311 VDDA.n1308 0.135917
R4913 VDDA.n2256 VDDA.n459 0.135917
R4914 VDDA.n541 VDDA.n538 0.135917
R4915 VDDA.n545 VDDA.n525 0.135917
R4916 VDDA.n553 VDDA.n521 0.135917
R4917 VDDA.n557 VDDA.n554 0.135917
R4918 VDDA.n565 VDDA.n562 0.135917
R4919 VDDA.n569 VDDA.n513 0.135917
R4920 VDDA.n577 VDDA.n509 0.135917
R4921 VDDA.n581 VDDA.n578 0.135917
R4922 VDDA.n589 VDDA.n586 0.135917
R4923 VDDA.n593 VDDA.n501 0.135917
R4924 VDDA.n601 VDDA.n497 0.135917
R4925 VDDA.n605 VDDA.n602 0.135917
R4926 VDDA.n613 VDDA.n610 0.135917
R4927 VDDA.n617 VDDA.n489 0.135917
R4928 VDDA.n1156 VDDA.n487 0.135917
R4929 VDDA.n1038 VDDA.n1023 0.135917
R4930 VDDA.n1044 VDDA.n1021 0.135917
R4931 VDDA.n1054 VDDA.n1017 0.135917
R4932 VDDA.n1058 VDDA.n1015 0.135917
R4933 VDDA.n1068 VDDA.n1011 0.135917
R4934 VDDA.n1074 VDDA.n1009 0.135917
R4935 VDDA.n1084 VDDA.n1005 0.135917
R4936 VDDA.n1088 VDDA.n1003 0.135917
R4937 VDDA.n1098 VDDA.n999 0.135917
R4938 VDDA.n1104 VDDA.n997 0.135917
R4939 VDDA.n1114 VDDA.n993 0.135917
R4940 VDDA.n1118 VDDA.n991 0.135917
R4941 VDDA.n1128 VDDA.n987 0.135917
R4942 VDDA.n1134 VDDA.n985 0.135917
R4943 VDDA.n1143 VDDA.n981 0.135917
R4944 VDDA.n887 VDDA.n873 0.135917
R4945 VDDA.n891 VDDA.n888 0.135917
R4946 VDDA.n899 VDDA.n896 0.135917
R4947 VDDA.n903 VDDA.n865 0.135917
R4948 VDDA.n911 VDDA.n861 0.135917
R4949 VDDA.n915 VDDA.n912 0.135917
R4950 VDDA.n923 VDDA.n920 0.135917
R4951 VDDA.n927 VDDA.n853 0.135917
R4952 VDDA.n935 VDDA.n849 0.135917
R4953 VDDA.n939 VDDA.n936 0.135917
R4954 VDDA.n947 VDDA.n944 0.135917
R4955 VDDA.n951 VDDA.n841 0.135917
R4956 VDDA.n959 VDDA.n837 0.135917
R4957 VDDA.n963 VDDA.n960 0.135917
R4958 VDDA.n972 VDDA.n636 0.135917
R4959 VDDA.n697 VDDA.n694 0.135917
R4960 VDDA.n703 VDDA.n683 0.135917
R4961 VDDA.n713 VDDA.n681 0.135917
R4962 VDDA.n717 VDDA.n714 0.135917
R4963 VDDA.n727 VDDA.n724 0.135917
R4964 VDDA.n733 VDDA.n677 0.135917
R4965 VDDA.n743 VDDA.n675 0.135917
R4966 VDDA.n747 VDDA.n744 0.135917
R4967 VDDA.n757 VDDA.n754 0.135917
R4968 VDDA.n763 VDDA.n671 0.135917
R4969 VDDA.n773 VDDA.n669 0.135917
R4970 VDDA.n777 VDDA.n774 0.135917
R4971 VDDA.n787 VDDA.n784 0.135917
R4972 VDDA.n793 VDDA.n665 0.135917
R4973 VDDA.n808 VDDA.n663 0.135917
R4974 VDDA.n1474 VDDA.n1453 0.1255
R4975 VDDA.n1491 VDDA.n1490 0.1255
R4976 VDDA.n1504 VDDA.n1447 0.1255
R4977 VDDA.n1521 VDDA.n1520 0.1255
R4978 VDDA.n1534 VDDA.n1441 0.1255
R4979 VDDA.n1551 VDDA.n1550 0.1255
R4980 VDDA.n1564 VDDA.n1435 0.1255
R4981 VDDA.n2129 VDDA.n2128 0.1255
R4982 VDDA.n2128 VDDA.n2127 0.1255
R4983 VDDA.n2002 VDDA.n1950 0.1255
R4984 VDDA.n1953 VDDA.n1950 0.1255
R4985 VDDA.n1955 VDDA.n1953 0.1255
R4986 VDDA.n1957 VDDA.n1955 0.1255
R4987 VDDA.n1959 VDDA.n1957 0.1255
R4988 VDDA.n1961 VDDA.n1959 0.1255
R4989 VDDA.n1963 VDDA.n1961 0.1255
R4990 VDDA.n1965 VDDA.n1963 0.1255
R4991 VDDA.n1967 VDDA.n1965 0.1255
R4992 VDDA.n1996 VDDA.n1967 0.1255
R4993 VDDA.n1995 VDDA.n1969 0.1255
R4994 VDDA.n1973 VDDA.n1969 0.1255
R4995 VDDA.n1975 VDDA.n1973 0.1255
R4996 VDDA.n1977 VDDA.n1975 0.1255
R4997 VDDA.n1979 VDDA.n1977 0.1255
R4998 VDDA.n1981 VDDA.n1979 0.1255
R4999 VDDA.n1983 VDDA.n1981 0.1255
R5000 VDDA.n1985 VDDA.n1983 0.1255
R5001 VDDA.n1987 VDDA.n1985 0.1255
R5002 VDDA.n2149 VDDA.n1928 0.1255
R5003 VDDA.n2166 VDDA.n2165 0.1255
R5004 VDDA.n2179 VDDA.n1922 0.1255
R5005 VDDA.n2196 VDDA.n2195 0.1255
R5006 VDDA.n2209 VDDA.n1916 0.1255
R5007 VDDA.n2226 VDDA.n2225 0.1255
R5008 VDDA.n2239 VDDA.n1910 0.1255
R5009 VDDA.n97 VDDA.n81 0.1255
R5010 VDDA.n110 VDDA.n109 0.1255
R5011 VDDA.n121 VDDA.n69 0.1255
R5012 VDDA.n134 VDDA.n133 0.1255
R5013 VDDA.n145 VDDA.n57 0.1255
R5014 VDDA.n158 VDDA.n157 0.1255
R5015 VDDA.n169 VDDA.n45 0.1255
R5016 VDDA.n2826 VDDA.n2809 0.1255
R5017 VDDA.n2842 VDDA.n2803 0.1255
R5018 VDDA.n2856 VDDA.n2797 0.1255
R5019 VDDA.n2872 VDDA.n2791 0.1255
R5020 VDDA.n2886 VDDA.n2785 0.1255
R5021 VDDA.n2902 VDDA.n2779 0.1255
R5022 VDDA.n2916 VDDA.n2773 0.1255
R5023 VDDA.n2676 VDDA.n2675 0.1255
R5024 VDDA.n2687 VDDA.n2653 0.1255
R5025 VDDA.n2700 VDDA.n2699 0.1255
R5026 VDDA.n2711 VDDA.n2641 0.1255
R5027 VDDA.n2724 VDDA.n2723 0.1255
R5028 VDDA.n2735 VDDA.n2629 0.1255
R5029 VDDA.n2748 VDDA.n2747 0.1255
R5030 VDDA.n275 VDDA.n259 0.1255
R5031 VDDA.n288 VDDA.n287 0.1255
R5032 VDDA.n299 VDDA.n247 0.1255
R5033 VDDA.n312 VDDA.n311 0.1255
R5034 VDDA.n323 VDDA.n235 0.1255
R5035 VDDA.n336 VDDA.n335 0.1255
R5036 VDDA.n347 VDDA.n223 0.1255
R5037 VDDA.n2478 VDDA.n2461 0.1255
R5038 VDDA.n2494 VDDA.n2455 0.1255
R5039 VDDA.n2508 VDDA.n2449 0.1255
R5040 VDDA.n2524 VDDA.n2443 0.1255
R5041 VDDA.n2538 VDDA.n2437 0.1255
R5042 VDDA.n2554 VDDA.n2431 0.1255
R5043 VDDA.n2568 VDDA.n2425 0.1255
R5044 VDDA.n1236 VDDA.n1235 0.1255
R5045 VDDA.n1247 VDDA.n1213 0.1255
R5046 VDDA.n1260 VDDA.n1259 0.1255
R5047 VDDA.n1271 VDDA.n1201 0.1255
R5048 VDDA.n1284 VDDA.n1283 0.1255
R5049 VDDA.n1295 VDDA.n1189 0.1255
R5050 VDDA.n1308 VDDA.n1307 0.1255
R5051 VDDA.n375 VDDA.n370 0.1255
R5052 VDDA.n382 VDDA.n376 0.1255
R5053 VDDA.n541 VDDA.n525 0.1255
R5054 VDDA.n554 VDDA.n553 0.1255
R5055 VDDA.n565 VDDA.n513 0.1255
R5056 VDDA.n578 VDDA.n577 0.1255
R5057 VDDA.n589 VDDA.n501 0.1255
R5058 VDDA.n602 VDDA.n601 0.1255
R5059 VDDA.n613 VDDA.n489 0.1255
R5060 VDDA.n1038 VDDA.n1021 0.1255
R5061 VDDA.n1054 VDDA.n1015 0.1255
R5062 VDDA.n1068 VDDA.n1009 0.1255
R5063 VDDA.n1084 VDDA.n1003 0.1255
R5064 VDDA.n1098 VDDA.n997 0.1255
R5065 VDDA.n1114 VDDA.n991 0.1255
R5066 VDDA.n1128 VDDA.n985 0.1255
R5067 VDDA.n888 VDDA.n887 0.1255
R5068 VDDA.n899 VDDA.n865 0.1255
R5069 VDDA.n912 VDDA.n911 0.1255
R5070 VDDA.n923 VDDA.n853 0.1255
R5071 VDDA.n936 VDDA.n935 0.1255
R5072 VDDA.n947 VDDA.n841 0.1255
R5073 VDDA.n960 VDDA.n959 0.1255
R5074 VDDA.n697 VDDA.n683 0.1255
R5075 VDDA.n714 VDDA.n713 0.1255
R5076 VDDA.n727 VDDA.n677 0.1255
R5077 VDDA.n744 VDDA.n743 0.1255
R5078 VDDA.n757 VDDA.n671 0.1255
R5079 VDDA.n774 VDDA.n773 0.1255
R5080 VDDA.n787 VDDA.n665 0.1255
R5081 VDDA.n1766 VDDA.n1765 0.123287
R5082 VDDA.n1788 VDDA.n1787 0.123287
R5083 VDDA.n2126 VDDA.n2125 0.115083
R5084 VDDA.n2125 VDDA.n2124 0.115083
R5085 VDDA.n2124 VDDA.n2123 0.115083
R5086 VDDA.n2121 VDDA.n2120 0.115083
R5087 VDDA.n2120 VDDA.n2119 0.115083
R5088 VDDA.n2119 VDDA.n2118 0.115083
R5089 VDDA.n2118 VDDA.n2117 0.115083
R5090 VDDA.n2115 VDDA.n2114 0.115083
R5091 VDDA.n2114 VDDA.n2113 0.115083
R5092 VDDA.n2313 VDDA.n2311 0.115083
R5093 VDDA.n2315 VDDA.n2313 0.115083
R5094 VDDA.n2317 VDDA.n2315 0.115083
R5095 VDDA.n2319 VDDA.n2317 0.115083
R5096 VDDA.n423 VDDA.n421 0.115083
R5097 VDDA.n421 VDDA.n419 0.115083
R5098 VDDA.n419 VDDA.n417 0.115083
R5099 VDDA.n417 VDDA.n415 0.115083
R5100 VDDA.n2297 VDDA.n2295 0.115083
R5101 VDDA.n2295 VDDA.n2293 0.115083
R5102 VDDA.n2293 VDDA.n2291 0.115083
R5103 VDDA.n2291 VDDA.n2289 0.115083
R5104 VDDA.n2302 VDDA.n2289 0.115083
R5105 VDDA.n403 VDDA.n390 0.115083
R5106 VDDA.n392 VDDA.n390 0.115083
R5107 VDDA.n394 VDDA.n392 0.115083
R5108 VDDA.n396 VDDA.n394 0.115083
R5109 VDDA.n398 VDDA.n396 0.115083
R5110 VDDA.n2362 VDDA.n2361 0.0838333
R5111 VDDA.n1761 VDDA.n1405 0.076587
R5112 VDDA.n1580 VDDA.n1405 0.076587
R5113 VDDA.n1753 VDDA.n1580 0.076587
R5114 VDDA.n1743 VDDA.n1585 0.076587
R5115 VDDA.n1743 VDDA.n1589 0.076587
R5116 VDDA.n1739 VDDA.n1589 0.076587
R5117 VDDA.n1729 VDDA.n1595 0.076587
R5118 VDDA.n1729 VDDA.n1597 0.076587
R5119 VDDA.n1723 VDDA.n1597 0.076587
R5120 VDDA.n1713 VDDA.n1603 0.076587
R5121 VDDA.n1713 VDDA.n1607 0.076587
R5122 VDDA.n1709 VDDA.n1607 0.076587
R5123 VDDA.n1699 VDDA.n1613 0.076587
R5124 VDDA.n1699 VDDA.n1615 0.076587
R5125 VDDA.n1693 VDDA.n1615 0.076587
R5126 VDDA.n1683 VDDA.n1621 0.076587
R5127 VDDA.n1683 VDDA.n1625 0.076587
R5128 VDDA.n1679 VDDA.n1625 0.076587
R5129 VDDA.n1669 VDDA.n1631 0.076587
R5130 VDDA.n1669 VDDA.n1633 0.076587
R5131 VDDA.n1663 VDDA.n1633 0.076587
R5132 VDDA.n1653 VDDA.n1639 0.076587
R5133 VDDA.n1653 VDDA.n1643 0.076587
R5134 VDDA.n1649 VDDA.n1643 0.076587
R5135 VDDA.n1762 VDDA.n1404 0.076587
R5136 VDDA.n1583 VDDA.n1404 0.076587
R5137 VDDA.n1752 VDDA.n1583 0.076587
R5138 VDDA.n1742 VDDA.n1584 0.076587
R5139 VDDA.n1742 VDDA.n1741 0.076587
R5140 VDDA.n1741 VDDA.n1740 0.076587
R5141 VDDA.n1731 VDDA.n1730 0.076587
R5142 VDDA.n1730 VDDA.n1596 0.076587
R5143 VDDA.n1722 VDDA.n1596 0.076587
R5144 VDDA.n1712 VDDA.n1602 0.076587
R5145 VDDA.n1712 VDDA.n1711 0.076587
R5146 VDDA.n1711 VDDA.n1710 0.076587
R5147 VDDA.n1701 VDDA.n1700 0.076587
R5148 VDDA.n1700 VDDA.n1614 0.076587
R5149 VDDA.n1692 VDDA.n1614 0.076587
R5150 VDDA.n1682 VDDA.n1620 0.076587
R5151 VDDA.n1682 VDDA.n1681 0.076587
R5152 VDDA.n1681 VDDA.n1680 0.076587
R5153 VDDA.n1671 VDDA.n1670 0.076587
R5154 VDDA.n1670 VDDA.n1632 0.076587
R5155 VDDA.n1662 VDDA.n1632 0.076587
R5156 VDDA.n1652 VDDA.n1638 0.076587
R5157 VDDA.n1652 VDDA.n1651 0.076587
R5158 VDDA.n1904 VDDA.n1368 0.0751758
R5159 VDDA.n1466 VDDA.n1465 0.0734167
R5160 VDDA.n1467 VDDA.n1466 0.0734167
R5161 VDDA.n1467 VDDA.n1454 0.0734167
R5162 VDDA.n1477 VDDA.n1452 0.0734167
R5163 VDDA.n1485 VDDA.n1452 0.0734167
R5164 VDDA.n1486 VDDA.n1485 0.0734167
R5165 VDDA.n1496 VDDA.n1495 0.0734167
R5166 VDDA.n1497 VDDA.n1496 0.0734167
R5167 VDDA.n1497 VDDA.n1448 0.0734167
R5168 VDDA.n1507 VDDA.n1446 0.0734167
R5169 VDDA.n1515 VDDA.n1446 0.0734167
R5170 VDDA.n1516 VDDA.n1515 0.0734167
R5171 VDDA.n1526 VDDA.n1525 0.0734167
R5172 VDDA.n1527 VDDA.n1526 0.0734167
R5173 VDDA.n1527 VDDA.n1442 0.0734167
R5174 VDDA.n1537 VDDA.n1440 0.0734167
R5175 VDDA.n1545 VDDA.n1440 0.0734167
R5176 VDDA.n1546 VDDA.n1545 0.0734167
R5177 VDDA.n1556 VDDA.n1555 0.0734167
R5178 VDDA.n1557 VDDA.n1556 0.0734167
R5179 VDDA.n1557 VDDA.n1436 0.0734167
R5180 VDDA.n1567 VDDA.n1434 0.0734167
R5181 VDDA.n1575 VDDA.n1434 0.0734167
R5182 VDDA.n2141 VDDA.n2140 0.0734167
R5183 VDDA.n2142 VDDA.n2141 0.0734167
R5184 VDDA.n2142 VDDA.n1929 0.0734167
R5185 VDDA.n2152 VDDA.n1927 0.0734167
R5186 VDDA.n2160 VDDA.n1927 0.0734167
R5187 VDDA.n2161 VDDA.n2160 0.0734167
R5188 VDDA.n2171 VDDA.n2170 0.0734167
R5189 VDDA.n2172 VDDA.n2171 0.0734167
R5190 VDDA.n2172 VDDA.n1923 0.0734167
R5191 VDDA.n2182 VDDA.n1921 0.0734167
R5192 VDDA.n2190 VDDA.n1921 0.0734167
R5193 VDDA.n2191 VDDA.n2190 0.0734167
R5194 VDDA.n2201 VDDA.n2200 0.0734167
R5195 VDDA.n2202 VDDA.n2201 0.0734167
R5196 VDDA.n2202 VDDA.n1917 0.0734167
R5197 VDDA.n2212 VDDA.n1915 0.0734167
R5198 VDDA.n2220 VDDA.n1915 0.0734167
R5199 VDDA.n2221 VDDA.n2220 0.0734167
R5200 VDDA.n2231 VDDA.n2230 0.0734167
R5201 VDDA.n2232 VDDA.n2231 0.0734167
R5202 VDDA.n2232 VDDA.n1911 0.0734167
R5203 VDDA.n2242 VDDA.n1909 0.0734167
R5204 VDDA.n2250 VDDA.n1909 0.0734167
R5205 VDDA.n92 VDDA.n91 0.0734167
R5206 VDDA.n92 VDDA.n84 0.0734167
R5207 VDDA.n100 VDDA.n80 0.0734167
R5208 VDDA.n106 VDDA.n80 0.0734167
R5209 VDDA.n107 VDDA.n106 0.0734167
R5210 VDDA.n115 VDDA.n114 0.0734167
R5211 VDDA.n116 VDDA.n115 0.0734167
R5212 VDDA.n116 VDDA.n72 0.0734167
R5213 VDDA.n124 VDDA.n68 0.0734167
R5214 VDDA.n130 VDDA.n68 0.0734167
R5215 VDDA.n131 VDDA.n130 0.0734167
R5216 VDDA.n139 VDDA.n138 0.0734167
R5217 VDDA.n140 VDDA.n139 0.0734167
R5218 VDDA.n140 VDDA.n60 0.0734167
R5219 VDDA.n148 VDDA.n56 0.0734167
R5220 VDDA.n154 VDDA.n56 0.0734167
R5221 VDDA.n155 VDDA.n154 0.0734167
R5222 VDDA.n163 VDDA.n162 0.0734167
R5223 VDDA.n164 VDDA.n163 0.0734167
R5224 VDDA.n164 VDDA.n48 0.0734167
R5225 VDDA.n172 VDDA.n44 0.0734167
R5226 VDDA.n178 VDDA.n44 0.0734167
R5227 VDDA.n179 VDDA.n178 0.0734167
R5228 VDDA.n2823 VDDA.n2812 0.0734167
R5229 VDDA.n2824 VDDA.n2823 0.0734167
R5230 VDDA.n2834 VDDA.n2833 0.0734167
R5231 VDDA.n2835 VDDA.n2834 0.0734167
R5232 VDDA.n2835 VDDA.n2804 0.0734167
R5233 VDDA.n2845 VDDA.n2800 0.0734167
R5234 VDDA.n2853 VDDA.n2800 0.0734167
R5235 VDDA.n2854 VDDA.n2853 0.0734167
R5236 VDDA.n2864 VDDA.n2863 0.0734167
R5237 VDDA.n2865 VDDA.n2864 0.0734167
R5238 VDDA.n2865 VDDA.n2792 0.0734167
R5239 VDDA.n2875 VDDA.n2788 0.0734167
R5240 VDDA.n2883 VDDA.n2788 0.0734167
R5241 VDDA.n2884 VDDA.n2883 0.0734167
R5242 VDDA.n2894 VDDA.n2893 0.0734167
R5243 VDDA.n2895 VDDA.n2894 0.0734167
R5244 VDDA.n2895 VDDA.n2780 0.0734167
R5245 VDDA.n2905 VDDA.n2776 0.0734167
R5246 VDDA.n2913 VDDA.n2776 0.0734167
R5247 VDDA.n2914 VDDA.n2913 0.0734167
R5248 VDDA.n2924 VDDA.n2923 0.0734167
R5249 VDDA.n2925 VDDA.n2924 0.0734167
R5250 VDDA.n2925 VDDA.n2768 0.0734167
R5251 VDDA.n2672 VDDA.n2664 0.0734167
R5252 VDDA.n2673 VDDA.n2672 0.0734167
R5253 VDDA.n2681 VDDA.n2680 0.0734167
R5254 VDDA.n2682 VDDA.n2681 0.0734167
R5255 VDDA.n2682 VDDA.n2656 0.0734167
R5256 VDDA.n2690 VDDA.n2652 0.0734167
R5257 VDDA.n2696 VDDA.n2652 0.0734167
R5258 VDDA.n2697 VDDA.n2696 0.0734167
R5259 VDDA.n2705 VDDA.n2704 0.0734167
R5260 VDDA.n2706 VDDA.n2705 0.0734167
R5261 VDDA.n2706 VDDA.n2644 0.0734167
R5262 VDDA.n2714 VDDA.n2640 0.0734167
R5263 VDDA.n2720 VDDA.n2640 0.0734167
R5264 VDDA.n2721 VDDA.n2720 0.0734167
R5265 VDDA.n2729 VDDA.n2728 0.0734167
R5266 VDDA.n2730 VDDA.n2729 0.0734167
R5267 VDDA.n2730 VDDA.n2632 0.0734167
R5268 VDDA.n2738 VDDA.n2628 0.0734167
R5269 VDDA.n2744 VDDA.n2628 0.0734167
R5270 VDDA.n2745 VDDA.n2744 0.0734167
R5271 VDDA.n2753 VDDA.n2752 0.0734167
R5272 VDDA.n2754 VDDA.n2753 0.0734167
R5273 VDDA.n2754 VDDA.n192 0.0734167
R5274 VDDA.n270 VDDA.n269 0.0734167
R5275 VDDA.n270 VDDA.n262 0.0734167
R5276 VDDA.n278 VDDA.n258 0.0734167
R5277 VDDA.n284 VDDA.n258 0.0734167
R5278 VDDA.n285 VDDA.n284 0.0734167
R5279 VDDA.n293 VDDA.n292 0.0734167
R5280 VDDA.n294 VDDA.n293 0.0734167
R5281 VDDA.n294 VDDA.n250 0.0734167
R5282 VDDA.n302 VDDA.n246 0.0734167
R5283 VDDA.n308 VDDA.n246 0.0734167
R5284 VDDA.n309 VDDA.n308 0.0734167
R5285 VDDA.n317 VDDA.n316 0.0734167
R5286 VDDA.n318 VDDA.n317 0.0734167
R5287 VDDA.n318 VDDA.n238 0.0734167
R5288 VDDA.n326 VDDA.n234 0.0734167
R5289 VDDA.n332 VDDA.n234 0.0734167
R5290 VDDA.n333 VDDA.n332 0.0734167
R5291 VDDA.n341 VDDA.n340 0.0734167
R5292 VDDA.n342 VDDA.n341 0.0734167
R5293 VDDA.n342 VDDA.n226 0.0734167
R5294 VDDA.n350 VDDA.n222 0.0734167
R5295 VDDA.n356 VDDA.n222 0.0734167
R5296 VDDA.n357 VDDA.n356 0.0734167
R5297 VDDA.n2475 VDDA.n2464 0.0734167
R5298 VDDA.n2476 VDDA.n2475 0.0734167
R5299 VDDA.n2486 VDDA.n2485 0.0734167
R5300 VDDA.n2487 VDDA.n2486 0.0734167
R5301 VDDA.n2487 VDDA.n2456 0.0734167
R5302 VDDA.n2497 VDDA.n2452 0.0734167
R5303 VDDA.n2505 VDDA.n2452 0.0734167
R5304 VDDA.n2506 VDDA.n2505 0.0734167
R5305 VDDA.n2516 VDDA.n2515 0.0734167
R5306 VDDA.n2517 VDDA.n2516 0.0734167
R5307 VDDA.n2517 VDDA.n2444 0.0734167
R5308 VDDA.n2527 VDDA.n2440 0.0734167
R5309 VDDA.n2535 VDDA.n2440 0.0734167
R5310 VDDA.n2536 VDDA.n2535 0.0734167
R5311 VDDA.n2546 VDDA.n2545 0.0734167
R5312 VDDA.n2547 VDDA.n2546 0.0734167
R5313 VDDA.n2547 VDDA.n2432 0.0734167
R5314 VDDA.n2557 VDDA.n2428 0.0734167
R5315 VDDA.n2565 VDDA.n2428 0.0734167
R5316 VDDA.n2566 VDDA.n2565 0.0734167
R5317 VDDA.n2576 VDDA.n2575 0.0734167
R5318 VDDA.n2577 VDDA.n2576 0.0734167
R5319 VDDA.n2577 VDDA.n2420 0.0734167
R5320 VDDA.n1232 VDDA.n1224 0.0734167
R5321 VDDA.n1233 VDDA.n1232 0.0734167
R5322 VDDA.n1241 VDDA.n1240 0.0734167
R5323 VDDA.n1242 VDDA.n1241 0.0734167
R5324 VDDA.n1242 VDDA.n1216 0.0734167
R5325 VDDA.n1250 VDDA.n1212 0.0734167
R5326 VDDA.n1256 VDDA.n1212 0.0734167
R5327 VDDA.n1257 VDDA.n1256 0.0734167
R5328 VDDA.n1265 VDDA.n1264 0.0734167
R5329 VDDA.n1266 VDDA.n1265 0.0734167
R5330 VDDA.n1266 VDDA.n1204 0.0734167
R5331 VDDA.n1274 VDDA.n1200 0.0734167
R5332 VDDA.n1280 VDDA.n1200 0.0734167
R5333 VDDA.n1281 VDDA.n1280 0.0734167
R5334 VDDA.n1289 VDDA.n1288 0.0734167
R5335 VDDA.n1290 VDDA.n1289 0.0734167
R5336 VDDA.n1290 VDDA.n1192 0.0734167
R5337 VDDA.n1298 VDDA.n1188 0.0734167
R5338 VDDA.n1304 VDDA.n1188 0.0734167
R5339 VDDA.n1305 VDDA.n1304 0.0734167
R5340 VDDA.n1313 VDDA.n1312 0.0734167
R5341 VDDA.n1314 VDDA.n1313 0.0734167
R5342 VDDA.n1314 VDDA.n458 0.0734167
R5343 VDDA.n536 VDDA.n535 0.0734167
R5344 VDDA.n536 VDDA.n528 0.0734167
R5345 VDDA.n544 VDDA.n524 0.0734167
R5346 VDDA.n550 VDDA.n524 0.0734167
R5347 VDDA.n551 VDDA.n550 0.0734167
R5348 VDDA.n559 VDDA.n558 0.0734167
R5349 VDDA.n560 VDDA.n559 0.0734167
R5350 VDDA.n560 VDDA.n516 0.0734167
R5351 VDDA.n568 VDDA.n512 0.0734167
R5352 VDDA.n574 VDDA.n512 0.0734167
R5353 VDDA.n575 VDDA.n574 0.0734167
R5354 VDDA.n583 VDDA.n582 0.0734167
R5355 VDDA.n584 VDDA.n583 0.0734167
R5356 VDDA.n584 VDDA.n504 0.0734167
R5357 VDDA.n592 VDDA.n500 0.0734167
R5358 VDDA.n598 VDDA.n500 0.0734167
R5359 VDDA.n599 VDDA.n598 0.0734167
R5360 VDDA.n607 VDDA.n606 0.0734167
R5361 VDDA.n608 VDDA.n607 0.0734167
R5362 VDDA.n608 VDDA.n492 0.0734167
R5363 VDDA.n616 VDDA.n488 0.0734167
R5364 VDDA.n622 VDDA.n488 0.0734167
R5365 VDDA.n623 VDDA.n622 0.0734167
R5366 VDDA.n1035 VDDA.n1024 0.0734167
R5367 VDDA.n1036 VDDA.n1035 0.0734167
R5368 VDDA.n1046 VDDA.n1045 0.0734167
R5369 VDDA.n1047 VDDA.n1046 0.0734167
R5370 VDDA.n1047 VDDA.n1016 0.0734167
R5371 VDDA.n1057 VDDA.n1012 0.0734167
R5372 VDDA.n1065 VDDA.n1012 0.0734167
R5373 VDDA.n1066 VDDA.n1065 0.0734167
R5374 VDDA.n1076 VDDA.n1075 0.0734167
R5375 VDDA.n1077 VDDA.n1076 0.0734167
R5376 VDDA.n1077 VDDA.n1004 0.0734167
R5377 VDDA.n1087 VDDA.n1000 0.0734167
R5378 VDDA.n1095 VDDA.n1000 0.0734167
R5379 VDDA.n1096 VDDA.n1095 0.0734167
R5380 VDDA.n1106 VDDA.n1105 0.0734167
R5381 VDDA.n1107 VDDA.n1106 0.0734167
R5382 VDDA.n1107 VDDA.n992 0.0734167
R5383 VDDA.n1117 VDDA.n988 0.0734167
R5384 VDDA.n1125 VDDA.n988 0.0734167
R5385 VDDA.n1126 VDDA.n1125 0.0734167
R5386 VDDA.n1136 VDDA.n1135 0.0734167
R5387 VDDA.n1137 VDDA.n1136 0.0734167
R5388 VDDA.n1137 VDDA.n980 0.0734167
R5389 VDDA.n884 VDDA.n876 0.0734167
R5390 VDDA.n885 VDDA.n884 0.0734167
R5391 VDDA.n893 VDDA.n892 0.0734167
R5392 VDDA.n894 VDDA.n893 0.0734167
R5393 VDDA.n894 VDDA.n868 0.0734167
R5394 VDDA.n902 VDDA.n864 0.0734167
R5395 VDDA.n908 VDDA.n864 0.0734167
R5396 VDDA.n909 VDDA.n908 0.0734167
R5397 VDDA.n917 VDDA.n916 0.0734167
R5398 VDDA.n918 VDDA.n917 0.0734167
R5399 VDDA.n918 VDDA.n856 0.0734167
R5400 VDDA.n926 VDDA.n852 0.0734167
R5401 VDDA.n932 VDDA.n852 0.0734167
R5402 VDDA.n933 VDDA.n932 0.0734167
R5403 VDDA.n941 VDDA.n940 0.0734167
R5404 VDDA.n942 VDDA.n941 0.0734167
R5405 VDDA.n942 VDDA.n844 0.0734167
R5406 VDDA.n950 VDDA.n840 0.0734167
R5407 VDDA.n956 VDDA.n840 0.0734167
R5408 VDDA.n957 VDDA.n956 0.0734167
R5409 VDDA.n965 VDDA.n964 0.0734167
R5410 VDDA.n966 VDDA.n965 0.0734167
R5411 VDDA.n966 VDDA.n635 0.0734167
R5412 VDDA.n690 VDDA.n689 0.0734167
R5413 VDDA.n690 VDDA.n684 0.0734167
R5414 VDDA.n700 VDDA.n682 0.0734167
R5415 VDDA.n708 VDDA.n682 0.0734167
R5416 VDDA.n709 VDDA.n708 0.0734167
R5417 VDDA.n719 VDDA.n718 0.0734167
R5418 VDDA.n720 VDDA.n719 0.0734167
R5419 VDDA.n720 VDDA.n678 0.0734167
R5420 VDDA.n730 VDDA.n676 0.0734167
R5421 VDDA.n738 VDDA.n676 0.0734167
R5422 VDDA.n739 VDDA.n738 0.0734167
R5423 VDDA.n749 VDDA.n748 0.0734167
R5424 VDDA.n750 VDDA.n749 0.0734167
R5425 VDDA.n750 VDDA.n672 0.0734167
R5426 VDDA.n760 VDDA.n670 0.0734167
R5427 VDDA.n768 VDDA.n670 0.0734167
R5428 VDDA.n769 VDDA.n768 0.0734167
R5429 VDDA.n779 VDDA.n778 0.0734167
R5430 VDDA.n780 VDDA.n779 0.0734167
R5431 VDDA.n780 VDDA.n666 0.0734167
R5432 VDDA.n790 VDDA.n664 0.0734167
R5433 VDDA.n798 VDDA.n664 0.0734167
R5434 VDDA.n799 VDDA.n798 0.0734167
R5435 VDDA.n1761 VDDA.n1403 0.0711522
R5436 VDDA.n1753 VDDA.n1582 0.0711522
R5437 VDDA.n1749 VDDA.n1585 0.0711522
R5438 VDDA.n1739 VDDA.n1591 0.0711522
R5439 VDDA.n1733 VDDA.n1595 0.0711522
R5440 VDDA.n1723 VDDA.n1601 0.0711522
R5441 VDDA.n1719 VDDA.n1603 0.0711522
R5442 VDDA.n1709 VDDA.n1609 0.0711522
R5443 VDDA.n1703 VDDA.n1613 0.0711522
R5444 VDDA.n1693 VDDA.n1619 0.0711522
R5445 VDDA.n1689 VDDA.n1621 0.0711522
R5446 VDDA.n1679 VDDA.n1627 0.0711522
R5447 VDDA.n1673 VDDA.n1631 0.0711522
R5448 VDDA.n1663 VDDA.n1637 0.0711522
R5449 VDDA.n1659 VDDA.n1639 0.0711522
R5450 VDDA.n1763 VDDA.n1762 0.0711522
R5451 VDDA.n1752 VDDA.n1751 0.0711522
R5452 VDDA.n1750 VDDA.n1584 0.0711522
R5453 VDDA.n1740 VDDA.n1590 0.0711522
R5454 VDDA.n1732 VDDA.n1731 0.0711522
R5455 VDDA.n1722 VDDA.n1721 0.0711522
R5456 VDDA.n1720 VDDA.n1602 0.0711522
R5457 VDDA.n1710 VDDA.n1608 0.0711522
R5458 VDDA.n1702 VDDA.n1701 0.0711522
R5459 VDDA.n1692 VDDA.n1691 0.0711522
R5460 VDDA.n1690 VDDA.n1620 0.0711522
R5461 VDDA.n1680 VDDA.n1626 0.0711522
R5462 VDDA.n1672 VDDA.n1671 0.0711522
R5463 VDDA.n1662 VDDA.n1661 0.0711522
R5464 VDDA.n1660 VDDA.n1638 0.0711522
R5465 VDDA.n1465 VDDA.n1461 0.0682083
R5466 VDDA.n1475 VDDA.n1454 0.0682083
R5467 VDDA.n1477 VDDA.n1476 0.0682083
R5468 VDDA.n1487 VDDA.n1486 0.0682083
R5469 VDDA.n1495 VDDA.n1450 0.0682083
R5470 VDDA.n1505 VDDA.n1448 0.0682083
R5471 VDDA.n1507 VDDA.n1506 0.0682083
R5472 VDDA.n1517 VDDA.n1516 0.0682083
R5473 VDDA.n1525 VDDA.n1444 0.0682083
R5474 VDDA.n1535 VDDA.n1442 0.0682083
R5475 VDDA.n1537 VDDA.n1536 0.0682083
R5476 VDDA.n1547 VDDA.n1546 0.0682083
R5477 VDDA.n1555 VDDA.n1438 0.0682083
R5478 VDDA.n1565 VDDA.n1436 0.0682083
R5479 VDDA.n1567 VDDA.n1566 0.0682083
R5480 VDDA.n2122 VDDA.n2121 0.0682083
R5481 VDDA.n2117 VDDA.n2116 0.0682083
R5482 VDDA.n2140 VDDA.n2136 0.0682083
R5483 VDDA.n2150 VDDA.n1929 0.0682083
R5484 VDDA.n2152 VDDA.n2151 0.0682083
R5485 VDDA.n2162 VDDA.n2161 0.0682083
R5486 VDDA.n2170 VDDA.n1925 0.0682083
R5487 VDDA.n2180 VDDA.n1923 0.0682083
R5488 VDDA.n2182 VDDA.n2181 0.0682083
R5489 VDDA.n2192 VDDA.n2191 0.0682083
R5490 VDDA.n2200 VDDA.n1919 0.0682083
R5491 VDDA.n2210 VDDA.n1917 0.0682083
R5492 VDDA.n2212 VDDA.n2211 0.0682083
R5493 VDDA.n2222 VDDA.n2221 0.0682083
R5494 VDDA.n2230 VDDA.n1913 0.0682083
R5495 VDDA.n2240 VDDA.n1911 0.0682083
R5496 VDDA.n2242 VDDA.n2241 0.0682083
R5497 VDDA.n98 VDDA.n84 0.0682083
R5498 VDDA.n100 VDDA.n99 0.0682083
R5499 VDDA.n108 VDDA.n107 0.0682083
R5500 VDDA.n114 VDDA.n76 0.0682083
R5501 VDDA.n122 VDDA.n72 0.0682083
R5502 VDDA.n124 VDDA.n123 0.0682083
R5503 VDDA.n132 VDDA.n131 0.0682083
R5504 VDDA.n138 VDDA.n64 0.0682083
R5505 VDDA.n146 VDDA.n60 0.0682083
R5506 VDDA.n148 VDDA.n147 0.0682083
R5507 VDDA.n156 VDDA.n155 0.0682083
R5508 VDDA.n162 VDDA.n52 0.0682083
R5509 VDDA.n170 VDDA.n48 0.0682083
R5510 VDDA.n172 VDDA.n171 0.0682083
R5511 VDDA.n2943 VDDA.n179 0.0682083
R5512 VDDA.n2825 VDDA.n2824 0.0682083
R5513 VDDA.n2833 VDDA.n2808 0.0682083
R5514 VDDA.n2843 VDDA.n2804 0.0682083
R5515 VDDA.n2845 VDDA.n2844 0.0682083
R5516 VDDA.n2855 VDDA.n2854 0.0682083
R5517 VDDA.n2863 VDDA.n2796 0.0682083
R5518 VDDA.n2873 VDDA.n2792 0.0682083
R5519 VDDA.n2875 VDDA.n2874 0.0682083
R5520 VDDA.n2885 VDDA.n2884 0.0682083
R5521 VDDA.n2893 VDDA.n2784 0.0682083
R5522 VDDA.n2903 VDDA.n2780 0.0682083
R5523 VDDA.n2905 VDDA.n2904 0.0682083
R5524 VDDA.n2915 VDDA.n2914 0.0682083
R5525 VDDA.n2923 VDDA.n2772 0.0682083
R5526 VDDA.n2932 VDDA.n2768 0.0682083
R5527 VDDA.n2674 VDDA.n2673 0.0682083
R5528 VDDA.n2680 VDDA.n2660 0.0682083
R5529 VDDA.n2688 VDDA.n2656 0.0682083
R5530 VDDA.n2690 VDDA.n2689 0.0682083
R5531 VDDA.n2698 VDDA.n2697 0.0682083
R5532 VDDA.n2704 VDDA.n2648 0.0682083
R5533 VDDA.n2712 VDDA.n2644 0.0682083
R5534 VDDA.n2714 VDDA.n2713 0.0682083
R5535 VDDA.n2722 VDDA.n2721 0.0682083
R5536 VDDA.n2728 VDDA.n2636 0.0682083
R5537 VDDA.n2736 VDDA.n2632 0.0682083
R5538 VDDA.n2738 VDDA.n2737 0.0682083
R5539 VDDA.n2746 VDDA.n2745 0.0682083
R5540 VDDA.n2752 VDDA.n2624 0.0682083
R5541 VDDA.n2761 VDDA.n192 0.0682083
R5542 VDDA.n276 VDDA.n262 0.0682083
R5543 VDDA.n278 VDDA.n277 0.0682083
R5544 VDDA.n286 VDDA.n285 0.0682083
R5545 VDDA.n292 VDDA.n254 0.0682083
R5546 VDDA.n300 VDDA.n250 0.0682083
R5547 VDDA.n302 VDDA.n301 0.0682083
R5548 VDDA.n310 VDDA.n309 0.0682083
R5549 VDDA.n316 VDDA.n242 0.0682083
R5550 VDDA.n324 VDDA.n238 0.0682083
R5551 VDDA.n326 VDDA.n325 0.0682083
R5552 VDDA.n334 VDDA.n333 0.0682083
R5553 VDDA.n340 VDDA.n230 0.0682083
R5554 VDDA.n348 VDDA.n226 0.0682083
R5555 VDDA.n350 VDDA.n349 0.0682083
R5556 VDDA.n2595 VDDA.n357 0.0682083
R5557 VDDA.n2477 VDDA.n2476 0.0682083
R5558 VDDA.n2485 VDDA.n2460 0.0682083
R5559 VDDA.n2495 VDDA.n2456 0.0682083
R5560 VDDA.n2497 VDDA.n2496 0.0682083
R5561 VDDA.n2507 VDDA.n2506 0.0682083
R5562 VDDA.n2515 VDDA.n2448 0.0682083
R5563 VDDA.n2525 VDDA.n2444 0.0682083
R5564 VDDA.n2527 VDDA.n2526 0.0682083
R5565 VDDA.n2537 VDDA.n2536 0.0682083
R5566 VDDA.n2545 VDDA.n2436 0.0682083
R5567 VDDA.n2555 VDDA.n2432 0.0682083
R5568 VDDA.n2557 VDDA.n2556 0.0682083
R5569 VDDA.n2567 VDDA.n2566 0.0682083
R5570 VDDA.n2575 VDDA.n2424 0.0682083
R5571 VDDA.n2584 VDDA.n2420 0.0682083
R5572 VDDA.n1234 VDDA.n1233 0.0682083
R5573 VDDA.n1240 VDDA.n1220 0.0682083
R5574 VDDA.n1248 VDDA.n1216 0.0682083
R5575 VDDA.n1250 VDDA.n1249 0.0682083
R5576 VDDA.n1258 VDDA.n1257 0.0682083
R5577 VDDA.n1264 VDDA.n1208 0.0682083
R5578 VDDA.n1272 VDDA.n1204 0.0682083
R5579 VDDA.n1274 VDDA.n1273 0.0682083
R5580 VDDA.n1282 VDDA.n1281 0.0682083
R5581 VDDA.n1288 VDDA.n1196 0.0682083
R5582 VDDA.n1296 VDDA.n1192 0.0682083
R5583 VDDA.n1298 VDDA.n1297 0.0682083
R5584 VDDA.n1306 VDDA.n1305 0.0682083
R5585 VDDA.n1312 VDDA.n1184 0.0682083
R5586 VDDA.n2257 VDDA.n458 0.0682083
R5587 VDDA.n542 VDDA.n528 0.0682083
R5588 VDDA.n544 VDDA.n543 0.0682083
R5589 VDDA.n552 VDDA.n551 0.0682083
R5590 VDDA.n558 VDDA.n520 0.0682083
R5591 VDDA.n566 VDDA.n516 0.0682083
R5592 VDDA.n568 VDDA.n567 0.0682083
R5593 VDDA.n576 VDDA.n575 0.0682083
R5594 VDDA.n582 VDDA.n508 0.0682083
R5595 VDDA.n590 VDDA.n504 0.0682083
R5596 VDDA.n592 VDDA.n591 0.0682083
R5597 VDDA.n600 VDDA.n599 0.0682083
R5598 VDDA.n606 VDDA.n496 0.0682083
R5599 VDDA.n614 VDDA.n492 0.0682083
R5600 VDDA.n616 VDDA.n615 0.0682083
R5601 VDDA.n1155 VDDA.n623 0.0682083
R5602 VDDA.n1037 VDDA.n1036 0.0682083
R5603 VDDA.n1045 VDDA.n1020 0.0682083
R5604 VDDA.n1055 VDDA.n1016 0.0682083
R5605 VDDA.n1057 VDDA.n1056 0.0682083
R5606 VDDA.n1067 VDDA.n1066 0.0682083
R5607 VDDA.n1075 VDDA.n1008 0.0682083
R5608 VDDA.n1085 VDDA.n1004 0.0682083
R5609 VDDA.n1087 VDDA.n1086 0.0682083
R5610 VDDA.n1097 VDDA.n1096 0.0682083
R5611 VDDA.n1105 VDDA.n996 0.0682083
R5612 VDDA.n1115 VDDA.n992 0.0682083
R5613 VDDA.n1117 VDDA.n1116 0.0682083
R5614 VDDA.n1127 VDDA.n1126 0.0682083
R5615 VDDA.n1135 VDDA.n984 0.0682083
R5616 VDDA.n1144 VDDA.n980 0.0682083
R5617 VDDA.n886 VDDA.n885 0.0682083
R5618 VDDA.n892 VDDA.n872 0.0682083
R5619 VDDA.n900 VDDA.n868 0.0682083
R5620 VDDA.n902 VDDA.n901 0.0682083
R5621 VDDA.n910 VDDA.n909 0.0682083
R5622 VDDA.n916 VDDA.n860 0.0682083
R5623 VDDA.n924 VDDA.n856 0.0682083
R5624 VDDA.n926 VDDA.n925 0.0682083
R5625 VDDA.n934 VDDA.n933 0.0682083
R5626 VDDA.n940 VDDA.n848 0.0682083
R5627 VDDA.n948 VDDA.n844 0.0682083
R5628 VDDA.n950 VDDA.n949 0.0682083
R5629 VDDA.n958 VDDA.n957 0.0682083
R5630 VDDA.n964 VDDA.n836 0.0682083
R5631 VDDA.n973 VDDA.n635 0.0682083
R5632 VDDA.n698 VDDA.n684 0.0682083
R5633 VDDA.n700 VDDA.n699 0.0682083
R5634 VDDA.n710 VDDA.n709 0.0682083
R5635 VDDA.n718 VDDA.n680 0.0682083
R5636 VDDA.n728 VDDA.n678 0.0682083
R5637 VDDA.n730 VDDA.n729 0.0682083
R5638 VDDA.n740 VDDA.n739 0.0682083
R5639 VDDA.n748 VDDA.n674 0.0682083
R5640 VDDA.n758 VDDA.n672 0.0682083
R5641 VDDA.n760 VDDA.n759 0.0682083
R5642 VDDA.n770 VDDA.n769 0.0682083
R5643 VDDA.n778 VDDA.n668 0.0682083
R5644 VDDA.n788 VDDA.n666 0.0682083
R5645 VDDA.n790 VDDA.n789 0.0682083
R5646 VDDA.n807 VDDA.n799 0.0682083
R5647 VDDA.n90 VDDA.n89 0.0672139
R5648 VDDA.n2816 VDDA.n2815 0.0672139
R5649 VDDA.n2667 VDDA.n2665 0.0672139
R5650 VDDA.n268 VDDA.n267 0.0672139
R5651 VDDA.n2468 VDDA.n2467 0.0672139
R5652 VDDA.n1227 VDDA.n1225 0.0672139
R5653 VDDA.n534 VDDA.n533 0.0672139
R5654 VDDA.n1028 VDDA.n1027 0.0672139
R5655 VDDA.n879 VDDA.n877 0.0672139
R5656 VDDA.n1576 VDDA.n1433 0.0672139
R5657 VDDA.n2251 VDDA.n1908 0.0672139
R5658 VDDA.n688 VDDA.n687 0.0672139
R5659 VDDA.n1749 VDDA.n1582 0.0657174
R5660 VDDA.n1733 VDDA.n1591 0.0657174
R5661 VDDA.n1719 VDDA.n1601 0.0657174
R5662 VDDA.n1703 VDDA.n1609 0.0657174
R5663 VDDA.n1689 VDDA.n1619 0.0657174
R5664 VDDA.n1673 VDDA.n1627 0.0657174
R5665 VDDA.n1659 VDDA.n1637 0.0657174
R5666 VDDA.n1751 VDDA.n1750 0.0657174
R5667 VDDA.n1732 VDDA.n1590 0.0657174
R5668 VDDA.n1721 VDDA.n1720 0.0657174
R5669 VDDA.n1702 VDDA.n1608 0.0657174
R5670 VDDA.n1691 VDDA.n1690 0.0657174
R5671 VDDA.n1672 VDDA.n1626 0.0657174
R5672 VDDA.n1661 VDDA.n1660 0.0657174
R5673 VDDA.n1476 VDDA.n1475 0.063
R5674 VDDA.n1487 VDDA.n1450 0.063
R5675 VDDA.n1506 VDDA.n1505 0.063
R5676 VDDA.n1517 VDDA.n1444 0.063
R5677 VDDA.n1536 VDDA.n1535 0.063
R5678 VDDA.n1547 VDDA.n1438 0.063
R5679 VDDA.n1566 VDDA.n1565 0.063
R5680 VDDA.n2151 VDDA.n2150 0.063
R5681 VDDA.n2162 VDDA.n1925 0.063
R5682 VDDA.n2181 VDDA.n2180 0.063
R5683 VDDA.n2192 VDDA.n1919 0.063
R5684 VDDA.n2211 VDDA.n2210 0.063
R5685 VDDA.n2222 VDDA.n1913 0.063
R5686 VDDA.n2241 VDDA.n2240 0.063
R5687 VDDA.n99 VDDA.n98 0.063
R5688 VDDA.n108 VDDA.n76 0.063
R5689 VDDA.n123 VDDA.n122 0.063
R5690 VDDA.n132 VDDA.n64 0.063
R5691 VDDA.n147 VDDA.n146 0.063
R5692 VDDA.n156 VDDA.n52 0.063
R5693 VDDA.n171 VDDA.n170 0.063
R5694 VDDA.n2825 VDDA.n2808 0.063
R5695 VDDA.n2844 VDDA.n2843 0.063
R5696 VDDA.n2855 VDDA.n2796 0.063
R5697 VDDA.n2874 VDDA.n2873 0.063
R5698 VDDA.n2885 VDDA.n2784 0.063
R5699 VDDA.n2904 VDDA.n2903 0.063
R5700 VDDA.n2915 VDDA.n2772 0.063
R5701 VDDA.n2674 VDDA.n2660 0.063
R5702 VDDA.n2689 VDDA.n2688 0.063
R5703 VDDA.n2698 VDDA.n2648 0.063
R5704 VDDA.n2713 VDDA.n2712 0.063
R5705 VDDA.n2722 VDDA.n2636 0.063
R5706 VDDA.n2737 VDDA.n2736 0.063
R5707 VDDA.n2746 VDDA.n2624 0.063
R5708 VDDA.n277 VDDA.n276 0.063
R5709 VDDA.n286 VDDA.n254 0.063
R5710 VDDA.n301 VDDA.n300 0.063
R5711 VDDA.n310 VDDA.n242 0.063
R5712 VDDA.n325 VDDA.n324 0.063
R5713 VDDA.n334 VDDA.n230 0.063
R5714 VDDA.n349 VDDA.n348 0.063
R5715 VDDA.n2477 VDDA.n2460 0.063
R5716 VDDA.n2496 VDDA.n2495 0.063
R5717 VDDA.n2507 VDDA.n2448 0.063
R5718 VDDA.n2526 VDDA.n2525 0.063
R5719 VDDA.n2537 VDDA.n2436 0.063
R5720 VDDA.n2556 VDDA.n2555 0.063
R5721 VDDA.n2567 VDDA.n2424 0.063
R5722 VDDA.n1234 VDDA.n1220 0.063
R5723 VDDA.n1249 VDDA.n1248 0.063
R5724 VDDA.n1258 VDDA.n1208 0.063
R5725 VDDA.n1273 VDDA.n1272 0.063
R5726 VDDA.n1282 VDDA.n1196 0.063
R5727 VDDA.n1297 VDDA.n1296 0.063
R5728 VDDA.n1306 VDDA.n1184 0.063
R5729 VDDA.n543 VDDA.n542 0.063
R5730 VDDA.n552 VDDA.n520 0.063
R5731 VDDA.n567 VDDA.n566 0.063
R5732 VDDA.n576 VDDA.n508 0.063
R5733 VDDA.n591 VDDA.n590 0.063
R5734 VDDA.n600 VDDA.n496 0.063
R5735 VDDA.n615 VDDA.n614 0.063
R5736 VDDA.n1037 VDDA.n1020 0.063
R5737 VDDA.n1056 VDDA.n1055 0.063
R5738 VDDA.n1067 VDDA.n1008 0.063
R5739 VDDA.n1086 VDDA.n1085 0.063
R5740 VDDA.n1097 VDDA.n996 0.063
R5741 VDDA.n1116 VDDA.n1115 0.063
R5742 VDDA.n1127 VDDA.n984 0.063
R5743 VDDA.n886 VDDA.n872 0.063
R5744 VDDA.n901 VDDA.n900 0.063
R5745 VDDA.n910 VDDA.n860 0.063
R5746 VDDA.n925 VDDA.n924 0.063
R5747 VDDA.n934 VDDA.n848 0.063
R5748 VDDA.n949 VDDA.n948 0.063
R5749 VDDA.n958 VDDA.n836 0.063
R5750 VDDA.n699 VDDA.n698 0.063
R5751 VDDA.n710 VDDA.n680 0.063
R5752 VDDA.n729 VDDA.n728 0.063
R5753 VDDA.n740 VDDA.n674 0.063
R5754 VDDA.n759 VDDA.n758 0.063
R5755 VDDA.n770 VDDA.n668 0.063
R5756 VDDA.n789 VDDA.n788 0.063
R5757 VDDA.n1797 VDDA.n1796 0.0603182
R5758 VDDA.n1811 VDDA.n1810 0.0603182
R5759 VDDA.n1827 VDDA.n1826 0.0603182
R5760 VDDA.n1841 VDDA.n1840 0.0603182
R5761 VDDA.n1857 VDDA.n1856 0.0603182
R5762 VDDA.n1871 VDDA.n1870 0.0603182
R5763 VDDA.n1887 VDDA.n1886 0.0603182
R5764 VDDA.n1901 VDDA.n1900 0.0603182
R5765 VDDA.n1905 VDDA.n1367 0.0581818
R5766 VDDA.n1791 VDDA.n1342 0.0560455
R5767 VDDA.n1801 VDDA.n1800 0.0560455
R5768 VDDA.n1807 VDDA.n1806 0.0560455
R5769 VDDA.n1817 VDDA.n1816 0.0560455
R5770 VDDA.n1821 VDDA.n1820 0.0560455
R5771 VDDA.n1831 VDDA.n1830 0.0560455
R5772 VDDA.n1837 VDDA.n1836 0.0560455
R5773 VDDA.n1847 VDDA.n1846 0.0560455
R5774 VDDA.n1851 VDDA.n1850 0.0560455
R5775 VDDA.n1861 VDDA.n1860 0.0560455
R5776 VDDA.n1867 VDDA.n1866 0.0560455
R5777 VDDA.n1877 VDDA.n1876 0.0560455
R5778 VDDA.n1881 VDDA.n1880 0.0560455
R5779 VDDA.n1891 VDDA.n1890 0.0560455
R5780 VDDA.n1897 VDDA.n1896 0.0560455
R5781 VDDA.n1469 VDDA.n1468 0.0553333
R5782 VDDA.n1483 VDDA.n1482 0.0553333
R5783 VDDA.n1499 VDDA.n1498 0.0553333
R5784 VDDA.n1513 VDDA.n1512 0.0553333
R5785 VDDA.n1529 VDDA.n1528 0.0553333
R5786 VDDA.n1543 VDDA.n1542 0.0553333
R5787 VDDA.n1559 VDDA.n1558 0.0553333
R5788 VDDA.n1573 VDDA.n1572 0.0553333
R5789 VDDA.n2144 VDDA.n2143 0.0553333
R5790 VDDA.n2158 VDDA.n2157 0.0553333
R5791 VDDA.n2174 VDDA.n2173 0.0553333
R5792 VDDA.n2188 VDDA.n2187 0.0553333
R5793 VDDA.n2204 VDDA.n2203 0.0553333
R5794 VDDA.n2218 VDDA.n2217 0.0553333
R5795 VDDA.n2234 VDDA.n2233 0.0553333
R5796 VDDA.n2248 VDDA.n2247 0.0553333
R5797 VDDA.n87 VDDA.n86 0.0553333
R5798 VDDA.n104 VDDA.n103 0.0553333
R5799 VDDA.n75 VDDA.n74 0.0553333
R5800 VDDA.n128 VDDA.n127 0.0553333
R5801 VDDA.n63 VDDA.n62 0.0553333
R5802 VDDA.n152 VDDA.n151 0.0553333
R5803 VDDA.n51 VDDA.n50 0.0553333
R5804 VDDA.n176 VDDA.n175 0.0553333
R5805 VDDA.n2821 VDDA.n2819 0.0553333
R5806 VDDA.n2837 VDDA.n2806 0.0553333
R5807 VDDA.n2851 VDDA.n2849 0.0553333
R5808 VDDA.n2867 VDDA.n2794 0.0553333
R5809 VDDA.n2881 VDDA.n2879 0.0553333
R5810 VDDA.n2897 VDDA.n2782 0.0553333
R5811 VDDA.n2911 VDDA.n2909 0.0553333
R5812 VDDA.n2927 VDDA.n2770 0.0553333
R5813 VDDA.n2670 VDDA.n2669 0.0553333
R5814 VDDA.n2659 VDDA.n2658 0.0553333
R5815 VDDA.n2694 VDDA.n2693 0.0553333
R5816 VDDA.n2647 VDDA.n2646 0.0553333
R5817 VDDA.n2718 VDDA.n2717 0.0553333
R5818 VDDA.n2635 VDDA.n2634 0.0553333
R5819 VDDA.n2742 VDDA.n2741 0.0553333
R5820 VDDA.n2756 VDDA.n2622 0.0553333
R5821 VDDA.n265 VDDA.n264 0.0553333
R5822 VDDA.n282 VDDA.n281 0.0553333
R5823 VDDA.n253 VDDA.n252 0.0553333
R5824 VDDA.n306 VDDA.n305 0.0553333
R5825 VDDA.n241 VDDA.n240 0.0553333
R5826 VDDA.n330 VDDA.n329 0.0553333
R5827 VDDA.n229 VDDA.n228 0.0553333
R5828 VDDA.n354 VDDA.n353 0.0553333
R5829 VDDA.n2473 VDDA.n2471 0.0553333
R5830 VDDA.n2489 VDDA.n2458 0.0553333
R5831 VDDA.n2503 VDDA.n2501 0.0553333
R5832 VDDA.n2519 VDDA.n2446 0.0553333
R5833 VDDA.n2533 VDDA.n2531 0.0553333
R5834 VDDA.n2549 VDDA.n2434 0.0553333
R5835 VDDA.n2563 VDDA.n2561 0.0553333
R5836 VDDA.n2579 VDDA.n2422 0.0553333
R5837 VDDA.n1230 VDDA.n1229 0.0553333
R5838 VDDA.n1219 VDDA.n1218 0.0553333
R5839 VDDA.n1254 VDDA.n1253 0.0553333
R5840 VDDA.n1207 VDDA.n1206 0.0553333
R5841 VDDA.n1278 VDDA.n1277 0.0553333
R5842 VDDA.n1195 VDDA.n1194 0.0553333
R5843 VDDA.n1302 VDDA.n1301 0.0553333
R5844 VDDA.n1316 VDDA.n1182 0.0553333
R5845 VDDA.n531 VDDA.n530 0.0553333
R5846 VDDA.n548 VDDA.n547 0.0553333
R5847 VDDA.n519 VDDA.n518 0.0553333
R5848 VDDA.n572 VDDA.n571 0.0553333
R5849 VDDA.n507 VDDA.n506 0.0553333
R5850 VDDA.n596 VDDA.n595 0.0553333
R5851 VDDA.n495 VDDA.n494 0.0553333
R5852 VDDA.n620 VDDA.n619 0.0553333
R5853 VDDA.n1033 VDDA.n1031 0.0553333
R5854 VDDA.n1049 VDDA.n1018 0.0553333
R5855 VDDA.n1063 VDDA.n1061 0.0553333
R5856 VDDA.n1079 VDDA.n1006 0.0553333
R5857 VDDA.n1093 VDDA.n1091 0.0553333
R5858 VDDA.n1109 VDDA.n994 0.0553333
R5859 VDDA.n1123 VDDA.n1121 0.0553333
R5860 VDDA.n1139 VDDA.n982 0.0553333
R5861 VDDA.n882 VDDA.n881 0.0553333
R5862 VDDA.n871 VDDA.n870 0.0553333
R5863 VDDA.n906 VDDA.n905 0.0553333
R5864 VDDA.n859 VDDA.n858 0.0553333
R5865 VDDA.n930 VDDA.n929 0.0553333
R5866 VDDA.n847 VDDA.n846 0.0553333
R5867 VDDA.n954 VDDA.n953 0.0553333
R5868 VDDA.n968 VDDA.n834 0.0553333
R5869 VDDA.n692 VDDA.n691 0.0553333
R5870 VDDA.n706 VDDA.n705 0.0553333
R5871 VDDA.n722 VDDA.n721 0.0553333
R5872 VDDA.n736 VDDA.n735 0.0553333
R5873 VDDA.n752 VDDA.n751 0.0553333
R5874 VDDA.n766 VDDA.n765 0.0553333
R5875 VDDA.n782 VDDA.n781 0.0553333
R5876 VDDA.n796 VDDA.n795 0.0553333
R5877 VDDA.n1463 VDDA.n1408 0.0514167
R5878 VDDA.n1473 VDDA.n1472 0.0514167
R5879 VDDA.n1479 VDDA.n1478 0.0514167
R5880 VDDA.n1489 VDDA.n1488 0.0514167
R5881 VDDA.n1493 VDDA.n1492 0.0514167
R5882 VDDA.n1503 VDDA.n1502 0.0514167
R5883 VDDA.n1509 VDDA.n1508 0.0514167
R5884 VDDA.n1519 VDDA.n1518 0.0514167
R5885 VDDA.n1523 VDDA.n1522 0.0514167
R5886 VDDA.n1533 VDDA.n1532 0.0514167
R5887 VDDA.n1539 VDDA.n1538 0.0514167
R5888 VDDA.n1549 VDDA.n1548 0.0514167
R5889 VDDA.n1553 VDDA.n1552 0.0514167
R5890 VDDA.n1563 VDDA.n1562 0.0514167
R5891 VDDA.n1569 VDDA.n1568 0.0514167
R5892 VDDA.n1577 VDDA.n1432 0.0514167
R5893 VDDA.n2138 VDDA.n1318 0.0514167
R5894 VDDA.n2148 VDDA.n2147 0.0514167
R5895 VDDA.n2154 VDDA.n2153 0.0514167
R5896 VDDA.n2164 VDDA.n2163 0.0514167
R5897 VDDA.n2168 VDDA.n2167 0.0514167
R5898 VDDA.n2178 VDDA.n2177 0.0514167
R5899 VDDA.n2184 VDDA.n2183 0.0514167
R5900 VDDA.n2194 VDDA.n2193 0.0514167
R5901 VDDA.n2198 VDDA.n2197 0.0514167
R5902 VDDA.n2208 VDDA.n2207 0.0514167
R5903 VDDA.n2214 VDDA.n2213 0.0514167
R5904 VDDA.n2224 VDDA.n2223 0.0514167
R5905 VDDA.n2228 VDDA.n2227 0.0514167
R5906 VDDA.n2238 VDDA.n2237 0.0514167
R5907 VDDA.n2244 VDDA.n2243 0.0514167
R5908 VDDA.n2252 VDDA.n1907 0.0514167
R5909 VDDA.n88 VDDA.n18 0.0514167
R5910 VDDA.n96 VDDA.n95 0.0514167
R5911 VDDA.n83 VDDA.n82 0.0514167
R5912 VDDA.n79 VDDA.n78 0.0514167
R5913 VDDA.n112 VDDA.n111 0.0514167
R5914 VDDA.n120 VDDA.n119 0.0514167
R5915 VDDA.n71 VDDA.n70 0.0514167
R5916 VDDA.n67 VDDA.n66 0.0514167
R5917 VDDA.n136 VDDA.n135 0.0514167
R5918 VDDA.n144 VDDA.n143 0.0514167
R5919 VDDA.n59 VDDA.n58 0.0514167
R5920 VDDA.n55 VDDA.n54 0.0514167
R5921 VDDA.n160 VDDA.n159 0.0514167
R5922 VDDA.n168 VDDA.n167 0.0514167
R5923 VDDA.n47 VDDA.n46 0.0514167
R5924 VDDA.n2945 VDDA.n42 0.0514167
R5925 VDDA.n2817 VDDA.n2814 0.0514167
R5926 VDDA.n2827 VDDA.n2810 0.0514167
R5927 VDDA.n2831 VDDA.n2829 0.0514167
R5928 VDDA.n2841 VDDA.n2839 0.0514167
R5929 VDDA.n2847 VDDA.n2802 0.0514167
R5930 VDDA.n2857 VDDA.n2798 0.0514167
R5931 VDDA.n2861 VDDA.n2859 0.0514167
R5932 VDDA.n2871 VDDA.n2869 0.0514167
R5933 VDDA.n2877 VDDA.n2790 0.0514167
R5934 VDDA.n2887 VDDA.n2786 0.0514167
R5935 VDDA.n2891 VDDA.n2889 0.0514167
R5936 VDDA.n2901 VDDA.n2899 0.0514167
R5937 VDDA.n2907 VDDA.n2778 0.0514167
R5938 VDDA.n2917 VDDA.n2774 0.0514167
R5939 VDDA.n2921 VDDA.n2919 0.0514167
R5940 VDDA.n2930 VDDA.n2929 0.0514167
R5941 VDDA.n2666 VDDA.n2599 0.0514167
R5942 VDDA.n2663 VDDA.n2662 0.0514167
R5943 VDDA.n2678 VDDA.n2677 0.0514167
R5944 VDDA.n2686 VDDA.n2685 0.0514167
R5945 VDDA.n2655 VDDA.n2654 0.0514167
R5946 VDDA.n2651 VDDA.n2650 0.0514167
R5947 VDDA.n2702 VDDA.n2701 0.0514167
R5948 VDDA.n2710 VDDA.n2709 0.0514167
R5949 VDDA.n2643 VDDA.n2642 0.0514167
R5950 VDDA.n2639 VDDA.n2638 0.0514167
R5951 VDDA.n2726 VDDA.n2725 0.0514167
R5952 VDDA.n2734 VDDA.n2733 0.0514167
R5953 VDDA.n2631 VDDA.n2630 0.0514167
R5954 VDDA.n2627 VDDA.n2626 0.0514167
R5955 VDDA.n2750 VDDA.n2749 0.0514167
R5956 VDDA.n2759 VDDA.n194 0.0514167
R5957 VDDA.n266 VDDA.n196 0.0514167
R5958 VDDA.n274 VDDA.n273 0.0514167
R5959 VDDA.n261 VDDA.n260 0.0514167
R5960 VDDA.n257 VDDA.n256 0.0514167
R5961 VDDA.n290 VDDA.n289 0.0514167
R5962 VDDA.n298 VDDA.n297 0.0514167
R5963 VDDA.n249 VDDA.n248 0.0514167
R5964 VDDA.n245 VDDA.n244 0.0514167
R5965 VDDA.n314 VDDA.n313 0.0514167
R5966 VDDA.n322 VDDA.n321 0.0514167
R5967 VDDA.n237 VDDA.n236 0.0514167
R5968 VDDA.n233 VDDA.n232 0.0514167
R5969 VDDA.n338 VDDA.n337 0.0514167
R5970 VDDA.n346 VDDA.n345 0.0514167
R5971 VDDA.n225 VDDA.n224 0.0514167
R5972 VDDA.n2597 VDDA.n220 0.0514167
R5973 VDDA.n2469 VDDA.n2466 0.0514167
R5974 VDDA.n2479 VDDA.n2462 0.0514167
R5975 VDDA.n2483 VDDA.n2481 0.0514167
R5976 VDDA.n2493 VDDA.n2491 0.0514167
R5977 VDDA.n2499 VDDA.n2454 0.0514167
R5978 VDDA.n2509 VDDA.n2450 0.0514167
R5979 VDDA.n2513 VDDA.n2511 0.0514167
R5980 VDDA.n2523 VDDA.n2521 0.0514167
R5981 VDDA.n2529 VDDA.n2442 0.0514167
R5982 VDDA.n2539 VDDA.n2438 0.0514167
R5983 VDDA.n2543 VDDA.n2541 0.0514167
R5984 VDDA.n2553 VDDA.n2551 0.0514167
R5985 VDDA.n2559 VDDA.n2430 0.0514167
R5986 VDDA.n2569 VDDA.n2426 0.0514167
R5987 VDDA.n2573 VDDA.n2571 0.0514167
R5988 VDDA.n2582 VDDA.n2581 0.0514167
R5989 VDDA.n1226 VDDA.n1159 0.0514167
R5990 VDDA.n1223 VDDA.n1222 0.0514167
R5991 VDDA.n1238 VDDA.n1237 0.0514167
R5992 VDDA.n1246 VDDA.n1245 0.0514167
R5993 VDDA.n1215 VDDA.n1214 0.0514167
R5994 VDDA.n1211 VDDA.n1210 0.0514167
R5995 VDDA.n1262 VDDA.n1261 0.0514167
R5996 VDDA.n1270 VDDA.n1269 0.0514167
R5997 VDDA.n1203 VDDA.n1202 0.0514167
R5998 VDDA.n1199 VDDA.n1198 0.0514167
R5999 VDDA.n1286 VDDA.n1285 0.0514167
R6000 VDDA.n1294 VDDA.n1293 0.0514167
R6001 VDDA.n1191 VDDA.n1190 0.0514167
R6002 VDDA.n1187 VDDA.n1186 0.0514167
R6003 VDDA.n1310 VDDA.n1309 0.0514167
R6004 VDDA.n2255 VDDA.n460 0.0514167
R6005 VDDA.n532 VDDA.n462 0.0514167
R6006 VDDA.n540 VDDA.n539 0.0514167
R6007 VDDA.n527 VDDA.n526 0.0514167
R6008 VDDA.n523 VDDA.n522 0.0514167
R6009 VDDA.n556 VDDA.n555 0.0514167
R6010 VDDA.n564 VDDA.n563 0.0514167
R6011 VDDA.n515 VDDA.n514 0.0514167
R6012 VDDA.n511 VDDA.n510 0.0514167
R6013 VDDA.n580 VDDA.n579 0.0514167
R6014 VDDA.n588 VDDA.n587 0.0514167
R6015 VDDA.n503 VDDA.n502 0.0514167
R6016 VDDA.n499 VDDA.n498 0.0514167
R6017 VDDA.n604 VDDA.n603 0.0514167
R6018 VDDA.n612 VDDA.n611 0.0514167
R6019 VDDA.n491 VDDA.n490 0.0514167
R6020 VDDA.n1157 VDDA.n486 0.0514167
R6021 VDDA.n1029 VDDA.n1026 0.0514167
R6022 VDDA.n1039 VDDA.n1022 0.0514167
R6023 VDDA.n1043 VDDA.n1041 0.0514167
R6024 VDDA.n1053 VDDA.n1051 0.0514167
R6025 VDDA.n1059 VDDA.n1014 0.0514167
R6026 VDDA.n1069 VDDA.n1010 0.0514167
R6027 VDDA.n1073 VDDA.n1071 0.0514167
R6028 VDDA.n1083 VDDA.n1081 0.0514167
R6029 VDDA.n1089 VDDA.n1002 0.0514167
R6030 VDDA.n1099 VDDA.n998 0.0514167
R6031 VDDA.n1103 VDDA.n1101 0.0514167
R6032 VDDA.n1113 VDDA.n1111 0.0514167
R6033 VDDA.n1119 VDDA.n990 0.0514167
R6034 VDDA.n1129 VDDA.n986 0.0514167
R6035 VDDA.n1133 VDDA.n1131 0.0514167
R6036 VDDA.n1142 VDDA.n1141 0.0514167
R6037 VDDA.n878 VDDA.n811 0.0514167
R6038 VDDA.n875 VDDA.n874 0.0514167
R6039 VDDA.n890 VDDA.n889 0.0514167
R6040 VDDA.n898 VDDA.n897 0.0514167
R6041 VDDA.n867 VDDA.n866 0.0514167
R6042 VDDA.n863 VDDA.n862 0.0514167
R6043 VDDA.n914 VDDA.n913 0.0514167
R6044 VDDA.n922 VDDA.n921 0.0514167
R6045 VDDA.n855 VDDA.n854 0.0514167
R6046 VDDA.n851 VDDA.n850 0.0514167
R6047 VDDA.n938 VDDA.n937 0.0514167
R6048 VDDA.n946 VDDA.n945 0.0514167
R6049 VDDA.n843 VDDA.n842 0.0514167
R6050 VDDA.n839 VDDA.n838 0.0514167
R6051 VDDA.n962 VDDA.n961 0.0514167
R6052 VDDA.n971 VDDA.n637 0.0514167
R6053 VDDA.n686 VDDA.n638 0.0514167
R6054 VDDA.n696 VDDA.n695 0.0514167
R6055 VDDA.n702 VDDA.n701 0.0514167
R6056 VDDA.n712 VDDA.n711 0.0514167
R6057 VDDA.n716 VDDA.n715 0.0514167
R6058 VDDA.n726 VDDA.n725 0.0514167
R6059 VDDA.n732 VDDA.n731 0.0514167
R6060 VDDA.n742 VDDA.n741 0.0514167
R6061 VDDA.n746 VDDA.n745 0.0514167
R6062 VDDA.n756 VDDA.n755 0.0514167
R6063 VDDA.n762 VDDA.n761 0.0514167
R6064 VDDA.n772 VDDA.n771 0.0514167
R6065 VDDA.n776 VDDA.n775 0.0514167
R6066 VDDA.n786 VDDA.n785 0.0514167
R6067 VDDA.n792 VDDA.n791 0.0514167
R6068 VDDA.n809 VDDA.n662 0.0514167
R6069 VDDA.n2253 VDDA.n1906 0.0487484
R6070 VDDA.n2393 VDDA.n388 0.0421667
R6071 VDDA.n978 VDDA.n630 0.0421667
R6072 VDDA.n1149 VDDA.n627 0.0421667
R6073 VDDA.n625 VDDA.n456 0.0421667
R6074 VDDA.n2262 VDDA.n453 0.0421667
R6075 VDDA.n2282 VDDA.n450 0.0421667
R6076 VDDA.n2400 VDDA.n366 0.0421667
R6077 VDDA.n2589 VDDA.n361 0.0421667
R6078 VDDA.n359 VDDA.n190 0.0421667
R6079 VDDA.n2766 VDDA.n187 0.0421667
R6080 VDDA.n2937 VDDA.n184 0.0421667
R6081 VDDA.n2940 VDDA.n182 0.0421667
R6082 VDDA.n1650 VDDA.n1649 0.0352506
R6083 VDDA.n1764 VDDA.n1763 0.0331087
R6084 VDDA.n1796 VDDA.n1343 0.030649
R6085 VDDA.n1800 VDDA.n1344 0.030649
R6086 VDDA.n1810 VDDA.n1346 0.030649
R6087 VDDA.n1816 VDDA.n1347 0.030649
R6088 VDDA.n1826 VDDA.n1349 0.030649
R6089 VDDA.n1830 VDDA.n1350 0.030649
R6090 VDDA.n1840 VDDA.n1352 0.030649
R6091 VDDA.n1846 VDDA.n1353 0.030649
R6092 VDDA.n1856 VDDA.n1355 0.030649
R6093 VDDA.n1860 VDDA.n1356 0.030649
R6094 VDDA.n1870 VDDA.n1358 0.030649
R6095 VDDA.n1876 VDDA.n1359 0.030649
R6096 VDDA.n1886 VDDA.n1361 0.030649
R6097 VDDA.n1890 VDDA.n1362 0.030649
R6098 VDDA.n1900 VDDA.n1364 0.030649
R6099 VDDA.n1367 VDDA.n1365 0.030649
R6100 VDDA.n1901 VDDA.n1365 0.030649
R6101 VDDA.n1897 VDDA.n1364 0.030649
R6102 VDDA.n1887 VDDA.n1362 0.030649
R6103 VDDA.n1881 VDDA.n1361 0.030649
R6104 VDDA.n1871 VDDA.n1359 0.030649
R6105 VDDA.n1867 VDDA.n1358 0.030649
R6106 VDDA.n1857 VDDA.n1356 0.030649
R6107 VDDA.n1851 VDDA.n1355 0.030649
R6108 VDDA.n1841 VDDA.n1353 0.030649
R6109 VDDA.n1837 VDDA.n1352 0.030649
R6110 VDDA.n1827 VDDA.n1350 0.030649
R6111 VDDA.n1821 VDDA.n1349 0.030649
R6112 VDDA.n1811 VDDA.n1347 0.030649
R6113 VDDA.n1807 VDDA.n1346 0.030649
R6114 VDDA.n1797 VDDA.n1344 0.030649
R6115 VDDA.n1791 VDDA.n1343 0.030649
R6116 VDDA.n1468 VDDA.n1409 0.028198
R6117 VDDA.n1472 VDDA.n1410 0.028198
R6118 VDDA.n1482 VDDA.n1412 0.028198
R6119 VDDA.n1488 VDDA.n1413 0.028198
R6120 VDDA.n1498 VDDA.n1415 0.028198
R6121 VDDA.n1502 VDDA.n1416 0.028198
R6122 VDDA.n1512 VDDA.n1418 0.028198
R6123 VDDA.n1518 VDDA.n1419 0.028198
R6124 VDDA.n1528 VDDA.n1421 0.028198
R6125 VDDA.n1532 VDDA.n1422 0.028198
R6126 VDDA.n1542 VDDA.n1424 0.028198
R6127 VDDA.n1548 VDDA.n1425 0.028198
R6128 VDDA.n1558 VDDA.n1427 0.028198
R6129 VDDA.n1562 VDDA.n1428 0.028198
R6130 VDDA.n1572 VDDA.n1430 0.028198
R6131 VDDA.n1432 VDDA.n1431 0.028198
R6132 VDDA.n2143 VDDA.n1319 0.028198
R6133 VDDA.n2147 VDDA.n1320 0.028198
R6134 VDDA.n2157 VDDA.n1322 0.028198
R6135 VDDA.n2163 VDDA.n1323 0.028198
R6136 VDDA.n2173 VDDA.n1325 0.028198
R6137 VDDA.n2177 VDDA.n1326 0.028198
R6138 VDDA.n2187 VDDA.n1328 0.028198
R6139 VDDA.n2193 VDDA.n1329 0.028198
R6140 VDDA.n2203 VDDA.n1331 0.028198
R6141 VDDA.n2207 VDDA.n1332 0.028198
R6142 VDDA.n2217 VDDA.n1334 0.028198
R6143 VDDA.n2223 VDDA.n1335 0.028198
R6144 VDDA.n2233 VDDA.n1337 0.028198
R6145 VDDA.n2237 VDDA.n1338 0.028198
R6146 VDDA.n2247 VDDA.n1340 0.028198
R6147 VDDA.n1907 VDDA.n1341 0.028198
R6148 VDDA.n86 VDDA.n19 0.028198
R6149 VDDA.n95 VDDA.n20 0.028198
R6150 VDDA.n103 VDDA.n22 0.028198
R6151 VDDA.n78 VDDA.n23 0.028198
R6152 VDDA.n74 VDDA.n25 0.028198
R6153 VDDA.n119 VDDA.n26 0.028198
R6154 VDDA.n127 VDDA.n28 0.028198
R6155 VDDA.n66 VDDA.n29 0.028198
R6156 VDDA.n62 VDDA.n31 0.028198
R6157 VDDA.n143 VDDA.n32 0.028198
R6158 VDDA.n151 VDDA.n34 0.028198
R6159 VDDA.n54 VDDA.n35 0.028198
R6160 VDDA.n50 VDDA.n37 0.028198
R6161 VDDA.n167 VDDA.n38 0.028198
R6162 VDDA.n175 VDDA.n40 0.028198
R6163 VDDA.n42 VDDA.n41 0.028198
R6164 VDDA.n2819 VDDA.n2818 0.028198
R6165 VDDA.n2820 VDDA.n2810 0.028198
R6166 VDDA.n2830 VDDA.n2806 0.028198
R6167 VDDA.n2839 VDDA.n2838 0.028198
R6168 VDDA.n2849 VDDA.n2848 0.028198
R6169 VDDA.n2850 VDDA.n2798 0.028198
R6170 VDDA.n2860 VDDA.n2794 0.028198
R6171 VDDA.n2869 VDDA.n2868 0.028198
R6172 VDDA.n2879 VDDA.n2878 0.028198
R6173 VDDA.n2880 VDDA.n2786 0.028198
R6174 VDDA.n2890 VDDA.n2782 0.028198
R6175 VDDA.n2899 VDDA.n2898 0.028198
R6176 VDDA.n2909 VDDA.n2908 0.028198
R6177 VDDA.n2910 VDDA.n2774 0.028198
R6178 VDDA.n2920 VDDA.n2770 0.028198
R6179 VDDA.n2929 VDDA.n2928 0.028198
R6180 VDDA.n2669 VDDA.n2600 0.028198
R6181 VDDA.n2662 VDDA.n2601 0.028198
R6182 VDDA.n2658 VDDA.n2603 0.028198
R6183 VDDA.n2685 VDDA.n2604 0.028198
R6184 VDDA.n2693 VDDA.n2606 0.028198
R6185 VDDA.n2650 VDDA.n2607 0.028198
R6186 VDDA.n2646 VDDA.n2609 0.028198
R6187 VDDA.n2709 VDDA.n2610 0.028198
R6188 VDDA.n2717 VDDA.n2612 0.028198
R6189 VDDA.n2638 VDDA.n2613 0.028198
R6190 VDDA.n2634 VDDA.n2615 0.028198
R6191 VDDA.n2733 VDDA.n2616 0.028198
R6192 VDDA.n2741 VDDA.n2618 0.028198
R6193 VDDA.n2626 VDDA.n2619 0.028198
R6194 VDDA.n2622 VDDA.n2621 0.028198
R6195 VDDA.n2757 VDDA.n194 0.028198
R6196 VDDA.n264 VDDA.n197 0.028198
R6197 VDDA.n273 VDDA.n198 0.028198
R6198 VDDA.n281 VDDA.n200 0.028198
R6199 VDDA.n256 VDDA.n201 0.028198
R6200 VDDA.n252 VDDA.n203 0.028198
R6201 VDDA.n297 VDDA.n204 0.028198
R6202 VDDA.n305 VDDA.n206 0.028198
R6203 VDDA.n244 VDDA.n207 0.028198
R6204 VDDA.n240 VDDA.n209 0.028198
R6205 VDDA.n321 VDDA.n210 0.028198
R6206 VDDA.n329 VDDA.n212 0.028198
R6207 VDDA.n232 VDDA.n213 0.028198
R6208 VDDA.n228 VDDA.n215 0.028198
R6209 VDDA.n345 VDDA.n216 0.028198
R6210 VDDA.n353 VDDA.n218 0.028198
R6211 VDDA.n220 VDDA.n219 0.028198
R6212 VDDA.n2471 VDDA.n2470 0.028198
R6213 VDDA.n2472 VDDA.n2462 0.028198
R6214 VDDA.n2482 VDDA.n2458 0.028198
R6215 VDDA.n2491 VDDA.n2490 0.028198
R6216 VDDA.n2501 VDDA.n2500 0.028198
R6217 VDDA.n2502 VDDA.n2450 0.028198
R6218 VDDA.n2512 VDDA.n2446 0.028198
R6219 VDDA.n2521 VDDA.n2520 0.028198
R6220 VDDA.n2531 VDDA.n2530 0.028198
R6221 VDDA.n2532 VDDA.n2438 0.028198
R6222 VDDA.n2542 VDDA.n2434 0.028198
R6223 VDDA.n2551 VDDA.n2550 0.028198
R6224 VDDA.n2561 VDDA.n2560 0.028198
R6225 VDDA.n2562 VDDA.n2426 0.028198
R6226 VDDA.n2572 VDDA.n2422 0.028198
R6227 VDDA.n2581 VDDA.n2580 0.028198
R6228 VDDA.n1229 VDDA.n1160 0.028198
R6229 VDDA.n1222 VDDA.n1161 0.028198
R6230 VDDA.n1218 VDDA.n1163 0.028198
R6231 VDDA.n1245 VDDA.n1164 0.028198
R6232 VDDA.n1253 VDDA.n1166 0.028198
R6233 VDDA.n1210 VDDA.n1167 0.028198
R6234 VDDA.n1206 VDDA.n1169 0.028198
R6235 VDDA.n1269 VDDA.n1170 0.028198
R6236 VDDA.n1277 VDDA.n1172 0.028198
R6237 VDDA.n1198 VDDA.n1173 0.028198
R6238 VDDA.n1194 VDDA.n1175 0.028198
R6239 VDDA.n1293 VDDA.n1176 0.028198
R6240 VDDA.n1301 VDDA.n1178 0.028198
R6241 VDDA.n1186 VDDA.n1179 0.028198
R6242 VDDA.n1182 VDDA.n1181 0.028198
R6243 VDDA.n1317 VDDA.n460 0.028198
R6244 VDDA.n530 VDDA.n463 0.028198
R6245 VDDA.n539 VDDA.n464 0.028198
R6246 VDDA.n547 VDDA.n466 0.028198
R6247 VDDA.n522 VDDA.n467 0.028198
R6248 VDDA.n518 VDDA.n469 0.028198
R6249 VDDA.n563 VDDA.n470 0.028198
R6250 VDDA.n571 VDDA.n472 0.028198
R6251 VDDA.n510 VDDA.n473 0.028198
R6252 VDDA.n506 VDDA.n475 0.028198
R6253 VDDA.n587 VDDA.n476 0.028198
R6254 VDDA.n595 VDDA.n478 0.028198
R6255 VDDA.n498 VDDA.n479 0.028198
R6256 VDDA.n494 VDDA.n481 0.028198
R6257 VDDA.n611 VDDA.n482 0.028198
R6258 VDDA.n619 VDDA.n484 0.028198
R6259 VDDA.n486 VDDA.n485 0.028198
R6260 VDDA.n1031 VDDA.n1030 0.028198
R6261 VDDA.n1032 VDDA.n1022 0.028198
R6262 VDDA.n1042 VDDA.n1018 0.028198
R6263 VDDA.n1051 VDDA.n1050 0.028198
R6264 VDDA.n1061 VDDA.n1060 0.028198
R6265 VDDA.n1062 VDDA.n1010 0.028198
R6266 VDDA.n1072 VDDA.n1006 0.028198
R6267 VDDA.n1081 VDDA.n1080 0.028198
R6268 VDDA.n1091 VDDA.n1090 0.028198
R6269 VDDA.n1092 VDDA.n998 0.028198
R6270 VDDA.n1102 VDDA.n994 0.028198
R6271 VDDA.n1111 VDDA.n1110 0.028198
R6272 VDDA.n1121 VDDA.n1120 0.028198
R6273 VDDA.n1122 VDDA.n986 0.028198
R6274 VDDA.n1132 VDDA.n982 0.028198
R6275 VDDA.n1141 VDDA.n1140 0.028198
R6276 VDDA.n881 VDDA.n812 0.028198
R6277 VDDA.n874 VDDA.n813 0.028198
R6278 VDDA.n870 VDDA.n815 0.028198
R6279 VDDA.n897 VDDA.n816 0.028198
R6280 VDDA.n905 VDDA.n818 0.028198
R6281 VDDA.n862 VDDA.n819 0.028198
R6282 VDDA.n858 VDDA.n821 0.028198
R6283 VDDA.n921 VDDA.n822 0.028198
R6284 VDDA.n929 VDDA.n824 0.028198
R6285 VDDA.n850 VDDA.n825 0.028198
R6286 VDDA.n846 VDDA.n827 0.028198
R6287 VDDA.n945 VDDA.n828 0.028198
R6288 VDDA.n953 VDDA.n830 0.028198
R6289 VDDA.n838 VDDA.n831 0.028198
R6290 VDDA.n834 VDDA.n833 0.028198
R6291 VDDA.n969 VDDA.n637 0.028198
R6292 VDDA.n691 VDDA.n639 0.028198
R6293 VDDA.n695 VDDA.n640 0.028198
R6294 VDDA.n705 VDDA.n642 0.028198
R6295 VDDA.n711 VDDA.n643 0.028198
R6296 VDDA.n721 VDDA.n645 0.028198
R6297 VDDA.n725 VDDA.n646 0.028198
R6298 VDDA.n735 VDDA.n648 0.028198
R6299 VDDA.n741 VDDA.n649 0.028198
R6300 VDDA.n751 VDDA.n651 0.028198
R6301 VDDA.n755 VDDA.n652 0.028198
R6302 VDDA.n765 VDDA.n654 0.028198
R6303 VDDA.n771 VDDA.n655 0.028198
R6304 VDDA.n781 VDDA.n657 0.028198
R6305 VDDA.n785 VDDA.n658 0.028198
R6306 VDDA.n795 VDDA.n660 0.028198
R6307 VDDA.n662 VDDA.n661 0.028198
R6308 VDDA.n796 VDDA.n661 0.028198
R6309 VDDA.n792 VDDA.n660 0.028198
R6310 VDDA.n782 VDDA.n658 0.028198
R6311 VDDA.n776 VDDA.n657 0.028198
R6312 VDDA.n766 VDDA.n655 0.028198
R6313 VDDA.n762 VDDA.n654 0.028198
R6314 VDDA.n752 VDDA.n652 0.028198
R6315 VDDA.n746 VDDA.n651 0.028198
R6316 VDDA.n736 VDDA.n649 0.028198
R6317 VDDA.n732 VDDA.n648 0.028198
R6318 VDDA.n722 VDDA.n646 0.028198
R6319 VDDA.n716 VDDA.n645 0.028198
R6320 VDDA.n706 VDDA.n643 0.028198
R6321 VDDA.n702 VDDA.n642 0.028198
R6322 VDDA.n692 VDDA.n640 0.028198
R6323 VDDA.n686 VDDA.n639 0.028198
R6324 VDDA.n969 VDDA.n968 0.028198
R6325 VDDA.n962 VDDA.n833 0.028198
R6326 VDDA.n954 VDDA.n831 0.028198
R6327 VDDA.n843 VDDA.n830 0.028198
R6328 VDDA.n847 VDDA.n828 0.028198
R6329 VDDA.n938 VDDA.n827 0.028198
R6330 VDDA.n930 VDDA.n825 0.028198
R6331 VDDA.n855 VDDA.n824 0.028198
R6332 VDDA.n859 VDDA.n822 0.028198
R6333 VDDA.n914 VDDA.n821 0.028198
R6334 VDDA.n906 VDDA.n819 0.028198
R6335 VDDA.n867 VDDA.n818 0.028198
R6336 VDDA.n871 VDDA.n816 0.028198
R6337 VDDA.n890 VDDA.n815 0.028198
R6338 VDDA.n882 VDDA.n813 0.028198
R6339 VDDA.n878 VDDA.n812 0.028198
R6340 VDDA.n1140 VDDA.n1139 0.028198
R6341 VDDA.n1133 VDDA.n1132 0.028198
R6342 VDDA.n1123 VDDA.n1122 0.028198
R6343 VDDA.n1120 VDDA.n1119 0.028198
R6344 VDDA.n1110 VDDA.n1109 0.028198
R6345 VDDA.n1103 VDDA.n1102 0.028198
R6346 VDDA.n1093 VDDA.n1092 0.028198
R6347 VDDA.n1090 VDDA.n1089 0.028198
R6348 VDDA.n1080 VDDA.n1079 0.028198
R6349 VDDA.n1073 VDDA.n1072 0.028198
R6350 VDDA.n1063 VDDA.n1062 0.028198
R6351 VDDA.n1060 VDDA.n1059 0.028198
R6352 VDDA.n1050 VDDA.n1049 0.028198
R6353 VDDA.n1043 VDDA.n1042 0.028198
R6354 VDDA.n1033 VDDA.n1032 0.028198
R6355 VDDA.n1030 VDDA.n1029 0.028198
R6356 VDDA.n620 VDDA.n485 0.028198
R6357 VDDA.n491 VDDA.n484 0.028198
R6358 VDDA.n495 VDDA.n482 0.028198
R6359 VDDA.n604 VDDA.n481 0.028198
R6360 VDDA.n596 VDDA.n479 0.028198
R6361 VDDA.n503 VDDA.n478 0.028198
R6362 VDDA.n507 VDDA.n476 0.028198
R6363 VDDA.n580 VDDA.n475 0.028198
R6364 VDDA.n572 VDDA.n473 0.028198
R6365 VDDA.n515 VDDA.n472 0.028198
R6366 VDDA.n519 VDDA.n470 0.028198
R6367 VDDA.n556 VDDA.n469 0.028198
R6368 VDDA.n548 VDDA.n467 0.028198
R6369 VDDA.n527 VDDA.n466 0.028198
R6370 VDDA.n531 VDDA.n464 0.028198
R6371 VDDA.n532 VDDA.n463 0.028198
R6372 VDDA.n1317 VDDA.n1316 0.028198
R6373 VDDA.n1310 VDDA.n1181 0.028198
R6374 VDDA.n1302 VDDA.n1179 0.028198
R6375 VDDA.n1191 VDDA.n1178 0.028198
R6376 VDDA.n1195 VDDA.n1176 0.028198
R6377 VDDA.n1286 VDDA.n1175 0.028198
R6378 VDDA.n1278 VDDA.n1173 0.028198
R6379 VDDA.n1203 VDDA.n1172 0.028198
R6380 VDDA.n1207 VDDA.n1170 0.028198
R6381 VDDA.n1262 VDDA.n1169 0.028198
R6382 VDDA.n1254 VDDA.n1167 0.028198
R6383 VDDA.n1215 VDDA.n1166 0.028198
R6384 VDDA.n1219 VDDA.n1164 0.028198
R6385 VDDA.n1238 VDDA.n1163 0.028198
R6386 VDDA.n1230 VDDA.n1161 0.028198
R6387 VDDA.n1226 VDDA.n1160 0.028198
R6388 VDDA.n2248 VDDA.n1341 0.028198
R6389 VDDA.n2244 VDDA.n1340 0.028198
R6390 VDDA.n2234 VDDA.n1338 0.028198
R6391 VDDA.n2228 VDDA.n1337 0.028198
R6392 VDDA.n2218 VDDA.n1335 0.028198
R6393 VDDA.n2214 VDDA.n1334 0.028198
R6394 VDDA.n2204 VDDA.n1332 0.028198
R6395 VDDA.n2198 VDDA.n1331 0.028198
R6396 VDDA.n2188 VDDA.n1329 0.028198
R6397 VDDA.n2184 VDDA.n1328 0.028198
R6398 VDDA.n2174 VDDA.n1326 0.028198
R6399 VDDA.n2168 VDDA.n1325 0.028198
R6400 VDDA.n2158 VDDA.n1323 0.028198
R6401 VDDA.n2154 VDDA.n1322 0.028198
R6402 VDDA.n2144 VDDA.n1320 0.028198
R6403 VDDA.n2138 VDDA.n1319 0.028198
R6404 VDDA.n2580 VDDA.n2579 0.028198
R6405 VDDA.n2573 VDDA.n2572 0.028198
R6406 VDDA.n2563 VDDA.n2562 0.028198
R6407 VDDA.n2560 VDDA.n2559 0.028198
R6408 VDDA.n2550 VDDA.n2549 0.028198
R6409 VDDA.n2543 VDDA.n2542 0.028198
R6410 VDDA.n2533 VDDA.n2532 0.028198
R6411 VDDA.n2530 VDDA.n2529 0.028198
R6412 VDDA.n2520 VDDA.n2519 0.028198
R6413 VDDA.n2513 VDDA.n2512 0.028198
R6414 VDDA.n2503 VDDA.n2502 0.028198
R6415 VDDA.n2500 VDDA.n2499 0.028198
R6416 VDDA.n2490 VDDA.n2489 0.028198
R6417 VDDA.n2483 VDDA.n2482 0.028198
R6418 VDDA.n2473 VDDA.n2472 0.028198
R6419 VDDA.n2470 VDDA.n2469 0.028198
R6420 VDDA.n354 VDDA.n219 0.028198
R6421 VDDA.n225 VDDA.n218 0.028198
R6422 VDDA.n229 VDDA.n216 0.028198
R6423 VDDA.n338 VDDA.n215 0.028198
R6424 VDDA.n330 VDDA.n213 0.028198
R6425 VDDA.n237 VDDA.n212 0.028198
R6426 VDDA.n241 VDDA.n210 0.028198
R6427 VDDA.n314 VDDA.n209 0.028198
R6428 VDDA.n306 VDDA.n207 0.028198
R6429 VDDA.n249 VDDA.n206 0.028198
R6430 VDDA.n253 VDDA.n204 0.028198
R6431 VDDA.n290 VDDA.n203 0.028198
R6432 VDDA.n282 VDDA.n201 0.028198
R6433 VDDA.n261 VDDA.n200 0.028198
R6434 VDDA.n265 VDDA.n198 0.028198
R6435 VDDA.n266 VDDA.n197 0.028198
R6436 VDDA.n2757 VDDA.n2756 0.028198
R6437 VDDA.n2750 VDDA.n2621 0.028198
R6438 VDDA.n2742 VDDA.n2619 0.028198
R6439 VDDA.n2631 VDDA.n2618 0.028198
R6440 VDDA.n2635 VDDA.n2616 0.028198
R6441 VDDA.n2726 VDDA.n2615 0.028198
R6442 VDDA.n2718 VDDA.n2613 0.028198
R6443 VDDA.n2643 VDDA.n2612 0.028198
R6444 VDDA.n2647 VDDA.n2610 0.028198
R6445 VDDA.n2702 VDDA.n2609 0.028198
R6446 VDDA.n2694 VDDA.n2607 0.028198
R6447 VDDA.n2655 VDDA.n2606 0.028198
R6448 VDDA.n2659 VDDA.n2604 0.028198
R6449 VDDA.n2678 VDDA.n2603 0.028198
R6450 VDDA.n2670 VDDA.n2601 0.028198
R6451 VDDA.n2666 VDDA.n2600 0.028198
R6452 VDDA.n2928 VDDA.n2927 0.028198
R6453 VDDA.n2921 VDDA.n2920 0.028198
R6454 VDDA.n2911 VDDA.n2910 0.028198
R6455 VDDA.n2908 VDDA.n2907 0.028198
R6456 VDDA.n2898 VDDA.n2897 0.028198
R6457 VDDA.n2891 VDDA.n2890 0.028198
R6458 VDDA.n2881 VDDA.n2880 0.028198
R6459 VDDA.n2878 VDDA.n2877 0.028198
R6460 VDDA.n2868 VDDA.n2867 0.028198
R6461 VDDA.n2861 VDDA.n2860 0.028198
R6462 VDDA.n2851 VDDA.n2850 0.028198
R6463 VDDA.n2848 VDDA.n2847 0.028198
R6464 VDDA.n2838 VDDA.n2837 0.028198
R6465 VDDA.n2831 VDDA.n2830 0.028198
R6466 VDDA.n2821 VDDA.n2820 0.028198
R6467 VDDA.n2818 VDDA.n2817 0.028198
R6468 VDDA.n176 VDDA.n41 0.028198
R6469 VDDA.n47 VDDA.n40 0.028198
R6470 VDDA.n51 VDDA.n38 0.028198
R6471 VDDA.n160 VDDA.n37 0.028198
R6472 VDDA.n152 VDDA.n35 0.028198
R6473 VDDA.n59 VDDA.n34 0.028198
R6474 VDDA.n63 VDDA.n32 0.028198
R6475 VDDA.n136 VDDA.n31 0.028198
R6476 VDDA.n128 VDDA.n29 0.028198
R6477 VDDA.n71 VDDA.n28 0.028198
R6478 VDDA.n75 VDDA.n26 0.028198
R6479 VDDA.n112 VDDA.n25 0.028198
R6480 VDDA.n104 VDDA.n23 0.028198
R6481 VDDA.n83 VDDA.n22 0.028198
R6482 VDDA.n87 VDDA.n20 0.028198
R6483 VDDA.n88 VDDA.n19 0.028198
R6484 VDDA.n1573 VDDA.n1431 0.028198
R6485 VDDA.n1569 VDDA.n1430 0.028198
R6486 VDDA.n1559 VDDA.n1428 0.028198
R6487 VDDA.n1553 VDDA.n1427 0.028198
R6488 VDDA.n1543 VDDA.n1425 0.028198
R6489 VDDA.n1539 VDDA.n1424 0.028198
R6490 VDDA.n1529 VDDA.n1422 0.028198
R6491 VDDA.n1523 VDDA.n1421 0.028198
R6492 VDDA.n1513 VDDA.n1419 0.028198
R6493 VDDA.n1509 VDDA.n1418 0.028198
R6494 VDDA.n1499 VDDA.n1416 0.028198
R6495 VDDA.n1493 VDDA.n1415 0.028198
R6496 VDDA.n1483 VDDA.n1413 0.028198
R6497 VDDA.n1479 VDDA.n1412 0.028198
R6498 VDDA.n1469 VDDA.n1410 0.028198
R6499 VDDA.n1463 VDDA.n1409 0.028198
R6500 VDDA.n1806 VDDA.n1345 0.0264451
R6501 VDDA.n1820 VDDA.n1348 0.0264451
R6502 VDDA.n1836 VDDA.n1351 0.0264451
R6503 VDDA.n1850 VDDA.n1354 0.0264451
R6504 VDDA.n1866 VDDA.n1357 0.0264451
R6505 VDDA.n1880 VDDA.n1360 0.0264451
R6506 VDDA.n1896 VDDA.n1363 0.0264451
R6507 VDDA.n1891 VDDA.n1363 0.0264451
R6508 VDDA.n1877 VDDA.n1360 0.0264451
R6509 VDDA.n1861 VDDA.n1357 0.0264451
R6510 VDDA.n1847 VDDA.n1354 0.0264451
R6511 VDDA.n1831 VDDA.n1351 0.0264451
R6512 VDDA.n1817 VDDA.n1348 0.0264451
R6513 VDDA.n1801 VDDA.n1345 0.0264451
R6514 VDDA.n3052 VDDA.n2946 0.0245875
R6515 VDDA.n1478 VDDA.n1411 0.0243392
R6516 VDDA.n1492 VDDA.n1414 0.0243392
R6517 VDDA.n1508 VDDA.n1417 0.0243392
R6518 VDDA.n1522 VDDA.n1420 0.0243392
R6519 VDDA.n1538 VDDA.n1423 0.0243392
R6520 VDDA.n1552 VDDA.n1426 0.0243392
R6521 VDDA.n1568 VDDA.n1429 0.0243392
R6522 VDDA.n2153 VDDA.n1321 0.0243392
R6523 VDDA.n2167 VDDA.n1324 0.0243392
R6524 VDDA.n2183 VDDA.n1327 0.0243392
R6525 VDDA.n2197 VDDA.n1330 0.0243392
R6526 VDDA.n2213 VDDA.n1333 0.0243392
R6527 VDDA.n2227 VDDA.n1336 0.0243392
R6528 VDDA.n2243 VDDA.n1339 0.0243392
R6529 VDDA.n82 VDDA.n21 0.0243392
R6530 VDDA.n111 VDDA.n24 0.0243392
R6531 VDDA.n70 VDDA.n27 0.0243392
R6532 VDDA.n135 VDDA.n30 0.0243392
R6533 VDDA.n58 VDDA.n33 0.0243392
R6534 VDDA.n159 VDDA.n36 0.0243392
R6535 VDDA.n46 VDDA.n39 0.0243392
R6536 VDDA.n2829 VDDA.n2828 0.0243392
R6537 VDDA.n2840 VDDA.n2802 0.0243392
R6538 VDDA.n2859 VDDA.n2858 0.0243392
R6539 VDDA.n2870 VDDA.n2790 0.0243392
R6540 VDDA.n2889 VDDA.n2888 0.0243392
R6541 VDDA.n2900 VDDA.n2778 0.0243392
R6542 VDDA.n2919 VDDA.n2918 0.0243392
R6543 VDDA.n2677 VDDA.n2602 0.0243392
R6544 VDDA.n2654 VDDA.n2605 0.0243392
R6545 VDDA.n2701 VDDA.n2608 0.0243392
R6546 VDDA.n2642 VDDA.n2611 0.0243392
R6547 VDDA.n2725 VDDA.n2614 0.0243392
R6548 VDDA.n2630 VDDA.n2617 0.0243392
R6549 VDDA.n2749 VDDA.n2620 0.0243392
R6550 VDDA.n260 VDDA.n199 0.0243392
R6551 VDDA.n289 VDDA.n202 0.0243392
R6552 VDDA.n248 VDDA.n205 0.0243392
R6553 VDDA.n313 VDDA.n208 0.0243392
R6554 VDDA.n236 VDDA.n211 0.0243392
R6555 VDDA.n337 VDDA.n214 0.0243392
R6556 VDDA.n224 VDDA.n217 0.0243392
R6557 VDDA.n2481 VDDA.n2480 0.0243392
R6558 VDDA.n2492 VDDA.n2454 0.0243392
R6559 VDDA.n2511 VDDA.n2510 0.0243392
R6560 VDDA.n2522 VDDA.n2442 0.0243392
R6561 VDDA.n2541 VDDA.n2540 0.0243392
R6562 VDDA.n2552 VDDA.n2430 0.0243392
R6563 VDDA.n2571 VDDA.n2570 0.0243392
R6564 VDDA.n1237 VDDA.n1162 0.0243392
R6565 VDDA.n1214 VDDA.n1165 0.0243392
R6566 VDDA.n1261 VDDA.n1168 0.0243392
R6567 VDDA.n1202 VDDA.n1171 0.0243392
R6568 VDDA.n1285 VDDA.n1174 0.0243392
R6569 VDDA.n1190 VDDA.n1177 0.0243392
R6570 VDDA.n1309 VDDA.n1180 0.0243392
R6571 VDDA.n526 VDDA.n465 0.0243392
R6572 VDDA.n555 VDDA.n468 0.0243392
R6573 VDDA.n514 VDDA.n471 0.0243392
R6574 VDDA.n579 VDDA.n474 0.0243392
R6575 VDDA.n502 VDDA.n477 0.0243392
R6576 VDDA.n603 VDDA.n480 0.0243392
R6577 VDDA.n490 VDDA.n483 0.0243392
R6578 VDDA.n1041 VDDA.n1040 0.0243392
R6579 VDDA.n1052 VDDA.n1014 0.0243392
R6580 VDDA.n1071 VDDA.n1070 0.0243392
R6581 VDDA.n1082 VDDA.n1002 0.0243392
R6582 VDDA.n1101 VDDA.n1100 0.0243392
R6583 VDDA.n1112 VDDA.n990 0.0243392
R6584 VDDA.n1131 VDDA.n1130 0.0243392
R6585 VDDA.n889 VDDA.n814 0.0243392
R6586 VDDA.n866 VDDA.n817 0.0243392
R6587 VDDA.n913 VDDA.n820 0.0243392
R6588 VDDA.n854 VDDA.n823 0.0243392
R6589 VDDA.n937 VDDA.n826 0.0243392
R6590 VDDA.n842 VDDA.n829 0.0243392
R6591 VDDA.n961 VDDA.n832 0.0243392
R6592 VDDA.n701 VDDA.n641 0.0243392
R6593 VDDA.n715 VDDA.n644 0.0243392
R6594 VDDA.n731 VDDA.n647 0.0243392
R6595 VDDA.n745 VDDA.n650 0.0243392
R6596 VDDA.n761 VDDA.n653 0.0243392
R6597 VDDA.n775 VDDA.n656 0.0243392
R6598 VDDA.n791 VDDA.n659 0.0243392
R6599 VDDA.n786 VDDA.n659 0.0243392
R6600 VDDA.n772 VDDA.n656 0.0243392
R6601 VDDA.n756 VDDA.n653 0.0243392
R6602 VDDA.n742 VDDA.n650 0.0243392
R6603 VDDA.n726 VDDA.n647 0.0243392
R6604 VDDA.n712 VDDA.n644 0.0243392
R6605 VDDA.n696 VDDA.n641 0.0243392
R6606 VDDA.n839 VDDA.n832 0.0243392
R6607 VDDA.n946 VDDA.n829 0.0243392
R6608 VDDA.n851 VDDA.n826 0.0243392
R6609 VDDA.n922 VDDA.n823 0.0243392
R6610 VDDA.n863 VDDA.n820 0.0243392
R6611 VDDA.n898 VDDA.n817 0.0243392
R6612 VDDA.n875 VDDA.n814 0.0243392
R6613 VDDA.n1130 VDDA.n1129 0.0243392
R6614 VDDA.n1113 VDDA.n1112 0.0243392
R6615 VDDA.n1100 VDDA.n1099 0.0243392
R6616 VDDA.n1083 VDDA.n1082 0.0243392
R6617 VDDA.n1070 VDDA.n1069 0.0243392
R6618 VDDA.n1053 VDDA.n1052 0.0243392
R6619 VDDA.n1040 VDDA.n1039 0.0243392
R6620 VDDA.n612 VDDA.n483 0.0243392
R6621 VDDA.n499 VDDA.n480 0.0243392
R6622 VDDA.n588 VDDA.n477 0.0243392
R6623 VDDA.n511 VDDA.n474 0.0243392
R6624 VDDA.n564 VDDA.n471 0.0243392
R6625 VDDA.n523 VDDA.n468 0.0243392
R6626 VDDA.n540 VDDA.n465 0.0243392
R6627 VDDA.n1187 VDDA.n1180 0.0243392
R6628 VDDA.n1294 VDDA.n1177 0.0243392
R6629 VDDA.n1199 VDDA.n1174 0.0243392
R6630 VDDA.n1270 VDDA.n1171 0.0243392
R6631 VDDA.n1211 VDDA.n1168 0.0243392
R6632 VDDA.n1246 VDDA.n1165 0.0243392
R6633 VDDA.n1223 VDDA.n1162 0.0243392
R6634 VDDA.n2238 VDDA.n1339 0.0243392
R6635 VDDA.n2224 VDDA.n1336 0.0243392
R6636 VDDA.n2208 VDDA.n1333 0.0243392
R6637 VDDA.n2194 VDDA.n1330 0.0243392
R6638 VDDA.n2178 VDDA.n1327 0.0243392
R6639 VDDA.n2164 VDDA.n1324 0.0243392
R6640 VDDA.n2148 VDDA.n1321 0.0243392
R6641 VDDA.n2570 VDDA.n2569 0.0243392
R6642 VDDA.n2553 VDDA.n2552 0.0243392
R6643 VDDA.n2540 VDDA.n2539 0.0243392
R6644 VDDA.n2523 VDDA.n2522 0.0243392
R6645 VDDA.n2510 VDDA.n2509 0.0243392
R6646 VDDA.n2493 VDDA.n2492 0.0243392
R6647 VDDA.n2480 VDDA.n2479 0.0243392
R6648 VDDA.n346 VDDA.n217 0.0243392
R6649 VDDA.n233 VDDA.n214 0.0243392
R6650 VDDA.n322 VDDA.n211 0.0243392
R6651 VDDA.n245 VDDA.n208 0.0243392
R6652 VDDA.n298 VDDA.n205 0.0243392
R6653 VDDA.n257 VDDA.n202 0.0243392
R6654 VDDA.n274 VDDA.n199 0.0243392
R6655 VDDA.n2627 VDDA.n2620 0.0243392
R6656 VDDA.n2734 VDDA.n2617 0.0243392
R6657 VDDA.n2639 VDDA.n2614 0.0243392
R6658 VDDA.n2710 VDDA.n2611 0.0243392
R6659 VDDA.n2651 VDDA.n2608 0.0243392
R6660 VDDA.n2686 VDDA.n2605 0.0243392
R6661 VDDA.n2663 VDDA.n2602 0.0243392
R6662 VDDA.n2918 VDDA.n2917 0.0243392
R6663 VDDA.n2901 VDDA.n2900 0.0243392
R6664 VDDA.n2888 VDDA.n2887 0.0243392
R6665 VDDA.n2871 VDDA.n2870 0.0243392
R6666 VDDA.n2858 VDDA.n2857 0.0243392
R6667 VDDA.n2841 VDDA.n2840 0.0243392
R6668 VDDA.n2828 VDDA.n2827 0.0243392
R6669 VDDA.n168 VDDA.n39 0.0243392
R6670 VDDA.n55 VDDA.n36 0.0243392
R6671 VDDA.n144 VDDA.n33 0.0243392
R6672 VDDA.n67 VDDA.n30 0.0243392
R6673 VDDA.n120 VDDA.n27 0.0243392
R6674 VDDA.n79 VDDA.n24 0.0243392
R6675 VDDA.n96 VDDA.n21 0.0243392
R6676 VDDA.n1563 VDDA.n1429 0.0243392
R6677 VDDA.n1549 VDDA.n1426 0.0243392
R6678 VDDA.n1533 VDDA.n1423 0.0243392
R6679 VDDA.n1519 VDDA.n1420 0.0243392
R6680 VDDA.n1503 VDDA.n1417 0.0243392
R6681 VDDA.n1489 VDDA.n1414 0.0243392
R6682 VDDA.n1473 VDDA.n1411 0.0243392
R6683 VDDA.n2130 VDDA.n1931 0.0217373
R6684 VDDA.n2080 VDDA.n1933 0.0217373
R6685 VDDA.n2003 VDDA.n1935 0.0217373
R6686 VDDA.n1942 VDDA.n1937 0.0217373
R6687 VDDA.n1946 VDDA.n1945 0.0217373
R6688 VDDA.n2007 VDDA.n2006 0.0217373
R6689 VDDA.n2084 VDDA.n2083 0.0217373
R6690 VDDA.n2134 VDDA.n2133 0.0217373
R6691 VDDA.n1944 VDDA.n1937 0.0217373
R6692 VDDA.n1947 VDDA.n1946 0.0217373
R6693 VDDA.n2005 VDDA.n1935 0.0217373
R6694 VDDA.n2008 VDDA.n2007 0.0217373
R6695 VDDA.n2082 VDDA.n1933 0.0217373
R6696 VDDA.n2085 VDDA.n2084 0.0217373
R6697 VDDA.n2132 VDDA.n1931 0.0217373
R6698 VDDA.n2135 VDDA.n2134 0.0217373
R6699 VDDA.n2942 VDDA.n2941 0.0217373
R6700 VDDA.n2939 VDDA.n183 0.0217373
R6701 VDDA.n2933 VDDA.n185 0.0217373
R6702 VDDA.n2936 VDDA.n186 0.0217373
R6703 VDDA.n2762 VDDA.n188 0.0217373
R6704 VDDA.n2765 VDDA.n189 0.0217373
R6705 VDDA.n2594 VDDA.n2593 0.0217373
R6706 VDDA.n2590 VDDA.n360 0.0217373
R6707 VDDA.n2585 VDDA.n362 0.0217373
R6708 VDDA.n2588 VDDA.n363 0.0217373
R6709 VDDA.n2258 VDDA.n454 0.0217373
R6710 VDDA.n2261 VDDA.n455 0.0217373
R6711 VDDA.n424 VDDA.n412 0.0217373
R6712 VDDA.n435 VDDA.n429 0.0217373
R6713 VDDA.n385 VDDA.n368 0.0217373
R6714 VDDA.n385 VDDA.n367 0.0217373
R6715 VDDA.n2395 VDDA.n2394 0.0217373
R6716 VDDA.n2392 VDDA.n404 0.0217373
R6717 VDDA.n427 VDDA.n406 0.0217373
R6718 VDDA.n411 VDDA.n409 0.0217373
R6719 VDDA.n429 VDDA.n407 0.0217373
R6720 VDDA.n428 VDDA.n427 0.0217373
R6721 VDDA.n412 VDDA.n410 0.0217373
R6722 VDDA.n2342 VDDA.n447 0.0217373
R6723 VDDA.n2394 VDDA.n387 0.0217373
R6724 VDDA.n404 VDDA.n387 0.0217373
R6725 VDDA.n2286 VDDA.n449 0.0217373
R6726 VDDA.n2337 VDDA.n448 0.0217373
R6727 VDDA.n2331 VDDA.n2304 0.0217373
R6728 VDDA.n2321 VDDA.n2307 0.0217373
R6729 VDDA.n2287 VDDA.n447 0.0217373
R6730 VDDA.n2337 VDDA.n2336 0.0217373
R6731 VDDA.n2333 VDDA.n2305 0.0217373
R6732 VDDA.n2332 VDDA.n2331 0.0217373
R6733 VDDA.n2322 VDDA.n2308 0.0217373
R6734 VDDA.n1154 VDDA.n1153 0.0217373
R6735 VDDA.n1150 VDDA.n626 0.0217373
R6736 VDDA.n1145 VDDA.n628 0.0217373
R6737 VDDA.n1148 VDDA.n629 0.0217373
R6738 VDDA.n974 VDDA.n631 0.0217373
R6739 VDDA.n977 VDDA.n632 0.0217373
R6740 VDDA.n802 VDDA.n633 0.0217373
R6741 VDDA.n2397 VDDA.n366 0.0217373
R6742 VDDA.n634 VDDA.n631 0.0217373
R6743 VDDA.n634 VDDA.n632 0.0217373
R6744 VDDA.n979 VDDA.n628 0.0217373
R6745 VDDA.n979 VDDA.n629 0.0217373
R6746 VDDA.n1153 VDDA.n1152 0.0217373
R6747 VDDA.n1152 VDDA.n626 0.0217373
R6748 VDDA.n2283 VDDA.n2281 0.0217373
R6749 VDDA.n2281 VDDA.n449 0.0217373
R6750 VDDA.n2399 VDDA.n368 0.0217373
R6751 VDDA.n2396 VDDA.n367 0.0217373
R6752 VDDA.n2398 VDDA.n2397 0.0217373
R6753 VDDA.n457 VDDA.n454 0.0217373
R6754 VDDA.n457 VDDA.n455 0.0217373
R6755 VDDA.n2419 VDDA.n362 0.0217373
R6756 VDDA.n2419 VDDA.n363 0.0217373
R6757 VDDA.n2593 VDDA.n2592 0.0217373
R6758 VDDA.n2592 VDDA.n360 0.0217373
R6759 VDDA.n191 VDDA.n188 0.0217373
R6760 VDDA.n191 VDDA.n189 0.0217373
R6761 VDDA.n2767 VDDA.n185 0.0217373
R6762 VDDA.n2767 VDDA.n186 0.0217373
R6763 VDDA.n2941 VDDA.n181 0.0217373
R6764 VDDA.n183 VDDA.n181 0.0217373
R6765 VDDA.n804 VDDA.n803 0.0217373
R6766 VDDA.n802 VDDA.n801 0.0217373
R6767 VDDA.n2132 VDDA.n1932 0.0217373
R6768 VDDA.n2082 VDDA.n1934 0.0217373
R6769 VDDA.n2005 VDDA.n1936 0.0217373
R6770 VDDA.n1944 VDDA.n1938 0.0217373
R6771 VDDA.n1945 VDDA.n1943 0.0217373
R6772 VDDA.n2006 VDDA.n2004 0.0217373
R6773 VDDA.n2083 VDDA.n2081 0.0217373
R6774 VDDA.n2133 VDDA.n2131 0.0217373
R6775 VDDA.n2004 VDDA.n1948 0.0217373
R6776 VDDA.n2081 VDDA.n2009 0.0217373
R6777 VDDA.n2131 VDDA.n2086 0.0217373
R6778 VDDA.n2308 VDDA.n2306 0.0217373
R6779 VDDA.n2305 VDDA.n2303 0.0217373
R6780 VDDA.n410 VDDA.n408 0.0217373
R6781 VDDA.n407 VDDA.n405 0.0217373
R6782 VDDA.n436 VDDA.n406 0.0217373
R6783 VDDA.n425 VDDA.n409 0.0217373
R6784 VDDA.n437 VDDA.n436 0.0217373
R6785 VDDA.n426 VDDA.n425 0.0217373
R6786 VDDA.n2339 VDDA.n2287 0.0217373
R6787 VDDA.n2391 VDDA.n386 0.0217373
R6788 VDDA.n388 VDDA.n386 0.0217373
R6789 VDDA.n2341 VDDA.n448 0.0217373
R6790 VDDA.n2334 VDDA.n2304 0.0217373
R6791 VDDA.n2323 VDDA.n2307 0.0217373
R6792 VDDA.n2341 VDDA.n2340 0.0217373
R6793 VDDA.n2339 VDDA.n2338 0.0217373
R6794 VDDA.n2335 VDDA.n2334 0.0217373
R6795 VDDA.n2330 VDDA.n2303 0.0217373
R6796 VDDA.n2324 VDDA.n2323 0.0217373
R6797 VDDA.n2320 VDDA.n2306 0.0217373
R6798 VDDA.n801 VDDA.n800 0.0217373
R6799 VDDA.n976 VDDA.n975 0.0217373
R6800 VDDA.n1147 VDDA.n1146 0.0217373
R6801 VDDA.n1151 VDDA.n624 0.0217373
R6802 VDDA.n2260 VDDA.n2259 0.0217373
R6803 VDDA.n2285 VDDA.n2284 0.0217373
R6804 VDDA.n2587 VDDA.n2586 0.0217373
R6805 VDDA.n2591 VDDA.n358 0.0217373
R6806 VDDA.n2764 VDDA.n2763 0.0217373
R6807 VDDA.n2935 VDDA.n2934 0.0217373
R6808 VDDA.n2938 VDDA.n180 0.0217373
R6809 VDDA.n975 VDDA.n630 0.0217373
R6810 VDDA.n1146 VDDA.n627 0.0217373
R6811 VDDA.n625 VDDA.n624 0.0217373
R6812 VDDA.n2284 VDDA.n2282 0.0217373
R6813 VDDA.n2259 VDDA.n453 0.0217373
R6814 VDDA.n2586 VDDA.n361 0.0217373
R6815 VDDA.n359 VDDA.n358 0.0217373
R6816 VDDA.n2763 VDDA.n187 0.0217373
R6817 VDDA.n2934 VDDA.n184 0.0217373
R6818 VDDA.n182 VDDA.n180 0.0217373
R6819 VDDA.n805 VDDA.n804 0.0217373
R6820 VDDA.n806 VDDA.n805 0.0217373
R6821 VDDA.n1759 VDDA.n1758 0.0152446
R6822 VDDA.n1757 VDDA.n1756 0.0152446
R6823 VDDA.n1755 VDDA.n1754 0.0152446
R6824 VDDA.n1745 VDDA.n1744 0.0152446
R6825 VDDA.n1592 VDDA.n1588 0.0152446
R6826 VDDA.n1738 VDDA.n1593 0.0152446
R6827 VDDA.n1728 VDDA.n1599 0.0152446
R6828 VDDA.n1727 VDDA.n1726 0.0152446
R6829 VDDA.n1725 VDDA.n1724 0.0152446
R6830 VDDA.n1715 VDDA.n1714 0.0152446
R6831 VDDA.n1610 VDDA.n1606 0.0152446
R6832 VDDA.n1708 VDDA.n1611 0.0152446
R6833 VDDA.n1698 VDDA.n1617 0.0152446
R6834 VDDA.n1697 VDDA.n1696 0.0152446
R6835 VDDA.n1695 VDDA.n1694 0.0152446
R6836 VDDA.n1685 VDDA.n1684 0.0152446
R6837 VDDA.n1628 VDDA.n1624 0.0152446
R6838 VDDA.n1678 VDDA.n1629 0.0152446
R6839 VDDA.n1668 VDDA.n1635 0.0152446
R6840 VDDA.n1667 VDDA.n1666 0.0152446
R6841 VDDA.n1665 VDDA.n1664 0.0152446
R6842 VDDA.n1655 VDDA.n1654 0.0152446
R6843 VDDA.n1645 VDDA.n1642 0.0152446
R6844 VDDA.n1648 VDDA.n1646 0.0152446
R6845 VDDA.n1646 VDDA.n1645 0.0152446
R6846 VDDA.n1654 VDDA.n1642 0.0152446
R6847 VDDA.n1656 VDDA.n1655 0.0152446
R6848 VDDA.n1666 VDDA.n1665 0.0152446
R6849 VDDA.n1668 VDDA.n1667 0.0152446
R6850 VDDA.n1635 VDDA.n1634 0.0152446
R6851 VDDA.n1629 VDDA.n1628 0.0152446
R6852 VDDA.n1684 VDDA.n1624 0.0152446
R6853 VDDA.n1686 VDDA.n1685 0.0152446
R6854 VDDA.n1696 VDDA.n1695 0.0152446
R6855 VDDA.n1698 VDDA.n1697 0.0152446
R6856 VDDA.n1617 VDDA.n1616 0.0152446
R6857 VDDA.n1611 VDDA.n1610 0.0152446
R6858 VDDA.n1714 VDDA.n1606 0.0152446
R6859 VDDA.n1716 VDDA.n1715 0.0152446
R6860 VDDA.n1726 VDDA.n1725 0.0152446
R6861 VDDA.n1728 VDDA.n1727 0.0152446
R6862 VDDA.n1599 VDDA.n1598 0.0152446
R6863 VDDA.n1593 VDDA.n1592 0.0152446
R6864 VDDA.n1744 VDDA.n1588 0.0152446
R6865 VDDA.n1746 VDDA.n1745 0.0152446
R6866 VDDA.n1756 VDDA.n1755 0.0152446
R6867 VDDA.n1758 VDDA.n1757 0.0152446
R6868 VDDA.n1760 VDDA.n1759 0.0152446
R6869 VDDA.n1760 VDDA.n1406 0.0142311
R6870 VDDA.n1586 VDDA.n1581 0.0142311
R6871 VDDA.n1747 VDDA.n1746 0.0142311
R6872 VDDA.n1737 VDDA.n1736 0.0142311
R6873 VDDA.n1598 VDDA.n1594 0.0142311
R6874 VDDA.n1604 VDDA.n1600 0.0142311
R6875 VDDA.n1717 VDDA.n1716 0.0142311
R6876 VDDA.n1707 VDDA.n1706 0.0142311
R6877 VDDA.n1616 VDDA.n1612 0.0142311
R6878 VDDA.n1622 VDDA.n1618 0.0142311
R6879 VDDA.n1687 VDDA.n1686 0.0142311
R6880 VDDA.n1677 VDDA.n1676 0.0142311
R6881 VDDA.n1634 VDDA.n1630 0.0142311
R6882 VDDA.n1640 VDDA.n1636 0.0142311
R6883 VDDA.n1657 VDDA.n1656 0.0142311
R6884 VDDA.n1647 VDDA.n1644 0.0142311
R6885 VDDA.n1648 VDDA.n1647 0.0142311
R6886 VDDA.n1658 VDDA.n1657 0.0142311
R6887 VDDA.n1664 VDDA.n1636 0.0142311
R6888 VDDA.n1674 VDDA.n1630 0.0142311
R6889 VDDA.n1678 VDDA.n1677 0.0142311
R6890 VDDA.n1688 VDDA.n1687 0.0142311
R6891 VDDA.n1694 VDDA.n1618 0.0142311
R6892 VDDA.n1704 VDDA.n1612 0.0142311
R6893 VDDA.n1708 VDDA.n1707 0.0142311
R6894 VDDA.n1718 VDDA.n1717 0.0142311
R6895 VDDA.n1724 VDDA.n1600 0.0142311
R6896 VDDA.n1734 VDDA.n1594 0.0142311
R6897 VDDA.n1738 VDDA.n1737 0.0142311
R6898 VDDA.n1748 VDDA.n1747 0.0142311
R6899 VDDA.n1754 VDDA.n1581 0.0142311
R6900 VDDA.n1407 VDDA.n1406 0.0142311
R6901 VDDA.n1748 VDDA.n1587 0.0132169
R6902 VDDA.n1735 VDDA.n1734 0.0132169
R6903 VDDA.n1718 VDDA.n1605 0.0132169
R6904 VDDA.n1705 VDDA.n1704 0.0132169
R6905 VDDA.n1688 VDDA.n1623 0.0132169
R6906 VDDA.n1675 VDDA.n1674 0.0132169
R6907 VDDA.n1658 VDDA.n1641 0.0132169
R6908 VDDA.n1641 VDDA.n1640 0.0132169
R6909 VDDA.n1676 VDDA.n1675 0.0132169
R6910 VDDA.n1623 VDDA.n1622 0.0132169
R6911 VDDA.n1706 VDDA.n1705 0.0132169
R6912 VDDA.n1605 VDDA.n1604 0.0132169
R6913 VDDA.n1736 VDDA.n1735 0.0132169
R6914 VDDA.n1587 VDDA.n1586 0.0132169
R6915 VDDA.n1579 VDDA.n1578 0.0129844
R6916 VDDA.n2254 VDDA.n1158 0.0107812
R6917 VDDA.n2598 VDDA.n195 0.0107812
R6918 VDDA.n1578 VDDA.n195 0.0101203
R6919 VDDA.n2254 VDDA.n2253 0.0099
R6920 VDDA VDDA.n3053 0.00879844
R6921 VDDA.n970 VDDA.n810 0.00564062
R6922 VDDA.n970 VDDA.n461 0.00564062
R6923 VDDA.n1158 VDDA.n461 0.00564062
R6924 VDDA.n2758 VDDA.n2598 0.00564062
R6925 VDDA.n2758 VDDA.n17 0.00564062
R6926 VDDA.n2946 VDDA.n17 0.00564062
R6927 VDDA.n1906 VDDA.n1366 0.00211562
R6928 VDDA.n3052 VDDA.n2962 0.00189531
R6929 VDDA.n2962 VDDA.n16 0.00189531
R6930 VDDA.n3011 VDDA.n3 0.00188102
R6931 VDDA.n3015 VDDA.n7 0.00188102
R6932 VDDA.n3019 VDDA.n11 0.00188102
R6933 VDDA.n2966 VDDA.n2960 0.00188102
R6934 VDDA.n2972 VDDA.n2958 0.00188102
R6935 VDDA.n2978 VDDA.n2956 0.00188102
R6936 VDDA.n2984 VDDA.n2954 0.00188102
R6937 VDDA.n2990 VDDA.n2952 0.00188102
R6938 VDDA.n2996 VDDA.n2950 0.00188102
R6939 VDDA.n3002 VDDA.n2948 0.00188102
R6940 VDDA.n3030 VDDA.n11 0.00188102
R6941 VDDA.n3038 VDDA.n7 0.00188102
R6942 VDDA.n3046 VDDA.n3 0.00188102
R6943 VDDA.n2967 VDDA.n2966 0.00188102
R6944 VDDA.n2973 VDDA.n2972 0.00188102
R6945 VDDA.n2979 VDDA.n2978 0.00188102
R6946 VDDA.n2985 VDDA.n2984 0.00188102
R6947 VDDA.n2991 VDDA.n2990 0.00188102
R6948 VDDA.n2997 VDDA.n2996 0.00188102
R6949 VDDA.n3003 VDDA.n3002 0.00188102
R6950 VDDA.n3009 VDDA.n3008 0.00173422
R6951 VDDA.n3009 VDDA.n1 0.00173422
R6952 VDDA.n3049 VDDA.n3010 0.00173422
R6953 VDDA.n3043 VDDA.n3013 0.00173422
R6954 VDDA.n3013 VDDA.n5 0.00173422
R6955 VDDA.n3041 VDDA.n3014 0.00173422
R6956 VDDA.n3035 VDDA.n3017 0.00173422
R6957 VDDA.n3017 VDDA.n9 0.00173422
R6958 VDDA.n3033 VDDA.n3018 0.00173422
R6959 VDDA.n3027 VDDA.n3021 0.00173422
R6960 VDDA.n3021 VDDA.n13 0.00173422
R6961 VDDA.n3025 VDDA.n3022 0.00173422
R6962 VDDA.n2963 VDDA.n2961 0.00173422
R6963 VDDA.n2969 VDDA.n2959 0.00173422
R6964 VDDA.n2975 VDDA.n2957 0.00173422
R6965 VDDA.n2981 VDDA.n2955 0.00173422
R6966 VDDA.n2987 VDDA.n2953 0.00173422
R6967 VDDA.n2993 VDDA.n2951 0.00173422
R6968 VDDA.n2999 VDDA.n2949 0.00173422
R6969 VDDA.n3005 VDDA.n2947 0.00173422
R6970 VDDA.n3026 VDDA.n13 0.00173422
R6971 VDDA.n3034 VDDA.n9 0.00173422
R6972 VDDA.n3042 VDDA.n5 0.00173422
R6973 VDDA.n3050 VDDA.n1 0.00173422
R6974 VDDA.n2964 VDDA.n2963 0.00173422
R6975 VDDA.n3026 VDDA.n3025 0.00173422
R6976 VDDA.n3028 VDDA.n3027 0.00173422
R6977 VDDA.n3034 VDDA.n3033 0.00173422
R6978 VDDA.n3036 VDDA.n3035 0.00173422
R6979 VDDA.n3042 VDDA.n3041 0.00173422
R6980 VDDA.n3044 VDDA.n3043 0.00173422
R6981 VDDA.n3050 VDDA.n3049 0.00173422
R6982 VDDA.n3008 VDDA.n16 0.00173422
R6983 VDDA.n2970 VDDA.n2969 0.00173422
R6984 VDDA.n2976 VDDA.n2975 0.00173422
R6985 VDDA.n2982 VDDA.n2981 0.00173422
R6986 VDDA.n2988 VDDA.n2987 0.00173422
R6987 VDDA.n2994 VDDA.n2993 0.00173422
R6988 VDDA.n3000 VDDA.n2999 0.00173422
R6989 VDDA.n3006 VDDA.n3005 0.00173422
R6990 VDDA.n3010 VDDA.n2 0.00169751
R6991 VDDA.n3047 VDDA.n3011 0.00169751
R6992 VDDA.n3045 VDDA.n3012 0.00169751
R6993 VDDA.n3012 VDDA.n4 0.00169751
R6994 VDDA.n3014 VDDA.n6 0.00169751
R6995 VDDA.n3039 VDDA.n3015 0.00169751
R6996 VDDA.n3037 VDDA.n3016 0.00169751
R6997 VDDA.n3016 VDDA.n8 0.00169751
R6998 VDDA.n3018 VDDA.n10 0.00169751
R6999 VDDA.n3031 VDDA.n3019 0.00169751
R7000 VDDA.n3029 VDDA.n3020 0.00169751
R7001 VDDA.n3020 VDDA.n12 0.00169751
R7002 VDDA.n3022 VDDA.n14 0.00169751
R7003 VDDA.n3024 VDDA.n15 0.00169751
R7004 VDDA.n3023 VDDA.n14 0.00169751
R7005 VDDA.n3028 VDDA.n12 0.00169751
R7006 VDDA.n3032 VDDA.n10 0.00169751
R7007 VDDA.n3036 VDDA.n8 0.00169751
R7008 VDDA.n3040 VDDA.n6 0.00169751
R7009 VDDA.n3044 VDDA.n4 0.00169751
R7010 VDDA.n3048 VDDA.n2 0.00169751
R7011 VDDA.n3030 VDDA.n3029 0.00169751
R7012 VDDA.n3032 VDDA.n3031 0.00169751
R7013 VDDA.n3038 VDDA.n3037 0.00169751
R7014 VDDA.n3040 VDDA.n3039 0.00169751
R7015 VDDA.n3046 VDDA.n3045 0.00169751
R7016 VDDA.n3048 VDDA.n3047 0.00169751
R7017 VDDA.n3024 VDDA.n3023 0.00169751
R7018 VDDA.n2964 VDDA.n0 0.00166081
R7019 VDDA.n2967 VDDA.n2965 0.00166081
R7020 VDDA.n2970 VDDA.n2968 0.00166081
R7021 VDDA.n2973 VDDA.n2971 0.00166081
R7022 VDDA.n2976 VDDA.n2974 0.00166081
R7023 VDDA.n2979 VDDA.n2977 0.00166081
R7024 VDDA.n2982 VDDA.n2980 0.00166081
R7025 VDDA.n2985 VDDA.n2983 0.00166081
R7026 VDDA.n2988 VDDA.n2986 0.00166081
R7027 VDDA.n2991 VDDA.n2989 0.00166081
R7028 VDDA.n2994 VDDA.n2992 0.00166081
R7029 VDDA.n2997 VDDA.n2995 0.00166081
R7030 VDDA.n3000 VDDA.n2998 0.00166081
R7031 VDDA.n3003 VDDA.n3001 0.00166081
R7032 VDDA.n3006 VDDA.n3004 0.00166081
R7033 VDDA.n3051 VDDA.n3007 0.00166081
R7034 VDDA.n3053 VDDA.n0 0.00166081
R7035 VDDA.n2965 VDDA.n2961 0.00166081
R7036 VDDA.n2968 VDDA.n2960 0.00166081
R7037 VDDA.n2971 VDDA.n2959 0.00166081
R7038 VDDA.n2974 VDDA.n2958 0.00166081
R7039 VDDA.n2977 VDDA.n2957 0.00166081
R7040 VDDA.n2980 VDDA.n2956 0.00166081
R7041 VDDA.n2983 VDDA.n2955 0.00166081
R7042 VDDA.n2986 VDDA.n2954 0.00166081
R7043 VDDA.n2989 VDDA.n2953 0.00166081
R7044 VDDA.n2992 VDDA.n2952 0.00166081
R7045 VDDA.n2995 VDDA.n2951 0.00166081
R7046 VDDA.n2998 VDDA.n2950 0.00166081
R7047 VDDA.n3001 VDDA.n2949 0.00166081
R7048 VDDA.n3004 VDDA.n2948 0.00166081
R7049 VDDA.n3007 VDDA.n2947 0.00166081
R7050 VDDA.t91 VDDA.n1456 0.00152174
R7051 VDDA.t62 VDDA.n1457 0.00152174
R7052 VDDA.t147 VDDA.n1458 0.00152174
R7053 VDDA.t145 VDDA.n1459 0.00152174
R7054 VDDA.t124 VDDA.n1460 0.00152174
R7055 VDDA.n1579 VDDA.n1366 0.00138125
R7056 two_stage_opamp_dummy_magic_25_0.VD3.n32 two_stage_opamp_dummy_magic_25_0.VD3.t13 672.293
R7057 two_stage_opamp_dummy_magic_25_0.VD3.n42 two_stage_opamp_dummy_magic_25_0.VD3.t10 672.293
R7058 two_stage_opamp_dummy_magic_25_0.VD3.t14 two_stage_opamp_dummy_magic_25_0.VD3.n40 213.131
R7059 two_stage_opamp_dummy_magic_25_0.VD3.n41 two_stage_opamp_dummy_magic_25_0.VD3.t11 213.131
R7060 two_stage_opamp_dummy_magic_25_0.VD3.t20 two_stage_opamp_dummy_magic_25_0.VD3.t14 146.155
R7061 two_stage_opamp_dummy_magic_25_0.VD3.t36 two_stage_opamp_dummy_magic_25_0.VD3.t20 146.155
R7062 two_stage_opamp_dummy_magic_25_0.VD3.t34 two_stage_opamp_dummy_magic_25_0.VD3.t36 146.155
R7063 two_stage_opamp_dummy_magic_25_0.VD3.t4 two_stage_opamp_dummy_magic_25_0.VD3.t34 146.155
R7064 two_stage_opamp_dummy_magic_25_0.VD3.t2 two_stage_opamp_dummy_magic_25_0.VD3.t4 146.155
R7065 two_stage_opamp_dummy_magic_25_0.VD3.t8 two_stage_opamp_dummy_magic_25_0.VD3.t2 146.155
R7066 two_stage_opamp_dummy_magic_25_0.VD3.t18 two_stage_opamp_dummy_magic_25_0.VD3.t8 146.155
R7067 two_stage_opamp_dummy_magic_25_0.VD3.t0 two_stage_opamp_dummy_magic_25_0.VD3.t18 146.155
R7068 two_stage_opamp_dummy_magic_25_0.VD3.t6 two_stage_opamp_dummy_magic_25_0.VD3.t0 146.155
R7069 two_stage_opamp_dummy_magic_25_0.VD3.t16 two_stage_opamp_dummy_magic_25_0.VD3.t6 146.155
R7070 two_stage_opamp_dummy_magic_25_0.VD3.t11 two_stage_opamp_dummy_magic_25_0.VD3.t16 146.155
R7071 two_stage_opamp_dummy_magic_25_0.VD3.n40 two_stage_opamp_dummy_magic_25_0.VD3.t15 76.2576
R7072 two_stage_opamp_dummy_magic_25_0.VD3.n41 two_stage_opamp_dummy_magic_25_0.VD3.t12 76.2576
R7073 two_stage_opamp_dummy_magic_25_0.VD3.n34 two_stage_opamp_dummy_magic_25_0.VD3.n33 66.9922
R7074 two_stage_opamp_dummy_magic_25_0.VD3.n46 two_stage_opamp_dummy_magic_25_0.VD3.n35 66.9922
R7075 two_stage_opamp_dummy_magic_25_0.VD3.n45 two_stage_opamp_dummy_magic_25_0.VD3.n36 66.9922
R7076 two_stage_opamp_dummy_magic_25_0.VD3.n44 two_stage_opamp_dummy_magic_25_0.VD3.n37 66.9922
R7077 two_stage_opamp_dummy_magic_25_0.VD3.n39 two_stage_opamp_dummy_magic_25_0.VD3.n38 66.9922
R7078 two_stage_opamp_dummy_magic_25_0.VD3.n29 two_stage_opamp_dummy_magic_25_0.VD3.n28 66.0338
R7079 two_stage_opamp_dummy_magic_25_0.VD3.n27 two_stage_opamp_dummy_magic_25_0.VD3.n26 66.0338
R7080 two_stage_opamp_dummy_magic_25_0.VD3.n50 two_stage_opamp_dummy_magic_25_0.VD3.n49 66.0338
R7081 two_stage_opamp_dummy_magic_25_0.VD3.n31 two_stage_opamp_dummy_magic_25_0.VD3.n30 66.0338
R7082 two_stage_opamp_dummy_magic_25_0.VD3.n55 two_stage_opamp_dummy_magic_25_0.VD3.n54 66.0338
R7083 two_stage_opamp_dummy_magic_25_0.VD3.n59 two_stage_opamp_dummy_magic_25_0.VD3.n58 66.0338
R7084 two_stage_opamp_dummy_magic_25_0.VD3.n28 two_stage_opamp_dummy_magic_25_0.VD3.t32 11.2576
R7085 two_stage_opamp_dummy_magic_25_0.VD3.n28 two_stage_opamp_dummy_magic_25_0.VD3.t24 11.2576
R7086 two_stage_opamp_dummy_magic_25_0.VD3.n26 two_stage_opamp_dummy_magic_25_0.VD3.t26 11.2576
R7087 two_stage_opamp_dummy_magic_25_0.VD3.n26 two_stage_opamp_dummy_magic_25_0.VD3.t29 11.2576
R7088 two_stage_opamp_dummy_magic_25_0.VD3.n33 two_stage_opamp_dummy_magic_25_0.VD3.t21 11.2576
R7089 two_stage_opamp_dummy_magic_25_0.VD3.n33 two_stage_opamp_dummy_magic_25_0.VD3.t37 11.2576
R7090 two_stage_opamp_dummy_magic_25_0.VD3.n35 two_stage_opamp_dummy_magic_25_0.VD3.t35 11.2576
R7091 two_stage_opamp_dummy_magic_25_0.VD3.n35 two_stage_opamp_dummy_magic_25_0.VD3.t5 11.2576
R7092 two_stage_opamp_dummy_magic_25_0.VD3.n36 two_stage_opamp_dummy_magic_25_0.VD3.t3 11.2576
R7093 two_stage_opamp_dummy_magic_25_0.VD3.n36 two_stage_opamp_dummy_magic_25_0.VD3.t9 11.2576
R7094 two_stage_opamp_dummy_magic_25_0.VD3.n37 two_stage_opamp_dummy_magic_25_0.VD3.t19 11.2576
R7095 two_stage_opamp_dummy_magic_25_0.VD3.n37 two_stage_opamp_dummy_magic_25_0.VD3.t1 11.2576
R7096 two_stage_opamp_dummy_magic_25_0.VD3.n38 two_stage_opamp_dummy_magic_25_0.VD3.t7 11.2576
R7097 two_stage_opamp_dummy_magic_25_0.VD3.n38 two_stage_opamp_dummy_magic_25_0.VD3.t17 11.2576
R7098 two_stage_opamp_dummy_magic_25_0.VD3.n49 two_stage_opamp_dummy_magic_25_0.VD3.t28 11.2576
R7099 two_stage_opamp_dummy_magic_25_0.VD3.n49 two_stage_opamp_dummy_magic_25_0.VD3.t33 11.2576
R7100 two_stage_opamp_dummy_magic_25_0.VD3.n30 two_stage_opamp_dummy_magic_25_0.VD3.t27 11.2576
R7101 two_stage_opamp_dummy_magic_25_0.VD3.n30 two_stage_opamp_dummy_magic_25_0.VD3.t30 11.2576
R7102 two_stage_opamp_dummy_magic_25_0.VD3.n54 two_stage_opamp_dummy_magic_25_0.VD3.t23 11.2576
R7103 two_stage_opamp_dummy_magic_25_0.VD3.n54 two_stage_opamp_dummy_magic_25_0.VD3.t25 11.2576
R7104 two_stage_opamp_dummy_magic_25_0.VD3.t31 two_stage_opamp_dummy_magic_25_0.VD3.n59 11.2576
R7105 two_stage_opamp_dummy_magic_25_0.VD3.n59 two_stage_opamp_dummy_magic_25_0.VD3.t22 11.2576
R7106 two_stage_opamp_dummy_magic_25_0.VD3.n50 two_stage_opamp_dummy_magic_25_0.VD3.n25 5.91717
R7107 two_stage_opamp_dummy_magic_25_0.VD3.n29 two_stage_opamp_dummy_magic_25_0.VD3.n24 5.91717
R7108 two_stage_opamp_dummy_magic_25_0.VD3.n27 two_stage_opamp_dummy_magic_25_0.VD3.n24 5.29217
R7109 two_stage_opamp_dummy_magic_25_0.VD3.n31 two_stage_opamp_dummy_magic_25_0.VD3.n25 5.29217
R7110 two_stage_opamp_dummy_magic_25_0.VD3.n56 two_stage_opamp_dummy_magic_25_0.VD3.n55 5.29217
R7111 two_stage_opamp_dummy_magic_25_0.VD3.n58 two_stage_opamp_dummy_magic_25_0.VD3.n57 5.29217
R7112 two_stage_opamp_dummy_magic_25_0.VD3.n3 two_stage_opamp_dummy_magic_25_0.VD3.n5 0.740726
R7113 two_stage_opamp_dummy_magic_25_0.VD3.n4 two_stage_opamp_dummy_magic_25_0.VD3.n0 0.740726
R7114 two_stage_opamp_dummy_magic_25_0.VD3.n51 two_stage_opamp_dummy_magic_25_0.VD3.n4 0.0215479
R7115 two_stage_opamp_dummy_magic_25_0.VD3.n1 two_stage_opamp_dummy_magic_25_0.VD3.n2 0.740726
R7116 two_stage_opamp_dummy_magic_25_0.VD3.n53 two_stage_opamp_dummy_magic_25_0.VD3.n52 1.5005
R7117 two_stage_opamp_dummy_magic_25_0.VD3.n19 two_stage_opamp_dummy_magic_25_0.VD3.n17 0.740726
R7118 two_stage_opamp_dummy_magic_25_0.VD3.n15 two_stage_opamp_dummy_magic_25_0.VD3.n18 0.740726
R7119 two_stage_opamp_dummy_magic_25_0.VD3.n16 two_stage_opamp_dummy_magic_25_0.VD3.n13 0.740726
R7120 two_stage_opamp_dummy_magic_25_0.VD3.n45 two_stage_opamp_dummy_magic_25_0.VD3.n16 0.0215479
R7121 two_stage_opamp_dummy_magic_25_0.VD3.n11 two_stage_opamp_dummy_magic_25_0.VD3.n14 0.740726
R7122 two_stage_opamp_dummy_magic_25_0.VD3.n12 two_stage_opamp_dummy_magic_25_0.VD3.n9 0.740726
R7123 two_stage_opamp_dummy_magic_25_0.VD3.n6 two_stage_opamp_dummy_magic_25_0.VD3.n10 0.740726
R7124 two_stage_opamp_dummy_magic_25_0.VD3.n10 two_stage_opamp_dummy_magic_25_0.VD3.n34 0.0215479
R7125 two_stage_opamp_dummy_magic_25_0.VD3.n8 two_stage_opamp_dummy_magic_25_0.VD3.n7 0.740726
R7126 two_stage_opamp_dummy_magic_25_0.VD3.n48 two_stage_opamp_dummy_magic_25_0.VD3.n47 1.5005
R7127 two_stage_opamp_dummy_magic_25_0.VD3.n21 two_stage_opamp_dummy_magic_25_0.VD3.n20 0.740726
R7128 two_stage_opamp_dummy_magic_25_0.VD3.n23 two_stage_opamp_dummy_magic_25_0.VD3.n22 0.0749176
R7129 two_stage_opamp_dummy_magic_25_0.VD3.n40 two_stage_opamp_dummy_magic_25_0.VD3.n32 1.03383
R7130 two_stage_opamp_dummy_magic_25_0.VD3.n42 two_stage_opamp_dummy_magic_25_0.VD3.n41 1.03383
R7131 two_stage_opamp_dummy_magic_25_0.VD3.n22 two_stage_opamp_dummy_magic_25_0.VD3.n29 1.04479
R7132 two_stage_opamp_dummy_magic_25_0.VD3.n43 two_stage_opamp_dummy_magic_25_0.VD3.n42 1.02322
R7133 two_stage_opamp_dummy_magic_25_0.VD3.n23 two_stage_opamp_dummy_magic_25_0.VD3.n27 0.958833
R7134 two_stage_opamp_dummy_magic_25_0.VD3.n47 two_stage_opamp_dummy_magic_25_0.VD3.n32 0.958833
R7135 two_stage_opamp_dummy_magic_25_0.VD3.n51 two_stage_opamp_dummy_magic_25_0.VD3.n31 0.958833
R7136 two_stage_opamp_dummy_magic_25_0.VD3.n55 two_stage_opamp_dummy_magic_25_0.VD3.n53 0.958833
R7137 two_stage_opamp_dummy_magic_25_0.VD3.n5 two_stage_opamp_dummy_magic_25_0.VD3.n50 0.979881
R7138 two_stage_opamp_dummy_magic_25_0.VD3.n58 two_stage_opamp_dummy_magic_25_0.VD3.n20 0.958833
R7139 two_stage_opamp_dummy_magic_25_0.VD3.n3 two_stage_opamp_dummy_magic_25_0.VD3.n48 0.786958
R7140 two_stage_opamp_dummy_magic_25_0.VD3.n57 two_stage_opamp_dummy_magic_25_0.VD3.n56 0.6255
R7141 two_stage_opamp_dummy_magic_25_0.VD3.n56 two_stage_opamp_dummy_magic_25_0.VD3.n25 0.6255
R7142 two_stage_opamp_dummy_magic_25_0.VD3.n57 two_stage_opamp_dummy_magic_25_0.VD3.n24 0.6255
R7143 two_stage_opamp_dummy_magic_25_0.VD3.n22 two_stage_opamp_dummy_magic_25_0.VD3.n21 0.37999
R7144 two_stage_opamp_dummy_magic_25_0.VD3.n17 two_stage_opamp_dummy_magic_25_0.VD3.n43 0.427973
R7145 two_stage_opamp_dummy_magic_25_0.VD3.n20 two_stage_opamp_dummy_magic_25_0.VD3.n23 0.0838333
R7146 two_stage_opamp_dummy_magic_25_0.VD3.n43 two_stage_opamp_dummy_magic_25_0.VD3.n39 0.0587394
R7147 two_stage_opamp_dummy_magic_25_0.VD3.n47 two_stage_opamp_dummy_magic_25_0.VD3.n8 0.0632146
R7148 two_stage_opamp_dummy_magic_25_0.VD3.n8 two_stage_opamp_dummy_magic_25_0.VD3.n34 0.0632146
R7149 two_stage_opamp_dummy_magic_25_0.VD3.n12 two_stage_opamp_dummy_magic_25_0.VD3.n10 0.0842626
R7150 two_stage_opamp_dummy_magic_25_0.VD3.n12 two_stage_opamp_dummy_magic_25_0.VD3.n46 0.0215479
R7151 two_stage_opamp_dummy_magic_25_0.VD3.n46 two_stage_opamp_dummy_magic_25_0.VD3.n14 0.0632146
R7152 two_stage_opamp_dummy_magic_25_0.VD3.n45 two_stage_opamp_dummy_magic_25_0.VD3.n14 0.0632146
R7153 two_stage_opamp_dummy_magic_25_0.VD3.n16 two_stage_opamp_dummy_magic_25_0.VD3.n18 0.0842626
R7154 two_stage_opamp_dummy_magic_25_0.VD3.n44 two_stage_opamp_dummy_magic_25_0.VD3.n18 0.0215479
R7155 two_stage_opamp_dummy_magic_25_0.VD3.n44 two_stage_opamp_dummy_magic_25_0.VD3.n19 0.0632146
R7156 two_stage_opamp_dummy_magic_25_0.VD3.n19 two_stage_opamp_dummy_magic_25_0.VD3.n39 0.0632146
R7157 two_stage_opamp_dummy_magic_25_0.VD3.n53 two_stage_opamp_dummy_magic_25_0.VD3.n2 0.0632146
R7158 two_stage_opamp_dummy_magic_25_0.VD3.n51 two_stage_opamp_dummy_magic_25_0.VD3.n2 0.0632146
R7159 two_stage_opamp_dummy_magic_25_0.VD3.n4 two_stage_opamp_dummy_magic_25_0.VD3.n5 0.0842626
R7160 two_stage_opamp_dummy_magic_25_0.VD3.n52 two_stage_opamp_dummy_magic_25_0.VD3.n21 0.146548
R7161 two_stage_opamp_dummy_magic_25_0.VD3.n15 two_stage_opamp_dummy_magic_25_0.VD3.n17 0.0838333
R7162 two_stage_opamp_dummy_magic_25_0.VD3.n13 two_stage_opamp_dummy_magic_25_0.VD3.n15 0.0838333
R7163 two_stage_opamp_dummy_magic_25_0.VD3.n11 two_stage_opamp_dummy_magic_25_0.VD3.n13 0.0838333
R7164 two_stage_opamp_dummy_magic_25_0.VD3.n9 two_stage_opamp_dummy_magic_25_0.VD3.n11 0.0838333
R7165 two_stage_opamp_dummy_magic_25_0.VD3.n6 two_stage_opamp_dummy_magic_25_0.VD3.n9 0.0838333
R7166 two_stage_opamp_dummy_magic_25_0.VD3.n7 two_stage_opamp_dummy_magic_25_0.VD3.n6 0.0838333
R7167 two_stage_opamp_dummy_magic_25_0.VD3.n48 two_stage_opamp_dummy_magic_25_0.VD3.n7 0.0838333
R7168 two_stage_opamp_dummy_magic_25_0.VD3.n0 two_stage_opamp_dummy_magic_25_0.VD3.n3 0.0838333
R7169 two_stage_opamp_dummy_magic_25_0.VD3.n1 two_stage_opamp_dummy_magic_25_0.VD3.n0 0.0838333
R7170 two_stage_opamp_dummy_magic_25_0.VD3.n52 two_stage_opamp_dummy_magic_25_0.VD3.n1 0.0838333
R7171 VOUT+.n19 VOUT+.t1 110.191
R7172 VOUT+.n48 VOUT+.n47 34.9935
R7173 VOUT+.n46 VOUT+.n45 34.9935
R7174 VOUT+.n60 VOUT+.n59 34.9935
R7175 VOUT+.n56 VOUT+.n55 34.9935
R7176 VOUT+.n53 VOUT+.n52 34.9935
R7177 VOUT+.n50 VOUT+.n49 34.9935
R7178 VOUT+.n2 VOUT+.n1 9.73997
R7179 VOUT+.n6 VOUT+.n5 9.73997
R7180 VOUT+.n9 VOUT+.n8 9.73997
R7181 VOUT+.n7 VOUT+.n6 6.64633
R7182 VOUT+.n7 VOUT+.n2 6.64633
R7183 VOUT+.n47 VOUT+.t5 6.56717
R7184 VOUT+.n47 VOUT+.t15 6.56717
R7185 VOUT+.n45 VOUT+.t14 6.56717
R7186 VOUT+.n45 VOUT+.t18 6.56717
R7187 VOUT+.n59 VOUT+.t7 6.56717
R7188 VOUT+.n59 VOUT+.t6 6.56717
R7189 VOUT+.n55 VOUT+.t13 6.56717
R7190 VOUT+.n55 VOUT+.t2 6.56717
R7191 VOUT+.n52 VOUT+.t16 6.56717
R7192 VOUT+.n52 VOUT+.t8 6.56717
R7193 VOUT+.n49 VOUT+.t11 6.56717
R7194 VOUT+.n49 VOUT+.t17 6.56717
R7195 VOUT+.n58 VOUT+.n46 6.3755
R7196 VOUT+.n51 VOUT+.n48 6.3755
R7197 VOUT+.n9 VOUT+.n7 6.02133
R7198 VOUT+.n60 VOUT+.n58 5.813
R7199 VOUT+.n57 VOUT+.n56 5.813
R7200 VOUT+.n54 VOUT+.n53 5.813
R7201 VOUT+.n51 VOUT+.n50 5.813
R7202 VOUT+.n61 VOUT+.n37 5.063
R7203 VOUT+.n64 VOUT+.n44 5.063
R7204 VOUT+.n131 VOUT+.t52 4.8295
R7205 VOUT+.n132 VOUT+.t88 4.8295
R7206 VOUT+.n133 VOUT+.t123 4.8295
R7207 VOUT+.n134 VOUT+.t26 4.8295
R7208 VOUT+.n135 VOUT+.t68 4.8295
R7209 VOUT+.n136 VOUT+.t114 4.8295
R7210 VOUT+.n146 VOUT+.t144 4.8295
R7211 VOUT+.n148 VOUT+.t124 4.8295
R7212 VOUT+.n149 VOUT+.t33 4.8295
R7213 VOUT+.n151 VOUT+.t139 4.8295
R7214 VOUT+.n152 VOUT+.t27 4.8295
R7215 VOUT+.n154 VOUT+.t106 4.8295
R7216 VOUT+.n155 VOUT+.t132 4.8295
R7217 VOUT+.n157 VOUT+.t133 4.8295
R7218 VOUT+.n158 VOUT+.t21 4.8295
R7219 VOUT+.n160 VOUT+.t98 4.8295
R7220 VOUT+.n161 VOUT+.t126 4.8295
R7221 VOUT+.n163 VOUT+.t59 4.8295
R7222 VOUT+.n164 VOUT+.t90 4.8295
R7223 VOUT+.n166 VOUT+.t92 4.8295
R7224 VOUT+.n167 VOUT+.t125 4.8295
R7225 VOUT+.n169 VOUT+.t49 4.8295
R7226 VOUT+.n170 VOUT+.t82 4.8295
R7227 VOUT+.n172 VOUT+.t149 4.8295
R7228 VOUT+.n173 VOUT+.t39 4.8295
R7229 VOUT+.n175 VOUT+.t116 4.8295
R7230 VOUT+.n176 VOUT+.t143 4.8295
R7231 VOUT+.n98 VOUT+.t142 4.8295
R7232 VOUT+.n111 VOUT+.t109 4.8295
R7233 VOUT+.n113 VOUT+.t155 4.8295
R7234 VOUT+.n114 VOUT+.t47 4.8295
R7235 VOUT+.n116 VOUT+.t51 4.8295
R7236 VOUT+.n117 VOUT+.t84 4.8295
R7237 VOUT+.n119 VOUT+.t41 4.8295
R7238 VOUT+.n120 VOUT+.t48 4.8295
R7239 VOUT+.n122 VOUT+.t105 4.8295
R7240 VOUT+.n123 VOUT+.t131 4.8295
R7241 VOUT+.n125 VOUT+.t67 4.8295
R7242 VOUT+.n126 VOUT+.t101 4.8295
R7243 VOUT+.n128 VOUT+.t111 4.8295
R7244 VOUT+.n129 VOUT+.t137 4.8295
R7245 VOUT+.n178 VOUT+.t32 4.8295
R7246 VOUT+.n138 VOUT+.t91 4.8154
R7247 VOUT+.n110 VOUT+.t45 4.806
R7248 VOUT+.n109 VOUT+.t85 4.806
R7249 VOUT+.n108 VOUT+.t63 4.806
R7250 VOUT+.n107 VOUT+.t107 4.806
R7251 VOUT+.n106 VOUT+.t138 4.806
R7252 VOUT+.n105 VOUT+.t120 4.806
R7253 VOUT+.n104 VOUT+.t153 4.806
R7254 VOUT+.n103 VOUT+.t56 4.806
R7255 VOUT+.n102 VOUT+.t94 4.806
R7256 VOUT+.n101 VOUT+.t70 4.806
R7257 VOUT+.n100 VOUT+.t112 4.806
R7258 VOUT+.n131 VOUT+.t103 4.5005
R7259 VOUT+.n132 VOUT+.t136 4.5005
R7260 VOUT+.n133 VOUT+.t29 4.5005
R7261 VOUT+.n134 VOUT+.t151 4.5005
R7262 VOUT+.n135 VOUT+.t55 4.5005
R7263 VOUT+.n136 VOUT+.t72 4.5005
R7264 VOUT+.n137 VOUT+.t96 4.5005
R7265 VOUT+.n138 VOUT+.t57 4.5005
R7266 VOUT+.n139 VOUT+.t156 4.5005
R7267 VOUT+.n140 VOUT+.t121 4.5005
R7268 VOUT+.n141 VOUT+.t140 4.5005
R7269 VOUT+.n142 VOUT+.t108 4.5005
R7270 VOUT+.n143 VOUT+.t64 4.5005
R7271 VOUT+.n144 VOUT+.t89 4.5005
R7272 VOUT+.n145 VOUT+.t46 4.5005
R7273 VOUT+.n147 VOUT+.t40 4.5005
R7274 VOUT+.n146 VOUT+.t77 4.5005
R7275 VOUT+.n148 VOUT+.t83 4.5005
R7276 VOUT+.n150 VOUT+.t79 4.5005
R7277 VOUT+.n149 VOUT+.t117 4.5005
R7278 VOUT+.n151 VOUT+.t110 4.5005
R7279 VOUT+.n153 VOUT+.t80 4.5005
R7280 VOUT+.n152 VOUT+.t81 4.5005
R7281 VOUT+.n154 VOUT+.t66 4.5005
R7282 VOUT+.n156 VOUT+.t35 4.5005
R7283 VOUT+.n155 VOUT+.t37 4.5005
R7284 VOUT+.n157 VOUT+.t104 4.5005
R7285 VOUT+.n159 VOUT+.t75 4.5005
R7286 VOUT+.n158 VOUT+.t76 4.5005
R7287 VOUT+.n160 VOUT+.t61 4.5005
R7288 VOUT+.n162 VOUT+.t30 4.5005
R7289 VOUT+.n161 VOUT+.t31 4.5005
R7290 VOUT+.n163 VOUT+.t19 4.5005
R7291 VOUT+.n165 VOUT+.t134 4.5005
R7292 VOUT+.n164 VOUT+.t135 4.5005
R7293 VOUT+.n166 VOUT+.t58 4.5005
R7294 VOUT+.n168 VOUT+.t24 4.5005
R7295 VOUT+.n167 VOUT+.t25 4.5005
R7296 VOUT+.n169 VOUT+.t152 4.5005
R7297 VOUT+.n171 VOUT+.t127 4.5005
R7298 VOUT+.n170 VOUT+.t128 4.5005
R7299 VOUT+.n172 VOUT+.t118 4.5005
R7300 VOUT+.n174 VOUT+.t93 4.5005
R7301 VOUT+.n173 VOUT+.t95 4.5005
R7302 VOUT+.n175 VOUT+.t74 4.5005
R7303 VOUT+.n177 VOUT+.t50 4.5005
R7304 VOUT+.n176 VOUT+.t54 4.5005
R7305 VOUT+.n99 VOUT+.t38 4.5005
R7306 VOUT+.n98 VOUT+.t73 4.5005
R7307 VOUT+.n100 VOUT+.t69 4.5005
R7308 VOUT+.n101 VOUT+.t22 4.5005
R7309 VOUT+.n102 VOUT+.t53 4.5005
R7310 VOUT+.n103 VOUT+.t150 4.5005
R7311 VOUT+.n104 VOUT+.t119 4.5005
R7312 VOUT+.n105 VOUT+.t78 4.5005
R7313 VOUT+.n106 VOUT+.t102 4.5005
R7314 VOUT+.n107 VOUT+.t62 4.5005
R7315 VOUT+.n108 VOUT+.t20 4.5005
R7316 VOUT+.n109 VOUT+.t42 4.5005
R7317 VOUT+.n110 VOUT+.t148 4.5005
R7318 VOUT+.n112 VOUT+.t141 4.5005
R7319 VOUT+.n111 VOUT+.t28 4.5005
R7320 VOUT+.n113 VOUT+.t122 4.5005
R7321 VOUT+.n115 VOUT+.t99 4.5005
R7322 VOUT+.n114 VOUT+.t100 4.5005
R7323 VOUT+.n116 VOUT+.t154 4.5005
R7324 VOUT+.n118 VOUT+.t129 4.5005
R7325 VOUT+.n117 VOUT+.t130 4.5005
R7326 VOUT+.n119 VOUT+.t97 4.5005
R7327 VOUT+.n121 VOUT+.t60 4.5005
R7328 VOUT+.n120 VOUT+.t113 4.5005
R7329 VOUT+.n122 VOUT+.t65 4.5005
R7330 VOUT+.n124 VOUT+.t34 4.5005
R7331 VOUT+.n123 VOUT+.t36 4.5005
R7332 VOUT+.n125 VOUT+.t23 4.5005
R7333 VOUT+.n127 VOUT+.t146 4.5005
R7334 VOUT+.n126 VOUT+.t147 4.5005
R7335 VOUT+.n128 VOUT+.t71 4.5005
R7336 VOUT+.n130 VOUT+.t43 4.5005
R7337 VOUT+.n129 VOUT+.t44 4.5005
R7338 VOUT+.n180 VOUT+.t115 4.5005
R7339 VOUT+.n179 VOUT+.t86 4.5005
R7340 VOUT+.n178 VOUT+.t87 4.5005
R7341 VOUT+.n181 VOUT+.t145 4.5005
R7342 VOUT+.n61 VOUT+.n38 4.5005
R7343 VOUT+.n62 VOUT+.n41 4.5005
R7344 VOUT+.n63 VOUT+.n42 4.5005
R7345 VOUT+.n65 VOUT+.n64 4.5005
R7346 VOUT+.n88 VOUT+.n87 4.5005
R7347 VOUT+.n84 VOUT+.n81 4.5005
R7348 VOUT+.n88 VOUT+.n81 4.5005
R7349 VOUT+.n89 VOUT+.n33 4.5005
R7350 VOUT+.n89 VOUT+.n35 4.5005
R7351 VOUT+.n89 VOUT+.n88 4.5005
R7352 VOUT+.n186 VOUT+.n92 4.5005
R7353 VOUT+.n187 VOUT+.n186 4.5005
R7354 VOUT+.n187 VOUT+.n29 4.5005
R7355 VOUT+.n188 VOUT+.n28 4.5005
R7356 VOUT+.n188 VOUT+.n187 4.5005
R7357 VOUT+.n192 VOUT+.n191 4.5005
R7358 VOUT+.n191 VOUT+.n20 4.5005
R7359 VOUT+.n23 VOUT+.n20 4.5005
R7360 VOUT+.n194 VOUT+.n20 4.5005
R7361 VOUT+.n196 VOUT+.n20 4.5005
R7362 VOUT+.n195 VOUT+.n23 4.5005
R7363 VOUT+.n195 VOUT+.n194 4.5005
R7364 VOUT+.n196 VOUT+.n195 4.5005
R7365 VOUT+.n1 VOUT+.t12 3.42907
R7366 VOUT+.n1 VOUT+.t9 3.42907
R7367 VOUT+.n5 VOUT+.t4 3.42907
R7368 VOUT+.n5 VOUT+.t3 3.42907
R7369 VOUT+.n8 VOUT+.t0 3.42907
R7370 VOUT+.n8 VOUT+.t10 3.42907
R7371 VOUT+.n86 VOUT+.n34 2.26725
R7372 VOUT+.n82 VOUT+.n32 2.24601
R7373 VOUT+.n190 VOUT+.n189 2.24601
R7374 VOUT+.n25 VOUT+.n22 2.24601
R7375 VOUT+.n185 VOUT+.n184 2.24477
R7376 VOUT+.n31 VOUT+.n26 2.24477
R7377 VOUT+.n89 VOUT+.n34 2.24063
R7378 VOUT+.n188 VOUT+.n27 2.24063
R7379 VOUT+.n195 VOUT+.n24 2.24063
R7380 VOUT+.n81 VOUT+.n80 2.24063
R7381 VOUT+.n186 VOUT+.n90 2.24063
R7382 VOUT+.n91 VOUT+.n29 2.24063
R7383 VOUT+.n193 VOUT+.n192 2.24063
R7384 VOUT+.n192 VOUT+.n21 2.24063
R7385 VOUT+.n87 VOUT+.n85 2.23934
R7386 VOUT+.n87 VOUT+.n83 2.23934
R7387 VOUT+.n6 VOUT+.n4 1.62886
R7388 VOUT+.n10 VOUT+.n9 1.52133
R7389 VOUT+.n17 VOUT+.n2 1.52133
R7390 VOUT+.n79 VOUT+.n78 1.5005
R7391 VOUT+.n77 VOUT+.n36 1.5005
R7392 VOUT+.n76 VOUT+.n75 1.5005
R7393 VOUT+.n74 VOUT+.n39 1.5005
R7394 VOUT+.n73 VOUT+.n72 1.5005
R7395 VOUT+.n71 VOUT+.n40 1.5005
R7396 VOUT+.n70 VOUT+.n69 1.5005
R7397 VOUT+.n68 VOUT+.n43 1.5005
R7398 VOUT+.n18 VOUT+.n17 1.5005
R7399 VOUT+.n16 VOUT+.n0 1.5005
R7400 VOUT+.n15 VOUT+.n14 1.5005
R7401 VOUT+.n13 VOUT+.n3 1.5005
R7402 VOUT+.n12 VOUT+.n11 1.5005
R7403 VOUT+.n65 VOUT+.n60 1.313
R7404 VOUT+.n56 VOUT+.n42 1.313
R7405 VOUT+.n53 VOUT+.n41 1.313
R7406 VOUT+.n50 VOUT+.n38 1.313
R7407 VOUT+.n46 VOUT+.n44 1.313
R7408 VOUT+.n48 VOUT+.n37 1.313
R7409 VOUT+.n187 VOUT+.n30 1.1455
R7410 VOUT+.n96 VOUT+.n95 1.13717
R7411 VOUT+.n97 VOUT+.n93 1.13717
R7412 VOUT+.n183 VOUT+.n182 1.13717
R7413 VOUT+.n94 VOUT+.n31 1.13717
R7414 VOUT+.n95 VOUT+.n28 1.13717
R7415 VOUT+.n93 VOUT+.n92 1.13717
R7416 VOUT+.n184 VOUT+.n183 1.13717
R7417 VOUT+.n67 VOUT+.n44 0.715216
R7418 VOUT+.n66 VOUT+.n65 0.65675
R7419 VOUT+.n70 VOUT+.n42 0.65675
R7420 VOUT+.n72 VOUT+.n41 0.65675
R7421 VOUT+.n76 VOUT+.n38 0.65675
R7422 VOUT+.n78 VOUT+.n37 0.65675
R7423 VOUT+.n96 VOUT+.n30 0.585
R7424 VOUT+.n192 VOUT+.n188 0.5705
R7425 VOUT+.n68 VOUT+.n67 0.564601
R7426 VOUT+.n62 VOUT+.n61 0.563
R7427 VOUT+.n63 VOUT+.n62 0.563
R7428 VOUT+.n64 VOUT+.n63 0.563
R7429 VOUT+.n58 VOUT+.n57 0.563
R7430 VOUT+.n57 VOUT+.n54 0.563
R7431 VOUT+.n54 VOUT+.n51 0.563
R7432 VOUT+.n88 VOUT+.n79 0.495292
R7433 VOUT+.n19 VOUT+.n18 0.380708
R7434 VOUT+.n137 VOUT+.n136 0.3295
R7435 VOUT+.n138 VOUT+.n137 0.3295
R7436 VOUT+.n139 VOUT+.n138 0.3295
R7437 VOUT+.n140 VOUT+.n139 0.3295
R7438 VOUT+.n141 VOUT+.n140 0.3295
R7439 VOUT+.n142 VOUT+.n141 0.3295
R7440 VOUT+.n143 VOUT+.n142 0.3295
R7441 VOUT+.n144 VOUT+.n143 0.3295
R7442 VOUT+.n145 VOUT+.n144 0.3295
R7443 VOUT+.n147 VOUT+.n145 0.3295
R7444 VOUT+.n147 VOUT+.n146 0.3295
R7445 VOUT+.n150 VOUT+.n148 0.3295
R7446 VOUT+.n150 VOUT+.n149 0.3295
R7447 VOUT+.n153 VOUT+.n151 0.3295
R7448 VOUT+.n153 VOUT+.n152 0.3295
R7449 VOUT+.n156 VOUT+.n154 0.3295
R7450 VOUT+.n156 VOUT+.n155 0.3295
R7451 VOUT+.n159 VOUT+.n157 0.3295
R7452 VOUT+.n159 VOUT+.n158 0.3295
R7453 VOUT+.n162 VOUT+.n160 0.3295
R7454 VOUT+.n162 VOUT+.n161 0.3295
R7455 VOUT+.n165 VOUT+.n163 0.3295
R7456 VOUT+.n165 VOUT+.n164 0.3295
R7457 VOUT+.n168 VOUT+.n166 0.3295
R7458 VOUT+.n168 VOUT+.n167 0.3295
R7459 VOUT+.n171 VOUT+.n169 0.3295
R7460 VOUT+.n171 VOUT+.n170 0.3295
R7461 VOUT+.n174 VOUT+.n172 0.3295
R7462 VOUT+.n174 VOUT+.n173 0.3295
R7463 VOUT+.n177 VOUT+.n175 0.3295
R7464 VOUT+.n177 VOUT+.n176 0.3295
R7465 VOUT+.n99 VOUT+.n98 0.3295
R7466 VOUT+.n101 VOUT+.n100 0.3295
R7467 VOUT+.n102 VOUT+.n101 0.3295
R7468 VOUT+.n103 VOUT+.n102 0.3295
R7469 VOUT+.n104 VOUT+.n103 0.3295
R7470 VOUT+.n105 VOUT+.n104 0.3295
R7471 VOUT+.n106 VOUT+.n105 0.3295
R7472 VOUT+.n107 VOUT+.n106 0.3295
R7473 VOUT+.n108 VOUT+.n107 0.3295
R7474 VOUT+.n109 VOUT+.n108 0.3295
R7475 VOUT+.n110 VOUT+.n109 0.3295
R7476 VOUT+.n112 VOUT+.n110 0.3295
R7477 VOUT+.n112 VOUT+.n111 0.3295
R7478 VOUT+.n115 VOUT+.n113 0.3295
R7479 VOUT+.n115 VOUT+.n114 0.3295
R7480 VOUT+.n118 VOUT+.n116 0.3295
R7481 VOUT+.n118 VOUT+.n117 0.3295
R7482 VOUT+.n121 VOUT+.n119 0.3295
R7483 VOUT+.n121 VOUT+.n120 0.3295
R7484 VOUT+.n124 VOUT+.n122 0.3295
R7485 VOUT+.n124 VOUT+.n123 0.3295
R7486 VOUT+.n127 VOUT+.n125 0.3295
R7487 VOUT+.n127 VOUT+.n126 0.3295
R7488 VOUT+.n130 VOUT+.n128 0.3295
R7489 VOUT+.n130 VOUT+.n129 0.3295
R7490 VOUT+.n180 VOUT+.n179 0.3295
R7491 VOUT+.n179 VOUT+.n178 0.3295
R7492 VOUT+.n139 VOUT+.n135 0.3154
R7493 VOUT+.n12 VOUT+.n4 0.314966
R7494 VOUT+.n181 VOUT+.n180 0.313833
R7495 VOUT+.n143 VOUT+.n131 0.306
R7496 VOUT+.n142 VOUT+.n132 0.306
R7497 VOUT+.n141 VOUT+.n133 0.306
R7498 VOUT+.n140 VOUT+.n134 0.306
R7499 VOUT+.n150 VOUT+.n147 0.2825
R7500 VOUT+.n153 VOUT+.n150 0.2825
R7501 VOUT+.n156 VOUT+.n153 0.2825
R7502 VOUT+.n159 VOUT+.n156 0.2825
R7503 VOUT+.n162 VOUT+.n159 0.2825
R7504 VOUT+.n165 VOUT+.n162 0.2825
R7505 VOUT+.n168 VOUT+.n165 0.2825
R7506 VOUT+.n171 VOUT+.n168 0.2825
R7507 VOUT+.n174 VOUT+.n171 0.2825
R7508 VOUT+.n177 VOUT+.n174 0.2825
R7509 VOUT+.n112 VOUT+.n99 0.2825
R7510 VOUT+.n115 VOUT+.n112 0.2825
R7511 VOUT+.n118 VOUT+.n115 0.2825
R7512 VOUT+.n121 VOUT+.n118 0.2825
R7513 VOUT+.n124 VOUT+.n121 0.2825
R7514 VOUT+.n127 VOUT+.n124 0.2825
R7515 VOUT+.n130 VOUT+.n127 0.2825
R7516 VOUT+.n179 VOUT+.n130 0.2825
R7517 VOUT+.n179 VOUT+.n177 0.2825
R7518 VOUT+.n186 VOUT+.n89 0.2655
R7519 VOUT+ VOUT+.n196 0.15675
R7520 VOUT+.n182 VOUT+.n181 0.138367
R7521 VOUT+.n10 VOUT+.n4 0.0891864
R7522 VOUT+.n66 VOUT+.n43 0.0577917
R7523 VOUT+.n70 VOUT+.n43 0.0577917
R7524 VOUT+.n71 VOUT+.n70 0.0577917
R7525 VOUT+.n72 VOUT+.n71 0.0577917
R7526 VOUT+.n72 VOUT+.n39 0.0577917
R7527 VOUT+.n76 VOUT+.n39 0.0577917
R7528 VOUT+.n77 VOUT+.n76 0.0577917
R7529 VOUT+.n78 VOUT+.n77 0.0577917
R7530 VOUT+.n69 VOUT+.n68 0.0577917
R7531 VOUT+.n69 VOUT+.n40 0.0577917
R7532 VOUT+.n73 VOUT+.n40 0.0577917
R7533 VOUT+.n74 VOUT+.n73 0.0577917
R7534 VOUT+.n75 VOUT+.n74 0.0577917
R7535 VOUT+.n75 VOUT+.n36 0.0577917
R7536 VOUT+.n79 VOUT+.n36 0.0577917
R7537 VOUT+.n67 VOUT+.n66 0.054517
R7538 VOUT+.n194 VOUT+.n25 0.047375
R7539 VOUT+.n189 VOUT+.n23 0.047375
R7540 VOUT+.n187 VOUT+.n31 0.0421667
R7541 VOUT+.n88 VOUT+.n82 0.0421667
R7542 VOUT+.n11 VOUT+.n10 0.0421667
R7543 VOUT+.n11 VOUT+.n3 0.0421667
R7544 VOUT+.n15 VOUT+.n3 0.0421667
R7545 VOUT+.n16 VOUT+.n15 0.0421667
R7546 VOUT+.n17 VOUT+.n16 0.0421667
R7547 VOUT+.n13 VOUT+.n12 0.0421667
R7548 VOUT+.n14 VOUT+.n13 0.0421667
R7549 VOUT+.n14 VOUT+.n0 0.0421667
R7550 VOUT+.n18 VOUT+.n0 0.0421667
R7551 VOUT+ VOUT+.n19 0.0369583
R7552 VOUT+.n83 VOUT+.n82 0.0243161
R7553 VOUT+.n85 VOUT+.n33 0.0243161
R7554 VOUT+.n85 VOUT+.n84 0.0243161
R7555 VOUT+.n83 VOUT+.n35 0.0243161
R7556 VOUT+.n184 VOUT+.n27 0.0217373
R7557 VOUT+.n84 VOUT+.n34 0.0217373
R7558 VOUT+.n92 VOUT+.n27 0.0217373
R7559 VOUT+.n191 VOUT+.n24 0.0217373
R7560 VOUT+.n189 VOUT+.n24 0.0217373
R7561 VOUT+.n90 VOUT+.n31 0.0217373
R7562 VOUT+.n92 VOUT+.n91 0.0217373
R7563 VOUT+.n80 VOUT+.n33 0.0217373
R7564 VOUT+.n80 VOUT+.n35 0.0217373
R7565 VOUT+.n90 VOUT+.n28 0.0217373
R7566 VOUT+.n91 VOUT+.n28 0.0217373
R7567 VOUT+.n196 VOUT+.n21 0.0217373
R7568 VOUT+.n194 VOUT+.n193 0.0217373
R7569 VOUT+.n193 VOUT+.n23 0.0217373
R7570 VOUT+.n25 VOUT+.n21 0.0217373
R7571 VOUT+.n97 VOUT+.n96 0.0161667
R7572 VOUT+.n182 VOUT+.n97 0.0161667
R7573 VOUT+.n95 VOUT+.n94 0.0161667
R7574 VOUT+.n95 VOUT+.n93 0.0161667
R7575 VOUT+.n183 VOUT+.n93 0.0161667
R7576 VOUT+.n185 VOUT+.n29 0.0134654
R7577 VOUT+.n188 VOUT+.n26 0.0134654
R7578 VOUT+.n186 VOUT+.n185 0.0134654
R7579 VOUT+.n29 VOUT+.n26 0.0134654
R7580 VOUT+.n86 VOUT+.n81 0.0109778
R7581 VOUT+.n89 VOUT+.n32 0.0109778
R7582 VOUT+.n190 VOUT+.n20 0.0109778
R7583 VOUT+.n195 VOUT+.n22 0.0109778
R7584 VOUT+.n87 VOUT+.n86 0.0109778
R7585 VOUT+.n81 VOUT+.n32 0.0109778
R7586 VOUT+.n192 VOUT+.n190 0.0109778
R7587 VOUT+.n22 VOUT+.n20 0.0109778
R7588 VOUT+.n94 VOUT+.n30 0.00872683
R7589 two_stage_opamp_dummy_magic_25_0.cap_res_Y two_stage_opamp_dummy_magic_25_0.cap_res_Y.t0 49.4263
R7590 two_stage_opamp_dummy_magic_25_0.cap_res_Y two_stage_opamp_dummy_magic_25_0.cap_res_Y.t69 1.481
R7591 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t80 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t13 0.1603
R7592 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t124 0.1603
R7593 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t33 0.1603
R7594 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t130 0.1603
R7595 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t18 0.1603
R7596 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t25 0.1603
R7597 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t51 0.1603
R7598 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t136 0.1603
R7599 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t24 0.1603
R7600 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t31 0.1603
R7601 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t59 0.1603
R7602 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t67 0.1603
R7603 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t98 0.1603
R7604 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t32 0.1603
R7605 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t65 0.1603
R7606 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t75 0.1603
R7607 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t108 0.1603
R7608 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t118 0.1603
R7609 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t8 0.1603
R7610 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t14 0.1603
R7611 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t41 0.1603
R7612 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t125 0.1603
R7613 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t12 0.1603
R7614 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t20 0.1603
R7615 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t46 0.1603
R7616 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t56 0.1603
R7617 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t90 0.1603
R7618 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t26 0.1603
R7619 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t52 0.1603
R7620 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t109 0.1603
R7621 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t116 0.1603
R7622 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t73 0.1603
R7623 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t106 0.1603
R7624 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t110 0.1603
R7625 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t2 0.1603
R7626 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t48 0.1603
R7627 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t45 0.1603
R7628 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t87 0.1603
R7629 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t63 0.1603
R7630 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t101 0.1603
R7631 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t4 0.1603
R7632 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t37 0.1603
R7633 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t19 0.1603
R7634 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t50 0.1603
R7635 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t94 0.1603
R7636 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t72 0.1603
R7637 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t112 0.1603
R7638 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t15 0.1603
R7639 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t111 0.1603
R7640 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t105 0.1603
R7641 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t54 0.1603
R7642 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t43 0.1603
R7643 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t85 0.1603
R7644 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t66 0.1603
R7645 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t89 0.1603
R7646 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t102 0.1603
R7647 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t131 0.1603
R7648 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t6 0.1603
R7649 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t34 0.1603
R7650 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t128 0.1603
R7651 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t49 0.1603
R7652 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t21 0.1603
R7653 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n14 0.159278
R7654 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n15 0.159278
R7655 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n16 0.159278
R7656 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n17 0.159278
R7657 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n18 0.159278
R7658 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n19 0.159278
R7659 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n20 0.159278
R7660 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n21 0.159278
R7661 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n22 0.159278
R7662 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n23 0.159278
R7663 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n24 0.159278
R7664 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n25 0.159278
R7665 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n26 0.159278
R7666 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n27 0.159278
R7667 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n28 0.159278
R7668 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n29 0.159278
R7669 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n30 0.159278
R7670 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n31 0.159278
R7671 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n32 0.159278
R7672 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t80 0.1368
R7673 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t40 0.1368
R7674 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t74 0.1368
R7675 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t76 0.1368
R7676 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t47 0.1368
R7677 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t120 0.1368
R7678 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t91 0.1368
R7679 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t81 0.1368
R7680 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t53 0.1368
R7681 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t126 0.1368
R7682 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t96 0.1368
R7683 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t22 0.1368
R7684 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t138 0.1368
R7685 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t132 0.1368
R7686 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t99 0.1368
R7687 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t29 0.1368
R7688 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t5 0.1368
R7689 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t62 0.1368
R7690 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t39 0.1368
R7691 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t103 0.1368
R7692 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t83 0.1368
R7693 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t70 0.1368
R7694 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t42 0.1368
R7695 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t113 0.1368
R7696 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t86 0.1368
R7697 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t10 0.1368
R7698 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t134 0.1368
R7699 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t121 0.1368
R7700 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t92 0.1368
R7701 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t44 0.1368
R7702 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t60 0.1368
R7703 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t27 0.1368
R7704 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t3 0.1368
R7705 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t57 0.1368
R7706 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t35 0.1368
R7707 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t129 0.1368
R7708 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t84 0.1368
R7709 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n33 0.1368
R7710 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t68 0.1368
R7711 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t61 0.1368
R7712 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t88 0.114322
R7713 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n4 0.1133
R7714 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n5 0.1133
R7715 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n6 0.1133
R7716 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n7 0.1133
R7717 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n8 0.1133
R7718 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n9 0.1133
R7719 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n10 0.1133
R7720 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n11 0.1133
R7721 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n12 0.1133
R7722 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n13 0.1133
R7723 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n0 0.1133
R7724 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n1 0.1133
R7725 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n2 0.1133
R7726 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n3 0.1133
R7727 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n34 0.1133
R7728 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t135 0.00152174
R7729 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t104 0.00152174
R7730 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t7 0.00152174
R7731 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t38 0.00152174
R7732 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t79 0.00152174
R7733 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t55 0.00152174
R7734 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t95 0.00152174
R7735 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t137 0.00152174
R7736 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t115 0.00152174
R7737 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t9 0.00152174
R7738 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t119 0.00152174
R7739 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t16 0.00152174
R7740 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t58 0.00152174
R7741 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t28 0.00152174
R7742 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t97 0.00152174
R7743 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t123 0.00152174
R7744 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t11 0.00152174
R7745 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t114 0.00152174
R7746 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t71 0.00152174
R7747 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t107 0.00152174
R7748 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t64 0.00152174
R7749 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t30 0.00152174
R7750 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t133 0.00152174
R7751 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t23 0.00152174
R7752 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t127 0.00152174
R7753 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t82 0.00152174
R7754 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t122 0.00152174
R7755 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t77 0.00152174
R7756 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t78 0.00152174
R7757 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t117 0.00152174
R7758 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t93 0.00152174
R7759 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t100 0.00152174
R7760 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t1 0.00152174
R7761 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t36 0.00152174
R7762 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t17 0.00152174
R7763 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n35 0.00152174
R7764 two_stage_opamp_dummy_magic_25_0.Vb2.n7 two_stage_opamp_dummy_magic_25_0.Vb2.t22 746.673
R7765 two_stage_opamp_dummy_magic_25_0.Vb2.n29 two_stage_opamp_dummy_magic_25_0.Vb2.t3 721.625
R7766 two_stage_opamp_dummy_magic_25_0.Vb2.n21 two_stage_opamp_dummy_magic_25_0.Vb2.t27 611.739
R7767 two_stage_opamp_dummy_magic_25_0.Vb2.n17 two_stage_opamp_dummy_magic_25_0.Vb2.t20 611.739
R7768 two_stage_opamp_dummy_magic_25_0.Vb2.n12 two_stage_opamp_dummy_magic_25_0.Vb2.t15 611.739
R7769 two_stage_opamp_dummy_magic_25_0.Vb2.n8 two_stage_opamp_dummy_magic_25_0.Vb2.t12 611.739
R7770 two_stage_opamp_dummy_magic_25_0.Vb2.n28 two_stage_opamp_dummy_magic_25_0.Vb2.t31 563.451
R7771 two_stage_opamp_dummy_magic_25_0.Vb2.n21 two_stage_opamp_dummy_magic_25_0.Vb2.t24 421.75
R7772 two_stage_opamp_dummy_magic_25_0.Vb2.n22 two_stage_opamp_dummy_magic_25_0.Vb2.t18 421.75
R7773 two_stage_opamp_dummy_magic_25_0.Vb2.n23 two_stage_opamp_dummy_magic_25_0.Vb2.t14 421.75
R7774 two_stage_opamp_dummy_magic_25_0.Vb2.n24 two_stage_opamp_dummy_magic_25_0.Vb2.t30 421.75
R7775 two_stage_opamp_dummy_magic_25_0.Vb2.n17 two_stage_opamp_dummy_magic_25_0.Vb2.t16 421.75
R7776 two_stage_opamp_dummy_magic_25_0.Vb2.n18 two_stage_opamp_dummy_magic_25_0.Vb2.t21 421.75
R7777 two_stage_opamp_dummy_magic_25_0.Vb2.n19 two_stage_opamp_dummy_magic_25_0.Vb2.t26 421.75
R7778 two_stage_opamp_dummy_magic_25_0.Vb2.n20 two_stage_opamp_dummy_magic_25_0.Vb2.t28 421.75
R7779 two_stage_opamp_dummy_magic_25_0.Vb2.n12 two_stage_opamp_dummy_magic_25_0.Vb2.t11 421.75
R7780 two_stage_opamp_dummy_magic_25_0.Vb2.n13 two_stage_opamp_dummy_magic_25_0.Vb2.t13 421.75
R7781 two_stage_opamp_dummy_magic_25_0.Vb2.n14 two_stage_opamp_dummy_magic_25_0.Vb2.t32 421.75
R7782 two_stage_opamp_dummy_magic_25_0.Vb2.n15 two_stage_opamp_dummy_magic_25_0.Vb2.t29 421.75
R7783 two_stage_opamp_dummy_magic_25_0.Vb2.n8 two_stage_opamp_dummy_magic_25_0.Vb2.t17 421.75
R7784 two_stage_opamp_dummy_magic_25_0.Vb2.n9 two_stage_opamp_dummy_magic_25_0.Vb2.t23 421.75
R7785 two_stage_opamp_dummy_magic_25_0.Vb2.n10 two_stage_opamp_dummy_magic_25_0.Vb2.t19 421.75
R7786 two_stage_opamp_dummy_magic_25_0.Vb2.n11 two_stage_opamp_dummy_magic_25_0.Vb2.t25 421.75
R7787 two_stage_opamp_dummy_magic_25_0.Vb2.n26 two_stage_opamp_dummy_magic_25_0.Vb2.n16 313.776
R7788 two_stage_opamp_dummy_magic_25_0.Vb2.n26 two_stage_opamp_dummy_magic_25_0.Vb2.n25 313.212
R7789 two_stage_opamp_dummy_magic_25_0.Vb2.n22 two_stage_opamp_dummy_magic_25_0.Vb2.n21 167.094
R7790 two_stage_opamp_dummy_magic_25_0.Vb2.n23 two_stage_opamp_dummy_magic_25_0.Vb2.n22 167.094
R7791 two_stage_opamp_dummy_magic_25_0.Vb2.n24 two_stage_opamp_dummy_magic_25_0.Vb2.n23 167.094
R7792 two_stage_opamp_dummy_magic_25_0.Vb2.n18 two_stage_opamp_dummy_magic_25_0.Vb2.n17 167.094
R7793 two_stage_opamp_dummy_magic_25_0.Vb2.n19 two_stage_opamp_dummy_magic_25_0.Vb2.n18 167.094
R7794 two_stage_opamp_dummy_magic_25_0.Vb2.n20 two_stage_opamp_dummy_magic_25_0.Vb2.n19 167.094
R7795 two_stage_opamp_dummy_magic_25_0.Vb2.n13 two_stage_opamp_dummy_magic_25_0.Vb2.n12 167.094
R7796 two_stage_opamp_dummy_magic_25_0.Vb2.n14 two_stage_opamp_dummy_magic_25_0.Vb2.n13 167.094
R7797 two_stage_opamp_dummy_magic_25_0.Vb2.n15 two_stage_opamp_dummy_magic_25_0.Vb2.n14 167.094
R7798 two_stage_opamp_dummy_magic_25_0.Vb2.n9 two_stage_opamp_dummy_magic_25_0.Vb2.n8 167.094
R7799 two_stage_opamp_dummy_magic_25_0.Vb2.n10 two_stage_opamp_dummy_magic_25_0.Vb2.n9 167.094
R7800 two_stage_opamp_dummy_magic_25_0.Vb2.n11 two_stage_opamp_dummy_magic_25_0.Vb2.n10 167.094
R7801 two_stage_opamp_dummy_magic_25_0.Vb2.n2 two_stage_opamp_dummy_magic_25_0.Vb2.n0 140.546
R7802 two_stage_opamp_dummy_magic_25_0.Vb2.n6 two_stage_opamp_dummy_magic_25_0.Vb2.n5 139.297
R7803 two_stage_opamp_dummy_magic_25_0.Vb2.n4 two_stage_opamp_dummy_magic_25_0.Vb2.n3 139.297
R7804 two_stage_opamp_dummy_magic_25_0.Vb2.n2 two_stage_opamp_dummy_magic_25_0.Vb2.n1 139.297
R7805 two_stage_opamp_dummy_magic_25_0.Vb2.n7 two_stage_opamp_dummy_magic_25_0.Vb2.n6 82.6036
R7806 two_stage_opamp_dummy_magic_25_0.Vb2.n30 two_stage_opamp_dummy_magic_25_0.Vb2.n29 67.013
R7807 two_stage_opamp_dummy_magic_25_0.Vb2.n25 two_stage_opamp_dummy_magic_25_0.Vb2.n24 35.3472
R7808 two_stage_opamp_dummy_magic_25_0.Vb2.n25 two_stage_opamp_dummy_magic_25_0.Vb2.n20 35.3472
R7809 two_stage_opamp_dummy_magic_25_0.Vb2.n16 two_stage_opamp_dummy_magic_25_0.Vb2.n15 35.3472
R7810 two_stage_opamp_dummy_magic_25_0.Vb2.n16 two_stage_opamp_dummy_magic_25_0.Vb2.n11 35.3472
R7811 two_stage_opamp_dummy_magic_25_0.Vb2.n5 two_stage_opamp_dummy_magic_25_0.Vb2.t6 24.0005
R7812 two_stage_opamp_dummy_magic_25_0.Vb2.n5 two_stage_opamp_dummy_magic_25_0.Vb2.t2 24.0005
R7813 two_stage_opamp_dummy_magic_25_0.Vb2.n3 two_stage_opamp_dummy_magic_25_0.Vb2.t10 24.0005
R7814 two_stage_opamp_dummy_magic_25_0.Vb2.n3 two_stage_opamp_dummy_magic_25_0.Vb2.t9 24.0005
R7815 two_stage_opamp_dummy_magic_25_0.Vb2.n1 two_stage_opamp_dummy_magic_25_0.Vb2.t1 24.0005
R7816 two_stage_opamp_dummy_magic_25_0.Vb2.n1 two_stage_opamp_dummy_magic_25_0.Vb2.t0 24.0005
R7817 two_stage_opamp_dummy_magic_25_0.Vb2.n0 two_stage_opamp_dummy_magic_25_0.Vb2.t8 24.0005
R7818 two_stage_opamp_dummy_magic_25_0.Vb2.n0 two_stage_opamp_dummy_magic_25_0.Vb2.t5 24.0005
R7819 two_stage_opamp_dummy_magic_25_0.Vb2.n27 two_stage_opamp_dummy_magic_25_0.Vb2.n26 14.5005
R7820 two_stage_opamp_dummy_magic_25_0.Vb2.t4 two_stage_opamp_dummy_magic_25_0.Vb2.n30 11.2576
R7821 two_stage_opamp_dummy_magic_25_0.Vb2.n30 two_stage_opamp_dummy_magic_25_0.Vb2.t7 11.2576
R7822 two_stage_opamp_dummy_magic_25_0.Vb2.n29 two_stage_opamp_dummy_magic_25_0.Vb2.n28 7.35988
R7823 two_stage_opamp_dummy_magic_25_0.Vb2.n4 two_stage_opamp_dummy_magic_25_0.Vb2.n2 5.8755
R7824 two_stage_opamp_dummy_magic_25_0.Vb2.n27 two_stage_opamp_dummy_magic_25_0.Vb2.n7 4.55362
R7825 two_stage_opamp_dummy_magic_25_0.Vb2.n6 two_stage_opamp_dummy_magic_25_0.Vb2.n4 1.2505
R7826 two_stage_opamp_dummy_magic_25_0.Vb2.n28 two_stage_opamp_dummy_magic_25_0.Vb2.n27 1.14112
R7827 two_stage_opamp_dummy_magic_25_0.X.n51 two_stage_opamp_dummy_magic_25_0.X.t51 1172.87
R7828 two_stage_opamp_dummy_magic_25_0.X.n47 two_stage_opamp_dummy_magic_25_0.X.t46 1172.87
R7829 two_stage_opamp_dummy_magic_25_0.X.n51 two_stage_opamp_dummy_magic_25_0.X.t38 996.134
R7830 two_stage_opamp_dummy_magic_25_0.X.n52 two_stage_opamp_dummy_magic_25_0.X.t26 996.134
R7831 two_stage_opamp_dummy_magic_25_0.X.n53 two_stage_opamp_dummy_magic_25_0.X.t37 996.134
R7832 two_stage_opamp_dummy_magic_25_0.X.n54 two_stage_opamp_dummy_magic_25_0.X.t25 996.134
R7833 two_stage_opamp_dummy_magic_25_0.X.n50 two_stage_opamp_dummy_magic_25_0.X.t41 996.134
R7834 two_stage_opamp_dummy_magic_25_0.X.n49 two_stage_opamp_dummy_magic_25_0.X.t29 996.134
R7835 two_stage_opamp_dummy_magic_25_0.X.n48 two_stage_opamp_dummy_magic_25_0.X.t44 996.134
R7836 two_stage_opamp_dummy_magic_25_0.X.n47 two_stage_opamp_dummy_magic_25_0.X.t31 996.134
R7837 two_stage_opamp_dummy_magic_25_0.X.n18 two_stage_opamp_dummy_magic_25_0.X.t47 690.867
R7838 two_stage_opamp_dummy_magic_25_0.X.n17 two_stage_opamp_dummy_magic_25_0.X.t43 690.867
R7839 two_stage_opamp_dummy_magic_25_0.X.n27 two_stage_opamp_dummy_magic_25_0.X.t48 530.201
R7840 two_stage_opamp_dummy_magic_25_0.X.n26 two_stage_opamp_dummy_magic_25_0.X.t45 530.201
R7841 two_stage_opamp_dummy_magic_25_0.X.n24 two_stage_opamp_dummy_magic_25_0.X.t40 514.134
R7842 two_stage_opamp_dummy_magic_25_0.X.n23 two_stage_opamp_dummy_magic_25_0.X.t54 514.134
R7843 two_stage_opamp_dummy_magic_25_0.X.n22 two_stage_opamp_dummy_magic_25_0.X.t36 514.134
R7844 two_stage_opamp_dummy_magic_25_0.X.n21 two_stage_opamp_dummy_magic_25_0.X.t49 514.134
R7845 two_stage_opamp_dummy_magic_25_0.X.n20 two_stage_opamp_dummy_magic_25_0.X.t32 514.134
R7846 two_stage_opamp_dummy_magic_25_0.X.n19 two_stage_opamp_dummy_magic_25_0.X.t50 514.134
R7847 two_stage_opamp_dummy_magic_25_0.X.n18 two_stage_opamp_dummy_magic_25_0.X.t33 514.134
R7848 two_stage_opamp_dummy_magic_25_0.X.n17 two_stage_opamp_dummy_magic_25_0.X.t28 514.134
R7849 two_stage_opamp_dummy_magic_25_0.X.n27 two_stage_opamp_dummy_magic_25_0.X.t35 353.467
R7850 two_stage_opamp_dummy_magic_25_0.X.n28 two_stage_opamp_dummy_magic_25_0.X.t53 353.467
R7851 two_stage_opamp_dummy_magic_25_0.X.n29 two_stage_opamp_dummy_magic_25_0.X.t34 353.467
R7852 two_stage_opamp_dummy_magic_25_0.X.n30 two_stage_opamp_dummy_magic_25_0.X.t52 353.467
R7853 two_stage_opamp_dummy_magic_25_0.X.n31 two_stage_opamp_dummy_magic_25_0.X.t39 353.467
R7854 two_stage_opamp_dummy_magic_25_0.X.n32 two_stage_opamp_dummy_magic_25_0.X.t27 353.467
R7855 two_stage_opamp_dummy_magic_25_0.X.n33 two_stage_opamp_dummy_magic_25_0.X.t42 353.467
R7856 two_stage_opamp_dummy_magic_25_0.X.n26 two_stage_opamp_dummy_magic_25_0.X.t30 353.467
R7857 two_stage_opamp_dummy_magic_25_0.X.n50 two_stage_opamp_dummy_magic_25_0.X.n49 176.733
R7858 two_stage_opamp_dummy_magic_25_0.X.n49 two_stage_opamp_dummy_magic_25_0.X.n48 176.733
R7859 two_stage_opamp_dummy_magic_25_0.X.n48 two_stage_opamp_dummy_magic_25_0.X.n47 176.733
R7860 two_stage_opamp_dummy_magic_25_0.X.n52 two_stage_opamp_dummy_magic_25_0.X.n51 176.733
R7861 two_stage_opamp_dummy_magic_25_0.X.n53 two_stage_opamp_dummy_magic_25_0.X.n52 176.733
R7862 two_stage_opamp_dummy_magic_25_0.X.n54 two_stage_opamp_dummy_magic_25_0.X.n53 176.733
R7863 two_stage_opamp_dummy_magic_25_0.X.n28 two_stage_opamp_dummy_magic_25_0.X.n27 176.733
R7864 two_stage_opamp_dummy_magic_25_0.X.n29 two_stage_opamp_dummy_magic_25_0.X.n28 176.733
R7865 two_stage_opamp_dummy_magic_25_0.X.n30 two_stage_opamp_dummy_magic_25_0.X.n29 176.733
R7866 two_stage_opamp_dummy_magic_25_0.X.n31 two_stage_opamp_dummy_magic_25_0.X.n30 176.733
R7867 two_stage_opamp_dummy_magic_25_0.X.n32 two_stage_opamp_dummy_magic_25_0.X.n31 176.733
R7868 two_stage_opamp_dummy_magic_25_0.X.n33 two_stage_opamp_dummy_magic_25_0.X.n32 176.733
R7869 two_stage_opamp_dummy_magic_25_0.X.n19 two_stage_opamp_dummy_magic_25_0.X.n18 176.733
R7870 two_stage_opamp_dummy_magic_25_0.X.n20 two_stage_opamp_dummy_magic_25_0.X.n19 176.733
R7871 two_stage_opamp_dummy_magic_25_0.X.n21 two_stage_opamp_dummy_magic_25_0.X.n20 176.733
R7872 two_stage_opamp_dummy_magic_25_0.X.n22 two_stage_opamp_dummy_magic_25_0.X.n21 176.733
R7873 two_stage_opamp_dummy_magic_25_0.X.n23 two_stage_opamp_dummy_magic_25_0.X.n22 176.733
R7874 two_stage_opamp_dummy_magic_25_0.X.n24 two_stage_opamp_dummy_magic_25_0.X.n23 176.733
R7875 two_stage_opamp_dummy_magic_25_0.X.n35 two_stage_opamp_dummy_magic_25_0.X.n34 165.472
R7876 two_stage_opamp_dummy_magic_25_0.X.n35 two_stage_opamp_dummy_magic_25_0.X.n25 165.472
R7877 two_stage_opamp_dummy_magic_25_0.X.n57 two_stage_opamp_dummy_magic_25_0.X.n56 152
R7878 two_stage_opamp_dummy_magic_25_0.X.n58 two_stage_opamp_dummy_magic_25_0.X.n57 131.571
R7879 two_stage_opamp_dummy_magic_25_0.X.n57 two_stage_opamp_dummy_magic_25_0.X.n55 124.517
R7880 two_stage_opamp_dummy_magic_25_0.X.n125 two_stage_opamp_dummy_magic_25_0.X.n35 74.5362
R7881 two_stage_opamp_dummy_magic_25_0.X.n79 two_stage_opamp_dummy_magic_25_0.X.n78 66.0338
R7882 two_stage_opamp_dummy_magic_25_0.X.n77 two_stage_opamp_dummy_magic_25_0.X.n76 66.0338
R7883 two_stage_opamp_dummy_magic_25_0.X.n89 two_stage_opamp_dummy_magic_25_0.X.n88 66.0338
R7884 two_stage_opamp_dummy_magic_25_0.X.n85 two_stage_opamp_dummy_magic_25_0.X.n84 66.0338
R7885 two_stage_opamp_dummy_magic_25_0.X.n82 two_stage_opamp_dummy_magic_25_0.X.n81 66.0338
R7886 two_stage_opamp_dummy_magic_25_0.X.n75 two_stage_opamp_dummy_magic_25_0.X.n74 66.0338
R7887 two_stage_opamp_dummy_magic_25_0.X.n6 two_stage_opamp_dummy_magic_25_0.X.n5 49.3505
R7888 two_stage_opamp_dummy_magic_25_0.X.n10 two_stage_opamp_dummy_magic_25_0.X.n9 49.3505
R7889 two_stage_opamp_dummy_magic_25_0.X.n134 two_stage_opamp_dummy_magic_25_0.X.n133 49.3505
R7890 two_stage_opamp_dummy_magic_25_0.X.n140 two_stage_opamp_dummy_magic_25_0.X.n139 49.3505
R7891 two_stage_opamp_dummy_magic_25_0.X.n143 two_stage_opamp_dummy_magic_25_0.X.n142 49.3505
R7892 two_stage_opamp_dummy_magic_25_0.X.n147 two_stage_opamp_dummy_magic_25_0.X.n146 49.3505
R7893 two_stage_opamp_dummy_magic_25_0.X.n41 two_stage_opamp_dummy_magic_25_0.X.t23 41.0384
R7894 two_stage_opamp_dummy_magic_25_0.X.n55 two_stage_opamp_dummy_magic_25_0.X.n50 40.1672
R7895 two_stage_opamp_dummy_magic_25_0.X.n55 two_stage_opamp_dummy_magic_25_0.X.n54 40.1672
R7896 two_stage_opamp_dummy_magic_25_0.X.n34 two_stage_opamp_dummy_magic_25_0.X.n26 40.1672
R7897 two_stage_opamp_dummy_magic_25_0.X.n34 two_stage_opamp_dummy_magic_25_0.X.n33 40.1672
R7898 two_stage_opamp_dummy_magic_25_0.X.n25 two_stage_opamp_dummy_magic_25_0.X.n17 40.1672
R7899 two_stage_opamp_dummy_magic_25_0.X.n25 two_stage_opamp_dummy_magic_25_0.X.n24 40.1672
R7900 two_stage_opamp_dummy_magic_25_0.X.n59 two_stage_opamp_dummy_magic_25_0.X.n58 16.3217
R7901 two_stage_opamp_dummy_magic_25_0.X.n5 two_stage_opamp_dummy_magic_25_0.X.t24 16.0005
R7902 two_stage_opamp_dummy_magic_25_0.X.n5 two_stage_opamp_dummy_magic_25_0.X.t1 16.0005
R7903 two_stage_opamp_dummy_magic_25_0.X.n9 two_stage_opamp_dummy_magic_25_0.X.t2 16.0005
R7904 two_stage_opamp_dummy_magic_25_0.X.n9 two_stage_opamp_dummy_magic_25_0.X.t21 16.0005
R7905 two_stage_opamp_dummy_magic_25_0.X.n133 two_stage_opamp_dummy_magic_25_0.X.t18 16.0005
R7906 two_stage_opamp_dummy_magic_25_0.X.n133 two_stage_opamp_dummy_magic_25_0.X.t0 16.0005
R7907 two_stage_opamp_dummy_magic_25_0.X.n139 two_stage_opamp_dummy_magic_25_0.X.t22 16.0005
R7908 two_stage_opamp_dummy_magic_25_0.X.n139 two_stage_opamp_dummy_magic_25_0.X.t16 16.0005
R7909 two_stage_opamp_dummy_magic_25_0.X.n142 two_stage_opamp_dummy_magic_25_0.X.t19 16.0005
R7910 two_stage_opamp_dummy_magic_25_0.X.n142 two_stage_opamp_dummy_magic_25_0.X.t17 16.0005
R7911 two_stage_opamp_dummy_magic_25_0.X.n146 two_stage_opamp_dummy_magic_25_0.X.t20 16.0005
R7912 two_stage_opamp_dummy_magic_25_0.X.n146 two_stage_opamp_dummy_magic_25_0.X.t5 16.0005
R7913 two_stage_opamp_dummy_magic_25_0.X.n56 two_stage_opamp_dummy_magic_25_0.X.n46 12.8005
R7914 two_stage_opamp_dummy_magic_25_0.X.n78 two_stage_opamp_dummy_magic_25_0.X.t14 11.2576
R7915 two_stage_opamp_dummy_magic_25_0.X.n78 two_stage_opamp_dummy_magic_25_0.X.t3 11.2576
R7916 two_stage_opamp_dummy_magic_25_0.X.n76 two_stage_opamp_dummy_magic_25_0.X.t4 11.2576
R7917 two_stage_opamp_dummy_magic_25_0.X.n76 two_stage_opamp_dummy_magic_25_0.X.t12 11.2576
R7918 two_stage_opamp_dummy_magic_25_0.X.n88 two_stage_opamp_dummy_magic_25_0.X.t15 11.2576
R7919 two_stage_opamp_dummy_magic_25_0.X.n88 two_stage_opamp_dummy_magic_25_0.X.t13 11.2576
R7920 two_stage_opamp_dummy_magic_25_0.X.n84 two_stage_opamp_dummy_magic_25_0.X.t6 11.2576
R7921 two_stage_opamp_dummy_magic_25_0.X.n84 two_stage_opamp_dummy_magic_25_0.X.t7 11.2576
R7922 two_stage_opamp_dummy_magic_25_0.X.n81 two_stage_opamp_dummy_magic_25_0.X.t8 11.2576
R7923 two_stage_opamp_dummy_magic_25_0.X.n81 two_stage_opamp_dummy_magic_25_0.X.t10 11.2576
R7924 two_stage_opamp_dummy_magic_25_0.X.n74 two_stage_opamp_dummy_magic_25_0.X.t9 11.2576
R7925 two_stage_opamp_dummy_magic_25_0.X.n74 two_stage_opamp_dummy_magic_25_0.X.t11 11.2576
R7926 two_stage_opamp_dummy_magic_25_0.X.n56 two_stage_opamp_dummy_magic_25_0.X.n44 9.36264
R7927 two_stage_opamp_dummy_magic_25_0.X.n46 two_stage_opamp_dummy_magic_25_0.X.n45 9.3005
R7928 two_stage_opamp_dummy_magic_25_0.X.n87 two_stage_opamp_dummy_magic_25_0.X.n77 5.91717
R7929 two_stage_opamp_dummy_magic_25_0.X.n80 two_stage_opamp_dummy_magic_25_0.X.n79 5.91717
R7930 two_stage_opamp_dummy_magic_25_0.X.n10 two_stage_opamp_dummy_magic_25_0.X.n8 5.6255
R7931 two_stage_opamp_dummy_magic_25_0.X.n145 two_stage_opamp_dummy_magic_25_0.X.n6 5.6255
R7932 two_stage_opamp_dummy_magic_25_0.X.n58 two_stage_opamp_dummy_magic_25_0.X.n46 5.33141
R7933 two_stage_opamp_dummy_magic_25_0.X.n89 two_stage_opamp_dummy_magic_25_0.X.n87 5.29217
R7934 two_stage_opamp_dummy_magic_25_0.X.n86 two_stage_opamp_dummy_magic_25_0.X.n85 5.29217
R7935 two_stage_opamp_dummy_magic_25_0.X.n83 two_stage_opamp_dummy_magic_25_0.X.n82 5.29217
R7936 two_stage_opamp_dummy_magic_25_0.X.n80 two_stage_opamp_dummy_magic_25_0.X.n75 5.29217
R7937 two_stage_opamp_dummy_magic_25_0.X.n94 two_stage_opamp_dummy_magic_25_0.X.n73 5.1255
R7938 two_stage_opamp_dummy_magic_25_0.X.n91 two_stage_opamp_dummy_magic_25_0.X.n65 5.1255
R7939 two_stage_opamp_dummy_magic_25_0.X.n134 two_stage_opamp_dummy_magic_25_0.X.n8 5.063
R7940 two_stage_opamp_dummy_magic_25_0.X.n141 two_stage_opamp_dummy_magic_25_0.X.n140 5.063
R7941 two_stage_opamp_dummy_magic_25_0.X.n144 two_stage_opamp_dummy_magic_25_0.X.n143 5.063
R7942 two_stage_opamp_dummy_magic_25_0.X.n147 two_stage_opamp_dummy_magic_25_0.X.n145 5.063
R7943 two_stage_opamp_dummy_magic_25_0.X.n150 two_stage_opamp_dummy_magic_25_0.X.n149 5.063
R7944 two_stage_opamp_dummy_magic_25_0.X.n136 two_stage_opamp_dummy_magic_25_0.X.n11 5.063
R7945 two_stage_opamp_dummy_magic_25_0.X.n95 two_stage_opamp_dummy_magic_25_0.X.n94 4.5005
R7946 two_stage_opamp_dummy_magic_25_0.X.n93 two_stage_opamp_dummy_magic_25_0.X.n71 4.5005
R7947 two_stage_opamp_dummy_magic_25_0.X.n92 two_stage_opamp_dummy_magic_25_0.X.n68 4.5005
R7948 two_stage_opamp_dummy_magic_25_0.X.n91 two_stage_opamp_dummy_magic_25_0.X.n90 4.5005
R7949 two_stage_opamp_dummy_magic_25_0.X.n119 two_stage_opamp_dummy_magic_25_0.X.n118 4.5005
R7950 two_stage_opamp_dummy_magic_25_0.X.n149 two_stage_opamp_dummy_magic_25_0.X.n148 4.5005
R7951 two_stage_opamp_dummy_magic_25_0.X.n7 two_stage_opamp_dummy_magic_25_0.X.n3 4.5005
R7952 two_stage_opamp_dummy_magic_25_0.X.n138 two_stage_opamp_dummy_magic_25_0.X.n137 4.5005
R7953 two_stage_opamp_dummy_magic_25_0.X.n136 two_stage_opamp_dummy_magic_25_0.X.n135 4.5005
R7954 two_stage_opamp_dummy_magic_25_0.X.n124 two_stage_opamp_dummy_magic_25_0.X.n61 4.5005
R7955 two_stage_opamp_dummy_magic_25_0.X.n126 two_stage_opamp_dummy_magic_25_0.X.n125 4.5005
R7956 two_stage_opamp_dummy_magic_25_0.X.n125 two_stage_opamp_dummy_magic_25_0.X.n124 4.5005
R7957 two_stage_opamp_dummy_magic_25_0.X.n60 two_stage_opamp_dummy_magic_25_0.X.n59 4.5005
R7958 two_stage_opamp_dummy_magic_25_0.X.n38 two_stage_opamp_dummy_magic_25_0.X.n37 4.5005
R7959 two_stage_opamp_dummy_magic_25_0.X.n120 two_stage_opamp_dummy_magic_25_0.X.n63 2.26187
R7960 two_stage_opamp_dummy_magic_25_0.X.n40 two_stage_opamp_dummy_magic_25_0.X.n39 2.26187
R7961 two_stage_opamp_dummy_magic_25_0.X.n39 two_stage_opamp_dummy_magic_25_0.X.n36 2.26187
R7962 two_stage_opamp_dummy_magic_25_0.X.n117 two_stage_opamp_dummy_magic_25_0.X.n63 2.26187
R7963 two_stage_opamp_dummy_magic_25_0.X.n121 two_stage_opamp_dummy_magic_25_0.X.n62 2.24063
R7964 two_stage_opamp_dummy_magic_25_0.X.n126 two_stage_opamp_dummy_magic_25_0.X.n15 2.24063
R7965 two_stage_opamp_dummy_magic_25_0.X.n16 two_stage_opamp_dummy_magic_25_0.X.n14 2.24063
R7966 two_stage_opamp_dummy_magic_25_0.X.n117 two_stage_opamp_dummy_magic_25_0.X.n116 2.24063
R7967 two_stage_opamp_dummy_magic_25_0.X.n123 two_stage_opamp_dummy_magic_25_0.X.n122 2.24063
R7968 two_stage_opamp_dummy_magic_25_0.X.n41 two_stage_opamp_dummy_magic_25_0.X.n40 2.24063
R7969 two_stage_opamp_dummy_magic_25_0.X.n43 two_stage_opamp_dummy_magic_25_0.X.n42 2.24063
R7970 two_stage_opamp_dummy_magic_25_0.X.n60 two_stage_opamp_dummy_magic_25_0.X.n44 2.22018
R7971 two_stage_opamp_dummy_magic_25_0.X.n98 two_stage_opamp_dummy_magic_25_0.X.n72 1.5005
R7972 two_stage_opamp_dummy_magic_25_0.X.n100 two_stage_opamp_dummy_magic_25_0.X.n99 1.5005
R7973 two_stage_opamp_dummy_magic_25_0.X.n101 two_stage_opamp_dummy_magic_25_0.X.n70 1.5005
R7974 two_stage_opamp_dummy_magic_25_0.X.n103 two_stage_opamp_dummy_magic_25_0.X.n102 1.5005
R7975 two_stage_opamp_dummy_magic_25_0.X.n104 two_stage_opamp_dummy_magic_25_0.X.n69 1.5005
R7976 two_stage_opamp_dummy_magic_25_0.X.n106 two_stage_opamp_dummy_magic_25_0.X.n105 1.5005
R7977 two_stage_opamp_dummy_magic_25_0.X.n107 two_stage_opamp_dummy_magic_25_0.X.n67 1.5005
R7978 two_stage_opamp_dummy_magic_25_0.X.n109 two_stage_opamp_dummy_magic_25_0.X.n108 1.5005
R7979 two_stage_opamp_dummy_magic_25_0.X.n110 two_stage_opamp_dummy_magic_25_0.X.n66 1.5005
R7980 two_stage_opamp_dummy_magic_25_0.X.n112 two_stage_opamp_dummy_magic_25_0.X.n111 1.5005
R7981 two_stage_opamp_dummy_magic_25_0.X.n113 two_stage_opamp_dummy_magic_25_0.X.n64 1.5005
R7982 two_stage_opamp_dummy_magic_25_0.X.n115 two_stage_opamp_dummy_magic_25_0.X.n114 1.5005
R7983 two_stage_opamp_dummy_magic_25_0.X.n153 two_stage_opamp_dummy_magic_25_0.X.n152 1.5005
R7984 two_stage_opamp_dummy_magic_25_0.X.n154 two_stage_opamp_dummy_magic_25_0.X.n1 1.5005
R7985 two_stage_opamp_dummy_magic_25_0.X.n156 two_stage_opamp_dummy_magic_25_0.X.n155 1.5005
R7986 two_stage_opamp_dummy_magic_25_0.X.n2 two_stage_opamp_dummy_magic_25_0.X.n0 1.5005
R7987 two_stage_opamp_dummy_magic_25_0.X.n130 two_stage_opamp_dummy_magic_25_0.X.n13 1.5005
R7988 two_stage_opamp_dummy_magic_25_0.X.n132 two_stage_opamp_dummy_magic_25_0.X.n131 1.5005
R7989 two_stage_opamp_dummy_magic_25_0.X.n129 two_stage_opamp_dummy_magic_25_0.X.n12 1.5005
R7990 two_stage_opamp_dummy_magic_25_0.X.n128 two_stage_opamp_dummy_magic_25_0.X.n127 1.5005
R7991 two_stage_opamp_dummy_magic_25_0.X.n151 two_stage_opamp_dummy_magic_25_0.X.n150 1.43397
R7992 two_stage_opamp_dummy_magic_25_0.X.n135 two_stage_opamp_dummy_magic_25_0.X.n132 1.3755
R7993 two_stage_opamp_dummy_magic_25_0.X.n138 two_stage_opamp_dummy_magic_25_0.X.n2 1.3755
R7994 two_stage_opamp_dummy_magic_25_0.X.n154 two_stage_opamp_dummy_magic_25_0.X.n3 1.3755
R7995 two_stage_opamp_dummy_magic_25_0.X.n148 two_stage_opamp_dummy_magic_25_0.X.n4 1.3755
R7996 two_stage_opamp_dummy_magic_25_0.X.n127 two_stage_opamp_dummy_magic_25_0.X.n11 1.3755
R7997 two_stage_opamp_dummy_magic_25_0.X.n122 two_stage_opamp_dummy_magic_25_0.X.n121 0.979667
R7998 two_stage_opamp_dummy_magic_25_0.X.n90 two_stage_opamp_dummy_magic_25_0.X.n89 0.792167
R7999 two_stage_opamp_dummy_magic_25_0.X.n85 two_stage_opamp_dummy_magic_25_0.X.n68 0.792167
R8000 two_stage_opamp_dummy_magic_25_0.X.n82 two_stage_opamp_dummy_magic_25_0.X.n71 0.792167
R8001 two_stage_opamp_dummy_magic_25_0.X.n95 two_stage_opamp_dummy_magic_25_0.X.n75 0.792167
R8002 two_stage_opamp_dummy_magic_25_0.X.n77 two_stage_opamp_dummy_magic_25_0.X.n65 0.792167
R8003 two_stage_opamp_dummy_magic_25_0.X.n79 two_stage_opamp_dummy_magic_25_0.X.n73 0.792167
R8004 two_stage_opamp_dummy_magic_25_0.X.n60 two_stage_opamp_dummy_magic_25_0.X.n43 0.682792
R8005 two_stage_opamp_dummy_magic_25_0.X.n128 two_stage_opamp_dummy_magic_25_0.X.n126 0.630708
R8006 two_stage_opamp_dummy_magic_25_0.X.n94 two_stage_opamp_dummy_magic_25_0.X.n93 0.6255
R8007 two_stage_opamp_dummy_magic_25_0.X.n93 two_stage_opamp_dummy_magic_25_0.X.n92 0.6255
R8008 two_stage_opamp_dummy_magic_25_0.X.n92 two_stage_opamp_dummy_magic_25_0.X.n91 0.6255
R8009 two_stage_opamp_dummy_magic_25_0.X.n87 two_stage_opamp_dummy_magic_25_0.X.n86 0.6255
R8010 two_stage_opamp_dummy_magic_25_0.X.n86 two_stage_opamp_dummy_magic_25_0.X.n83 0.6255
R8011 two_stage_opamp_dummy_magic_25_0.X.n83 two_stage_opamp_dummy_magic_25_0.X.n80 0.6255
R8012 two_stage_opamp_dummy_magic_25_0.X.n116 two_stage_opamp_dummy_magic_25_0.X.n115 0.609875
R8013 two_stage_opamp_dummy_magic_25_0.X.n152 two_stage_opamp_dummy_magic_25_0.X.n151 0.564601
R8014 two_stage_opamp_dummy_magic_25_0.X.n149 two_stage_opamp_dummy_magic_25_0.X.n7 0.563
R8015 two_stage_opamp_dummy_magic_25_0.X.n137 two_stage_opamp_dummy_magic_25_0.X.n7 0.563
R8016 two_stage_opamp_dummy_magic_25_0.X.n137 two_stage_opamp_dummy_magic_25_0.X.n136 0.563
R8017 two_stage_opamp_dummy_magic_25_0.X.n141 two_stage_opamp_dummy_magic_25_0.X.n8 0.563
R8018 two_stage_opamp_dummy_magic_25_0.X.n144 two_stage_opamp_dummy_magic_25_0.X.n141 0.563
R8019 two_stage_opamp_dummy_magic_25_0.X.n145 two_stage_opamp_dummy_magic_25_0.X.n144 0.563
R8020 two_stage_opamp_dummy_magic_25_0.X.n97 two_stage_opamp_dummy_magic_25_0.X.n73 0.533638
R8021 two_stage_opamp_dummy_magic_25_0.X.n90 two_stage_opamp_dummy_magic_25_0.X.n66 0.46925
R8022 two_stage_opamp_dummy_magic_25_0.X.n106 two_stage_opamp_dummy_magic_25_0.X.n68 0.46925
R8023 two_stage_opamp_dummy_magic_25_0.X.n101 two_stage_opamp_dummy_magic_25_0.X.n71 0.46925
R8024 two_stage_opamp_dummy_magic_25_0.X.n96 two_stage_opamp_dummy_magic_25_0.X.n95 0.46925
R8025 two_stage_opamp_dummy_magic_25_0.X.n114 two_stage_opamp_dummy_magic_25_0.X.n65 0.46925
R8026 two_stage_opamp_dummy_magic_25_0.X.n124 two_stage_opamp_dummy_magic_25_0.X.n60 0.46925
R8027 two_stage_opamp_dummy_magic_25_0.X.n98 two_stage_opamp_dummy_magic_25_0.X.n97 0.427973
R8028 two_stage_opamp_dummy_magic_25_0.X.n135 two_stage_opamp_dummy_magic_25_0.X.n134 0.3755
R8029 two_stage_opamp_dummy_magic_25_0.X.n140 two_stage_opamp_dummy_magic_25_0.X.n138 0.3755
R8030 two_stage_opamp_dummy_magic_25_0.X.n143 two_stage_opamp_dummy_magic_25_0.X.n3 0.3755
R8031 two_stage_opamp_dummy_magic_25_0.X.n148 two_stage_opamp_dummy_magic_25_0.X.n147 0.3755
R8032 two_stage_opamp_dummy_magic_25_0.X.n11 two_stage_opamp_dummy_magic_25_0.X.n10 0.3755
R8033 two_stage_opamp_dummy_magic_25_0.X.n150 two_stage_opamp_dummy_magic_25_0.X.n6 0.3755
R8034 two_stage_opamp_dummy_magic_25_0.X.n59 two_stage_opamp_dummy_magic_25_0.X.n45 0.1255
R8035 two_stage_opamp_dummy_magic_25_0.X.n45 two_stage_opamp_dummy_magic_25_0.X.n44 0.0626438
R8036 two_stage_opamp_dummy_magic_25_0.X.n97 two_stage_opamp_dummy_magic_25_0.X.n96 0.0587394
R8037 two_stage_opamp_dummy_magic_25_0.X.n127 two_stage_opamp_dummy_magic_25_0.X.n12 0.0577917
R8038 two_stage_opamp_dummy_magic_25_0.X.n132 two_stage_opamp_dummy_magic_25_0.X.n12 0.0577917
R8039 two_stage_opamp_dummy_magic_25_0.X.n132 two_stage_opamp_dummy_magic_25_0.X.n13 0.0577917
R8040 two_stage_opamp_dummy_magic_25_0.X.n13 two_stage_opamp_dummy_magic_25_0.X.n2 0.0577917
R8041 two_stage_opamp_dummy_magic_25_0.X.n155 two_stage_opamp_dummy_magic_25_0.X.n2 0.0577917
R8042 two_stage_opamp_dummy_magic_25_0.X.n155 two_stage_opamp_dummy_magic_25_0.X.n154 0.0577917
R8043 two_stage_opamp_dummy_magic_25_0.X.n154 two_stage_opamp_dummy_magic_25_0.X.n153 0.0577917
R8044 two_stage_opamp_dummy_magic_25_0.X.n153 two_stage_opamp_dummy_magic_25_0.X.n4 0.0577917
R8045 two_stage_opamp_dummy_magic_25_0.X.n129 two_stage_opamp_dummy_magic_25_0.X.n128 0.0577917
R8046 two_stage_opamp_dummy_magic_25_0.X.n131 two_stage_opamp_dummy_magic_25_0.X.n129 0.0577917
R8047 two_stage_opamp_dummy_magic_25_0.X.n131 two_stage_opamp_dummy_magic_25_0.X.n130 0.0577917
R8048 two_stage_opamp_dummy_magic_25_0.X.n130 two_stage_opamp_dummy_magic_25_0.X.n0 0.0577917
R8049 two_stage_opamp_dummy_magic_25_0.X.n156 two_stage_opamp_dummy_magic_25_0.X.n1 0.0577917
R8050 two_stage_opamp_dummy_magic_25_0.X.n152 two_stage_opamp_dummy_magic_25_0.X.n1 0.0577917
R8051 two_stage_opamp_dummy_magic_25_0.X.n151 two_stage_opamp_dummy_magic_25_0.X.n4 0.054517
R8052 two_stage_opamp_dummy_magic_25_0.X.n114 two_stage_opamp_dummy_magic_25_0.X.n113 0.0421667
R8053 two_stage_opamp_dummy_magic_25_0.X.n113 two_stage_opamp_dummy_magic_25_0.X.n112 0.0421667
R8054 two_stage_opamp_dummy_magic_25_0.X.n112 two_stage_opamp_dummy_magic_25_0.X.n66 0.0421667
R8055 two_stage_opamp_dummy_magic_25_0.X.n108 two_stage_opamp_dummy_magic_25_0.X.n66 0.0421667
R8056 two_stage_opamp_dummy_magic_25_0.X.n108 two_stage_opamp_dummy_magic_25_0.X.n107 0.0421667
R8057 two_stage_opamp_dummy_magic_25_0.X.n107 two_stage_opamp_dummy_magic_25_0.X.n106 0.0421667
R8058 two_stage_opamp_dummy_magic_25_0.X.n106 two_stage_opamp_dummy_magic_25_0.X.n69 0.0421667
R8059 two_stage_opamp_dummy_magic_25_0.X.n102 two_stage_opamp_dummy_magic_25_0.X.n69 0.0421667
R8060 two_stage_opamp_dummy_magic_25_0.X.n102 two_stage_opamp_dummy_magic_25_0.X.n101 0.0421667
R8061 two_stage_opamp_dummy_magic_25_0.X.n101 two_stage_opamp_dummy_magic_25_0.X.n100 0.0421667
R8062 two_stage_opamp_dummy_magic_25_0.X.n100 two_stage_opamp_dummy_magic_25_0.X.n72 0.0421667
R8063 two_stage_opamp_dummy_magic_25_0.X.n96 two_stage_opamp_dummy_magic_25_0.X.n72 0.0421667
R8064 two_stage_opamp_dummy_magic_25_0.X.n115 two_stage_opamp_dummy_magic_25_0.X.n64 0.0421667
R8065 two_stage_opamp_dummy_magic_25_0.X.n111 two_stage_opamp_dummy_magic_25_0.X.n64 0.0421667
R8066 two_stage_opamp_dummy_magic_25_0.X.n111 two_stage_opamp_dummy_magic_25_0.X.n110 0.0421667
R8067 two_stage_opamp_dummy_magic_25_0.X.n110 two_stage_opamp_dummy_magic_25_0.X.n109 0.0421667
R8068 two_stage_opamp_dummy_magic_25_0.X.n109 two_stage_opamp_dummy_magic_25_0.X.n67 0.0421667
R8069 two_stage_opamp_dummy_magic_25_0.X.n105 two_stage_opamp_dummy_magic_25_0.X.n67 0.0421667
R8070 two_stage_opamp_dummy_magic_25_0.X.n105 two_stage_opamp_dummy_magic_25_0.X.n104 0.0421667
R8071 two_stage_opamp_dummy_magic_25_0.X.n104 two_stage_opamp_dummy_magic_25_0.X.n103 0.0421667
R8072 two_stage_opamp_dummy_magic_25_0.X.n103 two_stage_opamp_dummy_magic_25_0.X.n70 0.0421667
R8073 two_stage_opamp_dummy_magic_25_0.X.n99 two_stage_opamp_dummy_magic_25_0.X.n70 0.0421667
R8074 two_stage_opamp_dummy_magic_25_0.X.n99 two_stage_opamp_dummy_magic_25_0.X.n98 0.0421667
R8075 two_stage_opamp_dummy_magic_25_0.X.n126 two_stage_opamp_dummy_magic_25_0.X.n14 0.0421667
R8076 two_stage_opamp_dummy_magic_25_0.X two_stage_opamp_dummy_magic_25_0.X.n156 0.0369583
R8077 two_stage_opamp_dummy_magic_25_0.X.n116 two_stage_opamp_dummy_magic_25_0.X.n62 0.0217373
R8078 two_stage_opamp_dummy_magic_25_0.X.n120 two_stage_opamp_dummy_magic_25_0.X.n119 0.0217373
R8079 two_stage_opamp_dummy_magic_25_0.X.n122 two_stage_opamp_dummy_magic_25_0.X.n15 0.0217373
R8080 two_stage_opamp_dummy_magic_25_0.X.n125 two_stage_opamp_dummy_magic_25_0.X.n16 0.0217373
R8081 two_stage_opamp_dummy_magic_25_0.X.n118 two_stage_opamp_dummy_magic_25_0.X.n62 0.0217373
R8082 two_stage_opamp_dummy_magic_25_0.X.n121 two_stage_opamp_dummy_magic_25_0.X.n120 0.0217373
R8083 two_stage_opamp_dummy_magic_25_0.X.n43 two_stage_opamp_dummy_magic_25_0.X.n36 0.0217373
R8084 two_stage_opamp_dummy_magic_25_0.X.n61 two_stage_opamp_dummy_magic_25_0.X.n15 0.0217373
R8085 two_stage_opamp_dummy_magic_25_0.X.n61 two_stage_opamp_dummy_magic_25_0.X.n16 0.0217373
R8086 two_stage_opamp_dummy_magic_25_0.X.n39 two_stage_opamp_dummy_magic_25_0.X.n37 0.0217373
R8087 two_stage_opamp_dummy_magic_25_0.X.n38 two_stage_opamp_dummy_magic_25_0.X.n36 0.0217373
R8088 two_stage_opamp_dummy_magic_25_0.X.n118 two_stage_opamp_dummy_magic_25_0.X.n63 0.0217373
R8089 two_stage_opamp_dummy_magic_25_0.X.n119 two_stage_opamp_dummy_magic_25_0.X.n117 0.0217373
R8090 two_stage_opamp_dummy_magic_25_0.X.n40 two_stage_opamp_dummy_magic_25_0.X.n38 0.0217373
R8091 two_stage_opamp_dummy_magic_25_0.X.n124 two_stage_opamp_dummy_magic_25_0.X.n123 0.0217373
R8092 two_stage_opamp_dummy_magic_25_0.X.n123 two_stage_opamp_dummy_magic_25_0.X.n14 0.0217373
R8093 two_stage_opamp_dummy_magic_25_0.X.n42 two_stage_opamp_dummy_magic_25_0.X.n37 0.0217373
R8094 two_stage_opamp_dummy_magic_25_0.X.n42 two_stage_opamp_dummy_magic_25_0.X.n41 0.0217373
R8095 two_stage_opamp_dummy_magic_25_0.X two_stage_opamp_dummy_magic_25_0.X.n0 0.0213333
R8096 GNDA.n6987 GNDA.n6986 479844
R8097 GNDA.n5319 GNDA.n315 401768
R8098 GNDA.n5319 GNDA.n5318 145595
R8099 GNDA.n6986 GNDA.n314 103560
R8100 GNDA.n6986 GNDA.n6985 71285.5
R8101 GNDA.n6987 GNDA.t325 55309.3
R8102 GNDA.n6992 GNDA.n311 51271.7
R8103 GNDA.n6993 GNDA.n310 25810.5
R8104 GNDA.n1748 GNDA.n313 14443.6
R8105 GNDA.n312 GNDA.n311 13807.5
R8106 GNDA.n5320 GNDA.n312 13460.8
R8107 GNDA.n6984 GNDA.n310 11878.2
R8108 GNDA.n6985 GNDA.n6984 9755.2
R8109 GNDA.n311 GNDA.n310 8531.5
R8110 GNDA.n1752 GNDA.n1748 7511.38
R8111 GNDA.n1748 GNDA.n1747 7511.38
R8112 GNDA.n6991 GNDA.n312 7115.05
R8113 GNDA.n6989 GNDA.n6988 5032.34
R8114 GNDA.n6990 GNDA.n314 4738.46
R8115 GNDA.n6989 GNDA.n315 4544.93
R8116 GNDA.n6985 GNDA.n5320 4106.67
R8117 GNDA.n6984 GNDA.n6983 3974.19
R8118 GNDA.n1751 GNDA.n1749 3925.98
R8119 GNDA.n1751 GNDA.n1750 3882.89
R8120 GNDA.n6988 GNDA.t70 3252.41
R8121 GNDA.n6988 GNDA.t67 2442.21
R8122 GNDA.n6993 GNDA.n6992 2413.89
R8123 GNDA.t34 GNDA.n1749 1968.35
R8124 GNDA.n7413 GNDA.n7412 1518.49
R8125 GNDA.n6992 GNDA.n6991 1295.8
R8126 GNDA.n5320 GNDA.n314 1031.25
R8127 GNDA.n1749 GNDA.n313 970.167
R8128 GNDA.n5316 GNDA.t204 749.742
R8129 GNDA.n3403 GNDA.t151 747.734
R8130 GNDA.n3400 GNDA.t240 747.734
R8131 GNDA.n5313 GNDA.t225 747.734
R8132 GNDA.t283 GNDA.n6993 697.547
R8133 GNDA.n6776 GNDA.n6775 686.717
R8134 GNDA.n6793 GNDA.n6792 686.717
R8135 GNDA.n6785 GNDA.n6649 686.717
R8136 GNDA.n6767 GNDA.n6763 686.717
R8137 GNDA.n6938 GNDA.n6937 669.307
R8138 GNDA.n6954 GNDA.n6953 669.307
R8139 GNDA.n7239 GNDA.n7236 669.307
R8140 GNDA.n1707 GNDA.t237 659.367
R8141 GNDA.n1706 GNDA.t158 659.367
R8142 GNDA.n5282 GNDA.t171 659.367
R8143 GNDA.n5305 GNDA.t219 659.367
R8144 GNDA.n5408 GNDA.n5407 585.003
R8145 GNDA.n6645 GNDA.n6644 585.001
R8146 GNDA.n6648 GNDA.n6647 585.001
R8147 GNDA.n5386 GNDA.n5385 585.001
R8148 GNDA.n6957 GNDA.n6956 585.001
R8149 GNDA.n5363 GNDA.n5362 585.001
R8150 GNDA.n5365 GNDA.n5364 585.001
R8151 GNDA.n7033 GNDA.n7032 585.001
R8152 GNDA.n7238 GNDA.n7237 585
R8153 GNDA.n89 GNDA.n86 585
R8154 GNDA.t145 GNDA.n89 585
R8155 GNDA.n6300 GNDA.n6299 585
R8156 GNDA.n6300 GNDA.n77 585
R8157 GNDA.n6301 GNDA.n6267 585
R8158 GNDA.n6302 GNDA.n6301 585
R8159 GNDA.n6305 GNDA.n6304 585
R8160 GNDA.n6304 GNDA.n6303 585
R8161 GNDA.n6306 GNDA.n6266 585
R8162 GNDA.n6266 GNDA.n6265 585
R8163 GNDA.n6308 GNDA.n6307 585
R8164 GNDA.n6309 GNDA.n6308 585
R8165 GNDA.n6264 GNDA.n6263 585
R8166 GNDA.n6310 GNDA.n6264 585
R8167 GNDA.n6313 GNDA.n6312 585
R8168 GNDA.n6312 GNDA.n6311 585
R8169 GNDA.n6314 GNDA.n6262 585
R8170 GNDA.n6262 GNDA.n6261 585
R8171 GNDA.n6316 GNDA.n6315 585
R8172 GNDA.n6317 GNDA.n6316 585
R8173 GNDA.n6259 GNDA.n6258 585
R8174 GNDA.n6318 GNDA.n6259 585
R8175 GNDA.n6321 GNDA.n6320 585
R8176 GNDA.n6320 GNDA.n6319 585
R8177 GNDA.n6322 GNDA.n6257 585
R8178 GNDA.n6260 GNDA.n6257 585
R8179 GNDA.n7465 GNDA.n67 585
R8180 GNDA.n7468 GNDA.n7467 585
R8181 GNDA.n71 GNDA.n70 585
R8182 GNDA.n6281 GNDA.n6280 585
R8183 GNDA.n6282 GNDA.n6279 585
R8184 GNDA.n6276 GNDA.n6275 585
R8185 GNDA.n6288 GNDA.n6274 585
R8186 GNDA.n6289 GNDA.n6273 585
R8187 GNDA.n6290 GNDA.n6272 585
R8188 GNDA.n6270 GNDA.n6269 585
R8189 GNDA.n6296 GNDA.n6268 585
R8190 GNDA.n6298 GNDA.n6297 585
R8191 GNDA.n6297 GNDA.n79 585
R8192 GNDA.n6296 GNDA.n6295 585
R8193 GNDA.n6293 GNDA.n6270 585
R8194 GNDA.n6291 GNDA.n6290 585
R8195 GNDA.n6289 GNDA.n6271 585
R8196 GNDA.n6288 GNDA.n6287 585
R8197 GNDA.n6285 GNDA.n6276 585
R8198 GNDA.n6283 GNDA.n6282 585
R8199 GNDA.n6281 GNDA.n6278 585
R8200 GNDA.n70 GNDA.n69 585
R8201 GNDA.n7469 GNDA.n7468 585
R8202 GNDA.n7471 GNDA.n67 585
R8203 GNDA.n6100 GNDA.n6099 585
R8204 GNDA.n6101 GNDA.n6082 585
R8205 GNDA.n6103 GNDA.n6102 585
R8206 GNDA.n6105 GNDA.n6080 585
R8207 GNDA.n6107 GNDA.n6106 585
R8208 GNDA.n6108 GNDA.n6079 585
R8209 GNDA.n6110 GNDA.n6109 585
R8210 GNDA.n6112 GNDA.n6077 585
R8211 GNDA.n6114 GNDA.n6113 585
R8212 GNDA.n6115 GNDA.n6076 585
R8213 GNDA.n6117 GNDA.n6116 585
R8214 GNDA.n6119 GNDA.n6075 585
R8215 GNDA.n5997 GNDA.n5996 585
R8216 GNDA.n5994 GNDA.n5514 585
R8217 GNDA.n5885 GNDA.n5884 585
R8218 GNDA.n5989 GNDA.n5988 585
R8219 GNDA.n5987 GNDA.n5986 585
R8220 GNDA.n5913 GNDA.n5889 585
R8221 GNDA.n5915 GNDA.n5914 585
R8222 GNDA.n5920 GNDA.n5919 585
R8223 GNDA.n5918 GNDA.n5911 585
R8224 GNDA.n5926 GNDA.n5925 585
R8225 GNDA.n5928 GNDA.n5927 585
R8226 GNDA.n5909 GNDA.n5908 585
R8227 GNDA.n6068 GNDA.n6067 585
R8228 GNDA.n6065 GNDA.n6064 585
R8229 GNDA.n6063 GNDA.n6062 585
R8230 GNDA.n5487 GNDA.n5454 585
R8231 GNDA.n5507 GNDA.n5506 585
R8232 GNDA.n5503 GNDA.n5486 585
R8233 GNDA.n5490 GNDA.n5489 585
R8234 GNDA.n5498 GNDA.n5497 585
R8235 GNDA.n5496 GNDA.n5495 585
R8236 GNDA.n5475 GNDA.n5474 585
R8237 GNDA.n6002 GNDA.n6001 585
R8238 GNDA.n5477 GNDA.n5476 585
R8239 GNDA.n5716 GNDA.n5445 585
R8240 GNDA.n5740 GNDA.n5718 585
R8241 GNDA.n5742 GNDA.n5741 585
R8242 GNDA.n5738 GNDA.n5737 585
R8243 GNDA.n5736 GNDA.n5735 585
R8244 GNDA.n5731 GNDA.n5730 585
R8245 GNDA.n5729 GNDA.n5728 585
R8246 GNDA.n5724 GNDA.n5723 585
R8247 GNDA.n5722 GNDA.n5643 585
R8248 GNDA.n5750 GNDA.n5749 585
R8249 GNDA.n5752 GNDA.n5751 585
R8250 GNDA.n5755 GNDA.n5754 585
R8251 GNDA.n6153 GNDA.n6152 585
R8252 GNDA.n6154 GNDA.n5441 585
R8253 GNDA.n6156 GNDA.n6155 585
R8254 GNDA.n6158 GNDA.n5440 585
R8255 GNDA.n6161 GNDA.n6160 585
R8256 GNDA.n6162 GNDA.n5439 585
R8257 GNDA.n6164 GNDA.n6163 585
R8258 GNDA.n6166 GNDA.n5438 585
R8259 GNDA.n6169 GNDA.n6168 585
R8260 GNDA.n6170 GNDA.n5437 585
R8261 GNDA.n6172 GNDA.n6171 585
R8262 GNDA.n6174 GNDA.n5434 585
R8263 GNDA.n6212 GNDA.n6211 585
R8264 GNDA.n6214 GNDA.n5432 585
R8265 GNDA.n6217 GNDA.n6216 585
R8266 GNDA.n6218 GNDA.n5431 585
R8267 GNDA.n6220 GNDA.n6219 585
R8268 GNDA.n6222 GNDA.n5430 585
R8269 GNDA.n6225 GNDA.n6224 585
R8270 GNDA.n6226 GNDA.n5429 585
R8271 GNDA.n6228 GNDA.n6227 585
R8272 GNDA.n6230 GNDA.n5428 585
R8273 GNDA.n6233 GNDA.n6232 585
R8274 GNDA.n6234 GNDA.n5427 585
R8275 GNDA.n6914 GNDA.n5389 585
R8276 GNDA.n6917 GNDA.n6916 585
R8277 GNDA.n5392 GNDA.n5391 585
R8278 GNDA.n6191 GNDA.n6190 585
R8279 GNDA.n6196 GNDA.n6188 585
R8280 GNDA.n6197 GNDA.n6186 585
R8281 GNDA.n6198 GNDA.n6185 585
R8282 GNDA.n6183 GNDA.n6181 585
R8283 GNDA.n6203 GNDA.n6180 585
R8284 GNDA.n6204 GNDA.n6178 585
R8285 GNDA.n6177 GNDA.n5436 585
R8286 GNDA.n6209 GNDA.n5433 585
R8287 GNDA.n6209 GNDA.n6208 585
R8288 GNDA.n6206 GNDA.n5436 585
R8289 GNDA.n6205 GNDA.n6204 585
R8290 GNDA.n6203 GNDA.n6202 585
R8291 GNDA.n6201 GNDA.n6181 585
R8292 GNDA.n6199 GNDA.n6198 585
R8293 GNDA.n6197 GNDA.n6182 585
R8294 GNDA.n6196 GNDA.n6195 585
R8295 GNDA.n6193 GNDA.n6191 585
R8296 GNDA.n5391 GNDA.n5390 585
R8297 GNDA.n6918 GNDA.n6917 585
R8298 GNDA.n6920 GNDA.n5389 585
R8299 GNDA.n5447 GNDA.n5435 585
R8300 GNDA.n6070 GNDA.n5447 585
R8301 GNDA.n6069 GNDA.n5435 585
R8302 GNDA.n6070 GNDA.n6069 585
R8303 GNDA.n5550 GNDA.n5549 585
R8304 GNDA.n5551 GNDA.n5547 585
R8305 GNDA.n5554 GNDA.n5546 585
R8306 GNDA.n5555 GNDA.n5544 585
R8307 GNDA.n5558 GNDA.n5543 585
R8308 GNDA.n5559 GNDA.n5541 585
R8309 GNDA.n5562 GNDA.n5540 585
R8310 GNDA.n5563 GNDA.n5538 585
R8311 GNDA.n5564 GNDA.n5537 585
R8312 GNDA.n5529 GNDA.n5528 585
R8313 GNDA.n5835 GNDA.n5834 585
R8314 GNDA.n5837 GNDA.n5526 585
R8315 GNDA.n5831 GNDA.n5526 585
R8316 GNDA.n5834 GNDA.n5833 585
R8317 GNDA.n5530 GNDA.n5529 585
R8318 GNDA.n5565 GNDA.n5564 585
R8319 GNDA.n5563 GNDA.n5535 585
R8320 GNDA.n5562 GNDA.n5561 585
R8321 GNDA.n5560 GNDA.n5559 585
R8322 GNDA.n5558 GNDA.n5557 585
R8323 GNDA.n5556 GNDA.n5555 585
R8324 GNDA.n5554 GNDA.n5553 585
R8325 GNDA.n5552 GNDA.n5551 585
R8326 GNDA.n5550 GNDA.n5448 585
R8327 GNDA.n5839 GNDA.n5838 585
R8328 GNDA.n5840 GNDA.n5523 585
R8329 GNDA.n5842 GNDA.n5841 585
R8330 GNDA.n5844 GNDA.n5521 585
R8331 GNDA.n5846 GNDA.n5845 585
R8332 GNDA.n5847 GNDA.n5520 585
R8333 GNDA.n5849 GNDA.n5848 585
R8334 GNDA.n5851 GNDA.n5518 585
R8335 GNDA.n5853 GNDA.n5852 585
R8336 GNDA.n5854 GNDA.n5517 585
R8337 GNDA.n5856 GNDA.n5855 585
R8338 GNDA.n5858 GNDA.n5515 585
R8339 GNDA.n5811 GNDA.n5810 585
R8340 GNDA.n5812 GNDA.n5575 585
R8341 GNDA.n5814 GNDA.n5813 585
R8342 GNDA.n5816 GNDA.n5573 585
R8343 GNDA.n5818 GNDA.n5817 585
R8344 GNDA.n5819 GNDA.n5572 585
R8345 GNDA.n5821 GNDA.n5820 585
R8346 GNDA.n5823 GNDA.n5570 585
R8347 GNDA.n5825 GNDA.n5824 585
R8348 GNDA.n5826 GNDA.n5569 585
R8349 GNDA.n5828 GNDA.n5827 585
R8350 GNDA.n5830 GNDA.n5568 585
R8351 GNDA.n5783 GNDA.n5782 585
R8352 GNDA.n5784 GNDA.n5626 585
R8353 GNDA.n5786 GNDA.n5785 585
R8354 GNDA.n5788 GNDA.n5624 585
R8355 GNDA.n5790 GNDA.n5789 585
R8356 GNDA.n5791 GNDA.n5623 585
R8357 GNDA.n5793 GNDA.n5792 585
R8358 GNDA.n5795 GNDA.n5621 585
R8359 GNDA.n5797 GNDA.n5796 585
R8360 GNDA.n5798 GNDA.n5620 585
R8361 GNDA.n5800 GNDA.n5799 585
R8362 GNDA.n5802 GNDA.n5619 585
R8363 GNDA.n65 GNDA.n64 585
R8364 GNDA.n7473 GNDA.n64 585
R8365 GNDA.n6546 GNDA.n6545 585
R8366 GNDA.n6543 GNDA.n6542 585
R8367 GNDA.n6541 GNDA.n6540 585
R8368 GNDA.n6457 GNDA.n6325 585
R8369 GNDA.n6459 GNDA.n6458 585
R8370 GNDA.n6463 GNDA.n6462 585
R8371 GNDA.n6465 GNDA.n6464 585
R8372 GNDA.n6472 GNDA.n6471 585
R8373 GNDA.n6470 GNDA.n6455 585
R8374 GNDA.n6478 GNDA.n6477 585
R8375 GNDA.n6480 GNDA.n6479 585
R8376 GNDA.n6453 GNDA.n6452 585
R8377 GNDA.n7472 GNDA.n65 585
R8378 GNDA.n7473 GNDA.n7472 585
R8379 GNDA.n6450 GNDA.n66 585
R8380 GNDA.n6448 GNDA.n6447 585
R8381 GNDA.n6446 GNDA.n6445 585
R8382 GNDA.n6356 GNDA.n6346 585
R8383 GNDA.n6358 GNDA.n6357 585
R8384 GNDA.n6362 GNDA.n6361 585
R8385 GNDA.n6364 GNDA.n6363 585
R8386 GNDA.n6370 GNDA.n6369 585
R8387 GNDA.n6372 GNDA.n6371 585
R8388 GNDA.n6373 GNDA.n55 585
R8389 GNDA.n7480 GNDA.n7479 585
R8390 GNDA.n7477 GNDA.n54 585
R8391 GNDA.n63 GNDA.n58 585
R8392 GNDA.n24 GNDA.n22 585
R8393 GNDA.n7485 GNDA.n7484 585
R8394 GNDA.n32 GNDA.n25 585
R8395 GNDA.n40 GNDA.n39 585
R8396 GNDA.n35 GNDA.n31 585
R8397 GNDA.n30 GNDA.n0 585
R8398 GNDA.n7374 GNDA.n1 585
R8399 GNDA.n7376 GNDA.n7375 585
R8400 GNDA.n7380 GNDA.n7379 585
R8401 GNDA.n7382 GNDA.n7381 585
R8402 GNDA.n7385 GNDA.n7384 585
R8403 GNDA.n7304 GNDA.n7303 585
R8404 GNDA.n7413 GNDA.n7304 585
R8405 GNDA.n7416 GNDA.n7415 585
R8406 GNDA.n7415 GNDA.n7414 585
R8407 GNDA.n7417 GNDA.n7302 585
R8408 GNDA.n7302 GNDA.n7301 585
R8409 GNDA.n7419 GNDA.n7418 585
R8410 GNDA.n7420 GNDA.n7419 585
R8411 GNDA.n7300 GNDA.n7299 585
R8412 GNDA.n7421 GNDA.n7300 585
R8413 GNDA.n7424 GNDA.n7423 585
R8414 GNDA.n7423 GNDA.n7422 585
R8415 GNDA.n7425 GNDA.n7298 585
R8416 GNDA.n7298 GNDA.n7297 585
R8417 GNDA.n7427 GNDA.n7426 585
R8418 GNDA.n7428 GNDA.n7427 585
R8419 GNDA.n7296 GNDA.n7295 585
R8420 GNDA.n7429 GNDA.n7296 585
R8421 GNDA.n7432 GNDA.n7431 585
R8422 GNDA.n7431 GNDA.n7430 585
R8423 GNDA.n7433 GNDA.n7248 585
R8424 GNDA.n7248 GNDA.n7246 585
R8425 GNDA.n7435 GNDA.n7434 585
R8426 GNDA.n7436 GNDA.n7435 585
R8427 GNDA.n7243 GNDA.n7242 585
R8428 GNDA.n7438 GNDA.n7243 585
R8429 GNDA.n7441 GNDA.n7440 585
R8430 GNDA.n7440 GNDA.n7439 585
R8431 GNDA.n7442 GNDA.n7241 585
R8432 GNDA.n7241 GNDA.n7240 585
R8433 GNDA.n7444 GNDA.n7443 585
R8434 GNDA.n7445 GNDA.n7444 585
R8435 GNDA.n88 GNDA.n87 585
R8436 GNDA.n7446 GNDA.n88 585
R8437 GNDA.n7449 GNDA.n7448 585
R8438 GNDA.n7448 GNDA.n7447 585
R8439 GNDA.n7451 GNDA.n85 585
R8440 GNDA.n85 GNDA.n84 585
R8441 GNDA.n7453 GNDA.n7452 585
R8442 GNDA.n7454 GNDA.n7453 585
R8443 GNDA.n83 GNDA.n82 585
R8444 GNDA.n7455 GNDA.n83 585
R8445 GNDA.n7458 GNDA.n7457 585
R8446 GNDA.n7457 GNDA.n7456 585
R8447 GNDA.n7459 GNDA.n80 585
R8448 GNDA.n80 GNDA.n78 585
R8449 GNDA.n7461 GNDA.n7460 585
R8450 GNDA.n7462 GNDA.n7461 585
R8451 GNDA.n7268 GNDA.n59 585
R8452 GNDA.n7271 GNDA.n7270 585
R8453 GNDA.n7276 GNDA.n7267 585
R8454 GNDA.n7277 GNDA.n7265 585
R8455 GNDA.n7278 GNDA.n7264 585
R8456 GNDA.n7262 GNDA.n7260 585
R8457 GNDA.n7284 GNDA.n7259 585
R8458 GNDA.n7285 GNDA.n7257 585
R8459 GNDA.n7286 GNDA.n7256 585
R8460 GNDA.n7254 GNDA.n7252 585
R8461 GNDA.n7292 GNDA.n7251 585
R8462 GNDA.n7293 GNDA.n7249 585
R8463 GNDA.n7475 GNDA.n60 585
R8464 GNDA.n7473 GNDA.n60 585
R8465 GNDA.n7293 GNDA.n7247 585
R8466 GNDA.n7292 GNDA.n7291 585
R8467 GNDA.n7289 GNDA.n7252 585
R8468 GNDA.n7287 GNDA.n7286 585
R8469 GNDA.n7285 GNDA.n7253 585
R8470 GNDA.n7284 GNDA.n7283 585
R8471 GNDA.n7281 GNDA.n7260 585
R8472 GNDA.n7279 GNDA.n7278 585
R8473 GNDA.n7277 GNDA.n7261 585
R8474 GNDA.n7276 GNDA.n7275 585
R8475 GNDA.n7273 GNDA.n7271 585
R8476 GNDA.n62 GNDA.n59 585
R8477 GNDA.n7475 GNDA.n7474 585
R8478 GNDA.n7474 GNDA.n7473 585
R8479 GNDA.n5601 GNDA.n5600 585
R8480 GNDA.n5602 GNDA.n5598 585
R8481 GNDA.n5605 GNDA.n5597 585
R8482 GNDA.n5606 GNDA.n5595 585
R8483 GNDA.n5609 GNDA.n5594 585
R8484 GNDA.n5610 GNDA.n5592 585
R8485 GNDA.n5613 GNDA.n5591 585
R8486 GNDA.n5614 GNDA.n5589 585
R8487 GNDA.n5615 GNDA.n5588 585
R8488 GNDA.n5580 GNDA.n5579 585
R8489 GNDA.n5807 GNDA.n5806 585
R8490 GNDA.n5809 GNDA.n5577 585
R8491 GNDA.n6072 GNDA.n5443 585
R8492 GNDA.n6070 GNDA.n5443 585
R8493 GNDA.n5803 GNDA.n5577 585
R8494 GNDA.n5806 GNDA.n5805 585
R8495 GNDA.n5581 GNDA.n5580 585
R8496 GNDA.n5616 GNDA.n5615 585
R8497 GNDA.n5614 GNDA.n5586 585
R8498 GNDA.n5613 GNDA.n5612 585
R8499 GNDA.n5611 GNDA.n5610 585
R8500 GNDA.n5609 GNDA.n5608 585
R8501 GNDA.n5607 GNDA.n5606 585
R8502 GNDA.n5605 GNDA.n5604 585
R8503 GNDA.n5603 GNDA.n5602 585
R8504 GNDA.n5601 GNDA.n5444 585
R8505 GNDA.n6072 GNDA.n6071 585
R8506 GNDA.n6071 GNDA.n6070 585
R8507 GNDA.n6924 GNDA.n5370 585
R8508 GNDA.n6927 GNDA.n6926 585
R8509 GNDA.n5375 GNDA.n5374 585
R8510 GNDA.n6131 GNDA.n6130 585
R8511 GNDA.n6136 GNDA.n6129 585
R8512 GNDA.n6137 GNDA.n6128 585
R8513 GNDA.n6138 GNDA.n6127 585
R8514 GNDA.n6125 GNDA.n6124 585
R8515 GNDA.n6143 GNDA.n6123 585
R8516 GNDA.n6144 GNDA.n6122 585
R8517 GNDA.n6121 GNDA.n6074 585
R8518 GNDA.n6150 GNDA.n6149 585
R8519 GNDA.n6149 GNDA.n6148 585
R8520 GNDA.n6146 GNDA.n6074 585
R8521 GNDA.n6145 GNDA.n6144 585
R8522 GNDA.n6143 GNDA.n6142 585
R8523 GNDA.n6141 GNDA.n6125 585
R8524 GNDA.n6139 GNDA.n6138 585
R8525 GNDA.n6137 GNDA.n6126 585
R8526 GNDA.n6136 GNDA.n6135 585
R8527 GNDA.n6133 GNDA.n6131 585
R8528 GNDA.n5374 GNDA.n5373 585
R8529 GNDA.n6928 GNDA.n6927 585
R8530 GNDA.n6930 GNDA.n5370 585
R8531 GNDA.n6952 GNDA.n5350 585
R8532 GNDA.n5352 GNDA.n5349 585
R8533 GNDA.n6955 GNDA.n5349 585
R8534 GNDA.n5361 GNDA.n5360 585
R8535 GNDA.n6941 GNDA.n6940 585
R8536 GNDA.n6940 GNDA.n6939 585
R8537 GNDA.n6783 GNDA.n6651 585
R8538 GNDA.n6790 GNDA.n6650 585
R8539 GNDA.n6794 GNDA.n6650 585
R8540 GNDA.n6788 GNDA.n6787 585
R8541 GNDA.n6770 GNDA.n6665 585
R8542 GNDA.n6773 GNDA.n6772 585
R8543 GNDA.n6774 GNDA.n6773 585
R8544 GNDA.n6765 GNDA.n6764 585
R8545 GNDA.n6913 GNDA.n5387 585
R8546 GNDA.n6913 GNDA.n6912 585
R8547 GNDA.n6823 GNDA.n6822 585
R8548 GNDA.n6824 GNDA.n6823 585
R8549 GNDA.n6820 GNDA.n5404 585
R8550 GNDA.n5404 GNDA.n5402 585
R8551 GNDA.n6642 GNDA.n6576 585
R8552 GNDA.n6646 GNDA.n6642 585
R8553 GNDA.n6815 GNDA.n6814 585
R8554 GNDA.n6814 GNDA.n6813 585
R8555 GNDA.n6797 GNDA.n6643 585
R8556 GNDA.n6812 GNDA.n6643 585
R8557 GNDA.n6810 GNDA.n6809 585
R8558 GNDA.n6811 GNDA.n6810 585
R8559 GNDA.n6800 GNDA.n6796 585
R8560 GNDA.n6796 GNDA.n6795 585
R8561 GNDA.n6801 GNDA.n5400 585
R8562 GNDA.n5401 GNDA.n5400 585
R8563 GNDA.n6828 GNDA.n6827 585
R8564 GNDA.n6827 GNDA.n6826 585
R8565 GNDA.n6829 GNDA.n5394 585
R8566 GNDA.n6825 GNDA.n5394 585
R8567 GNDA.n6909 GNDA.n6908 585
R8568 GNDA.n6910 GNDA.n6909 585
R8569 GNDA.n6906 GNDA.n5393 585
R8570 GNDA.n6911 GNDA.n5393 585
R8571 GNDA.n6932 GNDA.n5367 585
R8572 GNDA.n5382 GNDA.n5367 585
R8573 GNDA.n6921 GNDA.n5387 585
R8574 GNDA.n6922 GNDA.n6921 585
R8575 GNDA.n6904 GNDA.n5388 585
R8576 GNDA.n5388 GNDA.n5348 585
R8577 GNDA.n5346 GNDA.n5344 585
R8578 GNDA.n6958 GNDA.n5346 585
R8579 GNDA.n6973 GNDA.n6972 585
R8580 GNDA.n6972 GNDA.n6971 585
R8581 GNDA.n6960 GNDA.n5347 585
R8582 GNDA.n6970 GNDA.n5347 585
R8583 GNDA.n6968 GNDA.n6967 585
R8584 GNDA.n6969 GNDA.n6968 585
R8585 GNDA.n6963 GNDA.n5321 585
R8586 GNDA.n6959 GNDA.n5321 585
R8587 GNDA.n6981 GNDA.n6980 585
R8588 GNDA.n6982 GNDA.n6981 585
R8589 GNDA.n5323 GNDA.n5322 585
R8590 GNDA.n6841 GNDA.n5322 585
R8591 GNDA.n6840 GNDA.n6839 585
R8592 GNDA.n6842 GNDA.n6840 585
R8593 GNDA.n6846 GNDA.n6845 585
R8594 GNDA.n6845 GNDA.n6844 585
R8595 GNDA.n6847 GNDA.n5366 585
R8596 GNDA.n6843 GNDA.n5366 585
R8597 GNDA.n6935 GNDA.n6934 585
R8598 GNDA.n6936 GNDA.n6935 585
R8599 GNDA.n6932 GNDA.n6931 585
R8600 GNDA.n6931 GNDA.n5371 585
R8601 GNDA.n5372 GNDA.n5369 585
R8602 GNDA.n6742 GNDA.n5372 585
R8603 GNDA.n6744 GNDA.n6741 585
R8604 GNDA.n6744 GNDA.n6743 585
R8605 GNDA.n6745 GNDA.n6670 585
R8606 GNDA.n6746 GNDA.n6745 585
R8607 GNDA.n6750 GNDA.n6749 585
R8608 GNDA.n6749 GNDA.n6748 585
R8609 GNDA.n6667 GNDA.n6666 585
R8610 GNDA.n6747 GNDA.n6666 585
R8611 GNDA.n6761 GNDA.n6760 585
R8612 GNDA.n6762 GNDA.n6761 585
R8613 GNDA.n6758 GNDA.n296 585
R8614 GNDA.n7017 GNDA.n296 585
R8615 GNDA.n7020 GNDA.n7019 585
R8616 GNDA.n7019 GNDA.n7018 585
R8617 GNDA.n293 GNDA.n288 585
R8618 GNDA.n288 GNDA.n286 585
R8619 GNDA.n7030 GNDA.n7029 585
R8620 GNDA.n7031 GNDA.n7030 585
R8621 GNDA.n291 GNDA.n289 585
R8622 GNDA.n289 GNDA.n287 585
R8623 GNDA.n308 GNDA.n307 585
R8624 GNDA.n309 GNDA.n308 585
R8625 GNDA.n7000 GNDA.n6999 585
R8626 GNDA.n7001 GNDA.n7000 585
R8627 GNDA.n6997 GNDA.n6996 585
R8628 GNDA.n6996 GNDA.n6995 585
R8629 GNDA.n306 GNDA.n305 585
R8630 GNDA.n7007 GNDA.n7006 585
R8631 GNDA.n7008 GNDA.n7007 585
R8632 GNDA.n304 GNDA.n303 585
R8633 GNDA.n7009 GNDA.n304 585
R8634 GNDA.n7012 GNDA.n7011 585
R8635 GNDA.n7011 GNDA.n7010 585
R8636 GNDA.n7013 GNDA.n301 585
R8637 GNDA.n301 GNDA.n299 585
R8638 GNDA.n7015 GNDA.n7014 585
R8639 GNDA.n7016 GNDA.n7015 585
R8640 GNDA.n302 GNDA.n300 585
R8641 GNDA.n300 GNDA.n298 585
R8642 GNDA.n6091 GNDA.n6090 585
R8643 GNDA.n6090 GNDA.n6089 585
R8644 GNDA.n6092 GNDA.n6087 585
R8645 GNDA.n6087 GNDA.n6086 585
R8646 GNDA.n6094 GNDA.n6093 585
R8647 GNDA.n6095 GNDA.n6094 585
R8648 GNDA.n6088 GNDA.n6085 585
R8649 GNDA.n6096 GNDA.n6085 585
R8650 GNDA.n6098 GNDA.n6083 585
R8651 GNDA.n6098 GNDA.n6097 585
R8652 GNDA.n7003 GNDA.n7002 585
R8653 GNDA.n5759 GNDA.n5640 585
R8654 GNDA.n5762 GNDA.n5761 585
R8655 GNDA.n5761 GNDA.n5760 585
R8656 GNDA.n5763 GNDA.n5637 585
R8657 GNDA.n5637 GNDA.n5636 585
R8658 GNDA.n5765 GNDA.n5764 585
R8659 GNDA.n5766 GNDA.n5765 585
R8660 GNDA.n5638 GNDA.n5634 585
R8661 GNDA.n5767 GNDA.n5634 585
R8662 GNDA.n5769 GNDA.n5635 585
R8663 GNDA.n5769 GNDA.n5768 585
R8664 GNDA.n5770 GNDA.n5633 585
R8665 GNDA.n5771 GNDA.n5770 585
R8666 GNDA.n5774 GNDA.n5773 585
R8667 GNDA.n5773 GNDA.n5772 585
R8668 GNDA.n5775 GNDA.n5631 585
R8669 GNDA.n5631 GNDA.n5630 585
R8670 GNDA.n5777 GNDA.n5776 585
R8671 GNDA.n5778 GNDA.n5777 585
R8672 GNDA.n5632 GNDA.n5629 585
R8673 GNDA.n5779 GNDA.n5629 585
R8674 GNDA.n5781 GNDA.n5627 585
R8675 GNDA.n5781 GNDA.n5780 585
R8676 GNDA.n5758 GNDA.n5757 585
R8677 GNDA.n7389 GNDA.n7316 585
R8678 GNDA.n7392 GNDA.n7391 585
R8679 GNDA.n7391 GNDA.n7390 585
R8680 GNDA.n7393 GNDA.n7314 585
R8681 GNDA.n7314 GNDA.n7313 585
R8682 GNDA.n7395 GNDA.n7394 585
R8683 GNDA.n7396 GNDA.n7395 585
R8684 GNDA.n7312 GNDA.n7311 585
R8685 GNDA.n7397 GNDA.n7312 585
R8686 GNDA.n7400 GNDA.n7399 585
R8687 GNDA.n7399 GNDA.n7398 585
R8688 GNDA.n7401 GNDA.n7310 585
R8689 GNDA.n7310 GNDA.n7309 585
R8690 GNDA.n7403 GNDA.n7402 585
R8691 GNDA.n7404 GNDA.n7403 585
R8692 GNDA.n7308 GNDA.n7307 585
R8693 GNDA.n7405 GNDA.n7308 585
R8694 GNDA.n7408 GNDA.n7407 585
R8695 GNDA.n7407 GNDA.n7406 585
R8696 GNDA.n7409 GNDA.n7306 585
R8697 GNDA.n7306 GNDA.n7305 585
R8698 GNDA.n7411 GNDA.n7410 585
R8699 GNDA.n7412 GNDA.n7411 585
R8700 GNDA.n7388 GNDA.n7387 585
R8701 GNDA.n6253 GNDA.n6252 585
R8702 GNDA.n6251 GNDA.n5426 585
R8703 GNDA.n6250 GNDA.n6249 585
R8704 GNDA.n6248 GNDA.n6247 585
R8705 GNDA.n6246 GNDA.n6245 585
R8706 GNDA.n6244 GNDA.n6243 585
R8707 GNDA.n6242 GNDA.n6241 585
R8708 GNDA.n6240 GNDA.n6239 585
R8709 GNDA.n6238 GNDA.n6237 585
R8710 GNDA.n6236 GNDA.n6235 585
R8711 GNDA.n5406 GNDA.n5405 585
R8712 GNDA.n6571 GNDA.n5406 585
R8713 GNDA.n6574 GNDA.n6573 585
R8714 GNDA.n6574 GNDA.n5403 585
R8715 GNDA.n5860 GNDA.n5859 585
R8716 GNDA.n5862 GNDA.n5861 585
R8717 GNDA.n5864 GNDA.n5863 585
R8718 GNDA.n5866 GNDA.n5865 585
R8719 GNDA.n5868 GNDA.n5867 585
R8720 GNDA.n5870 GNDA.n5869 585
R8721 GNDA.n5872 GNDA.n5871 585
R8722 GNDA.n5874 GNDA.n5873 585
R8723 GNDA.n5876 GNDA.n5875 585
R8724 GNDA.n5878 GNDA.n5877 585
R8725 GNDA.n5880 GNDA.n5879 585
R8726 GNDA.n6571 GNDA.n5421 585
R8727 GNDA.n6569 GNDA.n6568 585
R8728 GNDA.n6567 GNDA.n6256 585
R8729 GNDA.n6566 GNDA.n6255 585
R8730 GNDA.n6571 GNDA.n6255 585
R8731 GNDA.n6565 GNDA.n6564 585
R8732 GNDA.n6563 GNDA.n6562 585
R8733 GNDA.n6561 GNDA.n6560 585
R8734 GNDA.n6559 GNDA.n6558 585
R8735 GNDA.n6557 GNDA.n6556 585
R8736 GNDA.n6555 GNDA.n6554 585
R8737 GNDA.n6553 GNDA.n6552 585
R8738 GNDA.n6551 GNDA.n6550 585
R8739 GNDA.n6549 GNDA.n6548 585
R8740 GNDA.n6548 GNDA.n6547 585
R8741 GNDA.n1752 GNDA.n1751 577.346
R8742 GNDA.n6991 GNDA.n313 568.266
R8743 GNDA.n2108 GNDA.t201 524.808
R8744 GNDA.n4999 GNDA.t213 524.808
R8745 GNDA.n5004 GNDA.t228 524.808
R8746 GNDA.n659 GNDA.t189 524.808
R8747 GNDA.n1733 GNDA.t164 508.743
R8748 GNDA.n1741 GNDA.t161 508.743
R8749 GNDA.n3391 GNDA.t210 508.743
R8750 GNDA.n3381 GNDA.t183 508.743
R8751 GNDA.n3397 GNDA.t234 499.442
R8752 GNDA.n5308 GNDA.t222 499.442
R8753 GNDA.n1755 GNDA.t175 499.442
R8754 GNDA.n1744 GNDA.t168 499.442
R8755 GNDA.n3385 GNDA.t216 475.976
R8756 GNDA.n3385 GNDA.t198 475.976
R8757 GNDA.n1727 GNDA.t231 475.976
R8758 GNDA.n1727 GNDA.t207 475.976
R8759 GNDA.n5311 GNDA.n5310 471.68
R8760 GNDA.n3395 GNDA.n574 471.68
R8761 GNDA.n7002 GNDA.n7001 427.599
R8762 GNDA.n272 GNDA.t194 425.134
R8763 GNDA.n269 GNDA.t148 409.067
R8764 GNDA.n7034 GNDA.t243 409.067
R8765 GNDA.n282 GNDA.t178 409.067
R8766 GNDA.n281 GNDA.t141 409.067
R8767 GNDA.n278 GNDA.t186 409.067
R8768 GNDA.n277 GNDA.t154 409.067
R8769 GNDA.n273 GNDA.t246 409.067
R8770 GNDA.n7437 GNDA.n7245 370.214
R8771 GNDA.n7463 GNDA.n68 370.214
R8772 GNDA.n7437 GNDA.n7244 365.957
R8773 GNDA.n7464 GNDA.n7463 365.957
R8774 GNDA.n1747 GNDA.n1746 337.098
R8775 GNDA.n1753 GNDA.n1752 337.098
R8776 GNDA.n7244 GNDA.t145 327.661
R8777 GNDA.n7464 GNDA.t145 327.661
R8778 GNDA.n5381 GNDA.t145 172.876
R8779 GNDA.n6923 GNDA.t145 172.876
R8780 GNDA.n7245 GNDA.t145 323.404
R8781 GNDA.t145 GNDA.n68 323.404
R8782 GNDA.n5384 GNDA.t145 172.615
R8783 GNDA.t145 GNDA.n297 172.615
R8784 GNDA.n1736 GNDA.n1734 296.158
R8785 GNDA.n1740 GNDA.n1739 296.158
R8786 GNDA.n3393 GNDA.n3392 296.158
R8787 GNDA.n3383 GNDA.n3382 296.158
R8788 GNDA.n5310 GNDA.n5309 292.5
R8789 GNDA.n1732 GNDA.n1731 292.5
R8790 GNDA.n3390 GNDA.n3389 292.5
R8791 GNDA.n3396 GNDA.n3395 292.5
R8792 GNDA.n1746 GNDA.n1745 292.5
R8793 GNDA.n1754 GNDA.n1753 292.5
R8794 GNDA.n7005 GNDA.n7004 264.301
R8795 GNDA.n5756 GNDA.n5639 264.301
R8796 GNDA.n7386 GNDA.n7315 264.301
R8797 GNDA.n6572 GNDA.n6571 264.301
R8798 GNDA.n5882 GNDA.n5881 264.301
R8799 GNDA.n6571 GNDA.n5414 264.301
R8800 GNDA.n6999 GNDA.t1 260
R8801 GNDA.n6997 GNDA.t1 260
R8802 GNDA.n7411 GNDA.n7304 259.416
R8803 GNDA.n5782 GNDA.n5781 259.416
R8804 GNDA.n5810 GNDA.n5809 259.416
R8805 GNDA.n5838 GNDA.n5837 259.416
R8806 GNDA.n7249 GNDA.n7243 259.416
R8807 GNDA.n6300 GNDA.n6298 259.416
R8808 GNDA.n6212 GNDA.n5433 259.416
R8809 GNDA.n6099 GNDA.n6098 259.416
R8810 GNDA.n6152 GNDA.n6150 259.416
R8811 GNDA.n6519 GNDA.n6518 258.334
R8812 GNDA.n6424 GNDA.n6423 258.334
R8813 GNDA.n6886 GNDA.n6885 258.334
R8814 GNDA.n6623 GNDA.n6621 258.334
R8815 GNDA.n5699 GNDA.n5698 258.334
R8816 GNDA.n6041 GNDA.n6040 258.334
R8817 GNDA.n5965 GNDA.n5906 258.334
R8818 GNDA.n6721 GNDA.n6719 258.334
R8819 GNDA.n7335 GNDA.n7334 258.334
R8820 GNDA.n7466 GNDA.n7464 254.34
R8821 GNDA.n7464 GNDA.n76 254.34
R8822 GNDA.n7464 GNDA.n75 254.34
R8823 GNDA.n7464 GNDA.n74 254.34
R8824 GNDA.n7464 GNDA.n73 254.34
R8825 GNDA.n7464 GNDA.n72 254.34
R8826 GNDA.n6294 GNDA.n68 254.34
R8827 GNDA.n6292 GNDA.n68 254.34
R8828 GNDA.n6286 GNDA.n68 254.34
R8829 GNDA.n6284 GNDA.n68 254.34
R8830 GNDA.n6277 GNDA.n68 254.34
R8831 GNDA.n7470 GNDA.n68 254.34
R8832 GNDA.n6084 GNDA.n5383 254.34
R8833 GNDA.n6104 GNDA.n5383 254.34
R8834 GNDA.n6081 GNDA.n5383 254.34
R8835 GNDA.n6111 GNDA.n5383 254.34
R8836 GNDA.n6078 GNDA.n5383 254.34
R8837 GNDA.n6118 GNDA.n5383 254.34
R8838 GNDA.n5999 GNDA.n5998 254.34
R8839 GNDA.n5999 GNDA.n5513 254.34
R8840 GNDA.n5999 GNDA.n5512 254.34
R8841 GNDA.n5999 GNDA.n5511 254.34
R8842 GNDA.n5999 GNDA.n5510 254.34
R8843 GNDA.n5999 GNDA.n5509 254.34
R8844 GNDA.n5999 GNDA.n5449 254.34
R8845 GNDA.n5999 GNDA.n5453 254.34
R8846 GNDA.n5999 GNDA.n5508 254.34
R8847 GNDA.n5999 GNDA.n5485 254.34
R8848 GNDA.n5999 GNDA.n5484 254.34
R8849 GNDA.n6000 GNDA.n5999 254.34
R8850 GNDA.n5999 GNDA.n5483 254.34
R8851 GNDA.n5999 GNDA.n5482 254.34
R8852 GNDA.n5999 GNDA.n5481 254.34
R8853 GNDA.n5999 GNDA.n5480 254.34
R8854 GNDA.n5999 GNDA.n5479 254.34
R8855 GNDA.n5999 GNDA.n5478 254.34
R8856 GNDA.n6151 GNDA.n5383 254.34
R8857 GNDA.n6157 GNDA.n5383 254.34
R8858 GNDA.n6159 GNDA.n5383 254.34
R8859 GNDA.n6165 GNDA.n5383 254.34
R8860 GNDA.n6167 GNDA.n5383 254.34
R8861 GNDA.n6173 GNDA.n5383 254.34
R8862 GNDA.n6213 GNDA.n5383 254.34
R8863 GNDA.n6215 GNDA.n5383 254.34
R8864 GNDA.n6221 GNDA.n5383 254.34
R8865 GNDA.n6223 GNDA.n5383 254.34
R8866 GNDA.n6229 GNDA.n5383 254.34
R8867 GNDA.n6231 GNDA.n5383 254.34
R8868 GNDA.n6915 GNDA.n5381 254.34
R8869 GNDA.n6189 GNDA.n5381 254.34
R8870 GNDA.n6187 GNDA.n5381 254.34
R8871 GNDA.n6184 GNDA.n5381 254.34
R8872 GNDA.n6179 GNDA.n5381 254.34
R8873 GNDA.n6176 GNDA.n5381 254.34
R8874 GNDA.n6207 GNDA.n5384 254.34
R8875 GNDA.n6175 GNDA.n5384 254.34
R8876 GNDA.n6200 GNDA.n5384 254.34
R8877 GNDA.n6194 GNDA.n5384 254.34
R8878 GNDA.n6192 GNDA.n5384 254.34
R8879 GNDA.n6919 GNDA.n5384 254.34
R8880 GNDA.n5548 GNDA.n5527 254.34
R8881 GNDA.n5545 GNDA.n5527 254.34
R8882 GNDA.n5542 GNDA.n5527 254.34
R8883 GNDA.n5539 GNDA.n5527 254.34
R8884 GNDA.n5536 GNDA.n5527 254.34
R8885 GNDA.n5836 GNDA.n5527 254.34
R8886 GNDA.n5832 GNDA.n5567 254.34
R8887 GNDA.n5567 GNDA.n5566 254.34
R8888 GNDA.n5567 GNDA.n5534 254.34
R8889 GNDA.n5567 GNDA.n5533 254.34
R8890 GNDA.n5567 GNDA.n5532 254.34
R8891 GNDA.n5567 GNDA.n5531 254.34
R8892 GNDA.n5525 GNDA.n5516 254.34
R8893 GNDA.n5843 GNDA.n5516 254.34
R8894 GNDA.n5522 GNDA.n5516 254.34
R8895 GNDA.n5850 GNDA.n5516 254.34
R8896 GNDA.n5519 GNDA.n5516 254.34
R8897 GNDA.n5857 GNDA.n5516 254.34
R8898 GNDA.n5576 GNDA.n5516 254.34
R8899 GNDA.n5815 GNDA.n5516 254.34
R8900 GNDA.n5574 GNDA.n5516 254.34
R8901 GNDA.n5822 GNDA.n5516 254.34
R8902 GNDA.n5571 GNDA.n5516 254.34
R8903 GNDA.n5829 GNDA.n5516 254.34
R8904 GNDA.n5628 GNDA.n5516 254.34
R8905 GNDA.n5787 GNDA.n5516 254.34
R8906 GNDA.n5625 GNDA.n5516 254.34
R8907 GNDA.n5794 GNDA.n5516 254.34
R8908 GNDA.n5622 GNDA.n5516 254.34
R8909 GNDA.n5801 GNDA.n5516 254.34
R8910 GNDA.n7482 GNDA.n43 254.34
R8911 GNDA.n7482 GNDA.n44 254.34
R8912 GNDA.n7482 GNDA.n45 254.34
R8913 GNDA.n7482 GNDA.n46 254.34
R8914 GNDA.n7482 GNDA.n47 254.34
R8915 GNDA.n7482 GNDA.n48 254.34
R8916 GNDA.n7482 GNDA.n49 254.34
R8917 GNDA.n7482 GNDA.n50 254.34
R8918 GNDA.n7482 GNDA.n51 254.34
R8919 GNDA.n7482 GNDA.n52 254.34
R8920 GNDA.n7482 GNDA.n53 254.34
R8921 GNDA.n7482 GNDA.n7481 254.34
R8922 GNDA.n7482 GNDA.n42 254.34
R8923 GNDA.n7483 GNDA.n7482 254.34
R8924 GNDA.n7482 GNDA.n41 254.34
R8925 GNDA.n7482 GNDA.n29 254.34
R8926 GNDA.n7482 GNDA.n28 254.34
R8927 GNDA.n7482 GNDA.n27 254.34
R8928 GNDA.n7269 GNDA.n7244 254.34
R8929 GNDA.n7266 GNDA.n7244 254.34
R8930 GNDA.n7263 GNDA.n7244 254.34
R8931 GNDA.n7258 GNDA.n7244 254.34
R8932 GNDA.n7255 GNDA.n7244 254.34
R8933 GNDA.n7250 GNDA.n7244 254.34
R8934 GNDA.n7290 GNDA.n7245 254.34
R8935 GNDA.n7288 GNDA.n7245 254.34
R8936 GNDA.n7282 GNDA.n7245 254.34
R8937 GNDA.n7280 GNDA.n7245 254.34
R8938 GNDA.n7274 GNDA.n7245 254.34
R8939 GNDA.n7272 GNDA.n7245 254.34
R8940 GNDA.n5599 GNDA.n5578 254.34
R8941 GNDA.n5596 GNDA.n5578 254.34
R8942 GNDA.n5593 GNDA.n5578 254.34
R8943 GNDA.n5590 GNDA.n5578 254.34
R8944 GNDA.n5587 GNDA.n5578 254.34
R8945 GNDA.n5808 GNDA.n5578 254.34
R8946 GNDA.n5804 GNDA.n5618 254.34
R8947 GNDA.n5618 GNDA.n5617 254.34
R8948 GNDA.n5618 GNDA.n5585 254.34
R8949 GNDA.n5618 GNDA.n5584 254.34
R8950 GNDA.n5618 GNDA.n5583 254.34
R8951 GNDA.n5618 GNDA.n5582 254.34
R8952 GNDA.n6925 GNDA.n6923 254.34
R8953 GNDA.n6923 GNDA.n5380 254.34
R8954 GNDA.n6923 GNDA.n5379 254.34
R8955 GNDA.n6923 GNDA.n5378 254.34
R8956 GNDA.n6923 GNDA.n5377 254.34
R8957 GNDA.n6923 GNDA.n5376 254.34
R8958 GNDA.n6147 GNDA.n297 254.34
R8959 GNDA.n6120 GNDA.n297 254.34
R8960 GNDA.n6140 GNDA.n297 254.34
R8961 GNDA.n6134 GNDA.n297 254.34
R8962 GNDA.n6132 GNDA.n297 254.34
R8963 GNDA.n6929 GNDA.n297 254.34
R8964 GNDA.n6571 GNDA.n6254 254.34
R8965 GNDA.n6571 GNDA.n5425 254.34
R8966 GNDA.n6571 GNDA.n5424 254.34
R8967 GNDA.n6571 GNDA.n5423 254.34
R8968 GNDA.n6571 GNDA.n5422 254.34
R8969 GNDA.n6571 GNDA.n5415 254.34
R8970 GNDA.n6571 GNDA.n5416 254.34
R8971 GNDA.n6571 GNDA.n5417 254.34
R8972 GNDA.n6571 GNDA.n5418 254.34
R8973 GNDA.n6571 GNDA.n5419 254.34
R8974 GNDA.n6571 GNDA.n5420 254.34
R8975 GNDA.n6571 GNDA.n6570 254.34
R8976 GNDA.n6571 GNDA.n5410 254.34
R8977 GNDA.n6571 GNDA.n5411 254.34
R8978 GNDA.n6571 GNDA.n5412 254.34
R8979 GNDA.n6571 GNDA.n5413 254.34
R8980 GNDA.t145 GNDA.n7239 250.349
R8981 GNDA.n6955 GNDA.n6954 250.349
R8982 GNDA.n6939 GNDA.n6938 250.349
R8983 GNDA.n7435 GNDA.n7247 249.663
R8984 GNDA.n5803 GNDA.n5802 249.663
R8985 GNDA.n5831 GNDA.n5830 249.663
R8986 GNDA.n5859 GNDA.n5858 249.663
R8987 GNDA.n7461 GNDA.n79 249.663
R8988 GNDA.n6569 GNDA.n6257 249.663
R8989 GNDA.n6253 GNDA.n5427 249.663
R8990 GNDA.n6148 GNDA.n6119 249.663
R8991 GNDA.n6208 GNDA.n6174 249.663
R8992 GNDA.n7000 GNDA.n6996 246.25
R8993 GNDA.n6773 GNDA.n6665 246.25
R8994 GNDA.n6773 GNDA.n6764 246.25
R8995 GNDA.n6651 GNDA.n6650 246.25
R8996 GNDA.n6787 GNDA.n6650 246.25
R8997 GNDA.n6794 GNDA.n6793 241.643
R8998 GNDA.n6794 GNDA.n6649 241.643
R8999 GNDA.n6775 GNDA.n6774 241.643
R9000 GNDA.n6774 GNDA.n6763 241.643
R9001 GNDA.n1746 GNDA.t169 239.517
R9002 GNDA.n1739 GNDA.t162 239.517
R9003 GNDA.n1739 GNDA.t159 239.517
R9004 GNDA.t238 GNDA.n1736 239.517
R9005 GNDA.n1736 GNDA.t165 239.517
R9006 GNDA.n1753 GNDA.t176 239.517
R9007 GNDA.n1736 GNDA.n1735 197.133
R9008 GNDA.n1739 GNDA.n1738 197.133
R9009 GNDA.n5307 GNDA.n5306 197.133
R9010 GNDA.n3394 GNDA.n321 197.133
R9011 GNDA.n6940 GNDA.n5361 197
R9012 GNDA.n5350 GNDA.n5349 197
R9013 GNDA.n60 GNDA.n54 197
R9014 GNDA.n7238 GNDA.n89 197
R9015 GNDA.n6452 GNDA.n64 197
R9016 GNDA.n6913 GNDA.n5393 197
R9017 GNDA.n5757 GNDA.n5755 197
R9018 GNDA.n5477 GNDA.n5443 197
R9019 GNDA.n5908 GNDA.n5447 197
R9020 GNDA.n7003 GNDA.n308 197
R9021 GNDA.n6935 GNDA.n5367 197
R9022 GNDA.n7387 GNDA.n7385 197
R9023 GNDA.t303 GNDA.t169 195.161
R9024 GNDA.t82 GNDA.t303 195.161
R9025 GNDA.t42 GNDA.t82 195.161
R9026 GNDA.t309 GNDA.t42 195.161
R9027 GNDA.t64 GNDA.t309 195.161
R9028 GNDA.t88 GNDA.t64 195.161
R9029 GNDA.t69 GNDA.t88 195.161
R9030 GNDA.t130 GNDA.t69 195.161
R9031 GNDA.t57 GNDA.t130 195.161
R9032 GNDA.t336 GNDA.t57 195.161
R9033 GNDA.t162 GNDA.t336 195.161
R9034 GNDA.t159 GNDA.t11 195.161
R9035 GNDA.t299 GNDA.t238 195.161
R9036 GNDA.t165 GNDA.t321 195.161
R9037 GNDA.t321 GNDA.t89 195.161
R9038 GNDA.t89 GNDA.t98 195.161
R9039 GNDA.t98 GNDA.t22 195.161
R9040 GNDA.t22 GNDA.t333 195.161
R9041 GNDA.t333 GNDA.t87 195.161
R9042 GNDA.t87 GNDA.t76 195.161
R9043 GNDA.t76 GNDA.t326 195.161
R9044 GNDA.t326 GNDA.t51 195.161
R9045 GNDA.t51 GNDA.t83 195.161
R9046 GNDA.t83 GNDA.t176 195.161
R9047 GNDA.t137 GNDA.t195 187.597
R9048 GNDA.n7472 GNDA.n66 187.249
R9049 GNDA.n6547 GNDA.n6546 187.249
R9050 GNDA.n6823 GNDA.n5403 187.249
R9051 GNDA.n6071 GNDA.n5445 187.249
R9052 GNDA.n6069 GNDA.n6068 187.249
R9053 GNDA.n5997 GNDA.n5421 187.249
R9054 GNDA.n6931 GNDA.n5372 187.249
R9055 GNDA.n6921 GNDA.n5388 187.249
R9056 GNDA.n7474 GNDA.n63 187.249
R9057 GNDA.n6776 GNDA.n6664 185
R9058 GNDA.n6768 GNDA.n6767 185
R9059 GNDA.n6792 GNDA.n6791 185
R9060 GNDA.n6791 GNDA.n6790 185
R9061 GNDA.n6792 GNDA.n6782 185
R9062 GNDA.n6785 GNDA.n6782 185
R9063 GNDA.n6520 GNDA.n6519 185
R9064 GNDA.n6522 GNDA.n6521 185
R9065 GNDA.n6524 GNDA.n6523 185
R9066 GNDA.n6526 GNDA.n6525 185
R9067 GNDA.n6528 GNDA.n6527 185
R9068 GNDA.n6530 GNDA.n6529 185
R9069 GNDA.n6532 GNDA.n6531 185
R9070 GNDA.n6534 GNDA.n6533 185
R9071 GNDA.n6535 GNDA.n6323 185
R9072 GNDA.n6502 GNDA.n6501 185
R9073 GNDA.n6504 GNDA.n6503 185
R9074 GNDA.n6506 GNDA.n6505 185
R9075 GNDA.n6508 GNDA.n6507 185
R9076 GNDA.n6510 GNDA.n6509 185
R9077 GNDA.n6512 GNDA.n6511 185
R9078 GNDA.n6514 GNDA.n6513 185
R9079 GNDA.n6516 GNDA.n6515 185
R9080 GNDA.n6518 GNDA.n6517 185
R9081 GNDA.n6484 GNDA.n6483 185
R9082 GNDA.n6486 GNDA.n6485 185
R9083 GNDA.n6488 GNDA.n6487 185
R9084 GNDA.n6490 GNDA.n6489 185
R9085 GNDA.n6492 GNDA.n6491 185
R9086 GNDA.n6494 GNDA.n6493 185
R9087 GNDA.n6496 GNDA.n6495 185
R9088 GNDA.n6498 GNDA.n6497 185
R9089 GNDA.n6500 GNDA.n6499 185
R9090 GNDA.n6425 GNDA.n6424 185
R9091 GNDA.n6427 GNDA.n6426 185
R9092 GNDA.n6429 GNDA.n6428 185
R9093 GNDA.n6431 GNDA.n6430 185
R9094 GNDA.n6433 GNDA.n6432 185
R9095 GNDA.n6435 GNDA.n6434 185
R9096 GNDA.n6437 GNDA.n6436 185
R9097 GNDA.n6439 GNDA.n6438 185
R9098 GNDA.n6440 GNDA.n6344 185
R9099 GNDA.n6407 GNDA.n6406 185
R9100 GNDA.n6409 GNDA.n6408 185
R9101 GNDA.n6411 GNDA.n6410 185
R9102 GNDA.n6413 GNDA.n6412 185
R9103 GNDA.n6415 GNDA.n6414 185
R9104 GNDA.n6417 GNDA.n6416 185
R9105 GNDA.n6419 GNDA.n6418 185
R9106 GNDA.n6421 GNDA.n6420 185
R9107 GNDA.n6423 GNDA.n6422 185
R9108 GNDA.n6382 GNDA.n57 185
R9109 GNDA.n6391 GNDA.n6390 185
R9110 GNDA.n6393 GNDA.n6392 185
R9111 GNDA.n6395 GNDA.n6394 185
R9112 GNDA.n6397 GNDA.n6396 185
R9113 GNDA.n6399 GNDA.n6398 185
R9114 GNDA.n6401 GNDA.n6400 185
R9115 GNDA.n6403 GNDA.n6402 185
R9116 GNDA.n6405 GNDA.n6404 185
R9117 GNDA.n6381 GNDA.n56 185
R9118 GNDA.n6375 GNDA.n6374 185
R9119 GNDA.n6354 GNDA.n6353 185
R9120 GNDA.n6368 GNDA.n6367 185
R9121 GNDA.n6366 GNDA.n6365 185
R9122 GNDA.n6360 GNDA.n6359 185
R9123 GNDA.n6355 GNDA.n6348 185
R9124 GNDA.n6444 GNDA.n6443 185
R9125 GNDA.n6347 GNDA.n6345 185
R9126 GNDA.n6482 GNDA.n6481 185
R9127 GNDA.n6476 GNDA.n6475 185
R9128 GNDA.n6474 GNDA.n6473 185
R9129 GNDA.n6469 GNDA.n6468 185
R9130 GNDA.n6467 GNDA.n6466 185
R9131 GNDA.n6461 GNDA.n6460 185
R9132 GNDA.n6456 GNDA.n6327 185
R9133 GNDA.n6539 GNDA.n6538 185
R9134 GNDA.n6326 GNDA.n6324 185
R9135 GNDA.n6887 GNDA.n6886 185
R9136 GNDA.n6889 GNDA.n6888 185
R9137 GNDA.n6891 GNDA.n6890 185
R9138 GNDA.n6893 GNDA.n6892 185
R9139 GNDA.n6895 GNDA.n6894 185
R9140 GNDA.n6897 GNDA.n6896 185
R9141 GNDA.n6899 GNDA.n6898 185
R9142 GNDA.n6901 GNDA.n6900 185
R9143 GNDA.n6902 GNDA.n5342 185
R9144 GNDA.n6869 GNDA.n6868 185
R9145 GNDA.n6871 GNDA.n6870 185
R9146 GNDA.n6873 GNDA.n6872 185
R9147 GNDA.n6875 GNDA.n6874 185
R9148 GNDA.n6877 GNDA.n6876 185
R9149 GNDA.n6879 GNDA.n6878 185
R9150 GNDA.n6881 GNDA.n6880 185
R9151 GNDA.n6883 GNDA.n6882 185
R9152 GNDA.n6885 GNDA.n6884 185
R9153 GNDA.n6851 GNDA.n6850 185
R9154 GNDA.n6853 GNDA.n6852 185
R9155 GNDA.n6855 GNDA.n6854 185
R9156 GNDA.n6857 GNDA.n6856 185
R9157 GNDA.n6859 GNDA.n6858 185
R9158 GNDA.n6861 GNDA.n6860 185
R9159 GNDA.n6863 GNDA.n6862 185
R9160 GNDA.n6865 GNDA.n6864 185
R9161 GNDA.n6867 GNDA.n6866 185
R9162 GNDA.n6849 GNDA.n6848 185
R9163 GNDA.n6837 GNDA.n6836 185
R9164 GNDA.n6838 GNDA.n5325 185
R9165 GNDA.n6979 GNDA.n6978 185
R9166 GNDA.n6962 GNDA.n5324 185
R9167 GNDA.n6966 GNDA.n6965 185
R9168 GNDA.n6964 GNDA.n6961 185
R9169 GNDA.n5345 GNDA.n5343 185
R9170 GNDA.n6975 GNDA.n6974 185
R9171 GNDA.n6624 GNDA.n6623 185
R9172 GNDA.n6625 GNDA.n6580 185
R9173 GNDA.n6627 GNDA.n6626 185
R9174 GNDA.n6629 GNDA.n6579 185
R9175 GNDA.n6632 GNDA.n6631 185
R9176 GNDA.n6633 GNDA.n6578 185
R9177 GNDA.n6635 GNDA.n6634 185
R9178 GNDA.n6637 GNDA.n6577 185
R9179 GNDA.n6638 GNDA.n6575 185
R9180 GNDA.n6605 GNDA.n6585 185
R9181 GNDA.n6608 GNDA.n6607 185
R9182 GNDA.n6609 GNDA.n6584 185
R9183 GNDA.n6611 GNDA.n6610 185
R9184 GNDA.n6613 GNDA.n6583 185
R9185 GNDA.n6616 GNDA.n6615 185
R9186 GNDA.n6617 GNDA.n6582 185
R9187 GNDA.n6619 GNDA.n6618 185
R9188 GNDA.n6621 GNDA.n6581 185
R9189 GNDA.n6835 GNDA.n6834 185
R9190 GNDA.n6591 GNDA.n5396 185
R9191 GNDA.n6593 GNDA.n6592 185
R9192 GNDA.n6594 GNDA.n6589 185
R9193 GNDA.n6596 GNDA.n6595 185
R9194 GNDA.n6598 GNDA.n6587 185
R9195 GNDA.n6600 GNDA.n6599 185
R9196 GNDA.n6601 GNDA.n6586 185
R9197 GNDA.n6603 GNDA.n6602 185
R9198 GNDA.n6833 GNDA.n5395 185
R9199 GNDA.n6831 GNDA.n6830 185
R9200 GNDA.n5399 GNDA.n5398 185
R9201 GNDA.n6803 GNDA.n6802 185
R9202 GNDA.n6808 GNDA.n6807 185
R9203 GNDA.n6805 GNDA.n6798 185
R9204 GNDA.n6804 GNDA.n6641 185
R9205 GNDA.n6817 GNDA.n6816 185
R9206 GNDA.n6819 GNDA.n6818 185
R9207 GNDA.n5700 GNDA.n5699 185
R9208 GNDA.n5702 GNDA.n5701 185
R9209 GNDA.n5704 GNDA.n5703 185
R9210 GNDA.n5706 GNDA.n5705 185
R9211 GNDA.n5708 GNDA.n5707 185
R9212 GNDA.n5710 GNDA.n5709 185
R9213 GNDA.n5712 GNDA.n5711 185
R9214 GNDA.n5714 GNDA.n5713 185
R9215 GNDA.n5715 GNDA.n5663 185
R9216 GNDA.n5682 GNDA.n5681 185
R9217 GNDA.n5684 GNDA.n5683 185
R9218 GNDA.n5686 GNDA.n5685 185
R9219 GNDA.n5688 GNDA.n5687 185
R9220 GNDA.n5690 GNDA.n5689 185
R9221 GNDA.n5692 GNDA.n5691 185
R9222 GNDA.n5694 GNDA.n5693 185
R9223 GNDA.n5696 GNDA.n5695 185
R9224 GNDA.n5698 GNDA.n5697 185
R9225 GNDA.n5655 GNDA.n5641 185
R9226 GNDA.n5666 GNDA.n5665 185
R9227 GNDA.n5668 GNDA.n5667 185
R9228 GNDA.n5670 GNDA.n5669 185
R9229 GNDA.n5672 GNDA.n5671 185
R9230 GNDA.n5674 GNDA.n5673 185
R9231 GNDA.n5676 GNDA.n5675 185
R9232 GNDA.n5678 GNDA.n5677 185
R9233 GNDA.n5680 GNDA.n5679 185
R9234 GNDA.n5645 GNDA.n5642 185
R9235 GNDA.n5748 GNDA.n5747 185
R9236 GNDA.n5721 GNDA.n5644 185
R9237 GNDA.n5727 GNDA.n5726 185
R9238 GNDA.n5725 GNDA.n5720 185
R9239 GNDA.n5734 GNDA.n5733 185
R9240 GNDA.n5732 GNDA.n5719 185
R9241 GNDA.n5739 GNDA.n5664 185
R9242 GNDA.n5744 GNDA.n5743 185
R9243 GNDA.n6042 GNDA.n6041 185
R9244 GNDA.n6044 GNDA.n6043 185
R9245 GNDA.n6046 GNDA.n6045 185
R9246 GNDA.n6048 GNDA.n6047 185
R9247 GNDA.n6050 GNDA.n6049 185
R9248 GNDA.n6052 GNDA.n6051 185
R9249 GNDA.n6054 GNDA.n6053 185
R9250 GNDA.n6056 GNDA.n6055 185
R9251 GNDA.n6057 GNDA.n5451 185
R9252 GNDA.n6024 GNDA.n6023 185
R9253 GNDA.n6026 GNDA.n6025 185
R9254 GNDA.n6028 GNDA.n6027 185
R9255 GNDA.n6030 GNDA.n6029 185
R9256 GNDA.n6032 GNDA.n6031 185
R9257 GNDA.n6034 GNDA.n6033 185
R9258 GNDA.n6036 GNDA.n6035 185
R9259 GNDA.n6038 GNDA.n6037 185
R9260 GNDA.n6040 GNDA.n6039 185
R9261 GNDA.n6006 GNDA.n6005 185
R9262 GNDA.n6008 GNDA.n6007 185
R9263 GNDA.n6010 GNDA.n6009 185
R9264 GNDA.n6012 GNDA.n6011 185
R9265 GNDA.n6014 GNDA.n6013 185
R9266 GNDA.n6016 GNDA.n6015 185
R9267 GNDA.n6018 GNDA.n6017 185
R9268 GNDA.n6020 GNDA.n6019 185
R9269 GNDA.n6022 GNDA.n6021 185
R9270 GNDA.n6004 GNDA.n6003 185
R9271 GNDA.n5494 GNDA.n5493 185
R9272 GNDA.n5492 GNDA.n5491 185
R9273 GNDA.n5500 GNDA.n5499 185
R9274 GNDA.n5502 GNDA.n5501 185
R9275 GNDA.n5505 GNDA.n5504 185
R9276 GNDA.n5488 GNDA.n5456 185
R9277 GNDA.n6061 GNDA.n6060 185
R9278 GNDA.n5455 GNDA.n5452 185
R9279 GNDA.n5967 GNDA.n5906 185
R9280 GNDA.n5981 GNDA.n5980 185
R9281 GNDA.n5979 GNDA.n5907 185
R9282 GNDA.n5978 GNDA.n5977 185
R9283 GNDA.n5976 GNDA.n5975 185
R9284 GNDA.n5974 GNDA.n5973 185
R9285 GNDA.n5972 GNDA.n5971 185
R9286 GNDA.n5970 GNDA.n5969 185
R9287 GNDA.n5968 GNDA.n5883 185
R9288 GNDA.n5950 GNDA.n5949 185
R9289 GNDA.n5952 GNDA.n5951 185
R9290 GNDA.n5954 GNDA.n5953 185
R9291 GNDA.n5956 GNDA.n5955 185
R9292 GNDA.n5958 GNDA.n5957 185
R9293 GNDA.n5960 GNDA.n5959 185
R9294 GNDA.n5962 GNDA.n5961 185
R9295 GNDA.n5964 GNDA.n5963 185
R9296 GNDA.n5966 GNDA.n5965 185
R9297 GNDA.n5932 GNDA.n5931 185
R9298 GNDA.n5934 GNDA.n5933 185
R9299 GNDA.n5936 GNDA.n5935 185
R9300 GNDA.n5938 GNDA.n5937 185
R9301 GNDA.n5940 GNDA.n5939 185
R9302 GNDA.n5942 GNDA.n5941 185
R9303 GNDA.n5944 GNDA.n5943 185
R9304 GNDA.n5946 GNDA.n5945 185
R9305 GNDA.n5948 GNDA.n5947 185
R9306 GNDA.n5930 GNDA.n5929 185
R9307 GNDA.n5924 GNDA.n5923 185
R9308 GNDA.n5922 GNDA.n5921 185
R9309 GNDA.n5917 GNDA.n5916 185
R9310 GNDA.n5912 GNDA.n5891 185
R9311 GNDA.n5985 GNDA.n5984 185
R9312 GNDA.n5890 GNDA.n5888 185
R9313 GNDA.n5991 GNDA.n5990 185
R9314 GNDA.n5993 GNDA.n5992 185
R9315 GNDA.n6722 GNDA.n6721 185
R9316 GNDA.n6723 GNDA.n6674 185
R9317 GNDA.n6725 GNDA.n6724 185
R9318 GNDA.n6727 GNDA.n6673 185
R9319 GNDA.n6730 GNDA.n6729 185
R9320 GNDA.n6731 GNDA.n6672 185
R9321 GNDA.n6733 GNDA.n6732 185
R9322 GNDA.n6735 GNDA.n6671 185
R9323 GNDA.n6738 GNDA.n6737 185
R9324 GNDA.n6703 GNDA.n6679 185
R9325 GNDA.n6706 GNDA.n6705 185
R9326 GNDA.n6707 GNDA.n6678 185
R9327 GNDA.n6709 GNDA.n6708 185
R9328 GNDA.n6711 GNDA.n6677 185
R9329 GNDA.n6714 GNDA.n6713 185
R9330 GNDA.n6715 GNDA.n6676 185
R9331 GNDA.n6717 GNDA.n6716 185
R9332 GNDA.n6719 GNDA.n6675 185
R9333 GNDA.n6685 GNDA.n292 185
R9334 GNDA.n6689 GNDA.n6686 185
R9335 GNDA.n6691 GNDA.n6690 185
R9336 GNDA.n6692 GNDA.n6683 185
R9337 GNDA.n6694 GNDA.n6693 185
R9338 GNDA.n6696 GNDA.n6681 185
R9339 GNDA.n6698 GNDA.n6697 185
R9340 GNDA.n6699 GNDA.n6680 185
R9341 GNDA.n6701 GNDA.n6700 185
R9342 GNDA.n7028 GNDA.n7027 185
R9343 GNDA.n7025 GNDA.n290 185
R9344 GNDA.n7024 GNDA.n294 185
R9345 GNDA.n7022 GNDA.n7021 185
R9346 GNDA.n6759 GNDA.n295 185
R9347 GNDA.n6757 GNDA.n6756 185
R9348 GNDA.n6754 GNDA.n6668 185
R9349 GNDA.n6752 GNDA.n6751 185
R9350 GNDA.n6740 GNDA.n6669 185
R9351 GNDA.n7334 GNDA.n7333 185
R9352 GNDA.n7332 GNDA.n7331 185
R9353 GNDA.n7330 GNDA.n7329 185
R9354 GNDA.n7328 GNDA.n7327 185
R9355 GNDA.n7326 GNDA.n7325 185
R9356 GNDA.n7324 GNDA.n7323 185
R9357 GNDA.n7322 GNDA.n7321 185
R9358 GNDA.n7320 GNDA.n7319 185
R9359 GNDA.n7318 GNDA.n20 185
R9360 GNDA.n7352 GNDA.n7351 185
R9361 GNDA.n7350 GNDA.n7349 185
R9362 GNDA.n7348 GNDA.n7347 185
R9363 GNDA.n7346 GNDA.n7345 185
R9364 GNDA.n7344 GNDA.n7343 185
R9365 GNDA.n7342 GNDA.n7341 185
R9366 GNDA.n7340 GNDA.n7339 185
R9367 GNDA.n7338 GNDA.n7337 185
R9368 GNDA.n7336 GNDA.n7335 185
R9369 GNDA.n7370 GNDA.n7369 185
R9370 GNDA.n7368 GNDA.n7367 185
R9371 GNDA.n7366 GNDA.n7365 185
R9372 GNDA.n7364 GNDA.n7363 185
R9373 GNDA.n7362 GNDA.n7361 185
R9374 GNDA.n7360 GNDA.n7359 185
R9375 GNDA.n7358 GNDA.n7357 185
R9376 GNDA.n7356 GNDA.n7355 185
R9377 GNDA.n7354 GNDA.n7353 185
R9378 GNDA.n7372 GNDA.n7371 185
R9379 GNDA.n7378 GNDA.n7377 185
R9380 GNDA.n7373 GNDA.n3 185
R9381 GNDA.n7491 GNDA.n7490 185
R9382 GNDA.n34 GNDA.n2 185
R9383 GNDA.n38 GNDA.n37 185
R9384 GNDA.n36 GNDA.n33 185
R9385 GNDA.n23 GNDA.n21 185
R9386 GNDA.n7487 GNDA.n7486 185
R9387 GNDA.n7411 GNDA.n7306 175.546
R9388 GNDA.n7407 GNDA.n7306 175.546
R9389 GNDA.n7407 GNDA.n7308 175.546
R9390 GNDA.n7403 GNDA.n7308 175.546
R9391 GNDA.n7403 GNDA.n7310 175.546
R9392 GNDA.n7399 GNDA.n7310 175.546
R9393 GNDA.n7399 GNDA.n7312 175.546
R9394 GNDA.n7395 GNDA.n7312 175.546
R9395 GNDA.n7395 GNDA.n7314 175.546
R9396 GNDA.n7391 GNDA.n7314 175.546
R9397 GNDA.n7391 GNDA.n7316 175.546
R9398 GNDA.n7291 GNDA.n7289 175.546
R9399 GNDA.n7287 GNDA.n7253 175.546
R9400 GNDA.n7283 GNDA.n7281 175.546
R9401 GNDA.n7279 GNDA.n7261 175.546
R9402 GNDA.n7275 GNDA.n7273 175.546
R9403 GNDA.n7435 GNDA.n7248 175.546
R9404 GNDA.n7431 GNDA.n7248 175.546
R9405 GNDA.n7431 GNDA.n7296 175.546
R9406 GNDA.n7427 GNDA.n7296 175.546
R9407 GNDA.n7427 GNDA.n7298 175.546
R9408 GNDA.n7423 GNDA.n7298 175.546
R9409 GNDA.n7423 GNDA.n7300 175.546
R9410 GNDA.n7419 GNDA.n7300 175.546
R9411 GNDA.n7419 GNDA.n7302 175.546
R9412 GNDA.n7415 GNDA.n7302 175.546
R9413 GNDA.n7415 GNDA.n7304 175.546
R9414 GNDA.n5781 GNDA.n5629 175.546
R9415 GNDA.n5777 GNDA.n5629 175.546
R9416 GNDA.n5777 GNDA.n5631 175.546
R9417 GNDA.n5773 GNDA.n5631 175.546
R9418 GNDA.n5773 GNDA.n5770 175.546
R9419 GNDA.n5770 GNDA.n5769 175.546
R9420 GNDA.n5769 GNDA.n5634 175.546
R9421 GNDA.n5765 GNDA.n5634 175.546
R9422 GNDA.n5765 GNDA.n5637 175.546
R9423 GNDA.n5761 GNDA.n5637 175.546
R9424 GNDA.n5761 GNDA.n5640 175.546
R9425 GNDA.n5805 GNDA.n5581 175.546
R9426 GNDA.n5616 GNDA.n5586 175.546
R9427 GNDA.n5612 GNDA.n5611 175.546
R9428 GNDA.n5608 GNDA.n5607 175.546
R9429 GNDA.n5604 GNDA.n5603 175.546
R9430 GNDA.n5800 GNDA.n5620 175.546
R9431 GNDA.n5796 GNDA.n5795 175.546
R9432 GNDA.n5793 GNDA.n5623 175.546
R9433 GNDA.n5789 GNDA.n5788 175.546
R9434 GNDA.n5786 GNDA.n5626 175.546
R9435 GNDA.n5807 GNDA.n5579 175.546
R9436 GNDA.n5589 GNDA.n5588 175.546
R9437 GNDA.n5592 GNDA.n5591 175.546
R9438 GNDA.n5595 GNDA.n5594 175.546
R9439 GNDA.n5598 GNDA.n5597 175.546
R9440 GNDA.n5828 GNDA.n5569 175.546
R9441 GNDA.n5824 GNDA.n5823 175.546
R9442 GNDA.n5821 GNDA.n5572 175.546
R9443 GNDA.n5817 GNDA.n5816 175.546
R9444 GNDA.n5814 GNDA.n5575 175.546
R9445 GNDA.n5833 GNDA.n5530 175.546
R9446 GNDA.n5565 GNDA.n5535 175.546
R9447 GNDA.n5561 GNDA.n5560 175.546
R9448 GNDA.n5557 GNDA.n5556 175.546
R9449 GNDA.n5553 GNDA.n5552 175.546
R9450 GNDA.n5863 GNDA.n5862 175.546
R9451 GNDA.n5867 GNDA.n5866 175.546
R9452 GNDA.n5871 GNDA.n5870 175.546
R9453 GNDA.n5875 GNDA.n5874 175.546
R9454 GNDA.n5879 GNDA.n5878 175.546
R9455 GNDA.n5856 GNDA.n5517 175.546
R9456 GNDA.n5852 GNDA.n5851 175.546
R9457 GNDA.n5849 GNDA.n5520 175.546
R9458 GNDA.n5845 GNDA.n5844 175.546
R9459 GNDA.n5842 GNDA.n5523 175.546
R9460 GNDA.n5835 GNDA.n5528 175.546
R9461 GNDA.n5538 GNDA.n5537 175.546
R9462 GNDA.n5541 GNDA.n5540 175.546
R9463 GNDA.n5544 GNDA.n5543 175.546
R9464 GNDA.n5547 GNDA.n5546 175.546
R9465 GNDA.n7254 GNDA.n7251 175.546
R9466 GNDA.n7257 GNDA.n7256 175.546
R9467 GNDA.n7262 GNDA.n7259 175.546
R9468 GNDA.n7265 GNDA.n7264 175.546
R9469 GNDA.n7270 GNDA.n7267 175.546
R9470 GNDA.n7461 GNDA.n80 175.546
R9471 GNDA.n7457 GNDA.n80 175.546
R9472 GNDA.n7457 GNDA.n83 175.546
R9473 GNDA.n7453 GNDA.n83 175.546
R9474 GNDA.n7453 GNDA.n85 175.546
R9475 GNDA.n7448 GNDA.n85 175.546
R9476 GNDA.n7448 GNDA.n88 175.546
R9477 GNDA.n7444 GNDA.n88 175.546
R9478 GNDA.n7444 GNDA.n7241 175.546
R9479 GNDA.n7440 GNDA.n7241 175.546
R9480 GNDA.n7440 GNDA.n7243 175.546
R9481 GNDA.n6447 GNDA.n6446 175.546
R9482 GNDA.n6357 GNDA.n6356 175.546
R9483 GNDA.n6363 GNDA.n6362 175.546
R9484 GNDA.n6371 GNDA.n6370 175.546
R9485 GNDA.n7480 GNDA.n55 175.546
R9486 GNDA.n6295 GNDA.n6293 175.546
R9487 GNDA.n6291 GNDA.n6271 175.546
R9488 GNDA.n6287 GNDA.n6285 175.546
R9489 GNDA.n6283 GNDA.n6278 175.546
R9490 GNDA.n7469 GNDA.n69 175.546
R9491 GNDA.n6269 GNDA.n6268 175.546
R9492 GNDA.n6273 GNDA.n6272 175.546
R9493 GNDA.n6275 GNDA.n6274 175.546
R9494 GNDA.n6280 GNDA.n6279 175.546
R9495 GNDA.n7467 GNDA.n71 175.546
R9496 GNDA.n6542 GNDA.n6541 175.546
R9497 GNDA.n6458 GNDA.n6457 175.546
R9498 GNDA.n6464 GNDA.n6463 175.546
R9499 GNDA.n6471 GNDA.n6470 175.546
R9500 GNDA.n6479 GNDA.n6478 175.546
R9501 GNDA.n6256 GNDA.n6255 175.546
R9502 GNDA.n6564 GNDA.n6255 175.546
R9503 GNDA.n6562 GNDA.n6561 175.546
R9504 GNDA.n6558 GNDA.n6557 175.546
R9505 GNDA.n6554 GNDA.n6553 175.546
R9506 GNDA.n6550 GNDA.n6549 175.546
R9507 GNDA.n6320 GNDA.n6257 175.546
R9508 GNDA.n6320 GNDA.n6259 175.546
R9509 GNDA.n6316 GNDA.n6259 175.546
R9510 GNDA.n6316 GNDA.n6262 175.546
R9511 GNDA.n6312 GNDA.n6262 175.546
R9512 GNDA.n6312 GNDA.n6264 175.546
R9513 GNDA.n6308 GNDA.n6264 175.546
R9514 GNDA.n6308 GNDA.n6266 175.546
R9515 GNDA.n6304 GNDA.n6266 175.546
R9516 GNDA.n6304 GNDA.n6301 175.546
R9517 GNDA.n6301 GNDA.n6300 175.546
R9518 GNDA.n6178 GNDA.n6177 175.546
R9519 GNDA.n6183 GNDA.n6180 175.546
R9520 GNDA.n6186 GNDA.n6185 175.546
R9521 GNDA.n6190 GNDA.n6188 175.546
R9522 GNDA.n6916 GNDA.n5392 175.546
R9523 GNDA.n6823 GNDA.n5404 175.546
R9524 GNDA.n6642 GNDA.n5404 175.546
R9525 GNDA.n6814 GNDA.n6642 175.546
R9526 GNDA.n6814 GNDA.n6643 175.546
R9527 GNDA.n6810 GNDA.n6643 175.546
R9528 GNDA.n6810 GNDA.n6796 175.546
R9529 GNDA.n6796 GNDA.n5400 175.546
R9530 GNDA.n6827 GNDA.n5400 175.546
R9531 GNDA.n6827 GNDA.n5394 175.546
R9532 GNDA.n6909 GNDA.n5394 175.546
R9533 GNDA.n6909 GNDA.n5393 175.546
R9534 GNDA.n6249 GNDA.n5426 175.546
R9535 GNDA.n6247 GNDA.n6246 175.546
R9536 GNDA.n6243 GNDA.n6242 175.546
R9537 GNDA.n6239 GNDA.n6238 175.546
R9538 GNDA.n6235 GNDA.n5406 175.546
R9539 GNDA.n6573 GNDA.n5406 175.546
R9540 GNDA.n6232 GNDA.n6230 175.546
R9541 GNDA.n6228 GNDA.n5429 175.546
R9542 GNDA.n6224 GNDA.n6222 175.546
R9543 GNDA.n6220 GNDA.n5431 175.546
R9544 GNDA.n6216 GNDA.n6214 175.546
R9545 GNDA.n5741 GNDA.n5740 175.546
R9546 GNDA.n5737 GNDA.n5736 175.546
R9547 GNDA.n5730 GNDA.n5729 175.546
R9548 GNDA.n5723 GNDA.n5722 175.546
R9549 GNDA.n5751 GNDA.n5750 175.546
R9550 GNDA.n6064 GNDA.n6063 175.546
R9551 GNDA.n5507 GNDA.n5487 175.546
R9552 GNDA.n5489 GNDA.n5486 175.546
R9553 GNDA.n5497 GNDA.n5496 175.546
R9554 GNDA.n6001 GNDA.n5475 175.546
R9555 GNDA.n5884 GNDA.n5514 175.546
R9556 GNDA.n5988 GNDA.n5987 175.546
R9557 GNDA.n5914 GNDA.n5913 175.546
R9558 GNDA.n5919 GNDA.n5918 175.546
R9559 GNDA.n5927 GNDA.n5926 175.546
R9560 GNDA.n6098 GNDA.n6085 175.546
R9561 GNDA.n6094 GNDA.n6085 175.546
R9562 GNDA.n6094 GNDA.n6087 175.546
R9563 GNDA.n6090 GNDA.n6087 175.546
R9564 GNDA.n6090 GNDA.n300 175.546
R9565 GNDA.n7015 GNDA.n300 175.546
R9566 GNDA.n7015 GNDA.n301 175.546
R9567 GNDA.n7011 GNDA.n301 175.546
R9568 GNDA.n7011 GNDA.n304 175.546
R9569 GNDA.n7007 GNDA.n304 175.546
R9570 GNDA.n7007 GNDA.n306 175.546
R9571 GNDA.n6744 GNDA.n5372 175.546
R9572 GNDA.n6745 GNDA.n6744 175.546
R9573 GNDA.n6749 GNDA.n6745 175.546
R9574 GNDA.n6749 GNDA.n6666 175.546
R9575 GNDA.n6761 GNDA.n6666 175.546
R9576 GNDA.n6761 GNDA.n296 175.546
R9577 GNDA.n7019 GNDA.n296 175.546
R9578 GNDA.n7019 GNDA.n288 175.546
R9579 GNDA.n7030 GNDA.n288 175.546
R9580 GNDA.n7030 GNDA.n289 175.546
R9581 GNDA.n308 GNDA.n289 175.546
R9582 GNDA.n6146 GNDA.n6145 175.546
R9583 GNDA.n6142 GNDA.n6141 175.546
R9584 GNDA.n6139 GNDA.n6126 175.546
R9585 GNDA.n6135 GNDA.n6133 175.546
R9586 GNDA.n6928 GNDA.n5373 175.546
R9587 GNDA.n6117 GNDA.n6076 175.546
R9588 GNDA.n6113 GNDA.n6112 175.546
R9589 GNDA.n6110 GNDA.n6079 175.546
R9590 GNDA.n6106 GNDA.n6105 175.546
R9591 GNDA.n6103 GNDA.n6082 175.546
R9592 GNDA.n6122 GNDA.n6121 175.546
R9593 GNDA.n6124 GNDA.n6123 175.546
R9594 GNDA.n6128 GNDA.n6127 175.546
R9595 GNDA.n6130 GNDA.n6129 175.546
R9596 GNDA.n6926 GNDA.n5375 175.546
R9597 GNDA.n5388 GNDA.n5346 175.546
R9598 GNDA.n6972 GNDA.n5346 175.546
R9599 GNDA.n6972 GNDA.n5347 175.546
R9600 GNDA.n6968 GNDA.n5347 175.546
R9601 GNDA.n6968 GNDA.n5321 175.546
R9602 GNDA.n6981 GNDA.n5321 175.546
R9603 GNDA.n6981 GNDA.n5322 175.546
R9604 GNDA.n6840 GNDA.n5322 175.546
R9605 GNDA.n6845 GNDA.n6840 175.546
R9606 GNDA.n6845 GNDA.n5366 175.546
R9607 GNDA.n6935 GNDA.n5366 175.546
R9608 GNDA.n6206 GNDA.n6205 175.546
R9609 GNDA.n6202 GNDA.n6201 175.546
R9610 GNDA.n6199 GNDA.n6182 175.546
R9611 GNDA.n6195 GNDA.n6193 175.546
R9612 GNDA.n6918 GNDA.n5390 175.546
R9613 GNDA.n6172 GNDA.n5437 175.546
R9614 GNDA.n6168 GNDA.n6166 175.546
R9615 GNDA.n6164 GNDA.n5439 175.546
R9616 GNDA.n6160 GNDA.n6158 175.546
R9617 GNDA.n6156 GNDA.n5441 175.546
R9618 GNDA.n7484 GNDA.n24 175.546
R9619 GNDA.n40 GNDA.n25 175.546
R9620 GNDA.n31 GNDA.n30 175.546
R9621 GNDA.n7375 GNDA.n7374 175.546
R9622 GNDA.n7381 GNDA.n7380 175.546
R9623 GNDA.n5527 GNDA.t145 172.876
R9624 GNDA.n5578 GNDA.t145 172.876
R9625 GNDA.n5567 GNDA.t145 172.615
R9626 GNDA.n5618 GNDA.t145 172.615
R9627 GNDA.n6483 GNDA.n6482 163.333
R9628 GNDA.n6382 GNDA.n6381 163.333
R9629 GNDA.n6850 GNDA.n6849 163.333
R9630 GNDA.n6834 GNDA.n6833 163.333
R9631 GNDA.n5655 GNDA.n5645 163.333
R9632 GNDA.n6005 GNDA.n6004 163.333
R9633 GNDA.n5931 GNDA.n5930 163.333
R9634 GNDA.n7027 GNDA.n292 163.333
R9635 GNDA.n7371 GNDA.n7370 163.333
R9636 GNDA.n3386 GNDA.n3385 161.3
R9637 GNDA.n1728 GNDA.n1727 161.3
R9638 GNDA.n6515 GNDA.n6514 150
R9639 GNDA.n6511 GNDA.n6510 150
R9640 GNDA.n6507 GNDA.n6506 150
R9641 GNDA.n6503 GNDA.n6502 150
R9642 GNDA.n6499 GNDA.n6498 150
R9643 GNDA.n6495 GNDA.n6494 150
R9644 GNDA.n6491 GNDA.n6490 150
R9645 GNDA.n6487 GNDA.n6486 150
R9646 GNDA.n6538 GNDA.n6326 150
R9647 GNDA.n6460 GNDA.n6327 150
R9648 GNDA.n6468 GNDA.n6467 150
R9649 GNDA.n6475 GNDA.n6474 150
R9650 GNDA.n6523 GNDA.n6522 150
R9651 GNDA.n6527 GNDA.n6526 150
R9652 GNDA.n6531 GNDA.n6530 150
R9653 GNDA.n6535 GNDA.n6534 150
R9654 GNDA.n6420 GNDA.n6419 150
R9655 GNDA.n6416 GNDA.n6415 150
R9656 GNDA.n6412 GNDA.n6411 150
R9657 GNDA.n6408 GNDA.n6407 150
R9658 GNDA.n6404 GNDA.n6403 150
R9659 GNDA.n6400 GNDA.n6399 150
R9660 GNDA.n6396 GNDA.n6395 150
R9661 GNDA.n6392 GNDA.n6391 150
R9662 GNDA.n6443 GNDA.n6347 150
R9663 GNDA.n6359 GNDA.n6348 150
R9664 GNDA.n6367 GNDA.n6366 150
R9665 GNDA.n6375 GNDA.n6353 150
R9666 GNDA.n6428 GNDA.n6427 150
R9667 GNDA.n6432 GNDA.n6431 150
R9668 GNDA.n6436 GNDA.n6435 150
R9669 GNDA.n6440 GNDA.n6439 150
R9670 GNDA.n6882 GNDA.n6881 150
R9671 GNDA.n6878 GNDA.n6877 150
R9672 GNDA.n6874 GNDA.n6873 150
R9673 GNDA.n6870 GNDA.n6869 150
R9674 GNDA.n6866 GNDA.n6865 150
R9675 GNDA.n6862 GNDA.n6861 150
R9676 GNDA.n6858 GNDA.n6857 150
R9677 GNDA.n6854 GNDA.n6853 150
R9678 GNDA.n6975 GNDA.n5343 150
R9679 GNDA.n6965 GNDA.n6964 150
R9680 GNDA.n6978 GNDA.n5324 150
R9681 GNDA.n6836 GNDA.n5325 150
R9682 GNDA.n6890 GNDA.n6889 150
R9683 GNDA.n6894 GNDA.n6893 150
R9684 GNDA.n6898 GNDA.n6897 150
R9685 GNDA.n6900 GNDA.n5342 150
R9686 GNDA.n6619 GNDA.n6582 150
R9687 GNDA.n6615 GNDA.n6613 150
R9688 GNDA.n6611 GNDA.n6584 150
R9689 GNDA.n6607 GNDA.n6605 150
R9690 GNDA.n6603 GNDA.n6586 150
R9691 GNDA.n6599 GNDA.n6598 150
R9692 GNDA.n6596 GNDA.n6589 150
R9693 GNDA.n6592 GNDA.n6591 150
R9694 GNDA.n6818 GNDA.n6817 150
R9695 GNDA.n6805 GNDA.n6804 150
R9696 GNDA.n6807 GNDA.n6803 150
R9697 GNDA.n6831 GNDA.n5398 150
R9698 GNDA.n6627 GNDA.n6580 150
R9699 GNDA.n6631 GNDA.n6629 150
R9700 GNDA.n6635 GNDA.n6578 150
R9701 GNDA.n6638 GNDA.n6637 150
R9702 GNDA.n5695 GNDA.n5694 150
R9703 GNDA.n5691 GNDA.n5690 150
R9704 GNDA.n5687 GNDA.n5686 150
R9705 GNDA.n5683 GNDA.n5682 150
R9706 GNDA.n5679 GNDA.n5678 150
R9707 GNDA.n5675 GNDA.n5674 150
R9708 GNDA.n5671 GNDA.n5670 150
R9709 GNDA.n5667 GNDA.n5666 150
R9710 GNDA.n5744 GNDA.n5664 150
R9711 GNDA.n5733 GNDA.n5732 150
R9712 GNDA.n5726 GNDA.n5725 150
R9713 GNDA.n5747 GNDA.n5644 150
R9714 GNDA.n5703 GNDA.n5702 150
R9715 GNDA.n5707 GNDA.n5706 150
R9716 GNDA.n5711 GNDA.n5710 150
R9717 GNDA.n5713 GNDA.n5663 150
R9718 GNDA.n6037 GNDA.n6036 150
R9719 GNDA.n6033 GNDA.n6032 150
R9720 GNDA.n6029 GNDA.n6028 150
R9721 GNDA.n6025 GNDA.n6024 150
R9722 GNDA.n6021 GNDA.n6020 150
R9723 GNDA.n6017 GNDA.n6016 150
R9724 GNDA.n6013 GNDA.n6012 150
R9725 GNDA.n6009 GNDA.n6008 150
R9726 GNDA.n6060 GNDA.n5455 150
R9727 GNDA.n5504 GNDA.n5456 150
R9728 GNDA.n5501 GNDA.n5500 150
R9729 GNDA.n5493 GNDA.n5492 150
R9730 GNDA.n6045 GNDA.n6044 150
R9731 GNDA.n6049 GNDA.n6048 150
R9732 GNDA.n6053 GNDA.n6052 150
R9733 GNDA.n6057 GNDA.n6056 150
R9734 GNDA.n5963 GNDA.n5962 150
R9735 GNDA.n5959 GNDA.n5958 150
R9736 GNDA.n5955 GNDA.n5954 150
R9737 GNDA.n5951 GNDA.n5950 150
R9738 GNDA.n5947 GNDA.n5946 150
R9739 GNDA.n5943 GNDA.n5942 150
R9740 GNDA.n5939 GNDA.n5938 150
R9741 GNDA.n5935 GNDA.n5934 150
R9742 GNDA.n5992 GNDA.n5991 150
R9743 GNDA.n5984 GNDA.n5890 150
R9744 GNDA.n5916 GNDA.n5891 150
R9745 GNDA.n5923 GNDA.n5922 150
R9746 GNDA.n5981 GNDA.n5907 150
R9747 GNDA.n5977 GNDA.n5976 150
R9748 GNDA.n5973 GNDA.n5972 150
R9749 GNDA.n5969 GNDA.n5968 150
R9750 GNDA.n6717 GNDA.n6676 150
R9751 GNDA.n6713 GNDA.n6711 150
R9752 GNDA.n6709 GNDA.n6678 150
R9753 GNDA.n6705 GNDA.n6703 150
R9754 GNDA.n6701 GNDA.n6680 150
R9755 GNDA.n6697 GNDA.n6696 150
R9756 GNDA.n6694 GNDA.n6683 150
R9757 GNDA.n6690 GNDA.n6689 150
R9758 GNDA.n6752 GNDA.n6669 150
R9759 GNDA.n6756 GNDA.n6754 150
R9760 GNDA.n7022 GNDA.n295 150
R9761 GNDA.n7025 GNDA.n7024 150
R9762 GNDA.n6725 GNDA.n6674 150
R9763 GNDA.n6729 GNDA.n6727 150
R9764 GNDA.n6733 GNDA.n6672 150
R9765 GNDA.n6737 GNDA.n6735 150
R9766 GNDA.n7339 GNDA.n7338 150
R9767 GNDA.n7343 GNDA.n7342 150
R9768 GNDA.n7347 GNDA.n7346 150
R9769 GNDA.n7351 GNDA.n7350 150
R9770 GNDA.n7355 GNDA.n7354 150
R9771 GNDA.n7359 GNDA.n7358 150
R9772 GNDA.n7363 GNDA.n7362 150
R9773 GNDA.n7367 GNDA.n7366 150
R9774 GNDA.n7487 GNDA.n21 150
R9775 GNDA.n37 GNDA.n36 150
R9776 GNDA.n7490 GNDA.n2 150
R9777 GNDA.n7377 GNDA.n3 150
R9778 GNDA.n7331 GNDA.n7330 150
R9779 GNDA.n7327 GNDA.n7326 150
R9780 GNDA.n7323 GNDA.n7322 150
R9781 GNDA.n7319 GNDA.n20 150
R9782 GNDA.n3402 GNDA.n575 148.017
R9783 GNDA.n3399 GNDA.n574 148.017
R9784 GNDA.n5312 GNDA.n5311 148.017
R9785 GNDA.n5318 GNDA.n5317 148.017
R9786 GNDA.n6990 GNDA.n6989 137.382
R9787 GNDA.n7035 GNDA.n285 136.145
R9788 GNDA.n7036 GNDA.n284 136.145
R9789 GNDA.n7037 GNDA.n283 136.145
R9790 GNDA.n7040 GNDA.n280 136.145
R9791 GNDA.n7041 GNDA.n279 136.145
R9792 GNDA.n7044 GNDA.n276 136.145
R9793 GNDA.n7045 GNDA.n275 136.145
R9794 GNDA.n7046 GNDA.n274 136.145
R9795 GNDA.n7049 GNDA.n271 136.145
R9796 GNDA.n7050 GNDA.n270 136.145
R9797 GNDA.n6791 GNDA.n6784 134.268
R9798 GNDA.n6784 GNDA.n6782 134.268
R9799 GNDA.n5881 GNDA.n5420 132.721
R9800 GNDA.n7033 GNDA.t245 130.001
R9801 GNDA.n5364 GNDA.t180 130.001
R9802 GNDA.n5362 GNDA.t143 130.001
R9803 GNDA.n6956 GNDA.t188 130.001
R9804 GNDA.n5385 GNDA.t156 130.001
R9805 GNDA.n6647 GNDA.t248 130.001
R9806 GNDA.n6644 GNDA.t197 130.001
R9807 GNDA.n5407 GNDA.t150 130
R9808 GNDA.n7474 GNDA.n62 124.832
R9809 GNDA.n6071 GNDA.n5444 124.832
R9810 GNDA.n5600 GNDA.n5443 124.832
R9811 GNDA.n6069 GNDA.n5448 124.832
R9812 GNDA.n5549 GNDA.n5447 124.832
R9813 GNDA.n7268 GNDA.n60 124.832
R9814 GNDA.n7472 GNDA.n7471 124.832
R9815 GNDA.n7465 GNDA.n64 124.832
R9816 GNDA.n6914 GNDA.n6913 124.832
R9817 GNDA.n6931 GNDA.n6930 124.832
R9818 GNDA.n6924 GNDA.n5367 124.832
R9819 GNDA.n6921 GNDA.n6920 124.832
R9820 GNDA.n6991 GNDA.n6990 124.21
R9821 GNDA.n3410 GNDA.n3408 121.251
R9822 GNDA.n3418 GNDA.n3417 121.136
R9823 GNDA.n3416 GNDA.n3415 121.136
R9824 GNDA.n3414 GNDA.n3413 121.136
R9825 GNDA.n3412 GNDA.n3411 121.136
R9826 GNDA.n3410 GNDA.n3409 121.136
R9827 GNDA.n1788 GNDA.n1787 121.136
R9828 GNDA.n1790 GNDA.n1789 121.136
R9829 GNDA.n1792 GNDA.n1791 121.136
R9830 GNDA.n1794 GNDA.n1793 121.136
R9831 GNDA.n1796 GNDA.n1795 121.136
R9832 GNDA.n1798 GNDA.n1797 121.136
R9833 GNDA.n7234 GNDA.t315 111.674
R9834 GNDA.n7235 GNDA.t3 111.206
R9835 GNDA.n7058 GNDA.t307 111.206
R9836 GNDA.n7058 GNDA.t20 111.076
R9837 GNDA.n6764 GNDA.n6763 101.718
R9838 GNDA.n6787 GNDA.n6649 101.718
R9839 GNDA.n6793 GNDA.n6651 101.718
R9840 GNDA.n6775 GNDA.n6665 101.718
R9841 GNDA.n5383 GNDA.t145 47.6748
R9842 GNDA.t11 GNDA.n1737 97.5812
R9843 GNDA.n1737 GNDA.t299 97.5812
R9844 GNDA.n6824 GNDA.n5402 96.751
R9845 GNDA.n6826 GNDA.n5401 96.751
R9846 GNDA.n6971 GNDA.n6958 96.751
R9847 GNDA.n6844 GNDA.n6843 96.751
R9848 GNDA.n6748 GNDA.n6747 96.751
R9849 GNDA.n7031 GNDA.n287 96.751
R9850 GNDA.n309 GNDA.n287 96.751
R9851 GNDA.n6648 GNDA.n6646 93.526
R9852 GNDA.t145 GNDA.n6922 93.526
R9853 GNDA.n7018 GNDA.t29 93.526
R9854 GNDA.t145 GNDA.n5382 92.451
R9855 GNDA.n6771 GNDA.n6664 91.069
R9856 GNDA.n6766 GNDA.n6664 91.069
R9857 GNDA.n6768 GNDA.n6663 91.069
R9858 GNDA.n6769 GNDA.n6768 91.069
R9859 GNDA.n6791 GNDA.n6786 91.069
R9860 GNDA.n6789 GNDA.n6782 91.069
R9861 GNDA.t45 GNDA.n6812 89.226
R9862 GNDA.n7032 GNDA.n7031 89.226
R9863 GNDA.n6795 GNDA.t334 88.151
R9864 GNDA.n6969 GNDA.t286 88.151
R9865 GNDA.t293 GNDA.n6746 88.151
R9866 GNDA.t67 GNDA.t15 84.4226
R9867 GNDA.n7239 GNDA.n7238 84.306
R9868 GNDA.n6954 GNDA.n5350 84.306
R9869 GNDA.n6938 GNDA.n5361 84.306
R9870 GNDA.t251 GNDA.n6825 83.851
R9871 GNDA.n6841 GNDA.t58 83.851
R9872 GNDA.n6762 GNDA.t260 83.851
R9873 GNDA.t13 GNDA.n6911 77.4009
R9874 GNDA.n7290 GNDA.n7247 76.3222
R9875 GNDA.n7289 GNDA.n7288 76.3222
R9876 GNDA.n7282 GNDA.n7253 76.3222
R9877 GNDA.n7281 GNDA.n7280 76.3222
R9878 GNDA.n7274 GNDA.n7261 76.3222
R9879 GNDA.n7273 GNDA.n7272 76.3222
R9880 GNDA.n5804 GNDA.n5803 76.3222
R9881 GNDA.n5617 GNDA.n5581 76.3222
R9882 GNDA.n5586 GNDA.n5585 76.3222
R9883 GNDA.n5611 GNDA.n5584 76.3222
R9884 GNDA.n5607 GNDA.n5583 76.3222
R9885 GNDA.n5603 GNDA.n5582 76.3222
R9886 GNDA.n5801 GNDA.n5800 76.3222
R9887 GNDA.n5796 GNDA.n5622 76.3222
R9888 GNDA.n5794 GNDA.n5793 76.3222
R9889 GNDA.n5789 GNDA.n5625 76.3222
R9890 GNDA.n5787 GNDA.n5786 76.3222
R9891 GNDA.n5782 GNDA.n5628 76.3222
R9892 GNDA.n5808 GNDA.n5807 76.3222
R9893 GNDA.n5588 GNDA.n5587 76.3222
R9894 GNDA.n5591 GNDA.n5590 76.3222
R9895 GNDA.n5594 GNDA.n5593 76.3222
R9896 GNDA.n5597 GNDA.n5596 76.3222
R9897 GNDA.n5600 GNDA.n5599 76.3222
R9898 GNDA.n5829 GNDA.n5828 76.3222
R9899 GNDA.n5824 GNDA.n5571 76.3222
R9900 GNDA.n5822 GNDA.n5821 76.3222
R9901 GNDA.n5817 GNDA.n5574 76.3222
R9902 GNDA.n5815 GNDA.n5814 76.3222
R9903 GNDA.n5810 GNDA.n5576 76.3222
R9904 GNDA.n5832 GNDA.n5831 76.3222
R9905 GNDA.n5566 GNDA.n5530 76.3222
R9906 GNDA.n5535 GNDA.n5534 76.3222
R9907 GNDA.n5560 GNDA.n5533 76.3222
R9908 GNDA.n5556 GNDA.n5532 76.3222
R9909 GNDA.n5552 GNDA.n5531 76.3222
R9910 GNDA.n5859 GNDA.n5415 76.3222
R9911 GNDA.n5863 GNDA.n5416 76.3222
R9912 GNDA.n5867 GNDA.n5417 76.3222
R9913 GNDA.n5871 GNDA.n5418 76.3222
R9914 GNDA.n5875 GNDA.n5419 76.3222
R9915 GNDA.n5879 GNDA.n5420 76.3222
R9916 GNDA.n5857 GNDA.n5856 76.3222
R9917 GNDA.n5852 GNDA.n5519 76.3222
R9918 GNDA.n5850 GNDA.n5849 76.3222
R9919 GNDA.n5845 GNDA.n5522 76.3222
R9920 GNDA.n5843 GNDA.n5842 76.3222
R9921 GNDA.n5838 GNDA.n5525 76.3222
R9922 GNDA.n5836 GNDA.n5835 76.3222
R9923 GNDA.n5537 GNDA.n5536 76.3222
R9924 GNDA.n5540 GNDA.n5539 76.3222
R9925 GNDA.n5543 GNDA.n5542 76.3222
R9926 GNDA.n5546 GNDA.n5545 76.3222
R9927 GNDA.n5549 GNDA.n5548 76.3222
R9928 GNDA.n7251 GNDA.n7250 76.3222
R9929 GNDA.n7256 GNDA.n7255 76.3222
R9930 GNDA.n7259 GNDA.n7258 76.3222
R9931 GNDA.n7264 GNDA.n7263 76.3222
R9932 GNDA.n7267 GNDA.n7266 76.3222
R9933 GNDA.n7269 GNDA.n7268 76.3222
R9934 GNDA.n66 GNDA.n49 76.3222
R9935 GNDA.n6446 GNDA.n50 76.3222
R9936 GNDA.n6357 GNDA.n51 76.3222
R9937 GNDA.n6363 GNDA.n52 76.3222
R9938 GNDA.n6371 GNDA.n53 76.3222
R9939 GNDA.n7481 GNDA.n7480 76.3222
R9940 GNDA.n6294 GNDA.n79 76.3222
R9941 GNDA.n6293 GNDA.n6292 76.3222
R9942 GNDA.n6286 GNDA.n6271 76.3222
R9943 GNDA.n6285 GNDA.n6284 76.3222
R9944 GNDA.n6278 GNDA.n6277 76.3222
R9945 GNDA.n7470 GNDA.n7469 76.3222
R9946 GNDA.n6268 GNDA.n72 76.3222
R9947 GNDA.n6272 GNDA.n73 76.3222
R9948 GNDA.n6274 GNDA.n74 76.3222
R9949 GNDA.n6279 GNDA.n75 76.3222
R9950 GNDA.n76 GNDA.n71 76.3222
R9951 GNDA.n7466 GNDA.n7465 76.3222
R9952 GNDA.n6546 GNDA.n43 76.3222
R9953 GNDA.n6541 GNDA.n44 76.3222
R9954 GNDA.n6458 GNDA.n45 76.3222
R9955 GNDA.n6464 GNDA.n46 76.3222
R9956 GNDA.n6470 GNDA.n47 76.3222
R9957 GNDA.n6479 GNDA.n48 76.3222
R9958 GNDA.n6570 GNDA.n6569 76.3222
R9959 GNDA.n6564 GNDA.n5410 76.3222
R9960 GNDA.n6561 GNDA.n5411 76.3222
R9961 GNDA.n6557 GNDA.n5412 76.3222
R9962 GNDA.n6553 GNDA.n5413 76.3222
R9963 GNDA.n7467 GNDA.n7466 76.3222
R9964 GNDA.n6280 GNDA.n76 76.3222
R9965 GNDA.n6275 GNDA.n75 76.3222
R9966 GNDA.n6273 GNDA.n74 76.3222
R9967 GNDA.n6269 GNDA.n73 76.3222
R9968 GNDA.n6298 GNDA.n72 76.3222
R9969 GNDA.n6295 GNDA.n6294 76.3222
R9970 GNDA.n6292 GNDA.n6291 76.3222
R9971 GNDA.n6287 GNDA.n6286 76.3222
R9972 GNDA.n6284 GNDA.n6283 76.3222
R9973 GNDA.n6277 GNDA.n69 76.3222
R9974 GNDA.n7471 GNDA.n7470 76.3222
R9975 GNDA.n6176 GNDA.n5433 76.3222
R9976 GNDA.n6179 GNDA.n6178 76.3222
R9977 GNDA.n6184 GNDA.n6183 76.3222
R9978 GNDA.n6187 GNDA.n6186 76.3222
R9979 GNDA.n6190 GNDA.n6189 76.3222
R9980 GNDA.n6916 GNDA.n6915 76.3222
R9981 GNDA.n6254 GNDA.n6253 76.3222
R9982 GNDA.n6249 GNDA.n5425 76.3222
R9983 GNDA.n6246 GNDA.n5424 76.3222
R9984 GNDA.n6242 GNDA.n5423 76.3222
R9985 GNDA.n6238 GNDA.n5422 76.3222
R9986 GNDA.n6231 GNDA.n5427 76.3222
R9987 GNDA.n6230 GNDA.n6229 76.3222
R9988 GNDA.n6223 GNDA.n5429 76.3222
R9989 GNDA.n6222 GNDA.n6221 76.3222
R9990 GNDA.n6215 GNDA.n5431 76.3222
R9991 GNDA.n6213 GNDA.n6212 76.3222
R9992 GNDA.n5483 GNDA.n5445 76.3222
R9993 GNDA.n5741 GNDA.n5482 76.3222
R9994 GNDA.n5736 GNDA.n5481 76.3222
R9995 GNDA.n5729 GNDA.n5480 76.3222
R9996 GNDA.n5722 GNDA.n5479 76.3222
R9997 GNDA.n5751 GNDA.n5478 76.3222
R9998 GNDA.n6068 GNDA.n5449 76.3222
R9999 GNDA.n6063 GNDA.n5453 76.3222
R10000 GNDA.n5508 GNDA.n5507 76.3222
R10001 GNDA.n5489 GNDA.n5485 76.3222
R10002 GNDA.n5496 GNDA.n5484 76.3222
R10003 GNDA.n6001 GNDA.n6000 76.3222
R10004 GNDA.n5998 GNDA.n5997 76.3222
R10005 GNDA.n5884 GNDA.n5513 76.3222
R10006 GNDA.n5987 GNDA.n5512 76.3222
R10007 GNDA.n5914 GNDA.n5511 76.3222
R10008 GNDA.n5918 GNDA.n5510 76.3222
R10009 GNDA.n5927 GNDA.n5509 76.3222
R10010 GNDA.n6148 GNDA.n6147 76.3222
R10011 GNDA.n6145 GNDA.n6120 76.3222
R10012 GNDA.n6141 GNDA.n6140 76.3222
R10013 GNDA.n6134 GNDA.n6126 76.3222
R10014 GNDA.n6133 GNDA.n6132 76.3222
R10015 GNDA.n6929 GNDA.n6928 76.3222
R10016 GNDA.n6118 GNDA.n6117 76.3222
R10017 GNDA.n6113 GNDA.n6078 76.3222
R10018 GNDA.n6111 GNDA.n6110 76.3222
R10019 GNDA.n6106 GNDA.n6081 76.3222
R10020 GNDA.n6104 GNDA.n6103 76.3222
R10021 GNDA.n6099 GNDA.n6084 76.3222
R10022 GNDA.n6084 GNDA.n6082 76.3222
R10023 GNDA.n6105 GNDA.n6104 76.3222
R10024 GNDA.n6081 GNDA.n6079 76.3222
R10025 GNDA.n6112 GNDA.n6111 76.3222
R10026 GNDA.n6078 GNDA.n6076 76.3222
R10027 GNDA.n6119 GNDA.n6118 76.3222
R10028 GNDA.n5998 GNDA.n5514 76.3222
R10029 GNDA.n5988 GNDA.n5513 76.3222
R10030 GNDA.n5913 GNDA.n5512 76.3222
R10031 GNDA.n5919 GNDA.n5511 76.3222
R10032 GNDA.n5926 GNDA.n5510 76.3222
R10033 GNDA.n5908 GNDA.n5509 76.3222
R10034 GNDA.n6064 GNDA.n5449 76.3222
R10035 GNDA.n5487 GNDA.n5453 76.3222
R10036 GNDA.n5508 GNDA.n5486 76.3222
R10037 GNDA.n5497 GNDA.n5485 76.3222
R10038 GNDA.n5484 GNDA.n5475 76.3222
R10039 GNDA.n6000 GNDA.n5477 76.3222
R10040 GNDA.n5740 GNDA.n5483 76.3222
R10041 GNDA.n5737 GNDA.n5482 76.3222
R10042 GNDA.n5730 GNDA.n5481 76.3222
R10043 GNDA.n5723 GNDA.n5480 76.3222
R10044 GNDA.n5750 GNDA.n5479 76.3222
R10045 GNDA.n5755 GNDA.n5478 76.3222
R10046 GNDA.n6121 GNDA.n5376 76.3222
R10047 GNDA.n6123 GNDA.n5377 76.3222
R10048 GNDA.n6127 GNDA.n5378 76.3222
R10049 GNDA.n6129 GNDA.n5379 76.3222
R10050 GNDA.n5380 GNDA.n5375 76.3222
R10051 GNDA.n6925 GNDA.n6924 76.3222
R10052 GNDA.n6208 GNDA.n6207 76.3222
R10053 GNDA.n6205 GNDA.n6175 76.3222
R10054 GNDA.n6201 GNDA.n6200 76.3222
R10055 GNDA.n6194 GNDA.n6182 76.3222
R10056 GNDA.n6193 GNDA.n6192 76.3222
R10057 GNDA.n6919 GNDA.n6918 76.3222
R10058 GNDA.n6174 GNDA.n6173 76.3222
R10059 GNDA.n6167 GNDA.n5437 76.3222
R10060 GNDA.n6166 GNDA.n6165 76.3222
R10061 GNDA.n6159 GNDA.n5439 76.3222
R10062 GNDA.n6158 GNDA.n6157 76.3222
R10063 GNDA.n6151 GNDA.n5441 76.3222
R10064 GNDA.n6152 GNDA.n6151 76.3222
R10065 GNDA.n6157 GNDA.n6156 76.3222
R10066 GNDA.n6160 GNDA.n6159 76.3222
R10067 GNDA.n6165 GNDA.n6164 76.3222
R10068 GNDA.n6168 GNDA.n6167 76.3222
R10069 GNDA.n6173 GNDA.n6172 76.3222
R10070 GNDA.n6214 GNDA.n6213 76.3222
R10071 GNDA.n6216 GNDA.n6215 76.3222
R10072 GNDA.n6221 GNDA.n6220 76.3222
R10073 GNDA.n6224 GNDA.n6223 76.3222
R10074 GNDA.n6229 GNDA.n6228 76.3222
R10075 GNDA.n6232 GNDA.n6231 76.3222
R10076 GNDA.n6915 GNDA.n6914 76.3222
R10077 GNDA.n6189 GNDA.n5392 76.3222
R10078 GNDA.n6188 GNDA.n6187 76.3222
R10079 GNDA.n6185 GNDA.n6184 76.3222
R10080 GNDA.n6180 GNDA.n6179 76.3222
R10081 GNDA.n6177 GNDA.n6176 76.3222
R10082 GNDA.n6207 GNDA.n6206 76.3222
R10083 GNDA.n6202 GNDA.n6175 76.3222
R10084 GNDA.n6200 GNDA.n6199 76.3222
R10085 GNDA.n6195 GNDA.n6194 76.3222
R10086 GNDA.n6192 GNDA.n5390 76.3222
R10087 GNDA.n6920 GNDA.n6919 76.3222
R10088 GNDA.n5548 GNDA.n5547 76.3222
R10089 GNDA.n5545 GNDA.n5544 76.3222
R10090 GNDA.n5542 GNDA.n5541 76.3222
R10091 GNDA.n5539 GNDA.n5538 76.3222
R10092 GNDA.n5536 GNDA.n5528 76.3222
R10093 GNDA.n5837 GNDA.n5836 76.3222
R10094 GNDA.n5833 GNDA.n5832 76.3222
R10095 GNDA.n5566 GNDA.n5565 76.3222
R10096 GNDA.n5561 GNDA.n5534 76.3222
R10097 GNDA.n5557 GNDA.n5533 76.3222
R10098 GNDA.n5553 GNDA.n5532 76.3222
R10099 GNDA.n5531 GNDA.n5448 76.3222
R10100 GNDA.n5525 GNDA.n5523 76.3222
R10101 GNDA.n5844 GNDA.n5843 76.3222
R10102 GNDA.n5522 GNDA.n5520 76.3222
R10103 GNDA.n5851 GNDA.n5850 76.3222
R10104 GNDA.n5519 GNDA.n5517 76.3222
R10105 GNDA.n5858 GNDA.n5857 76.3222
R10106 GNDA.n5576 GNDA.n5575 76.3222
R10107 GNDA.n5816 GNDA.n5815 76.3222
R10108 GNDA.n5574 GNDA.n5572 76.3222
R10109 GNDA.n5823 GNDA.n5822 76.3222
R10110 GNDA.n5571 GNDA.n5569 76.3222
R10111 GNDA.n5830 GNDA.n5829 76.3222
R10112 GNDA.n5628 GNDA.n5626 76.3222
R10113 GNDA.n5788 GNDA.n5787 76.3222
R10114 GNDA.n5625 GNDA.n5623 76.3222
R10115 GNDA.n5795 GNDA.n5794 76.3222
R10116 GNDA.n5622 GNDA.n5620 76.3222
R10117 GNDA.n5802 GNDA.n5801 76.3222
R10118 GNDA.n6542 GNDA.n43 76.3222
R10119 GNDA.n6457 GNDA.n44 76.3222
R10120 GNDA.n6463 GNDA.n45 76.3222
R10121 GNDA.n6471 GNDA.n46 76.3222
R10122 GNDA.n6478 GNDA.n47 76.3222
R10123 GNDA.n6452 GNDA.n48 76.3222
R10124 GNDA.n6447 GNDA.n49 76.3222
R10125 GNDA.n6356 GNDA.n50 76.3222
R10126 GNDA.n6362 GNDA.n51 76.3222
R10127 GNDA.n6370 GNDA.n52 76.3222
R10128 GNDA.n55 GNDA.n53 76.3222
R10129 GNDA.n7481 GNDA.n54 76.3222
R10130 GNDA.n42 GNDA.n24 76.3222
R10131 GNDA.n7483 GNDA.n25 76.3222
R10132 GNDA.n41 GNDA.n31 76.3222
R10133 GNDA.n7374 GNDA.n29 76.3222
R10134 GNDA.n7380 GNDA.n28 76.3222
R10135 GNDA.n7385 GNDA.n27 76.3222
R10136 GNDA.n63 GNDA.n42 76.3222
R10137 GNDA.n7484 GNDA.n7483 76.3222
R10138 GNDA.n41 GNDA.n40 76.3222
R10139 GNDA.n30 GNDA.n29 76.3222
R10140 GNDA.n7375 GNDA.n28 76.3222
R10141 GNDA.n7381 GNDA.n27 76.3222
R10142 GNDA.n7270 GNDA.n7269 76.3222
R10143 GNDA.n7266 GNDA.n7265 76.3222
R10144 GNDA.n7263 GNDA.n7262 76.3222
R10145 GNDA.n7258 GNDA.n7257 76.3222
R10146 GNDA.n7255 GNDA.n7254 76.3222
R10147 GNDA.n7250 GNDA.n7249 76.3222
R10148 GNDA.n7291 GNDA.n7290 76.3222
R10149 GNDA.n7288 GNDA.n7287 76.3222
R10150 GNDA.n7283 GNDA.n7282 76.3222
R10151 GNDA.n7280 GNDA.n7279 76.3222
R10152 GNDA.n7275 GNDA.n7274 76.3222
R10153 GNDA.n7272 GNDA.n62 76.3222
R10154 GNDA.n5599 GNDA.n5598 76.3222
R10155 GNDA.n5596 GNDA.n5595 76.3222
R10156 GNDA.n5593 GNDA.n5592 76.3222
R10157 GNDA.n5590 GNDA.n5589 76.3222
R10158 GNDA.n5587 GNDA.n5579 76.3222
R10159 GNDA.n5809 GNDA.n5808 76.3222
R10160 GNDA.n5805 GNDA.n5804 76.3222
R10161 GNDA.n5617 GNDA.n5616 76.3222
R10162 GNDA.n5612 GNDA.n5585 76.3222
R10163 GNDA.n5608 GNDA.n5584 76.3222
R10164 GNDA.n5604 GNDA.n5583 76.3222
R10165 GNDA.n5582 GNDA.n5444 76.3222
R10166 GNDA.n6926 GNDA.n6925 76.3222
R10167 GNDA.n6130 GNDA.n5380 76.3222
R10168 GNDA.n6128 GNDA.n5379 76.3222
R10169 GNDA.n6124 GNDA.n5378 76.3222
R10170 GNDA.n6122 GNDA.n5377 76.3222
R10171 GNDA.n6150 GNDA.n5376 76.3222
R10172 GNDA.n6147 GNDA.n6146 76.3222
R10173 GNDA.n6142 GNDA.n6120 76.3222
R10174 GNDA.n6140 GNDA.n6139 76.3222
R10175 GNDA.n6135 GNDA.n6134 76.3222
R10176 GNDA.n6132 GNDA.n5373 76.3222
R10177 GNDA.n6930 GNDA.n6929 76.3222
R10178 GNDA.n6254 GNDA.n5426 76.3222
R10179 GNDA.n6247 GNDA.n5425 76.3222
R10180 GNDA.n6243 GNDA.n5424 76.3222
R10181 GNDA.n6239 GNDA.n5423 76.3222
R10182 GNDA.n6235 GNDA.n5422 76.3222
R10183 GNDA.n5862 GNDA.n5415 76.3222
R10184 GNDA.n5866 GNDA.n5416 76.3222
R10185 GNDA.n5870 GNDA.n5417 76.3222
R10186 GNDA.n5874 GNDA.n5418 76.3222
R10187 GNDA.n5878 GNDA.n5419 76.3222
R10188 GNDA.n6570 GNDA.n6256 76.3222
R10189 GNDA.n6562 GNDA.n5410 76.3222
R10190 GNDA.n6558 GNDA.n5411 76.3222
R10191 GNDA.n6554 GNDA.n5412 76.3222
R10192 GNDA.n6550 GNDA.n5413 76.3222
R10193 GNDA.n6502 GNDA.n6333 74.5978
R10194 GNDA.n6499 GNDA.n6333 74.5978
R10195 GNDA.n6407 GNDA.n6377 74.5978
R10196 GNDA.n6404 GNDA.n6377 74.5978
R10197 GNDA.n6869 GNDA.n5331 74.5978
R10198 GNDA.n6866 GNDA.n5331 74.5978
R10199 GNDA.n6605 GNDA.n6604 74.5978
R10200 GNDA.n6604 GNDA.n6603 74.5978
R10201 GNDA.n5682 GNDA.n5651 74.5978
R10202 GNDA.n5679 GNDA.n5651 74.5978
R10203 GNDA.n6024 GNDA.n5462 74.5978
R10204 GNDA.n6021 GNDA.n5462 74.5978
R10205 GNDA.n5950 GNDA.n5896 74.5978
R10206 GNDA.n5947 GNDA.n5896 74.5978
R10207 GNDA.n6703 GNDA.n6702 74.5978
R10208 GNDA.n6702 GNDA.n6701 74.5978
R10209 GNDA.n7351 GNDA.n9 74.5978
R10210 GNDA.n7354 GNDA.n9 74.5978
R10211 GNDA.n6742 GNDA.t80 73.1009
R10212 GNDA.n7463 GNDA.n77 71.5297
R10213 GNDA.n7438 GNDA.n7437 71.5297
R10214 GNDA.n7463 GNDA.n7462 69.9996
R10215 GNDA.n7437 GNDA.n7436 69.9996
R10216 GNDA.n6536 GNDA.n6326 69.3109
R10217 GNDA.n6536 GNDA.n6535 69.3109
R10218 GNDA.n6441 GNDA.n6347 69.3109
R10219 GNDA.n6441 GNDA.n6440 69.3109
R10220 GNDA.n6976 GNDA.n6975 69.3109
R10221 GNDA.n6976 GNDA.n5342 69.3109
R10222 GNDA.n6818 GNDA.n6639 69.3109
R10223 GNDA.n6639 GNDA.n6638 69.3109
R10224 GNDA.n5745 GNDA.n5744 69.3109
R10225 GNDA.n5745 GNDA.n5663 69.3109
R10226 GNDA.n6058 GNDA.n5455 69.3109
R10227 GNDA.n6058 GNDA.n6057 69.3109
R10228 GNDA.n5992 GNDA.n5886 69.3109
R10229 GNDA.n5968 GNDA.n5886 69.3109
R10230 GNDA.n6736 GNDA.n6669 69.3109
R10231 GNDA.n6737 GNDA.n6736 69.3109
R10232 GNDA.n7488 GNDA.n7487 69.3109
R10233 GNDA.n7488 GNDA.n20 69.3109
R10234 GNDA.n6995 GNDA.n6994 69.2134
R10235 GNDA.n6970 GNDA.t257 66.6509
R10236 GNDA.n6743 GNDA.t4 66.6509
R10237 GNDA.t192 GNDA.n6343 65.8183
R10238 GNDA.t192 GNDA.n6342 65.8183
R10239 GNDA.t192 GNDA.n6341 65.8183
R10240 GNDA.t192 GNDA.n6340 65.8183
R10241 GNDA.t192 GNDA.n6331 65.8183
R10242 GNDA.t192 GNDA.n6338 65.8183
R10243 GNDA.t192 GNDA.n6328 65.8183
R10244 GNDA.t192 GNDA.n6339 65.8183
R10245 GNDA.t192 GNDA.n6337 65.8183
R10246 GNDA.t192 GNDA.n6336 65.8183
R10247 GNDA.t192 GNDA.n6335 65.8183
R10248 GNDA.t192 GNDA.n6334 65.8183
R10249 GNDA.t147 GNDA.n6389 65.8183
R10250 GNDA.t147 GNDA.n6388 65.8183
R10251 GNDA.t147 GNDA.n6387 65.8183
R10252 GNDA.t147 GNDA.n6386 65.8183
R10253 GNDA.t147 GNDA.n6352 65.8183
R10254 GNDA.t147 GNDA.n6384 65.8183
R10255 GNDA.t147 GNDA.n6349 65.8183
R10256 GNDA.t147 GNDA.n6385 65.8183
R10257 GNDA.t147 GNDA.n6383 65.8183
R10258 GNDA.t147 GNDA.n6380 65.8183
R10259 GNDA.t147 GNDA.n6379 65.8183
R10260 GNDA.t147 GNDA.n6378 65.8183
R10261 GNDA.t147 GNDA.n6376 65.8183
R10262 GNDA.t147 GNDA.n6351 65.8183
R10263 GNDA.t147 GNDA.n6350 65.8183
R10264 GNDA.n6442 GNDA.t147 65.8183
R10265 GNDA.t192 GNDA.n6332 65.8183
R10266 GNDA.t192 GNDA.n6330 65.8183
R10267 GNDA.t192 GNDA.n6329 65.8183
R10268 GNDA.n6537 GNDA.t192 65.8183
R10269 GNDA.t144 GNDA.n5341 65.8183
R10270 GNDA.t144 GNDA.n5340 65.8183
R10271 GNDA.t144 GNDA.n5339 65.8183
R10272 GNDA.t144 GNDA.n5338 65.8183
R10273 GNDA.t144 GNDA.n5329 65.8183
R10274 GNDA.t144 GNDA.n5336 65.8183
R10275 GNDA.t144 GNDA.n5327 65.8183
R10276 GNDA.t144 GNDA.n5337 65.8183
R10277 GNDA.t144 GNDA.n5335 65.8183
R10278 GNDA.t144 GNDA.n5334 65.8183
R10279 GNDA.t144 GNDA.n5333 65.8183
R10280 GNDA.t144 GNDA.n5332 65.8183
R10281 GNDA.t144 GNDA.n5330 65.8183
R10282 GNDA.n6977 GNDA.t144 65.8183
R10283 GNDA.t144 GNDA.n5328 65.8183
R10284 GNDA.t144 GNDA.n5326 65.8183
R10285 GNDA.n6622 GNDA.t146 65.8183
R10286 GNDA.n6628 GNDA.t146 65.8183
R10287 GNDA.n6630 GNDA.t146 65.8183
R10288 GNDA.n6636 GNDA.t146 65.8183
R10289 GNDA.n6606 GNDA.t146 65.8183
R10290 GNDA.n6612 GNDA.t146 65.8183
R10291 GNDA.n6614 GNDA.t146 65.8183
R10292 GNDA.n6620 GNDA.t146 65.8183
R10293 GNDA.t146 GNDA.n5397 65.8183
R10294 GNDA.n6590 GNDA.t146 65.8183
R10295 GNDA.n6597 GNDA.t146 65.8183
R10296 GNDA.n6588 GNDA.t146 65.8183
R10297 GNDA.n6832 GNDA.t146 65.8183
R10298 GNDA.n6799 GNDA.t146 65.8183
R10299 GNDA.n6806 GNDA.t146 65.8183
R10300 GNDA.n6640 GNDA.t146 65.8183
R10301 GNDA.t181 GNDA.n5662 65.8183
R10302 GNDA.t181 GNDA.n5661 65.8183
R10303 GNDA.t181 GNDA.n5660 65.8183
R10304 GNDA.t181 GNDA.n5659 65.8183
R10305 GNDA.t181 GNDA.n5650 65.8183
R10306 GNDA.t181 GNDA.n5657 65.8183
R10307 GNDA.t181 GNDA.n5647 65.8183
R10308 GNDA.t181 GNDA.n5658 65.8183
R10309 GNDA.t181 GNDA.n5656 65.8183
R10310 GNDA.t181 GNDA.n5654 65.8183
R10311 GNDA.t181 GNDA.n5653 65.8183
R10312 GNDA.t181 GNDA.n5652 65.8183
R10313 GNDA.n5746 GNDA.t181 65.8183
R10314 GNDA.t181 GNDA.n5649 65.8183
R10315 GNDA.t181 GNDA.n5648 65.8183
R10316 GNDA.t181 GNDA.n5646 65.8183
R10317 GNDA.t157 GNDA.n5472 65.8183
R10318 GNDA.t157 GNDA.n5471 65.8183
R10319 GNDA.t157 GNDA.n5470 65.8183
R10320 GNDA.t157 GNDA.n5469 65.8183
R10321 GNDA.t157 GNDA.n5460 65.8183
R10322 GNDA.t157 GNDA.n5467 65.8183
R10323 GNDA.t157 GNDA.n5457 65.8183
R10324 GNDA.t157 GNDA.n5468 65.8183
R10325 GNDA.t157 GNDA.n5466 65.8183
R10326 GNDA.t157 GNDA.n5465 65.8183
R10327 GNDA.t157 GNDA.n5464 65.8183
R10328 GNDA.t157 GNDA.n5463 65.8183
R10329 GNDA.t157 GNDA.n5461 65.8183
R10330 GNDA.t157 GNDA.n5459 65.8183
R10331 GNDA.t157 GNDA.n5458 65.8183
R10332 GNDA.n6059 GNDA.t157 65.8183
R10333 GNDA.t193 GNDA.n5982 65.8183
R10334 GNDA.t193 GNDA.n5905 65.8183
R10335 GNDA.t193 GNDA.n5904 65.8183
R10336 GNDA.t193 GNDA.n5903 65.8183
R10337 GNDA.t193 GNDA.n5894 65.8183
R10338 GNDA.t193 GNDA.n5901 65.8183
R10339 GNDA.t193 GNDA.n5892 65.8183
R10340 GNDA.t193 GNDA.n5902 65.8183
R10341 GNDA.t193 GNDA.n5900 65.8183
R10342 GNDA.t193 GNDA.n5899 65.8183
R10343 GNDA.t193 GNDA.n5898 65.8183
R10344 GNDA.t193 GNDA.n5897 65.8183
R10345 GNDA.t193 GNDA.n5895 65.8183
R10346 GNDA.t193 GNDA.n5893 65.8183
R10347 GNDA.n5983 GNDA.t193 65.8183
R10348 GNDA.t193 GNDA.n5887 65.8183
R10349 GNDA.n6720 GNDA.t167 65.8183
R10350 GNDA.n6726 GNDA.t167 65.8183
R10351 GNDA.n6728 GNDA.t167 65.8183
R10352 GNDA.n6734 GNDA.t167 65.8183
R10353 GNDA.n6704 GNDA.t167 65.8183
R10354 GNDA.n6710 GNDA.t167 65.8183
R10355 GNDA.n6712 GNDA.t167 65.8183
R10356 GNDA.n6718 GNDA.t167 65.8183
R10357 GNDA.n6688 GNDA.t167 65.8183
R10358 GNDA.n6687 GNDA.t167 65.8183
R10359 GNDA.n6695 GNDA.t167 65.8183
R10360 GNDA.n6682 GNDA.t167 65.8183
R10361 GNDA.n7026 GNDA.t167 65.8183
R10362 GNDA.n7023 GNDA.t167 65.8183
R10363 GNDA.n6755 GNDA.t167 65.8183
R10364 GNDA.n6753 GNDA.t167 65.8183
R10365 GNDA.t182 GNDA.n19 65.8183
R10366 GNDA.t182 GNDA.n18 65.8183
R10367 GNDA.t182 GNDA.n17 65.8183
R10368 GNDA.t182 GNDA.n16 65.8183
R10369 GNDA.t182 GNDA.n7 65.8183
R10370 GNDA.t182 GNDA.n14 65.8183
R10371 GNDA.t182 GNDA.n5 65.8183
R10372 GNDA.t182 GNDA.n15 65.8183
R10373 GNDA.t182 GNDA.n13 65.8183
R10374 GNDA.t182 GNDA.n12 65.8183
R10375 GNDA.t182 GNDA.n11 65.8183
R10376 GNDA.t182 GNDA.n10 65.8183
R10377 GNDA.t182 GNDA.n8 65.8183
R10378 GNDA.n7489 GNDA.t182 65.8183
R10379 GNDA.t182 GNDA.n6 65.8183
R10380 GNDA.t182 GNDA.n4 65.8183
R10381 GNDA.n6910 GNDA.t327 62.3509
R10382 GNDA.n6842 GNDA.t249 62.3509
R10383 GNDA.n3388 GNDA.t218 62.2505
R10384 GNDA.n3384 GNDA.t200 62.2505
R10385 GNDA.n1730 GNDA.t233 62.2505
R10386 GNDA.n1725 GNDA.t209 62.2505
R10387 GNDA.n3396 GNDA.t236 62.2505
R10388 GNDA.n5309 GNDA.t224 62.2505
R10389 GNDA.n1734 GNDA.t166 62.2505
R10390 GNDA.n1740 GNDA.t163 62.2505
R10391 GNDA.n1754 GNDA.t177 62.2505
R10392 GNDA.n1745 GNDA.t170 62.2505
R10393 GNDA.n3392 GNDA.t212 62.2505
R10394 GNDA.n3382 GNDA.t185 62.2505
R10395 GNDA.n6955 GNDA.n5348 61.2758
R10396 GNDA.n6936 GNDA.n5365 61.2758
R10397 GNDA.n5001 GNDA.n5000 59.2425
R10398 GNDA.n5003 GNDA.n5002 59.2425
R10399 GNDA.n658 GNDA.n319 59.2425
R10400 GNDA.n2107 GNDA.n316 59.2425
R10401 GNDA.t147 GNDA.n6441 57.8461
R10402 GNDA.t192 GNDA.n6536 57.8461
R10403 GNDA.t144 GNDA.n6976 57.8461
R10404 GNDA.n6639 GNDA.t146 57.8461
R10405 GNDA.t181 GNDA.n5745 57.8461
R10406 GNDA.t157 GNDA.n6058 57.8461
R10407 GNDA.t193 GNDA.n5886 57.8461
R10408 GNDA.n6736 GNDA.t167 57.8461
R10409 GNDA.t182 GNDA.n7488 57.8461
R10410 GNDA.n1750 GNDA.t124 57.4383
R10411 GNDA.n6646 GNDA.n6645 56.9758
R10412 GNDA.n5386 GNDA.n5348 56.9758
R10413 GNDA.n6939 GNDA.n6936 56.9758
R10414 GNDA.n7386 GNDA.n7316 56.3995
R10415 GNDA.n5756 GNDA.n5640 56.3995
R10416 GNDA.n6549 GNDA.n5414 56.3995
R10417 GNDA.n6573 GNDA.n6572 56.3995
R10418 GNDA.n7004 GNDA.n306 56.3995
R10419 GNDA.n7004 GNDA.n7003 56.3995
R10420 GNDA.n5757 GNDA.n5756 56.3995
R10421 GNDA.n7387 GNDA.n7386 56.3995
R10422 GNDA.n6572 GNDA.n5403 56.3995
R10423 GNDA.n5881 GNDA.n5421 56.3995
R10424 GNDA.n6547 GNDA.n5414 56.3995
R10425 GNDA.t313 GNDA.n6910 55.9008
R10426 GNDA.t142 GNDA.n6842 55.9008
R10427 GNDA.t244 GNDA.n7017 55.9008
R10428 GNDA.t192 GNDA.n6333 55.2026
R10429 GNDA.t147 GNDA.n6377 55.2026
R10430 GNDA.t144 GNDA.n5331 55.2026
R10431 GNDA.n6604 GNDA.t146 55.2026
R10432 GNDA.t181 GNDA.n5651 55.2026
R10433 GNDA.t157 GNDA.n5462 55.2026
R10434 GNDA.t193 GNDA.n5896 55.2026
R10435 GNDA.n6702 GNDA.t167 55.2026
R10436 GNDA.t182 GNDA.n9 55.2026
R10437 GNDA.n1747 GNDA.n315 55.0564
R10438 GNDA.n6518 GNDA.n6339 53.3664
R10439 GNDA.n6514 GNDA.n6328 53.3664
R10440 GNDA.n6510 GNDA.n6338 53.3664
R10441 GNDA.n6506 GNDA.n6331 53.3664
R10442 GNDA.n6495 GNDA.n6334 53.3664
R10443 GNDA.n6491 GNDA.n6335 53.3664
R10444 GNDA.n6487 GNDA.n6336 53.3664
R10445 GNDA.n6483 GNDA.n6337 53.3664
R10446 GNDA.n6538 GNDA.n6537 53.3664
R10447 GNDA.n6460 GNDA.n6329 53.3664
R10448 GNDA.n6468 GNDA.n6330 53.3664
R10449 GNDA.n6475 GNDA.n6332 53.3664
R10450 GNDA.n6522 GNDA.n6343 53.3664
R10451 GNDA.n6523 GNDA.n6342 53.3664
R10452 GNDA.n6527 GNDA.n6341 53.3664
R10453 GNDA.n6531 GNDA.n6340 53.3664
R10454 GNDA.n6519 GNDA.n6343 53.3664
R10455 GNDA.n6526 GNDA.n6342 53.3664
R10456 GNDA.n6530 GNDA.n6341 53.3664
R10457 GNDA.n6534 GNDA.n6340 53.3664
R10458 GNDA.n6503 GNDA.n6331 53.3664
R10459 GNDA.n6507 GNDA.n6338 53.3664
R10460 GNDA.n6511 GNDA.n6328 53.3664
R10461 GNDA.n6515 GNDA.n6339 53.3664
R10462 GNDA.n6486 GNDA.n6337 53.3664
R10463 GNDA.n6490 GNDA.n6336 53.3664
R10464 GNDA.n6494 GNDA.n6335 53.3664
R10465 GNDA.n6498 GNDA.n6334 53.3664
R10466 GNDA.n6423 GNDA.n6385 53.3664
R10467 GNDA.n6419 GNDA.n6349 53.3664
R10468 GNDA.n6415 GNDA.n6384 53.3664
R10469 GNDA.n6411 GNDA.n6352 53.3664
R10470 GNDA.n6400 GNDA.n6378 53.3664
R10471 GNDA.n6396 GNDA.n6379 53.3664
R10472 GNDA.n6392 GNDA.n6380 53.3664
R10473 GNDA.n6383 GNDA.n6382 53.3664
R10474 GNDA.n6443 GNDA.n6442 53.3664
R10475 GNDA.n6359 GNDA.n6350 53.3664
R10476 GNDA.n6367 GNDA.n6351 53.3664
R10477 GNDA.n6376 GNDA.n6375 53.3664
R10478 GNDA.n6427 GNDA.n6389 53.3664
R10479 GNDA.n6428 GNDA.n6388 53.3664
R10480 GNDA.n6432 GNDA.n6387 53.3664
R10481 GNDA.n6436 GNDA.n6386 53.3664
R10482 GNDA.n6424 GNDA.n6389 53.3664
R10483 GNDA.n6431 GNDA.n6388 53.3664
R10484 GNDA.n6435 GNDA.n6387 53.3664
R10485 GNDA.n6439 GNDA.n6386 53.3664
R10486 GNDA.n6408 GNDA.n6352 53.3664
R10487 GNDA.n6412 GNDA.n6384 53.3664
R10488 GNDA.n6416 GNDA.n6349 53.3664
R10489 GNDA.n6420 GNDA.n6385 53.3664
R10490 GNDA.n6391 GNDA.n6383 53.3664
R10491 GNDA.n6395 GNDA.n6380 53.3664
R10492 GNDA.n6399 GNDA.n6379 53.3664
R10493 GNDA.n6403 GNDA.n6378 53.3664
R10494 GNDA.n6381 GNDA.n6376 53.3664
R10495 GNDA.n6353 GNDA.n6351 53.3664
R10496 GNDA.n6366 GNDA.n6350 53.3664
R10497 GNDA.n6442 GNDA.n6348 53.3664
R10498 GNDA.n6482 GNDA.n6332 53.3664
R10499 GNDA.n6474 GNDA.n6330 53.3664
R10500 GNDA.n6467 GNDA.n6329 53.3664
R10501 GNDA.n6537 GNDA.n6327 53.3664
R10502 GNDA.n6885 GNDA.n5337 53.3664
R10503 GNDA.n6881 GNDA.n5327 53.3664
R10504 GNDA.n6877 GNDA.n5336 53.3664
R10505 GNDA.n6873 GNDA.n5329 53.3664
R10506 GNDA.n6862 GNDA.n5332 53.3664
R10507 GNDA.n6858 GNDA.n5333 53.3664
R10508 GNDA.n6854 GNDA.n5334 53.3664
R10509 GNDA.n6850 GNDA.n5335 53.3664
R10510 GNDA.n5343 GNDA.n5326 53.3664
R10511 GNDA.n6965 GNDA.n5328 53.3664
R10512 GNDA.n6978 GNDA.n6977 53.3664
R10513 GNDA.n6836 GNDA.n5330 53.3664
R10514 GNDA.n6889 GNDA.n5341 53.3664
R10515 GNDA.n6890 GNDA.n5340 53.3664
R10516 GNDA.n6894 GNDA.n5339 53.3664
R10517 GNDA.n6898 GNDA.n5338 53.3664
R10518 GNDA.n6886 GNDA.n5341 53.3664
R10519 GNDA.n6893 GNDA.n5340 53.3664
R10520 GNDA.n6897 GNDA.n5339 53.3664
R10521 GNDA.n6900 GNDA.n5338 53.3664
R10522 GNDA.n6870 GNDA.n5329 53.3664
R10523 GNDA.n6874 GNDA.n5336 53.3664
R10524 GNDA.n6878 GNDA.n5327 53.3664
R10525 GNDA.n6882 GNDA.n5337 53.3664
R10526 GNDA.n6853 GNDA.n5335 53.3664
R10527 GNDA.n6857 GNDA.n5334 53.3664
R10528 GNDA.n6861 GNDA.n5333 53.3664
R10529 GNDA.n6865 GNDA.n5332 53.3664
R10530 GNDA.n6849 GNDA.n5330 53.3664
R10531 GNDA.n6977 GNDA.n5325 53.3664
R10532 GNDA.n5328 GNDA.n5324 53.3664
R10533 GNDA.n6964 GNDA.n5326 53.3664
R10534 GNDA.n6621 GNDA.n6620 53.3664
R10535 GNDA.n6614 GNDA.n6582 53.3664
R10536 GNDA.n6613 GNDA.n6612 53.3664
R10537 GNDA.n6606 GNDA.n6584 53.3664
R10538 GNDA.n6599 GNDA.n6588 53.3664
R10539 GNDA.n6597 GNDA.n6596 53.3664
R10540 GNDA.n6592 GNDA.n6590 53.3664
R10541 GNDA.n6834 GNDA.n5397 53.3664
R10542 GNDA.n6817 GNDA.n6640 53.3664
R10543 GNDA.n6806 GNDA.n6805 53.3664
R10544 GNDA.n6803 GNDA.n6799 53.3664
R10545 GNDA.n6832 GNDA.n6831 53.3664
R10546 GNDA.n6622 GNDA.n6580 53.3664
R10547 GNDA.n6628 GNDA.n6627 53.3664
R10548 GNDA.n6631 GNDA.n6630 53.3664
R10549 GNDA.n6636 GNDA.n6635 53.3664
R10550 GNDA.n6623 GNDA.n6622 53.3664
R10551 GNDA.n6629 GNDA.n6628 53.3664
R10552 GNDA.n6630 GNDA.n6578 53.3664
R10553 GNDA.n6637 GNDA.n6636 53.3664
R10554 GNDA.n6607 GNDA.n6606 53.3664
R10555 GNDA.n6612 GNDA.n6611 53.3664
R10556 GNDA.n6615 GNDA.n6614 53.3664
R10557 GNDA.n6620 GNDA.n6619 53.3664
R10558 GNDA.n6591 GNDA.n5397 53.3664
R10559 GNDA.n6590 GNDA.n6589 53.3664
R10560 GNDA.n6598 GNDA.n6597 53.3664
R10561 GNDA.n6588 GNDA.n6586 53.3664
R10562 GNDA.n6833 GNDA.n6832 53.3664
R10563 GNDA.n6799 GNDA.n5398 53.3664
R10564 GNDA.n6807 GNDA.n6806 53.3664
R10565 GNDA.n6804 GNDA.n6640 53.3664
R10566 GNDA.n5698 GNDA.n5658 53.3664
R10567 GNDA.n5694 GNDA.n5647 53.3664
R10568 GNDA.n5690 GNDA.n5657 53.3664
R10569 GNDA.n5686 GNDA.n5650 53.3664
R10570 GNDA.n5675 GNDA.n5652 53.3664
R10571 GNDA.n5671 GNDA.n5653 53.3664
R10572 GNDA.n5667 GNDA.n5654 53.3664
R10573 GNDA.n5656 GNDA.n5655 53.3664
R10574 GNDA.n5664 GNDA.n5646 53.3664
R10575 GNDA.n5733 GNDA.n5648 53.3664
R10576 GNDA.n5726 GNDA.n5649 53.3664
R10577 GNDA.n5747 GNDA.n5746 53.3664
R10578 GNDA.n5702 GNDA.n5662 53.3664
R10579 GNDA.n5703 GNDA.n5661 53.3664
R10580 GNDA.n5707 GNDA.n5660 53.3664
R10581 GNDA.n5711 GNDA.n5659 53.3664
R10582 GNDA.n5699 GNDA.n5662 53.3664
R10583 GNDA.n5706 GNDA.n5661 53.3664
R10584 GNDA.n5710 GNDA.n5660 53.3664
R10585 GNDA.n5713 GNDA.n5659 53.3664
R10586 GNDA.n5683 GNDA.n5650 53.3664
R10587 GNDA.n5687 GNDA.n5657 53.3664
R10588 GNDA.n5691 GNDA.n5647 53.3664
R10589 GNDA.n5695 GNDA.n5658 53.3664
R10590 GNDA.n5666 GNDA.n5656 53.3664
R10591 GNDA.n5670 GNDA.n5654 53.3664
R10592 GNDA.n5674 GNDA.n5653 53.3664
R10593 GNDA.n5678 GNDA.n5652 53.3664
R10594 GNDA.n5746 GNDA.n5645 53.3664
R10595 GNDA.n5649 GNDA.n5644 53.3664
R10596 GNDA.n5725 GNDA.n5648 53.3664
R10597 GNDA.n5732 GNDA.n5646 53.3664
R10598 GNDA.n6040 GNDA.n5468 53.3664
R10599 GNDA.n6036 GNDA.n5457 53.3664
R10600 GNDA.n6032 GNDA.n5467 53.3664
R10601 GNDA.n6028 GNDA.n5460 53.3664
R10602 GNDA.n6017 GNDA.n5463 53.3664
R10603 GNDA.n6013 GNDA.n5464 53.3664
R10604 GNDA.n6009 GNDA.n5465 53.3664
R10605 GNDA.n6005 GNDA.n5466 53.3664
R10606 GNDA.n6060 GNDA.n6059 53.3664
R10607 GNDA.n5504 GNDA.n5458 53.3664
R10608 GNDA.n5500 GNDA.n5459 53.3664
R10609 GNDA.n5493 GNDA.n5461 53.3664
R10610 GNDA.n6044 GNDA.n5472 53.3664
R10611 GNDA.n6045 GNDA.n5471 53.3664
R10612 GNDA.n6049 GNDA.n5470 53.3664
R10613 GNDA.n6053 GNDA.n5469 53.3664
R10614 GNDA.n6041 GNDA.n5472 53.3664
R10615 GNDA.n6048 GNDA.n5471 53.3664
R10616 GNDA.n6052 GNDA.n5470 53.3664
R10617 GNDA.n6056 GNDA.n5469 53.3664
R10618 GNDA.n6025 GNDA.n5460 53.3664
R10619 GNDA.n6029 GNDA.n5467 53.3664
R10620 GNDA.n6033 GNDA.n5457 53.3664
R10621 GNDA.n6037 GNDA.n5468 53.3664
R10622 GNDA.n6008 GNDA.n5466 53.3664
R10623 GNDA.n6012 GNDA.n5465 53.3664
R10624 GNDA.n6016 GNDA.n5464 53.3664
R10625 GNDA.n6020 GNDA.n5463 53.3664
R10626 GNDA.n6004 GNDA.n5461 53.3664
R10627 GNDA.n5492 GNDA.n5459 53.3664
R10628 GNDA.n5501 GNDA.n5458 53.3664
R10629 GNDA.n6059 GNDA.n5456 53.3664
R10630 GNDA.n5965 GNDA.n5902 53.3664
R10631 GNDA.n5962 GNDA.n5892 53.3664
R10632 GNDA.n5958 GNDA.n5901 53.3664
R10633 GNDA.n5954 GNDA.n5894 53.3664
R10634 GNDA.n5943 GNDA.n5897 53.3664
R10635 GNDA.n5939 GNDA.n5898 53.3664
R10636 GNDA.n5935 GNDA.n5899 53.3664
R10637 GNDA.n5931 GNDA.n5900 53.3664
R10638 GNDA.n5991 GNDA.n5887 53.3664
R10639 GNDA.n5984 GNDA.n5983 53.3664
R10640 GNDA.n5916 GNDA.n5893 53.3664
R10641 GNDA.n5923 GNDA.n5895 53.3664
R10642 GNDA.n5982 GNDA.n5981 53.3664
R10643 GNDA.n5907 GNDA.n5905 53.3664
R10644 GNDA.n5976 GNDA.n5904 53.3664
R10645 GNDA.n5972 GNDA.n5903 53.3664
R10646 GNDA.n5982 GNDA.n5906 53.3664
R10647 GNDA.n5977 GNDA.n5905 53.3664
R10648 GNDA.n5973 GNDA.n5904 53.3664
R10649 GNDA.n5969 GNDA.n5903 53.3664
R10650 GNDA.n5951 GNDA.n5894 53.3664
R10651 GNDA.n5955 GNDA.n5901 53.3664
R10652 GNDA.n5959 GNDA.n5892 53.3664
R10653 GNDA.n5963 GNDA.n5902 53.3664
R10654 GNDA.n5934 GNDA.n5900 53.3664
R10655 GNDA.n5938 GNDA.n5899 53.3664
R10656 GNDA.n5942 GNDA.n5898 53.3664
R10657 GNDA.n5946 GNDA.n5897 53.3664
R10658 GNDA.n5930 GNDA.n5895 53.3664
R10659 GNDA.n5922 GNDA.n5893 53.3664
R10660 GNDA.n5983 GNDA.n5891 53.3664
R10661 GNDA.n5890 GNDA.n5887 53.3664
R10662 GNDA.n6719 GNDA.n6718 53.3664
R10663 GNDA.n6712 GNDA.n6676 53.3664
R10664 GNDA.n6711 GNDA.n6710 53.3664
R10665 GNDA.n6704 GNDA.n6678 53.3664
R10666 GNDA.n6697 GNDA.n6682 53.3664
R10667 GNDA.n6695 GNDA.n6694 53.3664
R10668 GNDA.n6690 GNDA.n6687 53.3664
R10669 GNDA.n6688 GNDA.n292 53.3664
R10670 GNDA.n6753 GNDA.n6752 53.3664
R10671 GNDA.n6756 GNDA.n6755 53.3664
R10672 GNDA.n7023 GNDA.n7022 53.3664
R10673 GNDA.n7026 GNDA.n7025 53.3664
R10674 GNDA.n6720 GNDA.n6674 53.3664
R10675 GNDA.n6726 GNDA.n6725 53.3664
R10676 GNDA.n6729 GNDA.n6728 53.3664
R10677 GNDA.n6734 GNDA.n6733 53.3664
R10678 GNDA.n6721 GNDA.n6720 53.3664
R10679 GNDA.n6727 GNDA.n6726 53.3664
R10680 GNDA.n6728 GNDA.n6672 53.3664
R10681 GNDA.n6735 GNDA.n6734 53.3664
R10682 GNDA.n6705 GNDA.n6704 53.3664
R10683 GNDA.n6710 GNDA.n6709 53.3664
R10684 GNDA.n6713 GNDA.n6712 53.3664
R10685 GNDA.n6718 GNDA.n6717 53.3664
R10686 GNDA.n6689 GNDA.n6688 53.3664
R10687 GNDA.n6687 GNDA.n6683 53.3664
R10688 GNDA.n6696 GNDA.n6695 53.3664
R10689 GNDA.n6682 GNDA.n6680 53.3664
R10690 GNDA.n7027 GNDA.n7026 53.3664
R10691 GNDA.n7024 GNDA.n7023 53.3664
R10692 GNDA.n6755 GNDA.n295 53.3664
R10693 GNDA.n6754 GNDA.n6753 53.3664
R10694 GNDA.n7335 GNDA.n15 53.3664
R10695 GNDA.n7339 GNDA.n5 53.3664
R10696 GNDA.n7343 GNDA.n14 53.3664
R10697 GNDA.n7347 GNDA.n7 53.3664
R10698 GNDA.n7358 GNDA.n10 53.3664
R10699 GNDA.n7362 GNDA.n11 53.3664
R10700 GNDA.n7366 GNDA.n12 53.3664
R10701 GNDA.n7370 GNDA.n13 53.3664
R10702 GNDA.n21 GNDA.n4 53.3664
R10703 GNDA.n37 GNDA.n6 53.3664
R10704 GNDA.n7490 GNDA.n7489 53.3664
R10705 GNDA.n7377 GNDA.n8 53.3664
R10706 GNDA.n7331 GNDA.n19 53.3664
R10707 GNDA.n7330 GNDA.n18 53.3664
R10708 GNDA.n7326 GNDA.n17 53.3664
R10709 GNDA.n7322 GNDA.n16 53.3664
R10710 GNDA.n7334 GNDA.n19 53.3664
R10711 GNDA.n7327 GNDA.n18 53.3664
R10712 GNDA.n7323 GNDA.n17 53.3664
R10713 GNDA.n7319 GNDA.n16 53.3664
R10714 GNDA.n7350 GNDA.n7 53.3664
R10715 GNDA.n7346 GNDA.n14 53.3664
R10716 GNDA.n7342 GNDA.n5 53.3664
R10717 GNDA.n7338 GNDA.n15 53.3664
R10718 GNDA.n7367 GNDA.n13 53.3664
R10719 GNDA.n7363 GNDA.n12 53.3664
R10720 GNDA.n7359 GNDA.n11 53.3664
R10721 GNDA.n7355 GNDA.n10 53.3664
R10722 GNDA.n7371 GNDA.n8 53.3664
R10723 GNDA.n7489 GNDA.n3 53.3664
R10724 GNDA.n6 GNDA.n2 53.3664
R10725 GNDA.n36 GNDA.n4 53.3664
R10726 GNDA.t247 GNDA.n6811 51.6008
R10727 GNDA.t187 GNDA.n6970 51.6008
R10728 GNDA.n6743 GNDA.t30 51.6008
R10729 GNDA.n6994 GNDA.t283 50.6082
R10730 GNDA.n6811 GNDA.t145 50.5258
R10731 GNDA.t274 GNDA.n5371 50.5258
R10732 GNDA.n6912 GNDA.t281 49.4508
R10733 GNDA.n5516 GNDA.t145 47.6748
R10734 GNDA.n5310 GNDA.t223 47.5205
R10735 GNDA.n3395 GNDA.t235 47.5205
R10736 GNDA.n5382 GNDA.n5365 47.3008
R10737 GNDA.n6922 GNDA.n5386 46.2258
R10738 GNDA.n7017 GNDA.t145 46.2258
R10739 GNDA.n6971 GNDA.t187 45.1508
R10740 GNDA.t30 GNDA.n6742 45.1508
R10741 GNDA.n6097 GNDA.t145 44.3072
R10742 GNDA.n6959 GNDA.t97 44.0757
R10743 GNDA.n6911 GNDA.t313 40.8507
R10744 GNDA.n6983 GNDA.n6982 40.8507
R10745 GNDA.n6844 GNDA.t142 40.8507
R10746 GNDA.n1735 GNDA.t239 40.4338
R10747 GNDA.n1738 GNDA.t160 40.4338
R10748 GNDA.n5306 GNDA.t221 40.4338
R10749 GNDA.n321 GNDA.t174 40.4338
R10750 GNDA.n5780 GNDA.t2 40.1125
R10751 GNDA.n6645 GNDA.n5402 39.7757
R10752 GNDA.n6812 GNDA.t125 39.7757
R10753 GNDA.t323 GNDA.n5319 39.5367
R10754 GNDA.t119 GNDA.t111 38.7205
R10755 GNDA.t120 GNDA.t108 38.7205
R10756 GNDA.t115 GNDA.t109 38.7205
R10757 GNDA.t114 GNDA.t103 38.7205
R10758 GNDA.t112 GNDA.t121 38.7205
R10759 GNDA.t223 GNDA.t263 38.7205
R10760 GNDA.t263 GNDA.t25 38.7205
R10761 GNDA.t25 GNDA.t256 38.7205
R10762 GNDA.t232 GNDA.t40 38.7205
R10763 GNDA.t78 GNDA.t232 38.7205
R10764 GNDA.t301 GNDA.t199 38.7205
R10765 GNDA.t55 GNDA.t290 38.7205
R10766 GNDA.t235 GNDA.t55 38.7205
R10767 GNDA.t93 GNDA.t140 38.7205
R10768 GNDA.t316 GNDA.t94 38.7205
R10769 GNDA.t96 GNDA.t17 38.7205
R10770 GNDA.t92 GNDA.t320 38.7205
R10771 GNDA.t329 GNDA.t95 38.7205
R10772 GNDA.t281 GNDA.t155 37.6257
R10773 GNDA.t179 GNDA.t274 37.6257
R10774 GNDA.n5284 GNDA.n5283 37.5297
R10775 GNDA.n5286 GNDA.n5285 37.5297
R10776 GNDA.n5288 GNDA.n5287 37.5297
R10777 GNDA.n5290 GNDA.n5289 37.5297
R10778 GNDA.n5292 GNDA.n5291 37.5297
R10779 GNDA.n5294 GNDA.n5293 37.5297
R10780 GNDA.n5296 GNDA.n5295 37.5297
R10781 GNDA.n5298 GNDA.n5297 37.5297
R10782 GNDA.n5300 GNDA.n5299 37.5297
R10783 GNDA.n5302 GNDA.n5301 37.5297
R10784 GNDA.n5304 GNDA.n5303 37.5297
R10785 GNDA.t202 GNDA.t205 36.9605
R10786 GNDA.t226 GNDA.t190 36.9605
R10787 GNDA.n3383 GNDA.t39 36.9605
R10788 GNDA.t241 GNDA.t229 36.9605
R10789 GNDA.t214 GNDA.t152 36.9605
R10790 GNDA.n7018 GNDA.t26 35.4757
R10791 GNDA.n1774 GNDA.n1773 34.5991
R10792 GNDA.n6319 GNDA.n6260 34.4263
R10793 GNDA.n6319 GNDA.n6318 34.4263
R10794 GNDA.n6318 GNDA.n6317 34.4263
R10795 GNDA.n6317 GNDA.n6261 34.4263
R10796 GNDA.n6311 GNDA.n6261 34.4263
R10797 GNDA.n6310 GNDA.n6309 34.4263
R10798 GNDA.n6309 GNDA.n6265 34.4263
R10799 GNDA.n6303 GNDA.n6265 34.4263
R10800 GNDA.n6303 GNDA.n6302 34.4263
R10801 GNDA.n6302 GNDA.n77 34.4263
R10802 GNDA.n7462 GNDA.n78 34.4263
R10803 GNDA.n7456 GNDA.n78 34.4263
R10804 GNDA.n7456 GNDA.n7455 34.4263
R10805 GNDA.n7455 GNDA.n7454 34.4263
R10806 GNDA.n7454 GNDA.n84 34.4263
R10807 GNDA.n7447 GNDA.n7446 34.4263
R10808 GNDA.n7446 GNDA.n7445 34.4263
R10809 GNDA.n7445 GNDA.n7240 34.4263
R10810 GNDA.n7439 GNDA.n7240 34.4263
R10811 GNDA.n7439 GNDA.n7438 34.4263
R10812 GNDA.n7436 GNDA.n7246 34.4263
R10813 GNDA.n7430 GNDA.n7246 34.4263
R10814 GNDA.n7430 GNDA.n7429 34.4263
R10815 GNDA.n7429 GNDA.n7428 34.4263
R10816 GNDA.n7428 GNDA.n7297 34.4263
R10817 GNDA.n7422 GNDA.n7421 34.4263
R10818 GNDA.n7421 GNDA.n7420 34.4263
R10819 GNDA.n7420 GNDA.n7301 34.4263
R10820 GNDA.n7414 GNDA.n7301 34.4263
R10821 GNDA.n7414 GNDA.n7413 34.4263
R10822 GNDA.t249 GNDA.n6841 34.4007
R10823 GNDA.n6792 GNDA.n6781 33.0531
R10824 GNDA.t145 GNDA.n26 32.9056
R10825 GNDA.n5446 GNDA.t145 32.9056
R10826 GNDA.n6777 GNDA.n6776 32.3969
R10827 GNDA.n6957 GNDA.n6955 32.2507
R10828 GNDA.n6939 GNDA.n5363 32.2507
R10829 GNDA.n3397 GNDA.n3396 31.5738
R10830 GNDA.n6912 GNDA.t13 31.1757
R10831 GNDA.n3402 GNDA.t153 31.1255
R10832 GNDA.n3399 GNDA.t242 31.1255
R10833 GNDA.n5312 GNDA.t227 31.1255
R10834 GNDA.n5317 GNDA.t206 31.1255
R10835 GNDA.t44 GNDA.t126 30.9902
R10836 GNDA.t257 GNDA.n6969 30.1007
R10837 GNDA.t80 GNDA.n5371 30.1007
R10838 GNDA.t288 GNDA.t119 29.9205
R10839 GNDA.t121 GNDA.t62 29.9205
R10840 GNDA.n5307 GNDA.t9 29.9205
R10841 GNDA.t37 GNDA.n3390 29.9205
R10842 GNDA.n3394 GNDA.t129 29.9205
R10843 GNDA.t140 GNDA.t47 29.9205
R10844 GNDA.t127 GNDA.t329 29.9205
R10845 GNDA.n5309 GNDA.n5308 29.8672
R10846 GNDA.n1755 GNDA.n1754 29.8672
R10847 GNDA.n1745 GNDA.n1744 29.8672
R10848 GNDA.t332 GNDA.t86 29.5889
R10849 GNDA.n5758 GNDA.t145 29.1014
R10850 GNDA.n6774 GNDA.n6762 29.0257
R10851 GNDA.n1750 GNDA.n575 28.1605
R10852 GNDA.n6520 GNDA.n6517 27.5561
R10853 GNDA.n6425 GNDA.n6422 27.5561
R10854 GNDA.n6887 GNDA.n6884 27.5561
R10855 GNDA.n6624 GNDA.n6581 27.5561
R10856 GNDA.n5700 GNDA.n5697 27.5561
R10857 GNDA.n6042 GNDA.n6039 27.5561
R10858 GNDA.n5967 GNDA.n5966 27.5561
R10859 GNDA.n6722 GNDA.n6675 27.5561
R10860 GNDA.n7336 GNDA.n7333 27.5561
R10861 GNDA.t16 GNDA.t325 27.2873
R10862 GNDA.t137 GNDA.t327 26.8757
R10863 GNDA.t4 GNDA.t0 26.8757
R10864 GNDA.t124 GNDA.t43 26.7157
R10865 GNDA.t73 GNDA.t324 26.7157
R10866 GNDA.n6501 GNDA.n6500 26.6672
R10867 GNDA.n6406 GNDA.n6405 26.6672
R10868 GNDA.n6868 GNDA.n6867 26.6672
R10869 GNDA.n6602 GNDA.n6585 26.6672
R10870 GNDA.n5681 GNDA.n5680 26.6672
R10871 GNDA.n6023 GNDA.n6022 26.6672
R10872 GNDA.n5949 GNDA.n5948 26.6672
R10873 GNDA.n6700 GNDA.n6679 26.6672
R10874 GNDA.n7353 GNDA.n7352 26.6672
R10875 GNDA.t205 GNDA.n316 26.4005
R10876 GNDA.n319 GNDA.t226 26.4005
R10877 GNDA.n5002 GNDA.t241 26.4005
R10878 GNDA.t152 GNDA.n5001 26.4005
R10879 GNDA.n6994 GNDA.n309 25.8006
R10880 GNDA.t310 GNDA.t84 25.5077
R10881 GNDA.t102 GNDA.t323 25.5077
R10882 GNDA.n6784 GNDA.n6783 25.3679
R10883 GNDA.t27 GNDA.t149 25.0134
R10884 GNDA.t23 GNDA.t27 25.0134
R10885 GNDA.t32 GNDA.t23 25.0134
R10886 GNDA.n6795 GNDA.n6794 24.7256
R10887 GNDA.t15 GNDA.t68 24.1211
R10888 GNDA.t68 GNDA.t306 24.1211
R10889 GNDA.n285 GNDA.t261 24.0005
R10890 GNDA.n285 GNDA.t136 24.0005
R10891 GNDA.n284 GNDA.t5 24.0005
R10892 GNDA.n284 GNDA.t294 24.0005
R10893 GNDA.n283 GNDA.t81 24.0005
R10894 GNDA.n283 GNDA.t31 24.0005
R10895 GNDA.n280 GNDA.t59 24.0005
R10896 GNDA.n280 GNDA.t250 24.0005
R10897 GNDA.n279 GNDA.t258 24.0005
R10898 GNDA.n279 GNDA.t287 24.0005
R10899 GNDA.n276 GNDA.t314 24.0005
R10900 GNDA.n276 GNDA.t14 24.0005
R10901 GNDA.n275 GNDA.t252 24.0005
R10902 GNDA.n275 GNDA.t328 24.0005
R10903 GNDA.n274 GNDA.t53 24.0005
R10904 GNDA.n274 GNDA.t335 24.0005
R10905 GNDA.n271 GNDA.t33 24.0005
R10906 GNDA.n271 GNDA.t196 24.0005
R10907 GNDA.n270 GNDA.t28 24.0005
R10908 GNDA.n270 GNDA.t24 24.0005
R10909 GNDA.n7412 GNDA.n7305 23.5958
R10910 GNDA.n7406 GNDA.n7305 23.5958
R10911 GNDA.n7406 GNDA.n7405 23.5958
R10912 GNDA.n7405 GNDA.n7404 23.5958
R10913 GNDA.n7404 GNDA.n7309 23.5958
R10914 GNDA.n7398 GNDA.n7397 23.5958
R10915 GNDA.n7397 GNDA.n7396 23.5958
R10916 GNDA.n7396 GNDA.n7313 23.5958
R10917 GNDA.n7390 GNDA.n7313 23.5958
R10918 GNDA.n7390 GNDA.n7389 23.5958
R10919 GNDA.n7389 GNDA.n7388 23.5958
R10920 GNDA.n7388 GNDA.t322 23.5958
R10921 GNDA.n5780 GNDA.n5779 23.5958
R10922 GNDA.n5779 GNDA.n5778 23.5958
R10923 GNDA.n5778 GNDA.n5630 23.5958
R10924 GNDA.n5772 GNDA.n5630 23.5958
R10925 GNDA.n5772 GNDA.n5771 23.5958
R10926 GNDA.n5768 GNDA.n5767 23.5958
R10927 GNDA.n5767 GNDA.n5766 23.5958
R10928 GNDA.n5766 GNDA.n5636 23.5958
R10929 GNDA.n5760 GNDA.n5636 23.5958
R10930 GNDA.n5760 GNDA.n5759 23.5958
R10931 GNDA.n5759 GNDA.n5758 23.5958
R10932 GNDA.n6097 GNDA.n6096 23.5958
R10933 GNDA.n6096 GNDA.n6095 23.5958
R10934 GNDA.n6095 GNDA.n6086 23.5958
R10935 GNDA.n6089 GNDA.n6086 23.5958
R10936 GNDA.n6089 GNDA.n298 23.5958
R10937 GNDA.n7016 GNDA.n299 23.5958
R10938 GNDA.n7010 GNDA.n299 23.5958
R10939 GNDA.n7010 GNDA.n7009 23.5958
R10940 GNDA.n7009 GNDA.n7008 23.5958
R10941 GNDA.n7008 GNDA.n305 23.5958
R10942 GNDA.n7002 GNDA.n305 23.5958
R10943 GNDA.t264 GNDA.t120 22.8805
R10944 GNDA.t103 GNDA.t268 22.8805
R10945 GNDA.t90 GNDA.t60 22.8805
R10946 GNDA.t94 GNDA.t7 22.8805
R10947 GNDA.t99 GNDA.t92 22.8805
R10948 GNDA.n5318 GNDA.n316 21.1205
R10949 GNDA.n5311 GNDA.n319 21.1205
R10950 GNDA.t259 GNDA.t220 21.1205
R10951 GNDA.t262 GNDA.t49 21.1205
R10952 GNDA.t36 GNDA.t65 21.1205
R10953 GNDA.t308 GNDA.t297 21.1205
R10954 GNDA.t77 GNDA.t271 21.1205
R10955 GNDA.t273 GNDA.t304 21.1205
R10956 GNDA.t208 GNDA.t71 21.1205
R10957 GNDA.t138 GNDA.t217 21.1205
R10958 GNDA.t291 GNDA.t101 21.1205
R10959 GNDA.t337 GNDA.t295 21.1205
R10960 GNDA.t133 GNDA.t56 21.1205
R10961 GNDA.t311 GNDA.t254 21.1205
R10962 GNDA.t131 GNDA.t91 21.1205
R10963 GNDA.t266 GNDA.t255 21.1205
R10964 GNDA.t172 GNDA.t10 21.1205
R10965 GNDA.n5002 GNDA.n574 21.1205
R10966 GNDA.n5001 GNDA.n575 21.1205
R10967 GNDA.n7034 GNDA.n7033 20.8233
R10968 GNDA.n5364 GNDA.n282 20.8233
R10969 GNDA.n5362 GNDA.n281 20.8233
R10970 GNDA.n6956 GNDA.n278 20.8233
R10971 GNDA.n5385 GNDA.n277 20.8233
R10972 GNDA.n6647 GNDA.n273 20.8233
R10973 GNDA.n6644 GNDA.n272 20.8233
R10974 GNDA.n5407 GNDA.n269 20.8233
R10975 GNDA.n3417 GNDA.t319 19.7005
R10976 GNDA.n3417 GNDA.t285 19.7005
R10977 GNDA.n3415 GNDA.t18 19.7005
R10978 GNDA.n3415 GNDA.t85 19.7005
R10979 GNDA.n3413 GNDA.t35 19.7005
R10980 GNDA.n3413 GNDA.t317 19.7005
R10981 GNDA.n3411 GNDA.t318 19.7005
R10982 GNDA.n3411 GNDA.t74 19.7005
R10983 GNDA.n3409 GNDA.t330 19.7005
R10984 GNDA.n3409 GNDA.t331 19.7005
R10985 GNDA.n3408 GNDA.t278 19.7005
R10986 GNDA.n3408 GNDA.t6 19.7005
R10987 GNDA.n1787 GNDA.t105 19.7005
R10988 GNDA.n1787 GNDA.t277 19.7005
R10989 GNDA.n1789 GNDA.t113 19.7005
R10990 GNDA.n1789 GNDA.t116 19.7005
R10991 GNDA.n1791 GNDA.t104 19.7005
R10992 GNDA.n1791 GNDA.t122 19.7005
R10993 GNDA.n1793 GNDA.t117 19.7005
R10994 GNDA.n1793 GNDA.t107 19.7005
R10995 GNDA.n1795 GNDA.t118 19.7005
R10996 GNDA.n1795 GNDA.t106 19.7005
R10997 GNDA.n1797 GNDA.t276 19.7005
R10998 GNDA.n1797 GNDA.t110 19.7005
R10999 GNDA.n1737 GNDA.t78 19.3605
R11000 GNDA.n1737 GNDA.t39 19.3605
R11001 GNDA.t19 GNDA.n5408 19.3287
R11002 GNDA.n7450 GNDA.n86 18.5605
R11003 GNDA.n6311 GNDA.t145 17.9784
R11004 GNDA.t145 GNDA.n84 17.9784
R11005 GNDA.t145 GNDA.n7297 17.9784
R11006 GNDA.t220 GNDA.t9 17.6005
R11007 GNDA.t49 GNDA.t259 17.6005
R11008 GNDA.t65 GNDA.t262 17.6005
R11009 GNDA.t297 GNDA.t36 17.6005
R11010 GNDA.t271 GNDA.t308 17.6005
R11011 GNDA.t304 GNDA.t77 17.6005
R11012 GNDA.t71 GNDA.t273 17.6005
R11013 GNDA.t60 GNDA.t208 17.6005
R11014 GNDA.t255 GNDA.t131 17.6005
R11015 GNDA.t10 GNDA.t266 17.6005
R11016 GNDA.t129 GNDA.t172 17.6005
R11017 GNDA.n5783 GNDA.n5627 17.5843
R11018 GNDA.n6100 GNDA.n6083 17.5843
R11019 GNDA.n7410 GNDA.n7303 17.5843
R11020 GNDA.n6568 GNDA.n6322 16.9379
R11021 GNDA.n6252 GNDA.n6234 16.9379
R11022 GNDA.n5860 GNDA.n5515 16.9379
R11023 GNDA.n5524 GNDA.n65 16.7709
R11024 GNDA.n6210 GNDA.n5435 16.7709
R11025 GNDA.n7475 GNDA.n61 16.7709
R11026 GNDA.n6073 GNDA.n6072 16.7709
R11027 GNDA.t145 GNDA.n6310 16.4484
R11028 GNDA.n7447 GNDA.t145 16.4484
R11029 GNDA.n7422 GNDA.t145 16.4484
R11030 GNDA.t52 GNDA.t145 16.1256
R11031 GNDA.t145 GNDA.t135 16.1256
R11032 GNDA.n7237 GNDA.n7236 16.0005
R11033 GNDA.n7237 GNDA.n86 16.0005
R11034 GNDA.n6521 GNDA.n6520 16.0005
R11035 GNDA.n6524 GNDA.n6521 16.0005
R11036 GNDA.n6525 GNDA.n6524 16.0005
R11037 GNDA.n6528 GNDA.n6525 16.0005
R11038 GNDA.n6529 GNDA.n6528 16.0005
R11039 GNDA.n6532 GNDA.n6529 16.0005
R11040 GNDA.n6533 GNDA.n6532 16.0005
R11041 GNDA.n6533 GNDA.n6323 16.0005
R11042 GNDA.n6517 GNDA.n6516 16.0005
R11043 GNDA.n6516 GNDA.n6513 16.0005
R11044 GNDA.n6513 GNDA.n6512 16.0005
R11045 GNDA.n6512 GNDA.n6509 16.0005
R11046 GNDA.n6509 GNDA.n6508 16.0005
R11047 GNDA.n6508 GNDA.n6505 16.0005
R11048 GNDA.n6505 GNDA.n6504 16.0005
R11049 GNDA.n6504 GNDA.n6501 16.0005
R11050 GNDA.n6500 GNDA.n6497 16.0005
R11051 GNDA.n6497 GNDA.n6496 16.0005
R11052 GNDA.n6496 GNDA.n6493 16.0005
R11053 GNDA.n6493 GNDA.n6492 16.0005
R11054 GNDA.n6492 GNDA.n6489 16.0005
R11055 GNDA.n6489 GNDA.n6488 16.0005
R11056 GNDA.n6488 GNDA.n6485 16.0005
R11057 GNDA.n6485 GNDA.n6484 16.0005
R11058 GNDA.n6426 GNDA.n6425 16.0005
R11059 GNDA.n6429 GNDA.n6426 16.0005
R11060 GNDA.n6430 GNDA.n6429 16.0005
R11061 GNDA.n6433 GNDA.n6430 16.0005
R11062 GNDA.n6434 GNDA.n6433 16.0005
R11063 GNDA.n6437 GNDA.n6434 16.0005
R11064 GNDA.n6438 GNDA.n6437 16.0005
R11065 GNDA.n6438 GNDA.n6344 16.0005
R11066 GNDA.n6422 GNDA.n6421 16.0005
R11067 GNDA.n6421 GNDA.n6418 16.0005
R11068 GNDA.n6418 GNDA.n6417 16.0005
R11069 GNDA.n6417 GNDA.n6414 16.0005
R11070 GNDA.n6414 GNDA.n6413 16.0005
R11071 GNDA.n6413 GNDA.n6410 16.0005
R11072 GNDA.n6410 GNDA.n6409 16.0005
R11073 GNDA.n6409 GNDA.n6406 16.0005
R11074 GNDA.n6405 GNDA.n6402 16.0005
R11075 GNDA.n6402 GNDA.n6401 16.0005
R11076 GNDA.n6401 GNDA.n6398 16.0005
R11077 GNDA.n6398 GNDA.n6397 16.0005
R11078 GNDA.n6397 GNDA.n6394 16.0005
R11079 GNDA.n6394 GNDA.n6393 16.0005
R11080 GNDA.n6393 GNDA.n6390 16.0005
R11081 GNDA.n6390 GNDA.n57 16.0005
R11082 GNDA.n6888 GNDA.n6887 16.0005
R11083 GNDA.n6891 GNDA.n6888 16.0005
R11084 GNDA.n6892 GNDA.n6891 16.0005
R11085 GNDA.n6895 GNDA.n6892 16.0005
R11086 GNDA.n6896 GNDA.n6895 16.0005
R11087 GNDA.n6899 GNDA.n6896 16.0005
R11088 GNDA.n6901 GNDA.n6899 16.0005
R11089 GNDA.n6902 GNDA.n6901 16.0005
R11090 GNDA.n6884 GNDA.n6883 16.0005
R11091 GNDA.n6883 GNDA.n6880 16.0005
R11092 GNDA.n6880 GNDA.n6879 16.0005
R11093 GNDA.n6879 GNDA.n6876 16.0005
R11094 GNDA.n6876 GNDA.n6875 16.0005
R11095 GNDA.n6875 GNDA.n6872 16.0005
R11096 GNDA.n6872 GNDA.n6871 16.0005
R11097 GNDA.n6871 GNDA.n6868 16.0005
R11098 GNDA.n6867 GNDA.n6864 16.0005
R11099 GNDA.n6864 GNDA.n6863 16.0005
R11100 GNDA.n6863 GNDA.n6860 16.0005
R11101 GNDA.n6860 GNDA.n6859 16.0005
R11102 GNDA.n6859 GNDA.n6856 16.0005
R11103 GNDA.n6856 GNDA.n6855 16.0005
R11104 GNDA.n6855 GNDA.n6852 16.0005
R11105 GNDA.n6852 GNDA.n6851 16.0005
R11106 GNDA.n6625 GNDA.n6624 16.0005
R11107 GNDA.n6626 GNDA.n6625 16.0005
R11108 GNDA.n6626 GNDA.n6579 16.0005
R11109 GNDA.n6632 GNDA.n6579 16.0005
R11110 GNDA.n6633 GNDA.n6632 16.0005
R11111 GNDA.n6634 GNDA.n6633 16.0005
R11112 GNDA.n6634 GNDA.n6577 16.0005
R11113 GNDA.n6577 GNDA.n6575 16.0005
R11114 GNDA.n6618 GNDA.n6581 16.0005
R11115 GNDA.n6618 GNDA.n6617 16.0005
R11116 GNDA.n6617 GNDA.n6616 16.0005
R11117 GNDA.n6616 GNDA.n6583 16.0005
R11118 GNDA.n6610 GNDA.n6583 16.0005
R11119 GNDA.n6610 GNDA.n6609 16.0005
R11120 GNDA.n6609 GNDA.n6608 16.0005
R11121 GNDA.n6608 GNDA.n6585 16.0005
R11122 GNDA.n6602 GNDA.n6601 16.0005
R11123 GNDA.n6601 GNDA.n6600 16.0005
R11124 GNDA.n6600 GNDA.n6587 16.0005
R11125 GNDA.n6595 GNDA.n6587 16.0005
R11126 GNDA.n6595 GNDA.n6594 16.0005
R11127 GNDA.n6594 GNDA.n6593 16.0005
R11128 GNDA.n6593 GNDA.n5396 16.0005
R11129 GNDA.n6835 GNDA.n5396 16.0005
R11130 GNDA.n5701 GNDA.n5700 16.0005
R11131 GNDA.n5704 GNDA.n5701 16.0005
R11132 GNDA.n5705 GNDA.n5704 16.0005
R11133 GNDA.n5708 GNDA.n5705 16.0005
R11134 GNDA.n5709 GNDA.n5708 16.0005
R11135 GNDA.n5712 GNDA.n5709 16.0005
R11136 GNDA.n5714 GNDA.n5712 16.0005
R11137 GNDA.n5715 GNDA.n5714 16.0005
R11138 GNDA.n5697 GNDA.n5696 16.0005
R11139 GNDA.n5696 GNDA.n5693 16.0005
R11140 GNDA.n5693 GNDA.n5692 16.0005
R11141 GNDA.n5692 GNDA.n5689 16.0005
R11142 GNDA.n5689 GNDA.n5688 16.0005
R11143 GNDA.n5688 GNDA.n5685 16.0005
R11144 GNDA.n5685 GNDA.n5684 16.0005
R11145 GNDA.n5684 GNDA.n5681 16.0005
R11146 GNDA.n5680 GNDA.n5677 16.0005
R11147 GNDA.n5677 GNDA.n5676 16.0005
R11148 GNDA.n5676 GNDA.n5673 16.0005
R11149 GNDA.n5673 GNDA.n5672 16.0005
R11150 GNDA.n5672 GNDA.n5669 16.0005
R11151 GNDA.n5669 GNDA.n5668 16.0005
R11152 GNDA.n5668 GNDA.n5665 16.0005
R11153 GNDA.n5665 GNDA.n5641 16.0005
R11154 GNDA.n6043 GNDA.n6042 16.0005
R11155 GNDA.n6046 GNDA.n6043 16.0005
R11156 GNDA.n6047 GNDA.n6046 16.0005
R11157 GNDA.n6050 GNDA.n6047 16.0005
R11158 GNDA.n6051 GNDA.n6050 16.0005
R11159 GNDA.n6054 GNDA.n6051 16.0005
R11160 GNDA.n6055 GNDA.n6054 16.0005
R11161 GNDA.n6055 GNDA.n5451 16.0005
R11162 GNDA.n6039 GNDA.n6038 16.0005
R11163 GNDA.n6038 GNDA.n6035 16.0005
R11164 GNDA.n6035 GNDA.n6034 16.0005
R11165 GNDA.n6034 GNDA.n6031 16.0005
R11166 GNDA.n6031 GNDA.n6030 16.0005
R11167 GNDA.n6030 GNDA.n6027 16.0005
R11168 GNDA.n6027 GNDA.n6026 16.0005
R11169 GNDA.n6026 GNDA.n6023 16.0005
R11170 GNDA.n6022 GNDA.n6019 16.0005
R11171 GNDA.n6019 GNDA.n6018 16.0005
R11172 GNDA.n6018 GNDA.n6015 16.0005
R11173 GNDA.n6015 GNDA.n6014 16.0005
R11174 GNDA.n6014 GNDA.n6011 16.0005
R11175 GNDA.n6011 GNDA.n6010 16.0005
R11176 GNDA.n6010 GNDA.n6007 16.0005
R11177 GNDA.n6007 GNDA.n6006 16.0005
R11178 GNDA.n5980 GNDA.n5967 16.0005
R11179 GNDA.n5980 GNDA.n5979 16.0005
R11180 GNDA.n5979 GNDA.n5978 16.0005
R11181 GNDA.n5978 GNDA.n5975 16.0005
R11182 GNDA.n5975 GNDA.n5974 16.0005
R11183 GNDA.n5974 GNDA.n5971 16.0005
R11184 GNDA.n5971 GNDA.n5970 16.0005
R11185 GNDA.n5970 GNDA.n5883 16.0005
R11186 GNDA.n5966 GNDA.n5964 16.0005
R11187 GNDA.n5964 GNDA.n5961 16.0005
R11188 GNDA.n5961 GNDA.n5960 16.0005
R11189 GNDA.n5960 GNDA.n5957 16.0005
R11190 GNDA.n5957 GNDA.n5956 16.0005
R11191 GNDA.n5956 GNDA.n5953 16.0005
R11192 GNDA.n5953 GNDA.n5952 16.0005
R11193 GNDA.n5952 GNDA.n5949 16.0005
R11194 GNDA.n5948 GNDA.n5945 16.0005
R11195 GNDA.n5945 GNDA.n5944 16.0005
R11196 GNDA.n5944 GNDA.n5941 16.0005
R11197 GNDA.n5941 GNDA.n5940 16.0005
R11198 GNDA.n5940 GNDA.n5937 16.0005
R11199 GNDA.n5937 GNDA.n5936 16.0005
R11200 GNDA.n5936 GNDA.n5933 16.0005
R11201 GNDA.n5933 GNDA.n5932 16.0005
R11202 GNDA.n6723 GNDA.n6722 16.0005
R11203 GNDA.n6724 GNDA.n6723 16.0005
R11204 GNDA.n6724 GNDA.n6673 16.0005
R11205 GNDA.n6730 GNDA.n6673 16.0005
R11206 GNDA.n6731 GNDA.n6730 16.0005
R11207 GNDA.n6732 GNDA.n6731 16.0005
R11208 GNDA.n6732 GNDA.n6671 16.0005
R11209 GNDA.n6738 GNDA.n6671 16.0005
R11210 GNDA.n6716 GNDA.n6675 16.0005
R11211 GNDA.n6716 GNDA.n6715 16.0005
R11212 GNDA.n6715 GNDA.n6714 16.0005
R11213 GNDA.n6714 GNDA.n6677 16.0005
R11214 GNDA.n6708 GNDA.n6677 16.0005
R11215 GNDA.n6708 GNDA.n6707 16.0005
R11216 GNDA.n6707 GNDA.n6706 16.0005
R11217 GNDA.n6706 GNDA.n6679 16.0005
R11218 GNDA.n6700 GNDA.n6699 16.0005
R11219 GNDA.n6699 GNDA.n6698 16.0005
R11220 GNDA.n6698 GNDA.n6681 16.0005
R11221 GNDA.n6693 GNDA.n6681 16.0005
R11222 GNDA.n6693 GNDA.n6692 16.0005
R11223 GNDA.n6692 GNDA.n6691 16.0005
R11224 GNDA.n6691 GNDA.n6686 16.0005
R11225 GNDA.n6686 GNDA.n6685 16.0005
R11226 GNDA.n7333 GNDA.n7332 16.0005
R11227 GNDA.n7332 GNDA.n7329 16.0005
R11228 GNDA.n7329 GNDA.n7328 16.0005
R11229 GNDA.n7328 GNDA.n7325 16.0005
R11230 GNDA.n7325 GNDA.n7324 16.0005
R11231 GNDA.n7324 GNDA.n7321 16.0005
R11232 GNDA.n7321 GNDA.n7320 16.0005
R11233 GNDA.n7320 GNDA.n7318 16.0005
R11234 GNDA.n7337 GNDA.n7336 16.0005
R11235 GNDA.n7340 GNDA.n7337 16.0005
R11236 GNDA.n7341 GNDA.n7340 16.0005
R11237 GNDA.n7344 GNDA.n7341 16.0005
R11238 GNDA.n7345 GNDA.n7344 16.0005
R11239 GNDA.n7348 GNDA.n7345 16.0005
R11240 GNDA.n7349 GNDA.n7348 16.0005
R11241 GNDA.n7352 GNDA.n7349 16.0005
R11242 GNDA.n7356 GNDA.n7353 16.0005
R11243 GNDA.n7357 GNDA.n7356 16.0005
R11244 GNDA.n7360 GNDA.n7357 16.0005
R11245 GNDA.n7361 GNDA.n7360 16.0005
R11246 GNDA.n7364 GNDA.n7361 16.0005
R11247 GNDA.n7365 GNDA.n7364 16.0005
R11248 GNDA.n7368 GNDA.n7365 16.0005
R11249 GNDA.n7369 GNDA.n7368 16.0005
R11250 GNDA.n7309 GNDA.t145 15.9929
R11251 GNDA.n5771 GNDA.t145 15.9929
R11252 GNDA.t145 GNDA.n298 15.9929
R11253 GNDA.t109 GNDA.t264 15.8405
R11254 GNDA.t268 GNDA.t115 15.8405
R11255 GNDA.n3393 GNDA.t311 15.8405
R11256 GNDA.t7 GNDA.t96 15.8405
R11257 GNDA.t17 GNDA.t99 15.8405
R11258 GNDA.n7236 GNDA.n7235 15.1755
R11259 GNDA.n7482 GNDA.n26 14.555
R11260 GNDA.n5999 GNDA.n5446 14.555
R11261 GNDA.n5409 GNDA.t145 14.2654
R11262 GNDA.n7001 GNDA.t0 13.109
R11263 GNDA.n6995 GNDA.t0 13.109
R11264 GNDA.n6826 GNDA.t251 12.9006
R11265 GNDA.n6982 GNDA.t58 12.9006
R11266 GNDA.n6747 GNDA.t260 12.9006
R11267 GNDA.n6937 GNDA.n5360 12.8005
R11268 GNDA.n6941 GNDA.n5360 12.8005
R11269 GNDA.n6953 GNDA.n6952 12.8005
R11270 GNDA.n6952 GNDA.n5352 12.8005
R11271 GNDA.n2107 GNDA.t203 12.6791
R11272 GNDA.n5000 GNDA.t215 12.6791
R11273 GNDA.n5003 GNDA.t230 12.6791
R11274 GNDA.n658 GNDA.t191 12.6791
R11275 GNDA.n3678 GNDA.n3677 12.1358
R11276 GNDA.n715 GNDA.n714 12.1358
R11277 GNDA.n3681 GNDA.n3680 12.1114
R11278 GNDA.n2279 GNDA.n718 12.1114
R11279 GNDA.n5827 GNDA.n5568 11.6369
R11280 GNDA.n5827 GNDA.n5826 11.6369
R11281 GNDA.n5826 GNDA.n5825 11.6369
R11282 GNDA.n5825 GNDA.n5570 11.6369
R11283 GNDA.n5820 GNDA.n5570 11.6369
R11284 GNDA.n5820 GNDA.n5819 11.6369
R11285 GNDA.n5819 GNDA.n5818 11.6369
R11286 GNDA.n5818 GNDA.n5573 11.6369
R11287 GNDA.n5813 GNDA.n5573 11.6369
R11288 GNDA.n5813 GNDA.n5812 11.6369
R11289 GNDA.n5812 GNDA.n5811 11.6369
R11290 GNDA.n6322 GNDA.n6321 11.6369
R11291 GNDA.n6321 GNDA.n6258 11.6369
R11292 GNDA.n6315 GNDA.n6258 11.6369
R11293 GNDA.n6315 GNDA.n6314 11.6369
R11294 GNDA.n6314 GNDA.n6313 11.6369
R11295 GNDA.n6313 GNDA.n6263 11.6369
R11296 GNDA.n6307 GNDA.n6263 11.6369
R11297 GNDA.n6307 GNDA.n6306 11.6369
R11298 GNDA.n6306 GNDA.n6305 11.6369
R11299 GNDA.n6305 GNDA.n6267 11.6369
R11300 GNDA.n6299 GNDA.n6267 11.6369
R11301 GNDA.n6568 GNDA.n6567 11.6369
R11302 GNDA.n6567 GNDA.n6566 11.6369
R11303 GNDA.n6566 GNDA.n6565 11.6369
R11304 GNDA.n6565 GNDA.n6563 11.6369
R11305 GNDA.n6563 GNDA.n6560 11.6369
R11306 GNDA.n6560 GNDA.n6559 11.6369
R11307 GNDA.n6559 GNDA.n6556 11.6369
R11308 GNDA.n6556 GNDA.n6555 11.6369
R11309 GNDA.n6555 GNDA.n6552 11.6369
R11310 GNDA.n6552 GNDA.n6551 11.6369
R11311 GNDA.n6252 GNDA.n6251 11.6369
R11312 GNDA.n6251 GNDA.n6250 11.6369
R11313 GNDA.n6250 GNDA.n6248 11.6369
R11314 GNDA.n6248 GNDA.n6245 11.6369
R11315 GNDA.n6245 GNDA.n6244 11.6369
R11316 GNDA.n6244 GNDA.n6241 11.6369
R11317 GNDA.n6241 GNDA.n6240 11.6369
R11318 GNDA.n6240 GNDA.n6237 11.6369
R11319 GNDA.n6237 GNDA.n6236 11.6369
R11320 GNDA.n6236 GNDA.n5405 11.6369
R11321 GNDA.n5799 GNDA.n5619 11.6369
R11322 GNDA.n5799 GNDA.n5798 11.6369
R11323 GNDA.n5798 GNDA.n5797 11.6369
R11324 GNDA.n5797 GNDA.n5621 11.6369
R11325 GNDA.n5792 GNDA.n5621 11.6369
R11326 GNDA.n5792 GNDA.n5791 11.6369
R11327 GNDA.n5791 GNDA.n5790 11.6369
R11328 GNDA.n5790 GNDA.n5624 11.6369
R11329 GNDA.n5785 GNDA.n5624 11.6369
R11330 GNDA.n5785 GNDA.n5784 11.6369
R11331 GNDA.n5784 GNDA.n5783 11.6369
R11332 GNDA.n5632 GNDA.n5627 11.6369
R11333 GNDA.n5776 GNDA.n5632 11.6369
R11334 GNDA.n5776 GNDA.n5775 11.6369
R11335 GNDA.n5775 GNDA.n5774 11.6369
R11336 GNDA.n5774 GNDA.n5633 11.6369
R11337 GNDA.n5635 GNDA.n5633 11.6369
R11338 GNDA.n5638 GNDA.n5635 11.6369
R11339 GNDA.n5764 GNDA.n5638 11.6369
R11340 GNDA.n5764 GNDA.n5763 11.6369
R11341 GNDA.n5763 GNDA.n5762 11.6369
R11342 GNDA.n5855 GNDA.n5515 11.6369
R11343 GNDA.n5855 GNDA.n5854 11.6369
R11344 GNDA.n5854 GNDA.n5853 11.6369
R11345 GNDA.n5853 GNDA.n5518 11.6369
R11346 GNDA.n5848 GNDA.n5518 11.6369
R11347 GNDA.n5848 GNDA.n5847 11.6369
R11348 GNDA.n5847 GNDA.n5846 11.6369
R11349 GNDA.n5846 GNDA.n5521 11.6369
R11350 GNDA.n5841 GNDA.n5521 11.6369
R11351 GNDA.n5841 GNDA.n5840 11.6369
R11352 GNDA.n5840 GNDA.n5839 11.6369
R11353 GNDA.n5861 GNDA.n5860 11.6369
R11354 GNDA.n5864 GNDA.n5861 11.6369
R11355 GNDA.n5865 GNDA.n5864 11.6369
R11356 GNDA.n5868 GNDA.n5865 11.6369
R11357 GNDA.n5869 GNDA.n5868 11.6369
R11358 GNDA.n5872 GNDA.n5869 11.6369
R11359 GNDA.n5873 GNDA.n5872 11.6369
R11360 GNDA.n5876 GNDA.n5873 11.6369
R11361 GNDA.n5877 GNDA.n5876 11.6369
R11362 GNDA.n5880 GNDA.n5877 11.6369
R11363 GNDA.n6088 GNDA.n6083 11.6369
R11364 GNDA.n6093 GNDA.n6088 11.6369
R11365 GNDA.n6093 GNDA.n6092 11.6369
R11366 GNDA.n6092 GNDA.n6091 11.6369
R11367 GNDA.n6091 GNDA.n302 11.6369
R11368 GNDA.n7014 GNDA.n302 11.6369
R11369 GNDA.n7014 GNDA.n7013 11.6369
R11370 GNDA.n7013 GNDA.n7012 11.6369
R11371 GNDA.n7012 GNDA.n303 11.6369
R11372 GNDA.n7006 GNDA.n303 11.6369
R11373 GNDA.n6116 GNDA.n6075 11.6369
R11374 GNDA.n6116 GNDA.n6115 11.6369
R11375 GNDA.n6115 GNDA.n6114 11.6369
R11376 GNDA.n6114 GNDA.n6077 11.6369
R11377 GNDA.n6109 GNDA.n6077 11.6369
R11378 GNDA.n6109 GNDA.n6108 11.6369
R11379 GNDA.n6108 GNDA.n6107 11.6369
R11380 GNDA.n6107 GNDA.n6080 11.6369
R11381 GNDA.n6102 GNDA.n6080 11.6369
R11382 GNDA.n6102 GNDA.n6101 11.6369
R11383 GNDA.n6101 GNDA.n6100 11.6369
R11384 GNDA.n6171 GNDA.n5434 11.6369
R11385 GNDA.n6171 GNDA.n6170 11.6369
R11386 GNDA.n6170 GNDA.n6169 11.6369
R11387 GNDA.n6169 GNDA.n5438 11.6369
R11388 GNDA.n6163 GNDA.n5438 11.6369
R11389 GNDA.n6163 GNDA.n6162 11.6369
R11390 GNDA.n6162 GNDA.n6161 11.6369
R11391 GNDA.n6161 GNDA.n5440 11.6369
R11392 GNDA.n6155 GNDA.n5440 11.6369
R11393 GNDA.n6155 GNDA.n6154 11.6369
R11394 GNDA.n6154 GNDA.n6153 11.6369
R11395 GNDA.n6234 GNDA.n6233 11.6369
R11396 GNDA.n6233 GNDA.n5428 11.6369
R11397 GNDA.n6227 GNDA.n5428 11.6369
R11398 GNDA.n6227 GNDA.n6226 11.6369
R11399 GNDA.n6226 GNDA.n6225 11.6369
R11400 GNDA.n6225 GNDA.n5430 11.6369
R11401 GNDA.n6219 GNDA.n5430 11.6369
R11402 GNDA.n6219 GNDA.n6218 11.6369
R11403 GNDA.n6218 GNDA.n6217 11.6369
R11404 GNDA.n6217 GNDA.n5432 11.6369
R11405 GNDA.n6211 GNDA.n5432 11.6369
R11406 GNDA.n7410 GNDA.n7409 11.6369
R11407 GNDA.n7409 GNDA.n7408 11.6369
R11408 GNDA.n7408 GNDA.n7307 11.6369
R11409 GNDA.n7402 GNDA.n7307 11.6369
R11410 GNDA.n7402 GNDA.n7401 11.6369
R11411 GNDA.n7401 GNDA.n7400 11.6369
R11412 GNDA.n7400 GNDA.n7311 11.6369
R11413 GNDA.n7394 GNDA.n7311 11.6369
R11414 GNDA.n7394 GNDA.n7393 11.6369
R11415 GNDA.n7393 GNDA.n7392 11.6369
R11416 GNDA.n7434 GNDA.n7433 11.6369
R11417 GNDA.n7433 GNDA.n7432 11.6369
R11418 GNDA.n7432 GNDA.n7295 11.6369
R11419 GNDA.n7426 GNDA.n7295 11.6369
R11420 GNDA.n7426 GNDA.n7425 11.6369
R11421 GNDA.n7425 GNDA.n7424 11.6369
R11422 GNDA.n7424 GNDA.n7299 11.6369
R11423 GNDA.n7418 GNDA.n7299 11.6369
R11424 GNDA.n7418 GNDA.n7417 11.6369
R11425 GNDA.n7417 GNDA.n7416 11.6369
R11426 GNDA.n7416 GNDA.n7303 11.6369
R11427 GNDA.n7460 GNDA.n7459 11.6369
R11428 GNDA.n7459 GNDA.n7458 11.6369
R11429 GNDA.n7458 GNDA.n82 11.6369
R11430 GNDA.n7452 GNDA.n82 11.6369
R11431 GNDA.n7452 GNDA.n7451 11.6369
R11432 GNDA.n7449 GNDA.n87 11.6369
R11433 GNDA.n7443 GNDA.n87 11.6369
R11434 GNDA.n7443 GNDA.n7442 11.6369
R11435 GNDA.n7442 GNDA.n7441 11.6369
R11436 GNDA.n7441 GNDA.n7242 11.6369
R11437 GNDA.n3398 GNDA.n3397 11.4533
R11438 GNDA.n5308 GNDA.n318 11.4533
R11439 GNDA.t149 GNDA.t19 11.37
R11440 GNDA.n1756 GNDA.n1755 11.2033
R11441 GNDA.n1744 GNDA.n1743 11.2033
R11442 GNDA.n7035 GNDA.n7034 10.9846
R11443 GNDA.n7051 GNDA.n269 10.87
R11444 GNDA.n7048 GNDA.n272 10.87
R11445 GNDA.n7047 GNDA.n273 10.87
R11446 GNDA.n7043 GNDA.n277 10.87
R11447 GNDA.n7042 GNDA.n278 10.87
R11448 GNDA.n7039 GNDA.n281 10.87
R11449 GNDA.n7038 GNDA.n282 10.87
R11450 GNDA.t217 GNDA.t21 10.5605
R11451 GNDA.t101 GNDA.t123 10.5605
R11452 GNDA.t295 GNDA.t54 10.5605
R11453 GNDA.t56 GNDA.t75 10.5605
R11454 GNDA.t254 GNDA.t211 10.5605
R11455 GNDA.n1773 GNDA.t12 9.6005
R11456 GNDA.n1773 GNDA.t300 9.6005
R11457 GNDA.n5283 GNDA.t267 9.6005
R11458 GNDA.n5283 GNDA.t173 9.6005
R11459 GNDA.n5285 GNDA.t312 9.6005
R11460 GNDA.n5285 GNDA.t132 9.6005
R11461 GNDA.n5287 GNDA.t338 9.6005
R11462 GNDA.n5287 GNDA.t134 9.6005
R11463 GNDA.n5289 GNDA.t139 9.6005
R11464 GNDA.n5289 GNDA.t292 9.6005
R11465 GNDA.n5291 GNDA.t302 9.6005
R11466 GNDA.n5291 GNDA.t38 9.6005
R11467 GNDA.n5293 GNDA.t253 9.6005
R11468 GNDA.n5293 GNDA.t296 9.6005
R11469 GNDA.n5295 GNDA.t270 9.6005
R11470 GNDA.n5295 GNDA.t79 9.6005
R11471 GNDA.n5297 GNDA.t61 9.6005
R11472 GNDA.n5297 GNDA.t41 9.6005
R11473 GNDA.n5299 GNDA.t305 9.6005
R11474 GNDA.n5299 GNDA.t72 9.6005
R11475 GNDA.n5301 GNDA.t298 9.6005
R11476 GNDA.n5301 GNDA.t272 9.6005
R11477 GNDA.n5303 GNDA.t50 9.6005
R11478 GNDA.n5303 GNDA.t66 9.6005
R11479 GNDA.n6768 GNDA.t284 9.6005
R11480 GNDA.n6664 GNDA.t275 9.6005
R11481 GNDA.n6782 GNDA.t280 9.6005
R11482 GNDA.n6791 GNDA.t282 9.6005
R11483 GNDA.n6937 GNDA.n5358 9.36264
R11484 GNDA.n6953 GNDA.n5351 9.36264
R11485 GNDA.n5360 GNDA.n5359 9.3005
R11486 GNDA.n6942 GNDA.n6941 9.3005
R11487 GNDA.n6952 GNDA.n6951 9.3005
R11488 GNDA.n6950 GNDA.n5352 9.3005
R11489 GNDA.t108 GNDA.t288 8.8005
R11490 GNDA.t62 GNDA.t114 8.8005
R11491 GNDA.t256 GNDA.n5307 8.8005
R11492 GNDA.t40 GNDA.n1732 8.8005
R11493 GNDA.t290 GNDA.n3394 8.8005
R11494 GNDA.t47 GNDA.t316 8.8005
R11495 GNDA.t320 GNDA.t127 8.8005
R11496 GNDA.n7473 GNDA.n26 8.60107
R11497 GNDA.n6070 GNDA.n5446 8.60107
R11498 GNDA.t195 GNDA.n6824 8.60055
R11499 GNDA.t334 GNDA.n5401 8.60055
R11500 GNDA.t286 GNDA.n6959 8.60055
R11501 GNDA.n6748 GNDA.t293 8.60055
R11502 GNDA.n6998 GNDA.n93 8.50251
R11503 GNDA.n5408 GNDA.t16 7.95916
R11504 GNDA.n6260 GNDA.t145 7.65068
R11505 GNDA.n7398 GNDA.t145 7.60343
R11506 GNDA.n5768 GNDA.t145 7.60343
R11507 GNDA.t145 GNDA.n7016 7.60343
R11508 GNDA.n6813 GNDA.t45 7.52554
R11509 GNDA.n6825 GNDA.t137 7.52554
R11510 GNDA.n6843 GNDA.n5363 7.52554
R11511 GNDA.n7032 GNDA.n286 7.52554
R11512 GNDA.n1732 GNDA.t90 7.0405
R11513 GNDA.t184 GNDA.t301 7.0405
R11514 GNDA.t21 GNDA.t37 7.0405
R11515 GNDA.t123 GNDA.t138 7.0405
R11516 GNDA.t54 GNDA.t291 7.0405
R11517 GNDA.t75 GNDA.t337 7.0405
R11518 GNDA.t211 GNDA.t133 7.0405
R11519 GNDA.t306 GNDA.n6987 7.03568
R11520 GNDA.n5811 GNDA.n61 6.72373
R11521 GNDA.n6299 GNDA.n81 6.72373
R11522 GNDA.n5839 GNDA.n5524 6.72373
R11523 GNDA.n6153 GNDA.n6073 6.72373
R11524 GNDA.n6211 GNDA.n6210 6.72373
R11525 GNDA.n7294 GNDA.n7242 6.72373
R11526 GNDA.t97 GNDA.t145 6.45054
R11527 GNDA.n5568 GNDA.n5524 6.20656
R11528 GNDA.n5619 GNDA.n61 6.20656
R11529 GNDA.n6075 GNDA.n6073 6.20656
R11530 GNDA.n6210 GNDA.n5434 6.20656
R11531 GNDA.n7434 GNDA.n7294 6.20656
R11532 GNDA.n7460 GNDA.n81 6.20656
R11533 GNDA.n7451 GNDA.n7450 6.07727
R11534 GNDA.n6792 GNDA.n6783 5.81868
R11535 GNDA.n6790 GNDA.n6783 5.81868
R11536 GNDA.n7450 GNDA.n7449 5.5601
R11537 GNDA.n6484 GNDA.n6454 5.51161
R11538 GNDA.n7478 GNDA.n57 5.51161
R11539 GNDA.n6851 GNDA.n5368 5.51161
R11540 GNDA.n6907 GNDA.n6835 5.51161
R11541 GNDA.n5753 GNDA.n5641 5.51161
R11542 GNDA.n6006 GNDA.n5473 5.51161
R11543 GNDA.n5932 GNDA.n5910 5.51161
R11544 GNDA.n6685 GNDA.n6684 5.51161
R11545 GNDA.n7383 GNDA.n7369 5.51161
R11546 GNDA.t125 GNDA.t247 5.37553
R11547 GNDA.n6794 GNDA.t52 5.37553
R11548 GNDA.t145 GNDA.t155 5.37553
R11549 GNDA.n6983 GNDA.t145 5.37553
R11550 GNDA.t145 GNDA.t179 5.37553
R11551 GNDA.n6774 GNDA.t135 5.37553
R11552 GNDA.t26 GNDA.t244 5.37553
R11553 GNDA.t43 GNDA.t73 5.34355
R11554 GNDA.t324 GNDA.t44 5.34355
R11555 GNDA.n5754 GNDA.n5639 5.1717
R11556 GNDA.n7005 GNDA.n307 5.1717
R11557 GNDA.n7384 GNDA.n7315 5.1717
R11558 GNDA.t86 GNDA.t310 5.10195
R11559 GNDA.t84 GNDA.t102 5.10195
R11560 GNDA.n5305 GNDA.n5304 5.063
R11561 GNDA.n6548 GNDA.n6545 4.9157
R11562 GNDA.n6822 GNDA.n6574 4.9157
R11563 GNDA.n5996 GNDA.n5882 4.9157
R11564 GNDA.n5284 GNDA.n5282 4.71925
R11565 GNDA.n3423 GNDA.n3422 4.5005
R11566 GNDA.n3429 GNDA.n3405 4.5005
R11567 GNDA.n3430 GNDA.n589 4.5005
R11568 GNDA.n3430 GNDA.n3429 4.5005
R11569 GNDA.n1713 GNDA.n1712 4.5005
R11570 GNDA.n1716 GNDA.n1715 4.5005
R11571 GNDA.n1771 GNDA.n1708 4.5005
R11572 GNDA.n1770 GNDA.n1769 4.5005
R11573 GNDA.n1771 GNDA.n1770 4.5005
R11574 GNDA.n1779 GNDA.n1778 4.5005
R11575 GNDA.n1724 GNDA.n1702 4.5005
R11576 GNDA.n1721 GNDA.n1702 4.5005
R11577 GNDA.n1722 GNDA.n1721 4.5005
R11578 GNDA.n1786 GNDA.n1699 4.5005
R11579 GNDA.n1785 GNDA.n1784 4.5005
R11580 GNDA.n1786 GNDA.n1785 4.5005
R11581 GNDA.n1802 GNDA.n1801 4.5005
R11582 GNDA.n1808 GNDA.n1807 4.5005
R11583 GNDA.n5275 GNDA.n5274 4.5005
R11584 GNDA.n327 GNDA.n326 4.5005
R11585 GNDA.n5160 GNDA.n5159 4.5005
R11586 GNDA.n5164 GNDA.n5161 4.5005
R11587 GNDA.n5165 GNDA.n5158 4.5005
R11588 GNDA.n5169 GNDA.n5168 4.5005
R11589 GNDA.n5170 GNDA.n5157 4.5005
R11590 GNDA.n5174 GNDA.n5171 4.5005
R11591 GNDA.n5175 GNDA.n5156 4.5005
R11592 GNDA.n5179 GNDA.n5178 4.5005
R11593 GNDA.n5180 GNDA.n5155 4.5005
R11594 GNDA.n5184 GNDA.n5181 4.5005
R11595 GNDA.n5185 GNDA.n5154 4.5005
R11596 GNDA.n5189 GNDA.n5188 4.5005
R11597 GNDA.n5190 GNDA.n5153 4.5005
R11598 GNDA.n5194 GNDA.n5191 4.5005
R11599 GNDA.n5195 GNDA.n5152 4.5005
R11600 GNDA.n5199 GNDA.n5198 4.5005
R11601 GNDA.n5200 GNDA.n5151 4.5005
R11602 GNDA.n5204 GNDA.n5201 4.5005
R11603 GNDA.n5205 GNDA.n5150 4.5005
R11604 GNDA.n5209 GNDA.n5208 4.5005
R11605 GNDA.n5210 GNDA.n5149 4.5005
R11606 GNDA.n5214 GNDA.n5211 4.5005
R11607 GNDA.n5215 GNDA.n5148 4.5005
R11608 GNDA.n5219 GNDA.n5218 4.5005
R11609 GNDA.n5220 GNDA.n5147 4.5005
R11610 GNDA.n5224 GNDA.n5221 4.5005
R11611 GNDA.n5225 GNDA.n5146 4.5005
R11612 GNDA.n5229 GNDA.n5228 4.5005
R11613 GNDA.n5230 GNDA.n5145 4.5005
R11614 GNDA.n5234 GNDA.n5231 4.5005
R11615 GNDA.n5235 GNDA.n5144 4.5005
R11616 GNDA.n5239 GNDA.n5238 4.5005
R11617 GNDA.n5240 GNDA.n5143 4.5005
R11618 GNDA.n5244 GNDA.n5241 4.5005
R11619 GNDA.n5245 GNDA.n5142 4.5005
R11620 GNDA.n5249 GNDA.n5248 4.5005
R11621 GNDA.n5250 GNDA.n5141 4.5005
R11622 GNDA.n5254 GNDA.n5251 4.5005
R11623 GNDA.n5255 GNDA.n5140 4.5005
R11624 GNDA.n5259 GNDA.n5258 4.5005
R11625 GNDA.n5260 GNDA.n5139 4.5005
R11626 GNDA.n5264 GNDA.n5261 4.5005
R11627 GNDA.n5265 GNDA.n5138 4.5005
R11628 GNDA.n5269 GNDA.n5268 4.5005
R11629 GNDA.n4962 GNDA.n4961 4.5005
R11630 GNDA.n3457 GNDA.n3456 4.5005
R11631 GNDA.n4847 GNDA.n4846 4.5005
R11632 GNDA.n4851 GNDA.n4848 4.5005
R11633 GNDA.n4852 GNDA.n4845 4.5005
R11634 GNDA.n4856 GNDA.n4855 4.5005
R11635 GNDA.n4857 GNDA.n4844 4.5005
R11636 GNDA.n4861 GNDA.n4858 4.5005
R11637 GNDA.n4862 GNDA.n4843 4.5005
R11638 GNDA.n4866 GNDA.n4865 4.5005
R11639 GNDA.n4867 GNDA.n4842 4.5005
R11640 GNDA.n4871 GNDA.n4868 4.5005
R11641 GNDA.n4872 GNDA.n4841 4.5005
R11642 GNDA.n4876 GNDA.n4875 4.5005
R11643 GNDA.n4877 GNDA.n4840 4.5005
R11644 GNDA.n4881 GNDA.n4878 4.5005
R11645 GNDA.n4882 GNDA.n4839 4.5005
R11646 GNDA.n4886 GNDA.n4885 4.5005
R11647 GNDA.n4887 GNDA.n4838 4.5005
R11648 GNDA.n4891 GNDA.n4888 4.5005
R11649 GNDA.n4892 GNDA.n4837 4.5005
R11650 GNDA.n4896 GNDA.n4895 4.5005
R11651 GNDA.n4897 GNDA.n4836 4.5005
R11652 GNDA.n4901 GNDA.n4898 4.5005
R11653 GNDA.n4902 GNDA.n4835 4.5005
R11654 GNDA.n4906 GNDA.n4905 4.5005
R11655 GNDA.n4907 GNDA.n4834 4.5005
R11656 GNDA.n4911 GNDA.n4908 4.5005
R11657 GNDA.n4912 GNDA.n4833 4.5005
R11658 GNDA.n4916 GNDA.n4915 4.5005
R11659 GNDA.n4917 GNDA.n4832 4.5005
R11660 GNDA.n4921 GNDA.n4918 4.5005
R11661 GNDA.n4922 GNDA.n4831 4.5005
R11662 GNDA.n4926 GNDA.n4925 4.5005
R11663 GNDA.n4927 GNDA.n4830 4.5005
R11664 GNDA.n4931 GNDA.n4928 4.5005
R11665 GNDA.n4932 GNDA.n4829 4.5005
R11666 GNDA.n4936 GNDA.n4935 4.5005
R11667 GNDA.n4937 GNDA.n4828 4.5005
R11668 GNDA.n4941 GNDA.n4938 4.5005
R11669 GNDA.n4942 GNDA.n4827 4.5005
R11670 GNDA.n4946 GNDA.n4945 4.5005
R11671 GNDA.n4947 GNDA.n4826 4.5005
R11672 GNDA.n4951 GNDA.n4948 4.5005
R11673 GNDA.n4952 GNDA.n4825 4.5005
R11674 GNDA.n4956 GNDA.n4955 4.5005
R11675 GNDA.n4683 GNDA.n4682 4.5005
R11676 GNDA.n4686 GNDA.n4685 4.5005
R11677 GNDA.n4687 GNDA.n4681 4.5005
R11678 GNDA.n4691 GNDA.n4688 4.5005
R11679 GNDA.n4692 GNDA.n4680 4.5005
R11680 GNDA.n4696 GNDA.n4695 4.5005
R11681 GNDA.n4697 GNDA.n4679 4.5005
R11682 GNDA.n4701 GNDA.n4698 4.5005
R11683 GNDA.n4702 GNDA.n4678 4.5005
R11684 GNDA.n4706 GNDA.n4705 4.5005
R11685 GNDA.n4707 GNDA.n4677 4.5005
R11686 GNDA.n4711 GNDA.n4708 4.5005
R11687 GNDA.n4712 GNDA.n4676 4.5005
R11688 GNDA.n4716 GNDA.n4715 4.5005
R11689 GNDA.n4717 GNDA.n4675 4.5005
R11690 GNDA.n4721 GNDA.n4718 4.5005
R11691 GNDA.n4722 GNDA.n4674 4.5005
R11692 GNDA.n4726 GNDA.n4725 4.5005
R11693 GNDA.n4727 GNDA.n4673 4.5005
R11694 GNDA.n4731 GNDA.n4728 4.5005
R11695 GNDA.n4732 GNDA.n4672 4.5005
R11696 GNDA.n4736 GNDA.n4735 4.5005
R11697 GNDA.n4737 GNDA.n4671 4.5005
R11698 GNDA.n4741 GNDA.n4738 4.5005
R11699 GNDA.n4742 GNDA.n4670 4.5005
R11700 GNDA.n4746 GNDA.n4745 4.5005
R11701 GNDA.n4747 GNDA.n4669 4.5005
R11702 GNDA.n4751 GNDA.n4748 4.5005
R11703 GNDA.n4752 GNDA.n4668 4.5005
R11704 GNDA.n4756 GNDA.n4755 4.5005
R11705 GNDA.n4757 GNDA.n4667 4.5005
R11706 GNDA.n4761 GNDA.n4758 4.5005
R11707 GNDA.n4762 GNDA.n4666 4.5005
R11708 GNDA.n4766 GNDA.n4765 4.5005
R11709 GNDA.n4767 GNDA.n4665 4.5005
R11710 GNDA.n4771 GNDA.n4768 4.5005
R11711 GNDA.n4772 GNDA.n4664 4.5005
R11712 GNDA.n4776 GNDA.n4775 4.5005
R11713 GNDA.n4777 GNDA.n4663 4.5005
R11714 GNDA.n4781 GNDA.n4778 4.5005
R11715 GNDA.n4782 GNDA.n4662 4.5005
R11716 GNDA.n4786 GNDA.n4785 4.5005
R11717 GNDA.n4787 GNDA.n4661 4.5005
R11718 GNDA.n4791 GNDA.n4788 4.5005
R11719 GNDA.n4792 GNDA.n4660 4.5005
R11720 GNDA.n4796 GNDA.n4795 4.5005
R11721 GNDA.n4517 GNDA.n4516 4.5005
R11722 GNDA.n4520 GNDA.n4519 4.5005
R11723 GNDA.n4521 GNDA.n4515 4.5005
R11724 GNDA.n4525 GNDA.n4522 4.5005
R11725 GNDA.n4526 GNDA.n4514 4.5005
R11726 GNDA.n4530 GNDA.n4529 4.5005
R11727 GNDA.n4531 GNDA.n4513 4.5005
R11728 GNDA.n4535 GNDA.n4532 4.5005
R11729 GNDA.n4536 GNDA.n4512 4.5005
R11730 GNDA.n4540 GNDA.n4539 4.5005
R11731 GNDA.n4541 GNDA.n4511 4.5005
R11732 GNDA.n4545 GNDA.n4542 4.5005
R11733 GNDA.n4546 GNDA.n4510 4.5005
R11734 GNDA.n4550 GNDA.n4549 4.5005
R11735 GNDA.n4551 GNDA.n4509 4.5005
R11736 GNDA.n4555 GNDA.n4552 4.5005
R11737 GNDA.n4556 GNDA.n4508 4.5005
R11738 GNDA.n4560 GNDA.n4559 4.5005
R11739 GNDA.n4561 GNDA.n4507 4.5005
R11740 GNDA.n4565 GNDA.n4562 4.5005
R11741 GNDA.n4566 GNDA.n4506 4.5005
R11742 GNDA.n4570 GNDA.n4569 4.5005
R11743 GNDA.n4571 GNDA.n4505 4.5005
R11744 GNDA.n4575 GNDA.n4572 4.5005
R11745 GNDA.n4576 GNDA.n4504 4.5005
R11746 GNDA.n4580 GNDA.n4579 4.5005
R11747 GNDA.n4581 GNDA.n4503 4.5005
R11748 GNDA.n4585 GNDA.n4582 4.5005
R11749 GNDA.n4586 GNDA.n4502 4.5005
R11750 GNDA.n4590 GNDA.n4589 4.5005
R11751 GNDA.n4591 GNDA.n4501 4.5005
R11752 GNDA.n4595 GNDA.n4592 4.5005
R11753 GNDA.n4596 GNDA.n4500 4.5005
R11754 GNDA.n4600 GNDA.n4599 4.5005
R11755 GNDA.n4601 GNDA.n4499 4.5005
R11756 GNDA.n4605 GNDA.n4602 4.5005
R11757 GNDA.n4606 GNDA.n4498 4.5005
R11758 GNDA.n4610 GNDA.n4609 4.5005
R11759 GNDA.n4611 GNDA.n4497 4.5005
R11760 GNDA.n4615 GNDA.n4612 4.5005
R11761 GNDA.n4616 GNDA.n4496 4.5005
R11762 GNDA.n4620 GNDA.n4619 4.5005
R11763 GNDA.n4621 GNDA.n4495 4.5005
R11764 GNDA.n4625 GNDA.n4622 4.5005
R11765 GNDA.n4626 GNDA.n4494 4.5005
R11766 GNDA.n4630 GNDA.n4629 4.5005
R11767 GNDA.n4351 GNDA.n4350 4.5005
R11768 GNDA.n4354 GNDA.n4353 4.5005
R11769 GNDA.n4355 GNDA.n4349 4.5005
R11770 GNDA.n4359 GNDA.n4356 4.5005
R11771 GNDA.n4360 GNDA.n4348 4.5005
R11772 GNDA.n4364 GNDA.n4363 4.5005
R11773 GNDA.n4365 GNDA.n4347 4.5005
R11774 GNDA.n4369 GNDA.n4366 4.5005
R11775 GNDA.n4370 GNDA.n4346 4.5005
R11776 GNDA.n4374 GNDA.n4373 4.5005
R11777 GNDA.n4375 GNDA.n4345 4.5005
R11778 GNDA.n4379 GNDA.n4376 4.5005
R11779 GNDA.n4380 GNDA.n4344 4.5005
R11780 GNDA.n4384 GNDA.n4383 4.5005
R11781 GNDA.n4385 GNDA.n4343 4.5005
R11782 GNDA.n4389 GNDA.n4386 4.5005
R11783 GNDA.n4390 GNDA.n4342 4.5005
R11784 GNDA.n4394 GNDA.n4393 4.5005
R11785 GNDA.n4395 GNDA.n4341 4.5005
R11786 GNDA.n4399 GNDA.n4396 4.5005
R11787 GNDA.n4400 GNDA.n4340 4.5005
R11788 GNDA.n4404 GNDA.n4403 4.5005
R11789 GNDA.n4405 GNDA.n4339 4.5005
R11790 GNDA.n4409 GNDA.n4406 4.5005
R11791 GNDA.n4410 GNDA.n4338 4.5005
R11792 GNDA.n4414 GNDA.n4413 4.5005
R11793 GNDA.n4415 GNDA.n4337 4.5005
R11794 GNDA.n4419 GNDA.n4416 4.5005
R11795 GNDA.n4420 GNDA.n4336 4.5005
R11796 GNDA.n4424 GNDA.n4423 4.5005
R11797 GNDA.n4425 GNDA.n4335 4.5005
R11798 GNDA.n4429 GNDA.n4426 4.5005
R11799 GNDA.n4430 GNDA.n4334 4.5005
R11800 GNDA.n4434 GNDA.n4433 4.5005
R11801 GNDA.n4435 GNDA.n4333 4.5005
R11802 GNDA.n4439 GNDA.n4436 4.5005
R11803 GNDA.n4440 GNDA.n4332 4.5005
R11804 GNDA.n4444 GNDA.n4443 4.5005
R11805 GNDA.n4445 GNDA.n4331 4.5005
R11806 GNDA.n4449 GNDA.n4446 4.5005
R11807 GNDA.n4450 GNDA.n4330 4.5005
R11808 GNDA.n4454 GNDA.n4453 4.5005
R11809 GNDA.n4455 GNDA.n4329 4.5005
R11810 GNDA.n4459 GNDA.n4456 4.5005
R11811 GNDA.n4460 GNDA.n4328 4.5005
R11812 GNDA.n4464 GNDA.n4463 4.5005
R11813 GNDA.n4185 GNDA.n4184 4.5005
R11814 GNDA.n4188 GNDA.n4187 4.5005
R11815 GNDA.n4189 GNDA.n4183 4.5005
R11816 GNDA.n4193 GNDA.n4190 4.5005
R11817 GNDA.n4194 GNDA.n4182 4.5005
R11818 GNDA.n4198 GNDA.n4197 4.5005
R11819 GNDA.n4199 GNDA.n4181 4.5005
R11820 GNDA.n4203 GNDA.n4200 4.5005
R11821 GNDA.n4204 GNDA.n4180 4.5005
R11822 GNDA.n4208 GNDA.n4207 4.5005
R11823 GNDA.n4209 GNDA.n4179 4.5005
R11824 GNDA.n4213 GNDA.n4210 4.5005
R11825 GNDA.n4214 GNDA.n4178 4.5005
R11826 GNDA.n4218 GNDA.n4217 4.5005
R11827 GNDA.n4219 GNDA.n4177 4.5005
R11828 GNDA.n4223 GNDA.n4220 4.5005
R11829 GNDA.n4224 GNDA.n4176 4.5005
R11830 GNDA.n4228 GNDA.n4227 4.5005
R11831 GNDA.n4229 GNDA.n4175 4.5005
R11832 GNDA.n4233 GNDA.n4230 4.5005
R11833 GNDA.n4234 GNDA.n4174 4.5005
R11834 GNDA.n4238 GNDA.n4237 4.5005
R11835 GNDA.n4239 GNDA.n4173 4.5005
R11836 GNDA.n4243 GNDA.n4240 4.5005
R11837 GNDA.n4244 GNDA.n4172 4.5005
R11838 GNDA.n4248 GNDA.n4247 4.5005
R11839 GNDA.n4249 GNDA.n4171 4.5005
R11840 GNDA.n4253 GNDA.n4250 4.5005
R11841 GNDA.n4254 GNDA.n4170 4.5005
R11842 GNDA.n4258 GNDA.n4257 4.5005
R11843 GNDA.n4259 GNDA.n4169 4.5005
R11844 GNDA.n4263 GNDA.n4260 4.5005
R11845 GNDA.n4264 GNDA.n4168 4.5005
R11846 GNDA.n4268 GNDA.n4267 4.5005
R11847 GNDA.n4269 GNDA.n4167 4.5005
R11848 GNDA.n4273 GNDA.n4270 4.5005
R11849 GNDA.n4274 GNDA.n4166 4.5005
R11850 GNDA.n4278 GNDA.n4277 4.5005
R11851 GNDA.n4279 GNDA.n4165 4.5005
R11852 GNDA.n4283 GNDA.n4280 4.5005
R11853 GNDA.n4284 GNDA.n4164 4.5005
R11854 GNDA.n4288 GNDA.n4287 4.5005
R11855 GNDA.n4289 GNDA.n4163 4.5005
R11856 GNDA.n4293 GNDA.n4290 4.5005
R11857 GNDA.n4294 GNDA.n4162 4.5005
R11858 GNDA.n4298 GNDA.n4297 4.5005
R11859 GNDA.n3687 GNDA.n3686 4.5005
R11860 GNDA.n3690 GNDA.n3689 4.5005
R11861 GNDA.n3691 GNDA.n3507 4.5005
R11862 GNDA.n3695 GNDA.n3692 4.5005
R11863 GNDA.n3696 GNDA.n3506 4.5005
R11864 GNDA.n3700 GNDA.n3699 4.5005
R11865 GNDA.n3701 GNDA.n3505 4.5005
R11866 GNDA.n3705 GNDA.n3702 4.5005
R11867 GNDA.n3706 GNDA.n3504 4.5005
R11868 GNDA.n3710 GNDA.n3709 4.5005
R11869 GNDA.n3711 GNDA.n3503 4.5005
R11870 GNDA.n3715 GNDA.n3712 4.5005
R11871 GNDA.n3716 GNDA.n3502 4.5005
R11872 GNDA.n3720 GNDA.n3719 4.5005
R11873 GNDA.n3721 GNDA.n3501 4.5005
R11874 GNDA.n3725 GNDA.n3722 4.5005
R11875 GNDA.n3726 GNDA.n3500 4.5005
R11876 GNDA.n3730 GNDA.n3729 4.5005
R11877 GNDA.n3731 GNDA.n3499 4.5005
R11878 GNDA.n3735 GNDA.n3732 4.5005
R11879 GNDA.n3736 GNDA.n3498 4.5005
R11880 GNDA.n3740 GNDA.n3739 4.5005
R11881 GNDA.n3741 GNDA.n3497 4.5005
R11882 GNDA.n3745 GNDA.n3742 4.5005
R11883 GNDA.n3746 GNDA.n3496 4.5005
R11884 GNDA.n3750 GNDA.n3749 4.5005
R11885 GNDA.n3751 GNDA.n3495 4.5005
R11886 GNDA.n3755 GNDA.n3752 4.5005
R11887 GNDA.n3756 GNDA.n3494 4.5005
R11888 GNDA.n3760 GNDA.n3759 4.5005
R11889 GNDA.n3761 GNDA.n3493 4.5005
R11890 GNDA.n3765 GNDA.n3762 4.5005
R11891 GNDA.n3766 GNDA.n3492 4.5005
R11892 GNDA.n3770 GNDA.n3769 4.5005
R11893 GNDA.n3771 GNDA.n3491 4.5005
R11894 GNDA.n3775 GNDA.n3772 4.5005
R11895 GNDA.n3776 GNDA.n3490 4.5005
R11896 GNDA.n3780 GNDA.n3779 4.5005
R11897 GNDA.n3781 GNDA.n3489 4.5005
R11898 GNDA.n3785 GNDA.n3782 4.5005
R11899 GNDA.n3786 GNDA.n3488 4.5005
R11900 GNDA.n3790 GNDA.n3789 4.5005
R11901 GNDA.n3791 GNDA.n3487 4.5005
R11902 GNDA.n3795 GNDA.n3792 4.5005
R11903 GNDA.n3796 GNDA.n3486 4.5005
R11904 GNDA.n3800 GNDA.n3799 4.5005
R11905 GNDA.n4019 GNDA.n4018 4.5005
R11906 GNDA.n4022 GNDA.n4021 4.5005
R11907 GNDA.n4023 GNDA.n4017 4.5005
R11908 GNDA.n4027 GNDA.n4024 4.5005
R11909 GNDA.n4028 GNDA.n4016 4.5005
R11910 GNDA.n4032 GNDA.n4031 4.5005
R11911 GNDA.n4033 GNDA.n4015 4.5005
R11912 GNDA.n4037 GNDA.n4034 4.5005
R11913 GNDA.n4038 GNDA.n4014 4.5005
R11914 GNDA.n4042 GNDA.n4041 4.5005
R11915 GNDA.n4043 GNDA.n4013 4.5005
R11916 GNDA.n4047 GNDA.n4044 4.5005
R11917 GNDA.n4048 GNDA.n4012 4.5005
R11918 GNDA.n4052 GNDA.n4051 4.5005
R11919 GNDA.n4053 GNDA.n4011 4.5005
R11920 GNDA.n4057 GNDA.n4054 4.5005
R11921 GNDA.n4058 GNDA.n4010 4.5005
R11922 GNDA.n4062 GNDA.n4061 4.5005
R11923 GNDA.n4063 GNDA.n4009 4.5005
R11924 GNDA.n4067 GNDA.n4064 4.5005
R11925 GNDA.n4068 GNDA.n4008 4.5005
R11926 GNDA.n4072 GNDA.n4071 4.5005
R11927 GNDA.n4073 GNDA.n4007 4.5005
R11928 GNDA.n4077 GNDA.n4074 4.5005
R11929 GNDA.n4078 GNDA.n4006 4.5005
R11930 GNDA.n4082 GNDA.n4081 4.5005
R11931 GNDA.n4083 GNDA.n4005 4.5005
R11932 GNDA.n4087 GNDA.n4084 4.5005
R11933 GNDA.n4088 GNDA.n4004 4.5005
R11934 GNDA.n4092 GNDA.n4091 4.5005
R11935 GNDA.n4093 GNDA.n4003 4.5005
R11936 GNDA.n4097 GNDA.n4094 4.5005
R11937 GNDA.n4098 GNDA.n4002 4.5005
R11938 GNDA.n4102 GNDA.n4101 4.5005
R11939 GNDA.n4103 GNDA.n4001 4.5005
R11940 GNDA.n4107 GNDA.n4104 4.5005
R11941 GNDA.n4108 GNDA.n4000 4.5005
R11942 GNDA.n4112 GNDA.n4111 4.5005
R11943 GNDA.n4113 GNDA.n3999 4.5005
R11944 GNDA.n4117 GNDA.n4114 4.5005
R11945 GNDA.n4118 GNDA.n3998 4.5005
R11946 GNDA.n4122 GNDA.n4121 4.5005
R11947 GNDA.n4123 GNDA.n3997 4.5005
R11948 GNDA.n4127 GNDA.n4124 4.5005
R11949 GNDA.n4128 GNDA.n3996 4.5005
R11950 GNDA.n4132 GNDA.n4131 4.5005
R11951 GNDA.n3853 GNDA.n3852 4.5005
R11952 GNDA.n3856 GNDA.n3855 4.5005
R11953 GNDA.n3857 GNDA.n3851 4.5005
R11954 GNDA.n3861 GNDA.n3858 4.5005
R11955 GNDA.n3862 GNDA.n3850 4.5005
R11956 GNDA.n3866 GNDA.n3865 4.5005
R11957 GNDA.n3867 GNDA.n3849 4.5005
R11958 GNDA.n3871 GNDA.n3868 4.5005
R11959 GNDA.n3872 GNDA.n3848 4.5005
R11960 GNDA.n3876 GNDA.n3875 4.5005
R11961 GNDA.n3877 GNDA.n3847 4.5005
R11962 GNDA.n3881 GNDA.n3878 4.5005
R11963 GNDA.n3882 GNDA.n3846 4.5005
R11964 GNDA.n3886 GNDA.n3885 4.5005
R11965 GNDA.n3887 GNDA.n3845 4.5005
R11966 GNDA.n3891 GNDA.n3888 4.5005
R11967 GNDA.n3892 GNDA.n3844 4.5005
R11968 GNDA.n3896 GNDA.n3895 4.5005
R11969 GNDA.n3897 GNDA.n3843 4.5005
R11970 GNDA.n3901 GNDA.n3898 4.5005
R11971 GNDA.n3902 GNDA.n3842 4.5005
R11972 GNDA.n3906 GNDA.n3905 4.5005
R11973 GNDA.n3907 GNDA.n3841 4.5005
R11974 GNDA.n3911 GNDA.n3908 4.5005
R11975 GNDA.n3912 GNDA.n3840 4.5005
R11976 GNDA.n3916 GNDA.n3915 4.5005
R11977 GNDA.n3917 GNDA.n3839 4.5005
R11978 GNDA.n3921 GNDA.n3918 4.5005
R11979 GNDA.n3922 GNDA.n3838 4.5005
R11980 GNDA.n3926 GNDA.n3925 4.5005
R11981 GNDA.n3927 GNDA.n3837 4.5005
R11982 GNDA.n3931 GNDA.n3928 4.5005
R11983 GNDA.n3932 GNDA.n3836 4.5005
R11984 GNDA.n3936 GNDA.n3935 4.5005
R11985 GNDA.n3937 GNDA.n3835 4.5005
R11986 GNDA.n3941 GNDA.n3938 4.5005
R11987 GNDA.n3942 GNDA.n3834 4.5005
R11988 GNDA.n3946 GNDA.n3945 4.5005
R11989 GNDA.n3947 GNDA.n3833 4.5005
R11990 GNDA.n3951 GNDA.n3948 4.5005
R11991 GNDA.n3952 GNDA.n3832 4.5005
R11992 GNDA.n3956 GNDA.n3955 4.5005
R11993 GNDA.n3957 GNDA.n3831 4.5005
R11994 GNDA.n3961 GNDA.n3958 4.5005
R11995 GNDA.n3962 GNDA.n3830 4.5005
R11996 GNDA.n3966 GNDA.n3965 4.5005
R11997 GNDA.n3675 GNDA.n3674 4.5005
R11998 GNDA.n3512 GNDA.n3511 4.5005
R11999 GNDA.n3558 GNDA.n3513 4.5005
R12000 GNDA.n3559 GNDA.n3514 4.5005
R12001 GNDA.n3560 GNDA.n3515 4.5005
R12002 GNDA.n3561 GNDA.n3516 4.5005
R12003 GNDA.n3562 GNDA.n3517 4.5005
R12004 GNDA.n3563 GNDA.n3518 4.5005
R12005 GNDA.n3564 GNDA.n3519 4.5005
R12006 GNDA.n3565 GNDA.n3520 4.5005
R12007 GNDA.n3566 GNDA.n3521 4.5005
R12008 GNDA.n3567 GNDA.n3522 4.5005
R12009 GNDA.n3568 GNDA.n3523 4.5005
R12010 GNDA.n3569 GNDA.n3524 4.5005
R12011 GNDA.n3570 GNDA.n3525 4.5005
R12012 GNDA.n3571 GNDA.n3526 4.5005
R12013 GNDA.n3572 GNDA.n3527 4.5005
R12014 GNDA.n3573 GNDA.n3528 4.5005
R12015 GNDA.n3574 GNDA.n3529 4.5005
R12016 GNDA.n3575 GNDA.n3530 4.5005
R12017 GNDA.n3576 GNDA.n3531 4.5005
R12018 GNDA.n3577 GNDA.n3532 4.5005
R12019 GNDA.n3578 GNDA.n3533 4.5005
R12020 GNDA.n3579 GNDA.n3534 4.5005
R12021 GNDA.n3580 GNDA.n3535 4.5005
R12022 GNDA.n3581 GNDA.n3536 4.5005
R12023 GNDA.n3582 GNDA.n3537 4.5005
R12024 GNDA.n3583 GNDA.n3538 4.5005
R12025 GNDA.n3584 GNDA.n3539 4.5005
R12026 GNDA.n3585 GNDA.n3540 4.5005
R12027 GNDA.n3586 GNDA.n3541 4.5005
R12028 GNDA.n3587 GNDA.n3542 4.5005
R12029 GNDA.n3588 GNDA.n3543 4.5005
R12030 GNDA.n3589 GNDA.n3544 4.5005
R12031 GNDA.n3590 GNDA.n3545 4.5005
R12032 GNDA.n3591 GNDA.n3546 4.5005
R12033 GNDA.n3592 GNDA.n3547 4.5005
R12034 GNDA.n3593 GNDA.n3548 4.5005
R12035 GNDA.n3594 GNDA.n3549 4.5005
R12036 GNDA.n3595 GNDA.n3550 4.5005
R12037 GNDA.n3596 GNDA.n3551 4.5005
R12038 GNDA.n3597 GNDA.n3552 4.5005
R12039 GNDA.n3598 GNDA.n3553 4.5005
R12040 GNDA.n3599 GNDA.n3554 4.5005
R12041 GNDA.n3600 GNDA.n3555 4.5005
R12042 GNDA.n3601 GNDA.n3556 4.5005
R12043 GNDA.n569 GNDA.n568 4.5005
R12044 GNDA.n406 GNDA.n405 4.5005
R12045 GNDA.n452 GNDA.n407 4.5005
R12046 GNDA.n453 GNDA.n408 4.5005
R12047 GNDA.n454 GNDA.n409 4.5005
R12048 GNDA.n455 GNDA.n410 4.5005
R12049 GNDA.n456 GNDA.n411 4.5005
R12050 GNDA.n457 GNDA.n412 4.5005
R12051 GNDA.n458 GNDA.n413 4.5005
R12052 GNDA.n459 GNDA.n414 4.5005
R12053 GNDA.n460 GNDA.n415 4.5005
R12054 GNDA.n461 GNDA.n416 4.5005
R12055 GNDA.n462 GNDA.n417 4.5005
R12056 GNDA.n463 GNDA.n418 4.5005
R12057 GNDA.n464 GNDA.n419 4.5005
R12058 GNDA.n465 GNDA.n420 4.5005
R12059 GNDA.n466 GNDA.n421 4.5005
R12060 GNDA.n467 GNDA.n422 4.5005
R12061 GNDA.n468 GNDA.n423 4.5005
R12062 GNDA.n469 GNDA.n424 4.5005
R12063 GNDA.n470 GNDA.n425 4.5005
R12064 GNDA.n471 GNDA.n426 4.5005
R12065 GNDA.n472 GNDA.n427 4.5005
R12066 GNDA.n473 GNDA.n428 4.5005
R12067 GNDA.n474 GNDA.n429 4.5005
R12068 GNDA.n475 GNDA.n430 4.5005
R12069 GNDA.n476 GNDA.n431 4.5005
R12070 GNDA.n477 GNDA.n432 4.5005
R12071 GNDA.n478 GNDA.n433 4.5005
R12072 GNDA.n479 GNDA.n434 4.5005
R12073 GNDA.n480 GNDA.n435 4.5005
R12074 GNDA.n481 GNDA.n436 4.5005
R12075 GNDA.n482 GNDA.n437 4.5005
R12076 GNDA.n483 GNDA.n438 4.5005
R12077 GNDA.n484 GNDA.n439 4.5005
R12078 GNDA.n485 GNDA.n440 4.5005
R12079 GNDA.n486 GNDA.n441 4.5005
R12080 GNDA.n487 GNDA.n442 4.5005
R12081 GNDA.n488 GNDA.n443 4.5005
R12082 GNDA.n489 GNDA.n444 4.5005
R12083 GNDA.n490 GNDA.n445 4.5005
R12084 GNDA.n491 GNDA.n446 4.5005
R12085 GNDA.n492 GNDA.n447 4.5005
R12086 GNDA.n493 GNDA.n448 4.5005
R12087 GNDA.n494 GNDA.n449 4.5005
R12088 GNDA.n495 GNDA.n450 4.5005
R12089 GNDA.n5019 GNDA.n5018 4.5005
R12090 GNDA.n5022 GNDA.n5021 4.5005
R12091 GNDA.n5023 GNDA.n401 4.5005
R12092 GNDA.n5027 GNDA.n5024 4.5005
R12093 GNDA.n5028 GNDA.n400 4.5005
R12094 GNDA.n5032 GNDA.n5031 4.5005
R12095 GNDA.n5033 GNDA.n399 4.5005
R12096 GNDA.n5037 GNDA.n5034 4.5005
R12097 GNDA.n5038 GNDA.n398 4.5005
R12098 GNDA.n5042 GNDA.n5041 4.5005
R12099 GNDA.n5043 GNDA.n397 4.5005
R12100 GNDA.n5047 GNDA.n5044 4.5005
R12101 GNDA.n5048 GNDA.n396 4.5005
R12102 GNDA.n5052 GNDA.n5051 4.5005
R12103 GNDA.n5053 GNDA.n395 4.5005
R12104 GNDA.n5057 GNDA.n5054 4.5005
R12105 GNDA.n5058 GNDA.n394 4.5005
R12106 GNDA.n5062 GNDA.n5061 4.5005
R12107 GNDA.n5063 GNDA.n393 4.5005
R12108 GNDA.n5067 GNDA.n5064 4.5005
R12109 GNDA.n5068 GNDA.n392 4.5005
R12110 GNDA.n5072 GNDA.n5071 4.5005
R12111 GNDA.n5073 GNDA.n391 4.5005
R12112 GNDA.n5077 GNDA.n5074 4.5005
R12113 GNDA.n5078 GNDA.n390 4.5005
R12114 GNDA.n5082 GNDA.n5081 4.5005
R12115 GNDA.n5083 GNDA.n389 4.5005
R12116 GNDA.n5087 GNDA.n5084 4.5005
R12117 GNDA.n5088 GNDA.n388 4.5005
R12118 GNDA.n5092 GNDA.n5091 4.5005
R12119 GNDA.n5093 GNDA.n387 4.5005
R12120 GNDA.n5097 GNDA.n5094 4.5005
R12121 GNDA.n5098 GNDA.n386 4.5005
R12122 GNDA.n5102 GNDA.n5101 4.5005
R12123 GNDA.n5103 GNDA.n385 4.5005
R12124 GNDA.n5107 GNDA.n5104 4.5005
R12125 GNDA.n5108 GNDA.n384 4.5005
R12126 GNDA.n5112 GNDA.n5111 4.5005
R12127 GNDA.n5113 GNDA.n383 4.5005
R12128 GNDA.n5117 GNDA.n5114 4.5005
R12129 GNDA.n5118 GNDA.n382 4.5005
R12130 GNDA.n5122 GNDA.n5121 4.5005
R12131 GNDA.n5123 GNDA.n381 4.5005
R12132 GNDA.n5127 GNDA.n5124 4.5005
R12133 GNDA.n5128 GNDA.n380 4.5005
R12134 GNDA.n5132 GNDA.n5131 4.5005
R12135 GNDA.n3372 GNDA.n3371 4.5005
R12136 GNDA.n3209 GNDA.n3208 4.5005
R12137 GNDA.n3255 GNDA.n3210 4.5005
R12138 GNDA.n3256 GNDA.n3211 4.5005
R12139 GNDA.n3257 GNDA.n3212 4.5005
R12140 GNDA.n3258 GNDA.n3213 4.5005
R12141 GNDA.n3259 GNDA.n3214 4.5005
R12142 GNDA.n3260 GNDA.n3215 4.5005
R12143 GNDA.n3261 GNDA.n3216 4.5005
R12144 GNDA.n3262 GNDA.n3217 4.5005
R12145 GNDA.n3263 GNDA.n3218 4.5005
R12146 GNDA.n3264 GNDA.n3219 4.5005
R12147 GNDA.n3265 GNDA.n3220 4.5005
R12148 GNDA.n3266 GNDA.n3221 4.5005
R12149 GNDA.n3267 GNDA.n3222 4.5005
R12150 GNDA.n3268 GNDA.n3223 4.5005
R12151 GNDA.n3269 GNDA.n3224 4.5005
R12152 GNDA.n3270 GNDA.n3225 4.5005
R12153 GNDA.n3271 GNDA.n3226 4.5005
R12154 GNDA.n3272 GNDA.n3227 4.5005
R12155 GNDA.n3273 GNDA.n3228 4.5005
R12156 GNDA.n3274 GNDA.n3229 4.5005
R12157 GNDA.n3275 GNDA.n3230 4.5005
R12158 GNDA.n3276 GNDA.n3231 4.5005
R12159 GNDA.n3277 GNDA.n3232 4.5005
R12160 GNDA.n3278 GNDA.n3233 4.5005
R12161 GNDA.n3279 GNDA.n3234 4.5005
R12162 GNDA.n3280 GNDA.n3235 4.5005
R12163 GNDA.n3281 GNDA.n3236 4.5005
R12164 GNDA.n3282 GNDA.n3237 4.5005
R12165 GNDA.n3283 GNDA.n3238 4.5005
R12166 GNDA.n3284 GNDA.n3239 4.5005
R12167 GNDA.n3285 GNDA.n3240 4.5005
R12168 GNDA.n3286 GNDA.n3241 4.5005
R12169 GNDA.n3287 GNDA.n3242 4.5005
R12170 GNDA.n3288 GNDA.n3243 4.5005
R12171 GNDA.n3289 GNDA.n3244 4.5005
R12172 GNDA.n3290 GNDA.n3245 4.5005
R12173 GNDA.n3291 GNDA.n3246 4.5005
R12174 GNDA.n3292 GNDA.n3247 4.5005
R12175 GNDA.n3293 GNDA.n3248 4.5005
R12176 GNDA.n3294 GNDA.n3249 4.5005
R12177 GNDA.n3295 GNDA.n3250 4.5005
R12178 GNDA.n3296 GNDA.n3251 4.5005
R12179 GNDA.n3297 GNDA.n3252 4.5005
R12180 GNDA.n3298 GNDA.n3253 4.5005
R12181 GNDA.n3200 GNDA.n3199 4.5005
R12182 GNDA.n597 GNDA.n596 4.5005
R12183 GNDA.n3085 GNDA.n3084 4.5005
R12184 GNDA.n3089 GNDA.n3086 4.5005
R12185 GNDA.n3090 GNDA.n3083 4.5005
R12186 GNDA.n3094 GNDA.n3093 4.5005
R12187 GNDA.n3095 GNDA.n3082 4.5005
R12188 GNDA.n3099 GNDA.n3096 4.5005
R12189 GNDA.n3100 GNDA.n3081 4.5005
R12190 GNDA.n3104 GNDA.n3103 4.5005
R12191 GNDA.n3105 GNDA.n3080 4.5005
R12192 GNDA.n3109 GNDA.n3106 4.5005
R12193 GNDA.n3110 GNDA.n3079 4.5005
R12194 GNDA.n3114 GNDA.n3113 4.5005
R12195 GNDA.n3115 GNDA.n3078 4.5005
R12196 GNDA.n3119 GNDA.n3116 4.5005
R12197 GNDA.n3120 GNDA.n3077 4.5005
R12198 GNDA.n3124 GNDA.n3123 4.5005
R12199 GNDA.n3125 GNDA.n3076 4.5005
R12200 GNDA.n3129 GNDA.n3126 4.5005
R12201 GNDA.n3130 GNDA.n3075 4.5005
R12202 GNDA.n3134 GNDA.n3133 4.5005
R12203 GNDA.n3135 GNDA.n3074 4.5005
R12204 GNDA.n3139 GNDA.n3136 4.5005
R12205 GNDA.n3140 GNDA.n3073 4.5005
R12206 GNDA.n3144 GNDA.n3143 4.5005
R12207 GNDA.n3145 GNDA.n3072 4.5005
R12208 GNDA.n3149 GNDA.n3146 4.5005
R12209 GNDA.n3150 GNDA.n3071 4.5005
R12210 GNDA.n3154 GNDA.n3153 4.5005
R12211 GNDA.n3155 GNDA.n3070 4.5005
R12212 GNDA.n3159 GNDA.n3156 4.5005
R12213 GNDA.n3160 GNDA.n3069 4.5005
R12214 GNDA.n3164 GNDA.n3163 4.5005
R12215 GNDA.n3165 GNDA.n3068 4.5005
R12216 GNDA.n3169 GNDA.n3166 4.5005
R12217 GNDA.n3170 GNDA.n3067 4.5005
R12218 GNDA.n3174 GNDA.n3173 4.5005
R12219 GNDA.n3175 GNDA.n3066 4.5005
R12220 GNDA.n3179 GNDA.n3176 4.5005
R12221 GNDA.n3180 GNDA.n3065 4.5005
R12222 GNDA.n3184 GNDA.n3183 4.5005
R12223 GNDA.n3185 GNDA.n3064 4.5005
R12224 GNDA.n3189 GNDA.n3186 4.5005
R12225 GNDA.n3190 GNDA.n3063 4.5005
R12226 GNDA.n3194 GNDA.n3193 4.5005
R12227 GNDA.n2921 GNDA.n2920 4.5005
R12228 GNDA.n2924 GNDA.n2923 4.5005
R12229 GNDA.n2925 GNDA.n2911 4.5005
R12230 GNDA.n2929 GNDA.n2926 4.5005
R12231 GNDA.n2930 GNDA.n2910 4.5005
R12232 GNDA.n2934 GNDA.n2933 4.5005
R12233 GNDA.n2935 GNDA.n2909 4.5005
R12234 GNDA.n2939 GNDA.n2936 4.5005
R12235 GNDA.n2940 GNDA.n2908 4.5005
R12236 GNDA.n2944 GNDA.n2943 4.5005
R12237 GNDA.n2945 GNDA.n2907 4.5005
R12238 GNDA.n2949 GNDA.n2946 4.5005
R12239 GNDA.n2950 GNDA.n2906 4.5005
R12240 GNDA.n2954 GNDA.n2953 4.5005
R12241 GNDA.n2955 GNDA.n2905 4.5005
R12242 GNDA.n2959 GNDA.n2956 4.5005
R12243 GNDA.n2960 GNDA.n2904 4.5005
R12244 GNDA.n2964 GNDA.n2963 4.5005
R12245 GNDA.n2965 GNDA.n2903 4.5005
R12246 GNDA.n2969 GNDA.n2966 4.5005
R12247 GNDA.n2970 GNDA.n2902 4.5005
R12248 GNDA.n2974 GNDA.n2973 4.5005
R12249 GNDA.n2975 GNDA.n2901 4.5005
R12250 GNDA.n2979 GNDA.n2976 4.5005
R12251 GNDA.n2980 GNDA.n2900 4.5005
R12252 GNDA.n2984 GNDA.n2983 4.5005
R12253 GNDA.n2985 GNDA.n2899 4.5005
R12254 GNDA.n2989 GNDA.n2986 4.5005
R12255 GNDA.n2990 GNDA.n2898 4.5005
R12256 GNDA.n2994 GNDA.n2993 4.5005
R12257 GNDA.n2995 GNDA.n2897 4.5005
R12258 GNDA.n2999 GNDA.n2996 4.5005
R12259 GNDA.n3000 GNDA.n2896 4.5005
R12260 GNDA.n3004 GNDA.n3003 4.5005
R12261 GNDA.n3005 GNDA.n2895 4.5005
R12262 GNDA.n3009 GNDA.n3006 4.5005
R12263 GNDA.n3010 GNDA.n2894 4.5005
R12264 GNDA.n3014 GNDA.n3013 4.5005
R12265 GNDA.n3015 GNDA.n2893 4.5005
R12266 GNDA.n3019 GNDA.n3016 4.5005
R12267 GNDA.n3020 GNDA.n2892 4.5005
R12268 GNDA.n3024 GNDA.n3023 4.5005
R12269 GNDA.n3025 GNDA.n2891 4.5005
R12270 GNDA.n3029 GNDA.n3026 4.5005
R12271 GNDA.n3030 GNDA.n2890 4.5005
R12272 GNDA.n3034 GNDA.n3033 4.5005
R12273 GNDA.n2285 GNDA.n2284 4.5005
R12274 GNDA.n2288 GNDA.n2287 4.5005
R12275 GNDA.n2289 GNDA.n713 4.5005
R12276 GNDA.n2293 GNDA.n2290 4.5005
R12277 GNDA.n2294 GNDA.n712 4.5005
R12278 GNDA.n2298 GNDA.n2297 4.5005
R12279 GNDA.n2299 GNDA.n711 4.5005
R12280 GNDA.n2303 GNDA.n2300 4.5005
R12281 GNDA.n2304 GNDA.n710 4.5005
R12282 GNDA.n2308 GNDA.n2307 4.5005
R12283 GNDA.n2309 GNDA.n709 4.5005
R12284 GNDA.n2313 GNDA.n2310 4.5005
R12285 GNDA.n2314 GNDA.n708 4.5005
R12286 GNDA.n2318 GNDA.n2317 4.5005
R12287 GNDA.n2319 GNDA.n707 4.5005
R12288 GNDA.n2323 GNDA.n2320 4.5005
R12289 GNDA.n2324 GNDA.n706 4.5005
R12290 GNDA.n2328 GNDA.n2327 4.5005
R12291 GNDA.n2329 GNDA.n705 4.5005
R12292 GNDA.n2333 GNDA.n2330 4.5005
R12293 GNDA.n2334 GNDA.n704 4.5005
R12294 GNDA.n2338 GNDA.n2337 4.5005
R12295 GNDA.n2339 GNDA.n703 4.5005
R12296 GNDA.n2343 GNDA.n2340 4.5005
R12297 GNDA.n2344 GNDA.n702 4.5005
R12298 GNDA.n2348 GNDA.n2347 4.5005
R12299 GNDA.n2349 GNDA.n701 4.5005
R12300 GNDA.n2353 GNDA.n2350 4.5005
R12301 GNDA.n2354 GNDA.n700 4.5005
R12302 GNDA.n2358 GNDA.n2357 4.5005
R12303 GNDA.n2359 GNDA.n699 4.5005
R12304 GNDA.n2363 GNDA.n2360 4.5005
R12305 GNDA.n2364 GNDA.n698 4.5005
R12306 GNDA.n2368 GNDA.n2367 4.5005
R12307 GNDA.n2369 GNDA.n697 4.5005
R12308 GNDA.n2373 GNDA.n2370 4.5005
R12309 GNDA.n2374 GNDA.n696 4.5005
R12310 GNDA.n2378 GNDA.n2377 4.5005
R12311 GNDA.n2379 GNDA.n695 4.5005
R12312 GNDA.n2383 GNDA.n2380 4.5005
R12313 GNDA.n2384 GNDA.n694 4.5005
R12314 GNDA.n2388 GNDA.n2387 4.5005
R12315 GNDA.n2389 GNDA.n693 4.5005
R12316 GNDA.n2393 GNDA.n2390 4.5005
R12317 GNDA.n2394 GNDA.n692 4.5005
R12318 GNDA.n2398 GNDA.n2397 4.5005
R12319 GNDA.n2747 GNDA.n2746 4.5005
R12320 GNDA.n2750 GNDA.n2749 4.5005
R12321 GNDA.n2751 GNDA.n647 4.5005
R12322 GNDA.n2755 GNDA.n2752 4.5005
R12323 GNDA.n2756 GNDA.n646 4.5005
R12324 GNDA.n2760 GNDA.n2759 4.5005
R12325 GNDA.n2761 GNDA.n645 4.5005
R12326 GNDA.n2765 GNDA.n2762 4.5005
R12327 GNDA.n2766 GNDA.n644 4.5005
R12328 GNDA.n2770 GNDA.n2769 4.5005
R12329 GNDA.n2771 GNDA.n643 4.5005
R12330 GNDA.n2775 GNDA.n2772 4.5005
R12331 GNDA.n2776 GNDA.n642 4.5005
R12332 GNDA.n2780 GNDA.n2779 4.5005
R12333 GNDA.n2781 GNDA.n641 4.5005
R12334 GNDA.n2785 GNDA.n2782 4.5005
R12335 GNDA.n2786 GNDA.n640 4.5005
R12336 GNDA.n2790 GNDA.n2789 4.5005
R12337 GNDA.n2791 GNDA.n639 4.5005
R12338 GNDA.n2795 GNDA.n2792 4.5005
R12339 GNDA.n2796 GNDA.n638 4.5005
R12340 GNDA.n2800 GNDA.n2799 4.5005
R12341 GNDA.n2801 GNDA.n637 4.5005
R12342 GNDA.n2805 GNDA.n2802 4.5005
R12343 GNDA.n2806 GNDA.n636 4.5005
R12344 GNDA.n2810 GNDA.n2809 4.5005
R12345 GNDA.n2811 GNDA.n635 4.5005
R12346 GNDA.n2815 GNDA.n2812 4.5005
R12347 GNDA.n2816 GNDA.n634 4.5005
R12348 GNDA.n2820 GNDA.n2819 4.5005
R12349 GNDA.n2821 GNDA.n633 4.5005
R12350 GNDA.n2825 GNDA.n2822 4.5005
R12351 GNDA.n2826 GNDA.n632 4.5005
R12352 GNDA.n2830 GNDA.n2829 4.5005
R12353 GNDA.n2831 GNDA.n631 4.5005
R12354 GNDA.n2835 GNDA.n2832 4.5005
R12355 GNDA.n2836 GNDA.n630 4.5005
R12356 GNDA.n2840 GNDA.n2839 4.5005
R12357 GNDA.n2841 GNDA.n629 4.5005
R12358 GNDA.n2845 GNDA.n2842 4.5005
R12359 GNDA.n2846 GNDA.n628 4.5005
R12360 GNDA.n2850 GNDA.n2849 4.5005
R12361 GNDA.n2851 GNDA.n627 4.5005
R12362 GNDA.n2855 GNDA.n2852 4.5005
R12363 GNDA.n2856 GNDA.n626 4.5005
R12364 GNDA.n2860 GNDA.n2859 4.5005
R12365 GNDA.n2735 GNDA.n2734 4.5005
R12366 GNDA.n2572 GNDA.n2571 4.5005
R12367 GNDA.n2618 GNDA.n2573 4.5005
R12368 GNDA.n2619 GNDA.n2574 4.5005
R12369 GNDA.n2620 GNDA.n2575 4.5005
R12370 GNDA.n2621 GNDA.n2576 4.5005
R12371 GNDA.n2622 GNDA.n2577 4.5005
R12372 GNDA.n2623 GNDA.n2578 4.5005
R12373 GNDA.n2624 GNDA.n2579 4.5005
R12374 GNDA.n2625 GNDA.n2580 4.5005
R12375 GNDA.n2626 GNDA.n2581 4.5005
R12376 GNDA.n2627 GNDA.n2582 4.5005
R12377 GNDA.n2628 GNDA.n2583 4.5005
R12378 GNDA.n2629 GNDA.n2584 4.5005
R12379 GNDA.n2630 GNDA.n2585 4.5005
R12380 GNDA.n2631 GNDA.n2586 4.5005
R12381 GNDA.n2632 GNDA.n2587 4.5005
R12382 GNDA.n2633 GNDA.n2588 4.5005
R12383 GNDA.n2634 GNDA.n2589 4.5005
R12384 GNDA.n2635 GNDA.n2590 4.5005
R12385 GNDA.n2636 GNDA.n2591 4.5005
R12386 GNDA.n2637 GNDA.n2592 4.5005
R12387 GNDA.n2638 GNDA.n2593 4.5005
R12388 GNDA.n2639 GNDA.n2594 4.5005
R12389 GNDA.n2640 GNDA.n2595 4.5005
R12390 GNDA.n2641 GNDA.n2596 4.5005
R12391 GNDA.n2642 GNDA.n2597 4.5005
R12392 GNDA.n2643 GNDA.n2598 4.5005
R12393 GNDA.n2644 GNDA.n2599 4.5005
R12394 GNDA.n2645 GNDA.n2600 4.5005
R12395 GNDA.n2646 GNDA.n2601 4.5005
R12396 GNDA.n2647 GNDA.n2602 4.5005
R12397 GNDA.n2648 GNDA.n2603 4.5005
R12398 GNDA.n2649 GNDA.n2604 4.5005
R12399 GNDA.n2650 GNDA.n2605 4.5005
R12400 GNDA.n2651 GNDA.n2606 4.5005
R12401 GNDA.n2652 GNDA.n2607 4.5005
R12402 GNDA.n2653 GNDA.n2608 4.5005
R12403 GNDA.n2654 GNDA.n2609 4.5005
R12404 GNDA.n2655 GNDA.n2610 4.5005
R12405 GNDA.n2656 GNDA.n2611 4.5005
R12406 GNDA.n2657 GNDA.n2612 4.5005
R12407 GNDA.n2658 GNDA.n2613 4.5005
R12408 GNDA.n2659 GNDA.n2614 4.5005
R12409 GNDA.n2660 GNDA.n2615 4.5005
R12410 GNDA.n2661 GNDA.n2616 4.5005
R12411 GNDA.n2564 GNDA.n2563 4.5005
R12412 GNDA.n663 GNDA.n662 4.5005
R12413 GNDA.n2449 GNDA.n2448 4.5005
R12414 GNDA.n2453 GNDA.n2450 4.5005
R12415 GNDA.n2454 GNDA.n2447 4.5005
R12416 GNDA.n2458 GNDA.n2457 4.5005
R12417 GNDA.n2459 GNDA.n2446 4.5005
R12418 GNDA.n2463 GNDA.n2460 4.5005
R12419 GNDA.n2464 GNDA.n2445 4.5005
R12420 GNDA.n2468 GNDA.n2467 4.5005
R12421 GNDA.n2469 GNDA.n2444 4.5005
R12422 GNDA.n2473 GNDA.n2470 4.5005
R12423 GNDA.n2474 GNDA.n2443 4.5005
R12424 GNDA.n2478 GNDA.n2477 4.5005
R12425 GNDA.n2479 GNDA.n2442 4.5005
R12426 GNDA.n2483 GNDA.n2480 4.5005
R12427 GNDA.n2484 GNDA.n2441 4.5005
R12428 GNDA.n2488 GNDA.n2487 4.5005
R12429 GNDA.n2489 GNDA.n2440 4.5005
R12430 GNDA.n2493 GNDA.n2490 4.5005
R12431 GNDA.n2494 GNDA.n2439 4.5005
R12432 GNDA.n2498 GNDA.n2497 4.5005
R12433 GNDA.n2499 GNDA.n2438 4.5005
R12434 GNDA.n2503 GNDA.n2500 4.5005
R12435 GNDA.n2504 GNDA.n2437 4.5005
R12436 GNDA.n2508 GNDA.n2507 4.5005
R12437 GNDA.n2509 GNDA.n2436 4.5005
R12438 GNDA.n2513 GNDA.n2510 4.5005
R12439 GNDA.n2514 GNDA.n2435 4.5005
R12440 GNDA.n2518 GNDA.n2517 4.5005
R12441 GNDA.n2519 GNDA.n2434 4.5005
R12442 GNDA.n2523 GNDA.n2520 4.5005
R12443 GNDA.n2524 GNDA.n2433 4.5005
R12444 GNDA.n2528 GNDA.n2527 4.5005
R12445 GNDA.n2529 GNDA.n2432 4.5005
R12446 GNDA.n2533 GNDA.n2530 4.5005
R12447 GNDA.n2534 GNDA.n2431 4.5005
R12448 GNDA.n2538 GNDA.n2537 4.5005
R12449 GNDA.n2539 GNDA.n2430 4.5005
R12450 GNDA.n2543 GNDA.n2540 4.5005
R12451 GNDA.n2544 GNDA.n2429 4.5005
R12452 GNDA.n2548 GNDA.n2547 4.5005
R12453 GNDA.n2549 GNDA.n2428 4.5005
R12454 GNDA.n2553 GNDA.n2550 4.5005
R12455 GNDA.n2554 GNDA.n2427 4.5005
R12456 GNDA.n2558 GNDA.n2557 4.5005
R12457 GNDA.n2275 GNDA.n2274 4.5005
R12458 GNDA.n2112 GNDA.n2111 4.5005
R12459 GNDA.n2158 GNDA.n2113 4.5005
R12460 GNDA.n2159 GNDA.n2114 4.5005
R12461 GNDA.n2160 GNDA.n2115 4.5005
R12462 GNDA.n2161 GNDA.n2116 4.5005
R12463 GNDA.n2162 GNDA.n2117 4.5005
R12464 GNDA.n2163 GNDA.n2118 4.5005
R12465 GNDA.n2164 GNDA.n2119 4.5005
R12466 GNDA.n2165 GNDA.n2120 4.5005
R12467 GNDA.n2166 GNDA.n2121 4.5005
R12468 GNDA.n2167 GNDA.n2122 4.5005
R12469 GNDA.n2168 GNDA.n2123 4.5005
R12470 GNDA.n2169 GNDA.n2124 4.5005
R12471 GNDA.n2170 GNDA.n2125 4.5005
R12472 GNDA.n2171 GNDA.n2126 4.5005
R12473 GNDA.n2172 GNDA.n2127 4.5005
R12474 GNDA.n2173 GNDA.n2128 4.5005
R12475 GNDA.n2174 GNDA.n2129 4.5005
R12476 GNDA.n2175 GNDA.n2130 4.5005
R12477 GNDA.n2176 GNDA.n2131 4.5005
R12478 GNDA.n2177 GNDA.n2132 4.5005
R12479 GNDA.n2178 GNDA.n2133 4.5005
R12480 GNDA.n2179 GNDA.n2134 4.5005
R12481 GNDA.n2180 GNDA.n2135 4.5005
R12482 GNDA.n2181 GNDA.n2136 4.5005
R12483 GNDA.n2182 GNDA.n2137 4.5005
R12484 GNDA.n2183 GNDA.n2138 4.5005
R12485 GNDA.n2184 GNDA.n2139 4.5005
R12486 GNDA.n2185 GNDA.n2140 4.5005
R12487 GNDA.n2186 GNDA.n2141 4.5005
R12488 GNDA.n2187 GNDA.n2142 4.5005
R12489 GNDA.n2188 GNDA.n2143 4.5005
R12490 GNDA.n2189 GNDA.n2144 4.5005
R12491 GNDA.n2190 GNDA.n2145 4.5005
R12492 GNDA.n2191 GNDA.n2146 4.5005
R12493 GNDA.n2192 GNDA.n2147 4.5005
R12494 GNDA.n2193 GNDA.n2148 4.5005
R12495 GNDA.n2194 GNDA.n2149 4.5005
R12496 GNDA.n2195 GNDA.n2150 4.5005
R12497 GNDA.n2196 GNDA.n2151 4.5005
R12498 GNDA.n2197 GNDA.n2152 4.5005
R12499 GNDA.n2198 GNDA.n2153 4.5005
R12500 GNDA.n2199 GNDA.n2154 4.5005
R12501 GNDA.n2200 GNDA.n2155 4.5005
R12502 GNDA.n2201 GNDA.n2156 4.5005
R12503 GNDA.n2101 GNDA.n2100 4.5005
R12504 GNDA.n726 GNDA.n725 4.5005
R12505 GNDA.n1986 GNDA.n1985 4.5005
R12506 GNDA.n1990 GNDA.n1987 4.5005
R12507 GNDA.n1991 GNDA.n1984 4.5005
R12508 GNDA.n1995 GNDA.n1994 4.5005
R12509 GNDA.n1996 GNDA.n1983 4.5005
R12510 GNDA.n2000 GNDA.n1997 4.5005
R12511 GNDA.n2001 GNDA.n1982 4.5005
R12512 GNDA.n2005 GNDA.n2004 4.5005
R12513 GNDA.n2006 GNDA.n1981 4.5005
R12514 GNDA.n2010 GNDA.n2007 4.5005
R12515 GNDA.n2011 GNDA.n1980 4.5005
R12516 GNDA.n2015 GNDA.n2014 4.5005
R12517 GNDA.n2016 GNDA.n1979 4.5005
R12518 GNDA.n2020 GNDA.n2017 4.5005
R12519 GNDA.n2021 GNDA.n1978 4.5005
R12520 GNDA.n2025 GNDA.n2024 4.5005
R12521 GNDA.n2026 GNDA.n1977 4.5005
R12522 GNDA.n2030 GNDA.n2027 4.5005
R12523 GNDA.n2031 GNDA.n1976 4.5005
R12524 GNDA.n2035 GNDA.n2034 4.5005
R12525 GNDA.n2036 GNDA.n1975 4.5005
R12526 GNDA.n2040 GNDA.n2037 4.5005
R12527 GNDA.n2041 GNDA.n1974 4.5005
R12528 GNDA.n2045 GNDA.n2044 4.5005
R12529 GNDA.n2046 GNDA.n1973 4.5005
R12530 GNDA.n2050 GNDA.n2047 4.5005
R12531 GNDA.n2051 GNDA.n1972 4.5005
R12532 GNDA.n2055 GNDA.n2054 4.5005
R12533 GNDA.n2056 GNDA.n1971 4.5005
R12534 GNDA.n2060 GNDA.n2057 4.5005
R12535 GNDA.n2061 GNDA.n1970 4.5005
R12536 GNDA.n2065 GNDA.n2064 4.5005
R12537 GNDA.n2066 GNDA.n1969 4.5005
R12538 GNDA.n2070 GNDA.n2067 4.5005
R12539 GNDA.n2071 GNDA.n1968 4.5005
R12540 GNDA.n2075 GNDA.n2074 4.5005
R12541 GNDA.n2076 GNDA.n1967 4.5005
R12542 GNDA.n2080 GNDA.n2077 4.5005
R12543 GNDA.n2081 GNDA.n1966 4.5005
R12544 GNDA.n2085 GNDA.n2084 4.5005
R12545 GNDA.n2086 GNDA.n1965 4.5005
R12546 GNDA.n2090 GNDA.n2087 4.5005
R12547 GNDA.n2091 GNDA.n1964 4.5005
R12548 GNDA.n2095 GNDA.n2094 4.5005
R12549 GNDA.n1822 GNDA.n1821 4.5005
R12550 GNDA.n1825 GNDA.n1824 4.5005
R12551 GNDA.n1826 GNDA.n776 4.5005
R12552 GNDA.n1830 GNDA.n1827 4.5005
R12553 GNDA.n1831 GNDA.n775 4.5005
R12554 GNDA.n1835 GNDA.n1834 4.5005
R12555 GNDA.n1836 GNDA.n774 4.5005
R12556 GNDA.n1840 GNDA.n1837 4.5005
R12557 GNDA.n1841 GNDA.n773 4.5005
R12558 GNDA.n1845 GNDA.n1844 4.5005
R12559 GNDA.n1846 GNDA.n772 4.5005
R12560 GNDA.n1850 GNDA.n1847 4.5005
R12561 GNDA.n1851 GNDA.n771 4.5005
R12562 GNDA.n1855 GNDA.n1854 4.5005
R12563 GNDA.n1856 GNDA.n770 4.5005
R12564 GNDA.n1860 GNDA.n1857 4.5005
R12565 GNDA.n1861 GNDA.n769 4.5005
R12566 GNDA.n1865 GNDA.n1864 4.5005
R12567 GNDA.n1866 GNDA.n768 4.5005
R12568 GNDA.n1870 GNDA.n1867 4.5005
R12569 GNDA.n1871 GNDA.n767 4.5005
R12570 GNDA.n1875 GNDA.n1874 4.5005
R12571 GNDA.n1876 GNDA.n766 4.5005
R12572 GNDA.n1880 GNDA.n1877 4.5005
R12573 GNDA.n1881 GNDA.n765 4.5005
R12574 GNDA.n1885 GNDA.n1884 4.5005
R12575 GNDA.n1886 GNDA.n764 4.5005
R12576 GNDA.n1890 GNDA.n1887 4.5005
R12577 GNDA.n1891 GNDA.n763 4.5005
R12578 GNDA.n1895 GNDA.n1894 4.5005
R12579 GNDA.n1896 GNDA.n762 4.5005
R12580 GNDA.n1900 GNDA.n1897 4.5005
R12581 GNDA.n1901 GNDA.n761 4.5005
R12582 GNDA.n1905 GNDA.n1904 4.5005
R12583 GNDA.n1906 GNDA.n760 4.5005
R12584 GNDA.n1910 GNDA.n1907 4.5005
R12585 GNDA.n1911 GNDA.n759 4.5005
R12586 GNDA.n1915 GNDA.n1914 4.5005
R12587 GNDA.n1916 GNDA.n758 4.5005
R12588 GNDA.n1920 GNDA.n1917 4.5005
R12589 GNDA.n1921 GNDA.n757 4.5005
R12590 GNDA.n1925 GNDA.n1924 4.5005
R12591 GNDA.n1926 GNDA.n756 4.5005
R12592 GNDA.n1930 GNDA.n1927 4.5005
R12593 GNDA.n1931 GNDA.n755 4.5005
R12594 GNDA.n1935 GNDA.n1934 4.5005
R12595 GNDA.n1688 GNDA.n1687 4.5005
R12596 GNDA.n1525 GNDA.n1524 4.5005
R12597 GNDA.n1571 GNDA.n1526 4.5005
R12598 GNDA.n1572 GNDA.n1527 4.5005
R12599 GNDA.n1573 GNDA.n1528 4.5005
R12600 GNDA.n1574 GNDA.n1529 4.5005
R12601 GNDA.n1575 GNDA.n1530 4.5005
R12602 GNDA.n1576 GNDA.n1531 4.5005
R12603 GNDA.n1577 GNDA.n1532 4.5005
R12604 GNDA.n1578 GNDA.n1533 4.5005
R12605 GNDA.n1579 GNDA.n1534 4.5005
R12606 GNDA.n1580 GNDA.n1535 4.5005
R12607 GNDA.n1581 GNDA.n1536 4.5005
R12608 GNDA.n1582 GNDA.n1537 4.5005
R12609 GNDA.n1583 GNDA.n1538 4.5005
R12610 GNDA.n1584 GNDA.n1539 4.5005
R12611 GNDA.n1585 GNDA.n1540 4.5005
R12612 GNDA.n1586 GNDA.n1541 4.5005
R12613 GNDA.n1587 GNDA.n1542 4.5005
R12614 GNDA.n1588 GNDA.n1543 4.5005
R12615 GNDA.n1589 GNDA.n1544 4.5005
R12616 GNDA.n1590 GNDA.n1545 4.5005
R12617 GNDA.n1591 GNDA.n1546 4.5005
R12618 GNDA.n1592 GNDA.n1547 4.5005
R12619 GNDA.n1593 GNDA.n1548 4.5005
R12620 GNDA.n1594 GNDA.n1549 4.5005
R12621 GNDA.n1595 GNDA.n1550 4.5005
R12622 GNDA.n1596 GNDA.n1551 4.5005
R12623 GNDA.n1597 GNDA.n1552 4.5005
R12624 GNDA.n1598 GNDA.n1553 4.5005
R12625 GNDA.n1599 GNDA.n1554 4.5005
R12626 GNDA.n1600 GNDA.n1555 4.5005
R12627 GNDA.n1601 GNDA.n1556 4.5005
R12628 GNDA.n1602 GNDA.n1557 4.5005
R12629 GNDA.n1603 GNDA.n1558 4.5005
R12630 GNDA.n1604 GNDA.n1559 4.5005
R12631 GNDA.n1605 GNDA.n1560 4.5005
R12632 GNDA.n1606 GNDA.n1561 4.5005
R12633 GNDA.n1607 GNDA.n1562 4.5005
R12634 GNDA.n1608 GNDA.n1563 4.5005
R12635 GNDA.n1609 GNDA.n1564 4.5005
R12636 GNDA.n1610 GNDA.n1565 4.5005
R12637 GNDA.n1611 GNDA.n1566 4.5005
R12638 GNDA.n1612 GNDA.n1567 4.5005
R12639 GNDA.n1613 GNDA.n1568 4.5005
R12640 GNDA.n1614 GNDA.n1569 4.5005
R12641 GNDA.n1517 GNDA.n1516 4.5005
R12642 GNDA.n792 GNDA.n791 4.5005
R12643 GNDA.n1402 GNDA.n1401 4.5005
R12644 GNDA.n1406 GNDA.n1403 4.5005
R12645 GNDA.n1407 GNDA.n1400 4.5005
R12646 GNDA.n1411 GNDA.n1410 4.5005
R12647 GNDA.n1412 GNDA.n1399 4.5005
R12648 GNDA.n1416 GNDA.n1413 4.5005
R12649 GNDA.n1417 GNDA.n1398 4.5005
R12650 GNDA.n1421 GNDA.n1420 4.5005
R12651 GNDA.n1422 GNDA.n1397 4.5005
R12652 GNDA.n1426 GNDA.n1423 4.5005
R12653 GNDA.n1427 GNDA.n1396 4.5005
R12654 GNDA.n1431 GNDA.n1430 4.5005
R12655 GNDA.n1432 GNDA.n1395 4.5005
R12656 GNDA.n1436 GNDA.n1433 4.5005
R12657 GNDA.n1437 GNDA.n1394 4.5005
R12658 GNDA.n1441 GNDA.n1440 4.5005
R12659 GNDA.n1442 GNDA.n1393 4.5005
R12660 GNDA.n1446 GNDA.n1443 4.5005
R12661 GNDA.n1447 GNDA.n1392 4.5005
R12662 GNDA.n1451 GNDA.n1450 4.5005
R12663 GNDA.n1452 GNDA.n1391 4.5005
R12664 GNDA.n1456 GNDA.n1453 4.5005
R12665 GNDA.n1457 GNDA.n1390 4.5005
R12666 GNDA.n1461 GNDA.n1460 4.5005
R12667 GNDA.n1462 GNDA.n1389 4.5005
R12668 GNDA.n1466 GNDA.n1463 4.5005
R12669 GNDA.n1467 GNDA.n1388 4.5005
R12670 GNDA.n1471 GNDA.n1470 4.5005
R12671 GNDA.n1472 GNDA.n1387 4.5005
R12672 GNDA.n1476 GNDA.n1473 4.5005
R12673 GNDA.n1477 GNDA.n1386 4.5005
R12674 GNDA.n1481 GNDA.n1480 4.5005
R12675 GNDA.n1482 GNDA.n1385 4.5005
R12676 GNDA.n1486 GNDA.n1483 4.5005
R12677 GNDA.n1487 GNDA.n1384 4.5005
R12678 GNDA.n1491 GNDA.n1490 4.5005
R12679 GNDA.n1492 GNDA.n1383 4.5005
R12680 GNDA.n1496 GNDA.n1493 4.5005
R12681 GNDA.n1497 GNDA.n1382 4.5005
R12682 GNDA.n1501 GNDA.n1500 4.5005
R12683 GNDA.n1502 GNDA.n1381 4.5005
R12684 GNDA.n1506 GNDA.n1503 4.5005
R12685 GNDA.n1507 GNDA.n1380 4.5005
R12686 GNDA.n1511 GNDA.n1510 4.5005
R12687 GNDA.n1239 GNDA.n1215 4.5005
R12688 GNDA.n1241 GNDA.n1240 4.5005
R12689 GNDA.n1244 GNDA.n1214 4.5005
R12690 GNDA.n1248 GNDA.n1247 4.5005
R12691 GNDA.n1249 GNDA.n1213 4.5005
R12692 GNDA.n1251 GNDA.n1250 4.5005
R12693 GNDA.n1254 GNDA.n1212 4.5005
R12694 GNDA.n1258 GNDA.n1257 4.5005
R12695 GNDA.n1259 GNDA.n1211 4.5005
R12696 GNDA.n1261 GNDA.n1260 4.5005
R12697 GNDA.n1264 GNDA.n1210 4.5005
R12698 GNDA.n1268 GNDA.n1267 4.5005
R12699 GNDA.n1269 GNDA.n1209 4.5005
R12700 GNDA.n1271 GNDA.n1270 4.5005
R12701 GNDA.n1274 GNDA.n1208 4.5005
R12702 GNDA.n1278 GNDA.n1277 4.5005
R12703 GNDA.n1279 GNDA.n1207 4.5005
R12704 GNDA.n1281 GNDA.n1280 4.5005
R12705 GNDA.n1284 GNDA.n1206 4.5005
R12706 GNDA.n1288 GNDA.n1287 4.5005
R12707 GNDA.n1289 GNDA.n1205 4.5005
R12708 GNDA.n1291 GNDA.n1290 4.5005
R12709 GNDA.n1294 GNDA.n1204 4.5005
R12710 GNDA.n1298 GNDA.n1297 4.5005
R12711 GNDA.n1299 GNDA.n1203 4.5005
R12712 GNDA.n1301 GNDA.n1300 4.5005
R12713 GNDA.n1304 GNDA.n1202 4.5005
R12714 GNDA.n1308 GNDA.n1307 4.5005
R12715 GNDA.n1309 GNDA.n1201 4.5005
R12716 GNDA.n1311 GNDA.n1310 4.5005
R12717 GNDA.n1314 GNDA.n1200 4.5005
R12718 GNDA.n1318 GNDA.n1317 4.5005
R12719 GNDA.n1319 GNDA.n1199 4.5005
R12720 GNDA.n1321 GNDA.n1320 4.5005
R12721 GNDA.n1324 GNDA.n1198 4.5005
R12722 GNDA.n1328 GNDA.n1327 4.5005
R12723 GNDA.n1329 GNDA.n1197 4.5005
R12724 GNDA.n1331 GNDA.n1330 4.5005
R12725 GNDA.n1334 GNDA.n1196 4.5005
R12726 GNDA.n1338 GNDA.n1337 4.5005
R12727 GNDA.n1339 GNDA.n1195 4.5005
R12728 GNDA.n1341 GNDA.n1340 4.5005
R12729 GNDA.n1344 GNDA.n1194 4.5005
R12730 GNDA.n1347 GNDA.n1346 4.5005
R12731 GNDA.n1348 GNDA.n1192 4.5005
R12732 GNDA.n1351 GNDA.n1350 4.5005
R12733 GNDA.n1225 GNDA.n1223 4.5005
R12734 GNDA.n1227 GNDA.n1226 4.5005
R12735 GNDA.n1226 GNDA.n1225 4.5005
R12736 GNDA.n1230 GNDA.n1228 4.5005
R12737 GNDA.n1232 GNDA.n1231 4.5005
R12738 GNDA.n1231 GNDA.n1230 4.5005
R12739 GNDA.n1237 GNDA.n1233 4.5005
R12740 GNDA.n1238 GNDA.n789 4.5005
R12741 GNDA.n1238 GNDA.n1237 4.5005
R12742 GNDA.n1522 GNDA.n1521 4.5005
R12743 GNDA.n1521 GNDA.n1520 4.5005
R12744 GNDA.n1520 GNDA.n790 4.5005
R12745 GNDA.n1693 GNDA.n1692 4.5005
R12746 GNDA.n1692 GNDA.n1691 4.5005
R12747 GNDA.n1691 GNDA.n1523 4.5005
R12748 GNDA.n1816 GNDA.n723 4.5005
R12749 GNDA.n1817 GNDA.n1816 4.5005
R12750 GNDA.n1818 GNDA.n1817 4.5005
R12751 GNDA.n2106 GNDA.n2105 4.5005
R12752 GNDA.n2105 GNDA.n2104 4.5005
R12753 GNDA.n2104 GNDA.n724 4.5005
R12754 GNDA.n2280 GNDA.n2279 4.5005
R12755 GNDA.n2279 GNDA.n2278 4.5005
R12756 GNDA.n2278 GNDA.n2110 4.5005
R12757 GNDA.n2569 GNDA.n2568 4.5005
R12758 GNDA.n2568 GNDA.n2567 4.5005
R12759 GNDA.n2567 GNDA.n661 4.5005
R12760 GNDA.n2740 GNDA.n2739 4.5005
R12761 GNDA.n2739 GNDA.n2738 4.5005
R12762 GNDA.n2738 GNDA.n2570 4.5005
R12763 GNDA.n2741 GNDA.n649 4.5005
R12764 GNDA.n2742 GNDA.n2741 4.5005
R12765 GNDA.n2743 GNDA.n2742 4.5005
R12766 GNDA.n2915 GNDA.n594 4.5005
R12767 GNDA.n2916 GNDA.n2915 4.5005
R12768 GNDA.n2917 GNDA.n2916 4.5005
R12769 GNDA.n3205 GNDA.n3204 4.5005
R12770 GNDA.n3204 GNDA.n3203 4.5005
R12771 GNDA.n3203 GNDA.n595 4.5005
R12772 GNDA.n3376 GNDA.n3207 4.5005
R12773 GNDA.n3379 GNDA.n3207 4.5005
R12774 GNDA.n3379 GNDA.n3206 4.5005
R12775 GNDA.n5013 GNDA.n5010 4.5005
R12776 GNDA.n5014 GNDA.n5013 4.5005
R12777 GNDA.n5015 GNDA.n5014 4.5005
R12778 GNDA.n5006 GNDA.n404 4.5005
R12779 GNDA.n5009 GNDA.n404 4.5005
R12780 GNDA.n5009 GNDA.n403 4.5005
R12781 GNDA.n4994 GNDA.n578 4.5005
R12782 GNDA.n4997 GNDA.n578 4.5005
R12783 GNDA.n4997 GNDA.n577 4.5005
R12784 GNDA.n4990 GNDA.n583 4.5005
R12785 GNDA.n4993 GNDA.n583 4.5005
R12786 GNDA.n4993 GNDA.n582 4.5005
R12787 GNDA.n3681 GNDA.n576 4.5005
R12788 GNDA.n3682 GNDA.n3681 4.5005
R12789 GNDA.n3683 GNDA.n3682 4.5005
R12790 GNDA.n4982 GNDA.n3435 4.5005
R12791 GNDA.n4985 GNDA.n3435 4.5005
R12792 GNDA.n4985 GNDA.n3434 4.5005
R12793 GNDA.n4978 GNDA.n3440 4.5005
R12794 GNDA.n4981 GNDA.n3440 4.5005
R12795 GNDA.n4981 GNDA.n3439 4.5005
R12796 GNDA.n4974 GNDA.n3445 4.5005
R12797 GNDA.n4977 GNDA.n3445 4.5005
R12798 GNDA.n4977 GNDA.n3444 4.5005
R12799 GNDA.n4970 GNDA.n3450 4.5005
R12800 GNDA.n4973 GNDA.n3450 4.5005
R12801 GNDA.n4973 GNDA.n3449 4.5005
R12802 GNDA.n4966 GNDA.n3455 4.5005
R12803 GNDA.n4969 GNDA.n3455 4.5005
R12804 GNDA.n4969 GNDA.n3454 4.5005
R12805 GNDA.n1813 GNDA.n1694 4.5005
R12806 GNDA.n1815 GNDA.n1814 4.5005
R12807 GNDA.n1814 GNDA.n1813 4.5005
R12808 GNDA.n4986 GNDA.n3431 4.5005
R12809 GNDA.n4989 GNDA.n3431 4.5005
R12810 GNDA.n4989 GNDA.n587 4.5005
R12811 GNDA.n5281 GNDA.n323 4.5005
R12812 GNDA.n5281 GNDA.n5280 4.5005
R12813 GNDA.n5280 GNDA.n325 4.5005
R12814 GNDA.n6950 GNDA.n6949 4.5005
R12815 GNDA.n6943 GNDA.n6942 4.5005
R12816 GNDA.n5356 GNDA.n5354 4.5005
R12817 GNDA.n6781 GNDA.n6652 4.5005
R12818 GNDA.n6778 GNDA.n5355 4.5005
R12819 GNDA.n6781 GNDA.n5355 4.5005
R12820 GNDA.n7135 GNDA.n7131 4.5005
R12821 GNDA.n7139 GNDA.n7138 4.5005
R12822 GNDA.n7140 GNDA.n7128 4.5005
R12823 GNDA.n7142 GNDA.n7141 4.5005
R12824 GNDA.n7143 GNDA.n7127 4.5005
R12825 GNDA.n7147 GNDA.n7146 4.5005
R12826 GNDA.n7148 GNDA.n7124 4.5005
R12827 GNDA.n7150 GNDA.n7149 4.5005
R12828 GNDA.n7151 GNDA.n7123 4.5005
R12829 GNDA.n7155 GNDA.n7154 4.5005
R12830 GNDA.n7156 GNDA.n7120 4.5005
R12831 GNDA.n7158 GNDA.n7157 4.5005
R12832 GNDA.n7159 GNDA.n7119 4.5005
R12833 GNDA.n7163 GNDA.n7162 4.5005
R12834 GNDA.n7164 GNDA.n7116 4.5005
R12835 GNDA.n7166 GNDA.n7165 4.5005
R12836 GNDA.n7167 GNDA.n7115 4.5005
R12837 GNDA.n7171 GNDA.n7170 4.5005
R12838 GNDA.n7172 GNDA.n7112 4.5005
R12839 GNDA.n7174 GNDA.n7173 4.5005
R12840 GNDA.n7175 GNDA.n7111 4.5005
R12841 GNDA.n7179 GNDA.n7178 4.5005
R12842 GNDA.n7180 GNDA.n7108 4.5005
R12843 GNDA.n7182 GNDA.n7181 4.5005
R12844 GNDA.n7183 GNDA.n7107 4.5005
R12845 GNDA.n7187 GNDA.n7186 4.5005
R12846 GNDA.n7188 GNDA.n7104 4.5005
R12847 GNDA.n7190 GNDA.n7189 4.5005
R12848 GNDA.n7191 GNDA.n7103 4.5005
R12849 GNDA.n7195 GNDA.n7194 4.5005
R12850 GNDA.n7196 GNDA.n7100 4.5005
R12851 GNDA.n7198 GNDA.n7197 4.5005
R12852 GNDA.n7199 GNDA.n7099 4.5005
R12853 GNDA.n7203 GNDA.n7202 4.5005
R12854 GNDA.n7204 GNDA.n7096 4.5005
R12855 GNDA.n7206 GNDA.n7205 4.5005
R12856 GNDA.n7207 GNDA.n7095 4.5005
R12857 GNDA.n7211 GNDA.n7210 4.5005
R12858 GNDA.n7212 GNDA.n7092 4.5005
R12859 GNDA.n7214 GNDA.n7213 4.5005
R12860 GNDA.n7215 GNDA.n7091 4.5005
R12861 GNDA.n7219 GNDA.n7218 4.5005
R12862 GNDA.n7220 GNDA.n7090 4.5005
R12863 GNDA.n7222 GNDA.n7221 4.5005
R12864 GNDA.n96 GNDA.n95 4.5005
R12865 GNDA.n7228 GNDA.n7227 4.5005
R12866 GNDA.n6657 GNDA.n6656 4.5005
R12867 GNDA.n7233 GNDA.n90 4.5005
R12868 GNDA.n7232 GNDA.n7231 4.5005
R12869 GNDA.n7233 GNDA.n7232 4.5005
R12870 GNDA.n263 GNDA.n262 4.5005
R12871 GNDA.n266 GNDA.n265 4.5005
R12872 GNDA.n150 GNDA.n146 4.5005
R12873 GNDA.n154 GNDA.n151 4.5005
R12874 GNDA.n155 GNDA.n145 4.5005
R12875 GNDA.n159 GNDA.n158 4.5005
R12876 GNDA.n160 GNDA.n144 4.5005
R12877 GNDA.n164 GNDA.n161 4.5005
R12878 GNDA.n165 GNDA.n143 4.5005
R12879 GNDA.n169 GNDA.n168 4.5005
R12880 GNDA.n170 GNDA.n142 4.5005
R12881 GNDA.n174 GNDA.n171 4.5005
R12882 GNDA.n175 GNDA.n141 4.5005
R12883 GNDA.n179 GNDA.n178 4.5005
R12884 GNDA.n180 GNDA.n140 4.5005
R12885 GNDA.n184 GNDA.n181 4.5005
R12886 GNDA.n185 GNDA.n139 4.5005
R12887 GNDA.n189 GNDA.n188 4.5005
R12888 GNDA.n190 GNDA.n138 4.5005
R12889 GNDA.n194 GNDA.n191 4.5005
R12890 GNDA.n195 GNDA.n137 4.5005
R12891 GNDA.n199 GNDA.n198 4.5005
R12892 GNDA.n200 GNDA.n136 4.5005
R12893 GNDA.n204 GNDA.n201 4.5005
R12894 GNDA.n205 GNDA.n135 4.5005
R12895 GNDA.n209 GNDA.n208 4.5005
R12896 GNDA.n210 GNDA.n134 4.5005
R12897 GNDA.n214 GNDA.n211 4.5005
R12898 GNDA.n215 GNDA.n133 4.5005
R12899 GNDA.n219 GNDA.n218 4.5005
R12900 GNDA.n220 GNDA.n132 4.5005
R12901 GNDA.n224 GNDA.n221 4.5005
R12902 GNDA.n225 GNDA.n131 4.5005
R12903 GNDA.n229 GNDA.n228 4.5005
R12904 GNDA.n230 GNDA.n130 4.5005
R12905 GNDA.n234 GNDA.n231 4.5005
R12906 GNDA.n235 GNDA.n129 4.5005
R12907 GNDA.n239 GNDA.n238 4.5005
R12908 GNDA.n240 GNDA.n128 4.5005
R12909 GNDA.n244 GNDA.n241 4.5005
R12910 GNDA.n245 GNDA.n127 4.5005
R12911 GNDA.n249 GNDA.n248 4.5005
R12912 GNDA.n250 GNDA.n126 4.5005
R12913 GNDA.n254 GNDA.n251 4.5005
R12914 GNDA.n255 GNDA.n125 4.5005
R12915 GNDA.n259 GNDA.n258 4.5005
R12916 GNDA.n260 GNDA.n124 4.5005
R12917 GNDA.n7063 GNDA.n7062 4.5005
R12918 GNDA.n6297 GNDA.n6296 4.26717
R12919 GNDA.n6296 GNDA.n6270 4.26717
R12920 GNDA.n6290 GNDA.n6270 4.26717
R12921 GNDA.n6290 GNDA.n6289 4.26717
R12922 GNDA.n6289 GNDA.n6288 4.26717
R12923 GNDA.n6288 GNDA.n6276 4.26717
R12924 GNDA.n6282 GNDA.n6276 4.26717
R12925 GNDA.n6282 GNDA.n6281 4.26717
R12926 GNDA.n6281 GNDA.n70 4.26717
R12927 GNDA.n7468 GNDA.n70 4.26717
R12928 GNDA.n7468 GNDA.n67 4.26717
R12929 GNDA.n6209 GNDA.n5436 4.26717
R12930 GNDA.n6204 GNDA.n5436 4.26717
R12931 GNDA.n6204 GNDA.n6203 4.26717
R12932 GNDA.n6203 GNDA.n6181 4.26717
R12933 GNDA.n6198 GNDA.n6181 4.26717
R12934 GNDA.n6198 GNDA.n6197 4.26717
R12935 GNDA.n6197 GNDA.n6196 4.26717
R12936 GNDA.n6196 GNDA.n6191 4.26717
R12937 GNDA.n6191 GNDA.n5391 4.26717
R12938 GNDA.n6917 GNDA.n5391 4.26717
R12939 GNDA.n6917 GNDA.n5389 4.26717
R12940 GNDA.n5834 GNDA.n5526 4.26717
R12941 GNDA.n5834 GNDA.n5529 4.26717
R12942 GNDA.n5564 GNDA.n5529 4.26717
R12943 GNDA.n5564 GNDA.n5563 4.26717
R12944 GNDA.n5563 GNDA.n5562 4.26717
R12945 GNDA.n5562 GNDA.n5559 4.26717
R12946 GNDA.n5559 GNDA.n5558 4.26717
R12947 GNDA.n5558 GNDA.n5555 4.26717
R12948 GNDA.n5555 GNDA.n5554 4.26717
R12949 GNDA.n5554 GNDA.n5551 4.26717
R12950 GNDA.n5551 GNDA.n5550 4.26717
R12951 GNDA.n7293 GNDA.n7292 4.26717
R12952 GNDA.n7292 GNDA.n7252 4.26717
R12953 GNDA.n7286 GNDA.n7252 4.26717
R12954 GNDA.n7286 GNDA.n7285 4.26717
R12955 GNDA.n7285 GNDA.n7284 4.26717
R12956 GNDA.n7284 GNDA.n7260 4.26717
R12957 GNDA.n7278 GNDA.n7260 4.26717
R12958 GNDA.n7278 GNDA.n7277 4.26717
R12959 GNDA.n7277 GNDA.n7276 4.26717
R12960 GNDA.n7276 GNDA.n7271 4.26717
R12961 GNDA.n7271 GNDA.n59 4.26717
R12962 GNDA.n5806 GNDA.n5577 4.26717
R12963 GNDA.n5806 GNDA.n5580 4.26717
R12964 GNDA.n5615 GNDA.n5580 4.26717
R12965 GNDA.n5615 GNDA.n5614 4.26717
R12966 GNDA.n5614 GNDA.n5613 4.26717
R12967 GNDA.n5613 GNDA.n5610 4.26717
R12968 GNDA.n5610 GNDA.n5609 4.26717
R12969 GNDA.n5609 GNDA.n5606 4.26717
R12970 GNDA.n5606 GNDA.n5605 4.26717
R12971 GNDA.n5605 GNDA.n5602 4.26717
R12972 GNDA.n5602 GNDA.n5601 4.26717
R12973 GNDA.n6149 GNDA.n6074 4.26717
R12974 GNDA.n6144 GNDA.n6074 4.26717
R12975 GNDA.n6144 GNDA.n6143 4.26717
R12976 GNDA.n6143 GNDA.n6125 4.26717
R12977 GNDA.n6138 GNDA.n6125 4.26717
R12978 GNDA.n6138 GNDA.n6137 4.26717
R12979 GNDA.n6137 GNDA.n6136 4.26717
R12980 GNDA.n6136 GNDA.n6131 4.26717
R12981 GNDA.n6131 GNDA.n5374 4.26717
R12982 GNDA.n6927 GNDA.n5374 4.26717
R12983 GNDA.n6927 GNDA.n5370 4.26717
R12984 GNDA.t2 GNDA.t145 4.19522
R12985 GNDA.n6297 GNDA.n81 3.93531
R12986 GNDA.n6210 GNDA.n6209 3.93531
R12987 GNDA.n5526 GNDA.n5524 3.93531
R12988 GNDA.n7294 GNDA.n7293 3.93531
R12989 GNDA.n5577 GNDA.n61 3.93531
R12990 GNDA.n6149 GNDA.n6073 3.93531
R12991 GNDA.t322 GNDA.t46 3.93305
R12992 GNDA.n5305 GNDA.n320 3.85122
R12993 GNDA.n6448 GNDA.n6345 3.7893
R12994 GNDA.n6445 GNDA.n6444 3.7893
R12995 GNDA.n6355 GNDA.n6346 3.7893
R12996 GNDA.n6360 GNDA.n6358 3.7893
R12997 GNDA.n6365 GNDA.n6361 3.7893
R12998 GNDA.n6369 GNDA.n6354 3.7893
R12999 GNDA.n6374 GNDA.n6372 3.7893
R13000 GNDA.n6373 GNDA.n56 3.7893
R13001 GNDA.n6543 GNDA.n6324 3.7893
R13002 GNDA.n6540 GNDA.n6539 3.7893
R13003 GNDA.n6456 GNDA.n6325 3.7893
R13004 GNDA.n6461 GNDA.n6459 3.7893
R13005 GNDA.n6466 GNDA.n6462 3.7893
R13006 GNDA.n6473 GNDA.n6472 3.7893
R13007 GNDA.n6476 GNDA.n6455 3.7893
R13008 GNDA.n6481 GNDA.n6477 3.7893
R13009 GNDA.n6974 GNDA.n5344 3.7893
R13010 GNDA.n6973 GNDA.n5345 3.7893
R13011 GNDA.n6961 GNDA.n6960 3.7893
R13012 GNDA.n6967 GNDA.n6966 3.7893
R13013 GNDA.n6963 GNDA.n6962 3.7893
R13014 GNDA.n6838 GNDA.n5323 3.7893
R13015 GNDA.n6839 GNDA.n6837 3.7893
R13016 GNDA.n6848 GNDA.n6846 3.7893
R13017 GNDA.n6820 GNDA.n6819 3.7893
R13018 GNDA.n6816 GNDA.n6576 3.7893
R13019 GNDA.n6815 GNDA.n6641 3.7893
R13020 GNDA.n6798 GNDA.n6797 3.7893
R13021 GNDA.n6809 GNDA.n6808 3.7893
R13022 GNDA.n6801 GNDA.n5399 3.7893
R13023 GNDA.n6830 GNDA.n6828 3.7893
R13024 GNDA.n6829 GNDA.n5395 3.7893
R13025 GNDA.n5743 GNDA.n5718 3.7893
R13026 GNDA.n5742 GNDA.n5739 3.7893
R13027 GNDA.n5738 GNDA.n5719 3.7893
R13028 GNDA.n5735 GNDA.n5734 3.7893
R13029 GNDA.n5731 GNDA.n5720 3.7893
R13030 GNDA.n5724 GNDA.n5721 3.7893
R13031 GNDA.n5748 GNDA.n5643 3.7893
R13032 GNDA.n5749 GNDA.n5642 3.7893
R13033 GNDA.n6065 GNDA.n5452 3.7893
R13034 GNDA.n6062 GNDA.n6061 3.7893
R13035 GNDA.n5488 GNDA.n5454 3.7893
R13036 GNDA.n5506 GNDA.n5505 3.7893
R13037 GNDA.n5503 GNDA.n5502 3.7893
R13038 GNDA.n5498 GNDA.n5491 3.7893
R13039 GNDA.n5495 GNDA.n5494 3.7893
R13040 GNDA.n6003 GNDA.n5474 3.7893
R13041 GNDA.n5994 GNDA.n5993 3.7893
R13042 GNDA.n5990 GNDA.n5885 3.7893
R13043 GNDA.n5989 GNDA.n5888 3.7893
R13044 GNDA.n5986 GNDA.n5985 3.7893
R13045 GNDA.n5912 GNDA.n5889 3.7893
R13046 GNDA.n5921 GNDA.n5920 3.7893
R13047 GNDA.n5924 GNDA.n5911 3.7893
R13048 GNDA.n5929 GNDA.n5925 3.7893
R13049 GNDA.n6741 GNDA.n6740 3.7893
R13050 GNDA.n6751 GNDA.n6670 3.7893
R13051 GNDA.n6750 GNDA.n6668 3.7893
R13052 GNDA.n6757 GNDA.n6667 3.7893
R13053 GNDA.n6760 GNDA.n6759 3.7893
R13054 GNDA.n7020 GNDA.n294 3.7893
R13055 GNDA.n293 GNDA.n290 3.7893
R13056 GNDA.n7029 GNDA.n7028 3.7893
R13057 GNDA.n7486 GNDA.n22 3.7893
R13058 GNDA.n7485 GNDA.n23 3.7893
R13059 GNDA.n33 GNDA.n32 3.7893
R13060 GNDA.n39 GNDA.n38 3.7893
R13061 GNDA.n35 GNDA.n34 3.7893
R13062 GNDA.n7373 GNDA.n1 3.7893
R13063 GNDA.n7378 GNDA.n7376 3.7893
R13064 GNDA.n7379 GNDA.n7372 3.7893
R13065 GNDA.n6368 GNDA 3.7381
R13066 GNDA.n6469 GNDA 3.7381
R13067 GNDA GNDA.n6979 3.7381
R13068 GNDA.n6802 GNDA 3.7381
R13069 GNDA GNDA.n5727 3.7381
R13070 GNDA.n5499 GNDA 3.7381
R13071 GNDA.n5917 GNDA 3.7381
R13072 GNDA.n7021 GNDA 3.7381
R13073 GNDA GNDA.n7491 3.7381
R13074 GNDA.n3389 GNDA.n3384 3.65764
R13075 GNDA.n3389 GNDA.n3388 3.65764
R13076 GNDA.n1731 GNDA.n1725 3.65764
R13077 GNDA.n1731 GNDA.n1730 3.65764
R13078 GNDA.n1349 GNDA.n1167 3.50398
R13079 GNDA.n149 GNDA.n99 3.47871
R13080 GNDA.n5271 GNDA.n5270 3.47821
R13081 GNDA.n4958 GNDA.n4957 3.47821
R13082 GNDA.n4798 GNDA.n4797 3.47821
R13083 GNDA.n4632 GNDA.n4631 3.47821
R13084 GNDA.n4466 GNDA.n4465 3.47821
R13085 GNDA.n4300 GNDA.n4299 3.47821
R13086 GNDA.n3802 GNDA.n3801 3.47821
R13087 GNDA.n4134 GNDA.n4133 3.47821
R13088 GNDA.n3968 GNDA.n3967 3.47821
R13089 GNDA.n3603 GNDA.n3602 3.47821
R13090 GNDA.n497 GNDA.n496 3.47821
R13091 GNDA.n5134 GNDA.n5133 3.47821
R13092 GNDA.n3300 GNDA.n3299 3.47821
R13093 GNDA.n3196 GNDA.n3195 3.47821
R13094 GNDA.n3036 GNDA.n3035 3.47821
R13095 GNDA.n2400 GNDA.n2399 3.47821
R13096 GNDA.n2862 GNDA.n2861 3.47821
R13097 GNDA.n2663 GNDA.n2662 3.47821
R13098 GNDA.n2560 GNDA.n2559 3.47821
R13099 GNDA.n2203 GNDA.n2202 3.47821
R13100 GNDA.n2097 GNDA.n2096 3.47821
R13101 GNDA.n1937 GNDA.n1936 3.47821
R13102 GNDA.n1616 GNDA.n1615 3.47821
R13103 GNDA.n1513 GNDA.n1512 3.47821
R13104 GNDA.n7132 GNDA.n7066 3.47821
R13105 GNDA.n1215 GNDA.n1168 3.43627
R13106 GNDA.n3680 GNDA.t100 3.42907
R13107 GNDA.n3680 GNDA.t128 3.42907
R13108 GNDA.n3677 GNDA.t48 3.42907
R13109 GNDA.n3677 GNDA.t8 3.42907
R13110 GNDA.n714 GNDA.t269 3.42907
R13111 GNDA.n714 GNDA.t63 3.42907
R13112 GNDA.n718 GNDA.t289 3.42907
R13113 GNDA.n718 GNDA.t265 3.42907
R13114 GNDA.t279 GNDA.t32 3.41135
R13115 GNDA.n5137 GNDA.n5136 3.4105
R13116 GNDA.n5268 GNDA.n5267 3.4105
R13117 GNDA.n5266 GNDA.n5265 3.4105
R13118 GNDA.n5264 GNDA.n5263 3.4105
R13119 GNDA.n5262 GNDA.n5139 3.4105
R13120 GNDA.n5258 GNDA.n5257 3.4105
R13121 GNDA.n5256 GNDA.n5255 3.4105
R13122 GNDA.n5254 GNDA.n5253 3.4105
R13123 GNDA.n5252 GNDA.n5141 3.4105
R13124 GNDA.n5248 GNDA.n5247 3.4105
R13125 GNDA.n5246 GNDA.n5245 3.4105
R13126 GNDA.n5244 GNDA.n5243 3.4105
R13127 GNDA.n5242 GNDA.n5143 3.4105
R13128 GNDA.n5238 GNDA.n5237 3.4105
R13129 GNDA.n5236 GNDA.n5235 3.4105
R13130 GNDA.n5234 GNDA.n5233 3.4105
R13131 GNDA.n5232 GNDA.n5145 3.4105
R13132 GNDA.n5228 GNDA.n5227 3.4105
R13133 GNDA.n5226 GNDA.n5225 3.4105
R13134 GNDA.n5224 GNDA.n5223 3.4105
R13135 GNDA.n5222 GNDA.n5147 3.4105
R13136 GNDA.n5218 GNDA.n5217 3.4105
R13137 GNDA.n5216 GNDA.n5215 3.4105
R13138 GNDA.n5214 GNDA.n5213 3.4105
R13139 GNDA.n5212 GNDA.n5149 3.4105
R13140 GNDA.n5208 GNDA.n5207 3.4105
R13141 GNDA.n5206 GNDA.n5205 3.4105
R13142 GNDA.n5204 GNDA.n5203 3.4105
R13143 GNDA.n5202 GNDA.n5151 3.4105
R13144 GNDA.n5198 GNDA.n5197 3.4105
R13145 GNDA.n5196 GNDA.n5195 3.4105
R13146 GNDA.n5194 GNDA.n5193 3.4105
R13147 GNDA.n5192 GNDA.n5153 3.4105
R13148 GNDA.n5188 GNDA.n5187 3.4105
R13149 GNDA.n5186 GNDA.n5185 3.4105
R13150 GNDA.n5184 GNDA.n5183 3.4105
R13151 GNDA.n5182 GNDA.n5155 3.4105
R13152 GNDA.n5178 GNDA.n5177 3.4105
R13153 GNDA.n5176 GNDA.n5175 3.4105
R13154 GNDA.n5174 GNDA.n5173 3.4105
R13155 GNDA.n5172 GNDA.n5157 3.4105
R13156 GNDA.n5168 GNDA.n5167 3.4105
R13157 GNDA.n5166 GNDA.n5165 3.4105
R13158 GNDA.n5164 GNDA.n5163 3.4105
R13159 GNDA.n5162 GNDA.n5159 3.4105
R13160 GNDA.n328 GNDA.n327 3.4105
R13161 GNDA.n5274 GNDA.n5273 3.4105
R13162 GNDA.n4824 GNDA.n4823 3.4105
R13163 GNDA.n4955 GNDA.n4954 3.4105
R13164 GNDA.n4953 GNDA.n4952 3.4105
R13165 GNDA.n4951 GNDA.n4950 3.4105
R13166 GNDA.n4949 GNDA.n4826 3.4105
R13167 GNDA.n4945 GNDA.n4944 3.4105
R13168 GNDA.n4943 GNDA.n4942 3.4105
R13169 GNDA.n4941 GNDA.n4940 3.4105
R13170 GNDA.n4939 GNDA.n4828 3.4105
R13171 GNDA.n4935 GNDA.n4934 3.4105
R13172 GNDA.n4933 GNDA.n4932 3.4105
R13173 GNDA.n4931 GNDA.n4930 3.4105
R13174 GNDA.n4929 GNDA.n4830 3.4105
R13175 GNDA.n4925 GNDA.n4924 3.4105
R13176 GNDA.n4923 GNDA.n4922 3.4105
R13177 GNDA.n4921 GNDA.n4920 3.4105
R13178 GNDA.n4919 GNDA.n4832 3.4105
R13179 GNDA.n4915 GNDA.n4914 3.4105
R13180 GNDA.n4913 GNDA.n4912 3.4105
R13181 GNDA.n4911 GNDA.n4910 3.4105
R13182 GNDA.n4909 GNDA.n4834 3.4105
R13183 GNDA.n4905 GNDA.n4904 3.4105
R13184 GNDA.n4903 GNDA.n4902 3.4105
R13185 GNDA.n4901 GNDA.n4900 3.4105
R13186 GNDA.n4899 GNDA.n4836 3.4105
R13187 GNDA.n4895 GNDA.n4894 3.4105
R13188 GNDA.n4893 GNDA.n4892 3.4105
R13189 GNDA.n4891 GNDA.n4890 3.4105
R13190 GNDA.n4889 GNDA.n4838 3.4105
R13191 GNDA.n4885 GNDA.n4884 3.4105
R13192 GNDA.n4883 GNDA.n4882 3.4105
R13193 GNDA.n4881 GNDA.n4880 3.4105
R13194 GNDA.n4879 GNDA.n4840 3.4105
R13195 GNDA.n4875 GNDA.n4874 3.4105
R13196 GNDA.n4873 GNDA.n4872 3.4105
R13197 GNDA.n4871 GNDA.n4870 3.4105
R13198 GNDA.n4869 GNDA.n4842 3.4105
R13199 GNDA.n4865 GNDA.n4864 3.4105
R13200 GNDA.n4863 GNDA.n4862 3.4105
R13201 GNDA.n4861 GNDA.n4860 3.4105
R13202 GNDA.n4859 GNDA.n4844 3.4105
R13203 GNDA.n4855 GNDA.n4854 3.4105
R13204 GNDA.n4853 GNDA.n4852 3.4105
R13205 GNDA.n4851 GNDA.n4850 3.4105
R13206 GNDA.n4849 GNDA.n4846 3.4105
R13207 GNDA.n3458 GNDA.n3457 3.4105
R13208 GNDA.n4961 GNDA.n4960 3.4105
R13209 GNDA.n4659 GNDA.n4658 3.4105
R13210 GNDA.n4795 GNDA.n4794 3.4105
R13211 GNDA.n4793 GNDA.n4792 3.4105
R13212 GNDA.n4791 GNDA.n4790 3.4105
R13213 GNDA.n4789 GNDA.n4661 3.4105
R13214 GNDA.n4785 GNDA.n4784 3.4105
R13215 GNDA.n4783 GNDA.n4782 3.4105
R13216 GNDA.n4781 GNDA.n4780 3.4105
R13217 GNDA.n4779 GNDA.n4663 3.4105
R13218 GNDA.n4775 GNDA.n4774 3.4105
R13219 GNDA.n4773 GNDA.n4772 3.4105
R13220 GNDA.n4771 GNDA.n4770 3.4105
R13221 GNDA.n4769 GNDA.n4665 3.4105
R13222 GNDA.n4765 GNDA.n4764 3.4105
R13223 GNDA.n4763 GNDA.n4762 3.4105
R13224 GNDA.n4761 GNDA.n4760 3.4105
R13225 GNDA.n4759 GNDA.n4667 3.4105
R13226 GNDA.n4755 GNDA.n4754 3.4105
R13227 GNDA.n4753 GNDA.n4752 3.4105
R13228 GNDA.n4751 GNDA.n4750 3.4105
R13229 GNDA.n4749 GNDA.n4669 3.4105
R13230 GNDA.n4745 GNDA.n4744 3.4105
R13231 GNDA.n4743 GNDA.n4742 3.4105
R13232 GNDA.n4741 GNDA.n4740 3.4105
R13233 GNDA.n4739 GNDA.n4671 3.4105
R13234 GNDA.n4735 GNDA.n4734 3.4105
R13235 GNDA.n4733 GNDA.n4732 3.4105
R13236 GNDA.n4731 GNDA.n4730 3.4105
R13237 GNDA.n4729 GNDA.n4673 3.4105
R13238 GNDA.n4725 GNDA.n4724 3.4105
R13239 GNDA.n4723 GNDA.n4722 3.4105
R13240 GNDA.n4721 GNDA.n4720 3.4105
R13241 GNDA.n4719 GNDA.n4675 3.4105
R13242 GNDA.n4715 GNDA.n4714 3.4105
R13243 GNDA.n4713 GNDA.n4712 3.4105
R13244 GNDA.n4711 GNDA.n4710 3.4105
R13245 GNDA.n4709 GNDA.n4677 3.4105
R13246 GNDA.n4705 GNDA.n4704 3.4105
R13247 GNDA.n4703 GNDA.n4702 3.4105
R13248 GNDA.n4701 GNDA.n4700 3.4105
R13249 GNDA.n4699 GNDA.n4679 3.4105
R13250 GNDA.n4695 GNDA.n4694 3.4105
R13251 GNDA.n4693 GNDA.n4692 3.4105
R13252 GNDA.n4691 GNDA.n4690 3.4105
R13253 GNDA.n4689 GNDA.n4681 3.4105
R13254 GNDA.n4685 GNDA.n4684 3.4105
R13255 GNDA.n4683 GNDA.n4634 3.4105
R13256 GNDA.n4493 GNDA.n4492 3.4105
R13257 GNDA.n4629 GNDA.n4628 3.4105
R13258 GNDA.n4627 GNDA.n4626 3.4105
R13259 GNDA.n4625 GNDA.n4624 3.4105
R13260 GNDA.n4623 GNDA.n4495 3.4105
R13261 GNDA.n4619 GNDA.n4618 3.4105
R13262 GNDA.n4617 GNDA.n4616 3.4105
R13263 GNDA.n4615 GNDA.n4614 3.4105
R13264 GNDA.n4613 GNDA.n4497 3.4105
R13265 GNDA.n4609 GNDA.n4608 3.4105
R13266 GNDA.n4607 GNDA.n4606 3.4105
R13267 GNDA.n4605 GNDA.n4604 3.4105
R13268 GNDA.n4603 GNDA.n4499 3.4105
R13269 GNDA.n4599 GNDA.n4598 3.4105
R13270 GNDA.n4597 GNDA.n4596 3.4105
R13271 GNDA.n4595 GNDA.n4594 3.4105
R13272 GNDA.n4593 GNDA.n4501 3.4105
R13273 GNDA.n4589 GNDA.n4588 3.4105
R13274 GNDA.n4587 GNDA.n4586 3.4105
R13275 GNDA.n4585 GNDA.n4584 3.4105
R13276 GNDA.n4583 GNDA.n4503 3.4105
R13277 GNDA.n4579 GNDA.n4578 3.4105
R13278 GNDA.n4577 GNDA.n4576 3.4105
R13279 GNDA.n4575 GNDA.n4574 3.4105
R13280 GNDA.n4573 GNDA.n4505 3.4105
R13281 GNDA.n4569 GNDA.n4568 3.4105
R13282 GNDA.n4567 GNDA.n4566 3.4105
R13283 GNDA.n4565 GNDA.n4564 3.4105
R13284 GNDA.n4563 GNDA.n4507 3.4105
R13285 GNDA.n4559 GNDA.n4558 3.4105
R13286 GNDA.n4557 GNDA.n4556 3.4105
R13287 GNDA.n4555 GNDA.n4554 3.4105
R13288 GNDA.n4553 GNDA.n4509 3.4105
R13289 GNDA.n4549 GNDA.n4548 3.4105
R13290 GNDA.n4547 GNDA.n4546 3.4105
R13291 GNDA.n4545 GNDA.n4544 3.4105
R13292 GNDA.n4543 GNDA.n4511 3.4105
R13293 GNDA.n4539 GNDA.n4538 3.4105
R13294 GNDA.n4537 GNDA.n4536 3.4105
R13295 GNDA.n4535 GNDA.n4534 3.4105
R13296 GNDA.n4533 GNDA.n4513 3.4105
R13297 GNDA.n4529 GNDA.n4528 3.4105
R13298 GNDA.n4527 GNDA.n4526 3.4105
R13299 GNDA.n4525 GNDA.n4524 3.4105
R13300 GNDA.n4523 GNDA.n4515 3.4105
R13301 GNDA.n4519 GNDA.n4518 3.4105
R13302 GNDA.n4517 GNDA.n4468 3.4105
R13303 GNDA.n4327 GNDA.n4326 3.4105
R13304 GNDA.n4463 GNDA.n4462 3.4105
R13305 GNDA.n4461 GNDA.n4460 3.4105
R13306 GNDA.n4459 GNDA.n4458 3.4105
R13307 GNDA.n4457 GNDA.n4329 3.4105
R13308 GNDA.n4453 GNDA.n4452 3.4105
R13309 GNDA.n4451 GNDA.n4450 3.4105
R13310 GNDA.n4449 GNDA.n4448 3.4105
R13311 GNDA.n4447 GNDA.n4331 3.4105
R13312 GNDA.n4443 GNDA.n4442 3.4105
R13313 GNDA.n4441 GNDA.n4440 3.4105
R13314 GNDA.n4439 GNDA.n4438 3.4105
R13315 GNDA.n4437 GNDA.n4333 3.4105
R13316 GNDA.n4433 GNDA.n4432 3.4105
R13317 GNDA.n4431 GNDA.n4430 3.4105
R13318 GNDA.n4429 GNDA.n4428 3.4105
R13319 GNDA.n4427 GNDA.n4335 3.4105
R13320 GNDA.n4423 GNDA.n4422 3.4105
R13321 GNDA.n4421 GNDA.n4420 3.4105
R13322 GNDA.n4419 GNDA.n4418 3.4105
R13323 GNDA.n4417 GNDA.n4337 3.4105
R13324 GNDA.n4413 GNDA.n4412 3.4105
R13325 GNDA.n4411 GNDA.n4410 3.4105
R13326 GNDA.n4409 GNDA.n4408 3.4105
R13327 GNDA.n4407 GNDA.n4339 3.4105
R13328 GNDA.n4403 GNDA.n4402 3.4105
R13329 GNDA.n4401 GNDA.n4400 3.4105
R13330 GNDA.n4399 GNDA.n4398 3.4105
R13331 GNDA.n4397 GNDA.n4341 3.4105
R13332 GNDA.n4393 GNDA.n4392 3.4105
R13333 GNDA.n4391 GNDA.n4390 3.4105
R13334 GNDA.n4389 GNDA.n4388 3.4105
R13335 GNDA.n4387 GNDA.n4343 3.4105
R13336 GNDA.n4383 GNDA.n4382 3.4105
R13337 GNDA.n4381 GNDA.n4380 3.4105
R13338 GNDA.n4379 GNDA.n4378 3.4105
R13339 GNDA.n4377 GNDA.n4345 3.4105
R13340 GNDA.n4373 GNDA.n4372 3.4105
R13341 GNDA.n4371 GNDA.n4370 3.4105
R13342 GNDA.n4369 GNDA.n4368 3.4105
R13343 GNDA.n4367 GNDA.n4347 3.4105
R13344 GNDA.n4363 GNDA.n4362 3.4105
R13345 GNDA.n4361 GNDA.n4360 3.4105
R13346 GNDA.n4359 GNDA.n4358 3.4105
R13347 GNDA.n4357 GNDA.n4349 3.4105
R13348 GNDA.n4353 GNDA.n4352 3.4105
R13349 GNDA.n4351 GNDA.n4302 3.4105
R13350 GNDA.n4161 GNDA.n4160 3.4105
R13351 GNDA.n4297 GNDA.n4296 3.4105
R13352 GNDA.n4295 GNDA.n4294 3.4105
R13353 GNDA.n4293 GNDA.n4292 3.4105
R13354 GNDA.n4291 GNDA.n4163 3.4105
R13355 GNDA.n4287 GNDA.n4286 3.4105
R13356 GNDA.n4285 GNDA.n4284 3.4105
R13357 GNDA.n4283 GNDA.n4282 3.4105
R13358 GNDA.n4281 GNDA.n4165 3.4105
R13359 GNDA.n4277 GNDA.n4276 3.4105
R13360 GNDA.n4275 GNDA.n4274 3.4105
R13361 GNDA.n4273 GNDA.n4272 3.4105
R13362 GNDA.n4271 GNDA.n4167 3.4105
R13363 GNDA.n4267 GNDA.n4266 3.4105
R13364 GNDA.n4265 GNDA.n4264 3.4105
R13365 GNDA.n4263 GNDA.n4262 3.4105
R13366 GNDA.n4261 GNDA.n4169 3.4105
R13367 GNDA.n4257 GNDA.n4256 3.4105
R13368 GNDA.n4255 GNDA.n4254 3.4105
R13369 GNDA.n4253 GNDA.n4252 3.4105
R13370 GNDA.n4251 GNDA.n4171 3.4105
R13371 GNDA.n4247 GNDA.n4246 3.4105
R13372 GNDA.n4245 GNDA.n4244 3.4105
R13373 GNDA.n4243 GNDA.n4242 3.4105
R13374 GNDA.n4241 GNDA.n4173 3.4105
R13375 GNDA.n4237 GNDA.n4236 3.4105
R13376 GNDA.n4235 GNDA.n4234 3.4105
R13377 GNDA.n4233 GNDA.n4232 3.4105
R13378 GNDA.n4231 GNDA.n4175 3.4105
R13379 GNDA.n4227 GNDA.n4226 3.4105
R13380 GNDA.n4225 GNDA.n4224 3.4105
R13381 GNDA.n4223 GNDA.n4222 3.4105
R13382 GNDA.n4221 GNDA.n4177 3.4105
R13383 GNDA.n4217 GNDA.n4216 3.4105
R13384 GNDA.n4215 GNDA.n4214 3.4105
R13385 GNDA.n4213 GNDA.n4212 3.4105
R13386 GNDA.n4211 GNDA.n4179 3.4105
R13387 GNDA.n4207 GNDA.n4206 3.4105
R13388 GNDA.n4205 GNDA.n4204 3.4105
R13389 GNDA.n4203 GNDA.n4202 3.4105
R13390 GNDA.n4201 GNDA.n4181 3.4105
R13391 GNDA.n4197 GNDA.n4196 3.4105
R13392 GNDA.n4195 GNDA.n4194 3.4105
R13393 GNDA.n4193 GNDA.n4192 3.4105
R13394 GNDA.n4191 GNDA.n4183 3.4105
R13395 GNDA.n4187 GNDA.n4186 3.4105
R13396 GNDA.n4185 GNDA.n4136 3.4105
R13397 GNDA.n3485 GNDA.n3484 3.4105
R13398 GNDA.n3799 GNDA.n3798 3.4105
R13399 GNDA.n3797 GNDA.n3796 3.4105
R13400 GNDA.n3795 GNDA.n3794 3.4105
R13401 GNDA.n3793 GNDA.n3487 3.4105
R13402 GNDA.n3789 GNDA.n3788 3.4105
R13403 GNDA.n3787 GNDA.n3786 3.4105
R13404 GNDA.n3785 GNDA.n3784 3.4105
R13405 GNDA.n3783 GNDA.n3489 3.4105
R13406 GNDA.n3779 GNDA.n3778 3.4105
R13407 GNDA.n3777 GNDA.n3776 3.4105
R13408 GNDA.n3775 GNDA.n3774 3.4105
R13409 GNDA.n3773 GNDA.n3491 3.4105
R13410 GNDA.n3769 GNDA.n3768 3.4105
R13411 GNDA.n3767 GNDA.n3766 3.4105
R13412 GNDA.n3765 GNDA.n3764 3.4105
R13413 GNDA.n3763 GNDA.n3493 3.4105
R13414 GNDA.n3759 GNDA.n3758 3.4105
R13415 GNDA.n3757 GNDA.n3756 3.4105
R13416 GNDA.n3755 GNDA.n3754 3.4105
R13417 GNDA.n3753 GNDA.n3495 3.4105
R13418 GNDA.n3749 GNDA.n3748 3.4105
R13419 GNDA.n3747 GNDA.n3746 3.4105
R13420 GNDA.n3745 GNDA.n3744 3.4105
R13421 GNDA.n3743 GNDA.n3497 3.4105
R13422 GNDA.n3739 GNDA.n3738 3.4105
R13423 GNDA.n3737 GNDA.n3736 3.4105
R13424 GNDA.n3735 GNDA.n3734 3.4105
R13425 GNDA.n3733 GNDA.n3499 3.4105
R13426 GNDA.n3729 GNDA.n3728 3.4105
R13427 GNDA.n3727 GNDA.n3726 3.4105
R13428 GNDA.n3725 GNDA.n3724 3.4105
R13429 GNDA.n3723 GNDA.n3501 3.4105
R13430 GNDA.n3719 GNDA.n3718 3.4105
R13431 GNDA.n3717 GNDA.n3716 3.4105
R13432 GNDA.n3715 GNDA.n3714 3.4105
R13433 GNDA.n3713 GNDA.n3503 3.4105
R13434 GNDA.n3709 GNDA.n3708 3.4105
R13435 GNDA.n3707 GNDA.n3706 3.4105
R13436 GNDA.n3705 GNDA.n3704 3.4105
R13437 GNDA.n3703 GNDA.n3505 3.4105
R13438 GNDA.n3699 GNDA.n3698 3.4105
R13439 GNDA.n3697 GNDA.n3696 3.4105
R13440 GNDA.n3695 GNDA.n3694 3.4105
R13441 GNDA.n3693 GNDA.n3507 3.4105
R13442 GNDA.n3689 GNDA.n3688 3.4105
R13443 GNDA.n3687 GNDA.n3460 3.4105
R13444 GNDA.n3995 GNDA.n3994 3.4105
R13445 GNDA.n4131 GNDA.n4130 3.4105
R13446 GNDA.n4129 GNDA.n4128 3.4105
R13447 GNDA.n4127 GNDA.n4126 3.4105
R13448 GNDA.n4125 GNDA.n3997 3.4105
R13449 GNDA.n4121 GNDA.n4120 3.4105
R13450 GNDA.n4119 GNDA.n4118 3.4105
R13451 GNDA.n4117 GNDA.n4116 3.4105
R13452 GNDA.n4115 GNDA.n3999 3.4105
R13453 GNDA.n4111 GNDA.n4110 3.4105
R13454 GNDA.n4109 GNDA.n4108 3.4105
R13455 GNDA.n4107 GNDA.n4106 3.4105
R13456 GNDA.n4105 GNDA.n4001 3.4105
R13457 GNDA.n4101 GNDA.n4100 3.4105
R13458 GNDA.n4099 GNDA.n4098 3.4105
R13459 GNDA.n4097 GNDA.n4096 3.4105
R13460 GNDA.n4095 GNDA.n4003 3.4105
R13461 GNDA.n4091 GNDA.n4090 3.4105
R13462 GNDA.n4089 GNDA.n4088 3.4105
R13463 GNDA.n4087 GNDA.n4086 3.4105
R13464 GNDA.n4085 GNDA.n4005 3.4105
R13465 GNDA.n4081 GNDA.n4080 3.4105
R13466 GNDA.n4079 GNDA.n4078 3.4105
R13467 GNDA.n4077 GNDA.n4076 3.4105
R13468 GNDA.n4075 GNDA.n4007 3.4105
R13469 GNDA.n4071 GNDA.n4070 3.4105
R13470 GNDA.n4069 GNDA.n4068 3.4105
R13471 GNDA.n4067 GNDA.n4066 3.4105
R13472 GNDA.n4065 GNDA.n4009 3.4105
R13473 GNDA.n4061 GNDA.n4060 3.4105
R13474 GNDA.n4059 GNDA.n4058 3.4105
R13475 GNDA.n4057 GNDA.n4056 3.4105
R13476 GNDA.n4055 GNDA.n4011 3.4105
R13477 GNDA.n4051 GNDA.n4050 3.4105
R13478 GNDA.n4049 GNDA.n4048 3.4105
R13479 GNDA.n4047 GNDA.n4046 3.4105
R13480 GNDA.n4045 GNDA.n4013 3.4105
R13481 GNDA.n4041 GNDA.n4040 3.4105
R13482 GNDA.n4039 GNDA.n4038 3.4105
R13483 GNDA.n4037 GNDA.n4036 3.4105
R13484 GNDA.n4035 GNDA.n4015 3.4105
R13485 GNDA.n4031 GNDA.n4030 3.4105
R13486 GNDA.n4029 GNDA.n4028 3.4105
R13487 GNDA.n4027 GNDA.n4026 3.4105
R13488 GNDA.n4025 GNDA.n4017 3.4105
R13489 GNDA.n4021 GNDA.n4020 3.4105
R13490 GNDA.n4019 GNDA.n3970 3.4105
R13491 GNDA.n3829 GNDA.n3828 3.4105
R13492 GNDA.n3965 GNDA.n3964 3.4105
R13493 GNDA.n3963 GNDA.n3962 3.4105
R13494 GNDA.n3961 GNDA.n3960 3.4105
R13495 GNDA.n3959 GNDA.n3831 3.4105
R13496 GNDA.n3955 GNDA.n3954 3.4105
R13497 GNDA.n3953 GNDA.n3952 3.4105
R13498 GNDA.n3951 GNDA.n3950 3.4105
R13499 GNDA.n3949 GNDA.n3833 3.4105
R13500 GNDA.n3945 GNDA.n3944 3.4105
R13501 GNDA.n3943 GNDA.n3942 3.4105
R13502 GNDA.n3941 GNDA.n3940 3.4105
R13503 GNDA.n3939 GNDA.n3835 3.4105
R13504 GNDA.n3935 GNDA.n3934 3.4105
R13505 GNDA.n3933 GNDA.n3932 3.4105
R13506 GNDA.n3931 GNDA.n3930 3.4105
R13507 GNDA.n3929 GNDA.n3837 3.4105
R13508 GNDA.n3925 GNDA.n3924 3.4105
R13509 GNDA.n3923 GNDA.n3922 3.4105
R13510 GNDA.n3921 GNDA.n3920 3.4105
R13511 GNDA.n3919 GNDA.n3839 3.4105
R13512 GNDA.n3915 GNDA.n3914 3.4105
R13513 GNDA.n3913 GNDA.n3912 3.4105
R13514 GNDA.n3911 GNDA.n3910 3.4105
R13515 GNDA.n3909 GNDA.n3841 3.4105
R13516 GNDA.n3905 GNDA.n3904 3.4105
R13517 GNDA.n3903 GNDA.n3902 3.4105
R13518 GNDA.n3901 GNDA.n3900 3.4105
R13519 GNDA.n3899 GNDA.n3843 3.4105
R13520 GNDA.n3895 GNDA.n3894 3.4105
R13521 GNDA.n3893 GNDA.n3892 3.4105
R13522 GNDA.n3891 GNDA.n3890 3.4105
R13523 GNDA.n3889 GNDA.n3845 3.4105
R13524 GNDA.n3885 GNDA.n3884 3.4105
R13525 GNDA.n3883 GNDA.n3882 3.4105
R13526 GNDA.n3881 GNDA.n3880 3.4105
R13527 GNDA.n3879 GNDA.n3847 3.4105
R13528 GNDA.n3875 GNDA.n3874 3.4105
R13529 GNDA.n3873 GNDA.n3872 3.4105
R13530 GNDA.n3871 GNDA.n3870 3.4105
R13531 GNDA.n3869 GNDA.n3849 3.4105
R13532 GNDA.n3865 GNDA.n3864 3.4105
R13533 GNDA.n3863 GNDA.n3862 3.4105
R13534 GNDA.n3861 GNDA.n3860 3.4105
R13535 GNDA.n3859 GNDA.n3851 3.4105
R13536 GNDA.n3855 GNDA.n3854 3.4105
R13537 GNDA.n3853 GNDA.n3804 3.4105
R13538 GNDA.n3604 GNDA.n3557 3.4105
R13539 GNDA.n3606 GNDA.n3556 3.4105
R13540 GNDA.n3607 GNDA.n3555 3.4105
R13541 GNDA.n3609 GNDA.n3554 3.4105
R13542 GNDA.n3610 GNDA.n3553 3.4105
R13543 GNDA.n3612 GNDA.n3552 3.4105
R13544 GNDA.n3613 GNDA.n3551 3.4105
R13545 GNDA.n3615 GNDA.n3550 3.4105
R13546 GNDA.n3616 GNDA.n3549 3.4105
R13547 GNDA.n3618 GNDA.n3548 3.4105
R13548 GNDA.n3619 GNDA.n3547 3.4105
R13549 GNDA.n3621 GNDA.n3546 3.4105
R13550 GNDA.n3622 GNDA.n3545 3.4105
R13551 GNDA.n3624 GNDA.n3544 3.4105
R13552 GNDA.n3625 GNDA.n3543 3.4105
R13553 GNDA.n3627 GNDA.n3542 3.4105
R13554 GNDA.n3628 GNDA.n3541 3.4105
R13555 GNDA.n3630 GNDA.n3540 3.4105
R13556 GNDA.n3631 GNDA.n3539 3.4105
R13557 GNDA.n3633 GNDA.n3538 3.4105
R13558 GNDA.n3634 GNDA.n3537 3.4105
R13559 GNDA.n3636 GNDA.n3536 3.4105
R13560 GNDA.n3637 GNDA.n3535 3.4105
R13561 GNDA.n3639 GNDA.n3534 3.4105
R13562 GNDA.n3640 GNDA.n3533 3.4105
R13563 GNDA.n3642 GNDA.n3532 3.4105
R13564 GNDA.n3643 GNDA.n3531 3.4105
R13565 GNDA.n3645 GNDA.n3530 3.4105
R13566 GNDA.n3646 GNDA.n3529 3.4105
R13567 GNDA.n3648 GNDA.n3528 3.4105
R13568 GNDA.n3649 GNDA.n3527 3.4105
R13569 GNDA.n3651 GNDA.n3526 3.4105
R13570 GNDA.n3652 GNDA.n3525 3.4105
R13571 GNDA.n3654 GNDA.n3524 3.4105
R13572 GNDA.n3655 GNDA.n3523 3.4105
R13573 GNDA.n3657 GNDA.n3522 3.4105
R13574 GNDA.n3658 GNDA.n3521 3.4105
R13575 GNDA.n3660 GNDA.n3520 3.4105
R13576 GNDA.n3661 GNDA.n3519 3.4105
R13577 GNDA.n3663 GNDA.n3518 3.4105
R13578 GNDA.n3664 GNDA.n3517 3.4105
R13579 GNDA.n3666 GNDA.n3516 3.4105
R13580 GNDA.n3667 GNDA.n3515 3.4105
R13581 GNDA.n3669 GNDA.n3514 3.4105
R13582 GNDA.n3670 GNDA.n3513 3.4105
R13583 GNDA.n3672 GNDA.n3512 3.4105
R13584 GNDA.n3674 GNDA.n3673 3.4105
R13585 GNDA.n498 GNDA.n451 3.4105
R13586 GNDA.n500 GNDA.n450 3.4105
R13587 GNDA.n501 GNDA.n449 3.4105
R13588 GNDA.n503 GNDA.n448 3.4105
R13589 GNDA.n504 GNDA.n447 3.4105
R13590 GNDA.n506 GNDA.n446 3.4105
R13591 GNDA.n507 GNDA.n445 3.4105
R13592 GNDA.n509 GNDA.n444 3.4105
R13593 GNDA.n510 GNDA.n443 3.4105
R13594 GNDA.n512 GNDA.n442 3.4105
R13595 GNDA.n513 GNDA.n441 3.4105
R13596 GNDA.n515 GNDA.n440 3.4105
R13597 GNDA.n516 GNDA.n439 3.4105
R13598 GNDA.n518 GNDA.n438 3.4105
R13599 GNDA.n519 GNDA.n437 3.4105
R13600 GNDA.n521 GNDA.n436 3.4105
R13601 GNDA.n522 GNDA.n435 3.4105
R13602 GNDA.n524 GNDA.n434 3.4105
R13603 GNDA.n525 GNDA.n433 3.4105
R13604 GNDA.n527 GNDA.n432 3.4105
R13605 GNDA.n528 GNDA.n431 3.4105
R13606 GNDA.n530 GNDA.n430 3.4105
R13607 GNDA.n531 GNDA.n429 3.4105
R13608 GNDA.n533 GNDA.n428 3.4105
R13609 GNDA.n534 GNDA.n427 3.4105
R13610 GNDA.n536 GNDA.n426 3.4105
R13611 GNDA.n537 GNDA.n425 3.4105
R13612 GNDA.n539 GNDA.n424 3.4105
R13613 GNDA.n540 GNDA.n423 3.4105
R13614 GNDA.n542 GNDA.n422 3.4105
R13615 GNDA.n543 GNDA.n421 3.4105
R13616 GNDA.n545 GNDA.n420 3.4105
R13617 GNDA.n546 GNDA.n419 3.4105
R13618 GNDA.n548 GNDA.n418 3.4105
R13619 GNDA.n549 GNDA.n417 3.4105
R13620 GNDA.n551 GNDA.n416 3.4105
R13621 GNDA.n552 GNDA.n415 3.4105
R13622 GNDA.n554 GNDA.n414 3.4105
R13623 GNDA.n555 GNDA.n413 3.4105
R13624 GNDA.n557 GNDA.n412 3.4105
R13625 GNDA.n558 GNDA.n411 3.4105
R13626 GNDA.n560 GNDA.n410 3.4105
R13627 GNDA.n561 GNDA.n409 3.4105
R13628 GNDA.n563 GNDA.n408 3.4105
R13629 GNDA.n564 GNDA.n407 3.4105
R13630 GNDA.n566 GNDA.n406 3.4105
R13631 GNDA.n568 GNDA.n567 3.4105
R13632 GNDA.n379 GNDA.n378 3.4105
R13633 GNDA.n5131 GNDA.n5130 3.4105
R13634 GNDA.n5129 GNDA.n5128 3.4105
R13635 GNDA.n5127 GNDA.n5126 3.4105
R13636 GNDA.n5125 GNDA.n381 3.4105
R13637 GNDA.n5121 GNDA.n5120 3.4105
R13638 GNDA.n5119 GNDA.n5118 3.4105
R13639 GNDA.n5117 GNDA.n5116 3.4105
R13640 GNDA.n5115 GNDA.n383 3.4105
R13641 GNDA.n5111 GNDA.n5110 3.4105
R13642 GNDA.n5109 GNDA.n5108 3.4105
R13643 GNDA.n5107 GNDA.n5106 3.4105
R13644 GNDA.n5105 GNDA.n385 3.4105
R13645 GNDA.n5101 GNDA.n5100 3.4105
R13646 GNDA.n5099 GNDA.n5098 3.4105
R13647 GNDA.n5097 GNDA.n5096 3.4105
R13648 GNDA.n5095 GNDA.n387 3.4105
R13649 GNDA.n5091 GNDA.n5090 3.4105
R13650 GNDA.n5089 GNDA.n5088 3.4105
R13651 GNDA.n5087 GNDA.n5086 3.4105
R13652 GNDA.n5085 GNDA.n389 3.4105
R13653 GNDA.n5081 GNDA.n5080 3.4105
R13654 GNDA.n5079 GNDA.n5078 3.4105
R13655 GNDA.n5077 GNDA.n5076 3.4105
R13656 GNDA.n5075 GNDA.n391 3.4105
R13657 GNDA.n5071 GNDA.n5070 3.4105
R13658 GNDA.n5069 GNDA.n5068 3.4105
R13659 GNDA.n5067 GNDA.n5066 3.4105
R13660 GNDA.n5065 GNDA.n393 3.4105
R13661 GNDA.n5061 GNDA.n5060 3.4105
R13662 GNDA.n5059 GNDA.n5058 3.4105
R13663 GNDA.n5057 GNDA.n5056 3.4105
R13664 GNDA.n5055 GNDA.n395 3.4105
R13665 GNDA.n5051 GNDA.n5050 3.4105
R13666 GNDA.n5049 GNDA.n5048 3.4105
R13667 GNDA.n5047 GNDA.n5046 3.4105
R13668 GNDA.n5045 GNDA.n397 3.4105
R13669 GNDA.n5041 GNDA.n5040 3.4105
R13670 GNDA.n5039 GNDA.n5038 3.4105
R13671 GNDA.n5037 GNDA.n5036 3.4105
R13672 GNDA.n5035 GNDA.n399 3.4105
R13673 GNDA.n5031 GNDA.n5030 3.4105
R13674 GNDA.n5029 GNDA.n5028 3.4105
R13675 GNDA.n5027 GNDA.n5026 3.4105
R13676 GNDA.n5025 GNDA.n401 3.4105
R13677 GNDA.n5021 GNDA.n5020 3.4105
R13678 GNDA.n5019 GNDA.n353 3.4105
R13679 GNDA.n3301 GNDA.n3254 3.4105
R13680 GNDA.n3303 GNDA.n3253 3.4105
R13681 GNDA.n3304 GNDA.n3252 3.4105
R13682 GNDA.n3306 GNDA.n3251 3.4105
R13683 GNDA.n3307 GNDA.n3250 3.4105
R13684 GNDA.n3309 GNDA.n3249 3.4105
R13685 GNDA.n3310 GNDA.n3248 3.4105
R13686 GNDA.n3312 GNDA.n3247 3.4105
R13687 GNDA.n3313 GNDA.n3246 3.4105
R13688 GNDA.n3315 GNDA.n3245 3.4105
R13689 GNDA.n3316 GNDA.n3244 3.4105
R13690 GNDA.n3318 GNDA.n3243 3.4105
R13691 GNDA.n3319 GNDA.n3242 3.4105
R13692 GNDA.n3321 GNDA.n3241 3.4105
R13693 GNDA.n3322 GNDA.n3240 3.4105
R13694 GNDA.n3324 GNDA.n3239 3.4105
R13695 GNDA.n3325 GNDA.n3238 3.4105
R13696 GNDA.n3327 GNDA.n3237 3.4105
R13697 GNDA.n3328 GNDA.n3236 3.4105
R13698 GNDA.n3330 GNDA.n3235 3.4105
R13699 GNDA.n3331 GNDA.n3234 3.4105
R13700 GNDA.n3333 GNDA.n3233 3.4105
R13701 GNDA.n3334 GNDA.n3232 3.4105
R13702 GNDA.n3336 GNDA.n3231 3.4105
R13703 GNDA.n3337 GNDA.n3230 3.4105
R13704 GNDA.n3339 GNDA.n3229 3.4105
R13705 GNDA.n3340 GNDA.n3228 3.4105
R13706 GNDA.n3342 GNDA.n3227 3.4105
R13707 GNDA.n3343 GNDA.n3226 3.4105
R13708 GNDA.n3345 GNDA.n3225 3.4105
R13709 GNDA.n3346 GNDA.n3224 3.4105
R13710 GNDA.n3348 GNDA.n3223 3.4105
R13711 GNDA.n3349 GNDA.n3222 3.4105
R13712 GNDA.n3351 GNDA.n3221 3.4105
R13713 GNDA.n3352 GNDA.n3220 3.4105
R13714 GNDA.n3354 GNDA.n3219 3.4105
R13715 GNDA.n3355 GNDA.n3218 3.4105
R13716 GNDA.n3357 GNDA.n3217 3.4105
R13717 GNDA.n3358 GNDA.n3216 3.4105
R13718 GNDA.n3360 GNDA.n3215 3.4105
R13719 GNDA.n3361 GNDA.n3214 3.4105
R13720 GNDA.n3363 GNDA.n3213 3.4105
R13721 GNDA.n3364 GNDA.n3212 3.4105
R13722 GNDA.n3366 GNDA.n3211 3.4105
R13723 GNDA.n3367 GNDA.n3210 3.4105
R13724 GNDA.n3369 GNDA.n3209 3.4105
R13725 GNDA.n3371 GNDA.n3370 3.4105
R13726 GNDA.n3062 GNDA.n3061 3.4105
R13727 GNDA.n3193 GNDA.n3192 3.4105
R13728 GNDA.n3191 GNDA.n3190 3.4105
R13729 GNDA.n3189 GNDA.n3188 3.4105
R13730 GNDA.n3187 GNDA.n3064 3.4105
R13731 GNDA.n3183 GNDA.n3182 3.4105
R13732 GNDA.n3181 GNDA.n3180 3.4105
R13733 GNDA.n3179 GNDA.n3178 3.4105
R13734 GNDA.n3177 GNDA.n3066 3.4105
R13735 GNDA.n3173 GNDA.n3172 3.4105
R13736 GNDA.n3171 GNDA.n3170 3.4105
R13737 GNDA.n3169 GNDA.n3168 3.4105
R13738 GNDA.n3167 GNDA.n3068 3.4105
R13739 GNDA.n3163 GNDA.n3162 3.4105
R13740 GNDA.n3161 GNDA.n3160 3.4105
R13741 GNDA.n3159 GNDA.n3158 3.4105
R13742 GNDA.n3157 GNDA.n3070 3.4105
R13743 GNDA.n3153 GNDA.n3152 3.4105
R13744 GNDA.n3151 GNDA.n3150 3.4105
R13745 GNDA.n3149 GNDA.n3148 3.4105
R13746 GNDA.n3147 GNDA.n3072 3.4105
R13747 GNDA.n3143 GNDA.n3142 3.4105
R13748 GNDA.n3141 GNDA.n3140 3.4105
R13749 GNDA.n3139 GNDA.n3138 3.4105
R13750 GNDA.n3137 GNDA.n3074 3.4105
R13751 GNDA.n3133 GNDA.n3132 3.4105
R13752 GNDA.n3131 GNDA.n3130 3.4105
R13753 GNDA.n3129 GNDA.n3128 3.4105
R13754 GNDA.n3127 GNDA.n3076 3.4105
R13755 GNDA.n3123 GNDA.n3122 3.4105
R13756 GNDA.n3121 GNDA.n3120 3.4105
R13757 GNDA.n3119 GNDA.n3118 3.4105
R13758 GNDA.n3117 GNDA.n3078 3.4105
R13759 GNDA.n3113 GNDA.n3112 3.4105
R13760 GNDA.n3111 GNDA.n3110 3.4105
R13761 GNDA.n3109 GNDA.n3108 3.4105
R13762 GNDA.n3107 GNDA.n3080 3.4105
R13763 GNDA.n3103 GNDA.n3102 3.4105
R13764 GNDA.n3101 GNDA.n3100 3.4105
R13765 GNDA.n3099 GNDA.n3098 3.4105
R13766 GNDA.n3097 GNDA.n3082 3.4105
R13767 GNDA.n3093 GNDA.n3092 3.4105
R13768 GNDA.n3091 GNDA.n3090 3.4105
R13769 GNDA.n3089 GNDA.n3088 3.4105
R13770 GNDA.n3087 GNDA.n3084 3.4105
R13771 GNDA.n598 GNDA.n597 3.4105
R13772 GNDA.n3199 GNDA.n3198 3.4105
R13773 GNDA.n2889 GNDA.n2888 3.4105
R13774 GNDA.n3033 GNDA.n3032 3.4105
R13775 GNDA.n3031 GNDA.n3030 3.4105
R13776 GNDA.n3029 GNDA.n3028 3.4105
R13777 GNDA.n3027 GNDA.n2891 3.4105
R13778 GNDA.n3023 GNDA.n3022 3.4105
R13779 GNDA.n3021 GNDA.n3020 3.4105
R13780 GNDA.n3019 GNDA.n3018 3.4105
R13781 GNDA.n3017 GNDA.n2893 3.4105
R13782 GNDA.n3013 GNDA.n3012 3.4105
R13783 GNDA.n3011 GNDA.n3010 3.4105
R13784 GNDA.n3009 GNDA.n3008 3.4105
R13785 GNDA.n3007 GNDA.n2895 3.4105
R13786 GNDA.n3003 GNDA.n3002 3.4105
R13787 GNDA.n3001 GNDA.n3000 3.4105
R13788 GNDA.n2999 GNDA.n2998 3.4105
R13789 GNDA.n2997 GNDA.n2897 3.4105
R13790 GNDA.n2993 GNDA.n2992 3.4105
R13791 GNDA.n2991 GNDA.n2990 3.4105
R13792 GNDA.n2989 GNDA.n2988 3.4105
R13793 GNDA.n2987 GNDA.n2899 3.4105
R13794 GNDA.n2983 GNDA.n2982 3.4105
R13795 GNDA.n2981 GNDA.n2980 3.4105
R13796 GNDA.n2979 GNDA.n2978 3.4105
R13797 GNDA.n2977 GNDA.n2901 3.4105
R13798 GNDA.n2973 GNDA.n2972 3.4105
R13799 GNDA.n2971 GNDA.n2970 3.4105
R13800 GNDA.n2969 GNDA.n2968 3.4105
R13801 GNDA.n2967 GNDA.n2903 3.4105
R13802 GNDA.n2963 GNDA.n2962 3.4105
R13803 GNDA.n2961 GNDA.n2960 3.4105
R13804 GNDA.n2959 GNDA.n2958 3.4105
R13805 GNDA.n2957 GNDA.n2905 3.4105
R13806 GNDA.n2953 GNDA.n2952 3.4105
R13807 GNDA.n2951 GNDA.n2950 3.4105
R13808 GNDA.n2949 GNDA.n2948 3.4105
R13809 GNDA.n2947 GNDA.n2907 3.4105
R13810 GNDA.n2943 GNDA.n2942 3.4105
R13811 GNDA.n2941 GNDA.n2940 3.4105
R13812 GNDA.n2939 GNDA.n2938 3.4105
R13813 GNDA.n2937 GNDA.n2909 3.4105
R13814 GNDA.n2933 GNDA.n2932 3.4105
R13815 GNDA.n2931 GNDA.n2930 3.4105
R13816 GNDA.n2929 GNDA.n2928 3.4105
R13817 GNDA.n2927 GNDA.n2911 3.4105
R13818 GNDA.n2923 GNDA.n2922 3.4105
R13819 GNDA.n2921 GNDA.n2864 3.4105
R13820 GNDA.n691 GNDA.n690 3.4105
R13821 GNDA.n2397 GNDA.n2396 3.4105
R13822 GNDA.n2395 GNDA.n2394 3.4105
R13823 GNDA.n2393 GNDA.n2392 3.4105
R13824 GNDA.n2391 GNDA.n693 3.4105
R13825 GNDA.n2387 GNDA.n2386 3.4105
R13826 GNDA.n2385 GNDA.n2384 3.4105
R13827 GNDA.n2383 GNDA.n2382 3.4105
R13828 GNDA.n2381 GNDA.n695 3.4105
R13829 GNDA.n2377 GNDA.n2376 3.4105
R13830 GNDA.n2375 GNDA.n2374 3.4105
R13831 GNDA.n2373 GNDA.n2372 3.4105
R13832 GNDA.n2371 GNDA.n697 3.4105
R13833 GNDA.n2367 GNDA.n2366 3.4105
R13834 GNDA.n2365 GNDA.n2364 3.4105
R13835 GNDA.n2363 GNDA.n2362 3.4105
R13836 GNDA.n2361 GNDA.n699 3.4105
R13837 GNDA.n2357 GNDA.n2356 3.4105
R13838 GNDA.n2355 GNDA.n2354 3.4105
R13839 GNDA.n2353 GNDA.n2352 3.4105
R13840 GNDA.n2351 GNDA.n701 3.4105
R13841 GNDA.n2347 GNDA.n2346 3.4105
R13842 GNDA.n2345 GNDA.n2344 3.4105
R13843 GNDA.n2343 GNDA.n2342 3.4105
R13844 GNDA.n2341 GNDA.n703 3.4105
R13845 GNDA.n2337 GNDA.n2336 3.4105
R13846 GNDA.n2335 GNDA.n2334 3.4105
R13847 GNDA.n2333 GNDA.n2332 3.4105
R13848 GNDA.n2331 GNDA.n705 3.4105
R13849 GNDA.n2327 GNDA.n2326 3.4105
R13850 GNDA.n2325 GNDA.n2324 3.4105
R13851 GNDA.n2323 GNDA.n2322 3.4105
R13852 GNDA.n2321 GNDA.n707 3.4105
R13853 GNDA.n2317 GNDA.n2316 3.4105
R13854 GNDA.n2315 GNDA.n2314 3.4105
R13855 GNDA.n2313 GNDA.n2312 3.4105
R13856 GNDA.n2311 GNDA.n709 3.4105
R13857 GNDA.n2307 GNDA.n2306 3.4105
R13858 GNDA.n2305 GNDA.n2304 3.4105
R13859 GNDA.n2303 GNDA.n2302 3.4105
R13860 GNDA.n2301 GNDA.n711 3.4105
R13861 GNDA.n2297 GNDA.n2296 3.4105
R13862 GNDA.n2295 GNDA.n2294 3.4105
R13863 GNDA.n2293 GNDA.n2292 3.4105
R13864 GNDA.n2291 GNDA.n713 3.4105
R13865 GNDA.n2287 GNDA.n2286 3.4105
R13866 GNDA.n2285 GNDA.n666 3.4105
R13867 GNDA.n625 GNDA.n624 3.4105
R13868 GNDA.n2859 GNDA.n2858 3.4105
R13869 GNDA.n2857 GNDA.n2856 3.4105
R13870 GNDA.n2855 GNDA.n2854 3.4105
R13871 GNDA.n2853 GNDA.n627 3.4105
R13872 GNDA.n2849 GNDA.n2848 3.4105
R13873 GNDA.n2847 GNDA.n2846 3.4105
R13874 GNDA.n2845 GNDA.n2844 3.4105
R13875 GNDA.n2843 GNDA.n629 3.4105
R13876 GNDA.n2839 GNDA.n2838 3.4105
R13877 GNDA.n2837 GNDA.n2836 3.4105
R13878 GNDA.n2835 GNDA.n2834 3.4105
R13879 GNDA.n2833 GNDA.n631 3.4105
R13880 GNDA.n2829 GNDA.n2828 3.4105
R13881 GNDA.n2827 GNDA.n2826 3.4105
R13882 GNDA.n2825 GNDA.n2824 3.4105
R13883 GNDA.n2823 GNDA.n633 3.4105
R13884 GNDA.n2819 GNDA.n2818 3.4105
R13885 GNDA.n2817 GNDA.n2816 3.4105
R13886 GNDA.n2815 GNDA.n2814 3.4105
R13887 GNDA.n2813 GNDA.n635 3.4105
R13888 GNDA.n2809 GNDA.n2808 3.4105
R13889 GNDA.n2807 GNDA.n2806 3.4105
R13890 GNDA.n2805 GNDA.n2804 3.4105
R13891 GNDA.n2803 GNDA.n637 3.4105
R13892 GNDA.n2799 GNDA.n2798 3.4105
R13893 GNDA.n2797 GNDA.n2796 3.4105
R13894 GNDA.n2795 GNDA.n2794 3.4105
R13895 GNDA.n2793 GNDA.n639 3.4105
R13896 GNDA.n2789 GNDA.n2788 3.4105
R13897 GNDA.n2787 GNDA.n2786 3.4105
R13898 GNDA.n2785 GNDA.n2784 3.4105
R13899 GNDA.n2783 GNDA.n641 3.4105
R13900 GNDA.n2779 GNDA.n2778 3.4105
R13901 GNDA.n2777 GNDA.n2776 3.4105
R13902 GNDA.n2775 GNDA.n2774 3.4105
R13903 GNDA.n2773 GNDA.n643 3.4105
R13904 GNDA.n2769 GNDA.n2768 3.4105
R13905 GNDA.n2767 GNDA.n2766 3.4105
R13906 GNDA.n2765 GNDA.n2764 3.4105
R13907 GNDA.n2763 GNDA.n645 3.4105
R13908 GNDA.n2759 GNDA.n2758 3.4105
R13909 GNDA.n2757 GNDA.n2756 3.4105
R13910 GNDA.n2755 GNDA.n2754 3.4105
R13911 GNDA.n2753 GNDA.n647 3.4105
R13912 GNDA.n2749 GNDA.n2748 3.4105
R13913 GNDA.n2747 GNDA.n600 3.4105
R13914 GNDA.n2664 GNDA.n2617 3.4105
R13915 GNDA.n2666 GNDA.n2616 3.4105
R13916 GNDA.n2667 GNDA.n2615 3.4105
R13917 GNDA.n2669 GNDA.n2614 3.4105
R13918 GNDA.n2670 GNDA.n2613 3.4105
R13919 GNDA.n2672 GNDA.n2612 3.4105
R13920 GNDA.n2673 GNDA.n2611 3.4105
R13921 GNDA.n2675 GNDA.n2610 3.4105
R13922 GNDA.n2676 GNDA.n2609 3.4105
R13923 GNDA.n2678 GNDA.n2608 3.4105
R13924 GNDA.n2679 GNDA.n2607 3.4105
R13925 GNDA.n2681 GNDA.n2606 3.4105
R13926 GNDA.n2682 GNDA.n2605 3.4105
R13927 GNDA.n2684 GNDA.n2604 3.4105
R13928 GNDA.n2685 GNDA.n2603 3.4105
R13929 GNDA.n2687 GNDA.n2602 3.4105
R13930 GNDA.n2688 GNDA.n2601 3.4105
R13931 GNDA.n2690 GNDA.n2600 3.4105
R13932 GNDA.n2691 GNDA.n2599 3.4105
R13933 GNDA.n2693 GNDA.n2598 3.4105
R13934 GNDA.n2694 GNDA.n2597 3.4105
R13935 GNDA.n2696 GNDA.n2596 3.4105
R13936 GNDA.n2697 GNDA.n2595 3.4105
R13937 GNDA.n2699 GNDA.n2594 3.4105
R13938 GNDA.n2700 GNDA.n2593 3.4105
R13939 GNDA.n2702 GNDA.n2592 3.4105
R13940 GNDA.n2703 GNDA.n2591 3.4105
R13941 GNDA.n2705 GNDA.n2590 3.4105
R13942 GNDA.n2706 GNDA.n2589 3.4105
R13943 GNDA.n2708 GNDA.n2588 3.4105
R13944 GNDA.n2709 GNDA.n2587 3.4105
R13945 GNDA.n2711 GNDA.n2586 3.4105
R13946 GNDA.n2712 GNDA.n2585 3.4105
R13947 GNDA.n2714 GNDA.n2584 3.4105
R13948 GNDA.n2715 GNDA.n2583 3.4105
R13949 GNDA.n2717 GNDA.n2582 3.4105
R13950 GNDA.n2718 GNDA.n2581 3.4105
R13951 GNDA.n2720 GNDA.n2580 3.4105
R13952 GNDA.n2721 GNDA.n2579 3.4105
R13953 GNDA.n2723 GNDA.n2578 3.4105
R13954 GNDA.n2724 GNDA.n2577 3.4105
R13955 GNDA.n2726 GNDA.n2576 3.4105
R13956 GNDA.n2727 GNDA.n2575 3.4105
R13957 GNDA.n2729 GNDA.n2574 3.4105
R13958 GNDA.n2730 GNDA.n2573 3.4105
R13959 GNDA.n2732 GNDA.n2572 3.4105
R13960 GNDA.n2734 GNDA.n2733 3.4105
R13961 GNDA.n2426 GNDA.n2425 3.4105
R13962 GNDA.n2557 GNDA.n2556 3.4105
R13963 GNDA.n2555 GNDA.n2554 3.4105
R13964 GNDA.n2553 GNDA.n2552 3.4105
R13965 GNDA.n2551 GNDA.n2428 3.4105
R13966 GNDA.n2547 GNDA.n2546 3.4105
R13967 GNDA.n2545 GNDA.n2544 3.4105
R13968 GNDA.n2543 GNDA.n2542 3.4105
R13969 GNDA.n2541 GNDA.n2430 3.4105
R13970 GNDA.n2537 GNDA.n2536 3.4105
R13971 GNDA.n2535 GNDA.n2534 3.4105
R13972 GNDA.n2533 GNDA.n2532 3.4105
R13973 GNDA.n2531 GNDA.n2432 3.4105
R13974 GNDA.n2527 GNDA.n2526 3.4105
R13975 GNDA.n2525 GNDA.n2524 3.4105
R13976 GNDA.n2523 GNDA.n2522 3.4105
R13977 GNDA.n2521 GNDA.n2434 3.4105
R13978 GNDA.n2517 GNDA.n2516 3.4105
R13979 GNDA.n2515 GNDA.n2514 3.4105
R13980 GNDA.n2513 GNDA.n2512 3.4105
R13981 GNDA.n2511 GNDA.n2436 3.4105
R13982 GNDA.n2507 GNDA.n2506 3.4105
R13983 GNDA.n2505 GNDA.n2504 3.4105
R13984 GNDA.n2503 GNDA.n2502 3.4105
R13985 GNDA.n2501 GNDA.n2438 3.4105
R13986 GNDA.n2497 GNDA.n2496 3.4105
R13987 GNDA.n2495 GNDA.n2494 3.4105
R13988 GNDA.n2493 GNDA.n2492 3.4105
R13989 GNDA.n2491 GNDA.n2440 3.4105
R13990 GNDA.n2487 GNDA.n2486 3.4105
R13991 GNDA.n2485 GNDA.n2484 3.4105
R13992 GNDA.n2483 GNDA.n2482 3.4105
R13993 GNDA.n2481 GNDA.n2442 3.4105
R13994 GNDA.n2477 GNDA.n2476 3.4105
R13995 GNDA.n2475 GNDA.n2474 3.4105
R13996 GNDA.n2473 GNDA.n2472 3.4105
R13997 GNDA.n2471 GNDA.n2444 3.4105
R13998 GNDA.n2467 GNDA.n2466 3.4105
R13999 GNDA.n2465 GNDA.n2464 3.4105
R14000 GNDA.n2463 GNDA.n2462 3.4105
R14001 GNDA.n2461 GNDA.n2446 3.4105
R14002 GNDA.n2457 GNDA.n2456 3.4105
R14003 GNDA.n2455 GNDA.n2454 3.4105
R14004 GNDA.n2453 GNDA.n2452 3.4105
R14005 GNDA.n2451 GNDA.n2448 3.4105
R14006 GNDA.n664 GNDA.n663 3.4105
R14007 GNDA.n2563 GNDA.n2562 3.4105
R14008 GNDA.n2204 GNDA.n2157 3.4105
R14009 GNDA.n2206 GNDA.n2156 3.4105
R14010 GNDA.n2207 GNDA.n2155 3.4105
R14011 GNDA.n2209 GNDA.n2154 3.4105
R14012 GNDA.n2210 GNDA.n2153 3.4105
R14013 GNDA.n2212 GNDA.n2152 3.4105
R14014 GNDA.n2213 GNDA.n2151 3.4105
R14015 GNDA.n2215 GNDA.n2150 3.4105
R14016 GNDA.n2216 GNDA.n2149 3.4105
R14017 GNDA.n2218 GNDA.n2148 3.4105
R14018 GNDA.n2219 GNDA.n2147 3.4105
R14019 GNDA.n2221 GNDA.n2146 3.4105
R14020 GNDA.n2222 GNDA.n2145 3.4105
R14021 GNDA.n2224 GNDA.n2144 3.4105
R14022 GNDA.n2225 GNDA.n2143 3.4105
R14023 GNDA.n2227 GNDA.n2142 3.4105
R14024 GNDA.n2228 GNDA.n2141 3.4105
R14025 GNDA.n2230 GNDA.n2140 3.4105
R14026 GNDA.n2231 GNDA.n2139 3.4105
R14027 GNDA.n2233 GNDA.n2138 3.4105
R14028 GNDA.n2234 GNDA.n2137 3.4105
R14029 GNDA.n2236 GNDA.n2136 3.4105
R14030 GNDA.n2237 GNDA.n2135 3.4105
R14031 GNDA.n2239 GNDA.n2134 3.4105
R14032 GNDA.n2240 GNDA.n2133 3.4105
R14033 GNDA.n2242 GNDA.n2132 3.4105
R14034 GNDA.n2243 GNDA.n2131 3.4105
R14035 GNDA.n2245 GNDA.n2130 3.4105
R14036 GNDA.n2246 GNDA.n2129 3.4105
R14037 GNDA.n2248 GNDA.n2128 3.4105
R14038 GNDA.n2249 GNDA.n2127 3.4105
R14039 GNDA.n2251 GNDA.n2126 3.4105
R14040 GNDA.n2252 GNDA.n2125 3.4105
R14041 GNDA.n2254 GNDA.n2124 3.4105
R14042 GNDA.n2255 GNDA.n2123 3.4105
R14043 GNDA.n2257 GNDA.n2122 3.4105
R14044 GNDA.n2258 GNDA.n2121 3.4105
R14045 GNDA.n2260 GNDA.n2120 3.4105
R14046 GNDA.n2261 GNDA.n2119 3.4105
R14047 GNDA.n2263 GNDA.n2118 3.4105
R14048 GNDA.n2264 GNDA.n2117 3.4105
R14049 GNDA.n2266 GNDA.n2116 3.4105
R14050 GNDA.n2267 GNDA.n2115 3.4105
R14051 GNDA.n2269 GNDA.n2114 3.4105
R14052 GNDA.n2270 GNDA.n2113 3.4105
R14053 GNDA.n2272 GNDA.n2112 3.4105
R14054 GNDA.n2274 GNDA.n2273 3.4105
R14055 GNDA.n1963 GNDA.n1962 3.4105
R14056 GNDA.n2094 GNDA.n2093 3.4105
R14057 GNDA.n2092 GNDA.n2091 3.4105
R14058 GNDA.n2090 GNDA.n2089 3.4105
R14059 GNDA.n2088 GNDA.n1965 3.4105
R14060 GNDA.n2084 GNDA.n2083 3.4105
R14061 GNDA.n2082 GNDA.n2081 3.4105
R14062 GNDA.n2080 GNDA.n2079 3.4105
R14063 GNDA.n2078 GNDA.n1967 3.4105
R14064 GNDA.n2074 GNDA.n2073 3.4105
R14065 GNDA.n2072 GNDA.n2071 3.4105
R14066 GNDA.n2070 GNDA.n2069 3.4105
R14067 GNDA.n2068 GNDA.n1969 3.4105
R14068 GNDA.n2064 GNDA.n2063 3.4105
R14069 GNDA.n2062 GNDA.n2061 3.4105
R14070 GNDA.n2060 GNDA.n2059 3.4105
R14071 GNDA.n2058 GNDA.n1971 3.4105
R14072 GNDA.n2054 GNDA.n2053 3.4105
R14073 GNDA.n2052 GNDA.n2051 3.4105
R14074 GNDA.n2050 GNDA.n2049 3.4105
R14075 GNDA.n2048 GNDA.n1973 3.4105
R14076 GNDA.n2044 GNDA.n2043 3.4105
R14077 GNDA.n2042 GNDA.n2041 3.4105
R14078 GNDA.n2040 GNDA.n2039 3.4105
R14079 GNDA.n2038 GNDA.n1975 3.4105
R14080 GNDA.n2034 GNDA.n2033 3.4105
R14081 GNDA.n2032 GNDA.n2031 3.4105
R14082 GNDA.n2030 GNDA.n2029 3.4105
R14083 GNDA.n2028 GNDA.n1977 3.4105
R14084 GNDA.n2024 GNDA.n2023 3.4105
R14085 GNDA.n2022 GNDA.n2021 3.4105
R14086 GNDA.n2020 GNDA.n2019 3.4105
R14087 GNDA.n2018 GNDA.n1979 3.4105
R14088 GNDA.n2014 GNDA.n2013 3.4105
R14089 GNDA.n2012 GNDA.n2011 3.4105
R14090 GNDA.n2010 GNDA.n2009 3.4105
R14091 GNDA.n2008 GNDA.n1981 3.4105
R14092 GNDA.n2004 GNDA.n2003 3.4105
R14093 GNDA.n2002 GNDA.n2001 3.4105
R14094 GNDA.n2000 GNDA.n1999 3.4105
R14095 GNDA.n1998 GNDA.n1983 3.4105
R14096 GNDA.n1994 GNDA.n1993 3.4105
R14097 GNDA.n1992 GNDA.n1991 3.4105
R14098 GNDA.n1990 GNDA.n1989 3.4105
R14099 GNDA.n1988 GNDA.n1985 3.4105
R14100 GNDA.n727 GNDA.n726 3.4105
R14101 GNDA.n2100 GNDA.n2099 3.4105
R14102 GNDA.n754 GNDA.n753 3.4105
R14103 GNDA.n1934 GNDA.n1933 3.4105
R14104 GNDA.n1932 GNDA.n1931 3.4105
R14105 GNDA.n1930 GNDA.n1929 3.4105
R14106 GNDA.n1928 GNDA.n756 3.4105
R14107 GNDA.n1924 GNDA.n1923 3.4105
R14108 GNDA.n1922 GNDA.n1921 3.4105
R14109 GNDA.n1920 GNDA.n1919 3.4105
R14110 GNDA.n1918 GNDA.n758 3.4105
R14111 GNDA.n1914 GNDA.n1913 3.4105
R14112 GNDA.n1912 GNDA.n1911 3.4105
R14113 GNDA.n1910 GNDA.n1909 3.4105
R14114 GNDA.n1908 GNDA.n760 3.4105
R14115 GNDA.n1904 GNDA.n1903 3.4105
R14116 GNDA.n1902 GNDA.n1901 3.4105
R14117 GNDA.n1900 GNDA.n1899 3.4105
R14118 GNDA.n1898 GNDA.n762 3.4105
R14119 GNDA.n1894 GNDA.n1893 3.4105
R14120 GNDA.n1892 GNDA.n1891 3.4105
R14121 GNDA.n1890 GNDA.n1889 3.4105
R14122 GNDA.n1888 GNDA.n764 3.4105
R14123 GNDA.n1884 GNDA.n1883 3.4105
R14124 GNDA.n1882 GNDA.n1881 3.4105
R14125 GNDA.n1880 GNDA.n1879 3.4105
R14126 GNDA.n1878 GNDA.n766 3.4105
R14127 GNDA.n1874 GNDA.n1873 3.4105
R14128 GNDA.n1872 GNDA.n1871 3.4105
R14129 GNDA.n1870 GNDA.n1869 3.4105
R14130 GNDA.n1868 GNDA.n768 3.4105
R14131 GNDA.n1864 GNDA.n1863 3.4105
R14132 GNDA.n1862 GNDA.n1861 3.4105
R14133 GNDA.n1860 GNDA.n1859 3.4105
R14134 GNDA.n1858 GNDA.n770 3.4105
R14135 GNDA.n1854 GNDA.n1853 3.4105
R14136 GNDA.n1852 GNDA.n1851 3.4105
R14137 GNDA.n1850 GNDA.n1849 3.4105
R14138 GNDA.n1848 GNDA.n772 3.4105
R14139 GNDA.n1844 GNDA.n1843 3.4105
R14140 GNDA.n1842 GNDA.n1841 3.4105
R14141 GNDA.n1840 GNDA.n1839 3.4105
R14142 GNDA.n1838 GNDA.n774 3.4105
R14143 GNDA.n1834 GNDA.n1833 3.4105
R14144 GNDA.n1832 GNDA.n1831 3.4105
R14145 GNDA.n1830 GNDA.n1829 3.4105
R14146 GNDA.n1828 GNDA.n776 3.4105
R14147 GNDA.n1824 GNDA.n1823 3.4105
R14148 GNDA.n1822 GNDA.n729 3.4105
R14149 GNDA.n1617 GNDA.n1570 3.4105
R14150 GNDA.n1619 GNDA.n1569 3.4105
R14151 GNDA.n1620 GNDA.n1568 3.4105
R14152 GNDA.n1622 GNDA.n1567 3.4105
R14153 GNDA.n1623 GNDA.n1566 3.4105
R14154 GNDA.n1625 GNDA.n1565 3.4105
R14155 GNDA.n1626 GNDA.n1564 3.4105
R14156 GNDA.n1628 GNDA.n1563 3.4105
R14157 GNDA.n1629 GNDA.n1562 3.4105
R14158 GNDA.n1631 GNDA.n1561 3.4105
R14159 GNDA.n1632 GNDA.n1560 3.4105
R14160 GNDA.n1634 GNDA.n1559 3.4105
R14161 GNDA.n1635 GNDA.n1558 3.4105
R14162 GNDA.n1637 GNDA.n1557 3.4105
R14163 GNDA.n1638 GNDA.n1556 3.4105
R14164 GNDA.n1640 GNDA.n1555 3.4105
R14165 GNDA.n1641 GNDA.n1554 3.4105
R14166 GNDA.n1643 GNDA.n1553 3.4105
R14167 GNDA.n1644 GNDA.n1552 3.4105
R14168 GNDA.n1646 GNDA.n1551 3.4105
R14169 GNDA.n1647 GNDA.n1550 3.4105
R14170 GNDA.n1649 GNDA.n1549 3.4105
R14171 GNDA.n1650 GNDA.n1548 3.4105
R14172 GNDA.n1652 GNDA.n1547 3.4105
R14173 GNDA.n1653 GNDA.n1546 3.4105
R14174 GNDA.n1655 GNDA.n1545 3.4105
R14175 GNDA.n1656 GNDA.n1544 3.4105
R14176 GNDA.n1658 GNDA.n1543 3.4105
R14177 GNDA.n1659 GNDA.n1542 3.4105
R14178 GNDA.n1661 GNDA.n1541 3.4105
R14179 GNDA.n1662 GNDA.n1540 3.4105
R14180 GNDA.n1664 GNDA.n1539 3.4105
R14181 GNDA.n1665 GNDA.n1538 3.4105
R14182 GNDA.n1667 GNDA.n1537 3.4105
R14183 GNDA.n1668 GNDA.n1536 3.4105
R14184 GNDA.n1670 GNDA.n1535 3.4105
R14185 GNDA.n1671 GNDA.n1534 3.4105
R14186 GNDA.n1673 GNDA.n1533 3.4105
R14187 GNDA.n1674 GNDA.n1532 3.4105
R14188 GNDA.n1676 GNDA.n1531 3.4105
R14189 GNDA.n1677 GNDA.n1530 3.4105
R14190 GNDA.n1679 GNDA.n1529 3.4105
R14191 GNDA.n1680 GNDA.n1528 3.4105
R14192 GNDA.n1682 GNDA.n1527 3.4105
R14193 GNDA.n1683 GNDA.n1526 3.4105
R14194 GNDA.n1685 GNDA.n1525 3.4105
R14195 GNDA.n1687 GNDA.n1686 3.4105
R14196 GNDA.n1379 GNDA.n1378 3.4105
R14197 GNDA.n1510 GNDA.n1509 3.4105
R14198 GNDA.n1508 GNDA.n1507 3.4105
R14199 GNDA.n1506 GNDA.n1505 3.4105
R14200 GNDA.n1504 GNDA.n1381 3.4105
R14201 GNDA.n1500 GNDA.n1499 3.4105
R14202 GNDA.n1498 GNDA.n1497 3.4105
R14203 GNDA.n1496 GNDA.n1495 3.4105
R14204 GNDA.n1494 GNDA.n1383 3.4105
R14205 GNDA.n1490 GNDA.n1489 3.4105
R14206 GNDA.n1488 GNDA.n1487 3.4105
R14207 GNDA.n1486 GNDA.n1485 3.4105
R14208 GNDA.n1484 GNDA.n1385 3.4105
R14209 GNDA.n1480 GNDA.n1479 3.4105
R14210 GNDA.n1478 GNDA.n1477 3.4105
R14211 GNDA.n1476 GNDA.n1475 3.4105
R14212 GNDA.n1474 GNDA.n1387 3.4105
R14213 GNDA.n1470 GNDA.n1469 3.4105
R14214 GNDA.n1468 GNDA.n1467 3.4105
R14215 GNDA.n1466 GNDA.n1465 3.4105
R14216 GNDA.n1464 GNDA.n1389 3.4105
R14217 GNDA.n1460 GNDA.n1459 3.4105
R14218 GNDA.n1458 GNDA.n1457 3.4105
R14219 GNDA.n1456 GNDA.n1455 3.4105
R14220 GNDA.n1454 GNDA.n1391 3.4105
R14221 GNDA.n1450 GNDA.n1449 3.4105
R14222 GNDA.n1448 GNDA.n1447 3.4105
R14223 GNDA.n1446 GNDA.n1445 3.4105
R14224 GNDA.n1444 GNDA.n1393 3.4105
R14225 GNDA.n1440 GNDA.n1439 3.4105
R14226 GNDA.n1438 GNDA.n1437 3.4105
R14227 GNDA.n1436 GNDA.n1435 3.4105
R14228 GNDA.n1434 GNDA.n1395 3.4105
R14229 GNDA.n1430 GNDA.n1429 3.4105
R14230 GNDA.n1428 GNDA.n1427 3.4105
R14231 GNDA.n1426 GNDA.n1425 3.4105
R14232 GNDA.n1424 GNDA.n1397 3.4105
R14233 GNDA.n1420 GNDA.n1419 3.4105
R14234 GNDA.n1418 GNDA.n1417 3.4105
R14235 GNDA.n1416 GNDA.n1415 3.4105
R14236 GNDA.n1414 GNDA.n1399 3.4105
R14237 GNDA.n1410 GNDA.n1409 3.4105
R14238 GNDA.n1408 GNDA.n1407 3.4105
R14239 GNDA.n1406 GNDA.n1405 3.4105
R14240 GNDA.n1404 GNDA.n1401 3.4105
R14241 GNDA.n793 GNDA.n792 3.4105
R14242 GNDA.n1516 GNDA.n1515 3.4105
R14243 GNDA.n1515 GNDA.n1514 3.4105
R14244 GNDA.n1514 GNDA.n1513 3.4105
R14245 GNDA.n1686 GNDA.n728 3.4105
R14246 GNDA.n1616 GNDA.n728 3.4105
R14247 GNDA.n1938 GNDA.n729 3.4105
R14248 GNDA.n1938 GNDA.n1937 3.4105
R14249 GNDA.n2099 GNDA.n2098 3.4105
R14250 GNDA.n2098 GNDA.n2097 3.4105
R14251 GNDA.n2273 GNDA.n665 3.4105
R14252 GNDA.n2203 GNDA.n665 3.4105
R14253 GNDA.n2562 GNDA.n2561 3.4105
R14254 GNDA.n2561 GNDA.n2560 3.4105
R14255 GNDA.n2733 GNDA.n599 3.4105
R14256 GNDA.n2663 GNDA.n599 3.4105
R14257 GNDA.n2863 GNDA.n600 3.4105
R14258 GNDA.n2863 GNDA.n2862 3.4105
R14259 GNDA.n2401 GNDA.n666 3.4105
R14260 GNDA.n2401 GNDA.n2400 3.4105
R14261 GNDA.n3037 GNDA.n2864 3.4105
R14262 GNDA.n3037 GNDA.n3036 3.4105
R14263 GNDA.n3198 GNDA.n3197 3.4105
R14264 GNDA.n3197 GNDA.n3196 3.4105
R14265 GNDA.n3370 GNDA.n329 3.4105
R14266 GNDA.n3300 GNDA.n329 3.4105
R14267 GNDA.n5135 GNDA.n353 3.4105
R14268 GNDA.n5135 GNDA.n5134 3.4105
R14269 GNDA.n567 GNDA.n377 3.4105
R14270 GNDA.n497 GNDA.n377 3.4105
R14271 GNDA.n3673 GNDA.n3459 3.4105
R14272 GNDA.n3603 GNDA.n3459 3.4105
R14273 GNDA.n3969 GNDA.n3804 3.4105
R14274 GNDA.n3969 GNDA.n3968 3.4105
R14275 GNDA.n4135 GNDA.n3970 3.4105
R14276 GNDA.n4135 GNDA.n4134 3.4105
R14277 GNDA.n3803 GNDA.n3460 3.4105
R14278 GNDA.n3803 GNDA.n3802 3.4105
R14279 GNDA.n4301 GNDA.n4136 3.4105
R14280 GNDA.n4301 GNDA.n4300 3.4105
R14281 GNDA.n4467 GNDA.n4302 3.4105
R14282 GNDA.n4467 GNDA.n4466 3.4105
R14283 GNDA.n4633 GNDA.n4468 3.4105
R14284 GNDA.n4633 GNDA.n4632 3.4105
R14285 GNDA.n4799 GNDA.n4634 3.4105
R14286 GNDA.n4799 GNDA.n4798 3.4105
R14287 GNDA.n4960 GNDA.n4959 3.4105
R14288 GNDA.n4959 GNDA.n4958 3.4105
R14289 GNDA.n5273 GNDA.n5272 3.4105
R14290 GNDA.n5272 GNDA.n5271 3.4105
R14291 GNDA.n1193 GNDA.n1191 3.4105
R14292 GNDA.n1352 GNDA.n1351 3.4105
R14293 GNDA.n1192 GNDA.n1190 3.4105
R14294 GNDA.n1346 GNDA.n1345 3.4105
R14295 GNDA.n1344 GNDA.n1343 3.4105
R14296 GNDA.n1342 GNDA.n1341 3.4105
R14297 GNDA.n1335 GNDA.n1195 3.4105
R14298 GNDA.n1337 GNDA.n1336 3.4105
R14299 GNDA.n1334 GNDA.n1333 3.4105
R14300 GNDA.n1332 GNDA.n1331 3.4105
R14301 GNDA.n1325 GNDA.n1197 3.4105
R14302 GNDA.n1327 GNDA.n1326 3.4105
R14303 GNDA.n1324 GNDA.n1323 3.4105
R14304 GNDA.n1322 GNDA.n1321 3.4105
R14305 GNDA.n1315 GNDA.n1199 3.4105
R14306 GNDA.n1317 GNDA.n1316 3.4105
R14307 GNDA.n1314 GNDA.n1313 3.4105
R14308 GNDA.n1312 GNDA.n1311 3.4105
R14309 GNDA.n1305 GNDA.n1201 3.4105
R14310 GNDA.n1307 GNDA.n1306 3.4105
R14311 GNDA.n1304 GNDA.n1303 3.4105
R14312 GNDA.n1302 GNDA.n1301 3.4105
R14313 GNDA.n1295 GNDA.n1203 3.4105
R14314 GNDA.n1297 GNDA.n1296 3.4105
R14315 GNDA.n1294 GNDA.n1293 3.4105
R14316 GNDA.n1292 GNDA.n1291 3.4105
R14317 GNDA.n1285 GNDA.n1205 3.4105
R14318 GNDA.n1287 GNDA.n1286 3.4105
R14319 GNDA.n1284 GNDA.n1283 3.4105
R14320 GNDA.n1282 GNDA.n1281 3.4105
R14321 GNDA.n1275 GNDA.n1207 3.4105
R14322 GNDA.n1277 GNDA.n1276 3.4105
R14323 GNDA.n1274 GNDA.n1273 3.4105
R14324 GNDA.n1272 GNDA.n1271 3.4105
R14325 GNDA.n1265 GNDA.n1209 3.4105
R14326 GNDA.n1267 GNDA.n1266 3.4105
R14327 GNDA.n1264 GNDA.n1263 3.4105
R14328 GNDA.n1262 GNDA.n1261 3.4105
R14329 GNDA.n1255 GNDA.n1211 3.4105
R14330 GNDA.n1257 GNDA.n1256 3.4105
R14331 GNDA.n1254 GNDA.n1253 3.4105
R14332 GNDA.n1252 GNDA.n1251 3.4105
R14333 GNDA.n1245 GNDA.n1213 3.4105
R14334 GNDA.n1247 GNDA.n1246 3.4105
R14335 GNDA.n1244 GNDA.n1243 3.4105
R14336 GNDA.n1242 GNDA.n1241 3.4105
R14337 GNDA.n97 GNDA.n96 3.4105
R14338 GNDA.n7223 GNDA.n7222 3.4105
R14339 GNDA.n7090 GNDA.n7089 3.4105
R14340 GNDA.n7218 GNDA.n7217 3.4105
R14341 GNDA.n7216 GNDA.n7215 3.4105
R14342 GNDA.n7214 GNDA.n7094 3.4105
R14343 GNDA.n7093 GNDA.n7092 3.4105
R14344 GNDA.n7210 GNDA.n7209 3.4105
R14345 GNDA.n7208 GNDA.n7207 3.4105
R14346 GNDA.n7206 GNDA.n7098 3.4105
R14347 GNDA.n7097 GNDA.n7096 3.4105
R14348 GNDA.n7202 GNDA.n7201 3.4105
R14349 GNDA.n7200 GNDA.n7199 3.4105
R14350 GNDA.n7198 GNDA.n7102 3.4105
R14351 GNDA.n7101 GNDA.n7100 3.4105
R14352 GNDA.n7194 GNDA.n7193 3.4105
R14353 GNDA.n7192 GNDA.n7191 3.4105
R14354 GNDA.n7190 GNDA.n7106 3.4105
R14355 GNDA.n7105 GNDA.n7104 3.4105
R14356 GNDA.n7186 GNDA.n7185 3.4105
R14357 GNDA.n7184 GNDA.n7183 3.4105
R14358 GNDA.n7182 GNDA.n7110 3.4105
R14359 GNDA.n7109 GNDA.n7108 3.4105
R14360 GNDA.n7178 GNDA.n7177 3.4105
R14361 GNDA.n7176 GNDA.n7175 3.4105
R14362 GNDA.n7174 GNDA.n7114 3.4105
R14363 GNDA.n7113 GNDA.n7112 3.4105
R14364 GNDA.n7170 GNDA.n7169 3.4105
R14365 GNDA.n7168 GNDA.n7167 3.4105
R14366 GNDA.n7166 GNDA.n7118 3.4105
R14367 GNDA.n7117 GNDA.n7116 3.4105
R14368 GNDA.n7162 GNDA.n7161 3.4105
R14369 GNDA.n7160 GNDA.n7159 3.4105
R14370 GNDA.n7158 GNDA.n7122 3.4105
R14371 GNDA.n7121 GNDA.n7120 3.4105
R14372 GNDA.n7154 GNDA.n7153 3.4105
R14373 GNDA.n7152 GNDA.n7151 3.4105
R14374 GNDA.n7150 GNDA.n7126 3.4105
R14375 GNDA.n7125 GNDA.n7124 3.4105
R14376 GNDA.n7146 GNDA.n7145 3.4105
R14377 GNDA.n7144 GNDA.n7143 3.4105
R14378 GNDA.n7142 GNDA.n7130 3.4105
R14379 GNDA.n7129 GNDA.n7128 3.4105
R14380 GNDA.n7138 GNDA.n7137 3.4105
R14381 GNDA.n7136 GNDA.n7135 3.4105
R14382 GNDA.n7134 GNDA.n7133 3.4105
R14383 GNDA.n7227 GNDA.n7226 3.4105
R14384 GNDA.n124 GNDA.n123 3.4105
R14385 GNDA.n258 GNDA.n257 3.4105
R14386 GNDA.n256 GNDA.n255 3.4105
R14387 GNDA.n254 GNDA.n253 3.4105
R14388 GNDA.n252 GNDA.n126 3.4105
R14389 GNDA.n248 GNDA.n247 3.4105
R14390 GNDA.n246 GNDA.n245 3.4105
R14391 GNDA.n244 GNDA.n243 3.4105
R14392 GNDA.n242 GNDA.n128 3.4105
R14393 GNDA.n238 GNDA.n237 3.4105
R14394 GNDA.n236 GNDA.n235 3.4105
R14395 GNDA.n234 GNDA.n233 3.4105
R14396 GNDA.n232 GNDA.n130 3.4105
R14397 GNDA.n228 GNDA.n227 3.4105
R14398 GNDA.n226 GNDA.n225 3.4105
R14399 GNDA.n224 GNDA.n223 3.4105
R14400 GNDA.n222 GNDA.n132 3.4105
R14401 GNDA.n218 GNDA.n217 3.4105
R14402 GNDA.n216 GNDA.n215 3.4105
R14403 GNDA.n214 GNDA.n213 3.4105
R14404 GNDA.n212 GNDA.n134 3.4105
R14405 GNDA.n208 GNDA.n207 3.4105
R14406 GNDA.n206 GNDA.n205 3.4105
R14407 GNDA.n204 GNDA.n203 3.4105
R14408 GNDA.n202 GNDA.n136 3.4105
R14409 GNDA.n198 GNDA.n197 3.4105
R14410 GNDA.n196 GNDA.n195 3.4105
R14411 GNDA.n194 GNDA.n193 3.4105
R14412 GNDA.n192 GNDA.n138 3.4105
R14413 GNDA.n188 GNDA.n187 3.4105
R14414 GNDA.n186 GNDA.n185 3.4105
R14415 GNDA.n184 GNDA.n183 3.4105
R14416 GNDA.n182 GNDA.n140 3.4105
R14417 GNDA.n178 GNDA.n177 3.4105
R14418 GNDA.n176 GNDA.n175 3.4105
R14419 GNDA.n174 GNDA.n173 3.4105
R14420 GNDA.n172 GNDA.n142 3.4105
R14421 GNDA.n168 GNDA.n167 3.4105
R14422 GNDA.n166 GNDA.n165 3.4105
R14423 GNDA.n164 GNDA.n163 3.4105
R14424 GNDA.n162 GNDA.n144 3.4105
R14425 GNDA.n158 GNDA.n157 3.4105
R14426 GNDA.n156 GNDA.n155 3.4105
R14427 GNDA.n154 GNDA.n153 3.4105
R14428 GNDA.n152 GNDA.n146 3.4105
R14429 GNDA.n148 GNDA.n147 3.4105
R14430 GNDA.n7064 GNDA.n7063 3.4105
R14431 GNDA.n7065 GNDA.n99 3.4105
R14432 GNDA.n7065 GNDA.n7064 3.4105
R14433 GNDA.n7225 GNDA.n7066 3.4105
R14434 GNDA.n7226 GNDA.n7225 3.4105
R14435 GNDA.n974 GNDA.n98 3.4105
R14436 GNDA.n974 GNDA.n945 3.4105
R14437 GNDA.n1037 GNDA.n974 3.4105
R14438 GNDA.n1035 GNDA.n992 3.4105
R14439 GNDA.n1037 GNDA.n992 3.4105
R14440 GNDA.n1035 GNDA.n960 3.4105
R14441 GNDA.n960 GNDA.n930 3.4105
R14442 GNDA.n960 GNDA.n932 3.4105
R14443 GNDA.n960 GNDA.n929 3.4105
R14444 GNDA.n960 GNDA.n933 3.4105
R14445 GNDA.n960 GNDA.n928 3.4105
R14446 GNDA.n960 GNDA.n934 3.4105
R14447 GNDA.n960 GNDA.n927 3.4105
R14448 GNDA.n960 GNDA.n935 3.4105
R14449 GNDA.n960 GNDA.n926 3.4105
R14450 GNDA.n960 GNDA.n936 3.4105
R14451 GNDA.n960 GNDA.n925 3.4105
R14452 GNDA.n960 GNDA.n937 3.4105
R14453 GNDA.n960 GNDA.n924 3.4105
R14454 GNDA.n960 GNDA.n938 3.4105
R14455 GNDA.n960 GNDA.n923 3.4105
R14456 GNDA.n960 GNDA.n939 3.4105
R14457 GNDA.n960 GNDA.n922 3.4105
R14458 GNDA.n960 GNDA.n940 3.4105
R14459 GNDA.n960 GNDA.n921 3.4105
R14460 GNDA.n960 GNDA.n941 3.4105
R14461 GNDA.n960 GNDA.n920 3.4105
R14462 GNDA.n960 GNDA.n942 3.4105
R14463 GNDA.n960 GNDA.n919 3.4105
R14464 GNDA.n960 GNDA.n943 3.4105
R14465 GNDA.n960 GNDA.n918 3.4105
R14466 GNDA.n960 GNDA.n944 3.4105
R14467 GNDA.n960 GNDA.n917 3.4105
R14468 GNDA.n960 GNDA.n945 3.4105
R14469 GNDA.n1037 GNDA.n960 3.4105
R14470 GNDA.n1035 GNDA.n995 3.4105
R14471 GNDA.n995 GNDA.n930 3.4105
R14472 GNDA.n995 GNDA.n932 3.4105
R14473 GNDA.n995 GNDA.n929 3.4105
R14474 GNDA.n995 GNDA.n933 3.4105
R14475 GNDA.n995 GNDA.n928 3.4105
R14476 GNDA.n995 GNDA.n934 3.4105
R14477 GNDA.n995 GNDA.n927 3.4105
R14478 GNDA.n995 GNDA.n935 3.4105
R14479 GNDA.n995 GNDA.n926 3.4105
R14480 GNDA.n995 GNDA.n936 3.4105
R14481 GNDA.n995 GNDA.n925 3.4105
R14482 GNDA.n995 GNDA.n937 3.4105
R14483 GNDA.n995 GNDA.n924 3.4105
R14484 GNDA.n995 GNDA.n938 3.4105
R14485 GNDA.n995 GNDA.n923 3.4105
R14486 GNDA.n995 GNDA.n939 3.4105
R14487 GNDA.n995 GNDA.n922 3.4105
R14488 GNDA.n995 GNDA.n940 3.4105
R14489 GNDA.n995 GNDA.n921 3.4105
R14490 GNDA.n995 GNDA.n941 3.4105
R14491 GNDA.n995 GNDA.n920 3.4105
R14492 GNDA.n995 GNDA.n942 3.4105
R14493 GNDA.n995 GNDA.n919 3.4105
R14494 GNDA.n995 GNDA.n943 3.4105
R14495 GNDA.n995 GNDA.n918 3.4105
R14496 GNDA.n995 GNDA.n944 3.4105
R14497 GNDA.n995 GNDA.n917 3.4105
R14498 GNDA.n995 GNDA.n945 3.4105
R14499 GNDA.n1037 GNDA.n995 3.4105
R14500 GNDA.n1035 GNDA.n959 3.4105
R14501 GNDA.n959 GNDA.n930 3.4105
R14502 GNDA.n959 GNDA.n932 3.4105
R14503 GNDA.n959 GNDA.n929 3.4105
R14504 GNDA.n959 GNDA.n933 3.4105
R14505 GNDA.n959 GNDA.n928 3.4105
R14506 GNDA.n959 GNDA.n934 3.4105
R14507 GNDA.n959 GNDA.n927 3.4105
R14508 GNDA.n959 GNDA.n935 3.4105
R14509 GNDA.n959 GNDA.n926 3.4105
R14510 GNDA.n959 GNDA.n936 3.4105
R14511 GNDA.n959 GNDA.n925 3.4105
R14512 GNDA.n959 GNDA.n937 3.4105
R14513 GNDA.n959 GNDA.n924 3.4105
R14514 GNDA.n959 GNDA.n938 3.4105
R14515 GNDA.n959 GNDA.n923 3.4105
R14516 GNDA.n959 GNDA.n939 3.4105
R14517 GNDA.n959 GNDA.n922 3.4105
R14518 GNDA.n959 GNDA.n940 3.4105
R14519 GNDA.n959 GNDA.n921 3.4105
R14520 GNDA.n959 GNDA.n941 3.4105
R14521 GNDA.n959 GNDA.n920 3.4105
R14522 GNDA.n959 GNDA.n942 3.4105
R14523 GNDA.n959 GNDA.n919 3.4105
R14524 GNDA.n959 GNDA.n943 3.4105
R14525 GNDA.n959 GNDA.n918 3.4105
R14526 GNDA.n959 GNDA.n944 3.4105
R14527 GNDA.n959 GNDA.n917 3.4105
R14528 GNDA.n959 GNDA.n945 3.4105
R14529 GNDA.n1037 GNDA.n959 3.4105
R14530 GNDA.n1035 GNDA.n998 3.4105
R14531 GNDA.n998 GNDA.n930 3.4105
R14532 GNDA.n998 GNDA.n932 3.4105
R14533 GNDA.n998 GNDA.n929 3.4105
R14534 GNDA.n998 GNDA.n933 3.4105
R14535 GNDA.n998 GNDA.n928 3.4105
R14536 GNDA.n998 GNDA.n934 3.4105
R14537 GNDA.n998 GNDA.n927 3.4105
R14538 GNDA.n998 GNDA.n935 3.4105
R14539 GNDA.n998 GNDA.n926 3.4105
R14540 GNDA.n998 GNDA.n936 3.4105
R14541 GNDA.n998 GNDA.n925 3.4105
R14542 GNDA.n998 GNDA.n937 3.4105
R14543 GNDA.n998 GNDA.n924 3.4105
R14544 GNDA.n998 GNDA.n938 3.4105
R14545 GNDA.n998 GNDA.n923 3.4105
R14546 GNDA.n998 GNDA.n939 3.4105
R14547 GNDA.n998 GNDA.n922 3.4105
R14548 GNDA.n998 GNDA.n940 3.4105
R14549 GNDA.n998 GNDA.n921 3.4105
R14550 GNDA.n998 GNDA.n941 3.4105
R14551 GNDA.n998 GNDA.n920 3.4105
R14552 GNDA.n998 GNDA.n942 3.4105
R14553 GNDA.n998 GNDA.n919 3.4105
R14554 GNDA.n998 GNDA.n943 3.4105
R14555 GNDA.n998 GNDA.n918 3.4105
R14556 GNDA.n998 GNDA.n944 3.4105
R14557 GNDA.n998 GNDA.n917 3.4105
R14558 GNDA.n998 GNDA.n945 3.4105
R14559 GNDA.n1037 GNDA.n998 3.4105
R14560 GNDA.n1035 GNDA.n958 3.4105
R14561 GNDA.n958 GNDA.n930 3.4105
R14562 GNDA.n958 GNDA.n932 3.4105
R14563 GNDA.n958 GNDA.n929 3.4105
R14564 GNDA.n958 GNDA.n933 3.4105
R14565 GNDA.n958 GNDA.n928 3.4105
R14566 GNDA.n958 GNDA.n934 3.4105
R14567 GNDA.n958 GNDA.n927 3.4105
R14568 GNDA.n958 GNDA.n935 3.4105
R14569 GNDA.n958 GNDA.n926 3.4105
R14570 GNDA.n958 GNDA.n936 3.4105
R14571 GNDA.n958 GNDA.n925 3.4105
R14572 GNDA.n958 GNDA.n937 3.4105
R14573 GNDA.n958 GNDA.n924 3.4105
R14574 GNDA.n958 GNDA.n938 3.4105
R14575 GNDA.n958 GNDA.n923 3.4105
R14576 GNDA.n958 GNDA.n939 3.4105
R14577 GNDA.n958 GNDA.n922 3.4105
R14578 GNDA.n958 GNDA.n940 3.4105
R14579 GNDA.n958 GNDA.n921 3.4105
R14580 GNDA.n958 GNDA.n941 3.4105
R14581 GNDA.n958 GNDA.n920 3.4105
R14582 GNDA.n958 GNDA.n942 3.4105
R14583 GNDA.n958 GNDA.n919 3.4105
R14584 GNDA.n958 GNDA.n943 3.4105
R14585 GNDA.n958 GNDA.n918 3.4105
R14586 GNDA.n958 GNDA.n944 3.4105
R14587 GNDA.n958 GNDA.n917 3.4105
R14588 GNDA.n958 GNDA.n945 3.4105
R14589 GNDA.n1037 GNDA.n958 3.4105
R14590 GNDA.n1035 GNDA.n1001 3.4105
R14591 GNDA.n1001 GNDA.n930 3.4105
R14592 GNDA.n1001 GNDA.n932 3.4105
R14593 GNDA.n1001 GNDA.n929 3.4105
R14594 GNDA.n1001 GNDA.n933 3.4105
R14595 GNDA.n1001 GNDA.n928 3.4105
R14596 GNDA.n1001 GNDA.n934 3.4105
R14597 GNDA.n1001 GNDA.n927 3.4105
R14598 GNDA.n1001 GNDA.n935 3.4105
R14599 GNDA.n1001 GNDA.n926 3.4105
R14600 GNDA.n1001 GNDA.n936 3.4105
R14601 GNDA.n1001 GNDA.n925 3.4105
R14602 GNDA.n1001 GNDA.n937 3.4105
R14603 GNDA.n1001 GNDA.n924 3.4105
R14604 GNDA.n1001 GNDA.n938 3.4105
R14605 GNDA.n1001 GNDA.n923 3.4105
R14606 GNDA.n1001 GNDA.n939 3.4105
R14607 GNDA.n1001 GNDA.n922 3.4105
R14608 GNDA.n1001 GNDA.n940 3.4105
R14609 GNDA.n1001 GNDA.n921 3.4105
R14610 GNDA.n1001 GNDA.n941 3.4105
R14611 GNDA.n1001 GNDA.n920 3.4105
R14612 GNDA.n1001 GNDA.n942 3.4105
R14613 GNDA.n1001 GNDA.n919 3.4105
R14614 GNDA.n1001 GNDA.n943 3.4105
R14615 GNDA.n1001 GNDA.n918 3.4105
R14616 GNDA.n1001 GNDA.n944 3.4105
R14617 GNDA.n1001 GNDA.n917 3.4105
R14618 GNDA.n1001 GNDA.n945 3.4105
R14619 GNDA.n1037 GNDA.n1001 3.4105
R14620 GNDA.n1035 GNDA.n957 3.4105
R14621 GNDA.n957 GNDA.n930 3.4105
R14622 GNDA.n957 GNDA.n932 3.4105
R14623 GNDA.n957 GNDA.n929 3.4105
R14624 GNDA.n957 GNDA.n933 3.4105
R14625 GNDA.n957 GNDA.n928 3.4105
R14626 GNDA.n957 GNDA.n934 3.4105
R14627 GNDA.n957 GNDA.n927 3.4105
R14628 GNDA.n957 GNDA.n935 3.4105
R14629 GNDA.n957 GNDA.n926 3.4105
R14630 GNDA.n957 GNDA.n936 3.4105
R14631 GNDA.n957 GNDA.n925 3.4105
R14632 GNDA.n957 GNDA.n937 3.4105
R14633 GNDA.n957 GNDA.n924 3.4105
R14634 GNDA.n957 GNDA.n938 3.4105
R14635 GNDA.n957 GNDA.n923 3.4105
R14636 GNDA.n957 GNDA.n939 3.4105
R14637 GNDA.n957 GNDA.n922 3.4105
R14638 GNDA.n957 GNDA.n940 3.4105
R14639 GNDA.n957 GNDA.n921 3.4105
R14640 GNDA.n957 GNDA.n941 3.4105
R14641 GNDA.n957 GNDA.n920 3.4105
R14642 GNDA.n957 GNDA.n942 3.4105
R14643 GNDA.n957 GNDA.n919 3.4105
R14644 GNDA.n957 GNDA.n943 3.4105
R14645 GNDA.n957 GNDA.n918 3.4105
R14646 GNDA.n957 GNDA.n944 3.4105
R14647 GNDA.n957 GNDA.n917 3.4105
R14648 GNDA.n957 GNDA.n945 3.4105
R14649 GNDA.n1037 GNDA.n957 3.4105
R14650 GNDA.n1035 GNDA.n1004 3.4105
R14651 GNDA.n1004 GNDA.n930 3.4105
R14652 GNDA.n1004 GNDA.n932 3.4105
R14653 GNDA.n1004 GNDA.n929 3.4105
R14654 GNDA.n1004 GNDA.n933 3.4105
R14655 GNDA.n1004 GNDA.n928 3.4105
R14656 GNDA.n1004 GNDA.n934 3.4105
R14657 GNDA.n1004 GNDA.n927 3.4105
R14658 GNDA.n1004 GNDA.n935 3.4105
R14659 GNDA.n1004 GNDA.n926 3.4105
R14660 GNDA.n1004 GNDA.n936 3.4105
R14661 GNDA.n1004 GNDA.n925 3.4105
R14662 GNDA.n1004 GNDA.n937 3.4105
R14663 GNDA.n1004 GNDA.n924 3.4105
R14664 GNDA.n1004 GNDA.n938 3.4105
R14665 GNDA.n1004 GNDA.n923 3.4105
R14666 GNDA.n1004 GNDA.n939 3.4105
R14667 GNDA.n1004 GNDA.n922 3.4105
R14668 GNDA.n1004 GNDA.n940 3.4105
R14669 GNDA.n1004 GNDA.n921 3.4105
R14670 GNDA.n1004 GNDA.n941 3.4105
R14671 GNDA.n1004 GNDA.n920 3.4105
R14672 GNDA.n1004 GNDA.n942 3.4105
R14673 GNDA.n1004 GNDA.n919 3.4105
R14674 GNDA.n1004 GNDA.n943 3.4105
R14675 GNDA.n1004 GNDA.n918 3.4105
R14676 GNDA.n1004 GNDA.n944 3.4105
R14677 GNDA.n1004 GNDA.n917 3.4105
R14678 GNDA.n1004 GNDA.n945 3.4105
R14679 GNDA.n1037 GNDA.n1004 3.4105
R14680 GNDA.n1035 GNDA.n956 3.4105
R14681 GNDA.n956 GNDA.n930 3.4105
R14682 GNDA.n956 GNDA.n932 3.4105
R14683 GNDA.n956 GNDA.n929 3.4105
R14684 GNDA.n956 GNDA.n933 3.4105
R14685 GNDA.n956 GNDA.n928 3.4105
R14686 GNDA.n956 GNDA.n934 3.4105
R14687 GNDA.n956 GNDA.n927 3.4105
R14688 GNDA.n956 GNDA.n935 3.4105
R14689 GNDA.n956 GNDA.n926 3.4105
R14690 GNDA.n956 GNDA.n936 3.4105
R14691 GNDA.n956 GNDA.n925 3.4105
R14692 GNDA.n956 GNDA.n937 3.4105
R14693 GNDA.n956 GNDA.n924 3.4105
R14694 GNDA.n956 GNDA.n938 3.4105
R14695 GNDA.n956 GNDA.n923 3.4105
R14696 GNDA.n956 GNDA.n939 3.4105
R14697 GNDA.n956 GNDA.n922 3.4105
R14698 GNDA.n956 GNDA.n940 3.4105
R14699 GNDA.n956 GNDA.n921 3.4105
R14700 GNDA.n956 GNDA.n941 3.4105
R14701 GNDA.n956 GNDA.n920 3.4105
R14702 GNDA.n956 GNDA.n942 3.4105
R14703 GNDA.n956 GNDA.n919 3.4105
R14704 GNDA.n956 GNDA.n943 3.4105
R14705 GNDA.n956 GNDA.n918 3.4105
R14706 GNDA.n956 GNDA.n944 3.4105
R14707 GNDA.n956 GNDA.n917 3.4105
R14708 GNDA.n956 GNDA.n945 3.4105
R14709 GNDA.n1037 GNDA.n956 3.4105
R14710 GNDA.n1035 GNDA.n1007 3.4105
R14711 GNDA.n1007 GNDA.n930 3.4105
R14712 GNDA.n1007 GNDA.n932 3.4105
R14713 GNDA.n1007 GNDA.n929 3.4105
R14714 GNDA.n1007 GNDA.n933 3.4105
R14715 GNDA.n1007 GNDA.n928 3.4105
R14716 GNDA.n1007 GNDA.n934 3.4105
R14717 GNDA.n1007 GNDA.n927 3.4105
R14718 GNDA.n1007 GNDA.n935 3.4105
R14719 GNDA.n1007 GNDA.n926 3.4105
R14720 GNDA.n1007 GNDA.n936 3.4105
R14721 GNDA.n1007 GNDA.n925 3.4105
R14722 GNDA.n1007 GNDA.n937 3.4105
R14723 GNDA.n1007 GNDA.n924 3.4105
R14724 GNDA.n1007 GNDA.n938 3.4105
R14725 GNDA.n1007 GNDA.n923 3.4105
R14726 GNDA.n1007 GNDA.n939 3.4105
R14727 GNDA.n1007 GNDA.n922 3.4105
R14728 GNDA.n1007 GNDA.n940 3.4105
R14729 GNDA.n1007 GNDA.n921 3.4105
R14730 GNDA.n1007 GNDA.n941 3.4105
R14731 GNDA.n1007 GNDA.n920 3.4105
R14732 GNDA.n1007 GNDA.n942 3.4105
R14733 GNDA.n1007 GNDA.n919 3.4105
R14734 GNDA.n1007 GNDA.n943 3.4105
R14735 GNDA.n1007 GNDA.n918 3.4105
R14736 GNDA.n1007 GNDA.n944 3.4105
R14737 GNDA.n1007 GNDA.n917 3.4105
R14738 GNDA.n1007 GNDA.n945 3.4105
R14739 GNDA.n1037 GNDA.n1007 3.4105
R14740 GNDA.n1035 GNDA.n955 3.4105
R14741 GNDA.n955 GNDA.n930 3.4105
R14742 GNDA.n955 GNDA.n932 3.4105
R14743 GNDA.n955 GNDA.n929 3.4105
R14744 GNDA.n955 GNDA.n933 3.4105
R14745 GNDA.n955 GNDA.n928 3.4105
R14746 GNDA.n955 GNDA.n934 3.4105
R14747 GNDA.n955 GNDA.n927 3.4105
R14748 GNDA.n955 GNDA.n935 3.4105
R14749 GNDA.n955 GNDA.n926 3.4105
R14750 GNDA.n955 GNDA.n936 3.4105
R14751 GNDA.n955 GNDA.n925 3.4105
R14752 GNDA.n955 GNDA.n937 3.4105
R14753 GNDA.n955 GNDA.n924 3.4105
R14754 GNDA.n955 GNDA.n938 3.4105
R14755 GNDA.n955 GNDA.n923 3.4105
R14756 GNDA.n955 GNDA.n939 3.4105
R14757 GNDA.n955 GNDA.n922 3.4105
R14758 GNDA.n955 GNDA.n940 3.4105
R14759 GNDA.n955 GNDA.n921 3.4105
R14760 GNDA.n955 GNDA.n941 3.4105
R14761 GNDA.n955 GNDA.n920 3.4105
R14762 GNDA.n955 GNDA.n942 3.4105
R14763 GNDA.n955 GNDA.n919 3.4105
R14764 GNDA.n955 GNDA.n943 3.4105
R14765 GNDA.n955 GNDA.n918 3.4105
R14766 GNDA.n955 GNDA.n944 3.4105
R14767 GNDA.n955 GNDA.n917 3.4105
R14768 GNDA.n955 GNDA.n945 3.4105
R14769 GNDA.n1037 GNDA.n955 3.4105
R14770 GNDA.n1035 GNDA.n1010 3.4105
R14771 GNDA.n1010 GNDA.n930 3.4105
R14772 GNDA.n1010 GNDA.n932 3.4105
R14773 GNDA.n1010 GNDA.n929 3.4105
R14774 GNDA.n1010 GNDA.n933 3.4105
R14775 GNDA.n1010 GNDA.n928 3.4105
R14776 GNDA.n1010 GNDA.n934 3.4105
R14777 GNDA.n1010 GNDA.n927 3.4105
R14778 GNDA.n1010 GNDA.n935 3.4105
R14779 GNDA.n1010 GNDA.n926 3.4105
R14780 GNDA.n1010 GNDA.n936 3.4105
R14781 GNDA.n1010 GNDA.n925 3.4105
R14782 GNDA.n1010 GNDA.n937 3.4105
R14783 GNDA.n1010 GNDA.n924 3.4105
R14784 GNDA.n1010 GNDA.n938 3.4105
R14785 GNDA.n1010 GNDA.n923 3.4105
R14786 GNDA.n1010 GNDA.n939 3.4105
R14787 GNDA.n1010 GNDA.n922 3.4105
R14788 GNDA.n1010 GNDA.n940 3.4105
R14789 GNDA.n1010 GNDA.n921 3.4105
R14790 GNDA.n1010 GNDA.n941 3.4105
R14791 GNDA.n1010 GNDA.n920 3.4105
R14792 GNDA.n1010 GNDA.n942 3.4105
R14793 GNDA.n1010 GNDA.n919 3.4105
R14794 GNDA.n1010 GNDA.n943 3.4105
R14795 GNDA.n1010 GNDA.n918 3.4105
R14796 GNDA.n1010 GNDA.n944 3.4105
R14797 GNDA.n1010 GNDA.n917 3.4105
R14798 GNDA.n1010 GNDA.n945 3.4105
R14799 GNDA.n1037 GNDA.n1010 3.4105
R14800 GNDA.n1035 GNDA.n954 3.4105
R14801 GNDA.n954 GNDA.n930 3.4105
R14802 GNDA.n954 GNDA.n932 3.4105
R14803 GNDA.n954 GNDA.n929 3.4105
R14804 GNDA.n954 GNDA.n933 3.4105
R14805 GNDA.n954 GNDA.n928 3.4105
R14806 GNDA.n954 GNDA.n934 3.4105
R14807 GNDA.n954 GNDA.n927 3.4105
R14808 GNDA.n954 GNDA.n935 3.4105
R14809 GNDA.n954 GNDA.n926 3.4105
R14810 GNDA.n954 GNDA.n936 3.4105
R14811 GNDA.n954 GNDA.n925 3.4105
R14812 GNDA.n954 GNDA.n937 3.4105
R14813 GNDA.n954 GNDA.n924 3.4105
R14814 GNDA.n954 GNDA.n938 3.4105
R14815 GNDA.n954 GNDA.n923 3.4105
R14816 GNDA.n954 GNDA.n939 3.4105
R14817 GNDA.n954 GNDA.n922 3.4105
R14818 GNDA.n954 GNDA.n940 3.4105
R14819 GNDA.n954 GNDA.n921 3.4105
R14820 GNDA.n954 GNDA.n941 3.4105
R14821 GNDA.n954 GNDA.n920 3.4105
R14822 GNDA.n954 GNDA.n942 3.4105
R14823 GNDA.n954 GNDA.n919 3.4105
R14824 GNDA.n954 GNDA.n943 3.4105
R14825 GNDA.n954 GNDA.n918 3.4105
R14826 GNDA.n954 GNDA.n944 3.4105
R14827 GNDA.n954 GNDA.n917 3.4105
R14828 GNDA.n954 GNDA.n945 3.4105
R14829 GNDA.n1037 GNDA.n954 3.4105
R14830 GNDA.n1035 GNDA.n1013 3.4105
R14831 GNDA.n1013 GNDA.n930 3.4105
R14832 GNDA.n1013 GNDA.n932 3.4105
R14833 GNDA.n1013 GNDA.n929 3.4105
R14834 GNDA.n1013 GNDA.n933 3.4105
R14835 GNDA.n1013 GNDA.n928 3.4105
R14836 GNDA.n1013 GNDA.n934 3.4105
R14837 GNDA.n1013 GNDA.n927 3.4105
R14838 GNDA.n1013 GNDA.n935 3.4105
R14839 GNDA.n1013 GNDA.n926 3.4105
R14840 GNDA.n1013 GNDA.n936 3.4105
R14841 GNDA.n1013 GNDA.n925 3.4105
R14842 GNDA.n1013 GNDA.n937 3.4105
R14843 GNDA.n1013 GNDA.n924 3.4105
R14844 GNDA.n1013 GNDA.n938 3.4105
R14845 GNDA.n1013 GNDA.n923 3.4105
R14846 GNDA.n1013 GNDA.n939 3.4105
R14847 GNDA.n1013 GNDA.n922 3.4105
R14848 GNDA.n1013 GNDA.n940 3.4105
R14849 GNDA.n1013 GNDA.n921 3.4105
R14850 GNDA.n1013 GNDA.n941 3.4105
R14851 GNDA.n1013 GNDA.n920 3.4105
R14852 GNDA.n1013 GNDA.n942 3.4105
R14853 GNDA.n1013 GNDA.n919 3.4105
R14854 GNDA.n1013 GNDA.n943 3.4105
R14855 GNDA.n1013 GNDA.n918 3.4105
R14856 GNDA.n1013 GNDA.n944 3.4105
R14857 GNDA.n1013 GNDA.n917 3.4105
R14858 GNDA.n1013 GNDA.n945 3.4105
R14859 GNDA.n1037 GNDA.n1013 3.4105
R14860 GNDA.n1035 GNDA.n953 3.4105
R14861 GNDA.n953 GNDA.n930 3.4105
R14862 GNDA.n953 GNDA.n932 3.4105
R14863 GNDA.n953 GNDA.n929 3.4105
R14864 GNDA.n953 GNDA.n933 3.4105
R14865 GNDA.n953 GNDA.n928 3.4105
R14866 GNDA.n953 GNDA.n934 3.4105
R14867 GNDA.n953 GNDA.n927 3.4105
R14868 GNDA.n953 GNDA.n935 3.4105
R14869 GNDA.n953 GNDA.n926 3.4105
R14870 GNDA.n953 GNDA.n936 3.4105
R14871 GNDA.n953 GNDA.n925 3.4105
R14872 GNDA.n953 GNDA.n937 3.4105
R14873 GNDA.n953 GNDA.n924 3.4105
R14874 GNDA.n953 GNDA.n938 3.4105
R14875 GNDA.n953 GNDA.n923 3.4105
R14876 GNDA.n953 GNDA.n939 3.4105
R14877 GNDA.n953 GNDA.n922 3.4105
R14878 GNDA.n953 GNDA.n940 3.4105
R14879 GNDA.n953 GNDA.n921 3.4105
R14880 GNDA.n953 GNDA.n941 3.4105
R14881 GNDA.n953 GNDA.n920 3.4105
R14882 GNDA.n953 GNDA.n942 3.4105
R14883 GNDA.n953 GNDA.n919 3.4105
R14884 GNDA.n953 GNDA.n943 3.4105
R14885 GNDA.n953 GNDA.n918 3.4105
R14886 GNDA.n953 GNDA.n944 3.4105
R14887 GNDA.n953 GNDA.n917 3.4105
R14888 GNDA.n953 GNDA.n945 3.4105
R14889 GNDA.n1037 GNDA.n953 3.4105
R14890 GNDA.n1035 GNDA.n1016 3.4105
R14891 GNDA.n1016 GNDA.n930 3.4105
R14892 GNDA.n1016 GNDA.n932 3.4105
R14893 GNDA.n1016 GNDA.n929 3.4105
R14894 GNDA.n1016 GNDA.n933 3.4105
R14895 GNDA.n1016 GNDA.n928 3.4105
R14896 GNDA.n1016 GNDA.n934 3.4105
R14897 GNDA.n1016 GNDA.n927 3.4105
R14898 GNDA.n1016 GNDA.n935 3.4105
R14899 GNDA.n1016 GNDA.n926 3.4105
R14900 GNDA.n1016 GNDA.n936 3.4105
R14901 GNDA.n1016 GNDA.n925 3.4105
R14902 GNDA.n1016 GNDA.n937 3.4105
R14903 GNDA.n1016 GNDA.n924 3.4105
R14904 GNDA.n1016 GNDA.n938 3.4105
R14905 GNDA.n1016 GNDA.n923 3.4105
R14906 GNDA.n1016 GNDA.n939 3.4105
R14907 GNDA.n1016 GNDA.n922 3.4105
R14908 GNDA.n1016 GNDA.n940 3.4105
R14909 GNDA.n1016 GNDA.n921 3.4105
R14910 GNDA.n1016 GNDA.n941 3.4105
R14911 GNDA.n1016 GNDA.n920 3.4105
R14912 GNDA.n1016 GNDA.n942 3.4105
R14913 GNDA.n1016 GNDA.n919 3.4105
R14914 GNDA.n1016 GNDA.n943 3.4105
R14915 GNDA.n1016 GNDA.n918 3.4105
R14916 GNDA.n1016 GNDA.n944 3.4105
R14917 GNDA.n1016 GNDA.n917 3.4105
R14918 GNDA.n1016 GNDA.n945 3.4105
R14919 GNDA.n1037 GNDA.n1016 3.4105
R14920 GNDA.n1035 GNDA.n952 3.4105
R14921 GNDA.n952 GNDA.n930 3.4105
R14922 GNDA.n952 GNDA.n932 3.4105
R14923 GNDA.n952 GNDA.n929 3.4105
R14924 GNDA.n952 GNDA.n933 3.4105
R14925 GNDA.n952 GNDA.n928 3.4105
R14926 GNDA.n952 GNDA.n934 3.4105
R14927 GNDA.n952 GNDA.n927 3.4105
R14928 GNDA.n952 GNDA.n935 3.4105
R14929 GNDA.n952 GNDA.n926 3.4105
R14930 GNDA.n952 GNDA.n936 3.4105
R14931 GNDA.n952 GNDA.n925 3.4105
R14932 GNDA.n952 GNDA.n937 3.4105
R14933 GNDA.n952 GNDA.n924 3.4105
R14934 GNDA.n952 GNDA.n938 3.4105
R14935 GNDA.n952 GNDA.n923 3.4105
R14936 GNDA.n952 GNDA.n939 3.4105
R14937 GNDA.n952 GNDA.n922 3.4105
R14938 GNDA.n952 GNDA.n940 3.4105
R14939 GNDA.n952 GNDA.n921 3.4105
R14940 GNDA.n952 GNDA.n941 3.4105
R14941 GNDA.n952 GNDA.n920 3.4105
R14942 GNDA.n952 GNDA.n942 3.4105
R14943 GNDA.n952 GNDA.n919 3.4105
R14944 GNDA.n952 GNDA.n943 3.4105
R14945 GNDA.n952 GNDA.n918 3.4105
R14946 GNDA.n952 GNDA.n944 3.4105
R14947 GNDA.n952 GNDA.n917 3.4105
R14948 GNDA.n952 GNDA.n945 3.4105
R14949 GNDA.n1037 GNDA.n952 3.4105
R14950 GNDA.n1035 GNDA.n1019 3.4105
R14951 GNDA.n1019 GNDA.n930 3.4105
R14952 GNDA.n1019 GNDA.n932 3.4105
R14953 GNDA.n1019 GNDA.n929 3.4105
R14954 GNDA.n1019 GNDA.n933 3.4105
R14955 GNDA.n1019 GNDA.n928 3.4105
R14956 GNDA.n1019 GNDA.n934 3.4105
R14957 GNDA.n1019 GNDA.n927 3.4105
R14958 GNDA.n1019 GNDA.n935 3.4105
R14959 GNDA.n1019 GNDA.n926 3.4105
R14960 GNDA.n1019 GNDA.n936 3.4105
R14961 GNDA.n1019 GNDA.n925 3.4105
R14962 GNDA.n1019 GNDA.n937 3.4105
R14963 GNDA.n1019 GNDA.n924 3.4105
R14964 GNDA.n1019 GNDA.n938 3.4105
R14965 GNDA.n1019 GNDA.n923 3.4105
R14966 GNDA.n1019 GNDA.n939 3.4105
R14967 GNDA.n1019 GNDA.n922 3.4105
R14968 GNDA.n1019 GNDA.n940 3.4105
R14969 GNDA.n1019 GNDA.n921 3.4105
R14970 GNDA.n1019 GNDA.n941 3.4105
R14971 GNDA.n1019 GNDA.n920 3.4105
R14972 GNDA.n1019 GNDA.n942 3.4105
R14973 GNDA.n1019 GNDA.n919 3.4105
R14974 GNDA.n1019 GNDA.n943 3.4105
R14975 GNDA.n1019 GNDA.n918 3.4105
R14976 GNDA.n1019 GNDA.n944 3.4105
R14977 GNDA.n1019 GNDA.n917 3.4105
R14978 GNDA.n1019 GNDA.n945 3.4105
R14979 GNDA.n1037 GNDA.n1019 3.4105
R14980 GNDA.n1035 GNDA.n951 3.4105
R14981 GNDA.n951 GNDA.n930 3.4105
R14982 GNDA.n951 GNDA.n932 3.4105
R14983 GNDA.n951 GNDA.n929 3.4105
R14984 GNDA.n951 GNDA.n933 3.4105
R14985 GNDA.n951 GNDA.n928 3.4105
R14986 GNDA.n951 GNDA.n934 3.4105
R14987 GNDA.n951 GNDA.n927 3.4105
R14988 GNDA.n951 GNDA.n935 3.4105
R14989 GNDA.n951 GNDA.n926 3.4105
R14990 GNDA.n951 GNDA.n936 3.4105
R14991 GNDA.n951 GNDA.n925 3.4105
R14992 GNDA.n951 GNDA.n937 3.4105
R14993 GNDA.n951 GNDA.n924 3.4105
R14994 GNDA.n951 GNDA.n938 3.4105
R14995 GNDA.n951 GNDA.n923 3.4105
R14996 GNDA.n951 GNDA.n939 3.4105
R14997 GNDA.n951 GNDA.n922 3.4105
R14998 GNDA.n951 GNDA.n940 3.4105
R14999 GNDA.n951 GNDA.n921 3.4105
R15000 GNDA.n951 GNDA.n941 3.4105
R15001 GNDA.n951 GNDA.n920 3.4105
R15002 GNDA.n951 GNDA.n942 3.4105
R15003 GNDA.n951 GNDA.n919 3.4105
R15004 GNDA.n951 GNDA.n943 3.4105
R15005 GNDA.n951 GNDA.n918 3.4105
R15006 GNDA.n951 GNDA.n944 3.4105
R15007 GNDA.n951 GNDA.n917 3.4105
R15008 GNDA.n951 GNDA.n945 3.4105
R15009 GNDA.n1037 GNDA.n951 3.4105
R15010 GNDA.n1035 GNDA.n1022 3.4105
R15011 GNDA.n1022 GNDA.n930 3.4105
R15012 GNDA.n1022 GNDA.n932 3.4105
R15013 GNDA.n1022 GNDA.n929 3.4105
R15014 GNDA.n1022 GNDA.n933 3.4105
R15015 GNDA.n1022 GNDA.n928 3.4105
R15016 GNDA.n1022 GNDA.n934 3.4105
R15017 GNDA.n1022 GNDA.n927 3.4105
R15018 GNDA.n1022 GNDA.n935 3.4105
R15019 GNDA.n1022 GNDA.n926 3.4105
R15020 GNDA.n1022 GNDA.n936 3.4105
R15021 GNDA.n1022 GNDA.n925 3.4105
R15022 GNDA.n1022 GNDA.n937 3.4105
R15023 GNDA.n1022 GNDA.n924 3.4105
R15024 GNDA.n1022 GNDA.n938 3.4105
R15025 GNDA.n1022 GNDA.n923 3.4105
R15026 GNDA.n1022 GNDA.n939 3.4105
R15027 GNDA.n1022 GNDA.n922 3.4105
R15028 GNDA.n1022 GNDA.n940 3.4105
R15029 GNDA.n1022 GNDA.n921 3.4105
R15030 GNDA.n1022 GNDA.n941 3.4105
R15031 GNDA.n1022 GNDA.n920 3.4105
R15032 GNDA.n1022 GNDA.n942 3.4105
R15033 GNDA.n1022 GNDA.n919 3.4105
R15034 GNDA.n1022 GNDA.n943 3.4105
R15035 GNDA.n1022 GNDA.n918 3.4105
R15036 GNDA.n1022 GNDA.n944 3.4105
R15037 GNDA.n1022 GNDA.n917 3.4105
R15038 GNDA.n1022 GNDA.n945 3.4105
R15039 GNDA.n1037 GNDA.n1022 3.4105
R15040 GNDA.n1035 GNDA.n950 3.4105
R15041 GNDA.n950 GNDA.n930 3.4105
R15042 GNDA.n950 GNDA.n932 3.4105
R15043 GNDA.n950 GNDA.n929 3.4105
R15044 GNDA.n950 GNDA.n933 3.4105
R15045 GNDA.n950 GNDA.n928 3.4105
R15046 GNDA.n950 GNDA.n934 3.4105
R15047 GNDA.n950 GNDA.n927 3.4105
R15048 GNDA.n950 GNDA.n935 3.4105
R15049 GNDA.n950 GNDA.n926 3.4105
R15050 GNDA.n950 GNDA.n936 3.4105
R15051 GNDA.n950 GNDA.n925 3.4105
R15052 GNDA.n950 GNDA.n937 3.4105
R15053 GNDA.n950 GNDA.n924 3.4105
R15054 GNDA.n950 GNDA.n938 3.4105
R15055 GNDA.n950 GNDA.n923 3.4105
R15056 GNDA.n950 GNDA.n939 3.4105
R15057 GNDA.n950 GNDA.n922 3.4105
R15058 GNDA.n950 GNDA.n940 3.4105
R15059 GNDA.n950 GNDA.n921 3.4105
R15060 GNDA.n950 GNDA.n941 3.4105
R15061 GNDA.n950 GNDA.n920 3.4105
R15062 GNDA.n950 GNDA.n942 3.4105
R15063 GNDA.n950 GNDA.n919 3.4105
R15064 GNDA.n950 GNDA.n943 3.4105
R15065 GNDA.n950 GNDA.n918 3.4105
R15066 GNDA.n950 GNDA.n944 3.4105
R15067 GNDA.n950 GNDA.n917 3.4105
R15068 GNDA.n950 GNDA.n945 3.4105
R15069 GNDA.n1037 GNDA.n950 3.4105
R15070 GNDA.n1035 GNDA.n1025 3.4105
R15071 GNDA.n1025 GNDA.n930 3.4105
R15072 GNDA.n1025 GNDA.n932 3.4105
R15073 GNDA.n1025 GNDA.n929 3.4105
R15074 GNDA.n1025 GNDA.n933 3.4105
R15075 GNDA.n1025 GNDA.n928 3.4105
R15076 GNDA.n1025 GNDA.n934 3.4105
R15077 GNDA.n1025 GNDA.n927 3.4105
R15078 GNDA.n1025 GNDA.n935 3.4105
R15079 GNDA.n1025 GNDA.n926 3.4105
R15080 GNDA.n1025 GNDA.n936 3.4105
R15081 GNDA.n1025 GNDA.n925 3.4105
R15082 GNDA.n1025 GNDA.n937 3.4105
R15083 GNDA.n1025 GNDA.n924 3.4105
R15084 GNDA.n1025 GNDA.n938 3.4105
R15085 GNDA.n1025 GNDA.n923 3.4105
R15086 GNDA.n1025 GNDA.n939 3.4105
R15087 GNDA.n1025 GNDA.n922 3.4105
R15088 GNDA.n1025 GNDA.n940 3.4105
R15089 GNDA.n1025 GNDA.n921 3.4105
R15090 GNDA.n1025 GNDA.n941 3.4105
R15091 GNDA.n1025 GNDA.n920 3.4105
R15092 GNDA.n1025 GNDA.n942 3.4105
R15093 GNDA.n1025 GNDA.n919 3.4105
R15094 GNDA.n1025 GNDA.n943 3.4105
R15095 GNDA.n1025 GNDA.n918 3.4105
R15096 GNDA.n1025 GNDA.n944 3.4105
R15097 GNDA.n1025 GNDA.n917 3.4105
R15098 GNDA.n1025 GNDA.n945 3.4105
R15099 GNDA.n1037 GNDA.n1025 3.4105
R15100 GNDA.n1035 GNDA.n949 3.4105
R15101 GNDA.n949 GNDA.n930 3.4105
R15102 GNDA.n949 GNDA.n932 3.4105
R15103 GNDA.n949 GNDA.n929 3.4105
R15104 GNDA.n949 GNDA.n933 3.4105
R15105 GNDA.n949 GNDA.n928 3.4105
R15106 GNDA.n949 GNDA.n934 3.4105
R15107 GNDA.n949 GNDA.n927 3.4105
R15108 GNDA.n949 GNDA.n935 3.4105
R15109 GNDA.n949 GNDA.n926 3.4105
R15110 GNDA.n949 GNDA.n936 3.4105
R15111 GNDA.n949 GNDA.n925 3.4105
R15112 GNDA.n949 GNDA.n937 3.4105
R15113 GNDA.n949 GNDA.n924 3.4105
R15114 GNDA.n949 GNDA.n938 3.4105
R15115 GNDA.n949 GNDA.n923 3.4105
R15116 GNDA.n949 GNDA.n939 3.4105
R15117 GNDA.n949 GNDA.n922 3.4105
R15118 GNDA.n949 GNDA.n940 3.4105
R15119 GNDA.n949 GNDA.n921 3.4105
R15120 GNDA.n949 GNDA.n941 3.4105
R15121 GNDA.n949 GNDA.n920 3.4105
R15122 GNDA.n949 GNDA.n942 3.4105
R15123 GNDA.n949 GNDA.n919 3.4105
R15124 GNDA.n949 GNDA.n943 3.4105
R15125 GNDA.n949 GNDA.n918 3.4105
R15126 GNDA.n949 GNDA.n944 3.4105
R15127 GNDA.n949 GNDA.n917 3.4105
R15128 GNDA.n949 GNDA.n945 3.4105
R15129 GNDA.n1037 GNDA.n949 3.4105
R15130 GNDA.n1035 GNDA.n1028 3.4105
R15131 GNDA.n1028 GNDA.n930 3.4105
R15132 GNDA.n1028 GNDA.n932 3.4105
R15133 GNDA.n1028 GNDA.n929 3.4105
R15134 GNDA.n1028 GNDA.n933 3.4105
R15135 GNDA.n1028 GNDA.n928 3.4105
R15136 GNDA.n1028 GNDA.n934 3.4105
R15137 GNDA.n1028 GNDA.n927 3.4105
R15138 GNDA.n1028 GNDA.n935 3.4105
R15139 GNDA.n1028 GNDA.n926 3.4105
R15140 GNDA.n1028 GNDA.n936 3.4105
R15141 GNDA.n1028 GNDA.n925 3.4105
R15142 GNDA.n1028 GNDA.n937 3.4105
R15143 GNDA.n1028 GNDA.n924 3.4105
R15144 GNDA.n1028 GNDA.n938 3.4105
R15145 GNDA.n1028 GNDA.n923 3.4105
R15146 GNDA.n1028 GNDA.n939 3.4105
R15147 GNDA.n1028 GNDA.n922 3.4105
R15148 GNDA.n1028 GNDA.n940 3.4105
R15149 GNDA.n1028 GNDA.n921 3.4105
R15150 GNDA.n1028 GNDA.n941 3.4105
R15151 GNDA.n1028 GNDA.n920 3.4105
R15152 GNDA.n1028 GNDA.n942 3.4105
R15153 GNDA.n1028 GNDA.n919 3.4105
R15154 GNDA.n1028 GNDA.n943 3.4105
R15155 GNDA.n1028 GNDA.n918 3.4105
R15156 GNDA.n1028 GNDA.n944 3.4105
R15157 GNDA.n1028 GNDA.n917 3.4105
R15158 GNDA.n1028 GNDA.n945 3.4105
R15159 GNDA.n1037 GNDA.n1028 3.4105
R15160 GNDA.n1035 GNDA.n948 3.4105
R15161 GNDA.n948 GNDA.n930 3.4105
R15162 GNDA.n948 GNDA.n932 3.4105
R15163 GNDA.n948 GNDA.n929 3.4105
R15164 GNDA.n948 GNDA.n933 3.4105
R15165 GNDA.n948 GNDA.n928 3.4105
R15166 GNDA.n948 GNDA.n934 3.4105
R15167 GNDA.n948 GNDA.n927 3.4105
R15168 GNDA.n948 GNDA.n935 3.4105
R15169 GNDA.n948 GNDA.n926 3.4105
R15170 GNDA.n948 GNDA.n936 3.4105
R15171 GNDA.n948 GNDA.n925 3.4105
R15172 GNDA.n948 GNDA.n937 3.4105
R15173 GNDA.n948 GNDA.n924 3.4105
R15174 GNDA.n948 GNDA.n938 3.4105
R15175 GNDA.n948 GNDA.n923 3.4105
R15176 GNDA.n948 GNDA.n939 3.4105
R15177 GNDA.n948 GNDA.n922 3.4105
R15178 GNDA.n948 GNDA.n940 3.4105
R15179 GNDA.n948 GNDA.n921 3.4105
R15180 GNDA.n948 GNDA.n941 3.4105
R15181 GNDA.n948 GNDA.n920 3.4105
R15182 GNDA.n948 GNDA.n942 3.4105
R15183 GNDA.n948 GNDA.n919 3.4105
R15184 GNDA.n948 GNDA.n943 3.4105
R15185 GNDA.n948 GNDA.n918 3.4105
R15186 GNDA.n948 GNDA.n944 3.4105
R15187 GNDA.n948 GNDA.n917 3.4105
R15188 GNDA.n948 GNDA.n945 3.4105
R15189 GNDA.n1037 GNDA.n948 3.4105
R15190 GNDA.n1035 GNDA.n1031 3.4105
R15191 GNDA.n1031 GNDA.n930 3.4105
R15192 GNDA.n1031 GNDA.n932 3.4105
R15193 GNDA.n1031 GNDA.n929 3.4105
R15194 GNDA.n1031 GNDA.n933 3.4105
R15195 GNDA.n1031 GNDA.n928 3.4105
R15196 GNDA.n1031 GNDA.n934 3.4105
R15197 GNDA.n1031 GNDA.n927 3.4105
R15198 GNDA.n1031 GNDA.n935 3.4105
R15199 GNDA.n1031 GNDA.n926 3.4105
R15200 GNDA.n1031 GNDA.n936 3.4105
R15201 GNDA.n1031 GNDA.n925 3.4105
R15202 GNDA.n1031 GNDA.n937 3.4105
R15203 GNDA.n1031 GNDA.n924 3.4105
R15204 GNDA.n1031 GNDA.n938 3.4105
R15205 GNDA.n1031 GNDA.n923 3.4105
R15206 GNDA.n1031 GNDA.n939 3.4105
R15207 GNDA.n1031 GNDA.n922 3.4105
R15208 GNDA.n1031 GNDA.n940 3.4105
R15209 GNDA.n1031 GNDA.n921 3.4105
R15210 GNDA.n1031 GNDA.n941 3.4105
R15211 GNDA.n1031 GNDA.n920 3.4105
R15212 GNDA.n1031 GNDA.n942 3.4105
R15213 GNDA.n1031 GNDA.n919 3.4105
R15214 GNDA.n1031 GNDA.n943 3.4105
R15215 GNDA.n1031 GNDA.n918 3.4105
R15216 GNDA.n1031 GNDA.n944 3.4105
R15217 GNDA.n1031 GNDA.n917 3.4105
R15218 GNDA.n1031 GNDA.n945 3.4105
R15219 GNDA.n1037 GNDA.n1031 3.4105
R15220 GNDA.n1035 GNDA.n947 3.4105
R15221 GNDA.n947 GNDA.n930 3.4105
R15222 GNDA.n947 GNDA.n932 3.4105
R15223 GNDA.n947 GNDA.n929 3.4105
R15224 GNDA.n947 GNDA.n933 3.4105
R15225 GNDA.n947 GNDA.n928 3.4105
R15226 GNDA.n947 GNDA.n934 3.4105
R15227 GNDA.n947 GNDA.n927 3.4105
R15228 GNDA.n947 GNDA.n935 3.4105
R15229 GNDA.n947 GNDA.n926 3.4105
R15230 GNDA.n947 GNDA.n936 3.4105
R15231 GNDA.n947 GNDA.n925 3.4105
R15232 GNDA.n947 GNDA.n937 3.4105
R15233 GNDA.n947 GNDA.n924 3.4105
R15234 GNDA.n947 GNDA.n938 3.4105
R15235 GNDA.n947 GNDA.n923 3.4105
R15236 GNDA.n947 GNDA.n939 3.4105
R15237 GNDA.n947 GNDA.n922 3.4105
R15238 GNDA.n947 GNDA.n940 3.4105
R15239 GNDA.n947 GNDA.n921 3.4105
R15240 GNDA.n947 GNDA.n941 3.4105
R15241 GNDA.n947 GNDA.n920 3.4105
R15242 GNDA.n947 GNDA.n942 3.4105
R15243 GNDA.n947 GNDA.n919 3.4105
R15244 GNDA.n947 GNDA.n943 3.4105
R15245 GNDA.n947 GNDA.n918 3.4105
R15246 GNDA.n947 GNDA.n944 3.4105
R15247 GNDA.n947 GNDA.n917 3.4105
R15248 GNDA.n947 GNDA.n945 3.4105
R15249 GNDA.n1037 GNDA.n947 3.4105
R15250 GNDA.n1036 GNDA.n1035 3.4105
R15251 GNDA.n1036 GNDA.n930 3.4105
R15252 GNDA.n1036 GNDA.n932 3.4105
R15253 GNDA.n1036 GNDA.n929 3.4105
R15254 GNDA.n1036 GNDA.n933 3.4105
R15255 GNDA.n1036 GNDA.n928 3.4105
R15256 GNDA.n1036 GNDA.n934 3.4105
R15257 GNDA.n1036 GNDA.n927 3.4105
R15258 GNDA.n1036 GNDA.n935 3.4105
R15259 GNDA.n1036 GNDA.n926 3.4105
R15260 GNDA.n1036 GNDA.n936 3.4105
R15261 GNDA.n1036 GNDA.n925 3.4105
R15262 GNDA.n1036 GNDA.n937 3.4105
R15263 GNDA.n1036 GNDA.n924 3.4105
R15264 GNDA.n1036 GNDA.n938 3.4105
R15265 GNDA.n1036 GNDA.n923 3.4105
R15266 GNDA.n1036 GNDA.n939 3.4105
R15267 GNDA.n1036 GNDA.n922 3.4105
R15268 GNDA.n1036 GNDA.n940 3.4105
R15269 GNDA.n1036 GNDA.n921 3.4105
R15270 GNDA.n1036 GNDA.n941 3.4105
R15271 GNDA.n1036 GNDA.n920 3.4105
R15272 GNDA.n1036 GNDA.n942 3.4105
R15273 GNDA.n1036 GNDA.n919 3.4105
R15274 GNDA.n1036 GNDA.n943 3.4105
R15275 GNDA.n1036 GNDA.n918 3.4105
R15276 GNDA.n1036 GNDA.n944 3.4105
R15277 GNDA.n1036 GNDA.n917 3.4105
R15278 GNDA.n1036 GNDA.n945 3.4105
R15279 GNDA.n1037 GNDA.n1036 3.4105
R15280 GNDA.n1035 GNDA.n946 3.4105
R15281 GNDA.n946 GNDA.n930 3.4105
R15282 GNDA.n946 GNDA.n932 3.4105
R15283 GNDA.n946 GNDA.n929 3.4105
R15284 GNDA.n946 GNDA.n933 3.4105
R15285 GNDA.n946 GNDA.n928 3.4105
R15286 GNDA.n946 GNDA.n934 3.4105
R15287 GNDA.n946 GNDA.n927 3.4105
R15288 GNDA.n946 GNDA.n935 3.4105
R15289 GNDA.n946 GNDA.n926 3.4105
R15290 GNDA.n946 GNDA.n936 3.4105
R15291 GNDA.n946 GNDA.n925 3.4105
R15292 GNDA.n946 GNDA.n937 3.4105
R15293 GNDA.n946 GNDA.n924 3.4105
R15294 GNDA.n946 GNDA.n938 3.4105
R15295 GNDA.n946 GNDA.n923 3.4105
R15296 GNDA.n946 GNDA.n939 3.4105
R15297 GNDA.n946 GNDA.n922 3.4105
R15298 GNDA.n946 GNDA.n940 3.4105
R15299 GNDA.n946 GNDA.n921 3.4105
R15300 GNDA.n946 GNDA.n941 3.4105
R15301 GNDA.n946 GNDA.n920 3.4105
R15302 GNDA.n946 GNDA.n942 3.4105
R15303 GNDA.n946 GNDA.n919 3.4105
R15304 GNDA.n946 GNDA.n943 3.4105
R15305 GNDA.n946 GNDA.n918 3.4105
R15306 GNDA.n946 GNDA.n944 3.4105
R15307 GNDA.n946 GNDA.n917 3.4105
R15308 GNDA.n946 GNDA.n945 3.4105
R15309 GNDA.n1037 GNDA.n946 3.4105
R15310 GNDA.n1038 GNDA.n930 3.4105
R15311 GNDA.n1038 GNDA.n932 3.4105
R15312 GNDA.n1038 GNDA.n929 3.4105
R15313 GNDA.n1038 GNDA.n933 3.4105
R15314 GNDA.n1038 GNDA.n928 3.4105
R15315 GNDA.n1038 GNDA.n934 3.4105
R15316 GNDA.n1038 GNDA.n927 3.4105
R15317 GNDA.n1038 GNDA.n935 3.4105
R15318 GNDA.n1038 GNDA.n926 3.4105
R15319 GNDA.n1038 GNDA.n936 3.4105
R15320 GNDA.n1038 GNDA.n925 3.4105
R15321 GNDA.n1038 GNDA.n937 3.4105
R15322 GNDA.n1038 GNDA.n924 3.4105
R15323 GNDA.n1038 GNDA.n938 3.4105
R15324 GNDA.n1038 GNDA.n923 3.4105
R15325 GNDA.n1038 GNDA.n939 3.4105
R15326 GNDA.n1038 GNDA.n922 3.4105
R15327 GNDA.n1038 GNDA.n940 3.4105
R15328 GNDA.n1038 GNDA.n921 3.4105
R15329 GNDA.n1038 GNDA.n941 3.4105
R15330 GNDA.n1038 GNDA.n920 3.4105
R15331 GNDA.n1038 GNDA.n942 3.4105
R15332 GNDA.n1038 GNDA.n919 3.4105
R15333 GNDA.n1038 GNDA.n943 3.4105
R15334 GNDA.n1038 GNDA.n918 3.4105
R15335 GNDA.n1038 GNDA.n944 3.4105
R15336 GNDA.n1038 GNDA.n917 3.4105
R15337 GNDA.n1038 GNDA.n945 3.4105
R15338 GNDA.n1038 GNDA.n1037 3.4105
R15339 GNDA.n1166 GNDA.n1059 3.4105
R15340 GNDA.n1162 GNDA.n1059 3.4105
R15341 GNDA.n1164 GNDA.n1059 3.4105
R15342 GNDA.n1163 GNDA.n1162 3.4105
R15343 GNDA.n1164 GNDA.n1163 3.4105
R15344 GNDA.n1166 GNDA.n809 3.4105
R15345 GNDA.n1090 GNDA.n809 3.4105
R15346 GNDA.n1088 GNDA.n809 3.4105
R15347 GNDA.n1092 GNDA.n809 3.4105
R15348 GNDA.n1087 GNDA.n809 3.4105
R15349 GNDA.n1094 GNDA.n809 3.4105
R15350 GNDA.n1086 GNDA.n809 3.4105
R15351 GNDA.n1096 GNDA.n809 3.4105
R15352 GNDA.n1085 GNDA.n809 3.4105
R15353 GNDA.n1098 GNDA.n809 3.4105
R15354 GNDA.n1084 GNDA.n809 3.4105
R15355 GNDA.n1100 GNDA.n809 3.4105
R15356 GNDA.n1083 GNDA.n809 3.4105
R15357 GNDA.n1102 GNDA.n809 3.4105
R15358 GNDA.n1082 GNDA.n809 3.4105
R15359 GNDA.n1104 GNDA.n809 3.4105
R15360 GNDA.n1081 GNDA.n809 3.4105
R15361 GNDA.n1106 GNDA.n809 3.4105
R15362 GNDA.n1080 GNDA.n809 3.4105
R15363 GNDA.n1108 GNDA.n809 3.4105
R15364 GNDA.n1079 GNDA.n809 3.4105
R15365 GNDA.n1110 GNDA.n809 3.4105
R15366 GNDA.n1078 GNDA.n809 3.4105
R15367 GNDA.n1112 GNDA.n809 3.4105
R15368 GNDA.n1077 GNDA.n809 3.4105
R15369 GNDA.n1114 GNDA.n809 3.4105
R15370 GNDA.n1076 GNDA.n809 3.4105
R15371 GNDA.n1115 GNDA.n809 3.4105
R15372 GNDA.n1162 GNDA.n809 3.4105
R15373 GNDA.n1164 GNDA.n809 3.4105
R15374 GNDA.n1166 GNDA.n1060 3.4105
R15375 GNDA.n1090 GNDA.n1060 3.4105
R15376 GNDA.n1088 GNDA.n1060 3.4105
R15377 GNDA.n1092 GNDA.n1060 3.4105
R15378 GNDA.n1087 GNDA.n1060 3.4105
R15379 GNDA.n1094 GNDA.n1060 3.4105
R15380 GNDA.n1086 GNDA.n1060 3.4105
R15381 GNDA.n1096 GNDA.n1060 3.4105
R15382 GNDA.n1085 GNDA.n1060 3.4105
R15383 GNDA.n1098 GNDA.n1060 3.4105
R15384 GNDA.n1084 GNDA.n1060 3.4105
R15385 GNDA.n1100 GNDA.n1060 3.4105
R15386 GNDA.n1083 GNDA.n1060 3.4105
R15387 GNDA.n1102 GNDA.n1060 3.4105
R15388 GNDA.n1082 GNDA.n1060 3.4105
R15389 GNDA.n1104 GNDA.n1060 3.4105
R15390 GNDA.n1081 GNDA.n1060 3.4105
R15391 GNDA.n1106 GNDA.n1060 3.4105
R15392 GNDA.n1080 GNDA.n1060 3.4105
R15393 GNDA.n1108 GNDA.n1060 3.4105
R15394 GNDA.n1079 GNDA.n1060 3.4105
R15395 GNDA.n1110 GNDA.n1060 3.4105
R15396 GNDA.n1078 GNDA.n1060 3.4105
R15397 GNDA.n1112 GNDA.n1060 3.4105
R15398 GNDA.n1077 GNDA.n1060 3.4105
R15399 GNDA.n1114 GNDA.n1060 3.4105
R15400 GNDA.n1076 GNDA.n1060 3.4105
R15401 GNDA.n1115 GNDA.n1060 3.4105
R15402 GNDA.n1162 GNDA.n1060 3.4105
R15403 GNDA.n1164 GNDA.n1060 3.4105
R15404 GNDA.n1166 GNDA.n808 3.4105
R15405 GNDA.n1090 GNDA.n808 3.4105
R15406 GNDA.n1088 GNDA.n808 3.4105
R15407 GNDA.n1092 GNDA.n808 3.4105
R15408 GNDA.n1087 GNDA.n808 3.4105
R15409 GNDA.n1094 GNDA.n808 3.4105
R15410 GNDA.n1086 GNDA.n808 3.4105
R15411 GNDA.n1096 GNDA.n808 3.4105
R15412 GNDA.n1085 GNDA.n808 3.4105
R15413 GNDA.n1098 GNDA.n808 3.4105
R15414 GNDA.n1084 GNDA.n808 3.4105
R15415 GNDA.n1100 GNDA.n808 3.4105
R15416 GNDA.n1083 GNDA.n808 3.4105
R15417 GNDA.n1102 GNDA.n808 3.4105
R15418 GNDA.n1082 GNDA.n808 3.4105
R15419 GNDA.n1104 GNDA.n808 3.4105
R15420 GNDA.n1081 GNDA.n808 3.4105
R15421 GNDA.n1106 GNDA.n808 3.4105
R15422 GNDA.n1080 GNDA.n808 3.4105
R15423 GNDA.n1108 GNDA.n808 3.4105
R15424 GNDA.n1079 GNDA.n808 3.4105
R15425 GNDA.n1110 GNDA.n808 3.4105
R15426 GNDA.n1078 GNDA.n808 3.4105
R15427 GNDA.n1112 GNDA.n808 3.4105
R15428 GNDA.n1077 GNDA.n808 3.4105
R15429 GNDA.n1114 GNDA.n808 3.4105
R15430 GNDA.n1076 GNDA.n808 3.4105
R15431 GNDA.n1115 GNDA.n808 3.4105
R15432 GNDA.n1162 GNDA.n808 3.4105
R15433 GNDA.n1164 GNDA.n808 3.4105
R15434 GNDA.n1166 GNDA.n1061 3.4105
R15435 GNDA.n1090 GNDA.n1061 3.4105
R15436 GNDA.n1088 GNDA.n1061 3.4105
R15437 GNDA.n1092 GNDA.n1061 3.4105
R15438 GNDA.n1087 GNDA.n1061 3.4105
R15439 GNDA.n1094 GNDA.n1061 3.4105
R15440 GNDA.n1086 GNDA.n1061 3.4105
R15441 GNDA.n1096 GNDA.n1061 3.4105
R15442 GNDA.n1085 GNDA.n1061 3.4105
R15443 GNDA.n1098 GNDA.n1061 3.4105
R15444 GNDA.n1084 GNDA.n1061 3.4105
R15445 GNDA.n1100 GNDA.n1061 3.4105
R15446 GNDA.n1083 GNDA.n1061 3.4105
R15447 GNDA.n1102 GNDA.n1061 3.4105
R15448 GNDA.n1082 GNDA.n1061 3.4105
R15449 GNDA.n1104 GNDA.n1061 3.4105
R15450 GNDA.n1081 GNDA.n1061 3.4105
R15451 GNDA.n1106 GNDA.n1061 3.4105
R15452 GNDA.n1080 GNDA.n1061 3.4105
R15453 GNDA.n1108 GNDA.n1061 3.4105
R15454 GNDA.n1079 GNDA.n1061 3.4105
R15455 GNDA.n1110 GNDA.n1061 3.4105
R15456 GNDA.n1078 GNDA.n1061 3.4105
R15457 GNDA.n1112 GNDA.n1061 3.4105
R15458 GNDA.n1077 GNDA.n1061 3.4105
R15459 GNDA.n1114 GNDA.n1061 3.4105
R15460 GNDA.n1076 GNDA.n1061 3.4105
R15461 GNDA.n1115 GNDA.n1061 3.4105
R15462 GNDA.n1162 GNDA.n1061 3.4105
R15463 GNDA.n1164 GNDA.n1061 3.4105
R15464 GNDA.n1166 GNDA.n807 3.4105
R15465 GNDA.n1090 GNDA.n807 3.4105
R15466 GNDA.n1088 GNDA.n807 3.4105
R15467 GNDA.n1092 GNDA.n807 3.4105
R15468 GNDA.n1087 GNDA.n807 3.4105
R15469 GNDA.n1094 GNDA.n807 3.4105
R15470 GNDA.n1086 GNDA.n807 3.4105
R15471 GNDA.n1096 GNDA.n807 3.4105
R15472 GNDA.n1085 GNDA.n807 3.4105
R15473 GNDA.n1098 GNDA.n807 3.4105
R15474 GNDA.n1084 GNDA.n807 3.4105
R15475 GNDA.n1100 GNDA.n807 3.4105
R15476 GNDA.n1083 GNDA.n807 3.4105
R15477 GNDA.n1102 GNDA.n807 3.4105
R15478 GNDA.n1082 GNDA.n807 3.4105
R15479 GNDA.n1104 GNDA.n807 3.4105
R15480 GNDA.n1081 GNDA.n807 3.4105
R15481 GNDA.n1106 GNDA.n807 3.4105
R15482 GNDA.n1080 GNDA.n807 3.4105
R15483 GNDA.n1108 GNDA.n807 3.4105
R15484 GNDA.n1079 GNDA.n807 3.4105
R15485 GNDA.n1110 GNDA.n807 3.4105
R15486 GNDA.n1078 GNDA.n807 3.4105
R15487 GNDA.n1112 GNDA.n807 3.4105
R15488 GNDA.n1077 GNDA.n807 3.4105
R15489 GNDA.n1114 GNDA.n807 3.4105
R15490 GNDA.n1076 GNDA.n807 3.4105
R15491 GNDA.n1115 GNDA.n807 3.4105
R15492 GNDA.n1162 GNDA.n807 3.4105
R15493 GNDA.n1164 GNDA.n807 3.4105
R15494 GNDA.n1166 GNDA.n1062 3.4105
R15495 GNDA.n1090 GNDA.n1062 3.4105
R15496 GNDA.n1088 GNDA.n1062 3.4105
R15497 GNDA.n1092 GNDA.n1062 3.4105
R15498 GNDA.n1087 GNDA.n1062 3.4105
R15499 GNDA.n1094 GNDA.n1062 3.4105
R15500 GNDA.n1086 GNDA.n1062 3.4105
R15501 GNDA.n1096 GNDA.n1062 3.4105
R15502 GNDA.n1085 GNDA.n1062 3.4105
R15503 GNDA.n1098 GNDA.n1062 3.4105
R15504 GNDA.n1084 GNDA.n1062 3.4105
R15505 GNDA.n1100 GNDA.n1062 3.4105
R15506 GNDA.n1083 GNDA.n1062 3.4105
R15507 GNDA.n1102 GNDA.n1062 3.4105
R15508 GNDA.n1082 GNDA.n1062 3.4105
R15509 GNDA.n1104 GNDA.n1062 3.4105
R15510 GNDA.n1081 GNDA.n1062 3.4105
R15511 GNDA.n1106 GNDA.n1062 3.4105
R15512 GNDA.n1080 GNDA.n1062 3.4105
R15513 GNDA.n1108 GNDA.n1062 3.4105
R15514 GNDA.n1079 GNDA.n1062 3.4105
R15515 GNDA.n1110 GNDA.n1062 3.4105
R15516 GNDA.n1078 GNDA.n1062 3.4105
R15517 GNDA.n1112 GNDA.n1062 3.4105
R15518 GNDA.n1077 GNDA.n1062 3.4105
R15519 GNDA.n1114 GNDA.n1062 3.4105
R15520 GNDA.n1076 GNDA.n1062 3.4105
R15521 GNDA.n1115 GNDA.n1062 3.4105
R15522 GNDA.n1162 GNDA.n1062 3.4105
R15523 GNDA.n1164 GNDA.n1062 3.4105
R15524 GNDA.n1166 GNDA.n806 3.4105
R15525 GNDA.n1090 GNDA.n806 3.4105
R15526 GNDA.n1088 GNDA.n806 3.4105
R15527 GNDA.n1092 GNDA.n806 3.4105
R15528 GNDA.n1087 GNDA.n806 3.4105
R15529 GNDA.n1094 GNDA.n806 3.4105
R15530 GNDA.n1086 GNDA.n806 3.4105
R15531 GNDA.n1096 GNDA.n806 3.4105
R15532 GNDA.n1085 GNDA.n806 3.4105
R15533 GNDA.n1098 GNDA.n806 3.4105
R15534 GNDA.n1084 GNDA.n806 3.4105
R15535 GNDA.n1100 GNDA.n806 3.4105
R15536 GNDA.n1083 GNDA.n806 3.4105
R15537 GNDA.n1102 GNDA.n806 3.4105
R15538 GNDA.n1082 GNDA.n806 3.4105
R15539 GNDA.n1104 GNDA.n806 3.4105
R15540 GNDA.n1081 GNDA.n806 3.4105
R15541 GNDA.n1106 GNDA.n806 3.4105
R15542 GNDA.n1080 GNDA.n806 3.4105
R15543 GNDA.n1108 GNDA.n806 3.4105
R15544 GNDA.n1079 GNDA.n806 3.4105
R15545 GNDA.n1110 GNDA.n806 3.4105
R15546 GNDA.n1078 GNDA.n806 3.4105
R15547 GNDA.n1112 GNDA.n806 3.4105
R15548 GNDA.n1077 GNDA.n806 3.4105
R15549 GNDA.n1114 GNDA.n806 3.4105
R15550 GNDA.n1076 GNDA.n806 3.4105
R15551 GNDA.n1115 GNDA.n806 3.4105
R15552 GNDA.n1162 GNDA.n806 3.4105
R15553 GNDA.n1164 GNDA.n806 3.4105
R15554 GNDA.n1166 GNDA.n1063 3.4105
R15555 GNDA.n1090 GNDA.n1063 3.4105
R15556 GNDA.n1088 GNDA.n1063 3.4105
R15557 GNDA.n1092 GNDA.n1063 3.4105
R15558 GNDA.n1087 GNDA.n1063 3.4105
R15559 GNDA.n1094 GNDA.n1063 3.4105
R15560 GNDA.n1086 GNDA.n1063 3.4105
R15561 GNDA.n1096 GNDA.n1063 3.4105
R15562 GNDA.n1085 GNDA.n1063 3.4105
R15563 GNDA.n1098 GNDA.n1063 3.4105
R15564 GNDA.n1084 GNDA.n1063 3.4105
R15565 GNDA.n1100 GNDA.n1063 3.4105
R15566 GNDA.n1083 GNDA.n1063 3.4105
R15567 GNDA.n1102 GNDA.n1063 3.4105
R15568 GNDA.n1082 GNDA.n1063 3.4105
R15569 GNDA.n1104 GNDA.n1063 3.4105
R15570 GNDA.n1081 GNDA.n1063 3.4105
R15571 GNDA.n1106 GNDA.n1063 3.4105
R15572 GNDA.n1080 GNDA.n1063 3.4105
R15573 GNDA.n1108 GNDA.n1063 3.4105
R15574 GNDA.n1079 GNDA.n1063 3.4105
R15575 GNDA.n1110 GNDA.n1063 3.4105
R15576 GNDA.n1078 GNDA.n1063 3.4105
R15577 GNDA.n1112 GNDA.n1063 3.4105
R15578 GNDA.n1077 GNDA.n1063 3.4105
R15579 GNDA.n1114 GNDA.n1063 3.4105
R15580 GNDA.n1076 GNDA.n1063 3.4105
R15581 GNDA.n1115 GNDA.n1063 3.4105
R15582 GNDA.n1162 GNDA.n1063 3.4105
R15583 GNDA.n1164 GNDA.n1063 3.4105
R15584 GNDA.n1166 GNDA.n805 3.4105
R15585 GNDA.n1090 GNDA.n805 3.4105
R15586 GNDA.n1088 GNDA.n805 3.4105
R15587 GNDA.n1092 GNDA.n805 3.4105
R15588 GNDA.n1087 GNDA.n805 3.4105
R15589 GNDA.n1094 GNDA.n805 3.4105
R15590 GNDA.n1086 GNDA.n805 3.4105
R15591 GNDA.n1096 GNDA.n805 3.4105
R15592 GNDA.n1085 GNDA.n805 3.4105
R15593 GNDA.n1098 GNDA.n805 3.4105
R15594 GNDA.n1084 GNDA.n805 3.4105
R15595 GNDA.n1100 GNDA.n805 3.4105
R15596 GNDA.n1083 GNDA.n805 3.4105
R15597 GNDA.n1102 GNDA.n805 3.4105
R15598 GNDA.n1082 GNDA.n805 3.4105
R15599 GNDA.n1104 GNDA.n805 3.4105
R15600 GNDA.n1081 GNDA.n805 3.4105
R15601 GNDA.n1106 GNDA.n805 3.4105
R15602 GNDA.n1080 GNDA.n805 3.4105
R15603 GNDA.n1108 GNDA.n805 3.4105
R15604 GNDA.n1079 GNDA.n805 3.4105
R15605 GNDA.n1110 GNDA.n805 3.4105
R15606 GNDA.n1078 GNDA.n805 3.4105
R15607 GNDA.n1112 GNDA.n805 3.4105
R15608 GNDA.n1077 GNDA.n805 3.4105
R15609 GNDA.n1114 GNDA.n805 3.4105
R15610 GNDA.n1076 GNDA.n805 3.4105
R15611 GNDA.n1115 GNDA.n805 3.4105
R15612 GNDA.n1162 GNDA.n805 3.4105
R15613 GNDA.n1164 GNDA.n805 3.4105
R15614 GNDA.n1166 GNDA.n1064 3.4105
R15615 GNDA.n1090 GNDA.n1064 3.4105
R15616 GNDA.n1088 GNDA.n1064 3.4105
R15617 GNDA.n1092 GNDA.n1064 3.4105
R15618 GNDA.n1087 GNDA.n1064 3.4105
R15619 GNDA.n1094 GNDA.n1064 3.4105
R15620 GNDA.n1086 GNDA.n1064 3.4105
R15621 GNDA.n1096 GNDA.n1064 3.4105
R15622 GNDA.n1085 GNDA.n1064 3.4105
R15623 GNDA.n1098 GNDA.n1064 3.4105
R15624 GNDA.n1084 GNDA.n1064 3.4105
R15625 GNDA.n1100 GNDA.n1064 3.4105
R15626 GNDA.n1083 GNDA.n1064 3.4105
R15627 GNDA.n1102 GNDA.n1064 3.4105
R15628 GNDA.n1082 GNDA.n1064 3.4105
R15629 GNDA.n1104 GNDA.n1064 3.4105
R15630 GNDA.n1081 GNDA.n1064 3.4105
R15631 GNDA.n1106 GNDA.n1064 3.4105
R15632 GNDA.n1080 GNDA.n1064 3.4105
R15633 GNDA.n1108 GNDA.n1064 3.4105
R15634 GNDA.n1079 GNDA.n1064 3.4105
R15635 GNDA.n1110 GNDA.n1064 3.4105
R15636 GNDA.n1078 GNDA.n1064 3.4105
R15637 GNDA.n1112 GNDA.n1064 3.4105
R15638 GNDA.n1077 GNDA.n1064 3.4105
R15639 GNDA.n1114 GNDA.n1064 3.4105
R15640 GNDA.n1076 GNDA.n1064 3.4105
R15641 GNDA.n1115 GNDA.n1064 3.4105
R15642 GNDA.n1162 GNDA.n1064 3.4105
R15643 GNDA.n1164 GNDA.n1064 3.4105
R15644 GNDA.n1166 GNDA.n804 3.4105
R15645 GNDA.n1090 GNDA.n804 3.4105
R15646 GNDA.n1088 GNDA.n804 3.4105
R15647 GNDA.n1092 GNDA.n804 3.4105
R15648 GNDA.n1087 GNDA.n804 3.4105
R15649 GNDA.n1094 GNDA.n804 3.4105
R15650 GNDA.n1086 GNDA.n804 3.4105
R15651 GNDA.n1096 GNDA.n804 3.4105
R15652 GNDA.n1085 GNDA.n804 3.4105
R15653 GNDA.n1098 GNDA.n804 3.4105
R15654 GNDA.n1084 GNDA.n804 3.4105
R15655 GNDA.n1100 GNDA.n804 3.4105
R15656 GNDA.n1083 GNDA.n804 3.4105
R15657 GNDA.n1102 GNDA.n804 3.4105
R15658 GNDA.n1082 GNDA.n804 3.4105
R15659 GNDA.n1104 GNDA.n804 3.4105
R15660 GNDA.n1081 GNDA.n804 3.4105
R15661 GNDA.n1106 GNDA.n804 3.4105
R15662 GNDA.n1080 GNDA.n804 3.4105
R15663 GNDA.n1108 GNDA.n804 3.4105
R15664 GNDA.n1079 GNDA.n804 3.4105
R15665 GNDA.n1110 GNDA.n804 3.4105
R15666 GNDA.n1078 GNDA.n804 3.4105
R15667 GNDA.n1112 GNDA.n804 3.4105
R15668 GNDA.n1077 GNDA.n804 3.4105
R15669 GNDA.n1114 GNDA.n804 3.4105
R15670 GNDA.n1076 GNDA.n804 3.4105
R15671 GNDA.n1115 GNDA.n804 3.4105
R15672 GNDA.n1162 GNDA.n804 3.4105
R15673 GNDA.n1164 GNDA.n804 3.4105
R15674 GNDA.n1166 GNDA.n1065 3.4105
R15675 GNDA.n1090 GNDA.n1065 3.4105
R15676 GNDA.n1088 GNDA.n1065 3.4105
R15677 GNDA.n1092 GNDA.n1065 3.4105
R15678 GNDA.n1087 GNDA.n1065 3.4105
R15679 GNDA.n1094 GNDA.n1065 3.4105
R15680 GNDA.n1086 GNDA.n1065 3.4105
R15681 GNDA.n1096 GNDA.n1065 3.4105
R15682 GNDA.n1085 GNDA.n1065 3.4105
R15683 GNDA.n1098 GNDA.n1065 3.4105
R15684 GNDA.n1084 GNDA.n1065 3.4105
R15685 GNDA.n1100 GNDA.n1065 3.4105
R15686 GNDA.n1083 GNDA.n1065 3.4105
R15687 GNDA.n1102 GNDA.n1065 3.4105
R15688 GNDA.n1082 GNDA.n1065 3.4105
R15689 GNDA.n1104 GNDA.n1065 3.4105
R15690 GNDA.n1081 GNDA.n1065 3.4105
R15691 GNDA.n1106 GNDA.n1065 3.4105
R15692 GNDA.n1080 GNDA.n1065 3.4105
R15693 GNDA.n1108 GNDA.n1065 3.4105
R15694 GNDA.n1079 GNDA.n1065 3.4105
R15695 GNDA.n1110 GNDA.n1065 3.4105
R15696 GNDA.n1078 GNDA.n1065 3.4105
R15697 GNDA.n1112 GNDA.n1065 3.4105
R15698 GNDA.n1077 GNDA.n1065 3.4105
R15699 GNDA.n1114 GNDA.n1065 3.4105
R15700 GNDA.n1076 GNDA.n1065 3.4105
R15701 GNDA.n1115 GNDA.n1065 3.4105
R15702 GNDA.n1162 GNDA.n1065 3.4105
R15703 GNDA.n1164 GNDA.n1065 3.4105
R15704 GNDA.n1166 GNDA.n803 3.4105
R15705 GNDA.n1090 GNDA.n803 3.4105
R15706 GNDA.n1088 GNDA.n803 3.4105
R15707 GNDA.n1092 GNDA.n803 3.4105
R15708 GNDA.n1087 GNDA.n803 3.4105
R15709 GNDA.n1094 GNDA.n803 3.4105
R15710 GNDA.n1086 GNDA.n803 3.4105
R15711 GNDA.n1096 GNDA.n803 3.4105
R15712 GNDA.n1085 GNDA.n803 3.4105
R15713 GNDA.n1098 GNDA.n803 3.4105
R15714 GNDA.n1084 GNDA.n803 3.4105
R15715 GNDA.n1100 GNDA.n803 3.4105
R15716 GNDA.n1083 GNDA.n803 3.4105
R15717 GNDA.n1102 GNDA.n803 3.4105
R15718 GNDA.n1082 GNDA.n803 3.4105
R15719 GNDA.n1104 GNDA.n803 3.4105
R15720 GNDA.n1081 GNDA.n803 3.4105
R15721 GNDA.n1106 GNDA.n803 3.4105
R15722 GNDA.n1080 GNDA.n803 3.4105
R15723 GNDA.n1108 GNDA.n803 3.4105
R15724 GNDA.n1079 GNDA.n803 3.4105
R15725 GNDA.n1110 GNDA.n803 3.4105
R15726 GNDA.n1078 GNDA.n803 3.4105
R15727 GNDA.n1112 GNDA.n803 3.4105
R15728 GNDA.n1077 GNDA.n803 3.4105
R15729 GNDA.n1114 GNDA.n803 3.4105
R15730 GNDA.n1076 GNDA.n803 3.4105
R15731 GNDA.n1115 GNDA.n803 3.4105
R15732 GNDA.n1162 GNDA.n803 3.4105
R15733 GNDA.n1164 GNDA.n803 3.4105
R15734 GNDA.n1166 GNDA.n1066 3.4105
R15735 GNDA.n1090 GNDA.n1066 3.4105
R15736 GNDA.n1088 GNDA.n1066 3.4105
R15737 GNDA.n1092 GNDA.n1066 3.4105
R15738 GNDA.n1087 GNDA.n1066 3.4105
R15739 GNDA.n1094 GNDA.n1066 3.4105
R15740 GNDA.n1086 GNDA.n1066 3.4105
R15741 GNDA.n1096 GNDA.n1066 3.4105
R15742 GNDA.n1085 GNDA.n1066 3.4105
R15743 GNDA.n1098 GNDA.n1066 3.4105
R15744 GNDA.n1084 GNDA.n1066 3.4105
R15745 GNDA.n1100 GNDA.n1066 3.4105
R15746 GNDA.n1083 GNDA.n1066 3.4105
R15747 GNDA.n1102 GNDA.n1066 3.4105
R15748 GNDA.n1082 GNDA.n1066 3.4105
R15749 GNDA.n1104 GNDA.n1066 3.4105
R15750 GNDA.n1081 GNDA.n1066 3.4105
R15751 GNDA.n1106 GNDA.n1066 3.4105
R15752 GNDA.n1080 GNDA.n1066 3.4105
R15753 GNDA.n1108 GNDA.n1066 3.4105
R15754 GNDA.n1079 GNDA.n1066 3.4105
R15755 GNDA.n1110 GNDA.n1066 3.4105
R15756 GNDA.n1078 GNDA.n1066 3.4105
R15757 GNDA.n1112 GNDA.n1066 3.4105
R15758 GNDA.n1077 GNDA.n1066 3.4105
R15759 GNDA.n1114 GNDA.n1066 3.4105
R15760 GNDA.n1076 GNDA.n1066 3.4105
R15761 GNDA.n1115 GNDA.n1066 3.4105
R15762 GNDA.n1162 GNDA.n1066 3.4105
R15763 GNDA.n1164 GNDA.n1066 3.4105
R15764 GNDA.n1166 GNDA.n802 3.4105
R15765 GNDA.n1090 GNDA.n802 3.4105
R15766 GNDA.n1088 GNDA.n802 3.4105
R15767 GNDA.n1092 GNDA.n802 3.4105
R15768 GNDA.n1087 GNDA.n802 3.4105
R15769 GNDA.n1094 GNDA.n802 3.4105
R15770 GNDA.n1086 GNDA.n802 3.4105
R15771 GNDA.n1096 GNDA.n802 3.4105
R15772 GNDA.n1085 GNDA.n802 3.4105
R15773 GNDA.n1098 GNDA.n802 3.4105
R15774 GNDA.n1084 GNDA.n802 3.4105
R15775 GNDA.n1100 GNDA.n802 3.4105
R15776 GNDA.n1083 GNDA.n802 3.4105
R15777 GNDA.n1102 GNDA.n802 3.4105
R15778 GNDA.n1082 GNDA.n802 3.4105
R15779 GNDA.n1104 GNDA.n802 3.4105
R15780 GNDA.n1081 GNDA.n802 3.4105
R15781 GNDA.n1106 GNDA.n802 3.4105
R15782 GNDA.n1080 GNDA.n802 3.4105
R15783 GNDA.n1108 GNDA.n802 3.4105
R15784 GNDA.n1079 GNDA.n802 3.4105
R15785 GNDA.n1110 GNDA.n802 3.4105
R15786 GNDA.n1078 GNDA.n802 3.4105
R15787 GNDA.n1112 GNDA.n802 3.4105
R15788 GNDA.n1077 GNDA.n802 3.4105
R15789 GNDA.n1114 GNDA.n802 3.4105
R15790 GNDA.n1076 GNDA.n802 3.4105
R15791 GNDA.n1115 GNDA.n802 3.4105
R15792 GNDA.n1162 GNDA.n802 3.4105
R15793 GNDA.n1164 GNDA.n802 3.4105
R15794 GNDA.n1166 GNDA.n1067 3.4105
R15795 GNDA.n1090 GNDA.n1067 3.4105
R15796 GNDA.n1088 GNDA.n1067 3.4105
R15797 GNDA.n1092 GNDA.n1067 3.4105
R15798 GNDA.n1087 GNDA.n1067 3.4105
R15799 GNDA.n1094 GNDA.n1067 3.4105
R15800 GNDA.n1086 GNDA.n1067 3.4105
R15801 GNDA.n1096 GNDA.n1067 3.4105
R15802 GNDA.n1085 GNDA.n1067 3.4105
R15803 GNDA.n1098 GNDA.n1067 3.4105
R15804 GNDA.n1084 GNDA.n1067 3.4105
R15805 GNDA.n1100 GNDA.n1067 3.4105
R15806 GNDA.n1083 GNDA.n1067 3.4105
R15807 GNDA.n1102 GNDA.n1067 3.4105
R15808 GNDA.n1082 GNDA.n1067 3.4105
R15809 GNDA.n1104 GNDA.n1067 3.4105
R15810 GNDA.n1081 GNDA.n1067 3.4105
R15811 GNDA.n1106 GNDA.n1067 3.4105
R15812 GNDA.n1080 GNDA.n1067 3.4105
R15813 GNDA.n1108 GNDA.n1067 3.4105
R15814 GNDA.n1079 GNDA.n1067 3.4105
R15815 GNDA.n1110 GNDA.n1067 3.4105
R15816 GNDA.n1078 GNDA.n1067 3.4105
R15817 GNDA.n1112 GNDA.n1067 3.4105
R15818 GNDA.n1077 GNDA.n1067 3.4105
R15819 GNDA.n1114 GNDA.n1067 3.4105
R15820 GNDA.n1076 GNDA.n1067 3.4105
R15821 GNDA.n1115 GNDA.n1067 3.4105
R15822 GNDA.n1162 GNDA.n1067 3.4105
R15823 GNDA.n1164 GNDA.n1067 3.4105
R15824 GNDA.n1166 GNDA.n801 3.4105
R15825 GNDA.n1090 GNDA.n801 3.4105
R15826 GNDA.n1088 GNDA.n801 3.4105
R15827 GNDA.n1092 GNDA.n801 3.4105
R15828 GNDA.n1087 GNDA.n801 3.4105
R15829 GNDA.n1094 GNDA.n801 3.4105
R15830 GNDA.n1086 GNDA.n801 3.4105
R15831 GNDA.n1096 GNDA.n801 3.4105
R15832 GNDA.n1085 GNDA.n801 3.4105
R15833 GNDA.n1098 GNDA.n801 3.4105
R15834 GNDA.n1084 GNDA.n801 3.4105
R15835 GNDA.n1100 GNDA.n801 3.4105
R15836 GNDA.n1083 GNDA.n801 3.4105
R15837 GNDA.n1102 GNDA.n801 3.4105
R15838 GNDA.n1082 GNDA.n801 3.4105
R15839 GNDA.n1104 GNDA.n801 3.4105
R15840 GNDA.n1081 GNDA.n801 3.4105
R15841 GNDA.n1106 GNDA.n801 3.4105
R15842 GNDA.n1080 GNDA.n801 3.4105
R15843 GNDA.n1108 GNDA.n801 3.4105
R15844 GNDA.n1079 GNDA.n801 3.4105
R15845 GNDA.n1110 GNDA.n801 3.4105
R15846 GNDA.n1078 GNDA.n801 3.4105
R15847 GNDA.n1112 GNDA.n801 3.4105
R15848 GNDA.n1077 GNDA.n801 3.4105
R15849 GNDA.n1114 GNDA.n801 3.4105
R15850 GNDA.n1076 GNDA.n801 3.4105
R15851 GNDA.n1115 GNDA.n801 3.4105
R15852 GNDA.n1162 GNDA.n801 3.4105
R15853 GNDA.n1164 GNDA.n801 3.4105
R15854 GNDA.n1166 GNDA.n1068 3.4105
R15855 GNDA.n1090 GNDA.n1068 3.4105
R15856 GNDA.n1088 GNDA.n1068 3.4105
R15857 GNDA.n1092 GNDA.n1068 3.4105
R15858 GNDA.n1087 GNDA.n1068 3.4105
R15859 GNDA.n1094 GNDA.n1068 3.4105
R15860 GNDA.n1086 GNDA.n1068 3.4105
R15861 GNDA.n1096 GNDA.n1068 3.4105
R15862 GNDA.n1085 GNDA.n1068 3.4105
R15863 GNDA.n1098 GNDA.n1068 3.4105
R15864 GNDA.n1084 GNDA.n1068 3.4105
R15865 GNDA.n1100 GNDA.n1068 3.4105
R15866 GNDA.n1083 GNDA.n1068 3.4105
R15867 GNDA.n1102 GNDA.n1068 3.4105
R15868 GNDA.n1082 GNDA.n1068 3.4105
R15869 GNDA.n1104 GNDA.n1068 3.4105
R15870 GNDA.n1081 GNDA.n1068 3.4105
R15871 GNDA.n1106 GNDA.n1068 3.4105
R15872 GNDA.n1080 GNDA.n1068 3.4105
R15873 GNDA.n1108 GNDA.n1068 3.4105
R15874 GNDA.n1079 GNDA.n1068 3.4105
R15875 GNDA.n1110 GNDA.n1068 3.4105
R15876 GNDA.n1078 GNDA.n1068 3.4105
R15877 GNDA.n1112 GNDA.n1068 3.4105
R15878 GNDA.n1077 GNDA.n1068 3.4105
R15879 GNDA.n1114 GNDA.n1068 3.4105
R15880 GNDA.n1076 GNDA.n1068 3.4105
R15881 GNDA.n1115 GNDA.n1068 3.4105
R15882 GNDA.n1162 GNDA.n1068 3.4105
R15883 GNDA.n1164 GNDA.n1068 3.4105
R15884 GNDA.n1166 GNDA.n800 3.4105
R15885 GNDA.n1090 GNDA.n800 3.4105
R15886 GNDA.n1088 GNDA.n800 3.4105
R15887 GNDA.n1092 GNDA.n800 3.4105
R15888 GNDA.n1087 GNDA.n800 3.4105
R15889 GNDA.n1094 GNDA.n800 3.4105
R15890 GNDA.n1086 GNDA.n800 3.4105
R15891 GNDA.n1096 GNDA.n800 3.4105
R15892 GNDA.n1085 GNDA.n800 3.4105
R15893 GNDA.n1098 GNDA.n800 3.4105
R15894 GNDA.n1084 GNDA.n800 3.4105
R15895 GNDA.n1100 GNDA.n800 3.4105
R15896 GNDA.n1083 GNDA.n800 3.4105
R15897 GNDA.n1102 GNDA.n800 3.4105
R15898 GNDA.n1082 GNDA.n800 3.4105
R15899 GNDA.n1104 GNDA.n800 3.4105
R15900 GNDA.n1081 GNDA.n800 3.4105
R15901 GNDA.n1106 GNDA.n800 3.4105
R15902 GNDA.n1080 GNDA.n800 3.4105
R15903 GNDA.n1108 GNDA.n800 3.4105
R15904 GNDA.n1079 GNDA.n800 3.4105
R15905 GNDA.n1110 GNDA.n800 3.4105
R15906 GNDA.n1078 GNDA.n800 3.4105
R15907 GNDA.n1112 GNDA.n800 3.4105
R15908 GNDA.n1077 GNDA.n800 3.4105
R15909 GNDA.n1114 GNDA.n800 3.4105
R15910 GNDA.n1076 GNDA.n800 3.4105
R15911 GNDA.n1115 GNDA.n800 3.4105
R15912 GNDA.n1162 GNDA.n800 3.4105
R15913 GNDA.n1164 GNDA.n800 3.4105
R15914 GNDA.n1166 GNDA.n1069 3.4105
R15915 GNDA.n1090 GNDA.n1069 3.4105
R15916 GNDA.n1088 GNDA.n1069 3.4105
R15917 GNDA.n1092 GNDA.n1069 3.4105
R15918 GNDA.n1087 GNDA.n1069 3.4105
R15919 GNDA.n1094 GNDA.n1069 3.4105
R15920 GNDA.n1086 GNDA.n1069 3.4105
R15921 GNDA.n1096 GNDA.n1069 3.4105
R15922 GNDA.n1085 GNDA.n1069 3.4105
R15923 GNDA.n1098 GNDA.n1069 3.4105
R15924 GNDA.n1084 GNDA.n1069 3.4105
R15925 GNDA.n1100 GNDA.n1069 3.4105
R15926 GNDA.n1083 GNDA.n1069 3.4105
R15927 GNDA.n1102 GNDA.n1069 3.4105
R15928 GNDA.n1082 GNDA.n1069 3.4105
R15929 GNDA.n1104 GNDA.n1069 3.4105
R15930 GNDA.n1081 GNDA.n1069 3.4105
R15931 GNDA.n1106 GNDA.n1069 3.4105
R15932 GNDA.n1080 GNDA.n1069 3.4105
R15933 GNDA.n1108 GNDA.n1069 3.4105
R15934 GNDA.n1079 GNDA.n1069 3.4105
R15935 GNDA.n1110 GNDA.n1069 3.4105
R15936 GNDA.n1078 GNDA.n1069 3.4105
R15937 GNDA.n1112 GNDA.n1069 3.4105
R15938 GNDA.n1077 GNDA.n1069 3.4105
R15939 GNDA.n1114 GNDA.n1069 3.4105
R15940 GNDA.n1076 GNDA.n1069 3.4105
R15941 GNDA.n1115 GNDA.n1069 3.4105
R15942 GNDA.n1162 GNDA.n1069 3.4105
R15943 GNDA.n1164 GNDA.n1069 3.4105
R15944 GNDA.n1166 GNDA.n799 3.4105
R15945 GNDA.n1090 GNDA.n799 3.4105
R15946 GNDA.n1088 GNDA.n799 3.4105
R15947 GNDA.n1092 GNDA.n799 3.4105
R15948 GNDA.n1087 GNDA.n799 3.4105
R15949 GNDA.n1094 GNDA.n799 3.4105
R15950 GNDA.n1086 GNDA.n799 3.4105
R15951 GNDA.n1096 GNDA.n799 3.4105
R15952 GNDA.n1085 GNDA.n799 3.4105
R15953 GNDA.n1098 GNDA.n799 3.4105
R15954 GNDA.n1084 GNDA.n799 3.4105
R15955 GNDA.n1100 GNDA.n799 3.4105
R15956 GNDA.n1083 GNDA.n799 3.4105
R15957 GNDA.n1102 GNDA.n799 3.4105
R15958 GNDA.n1082 GNDA.n799 3.4105
R15959 GNDA.n1104 GNDA.n799 3.4105
R15960 GNDA.n1081 GNDA.n799 3.4105
R15961 GNDA.n1106 GNDA.n799 3.4105
R15962 GNDA.n1080 GNDA.n799 3.4105
R15963 GNDA.n1108 GNDA.n799 3.4105
R15964 GNDA.n1079 GNDA.n799 3.4105
R15965 GNDA.n1110 GNDA.n799 3.4105
R15966 GNDA.n1078 GNDA.n799 3.4105
R15967 GNDA.n1112 GNDA.n799 3.4105
R15968 GNDA.n1077 GNDA.n799 3.4105
R15969 GNDA.n1114 GNDA.n799 3.4105
R15970 GNDA.n1076 GNDA.n799 3.4105
R15971 GNDA.n1115 GNDA.n799 3.4105
R15972 GNDA.n1162 GNDA.n799 3.4105
R15973 GNDA.n1164 GNDA.n799 3.4105
R15974 GNDA.n1166 GNDA.n1070 3.4105
R15975 GNDA.n1090 GNDA.n1070 3.4105
R15976 GNDA.n1088 GNDA.n1070 3.4105
R15977 GNDA.n1092 GNDA.n1070 3.4105
R15978 GNDA.n1087 GNDA.n1070 3.4105
R15979 GNDA.n1094 GNDA.n1070 3.4105
R15980 GNDA.n1086 GNDA.n1070 3.4105
R15981 GNDA.n1096 GNDA.n1070 3.4105
R15982 GNDA.n1085 GNDA.n1070 3.4105
R15983 GNDA.n1098 GNDA.n1070 3.4105
R15984 GNDA.n1084 GNDA.n1070 3.4105
R15985 GNDA.n1100 GNDA.n1070 3.4105
R15986 GNDA.n1083 GNDA.n1070 3.4105
R15987 GNDA.n1102 GNDA.n1070 3.4105
R15988 GNDA.n1082 GNDA.n1070 3.4105
R15989 GNDA.n1104 GNDA.n1070 3.4105
R15990 GNDA.n1081 GNDA.n1070 3.4105
R15991 GNDA.n1106 GNDA.n1070 3.4105
R15992 GNDA.n1080 GNDA.n1070 3.4105
R15993 GNDA.n1108 GNDA.n1070 3.4105
R15994 GNDA.n1079 GNDA.n1070 3.4105
R15995 GNDA.n1110 GNDA.n1070 3.4105
R15996 GNDA.n1078 GNDA.n1070 3.4105
R15997 GNDA.n1112 GNDA.n1070 3.4105
R15998 GNDA.n1077 GNDA.n1070 3.4105
R15999 GNDA.n1114 GNDA.n1070 3.4105
R16000 GNDA.n1076 GNDA.n1070 3.4105
R16001 GNDA.n1115 GNDA.n1070 3.4105
R16002 GNDA.n1162 GNDA.n1070 3.4105
R16003 GNDA.n1164 GNDA.n1070 3.4105
R16004 GNDA.n1166 GNDA.n798 3.4105
R16005 GNDA.n1090 GNDA.n798 3.4105
R16006 GNDA.n1088 GNDA.n798 3.4105
R16007 GNDA.n1092 GNDA.n798 3.4105
R16008 GNDA.n1087 GNDA.n798 3.4105
R16009 GNDA.n1094 GNDA.n798 3.4105
R16010 GNDA.n1086 GNDA.n798 3.4105
R16011 GNDA.n1096 GNDA.n798 3.4105
R16012 GNDA.n1085 GNDA.n798 3.4105
R16013 GNDA.n1098 GNDA.n798 3.4105
R16014 GNDA.n1084 GNDA.n798 3.4105
R16015 GNDA.n1100 GNDA.n798 3.4105
R16016 GNDA.n1083 GNDA.n798 3.4105
R16017 GNDA.n1102 GNDA.n798 3.4105
R16018 GNDA.n1082 GNDA.n798 3.4105
R16019 GNDA.n1104 GNDA.n798 3.4105
R16020 GNDA.n1081 GNDA.n798 3.4105
R16021 GNDA.n1106 GNDA.n798 3.4105
R16022 GNDA.n1080 GNDA.n798 3.4105
R16023 GNDA.n1108 GNDA.n798 3.4105
R16024 GNDA.n1079 GNDA.n798 3.4105
R16025 GNDA.n1110 GNDA.n798 3.4105
R16026 GNDA.n1078 GNDA.n798 3.4105
R16027 GNDA.n1112 GNDA.n798 3.4105
R16028 GNDA.n1077 GNDA.n798 3.4105
R16029 GNDA.n1114 GNDA.n798 3.4105
R16030 GNDA.n1076 GNDA.n798 3.4105
R16031 GNDA.n1115 GNDA.n798 3.4105
R16032 GNDA.n1162 GNDA.n798 3.4105
R16033 GNDA.n1164 GNDA.n798 3.4105
R16034 GNDA.n1166 GNDA.n1071 3.4105
R16035 GNDA.n1090 GNDA.n1071 3.4105
R16036 GNDA.n1088 GNDA.n1071 3.4105
R16037 GNDA.n1092 GNDA.n1071 3.4105
R16038 GNDA.n1087 GNDA.n1071 3.4105
R16039 GNDA.n1094 GNDA.n1071 3.4105
R16040 GNDA.n1086 GNDA.n1071 3.4105
R16041 GNDA.n1096 GNDA.n1071 3.4105
R16042 GNDA.n1085 GNDA.n1071 3.4105
R16043 GNDA.n1098 GNDA.n1071 3.4105
R16044 GNDA.n1084 GNDA.n1071 3.4105
R16045 GNDA.n1100 GNDA.n1071 3.4105
R16046 GNDA.n1083 GNDA.n1071 3.4105
R16047 GNDA.n1102 GNDA.n1071 3.4105
R16048 GNDA.n1082 GNDA.n1071 3.4105
R16049 GNDA.n1104 GNDA.n1071 3.4105
R16050 GNDA.n1081 GNDA.n1071 3.4105
R16051 GNDA.n1106 GNDA.n1071 3.4105
R16052 GNDA.n1080 GNDA.n1071 3.4105
R16053 GNDA.n1108 GNDA.n1071 3.4105
R16054 GNDA.n1079 GNDA.n1071 3.4105
R16055 GNDA.n1110 GNDA.n1071 3.4105
R16056 GNDA.n1078 GNDA.n1071 3.4105
R16057 GNDA.n1112 GNDA.n1071 3.4105
R16058 GNDA.n1077 GNDA.n1071 3.4105
R16059 GNDA.n1114 GNDA.n1071 3.4105
R16060 GNDA.n1076 GNDA.n1071 3.4105
R16061 GNDA.n1115 GNDA.n1071 3.4105
R16062 GNDA.n1162 GNDA.n1071 3.4105
R16063 GNDA.n1164 GNDA.n1071 3.4105
R16064 GNDA.n1166 GNDA.n797 3.4105
R16065 GNDA.n1090 GNDA.n797 3.4105
R16066 GNDA.n1088 GNDA.n797 3.4105
R16067 GNDA.n1092 GNDA.n797 3.4105
R16068 GNDA.n1087 GNDA.n797 3.4105
R16069 GNDA.n1094 GNDA.n797 3.4105
R16070 GNDA.n1086 GNDA.n797 3.4105
R16071 GNDA.n1096 GNDA.n797 3.4105
R16072 GNDA.n1085 GNDA.n797 3.4105
R16073 GNDA.n1098 GNDA.n797 3.4105
R16074 GNDA.n1084 GNDA.n797 3.4105
R16075 GNDA.n1100 GNDA.n797 3.4105
R16076 GNDA.n1083 GNDA.n797 3.4105
R16077 GNDA.n1102 GNDA.n797 3.4105
R16078 GNDA.n1082 GNDA.n797 3.4105
R16079 GNDA.n1104 GNDA.n797 3.4105
R16080 GNDA.n1081 GNDA.n797 3.4105
R16081 GNDA.n1106 GNDA.n797 3.4105
R16082 GNDA.n1080 GNDA.n797 3.4105
R16083 GNDA.n1108 GNDA.n797 3.4105
R16084 GNDA.n1079 GNDA.n797 3.4105
R16085 GNDA.n1110 GNDA.n797 3.4105
R16086 GNDA.n1078 GNDA.n797 3.4105
R16087 GNDA.n1112 GNDA.n797 3.4105
R16088 GNDA.n1077 GNDA.n797 3.4105
R16089 GNDA.n1114 GNDA.n797 3.4105
R16090 GNDA.n1076 GNDA.n797 3.4105
R16091 GNDA.n1115 GNDA.n797 3.4105
R16092 GNDA.n1162 GNDA.n797 3.4105
R16093 GNDA.n1164 GNDA.n797 3.4105
R16094 GNDA.n1166 GNDA.n1072 3.4105
R16095 GNDA.n1090 GNDA.n1072 3.4105
R16096 GNDA.n1088 GNDA.n1072 3.4105
R16097 GNDA.n1092 GNDA.n1072 3.4105
R16098 GNDA.n1087 GNDA.n1072 3.4105
R16099 GNDA.n1094 GNDA.n1072 3.4105
R16100 GNDA.n1086 GNDA.n1072 3.4105
R16101 GNDA.n1096 GNDA.n1072 3.4105
R16102 GNDA.n1085 GNDA.n1072 3.4105
R16103 GNDA.n1098 GNDA.n1072 3.4105
R16104 GNDA.n1084 GNDA.n1072 3.4105
R16105 GNDA.n1100 GNDA.n1072 3.4105
R16106 GNDA.n1083 GNDA.n1072 3.4105
R16107 GNDA.n1102 GNDA.n1072 3.4105
R16108 GNDA.n1082 GNDA.n1072 3.4105
R16109 GNDA.n1104 GNDA.n1072 3.4105
R16110 GNDA.n1081 GNDA.n1072 3.4105
R16111 GNDA.n1106 GNDA.n1072 3.4105
R16112 GNDA.n1080 GNDA.n1072 3.4105
R16113 GNDA.n1108 GNDA.n1072 3.4105
R16114 GNDA.n1079 GNDA.n1072 3.4105
R16115 GNDA.n1110 GNDA.n1072 3.4105
R16116 GNDA.n1078 GNDA.n1072 3.4105
R16117 GNDA.n1112 GNDA.n1072 3.4105
R16118 GNDA.n1077 GNDA.n1072 3.4105
R16119 GNDA.n1114 GNDA.n1072 3.4105
R16120 GNDA.n1076 GNDA.n1072 3.4105
R16121 GNDA.n1115 GNDA.n1072 3.4105
R16122 GNDA.n1162 GNDA.n1072 3.4105
R16123 GNDA.n1164 GNDA.n1072 3.4105
R16124 GNDA.n1166 GNDA.n796 3.4105
R16125 GNDA.n1090 GNDA.n796 3.4105
R16126 GNDA.n1088 GNDA.n796 3.4105
R16127 GNDA.n1092 GNDA.n796 3.4105
R16128 GNDA.n1087 GNDA.n796 3.4105
R16129 GNDA.n1094 GNDA.n796 3.4105
R16130 GNDA.n1086 GNDA.n796 3.4105
R16131 GNDA.n1096 GNDA.n796 3.4105
R16132 GNDA.n1085 GNDA.n796 3.4105
R16133 GNDA.n1098 GNDA.n796 3.4105
R16134 GNDA.n1084 GNDA.n796 3.4105
R16135 GNDA.n1100 GNDA.n796 3.4105
R16136 GNDA.n1083 GNDA.n796 3.4105
R16137 GNDA.n1102 GNDA.n796 3.4105
R16138 GNDA.n1082 GNDA.n796 3.4105
R16139 GNDA.n1104 GNDA.n796 3.4105
R16140 GNDA.n1081 GNDA.n796 3.4105
R16141 GNDA.n1106 GNDA.n796 3.4105
R16142 GNDA.n1080 GNDA.n796 3.4105
R16143 GNDA.n1108 GNDA.n796 3.4105
R16144 GNDA.n1079 GNDA.n796 3.4105
R16145 GNDA.n1110 GNDA.n796 3.4105
R16146 GNDA.n1078 GNDA.n796 3.4105
R16147 GNDA.n1112 GNDA.n796 3.4105
R16148 GNDA.n1077 GNDA.n796 3.4105
R16149 GNDA.n1114 GNDA.n796 3.4105
R16150 GNDA.n1076 GNDA.n796 3.4105
R16151 GNDA.n1115 GNDA.n796 3.4105
R16152 GNDA.n1162 GNDA.n796 3.4105
R16153 GNDA.n1164 GNDA.n796 3.4105
R16154 GNDA.n1166 GNDA.n1073 3.4105
R16155 GNDA.n1090 GNDA.n1073 3.4105
R16156 GNDA.n1088 GNDA.n1073 3.4105
R16157 GNDA.n1092 GNDA.n1073 3.4105
R16158 GNDA.n1087 GNDA.n1073 3.4105
R16159 GNDA.n1094 GNDA.n1073 3.4105
R16160 GNDA.n1086 GNDA.n1073 3.4105
R16161 GNDA.n1096 GNDA.n1073 3.4105
R16162 GNDA.n1085 GNDA.n1073 3.4105
R16163 GNDA.n1098 GNDA.n1073 3.4105
R16164 GNDA.n1084 GNDA.n1073 3.4105
R16165 GNDA.n1100 GNDA.n1073 3.4105
R16166 GNDA.n1083 GNDA.n1073 3.4105
R16167 GNDA.n1102 GNDA.n1073 3.4105
R16168 GNDA.n1082 GNDA.n1073 3.4105
R16169 GNDA.n1104 GNDA.n1073 3.4105
R16170 GNDA.n1081 GNDA.n1073 3.4105
R16171 GNDA.n1106 GNDA.n1073 3.4105
R16172 GNDA.n1080 GNDA.n1073 3.4105
R16173 GNDA.n1108 GNDA.n1073 3.4105
R16174 GNDA.n1079 GNDA.n1073 3.4105
R16175 GNDA.n1110 GNDA.n1073 3.4105
R16176 GNDA.n1078 GNDA.n1073 3.4105
R16177 GNDA.n1112 GNDA.n1073 3.4105
R16178 GNDA.n1077 GNDA.n1073 3.4105
R16179 GNDA.n1114 GNDA.n1073 3.4105
R16180 GNDA.n1076 GNDA.n1073 3.4105
R16181 GNDA.n1115 GNDA.n1073 3.4105
R16182 GNDA.n1162 GNDA.n1073 3.4105
R16183 GNDA.n1164 GNDA.n1073 3.4105
R16184 GNDA.n1166 GNDA.n795 3.4105
R16185 GNDA.n1090 GNDA.n795 3.4105
R16186 GNDA.n1088 GNDA.n795 3.4105
R16187 GNDA.n1092 GNDA.n795 3.4105
R16188 GNDA.n1087 GNDA.n795 3.4105
R16189 GNDA.n1094 GNDA.n795 3.4105
R16190 GNDA.n1086 GNDA.n795 3.4105
R16191 GNDA.n1096 GNDA.n795 3.4105
R16192 GNDA.n1085 GNDA.n795 3.4105
R16193 GNDA.n1098 GNDA.n795 3.4105
R16194 GNDA.n1084 GNDA.n795 3.4105
R16195 GNDA.n1100 GNDA.n795 3.4105
R16196 GNDA.n1083 GNDA.n795 3.4105
R16197 GNDA.n1102 GNDA.n795 3.4105
R16198 GNDA.n1082 GNDA.n795 3.4105
R16199 GNDA.n1104 GNDA.n795 3.4105
R16200 GNDA.n1081 GNDA.n795 3.4105
R16201 GNDA.n1106 GNDA.n795 3.4105
R16202 GNDA.n1080 GNDA.n795 3.4105
R16203 GNDA.n1108 GNDA.n795 3.4105
R16204 GNDA.n1079 GNDA.n795 3.4105
R16205 GNDA.n1110 GNDA.n795 3.4105
R16206 GNDA.n1078 GNDA.n795 3.4105
R16207 GNDA.n1112 GNDA.n795 3.4105
R16208 GNDA.n1077 GNDA.n795 3.4105
R16209 GNDA.n1114 GNDA.n795 3.4105
R16210 GNDA.n1076 GNDA.n795 3.4105
R16211 GNDA.n1115 GNDA.n795 3.4105
R16212 GNDA.n1162 GNDA.n795 3.4105
R16213 GNDA.n1164 GNDA.n795 3.4105
R16214 GNDA.n1166 GNDA.n1165 3.4105
R16215 GNDA.n1165 GNDA.n1090 3.4105
R16216 GNDA.n1165 GNDA.n1088 3.4105
R16217 GNDA.n1165 GNDA.n1092 3.4105
R16218 GNDA.n1165 GNDA.n1087 3.4105
R16219 GNDA.n1165 GNDA.n1094 3.4105
R16220 GNDA.n1165 GNDA.n1086 3.4105
R16221 GNDA.n1165 GNDA.n1096 3.4105
R16222 GNDA.n1165 GNDA.n1085 3.4105
R16223 GNDA.n1165 GNDA.n1098 3.4105
R16224 GNDA.n1165 GNDA.n1084 3.4105
R16225 GNDA.n1165 GNDA.n1100 3.4105
R16226 GNDA.n1165 GNDA.n1083 3.4105
R16227 GNDA.n1165 GNDA.n1102 3.4105
R16228 GNDA.n1165 GNDA.n1082 3.4105
R16229 GNDA.n1165 GNDA.n1104 3.4105
R16230 GNDA.n1165 GNDA.n1081 3.4105
R16231 GNDA.n1165 GNDA.n1106 3.4105
R16232 GNDA.n1165 GNDA.n1080 3.4105
R16233 GNDA.n1165 GNDA.n1108 3.4105
R16234 GNDA.n1165 GNDA.n1079 3.4105
R16235 GNDA.n1165 GNDA.n1110 3.4105
R16236 GNDA.n1165 GNDA.n1078 3.4105
R16237 GNDA.n1165 GNDA.n1112 3.4105
R16238 GNDA.n1165 GNDA.n1077 3.4105
R16239 GNDA.n1165 GNDA.n1114 3.4105
R16240 GNDA.n1165 GNDA.n1076 3.4105
R16241 GNDA.n1165 GNDA.n1115 3.4105
R16242 GNDA.n1165 GNDA.n1164 3.4105
R16243 GNDA.n1053 GNDA.n824 3.4105
R16244 GNDA.n869 GNDA.n824 3.4105
R16245 GNDA.n869 GNDA.n823 3.4105
R16246 GNDA.n1055 GNDA.n869 3.4105
R16247 GNDA.n1057 GNDA.n869 3.4105
R16248 GNDA.n855 GNDA.n824 3.4105
R16249 GNDA.n855 GNDA.n826 3.4105
R16250 GNDA.n855 GNDA.n822 3.4105
R16251 GNDA.n855 GNDA.n827 3.4105
R16252 GNDA.n855 GNDA.n821 3.4105
R16253 GNDA.n855 GNDA.n828 3.4105
R16254 GNDA.n855 GNDA.n820 3.4105
R16255 GNDA.n855 GNDA.n829 3.4105
R16256 GNDA.n855 GNDA.n819 3.4105
R16257 GNDA.n855 GNDA.n830 3.4105
R16258 GNDA.n855 GNDA.n818 3.4105
R16259 GNDA.n855 GNDA.n831 3.4105
R16260 GNDA.n855 GNDA.n817 3.4105
R16261 GNDA.n855 GNDA.n832 3.4105
R16262 GNDA.n855 GNDA.n816 3.4105
R16263 GNDA.n855 GNDA.n833 3.4105
R16264 GNDA.n855 GNDA.n815 3.4105
R16265 GNDA.n855 GNDA.n834 3.4105
R16266 GNDA.n855 GNDA.n814 3.4105
R16267 GNDA.n855 GNDA.n835 3.4105
R16268 GNDA.n855 GNDA.n813 3.4105
R16269 GNDA.n855 GNDA.n836 3.4105
R16270 GNDA.n855 GNDA.n812 3.4105
R16271 GNDA.n855 GNDA.n837 3.4105
R16272 GNDA.n855 GNDA.n811 3.4105
R16273 GNDA.n855 GNDA.n838 3.4105
R16274 GNDA.n1055 GNDA.n855 3.4105
R16275 GNDA.n1057 GNDA.n855 3.4105
R16276 GNDA.n871 GNDA.n823 3.4105
R16277 GNDA.n871 GNDA.n826 3.4105
R16278 GNDA.n871 GNDA.n822 3.4105
R16279 GNDA.n871 GNDA.n827 3.4105
R16280 GNDA.n871 GNDA.n821 3.4105
R16281 GNDA.n871 GNDA.n828 3.4105
R16282 GNDA.n871 GNDA.n820 3.4105
R16283 GNDA.n871 GNDA.n829 3.4105
R16284 GNDA.n871 GNDA.n819 3.4105
R16285 GNDA.n871 GNDA.n830 3.4105
R16286 GNDA.n871 GNDA.n818 3.4105
R16287 GNDA.n871 GNDA.n831 3.4105
R16288 GNDA.n871 GNDA.n817 3.4105
R16289 GNDA.n871 GNDA.n832 3.4105
R16290 GNDA.n871 GNDA.n816 3.4105
R16291 GNDA.n871 GNDA.n833 3.4105
R16292 GNDA.n871 GNDA.n815 3.4105
R16293 GNDA.n871 GNDA.n834 3.4105
R16294 GNDA.n871 GNDA.n814 3.4105
R16295 GNDA.n871 GNDA.n835 3.4105
R16296 GNDA.n871 GNDA.n813 3.4105
R16297 GNDA.n871 GNDA.n836 3.4105
R16298 GNDA.n871 GNDA.n812 3.4105
R16299 GNDA.n871 GNDA.n837 3.4105
R16300 GNDA.n871 GNDA.n811 3.4105
R16301 GNDA.n871 GNDA.n838 3.4105
R16302 GNDA.n1055 GNDA.n871 3.4105
R16303 GNDA.n1057 GNDA.n871 3.4105
R16304 GNDA.n853 GNDA.n824 3.4105
R16305 GNDA.n853 GNDA.n825 3.4105
R16306 GNDA.n853 GNDA.n823 3.4105
R16307 GNDA.n853 GNDA.n826 3.4105
R16308 GNDA.n853 GNDA.n822 3.4105
R16309 GNDA.n853 GNDA.n827 3.4105
R16310 GNDA.n853 GNDA.n821 3.4105
R16311 GNDA.n853 GNDA.n828 3.4105
R16312 GNDA.n853 GNDA.n820 3.4105
R16313 GNDA.n853 GNDA.n829 3.4105
R16314 GNDA.n853 GNDA.n819 3.4105
R16315 GNDA.n853 GNDA.n830 3.4105
R16316 GNDA.n853 GNDA.n818 3.4105
R16317 GNDA.n853 GNDA.n831 3.4105
R16318 GNDA.n853 GNDA.n817 3.4105
R16319 GNDA.n853 GNDA.n832 3.4105
R16320 GNDA.n853 GNDA.n816 3.4105
R16321 GNDA.n853 GNDA.n833 3.4105
R16322 GNDA.n853 GNDA.n815 3.4105
R16323 GNDA.n853 GNDA.n834 3.4105
R16324 GNDA.n853 GNDA.n814 3.4105
R16325 GNDA.n853 GNDA.n835 3.4105
R16326 GNDA.n853 GNDA.n813 3.4105
R16327 GNDA.n853 GNDA.n836 3.4105
R16328 GNDA.n853 GNDA.n812 3.4105
R16329 GNDA.n853 GNDA.n837 3.4105
R16330 GNDA.n853 GNDA.n811 3.4105
R16331 GNDA.n853 GNDA.n838 3.4105
R16332 GNDA.n1055 GNDA.n853 3.4105
R16333 GNDA.n1057 GNDA.n853 3.4105
R16334 GNDA.n872 GNDA.n824 3.4105
R16335 GNDA.n872 GNDA.n825 3.4105
R16336 GNDA.n872 GNDA.n823 3.4105
R16337 GNDA.n872 GNDA.n826 3.4105
R16338 GNDA.n872 GNDA.n822 3.4105
R16339 GNDA.n872 GNDA.n827 3.4105
R16340 GNDA.n872 GNDA.n821 3.4105
R16341 GNDA.n872 GNDA.n828 3.4105
R16342 GNDA.n872 GNDA.n820 3.4105
R16343 GNDA.n872 GNDA.n829 3.4105
R16344 GNDA.n872 GNDA.n819 3.4105
R16345 GNDA.n872 GNDA.n830 3.4105
R16346 GNDA.n872 GNDA.n818 3.4105
R16347 GNDA.n872 GNDA.n831 3.4105
R16348 GNDA.n872 GNDA.n817 3.4105
R16349 GNDA.n872 GNDA.n832 3.4105
R16350 GNDA.n872 GNDA.n816 3.4105
R16351 GNDA.n872 GNDA.n833 3.4105
R16352 GNDA.n872 GNDA.n815 3.4105
R16353 GNDA.n872 GNDA.n834 3.4105
R16354 GNDA.n872 GNDA.n814 3.4105
R16355 GNDA.n872 GNDA.n835 3.4105
R16356 GNDA.n872 GNDA.n813 3.4105
R16357 GNDA.n872 GNDA.n836 3.4105
R16358 GNDA.n872 GNDA.n812 3.4105
R16359 GNDA.n872 GNDA.n837 3.4105
R16360 GNDA.n872 GNDA.n811 3.4105
R16361 GNDA.n872 GNDA.n838 3.4105
R16362 GNDA.n1055 GNDA.n872 3.4105
R16363 GNDA.n1057 GNDA.n872 3.4105
R16364 GNDA.n852 GNDA.n824 3.4105
R16365 GNDA.n852 GNDA.n825 3.4105
R16366 GNDA.n852 GNDA.n823 3.4105
R16367 GNDA.n852 GNDA.n826 3.4105
R16368 GNDA.n852 GNDA.n822 3.4105
R16369 GNDA.n852 GNDA.n827 3.4105
R16370 GNDA.n852 GNDA.n821 3.4105
R16371 GNDA.n852 GNDA.n828 3.4105
R16372 GNDA.n852 GNDA.n820 3.4105
R16373 GNDA.n852 GNDA.n829 3.4105
R16374 GNDA.n852 GNDA.n819 3.4105
R16375 GNDA.n852 GNDA.n830 3.4105
R16376 GNDA.n852 GNDA.n818 3.4105
R16377 GNDA.n852 GNDA.n831 3.4105
R16378 GNDA.n852 GNDA.n817 3.4105
R16379 GNDA.n852 GNDA.n832 3.4105
R16380 GNDA.n852 GNDA.n816 3.4105
R16381 GNDA.n852 GNDA.n833 3.4105
R16382 GNDA.n852 GNDA.n815 3.4105
R16383 GNDA.n852 GNDA.n834 3.4105
R16384 GNDA.n852 GNDA.n814 3.4105
R16385 GNDA.n852 GNDA.n835 3.4105
R16386 GNDA.n852 GNDA.n813 3.4105
R16387 GNDA.n852 GNDA.n836 3.4105
R16388 GNDA.n852 GNDA.n812 3.4105
R16389 GNDA.n852 GNDA.n837 3.4105
R16390 GNDA.n852 GNDA.n811 3.4105
R16391 GNDA.n852 GNDA.n838 3.4105
R16392 GNDA.n1055 GNDA.n852 3.4105
R16393 GNDA.n1057 GNDA.n852 3.4105
R16394 GNDA.n873 GNDA.n824 3.4105
R16395 GNDA.n873 GNDA.n825 3.4105
R16396 GNDA.n873 GNDA.n823 3.4105
R16397 GNDA.n873 GNDA.n826 3.4105
R16398 GNDA.n873 GNDA.n822 3.4105
R16399 GNDA.n873 GNDA.n827 3.4105
R16400 GNDA.n873 GNDA.n821 3.4105
R16401 GNDA.n873 GNDA.n828 3.4105
R16402 GNDA.n873 GNDA.n820 3.4105
R16403 GNDA.n873 GNDA.n829 3.4105
R16404 GNDA.n873 GNDA.n819 3.4105
R16405 GNDA.n873 GNDA.n830 3.4105
R16406 GNDA.n873 GNDA.n818 3.4105
R16407 GNDA.n873 GNDA.n831 3.4105
R16408 GNDA.n873 GNDA.n817 3.4105
R16409 GNDA.n873 GNDA.n832 3.4105
R16410 GNDA.n873 GNDA.n816 3.4105
R16411 GNDA.n873 GNDA.n833 3.4105
R16412 GNDA.n873 GNDA.n815 3.4105
R16413 GNDA.n873 GNDA.n834 3.4105
R16414 GNDA.n873 GNDA.n814 3.4105
R16415 GNDA.n873 GNDA.n835 3.4105
R16416 GNDA.n873 GNDA.n813 3.4105
R16417 GNDA.n873 GNDA.n836 3.4105
R16418 GNDA.n873 GNDA.n812 3.4105
R16419 GNDA.n873 GNDA.n837 3.4105
R16420 GNDA.n873 GNDA.n811 3.4105
R16421 GNDA.n873 GNDA.n838 3.4105
R16422 GNDA.n1055 GNDA.n873 3.4105
R16423 GNDA.n1057 GNDA.n873 3.4105
R16424 GNDA.n851 GNDA.n824 3.4105
R16425 GNDA.n851 GNDA.n825 3.4105
R16426 GNDA.n851 GNDA.n823 3.4105
R16427 GNDA.n851 GNDA.n826 3.4105
R16428 GNDA.n851 GNDA.n822 3.4105
R16429 GNDA.n851 GNDA.n827 3.4105
R16430 GNDA.n851 GNDA.n821 3.4105
R16431 GNDA.n851 GNDA.n828 3.4105
R16432 GNDA.n851 GNDA.n820 3.4105
R16433 GNDA.n851 GNDA.n829 3.4105
R16434 GNDA.n851 GNDA.n819 3.4105
R16435 GNDA.n851 GNDA.n830 3.4105
R16436 GNDA.n851 GNDA.n818 3.4105
R16437 GNDA.n851 GNDA.n831 3.4105
R16438 GNDA.n851 GNDA.n817 3.4105
R16439 GNDA.n851 GNDA.n832 3.4105
R16440 GNDA.n851 GNDA.n816 3.4105
R16441 GNDA.n851 GNDA.n833 3.4105
R16442 GNDA.n851 GNDA.n815 3.4105
R16443 GNDA.n851 GNDA.n834 3.4105
R16444 GNDA.n851 GNDA.n814 3.4105
R16445 GNDA.n851 GNDA.n835 3.4105
R16446 GNDA.n851 GNDA.n813 3.4105
R16447 GNDA.n851 GNDA.n836 3.4105
R16448 GNDA.n851 GNDA.n812 3.4105
R16449 GNDA.n851 GNDA.n837 3.4105
R16450 GNDA.n851 GNDA.n811 3.4105
R16451 GNDA.n851 GNDA.n838 3.4105
R16452 GNDA.n1055 GNDA.n851 3.4105
R16453 GNDA.n1057 GNDA.n851 3.4105
R16454 GNDA.n874 GNDA.n824 3.4105
R16455 GNDA.n874 GNDA.n825 3.4105
R16456 GNDA.n874 GNDA.n823 3.4105
R16457 GNDA.n874 GNDA.n826 3.4105
R16458 GNDA.n874 GNDA.n822 3.4105
R16459 GNDA.n874 GNDA.n827 3.4105
R16460 GNDA.n874 GNDA.n821 3.4105
R16461 GNDA.n874 GNDA.n828 3.4105
R16462 GNDA.n874 GNDA.n820 3.4105
R16463 GNDA.n874 GNDA.n829 3.4105
R16464 GNDA.n874 GNDA.n819 3.4105
R16465 GNDA.n874 GNDA.n830 3.4105
R16466 GNDA.n874 GNDA.n818 3.4105
R16467 GNDA.n874 GNDA.n831 3.4105
R16468 GNDA.n874 GNDA.n817 3.4105
R16469 GNDA.n874 GNDA.n832 3.4105
R16470 GNDA.n874 GNDA.n816 3.4105
R16471 GNDA.n874 GNDA.n833 3.4105
R16472 GNDA.n874 GNDA.n815 3.4105
R16473 GNDA.n874 GNDA.n834 3.4105
R16474 GNDA.n874 GNDA.n814 3.4105
R16475 GNDA.n874 GNDA.n835 3.4105
R16476 GNDA.n874 GNDA.n813 3.4105
R16477 GNDA.n874 GNDA.n836 3.4105
R16478 GNDA.n874 GNDA.n812 3.4105
R16479 GNDA.n874 GNDA.n837 3.4105
R16480 GNDA.n874 GNDA.n811 3.4105
R16481 GNDA.n874 GNDA.n838 3.4105
R16482 GNDA.n1055 GNDA.n874 3.4105
R16483 GNDA.n1057 GNDA.n874 3.4105
R16484 GNDA.n850 GNDA.n824 3.4105
R16485 GNDA.n850 GNDA.n825 3.4105
R16486 GNDA.n850 GNDA.n823 3.4105
R16487 GNDA.n850 GNDA.n826 3.4105
R16488 GNDA.n850 GNDA.n822 3.4105
R16489 GNDA.n850 GNDA.n827 3.4105
R16490 GNDA.n850 GNDA.n821 3.4105
R16491 GNDA.n850 GNDA.n828 3.4105
R16492 GNDA.n850 GNDA.n820 3.4105
R16493 GNDA.n850 GNDA.n829 3.4105
R16494 GNDA.n850 GNDA.n819 3.4105
R16495 GNDA.n850 GNDA.n830 3.4105
R16496 GNDA.n850 GNDA.n818 3.4105
R16497 GNDA.n850 GNDA.n831 3.4105
R16498 GNDA.n850 GNDA.n817 3.4105
R16499 GNDA.n850 GNDA.n832 3.4105
R16500 GNDA.n850 GNDA.n816 3.4105
R16501 GNDA.n850 GNDA.n833 3.4105
R16502 GNDA.n850 GNDA.n815 3.4105
R16503 GNDA.n850 GNDA.n834 3.4105
R16504 GNDA.n850 GNDA.n814 3.4105
R16505 GNDA.n850 GNDA.n835 3.4105
R16506 GNDA.n850 GNDA.n813 3.4105
R16507 GNDA.n850 GNDA.n836 3.4105
R16508 GNDA.n850 GNDA.n812 3.4105
R16509 GNDA.n850 GNDA.n837 3.4105
R16510 GNDA.n850 GNDA.n811 3.4105
R16511 GNDA.n850 GNDA.n838 3.4105
R16512 GNDA.n1055 GNDA.n850 3.4105
R16513 GNDA.n1057 GNDA.n850 3.4105
R16514 GNDA.n875 GNDA.n824 3.4105
R16515 GNDA.n875 GNDA.n825 3.4105
R16516 GNDA.n875 GNDA.n823 3.4105
R16517 GNDA.n875 GNDA.n826 3.4105
R16518 GNDA.n875 GNDA.n822 3.4105
R16519 GNDA.n875 GNDA.n827 3.4105
R16520 GNDA.n875 GNDA.n821 3.4105
R16521 GNDA.n875 GNDA.n828 3.4105
R16522 GNDA.n875 GNDA.n820 3.4105
R16523 GNDA.n875 GNDA.n829 3.4105
R16524 GNDA.n875 GNDA.n819 3.4105
R16525 GNDA.n875 GNDA.n830 3.4105
R16526 GNDA.n875 GNDA.n818 3.4105
R16527 GNDA.n875 GNDA.n831 3.4105
R16528 GNDA.n875 GNDA.n817 3.4105
R16529 GNDA.n875 GNDA.n832 3.4105
R16530 GNDA.n875 GNDA.n816 3.4105
R16531 GNDA.n875 GNDA.n833 3.4105
R16532 GNDA.n875 GNDA.n815 3.4105
R16533 GNDA.n875 GNDA.n834 3.4105
R16534 GNDA.n875 GNDA.n814 3.4105
R16535 GNDA.n875 GNDA.n835 3.4105
R16536 GNDA.n875 GNDA.n813 3.4105
R16537 GNDA.n875 GNDA.n836 3.4105
R16538 GNDA.n875 GNDA.n812 3.4105
R16539 GNDA.n875 GNDA.n837 3.4105
R16540 GNDA.n875 GNDA.n811 3.4105
R16541 GNDA.n875 GNDA.n838 3.4105
R16542 GNDA.n1055 GNDA.n875 3.4105
R16543 GNDA.n1057 GNDA.n875 3.4105
R16544 GNDA.n849 GNDA.n824 3.4105
R16545 GNDA.n849 GNDA.n825 3.4105
R16546 GNDA.n849 GNDA.n823 3.4105
R16547 GNDA.n849 GNDA.n826 3.4105
R16548 GNDA.n849 GNDA.n822 3.4105
R16549 GNDA.n849 GNDA.n827 3.4105
R16550 GNDA.n849 GNDA.n821 3.4105
R16551 GNDA.n849 GNDA.n828 3.4105
R16552 GNDA.n849 GNDA.n820 3.4105
R16553 GNDA.n849 GNDA.n829 3.4105
R16554 GNDA.n849 GNDA.n819 3.4105
R16555 GNDA.n849 GNDA.n830 3.4105
R16556 GNDA.n849 GNDA.n818 3.4105
R16557 GNDA.n849 GNDA.n831 3.4105
R16558 GNDA.n849 GNDA.n817 3.4105
R16559 GNDA.n849 GNDA.n832 3.4105
R16560 GNDA.n849 GNDA.n816 3.4105
R16561 GNDA.n849 GNDA.n833 3.4105
R16562 GNDA.n849 GNDA.n815 3.4105
R16563 GNDA.n849 GNDA.n834 3.4105
R16564 GNDA.n849 GNDA.n814 3.4105
R16565 GNDA.n849 GNDA.n835 3.4105
R16566 GNDA.n849 GNDA.n813 3.4105
R16567 GNDA.n849 GNDA.n836 3.4105
R16568 GNDA.n849 GNDA.n812 3.4105
R16569 GNDA.n849 GNDA.n837 3.4105
R16570 GNDA.n849 GNDA.n811 3.4105
R16571 GNDA.n849 GNDA.n838 3.4105
R16572 GNDA.n1055 GNDA.n849 3.4105
R16573 GNDA.n1057 GNDA.n849 3.4105
R16574 GNDA.n876 GNDA.n824 3.4105
R16575 GNDA.n876 GNDA.n825 3.4105
R16576 GNDA.n876 GNDA.n823 3.4105
R16577 GNDA.n876 GNDA.n826 3.4105
R16578 GNDA.n876 GNDA.n822 3.4105
R16579 GNDA.n876 GNDA.n827 3.4105
R16580 GNDA.n876 GNDA.n821 3.4105
R16581 GNDA.n876 GNDA.n828 3.4105
R16582 GNDA.n876 GNDA.n820 3.4105
R16583 GNDA.n876 GNDA.n829 3.4105
R16584 GNDA.n876 GNDA.n819 3.4105
R16585 GNDA.n876 GNDA.n830 3.4105
R16586 GNDA.n876 GNDA.n818 3.4105
R16587 GNDA.n876 GNDA.n831 3.4105
R16588 GNDA.n876 GNDA.n817 3.4105
R16589 GNDA.n876 GNDA.n832 3.4105
R16590 GNDA.n876 GNDA.n816 3.4105
R16591 GNDA.n876 GNDA.n833 3.4105
R16592 GNDA.n876 GNDA.n815 3.4105
R16593 GNDA.n876 GNDA.n834 3.4105
R16594 GNDA.n876 GNDA.n814 3.4105
R16595 GNDA.n876 GNDA.n835 3.4105
R16596 GNDA.n876 GNDA.n813 3.4105
R16597 GNDA.n876 GNDA.n836 3.4105
R16598 GNDA.n876 GNDA.n812 3.4105
R16599 GNDA.n876 GNDA.n837 3.4105
R16600 GNDA.n876 GNDA.n811 3.4105
R16601 GNDA.n876 GNDA.n838 3.4105
R16602 GNDA.n1055 GNDA.n876 3.4105
R16603 GNDA.n1057 GNDA.n876 3.4105
R16604 GNDA.n848 GNDA.n824 3.4105
R16605 GNDA.n848 GNDA.n825 3.4105
R16606 GNDA.n848 GNDA.n823 3.4105
R16607 GNDA.n848 GNDA.n826 3.4105
R16608 GNDA.n848 GNDA.n822 3.4105
R16609 GNDA.n848 GNDA.n827 3.4105
R16610 GNDA.n848 GNDA.n821 3.4105
R16611 GNDA.n848 GNDA.n828 3.4105
R16612 GNDA.n848 GNDA.n820 3.4105
R16613 GNDA.n848 GNDA.n829 3.4105
R16614 GNDA.n848 GNDA.n819 3.4105
R16615 GNDA.n848 GNDA.n830 3.4105
R16616 GNDA.n848 GNDA.n818 3.4105
R16617 GNDA.n848 GNDA.n831 3.4105
R16618 GNDA.n848 GNDA.n817 3.4105
R16619 GNDA.n848 GNDA.n832 3.4105
R16620 GNDA.n848 GNDA.n816 3.4105
R16621 GNDA.n848 GNDA.n833 3.4105
R16622 GNDA.n848 GNDA.n815 3.4105
R16623 GNDA.n848 GNDA.n834 3.4105
R16624 GNDA.n848 GNDA.n814 3.4105
R16625 GNDA.n848 GNDA.n835 3.4105
R16626 GNDA.n848 GNDA.n813 3.4105
R16627 GNDA.n848 GNDA.n836 3.4105
R16628 GNDA.n848 GNDA.n812 3.4105
R16629 GNDA.n848 GNDA.n837 3.4105
R16630 GNDA.n848 GNDA.n811 3.4105
R16631 GNDA.n848 GNDA.n838 3.4105
R16632 GNDA.n1055 GNDA.n848 3.4105
R16633 GNDA.n1057 GNDA.n848 3.4105
R16634 GNDA.n877 GNDA.n824 3.4105
R16635 GNDA.n877 GNDA.n825 3.4105
R16636 GNDA.n877 GNDA.n823 3.4105
R16637 GNDA.n877 GNDA.n826 3.4105
R16638 GNDA.n877 GNDA.n822 3.4105
R16639 GNDA.n877 GNDA.n827 3.4105
R16640 GNDA.n877 GNDA.n821 3.4105
R16641 GNDA.n877 GNDA.n828 3.4105
R16642 GNDA.n877 GNDA.n820 3.4105
R16643 GNDA.n877 GNDA.n829 3.4105
R16644 GNDA.n877 GNDA.n819 3.4105
R16645 GNDA.n877 GNDA.n830 3.4105
R16646 GNDA.n877 GNDA.n818 3.4105
R16647 GNDA.n877 GNDA.n831 3.4105
R16648 GNDA.n877 GNDA.n817 3.4105
R16649 GNDA.n877 GNDA.n832 3.4105
R16650 GNDA.n877 GNDA.n816 3.4105
R16651 GNDA.n877 GNDA.n833 3.4105
R16652 GNDA.n877 GNDA.n815 3.4105
R16653 GNDA.n877 GNDA.n834 3.4105
R16654 GNDA.n877 GNDA.n814 3.4105
R16655 GNDA.n877 GNDA.n835 3.4105
R16656 GNDA.n877 GNDA.n813 3.4105
R16657 GNDA.n877 GNDA.n836 3.4105
R16658 GNDA.n877 GNDA.n812 3.4105
R16659 GNDA.n877 GNDA.n837 3.4105
R16660 GNDA.n877 GNDA.n811 3.4105
R16661 GNDA.n877 GNDA.n838 3.4105
R16662 GNDA.n1055 GNDA.n877 3.4105
R16663 GNDA.n1057 GNDA.n877 3.4105
R16664 GNDA.n847 GNDA.n824 3.4105
R16665 GNDA.n847 GNDA.n825 3.4105
R16666 GNDA.n847 GNDA.n823 3.4105
R16667 GNDA.n847 GNDA.n826 3.4105
R16668 GNDA.n847 GNDA.n822 3.4105
R16669 GNDA.n847 GNDA.n827 3.4105
R16670 GNDA.n847 GNDA.n821 3.4105
R16671 GNDA.n847 GNDA.n828 3.4105
R16672 GNDA.n847 GNDA.n820 3.4105
R16673 GNDA.n847 GNDA.n829 3.4105
R16674 GNDA.n847 GNDA.n819 3.4105
R16675 GNDA.n847 GNDA.n830 3.4105
R16676 GNDA.n847 GNDA.n818 3.4105
R16677 GNDA.n847 GNDA.n831 3.4105
R16678 GNDA.n847 GNDA.n817 3.4105
R16679 GNDA.n847 GNDA.n832 3.4105
R16680 GNDA.n847 GNDA.n816 3.4105
R16681 GNDA.n847 GNDA.n833 3.4105
R16682 GNDA.n847 GNDA.n815 3.4105
R16683 GNDA.n847 GNDA.n834 3.4105
R16684 GNDA.n847 GNDA.n814 3.4105
R16685 GNDA.n847 GNDA.n835 3.4105
R16686 GNDA.n847 GNDA.n813 3.4105
R16687 GNDA.n847 GNDA.n836 3.4105
R16688 GNDA.n847 GNDA.n812 3.4105
R16689 GNDA.n847 GNDA.n837 3.4105
R16690 GNDA.n847 GNDA.n811 3.4105
R16691 GNDA.n847 GNDA.n838 3.4105
R16692 GNDA.n1055 GNDA.n847 3.4105
R16693 GNDA.n1057 GNDA.n847 3.4105
R16694 GNDA.n878 GNDA.n824 3.4105
R16695 GNDA.n878 GNDA.n825 3.4105
R16696 GNDA.n878 GNDA.n823 3.4105
R16697 GNDA.n878 GNDA.n826 3.4105
R16698 GNDA.n878 GNDA.n822 3.4105
R16699 GNDA.n878 GNDA.n827 3.4105
R16700 GNDA.n878 GNDA.n821 3.4105
R16701 GNDA.n878 GNDA.n828 3.4105
R16702 GNDA.n878 GNDA.n820 3.4105
R16703 GNDA.n878 GNDA.n829 3.4105
R16704 GNDA.n878 GNDA.n819 3.4105
R16705 GNDA.n878 GNDA.n830 3.4105
R16706 GNDA.n878 GNDA.n818 3.4105
R16707 GNDA.n878 GNDA.n831 3.4105
R16708 GNDA.n878 GNDA.n817 3.4105
R16709 GNDA.n878 GNDA.n832 3.4105
R16710 GNDA.n878 GNDA.n816 3.4105
R16711 GNDA.n878 GNDA.n833 3.4105
R16712 GNDA.n878 GNDA.n815 3.4105
R16713 GNDA.n878 GNDA.n834 3.4105
R16714 GNDA.n878 GNDA.n814 3.4105
R16715 GNDA.n878 GNDA.n835 3.4105
R16716 GNDA.n878 GNDA.n813 3.4105
R16717 GNDA.n878 GNDA.n836 3.4105
R16718 GNDA.n878 GNDA.n812 3.4105
R16719 GNDA.n878 GNDA.n837 3.4105
R16720 GNDA.n878 GNDA.n811 3.4105
R16721 GNDA.n878 GNDA.n838 3.4105
R16722 GNDA.n1055 GNDA.n878 3.4105
R16723 GNDA.n1057 GNDA.n878 3.4105
R16724 GNDA.n846 GNDA.n824 3.4105
R16725 GNDA.n846 GNDA.n825 3.4105
R16726 GNDA.n846 GNDA.n823 3.4105
R16727 GNDA.n846 GNDA.n826 3.4105
R16728 GNDA.n846 GNDA.n822 3.4105
R16729 GNDA.n846 GNDA.n827 3.4105
R16730 GNDA.n846 GNDA.n821 3.4105
R16731 GNDA.n846 GNDA.n828 3.4105
R16732 GNDA.n846 GNDA.n820 3.4105
R16733 GNDA.n846 GNDA.n829 3.4105
R16734 GNDA.n846 GNDA.n819 3.4105
R16735 GNDA.n846 GNDA.n830 3.4105
R16736 GNDA.n846 GNDA.n818 3.4105
R16737 GNDA.n846 GNDA.n831 3.4105
R16738 GNDA.n846 GNDA.n817 3.4105
R16739 GNDA.n846 GNDA.n832 3.4105
R16740 GNDA.n846 GNDA.n816 3.4105
R16741 GNDA.n846 GNDA.n833 3.4105
R16742 GNDA.n846 GNDA.n815 3.4105
R16743 GNDA.n846 GNDA.n834 3.4105
R16744 GNDA.n846 GNDA.n814 3.4105
R16745 GNDA.n846 GNDA.n835 3.4105
R16746 GNDA.n846 GNDA.n813 3.4105
R16747 GNDA.n846 GNDA.n836 3.4105
R16748 GNDA.n846 GNDA.n812 3.4105
R16749 GNDA.n846 GNDA.n837 3.4105
R16750 GNDA.n846 GNDA.n811 3.4105
R16751 GNDA.n846 GNDA.n838 3.4105
R16752 GNDA.n1055 GNDA.n846 3.4105
R16753 GNDA.n1057 GNDA.n846 3.4105
R16754 GNDA.n879 GNDA.n824 3.4105
R16755 GNDA.n879 GNDA.n825 3.4105
R16756 GNDA.n879 GNDA.n823 3.4105
R16757 GNDA.n879 GNDA.n826 3.4105
R16758 GNDA.n879 GNDA.n822 3.4105
R16759 GNDA.n879 GNDA.n827 3.4105
R16760 GNDA.n879 GNDA.n821 3.4105
R16761 GNDA.n879 GNDA.n828 3.4105
R16762 GNDA.n879 GNDA.n820 3.4105
R16763 GNDA.n879 GNDA.n829 3.4105
R16764 GNDA.n879 GNDA.n819 3.4105
R16765 GNDA.n879 GNDA.n830 3.4105
R16766 GNDA.n879 GNDA.n818 3.4105
R16767 GNDA.n879 GNDA.n831 3.4105
R16768 GNDA.n879 GNDA.n817 3.4105
R16769 GNDA.n879 GNDA.n832 3.4105
R16770 GNDA.n879 GNDA.n816 3.4105
R16771 GNDA.n879 GNDA.n833 3.4105
R16772 GNDA.n879 GNDA.n815 3.4105
R16773 GNDA.n879 GNDA.n834 3.4105
R16774 GNDA.n879 GNDA.n814 3.4105
R16775 GNDA.n879 GNDA.n835 3.4105
R16776 GNDA.n879 GNDA.n813 3.4105
R16777 GNDA.n879 GNDA.n836 3.4105
R16778 GNDA.n879 GNDA.n812 3.4105
R16779 GNDA.n879 GNDA.n837 3.4105
R16780 GNDA.n879 GNDA.n811 3.4105
R16781 GNDA.n879 GNDA.n838 3.4105
R16782 GNDA.n1055 GNDA.n879 3.4105
R16783 GNDA.n1057 GNDA.n879 3.4105
R16784 GNDA.n845 GNDA.n824 3.4105
R16785 GNDA.n845 GNDA.n825 3.4105
R16786 GNDA.n845 GNDA.n823 3.4105
R16787 GNDA.n845 GNDA.n826 3.4105
R16788 GNDA.n845 GNDA.n822 3.4105
R16789 GNDA.n845 GNDA.n827 3.4105
R16790 GNDA.n845 GNDA.n821 3.4105
R16791 GNDA.n845 GNDA.n828 3.4105
R16792 GNDA.n845 GNDA.n820 3.4105
R16793 GNDA.n845 GNDA.n829 3.4105
R16794 GNDA.n845 GNDA.n819 3.4105
R16795 GNDA.n845 GNDA.n830 3.4105
R16796 GNDA.n845 GNDA.n818 3.4105
R16797 GNDA.n845 GNDA.n831 3.4105
R16798 GNDA.n845 GNDA.n817 3.4105
R16799 GNDA.n845 GNDA.n832 3.4105
R16800 GNDA.n845 GNDA.n816 3.4105
R16801 GNDA.n845 GNDA.n833 3.4105
R16802 GNDA.n845 GNDA.n815 3.4105
R16803 GNDA.n845 GNDA.n834 3.4105
R16804 GNDA.n845 GNDA.n814 3.4105
R16805 GNDA.n845 GNDA.n835 3.4105
R16806 GNDA.n845 GNDA.n813 3.4105
R16807 GNDA.n845 GNDA.n836 3.4105
R16808 GNDA.n845 GNDA.n812 3.4105
R16809 GNDA.n845 GNDA.n837 3.4105
R16810 GNDA.n845 GNDA.n811 3.4105
R16811 GNDA.n845 GNDA.n838 3.4105
R16812 GNDA.n1055 GNDA.n845 3.4105
R16813 GNDA.n1057 GNDA.n845 3.4105
R16814 GNDA.n880 GNDA.n824 3.4105
R16815 GNDA.n880 GNDA.n825 3.4105
R16816 GNDA.n880 GNDA.n823 3.4105
R16817 GNDA.n880 GNDA.n826 3.4105
R16818 GNDA.n880 GNDA.n822 3.4105
R16819 GNDA.n880 GNDA.n827 3.4105
R16820 GNDA.n880 GNDA.n821 3.4105
R16821 GNDA.n880 GNDA.n828 3.4105
R16822 GNDA.n880 GNDA.n820 3.4105
R16823 GNDA.n880 GNDA.n829 3.4105
R16824 GNDA.n880 GNDA.n819 3.4105
R16825 GNDA.n880 GNDA.n830 3.4105
R16826 GNDA.n880 GNDA.n818 3.4105
R16827 GNDA.n880 GNDA.n831 3.4105
R16828 GNDA.n880 GNDA.n817 3.4105
R16829 GNDA.n880 GNDA.n832 3.4105
R16830 GNDA.n880 GNDA.n816 3.4105
R16831 GNDA.n880 GNDA.n833 3.4105
R16832 GNDA.n880 GNDA.n815 3.4105
R16833 GNDA.n880 GNDA.n834 3.4105
R16834 GNDA.n880 GNDA.n814 3.4105
R16835 GNDA.n880 GNDA.n835 3.4105
R16836 GNDA.n880 GNDA.n813 3.4105
R16837 GNDA.n880 GNDA.n836 3.4105
R16838 GNDA.n880 GNDA.n812 3.4105
R16839 GNDA.n880 GNDA.n837 3.4105
R16840 GNDA.n880 GNDA.n811 3.4105
R16841 GNDA.n880 GNDA.n838 3.4105
R16842 GNDA.n1055 GNDA.n880 3.4105
R16843 GNDA.n1057 GNDA.n880 3.4105
R16844 GNDA.n844 GNDA.n824 3.4105
R16845 GNDA.n844 GNDA.n825 3.4105
R16846 GNDA.n844 GNDA.n823 3.4105
R16847 GNDA.n844 GNDA.n826 3.4105
R16848 GNDA.n844 GNDA.n822 3.4105
R16849 GNDA.n844 GNDA.n827 3.4105
R16850 GNDA.n844 GNDA.n821 3.4105
R16851 GNDA.n844 GNDA.n828 3.4105
R16852 GNDA.n844 GNDA.n820 3.4105
R16853 GNDA.n844 GNDA.n829 3.4105
R16854 GNDA.n844 GNDA.n819 3.4105
R16855 GNDA.n844 GNDA.n830 3.4105
R16856 GNDA.n844 GNDA.n818 3.4105
R16857 GNDA.n844 GNDA.n831 3.4105
R16858 GNDA.n844 GNDA.n817 3.4105
R16859 GNDA.n844 GNDA.n832 3.4105
R16860 GNDA.n844 GNDA.n816 3.4105
R16861 GNDA.n844 GNDA.n833 3.4105
R16862 GNDA.n844 GNDA.n815 3.4105
R16863 GNDA.n844 GNDA.n834 3.4105
R16864 GNDA.n844 GNDA.n814 3.4105
R16865 GNDA.n844 GNDA.n835 3.4105
R16866 GNDA.n844 GNDA.n813 3.4105
R16867 GNDA.n844 GNDA.n836 3.4105
R16868 GNDA.n844 GNDA.n812 3.4105
R16869 GNDA.n844 GNDA.n837 3.4105
R16870 GNDA.n844 GNDA.n811 3.4105
R16871 GNDA.n844 GNDA.n838 3.4105
R16872 GNDA.n1055 GNDA.n844 3.4105
R16873 GNDA.n1057 GNDA.n844 3.4105
R16874 GNDA.n881 GNDA.n824 3.4105
R16875 GNDA.n881 GNDA.n825 3.4105
R16876 GNDA.n881 GNDA.n823 3.4105
R16877 GNDA.n881 GNDA.n826 3.4105
R16878 GNDA.n881 GNDA.n822 3.4105
R16879 GNDA.n881 GNDA.n827 3.4105
R16880 GNDA.n881 GNDA.n821 3.4105
R16881 GNDA.n881 GNDA.n828 3.4105
R16882 GNDA.n881 GNDA.n820 3.4105
R16883 GNDA.n881 GNDA.n829 3.4105
R16884 GNDA.n881 GNDA.n819 3.4105
R16885 GNDA.n881 GNDA.n830 3.4105
R16886 GNDA.n881 GNDA.n818 3.4105
R16887 GNDA.n881 GNDA.n831 3.4105
R16888 GNDA.n881 GNDA.n817 3.4105
R16889 GNDA.n881 GNDA.n832 3.4105
R16890 GNDA.n881 GNDA.n816 3.4105
R16891 GNDA.n881 GNDA.n833 3.4105
R16892 GNDA.n881 GNDA.n815 3.4105
R16893 GNDA.n881 GNDA.n834 3.4105
R16894 GNDA.n881 GNDA.n814 3.4105
R16895 GNDA.n881 GNDA.n835 3.4105
R16896 GNDA.n881 GNDA.n813 3.4105
R16897 GNDA.n881 GNDA.n836 3.4105
R16898 GNDA.n881 GNDA.n812 3.4105
R16899 GNDA.n881 GNDA.n837 3.4105
R16900 GNDA.n881 GNDA.n811 3.4105
R16901 GNDA.n881 GNDA.n838 3.4105
R16902 GNDA.n1055 GNDA.n881 3.4105
R16903 GNDA.n1057 GNDA.n881 3.4105
R16904 GNDA.n843 GNDA.n824 3.4105
R16905 GNDA.n843 GNDA.n825 3.4105
R16906 GNDA.n843 GNDA.n823 3.4105
R16907 GNDA.n843 GNDA.n826 3.4105
R16908 GNDA.n843 GNDA.n822 3.4105
R16909 GNDA.n843 GNDA.n827 3.4105
R16910 GNDA.n843 GNDA.n821 3.4105
R16911 GNDA.n843 GNDA.n828 3.4105
R16912 GNDA.n843 GNDA.n820 3.4105
R16913 GNDA.n843 GNDA.n829 3.4105
R16914 GNDA.n843 GNDA.n819 3.4105
R16915 GNDA.n843 GNDA.n830 3.4105
R16916 GNDA.n843 GNDA.n818 3.4105
R16917 GNDA.n843 GNDA.n831 3.4105
R16918 GNDA.n843 GNDA.n817 3.4105
R16919 GNDA.n843 GNDA.n832 3.4105
R16920 GNDA.n843 GNDA.n816 3.4105
R16921 GNDA.n843 GNDA.n833 3.4105
R16922 GNDA.n843 GNDA.n815 3.4105
R16923 GNDA.n843 GNDA.n834 3.4105
R16924 GNDA.n843 GNDA.n814 3.4105
R16925 GNDA.n843 GNDA.n835 3.4105
R16926 GNDA.n843 GNDA.n813 3.4105
R16927 GNDA.n843 GNDA.n836 3.4105
R16928 GNDA.n843 GNDA.n812 3.4105
R16929 GNDA.n843 GNDA.n837 3.4105
R16930 GNDA.n843 GNDA.n811 3.4105
R16931 GNDA.n843 GNDA.n838 3.4105
R16932 GNDA.n1055 GNDA.n843 3.4105
R16933 GNDA.n1057 GNDA.n843 3.4105
R16934 GNDA.n882 GNDA.n824 3.4105
R16935 GNDA.n882 GNDA.n825 3.4105
R16936 GNDA.n882 GNDA.n823 3.4105
R16937 GNDA.n882 GNDA.n826 3.4105
R16938 GNDA.n882 GNDA.n822 3.4105
R16939 GNDA.n882 GNDA.n827 3.4105
R16940 GNDA.n882 GNDA.n821 3.4105
R16941 GNDA.n882 GNDA.n828 3.4105
R16942 GNDA.n882 GNDA.n820 3.4105
R16943 GNDA.n882 GNDA.n829 3.4105
R16944 GNDA.n882 GNDA.n819 3.4105
R16945 GNDA.n882 GNDA.n830 3.4105
R16946 GNDA.n882 GNDA.n818 3.4105
R16947 GNDA.n882 GNDA.n831 3.4105
R16948 GNDA.n882 GNDA.n817 3.4105
R16949 GNDA.n882 GNDA.n832 3.4105
R16950 GNDA.n882 GNDA.n816 3.4105
R16951 GNDA.n882 GNDA.n833 3.4105
R16952 GNDA.n882 GNDA.n815 3.4105
R16953 GNDA.n882 GNDA.n834 3.4105
R16954 GNDA.n882 GNDA.n814 3.4105
R16955 GNDA.n882 GNDA.n835 3.4105
R16956 GNDA.n882 GNDA.n813 3.4105
R16957 GNDA.n882 GNDA.n836 3.4105
R16958 GNDA.n882 GNDA.n812 3.4105
R16959 GNDA.n882 GNDA.n837 3.4105
R16960 GNDA.n882 GNDA.n811 3.4105
R16961 GNDA.n882 GNDA.n838 3.4105
R16962 GNDA.n1055 GNDA.n882 3.4105
R16963 GNDA.n1057 GNDA.n882 3.4105
R16964 GNDA.n842 GNDA.n824 3.4105
R16965 GNDA.n842 GNDA.n825 3.4105
R16966 GNDA.n842 GNDA.n823 3.4105
R16967 GNDA.n842 GNDA.n826 3.4105
R16968 GNDA.n842 GNDA.n822 3.4105
R16969 GNDA.n842 GNDA.n827 3.4105
R16970 GNDA.n842 GNDA.n821 3.4105
R16971 GNDA.n842 GNDA.n828 3.4105
R16972 GNDA.n842 GNDA.n820 3.4105
R16973 GNDA.n842 GNDA.n829 3.4105
R16974 GNDA.n842 GNDA.n819 3.4105
R16975 GNDA.n842 GNDA.n830 3.4105
R16976 GNDA.n842 GNDA.n818 3.4105
R16977 GNDA.n842 GNDA.n831 3.4105
R16978 GNDA.n842 GNDA.n817 3.4105
R16979 GNDA.n842 GNDA.n832 3.4105
R16980 GNDA.n842 GNDA.n816 3.4105
R16981 GNDA.n842 GNDA.n833 3.4105
R16982 GNDA.n842 GNDA.n815 3.4105
R16983 GNDA.n842 GNDA.n834 3.4105
R16984 GNDA.n842 GNDA.n814 3.4105
R16985 GNDA.n842 GNDA.n835 3.4105
R16986 GNDA.n842 GNDA.n813 3.4105
R16987 GNDA.n842 GNDA.n836 3.4105
R16988 GNDA.n842 GNDA.n812 3.4105
R16989 GNDA.n842 GNDA.n837 3.4105
R16990 GNDA.n842 GNDA.n811 3.4105
R16991 GNDA.n842 GNDA.n838 3.4105
R16992 GNDA.n1055 GNDA.n842 3.4105
R16993 GNDA.n1057 GNDA.n842 3.4105
R16994 GNDA.n883 GNDA.n824 3.4105
R16995 GNDA.n883 GNDA.n825 3.4105
R16996 GNDA.n883 GNDA.n823 3.4105
R16997 GNDA.n883 GNDA.n826 3.4105
R16998 GNDA.n883 GNDA.n822 3.4105
R16999 GNDA.n883 GNDA.n827 3.4105
R17000 GNDA.n883 GNDA.n821 3.4105
R17001 GNDA.n883 GNDA.n828 3.4105
R17002 GNDA.n883 GNDA.n820 3.4105
R17003 GNDA.n883 GNDA.n829 3.4105
R17004 GNDA.n883 GNDA.n819 3.4105
R17005 GNDA.n883 GNDA.n830 3.4105
R17006 GNDA.n883 GNDA.n818 3.4105
R17007 GNDA.n883 GNDA.n831 3.4105
R17008 GNDA.n883 GNDA.n817 3.4105
R17009 GNDA.n883 GNDA.n832 3.4105
R17010 GNDA.n883 GNDA.n816 3.4105
R17011 GNDA.n883 GNDA.n833 3.4105
R17012 GNDA.n883 GNDA.n815 3.4105
R17013 GNDA.n883 GNDA.n834 3.4105
R17014 GNDA.n883 GNDA.n814 3.4105
R17015 GNDA.n883 GNDA.n835 3.4105
R17016 GNDA.n883 GNDA.n813 3.4105
R17017 GNDA.n883 GNDA.n836 3.4105
R17018 GNDA.n883 GNDA.n812 3.4105
R17019 GNDA.n883 GNDA.n837 3.4105
R17020 GNDA.n883 GNDA.n811 3.4105
R17021 GNDA.n883 GNDA.n838 3.4105
R17022 GNDA.n1055 GNDA.n883 3.4105
R17023 GNDA.n1057 GNDA.n883 3.4105
R17024 GNDA.n841 GNDA.n824 3.4105
R17025 GNDA.n841 GNDA.n825 3.4105
R17026 GNDA.n841 GNDA.n823 3.4105
R17027 GNDA.n841 GNDA.n826 3.4105
R17028 GNDA.n841 GNDA.n822 3.4105
R17029 GNDA.n841 GNDA.n827 3.4105
R17030 GNDA.n841 GNDA.n821 3.4105
R17031 GNDA.n841 GNDA.n828 3.4105
R17032 GNDA.n841 GNDA.n820 3.4105
R17033 GNDA.n841 GNDA.n829 3.4105
R17034 GNDA.n841 GNDA.n819 3.4105
R17035 GNDA.n841 GNDA.n830 3.4105
R17036 GNDA.n841 GNDA.n818 3.4105
R17037 GNDA.n841 GNDA.n831 3.4105
R17038 GNDA.n841 GNDA.n817 3.4105
R17039 GNDA.n841 GNDA.n832 3.4105
R17040 GNDA.n841 GNDA.n816 3.4105
R17041 GNDA.n841 GNDA.n833 3.4105
R17042 GNDA.n841 GNDA.n815 3.4105
R17043 GNDA.n841 GNDA.n834 3.4105
R17044 GNDA.n841 GNDA.n814 3.4105
R17045 GNDA.n841 GNDA.n835 3.4105
R17046 GNDA.n841 GNDA.n813 3.4105
R17047 GNDA.n841 GNDA.n836 3.4105
R17048 GNDA.n841 GNDA.n812 3.4105
R17049 GNDA.n841 GNDA.n837 3.4105
R17050 GNDA.n841 GNDA.n811 3.4105
R17051 GNDA.n841 GNDA.n838 3.4105
R17052 GNDA.n1055 GNDA.n841 3.4105
R17053 GNDA.n1057 GNDA.n841 3.4105
R17054 GNDA.n1056 GNDA.n824 3.4105
R17055 GNDA.n1056 GNDA.n825 3.4105
R17056 GNDA.n1056 GNDA.n823 3.4105
R17057 GNDA.n1056 GNDA.n826 3.4105
R17058 GNDA.n1056 GNDA.n822 3.4105
R17059 GNDA.n1056 GNDA.n827 3.4105
R17060 GNDA.n1056 GNDA.n821 3.4105
R17061 GNDA.n1056 GNDA.n828 3.4105
R17062 GNDA.n1056 GNDA.n820 3.4105
R17063 GNDA.n1056 GNDA.n829 3.4105
R17064 GNDA.n1056 GNDA.n819 3.4105
R17065 GNDA.n1056 GNDA.n830 3.4105
R17066 GNDA.n1056 GNDA.n818 3.4105
R17067 GNDA.n1056 GNDA.n831 3.4105
R17068 GNDA.n1056 GNDA.n817 3.4105
R17069 GNDA.n1056 GNDA.n832 3.4105
R17070 GNDA.n1056 GNDA.n816 3.4105
R17071 GNDA.n1056 GNDA.n833 3.4105
R17072 GNDA.n1056 GNDA.n815 3.4105
R17073 GNDA.n1056 GNDA.n834 3.4105
R17074 GNDA.n1056 GNDA.n814 3.4105
R17075 GNDA.n1056 GNDA.n835 3.4105
R17076 GNDA.n1056 GNDA.n813 3.4105
R17077 GNDA.n1056 GNDA.n836 3.4105
R17078 GNDA.n1056 GNDA.n812 3.4105
R17079 GNDA.n1056 GNDA.n837 3.4105
R17080 GNDA.n1056 GNDA.n811 3.4105
R17081 GNDA.n1056 GNDA.n838 3.4105
R17082 GNDA.n1056 GNDA.n1055 3.4105
R17083 GNDA.n1057 GNDA.n1056 3.4105
R17084 GNDA.n840 GNDA.n824 3.4105
R17085 GNDA.n840 GNDA.n825 3.4105
R17086 GNDA.n840 GNDA.n823 3.4105
R17087 GNDA.n840 GNDA.n826 3.4105
R17088 GNDA.n840 GNDA.n822 3.4105
R17089 GNDA.n840 GNDA.n827 3.4105
R17090 GNDA.n840 GNDA.n821 3.4105
R17091 GNDA.n840 GNDA.n828 3.4105
R17092 GNDA.n840 GNDA.n820 3.4105
R17093 GNDA.n840 GNDA.n829 3.4105
R17094 GNDA.n840 GNDA.n819 3.4105
R17095 GNDA.n840 GNDA.n830 3.4105
R17096 GNDA.n840 GNDA.n818 3.4105
R17097 GNDA.n840 GNDA.n831 3.4105
R17098 GNDA.n840 GNDA.n817 3.4105
R17099 GNDA.n840 GNDA.n832 3.4105
R17100 GNDA.n840 GNDA.n816 3.4105
R17101 GNDA.n840 GNDA.n833 3.4105
R17102 GNDA.n840 GNDA.n815 3.4105
R17103 GNDA.n840 GNDA.n834 3.4105
R17104 GNDA.n840 GNDA.n814 3.4105
R17105 GNDA.n840 GNDA.n835 3.4105
R17106 GNDA.n840 GNDA.n813 3.4105
R17107 GNDA.n840 GNDA.n836 3.4105
R17108 GNDA.n840 GNDA.n812 3.4105
R17109 GNDA.n840 GNDA.n837 3.4105
R17110 GNDA.n840 GNDA.n811 3.4105
R17111 GNDA.n840 GNDA.n838 3.4105
R17112 GNDA.n1055 GNDA.n840 3.4105
R17113 GNDA.n1057 GNDA.n840 3.4105
R17114 GNDA.n1058 GNDA.n824 3.4105
R17115 GNDA.n1058 GNDA.n825 3.4105
R17116 GNDA.n1058 GNDA.n823 3.4105
R17117 GNDA.n1058 GNDA.n826 3.4105
R17118 GNDA.n1058 GNDA.n822 3.4105
R17119 GNDA.n1058 GNDA.n827 3.4105
R17120 GNDA.n1058 GNDA.n821 3.4105
R17121 GNDA.n1058 GNDA.n828 3.4105
R17122 GNDA.n1058 GNDA.n820 3.4105
R17123 GNDA.n1058 GNDA.n829 3.4105
R17124 GNDA.n1058 GNDA.n819 3.4105
R17125 GNDA.n1058 GNDA.n830 3.4105
R17126 GNDA.n1058 GNDA.n818 3.4105
R17127 GNDA.n1058 GNDA.n831 3.4105
R17128 GNDA.n1058 GNDA.n817 3.4105
R17129 GNDA.n1058 GNDA.n832 3.4105
R17130 GNDA.n1058 GNDA.n816 3.4105
R17131 GNDA.n1058 GNDA.n833 3.4105
R17132 GNDA.n1058 GNDA.n815 3.4105
R17133 GNDA.n1058 GNDA.n834 3.4105
R17134 GNDA.n1058 GNDA.n814 3.4105
R17135 GNDA.n1058 GNDA.n835 3.4105
R17136 GNDA.n1058 GNDA.n813 3.4105
R17137 GNDA.n1058 GNDA.n836 3.4105
R17138 GNDA.n1058 GNDA.n812 3.4105
R17139 GNDA.n1058 GNDA.n837 3.4105
R17140 GNDA.n1058 GNDA.n811 3.4105
R17141 GNDA.n1058 GNDA.n838 3.4105
R17142 GNDA.n1058 GNDA.n1057 3.4105
R17143 GNDA.n1734 GNDA.n1733 3.39217
R17144 GNDA.n1741 GNDA.n1740 3.39217
R17145 GNDA.n3392 GNDA.n3391 3.39217
R17146 GNDA.n3382 GNDA.n3381 3.39217
R17147 GNDA.n6813 GNDA.n6648 3.22552
R17148 GNDA.n6958 GNDA.n6957 3.22552
R17149 GNDA.n6746 GNDA.t0 3.22552
R17150 GNDA.t29 GNDA.n286 3.22552
R17151 GNDA.n3387 GNDA.n3384 3.13621
R17152 GNDA.n3388 GNDA.n3387 3.13621
R17153 GNDA.n1729 GNDA.n1725 3.13621
R17154 GNDA.n1730 GNDA.n1729 3.13621
R17155 GNDA.n7232 GNDA.n93 3.007
R17156 GNDA.n6770 GNDA.n6663 2.86505
R17157 GNDA.n6771 GNDA.n6770 2.86505
R17158 GNDA.n6769 GNDA.n6765 2.86505
R17159 GNDA.n6766 GNDA.n6765 2.86505
R17160 GNDA.n6772 GNDA.n6771 2.86505
R17161 GNDA.n6767 GNDA.n6766 2.86505
R17162 GNDA.n6776 GNDA.n6663 2.86505
R17163 GNDA.n6772 GNDA.n6769 2.86505
R17164 GNDA.n6789 GNDA.n6788 2.86505
R17165 GNDA.n6788 GNDA.n6786 2.86505
R17166 GNDA.n6786 GNDA.n6785 2.86505
R17167 GNDA.n6790 GNDA.n6789 2.86505
R17168 GNDA.n7056 GNDA.n7054 2.68279
R17169 GNDA.n6450 GNDA.n6449 2.6629
R17170 GNDA.n7477 GNDA.n7476 2.6629
R17171 GNDA.n6545 GNDA.n6544 2.6629
R17172 GNDA.n6453 GNDA.n6451 2.6629
R17173 GNDA.n6904 GNDA.n6903 2.6629
R17174 GNDA.n6934 GNDA.n6933 2.6629
R17175 GNDA.n6822 GNDA.n6821 2.6629
R17176 GNDA.n6906 GNDA.n6905 2.6629
R17177 GNDA.n5717 GNDA.n5716 2.6629
R17178 GNDA.n6067 GNDA.n6066 2.6629
R17179 GNDA.n5476 GNDA.n5442 2.6629
R17180 GNDA.n5996 GNDA.n5995 2.6629
R17181 GNDA.n5909 GNDA.n5450 2.6629
R17182 GNDA.n6739 GNDA.n5369 2.6629
R17183 GNDA.n7317 GNDA.n58 2.6629
R17184 GNDA.n7062 GNDA.n7061 2.56821
R17185 GNDA.n7229 GNDA.n7228 2.45883
R17186 GNDA.n6451 GNDA.n6450 2.4581
R17187 GNDA.n7478 GNDA.n7477 2.4581
R17188 GNDA.n6454 GNDA.n6453 2.4581
R17189 GNDA.n6905 GNDA.n6904 2.4581
R17190 GNDA.n6934 GNDA.n5368 2.4581
R17191 GNDA.n6907 GNDA.n6906 2.4581
R17192 GNDA.n5716 GNDA.n5442 2.4581
R17193 GNDA.n5754 GNDA.n5753 2.4581
R17194 GNDA.n6067 GNDA.n5450 2.4581
R17195 GNDA.n5476 GNDA.n5473 2.4581
R17196 GNDA.n5910 GNDA.n5909 2.4581
R17197 GNDA.n6933 GNDA.n5369 2.4581
R17198 GNDA.n6684 GNDA.n307 2.4581
R17199 GNDA.n7476 GNDA.n58 2.4581
R17200 GNDA.n7384 GNDA.n7383 2.4581
R17201 GNDA.n6999 GNDA.n6998 2.44675
R17202 GNDA.n6998 GNDA.n6997 2.44675
R17203 GNDA.n150 GNDA.n149 2.39683
R17204 GNDA.n4999 GNDA.n4998 2.38247
R17205 GNDA.n5005 GNDA.n5004 2.38247
R17206 GNDA.n660 GNDA.n659 2.38247
R17207 GNDA.n2109 GNDA.n2108 2.38212
R17208 GNDA.n7132 GNDA.n7131 2.30736
R17209 GNDA.n5270 GNDA.n5269 2.30736
R17210 GNDA.n4957 GNDA.n4956 2.30736
R17211 GNDA.n4797 GNDA.n4796 2.30736
R17212 GNDA.n4631 GNDA.n4630 2.30736
R17213 GNDA.n4465 GNDA.n4464 2.30736
R17214 GNDA.n4299 GNDA.n4298 2.30736
R17215 GNDA.n3801 GNDA.n3800 2.30736
R17216 GNDA.n4133 GNDA.n4132 2.30736
R17217 GNDA.n3967 GNDA.n3966 2.30736
R17218 GNDA.n3602 GNDA.n3601 2.30736
R17219 GNDA.n496 GNDA.n495 2.30736
R17220 GNDA.n5133 GNDA.n5132 2.30736
R17221 GNDA.n3299 GNDA.n3298 2.30736
R17222 GNDA.n3195 GNDA.n3194 2.30736
R17223 GNDA.n3035 GNDA.n3034 2.30736
R17224 GNDA.n2399 GNDA.n2398 2.30736
R17225 GNDA.n2861 GNDA.n2860 2.30736
R17226 GNDA.n2662 GNDA.n2661 2.30736
R17227 GNDA.n2559 GNDA.n2558 2.30736
R17228 GNDA.n2202 GNDA.n2201 2.30736
R17229 GNDA.n2096 GNDA.n2095 2.30736
R17230 GNDA.n1936 GNDA.n1935 2.30736
R17231 GNDA.n1615 GNDA.n1614 2.30736
R17232 GNDA.n1512 GNDA.n1511 2.30736
R17233 GNDA.n1350 GNDA.n1349 2.30736
R17234 GNDA.n3404 GNDA.n3403 2.29914
R17235 GNDA.n3401 GNDA.n3400 2.29914
R17236 GNDA.n5314 GNDA.n5313 2.29914
R17237 GNDA.n5316 GNDA.n5315 2.29914
R17238 GNDA.n1762 GNDA.n1711 2.26187
R17239 GNDA.n1759 GNDA.n1758 2.26187
R17240 GNDA.n1780 GNDA.n1705 2.26187
R17241 GNDA.n1723 GNDA.n1719 2.26187
R17242 GNDA.n1803 GNDA.n1698 2.26187
R17243 GNDA.n1809 GNDA.n1696 2.26187
R17244 GNDA.n4988 GNDA.n3432 2.26187
R17245 GNDA.n5357 GNDA.n5353 2.26187
R17246 GNDA.n6658 GNDA.n6655 2.26187
R17247 GNDA.n7055 GNDA.n261 2.26187
R17248 GNDA.n267 GNDA.n264 2.26187
R17249 GNDA.n268 GNDA.n267 2.26187
R17250 GNDA.n3420 GNDA.n3407 2.26187
R17251 GNDA.n3421 GNDA.n3420 2.26187
R17252 GNDA.n1760 GNDA.n1759 2.26187
R17253 GNDA.n1765 GNDA.n1764 2.26187
R17254 GNDA.n1768 GNDA.n1709 2.26187
R17255 GNDA.n1777 GNDA.n1705 2.26187
R17256 GNDA.n1800 GNDA.n1698 2.26187
R17257 GNDA.n1224 GNDA.n1221 2.26187
R17258 GNDA.n1229 GNDA.n1218 2.26187
R17259 GNDA.n1236 GNDA.n1235 2.26187
R17260 GNDA.n6659 GNDA.n6658 2.26187
R17261 GNDA.n6780 GNDA.n6779 2.26187
R17262 GNDA.t195 GNDA.t145 2.25277
R17263 GNDA.n2280 GNDA.n717 2.24241
R17264 GNDA.n719 GNDA.n716 2.24241
R17265 GNDA.n3684 GNDA.n576 2.24241
R17266 GNDA.n3510 GNDA.n3509 2.24241
R17267 GNDA.n3424 GNDA.n3419 2.24063
R17268 GNDA.n3425 GNDA.n3407 2.24063
R17269 GNDA.n3426 GNDA.n589 2.24063
R17270 GNDA.n3406 GNDA.n588 2.24063
R17271 GNDA.n1764 GNDA.n1763 2.24063
R17272 GNDA.n1758 GNDA.n1757 2.24063
R17273 GNDA.n1769 GNDA.n1768 2.24063
R17274 GNDA.n1767 GNDA.n1710 2.24063
R17275 GNDA.n1781 GNDA.n1704 2.24063
R17276 GNDA.n1724 GNDA.n1723 2.24063
R17277 GNDA.n1720 GNDA.n1718 2.24063
R17278 GNDA.n1784 GNDA.n1783 2.24063
R17279 GNDA.n1703 GNDA.n1701 2.24063
R17280 GNDA.n1804 GNDA.n1697 2.24063
R17281 GNDA.n1810 GNDA.n1695 2.24063
R17282 GNDA.n1227 GNDA.n1221 2.24063
R17283 GNDA.n1222 GNDA.n1220 2.24063
R17284 GNDA.n1232 GNDA.n1218 2.24063
R17285 GNDA.n1219 GNDA.n1217 2.24063
R17286 GNDA.n1235 GNDA.n789 2.24063
R17287 GNDA.n1234 GNDA.n1216 2.24063
R17288 GNDA.n1522 GNDA.n787 2.24063
R17289 GNDA.n788 GNDA.n786 2.24063
R17290 GNDA.n1519 GNDA.n1518 2.24063
R17291 GNDA.n1693 GNDA.n784 2.24063
R17292 GNDA.n785 GNDA.n783 2.24063
R17293 GNDA.n1690 GNDA.n1689 2.24063
R17294 GNDA.n1819 GNDA.n723 2.24063
R17295 GNDA.n779 GNDA.n778 2.24063
R17296 GNDA.n1820 GNDA.n777 2.24063
R17297 GNDA.n2106 GNDA.n721 2.24063
R17298 GNDA.n722 GNDA.n720 2.24063
R17299 GNDA.n2103 GNDA.n2102 2.24063
R17300 GNDA.n2277 GNDA.n2276 2.24063
R17301 GNDA.n2569 GNDA.n656 2.24063
R17302 GNDA.n657 GNDA.n655 2.24063
R17303 GNDA.n2566 GNDA.n2565 2.24063
R17304 GNDA.n2740 GNDA.n653 2.24063
R17305 GNDA.n654 GNDA.n652 2.24063
R17306 GNDA.n2737 GNDA.n2736 2.24063
R17307 GNDA.n2744 GNDA.n649 2.24063
R17308 GNDA.n651 GNDA.n650 2.24063
R17309 GNDA.n2745 GNDA.n648 2.24063
R17310 GNDA.n2918 GNDA.n594 2.24063
R17311 GNDA.n2914 GNDA.n2913 2.24063
R17312 GNDA.n2919 GNDA.n2912 2.24063
R17313 GNDA.n3205 GNDA.n592 2.24063
R17314 GNDA.n593 GNDA.n591 2.24063
R17315 GNDA.n3202 GNDA.n3201 2.24063
R17316 GNDA.n3376 GNDA.n3375 2.24063
R17317 GNDA.n3377 GNDA.n3374 2.24063
R17318 GNDA.n3378 GNDA.n3373 2.24063
R17319 GNDA.n5016 GNDA.n5010 2.24063
R17320 GNDA.n5012 GNDA.n5011 2.24063
R17321 GNDA.n5017 GNDA.n402 2.24063
R17322 GNDA.n5006 GNDA.n572 2.24063
R17323 GNDA.n5007 GNDA.n571 2.24063
R17324 GNDA.n5008 GNDA.n570 2.24063
R17325 GNDA.n4994 GNDA.n581 2.24063
R17326 GNDA.n4995 GNDA.n580 2.24063
R17327 GNDA.n4996 GNDA.n579 2.24063
R17328 GNDA.n4990 GNDA.n586 2.24063
R17329 GNDA.n4991 GNDA.n585 2.24063
R17330 GNDA.n4992 GNDA.n584 2.24063
R17331 GNDA.n3685 GNDA.n3508 2.24063
R17332 GNDA.n4982 GNDA.n3438 2.24063
R17333 GNDA.n4983 GNDA.n3437 2.24063
R17334 GNDA.n4984 GNDA.n3436 2.24063
R17335 GNDA.n4978 GNDA.n3443 2.24063
R17336 GNDA.n4979 GNDA.n3442 2.24063
R17337 GNDA.n4980 GNDA.n3441 2.24063
R17338 GNDA.n4974 GNDA.n3448 2.24063
R17339 GNDA.n4975 GNDA.n3447 2.24063
R17340 GNDA.n4976 GNDA.n3446 2.24063
R17341 GNDA.n4970 GNDA.n3453 2.24063
R17342 GNDA.n4971 GNDA.n3452 2.24063
R17343 GNDA.n4972 GNDA.n3451 2.24063
R17344 GNDA.n4966 GNDA.n4965 2.24063
R17345 GNDA.n4967 GNDA.n4964 2.24063
R17346 GNDA.n4968 GNDA.n4963 2.24063
R17347 GNDA.n1815 GNDA.n781 2.24063
R17348 GNDA.n782 GNDA.n780 2.24063
R17349 GNDA.n4986 GNDA.n3432 2.24063
R17350 GNDA.n4987 GNDA.n3433 2.24063
R17351 GNDA.n5276 GNDA.n323 2.24063
R17352 GNDA.n5278 GNDA.n322 2.24063
R17353 GNDA.n5279 GNDA.n5277 2.24063
R17354 GNDA.n6948 GNDA.n5353 2.24063
R17355 GNDA.n6779 GNDA.n6778 2.24063
R17356 GNDA.n6654 GNDA.n6653 2.24063
R17357 GNDA.n6662 GNDA.n6655 2.24063
R17358 GNDA.n7231 GNDA.n7230 2.24063
R17359 GNDA.n94 GNDA.n92 2.24063
R17360 GNDA.n7057 GNDA.n7056 2.24063
R17361 GNDA.n3428 GNDA.n3427 2.24063
R17362 GNDA.n1766 GNDA.n1711 2.24063
R17363 GNDA.n1761 GNDA.n1714 2.24063
R17364 GNDA.n1777 GNDA.n1776 2.24063
R17365 GNDA.n1782 GNDA.n1700 2.24063
R17366 GNDA.n1800 GNDA.n1799 2.24063
R17367 GNDA.n1805 GNDA.n1696 2.24063
R17368 GNDA.n1806 GNDA.n317 2.24063
R17369 GNDA.n1812 GNDA.n1811 2.24063
R17370 GNDA.n6947 GNDA.n6946 2.24063
R17371 GNDA.n6945 GNDA.n6944 2.24063
R17372 GNDA.n6661 GNDA.n6660 2.24063
R17373 GNDA.n7229 GNDA.n91 2.24063
R17374 GNDA.n7061 GNDA.n261 2.24063
R17375 GNDA.n7060 GNDA.n7059 2.24063
R17376 GNDA.n7054 GNDA.n264 2.24063
R17377 GNDA.n7053 GNDA.n7052 2.24063
R17378 GNDA.n5282 GNDA.n5281 2.24008
R17379 GNDA.n6949 GNDA.n5351 2.22018
R17380 GNDA.n6943 GNDA.n5358 2.22018
R17381 GNDA.n1735 GNDA.n1707 2.19633
R17382 GNDA.n1738 GNDA.n1706 2.19633
R17383 GNDA.n5306 GNDA.n5305 2.19633
R17384 GNDA.n6451 GNDA.n67 2.18124
R17385 GNDA.n6905 GNDA.n5389 2.18124
R17386 GNDA.n5550 GNDA.n5450 2.18124
R17387 GNDA.n7476 GNDA.n59 2.18124
R17388 GNDA.n5601 GNDA.n5442 2.18124
R17389 GNDA.n6933 GNDA.n5370 2.18124
R17390 GNDA.n3386 GNDA.n590 2.15331
R17391 GNDA.n1728 GNDA.n1726 2.15331
R17392 GNDA.n7479 GNDA.n7478 2.1509
R17393 GNDA.n6480 GNDA.n6454 2.1509
R17394 GNDA.n6847 GNDA.n5368 2.1509
R17395 GNDA.n6908 GNDA.n6907 2.1509
R17396 GNDA.n5753 GNDA.n5752 2.1509
R17397 GNDA.n6002 GNDA.n5473 2.1509
R17398 GNDA.n5928 GNDA.n5910 2.1509
R17399 GNDA.n6684 GNDA.n291 2.1509
R17400 GNDA.n7383 GNDA.n7382 2.1509
R17401 GNDA.n6544 GNDA.n6323 2.13383
R17402 GNDA.n6449 GNDA.n6344 2.13383
R17403 GNDA.n6903 GNDA.n6902 2.13383
R17404 GNDA.n6821 GNDA.n6575 2.13383
R17405 GNDA.n5717 GNDA.n5715 2.13383
R17406 GNDA.n6066 GNDA.n5451 2.13383
R17407 GNDA.n5995 GNDA.n5883 2.13383
R17408 GNDA.n6739 GNDA.n6738 2.13383
R17409 GNDA.n7318 GNDA.n7317 2.13383
R17410 GNDA.n5000 GNDA.n4999 2.09414
R17411 GNDA.n5004 GNDA.n5003 2.09414
R17412 GNDA.n659 GNDA.n658 2.09414
R17413 GNDA.n2108 GNDA.n2107 2.09414
R17414 GNDA.n6451 GNDA.n65 2.08643
R17415 GNDA.n6905 GNDA.n5387 2.08643
R17416 GNDA.n5450 GNDA.n5435 2.08643
R17417 GNDA.n7476 GNDA.n7475 2.08643
R17418 GNDA.n6072 GNDA.n5442 2.08643
R17419 GNDA.n6933 GNDA.n6932 2.08643
R17420 GNDA.n3391 GNDA.n324 2.00747
R17421 GNDA.n3381 GNDA.n3380 2.00747
R17422 GNDA.n6449 GNDA.n6448 1.9461
R17423 GNDA.n6544 GNDA.n6543 1.9461
R17424 GNDA.n6903 GNDA.n5344 1.9461
R17425 GNDA.n6821 GNDA.n6820 1.9461
R17426 GNDA.n5718 GNDA.n5717 1.9461
R17427 GNDA.n6066 GNDA.n6065 1.9461
R17428 GNDA.n5995 GNDA.n5994 1.9461
R17429 GNDA.n6741 GNDA.n6739 1.9461
R17430 GNDA.n7317 GNDA.n22 1.9461
R17431 GNDA.n3403 GNDA.n3402 1.93383
R17432 GNDA.n3400 GNDA.n3399 1.93383
R17433 GNDA.n5313 GNDA.n5312 1.93383
R17434 GNDA.n5317 GNDA.n5316 1.93383
R17435 GNDA.n5282 GNDA.n321 1.91062
R17436 GNDA.n1733 GNDA.n1717 1.90331
R17437 GNDA.n1742 GNDA.n1741 1.90331
R17438 GNDA.t111 GNDA.t202 1.7605
R17439 GNDA.t190 GNDA.t112 1.7605
R17440 GNDA.t199 GNDA.n3383 1.7605
R17441 GNDA.n3390 GNDA.t184 1.7605
R17442 GNDA.t91 GNDA.n3393 1.7605
R17443 GNDA.t229 GNDA.t93 1.7605
R17444 GNDA.t95 GNDA.t214 1.7605
R17445 GNDA.n976 GNDA.n975 1.70567
R17446 GNDA.n993 GNDA.n975 1.70567
R17447 GNDA.n996 GNDA.n975 1.70567
R17448 GNDA.n999 GNDA.n975 1.70567
R17449 GNDA.n1002 GNDA.n975 1.70567
R17450 GNDA.n1005 GNDA.n975 1.70567
R17451 GNDA.n1008 GNDA.n975 1.70567
R17452 GNDA.n1011 GNDA.n975 1.70567
R17453 GNDA.n1014 GNDA.n975 1.70567
R17454 GNDA.n1017 GNDA.n975 1.70567
R17455 GNDA.n1020 GNDA.n975 1.70567
R17456 GNDA.n1023 GNDA.n975 1.70567
R17457 GNDA.n1026 GNDA.n975 1.70567
R17458 GNDA.n1029 GNDA.n975 1.70567
R17459 GNDA.n1032 GNDA.n975 1.70567
R17460 GNDA.n975 GNDA.n916 1.70567
R17461 GNDA.n1131 GNDA.n1130 1.70567
R17462 GNDA.n1130 GNDA.n1116 1.70567
R17463 GNDA.n1130 GNDA.n1117 1.70567
R17464 GNDA.n1130 GNDA.n1118 1.70567
R17465 GNDA.n1130 GNDA.n1119 1.70567
R17466 GNDA.n1130 GNDA.n1120 1.70567
R17467 GNDA.n1130 GNDA.n1121 1.70567
R17468 GNDA.n1130 GNDA.n1122 1.70567
R17469 GNDA.n1130 GNDA.n1123 1.70567
R17470 GNDA.n1130 GNDA.n1124 1.70567
R17471 GNDA.n1130 GNDA.n1125 1.70567
R17472 GNDA.n1130 GNDA.n1126 1.70567
R17473 GNDA.n1130 GNDA.n1127 1.70567
R17474 GNDA.n1130 GNDA.n1128 1.70567
R17475 GNDA.n1130 GNDA.n1129 1.70567
R17476 GNDA.n1130 GNDA.n1074 1.70567
R17477 GNDA.n1052 GNDA.n825 1.70567
R17478 GNDA.n915 GNDA.n902 1.70567
R17479 GNDA.n915 GNDA.n903 1.70567
R17480 GNDA.n915 GNDA.n904 1.70567
R17481 GNDA.n915 GNDA.n905 1.70567
R17482 GNDA.n915 GNDA.n906 1.70567
R17483 GNDA.n915 GNDA.n907 1.70567
R17484 GNDA.n915 GNDA.n908 1.70567
R17485 GNDA.n915 GNDA.n909 1.70567
R17486 GNDA.n915 GNDA.n910 1.70567
R17487 GNDA.n915 GNDA.n911 1.70567
R17488 GNDA.n915 GNDA.n912 1.70567
R17489 GNDA.n915 GNDA.n913 1.70567
R17490 GNDA.n915 GNDA.n914 1.70567
R17491 GNDA.n915 GNDA.n884 1.70567
R17492 GNDA.n915 GNDA.n810 1.70567
R17493 GNDA.n1034 GNDA.n974 1.70565
R17494 GNDA.n974 GNDA.n972 1.70565
R17495 GNDA.n974 GNDA.n970 1.70565
R17496 GNDA.n974 GNDA.n968 1.70565
R17497 GNDA.n974 GNDA.n966 1.70565
R17498 GNDA.n974 GNDA.n964 1.70565
R17499 GNDA.n974 GNDA.n962 1.70565
R17500 GNDA.n992 GNDA.n988 1.70565
R17501 GNDA.n992 GNDA.n987 1.70565
R17502 GNDA.n992 GNDA.n984 1.70565
R17503 GNDA.n992 GNDA.n983 1.70565
R17504 GNDA.n992 GNDA.n980 1.70565
R17505 GNDA.n992 GNDA.n979 1.70565
R17506 GNDA.n1038 GNDA.n931 1.70565
R17507 GNDA.n1089 GNDA.n1059 1.70565
R17508 GNDA.n1093 GNDA.n1059 1.70565
R17509 GNDA.n1097 GNDA.n1059 1.70565
R17510 GNDA.n1101 GNDA.n1059 1.70565
R17511 GNDA.n1105 GNDA.n1059 1.70565
R17512 GNDA.n1109 GNDA.n1059 1.70565
R17513 GNDA.n1113 GNDA.n1059 1.70565
R17514 GNDA.n1163 GNDA.n794 1.70565
R17515 GNDA.n1163 GNDA.n1159 1.70565
R17516 GNDA.n1163 GNDA.n1158 1.70565
R17517 GNDA.n1163 GNDA.n1155 1.70565
R17518 GNDA.n1163 GNDA.n1154 1.70565
R17519 GNDA.n1163 GNDA.n1151 1.70565
R17520 GNDA.n1163 GNDA.n1150 1.70565
R17521 GNDA.n1053 GNDA.n1049 1.70565
R17522 GNDA.n1053 GNDA.n1048 1.70565
R17523 GNDA.n1053 GNDA.n1045 1.70565
R17524 GNDA.n1053 GNDA.n1044 1.70565
R17525 GNDA.n1053 GNDA.n1041 1.70565
R17526 GNDA.n1053 GNDA.n1040 1.70565
R17527 GNDA.n1053 GNDA.n856 1.70565
R17528 GNDA.n869 GNDA.n867 1.70565
R17529 GNDA.n869 GNDA.n865 1.70565
R17530 GNDA.n869 GNDA.n863 1.70565
R17531 GNDA.n869 GNDA.n861 1.70565
R17532 GNDA.n869 GNDA.n859 1.70565
R17533 GNDA.n869 GNDA.n857 1.70565
R17534 GNDA.n855 GNDA.n854 1.70565
R17535 GNDA.n871 GNDA.n870 1.70565
R17536 GNDA.n1058 GNDA.n839 1.70565
R17537 GNDA.n974 GNDA.n973 1.70563
R17538 GNDA.n974 GNDA.n969 1.70563
R17539 GNDA.n974 GNDA.n965 1.70563
R17540 GNDA.n974 GNDA.n961 1.70563
R17541 GNDA.n992 GNDA.n990 1.70563
R17542 GNDA.n992 GNDA.n989 1.70563
R17543 GNDA.n992 GNDA.n986 1.70563
R17544 GNDA.n992 GNDA.n985 1.70563
R17545 GNDA.n992 GNDA.n982 1.70563
R17546 GNDA.n992 GNDA.n981 1.70563
R17547 GNDA.n992 GNDA.n978 1.70563
R17548 GNDA.n992 GNDA.n977 1.70563
R17549 GNDA.n991 GNDA.n98 1.70563
R17550 GNDA.n997 GNDA.n98 1.70563
R17551 GNDA.n1003 GNDA.n98 1.70563
R17552 GNDA.n1009 GNDA.n98 1.70563
R17553 GNDA.n1015 GNDA.n98 1.70563
R17554 GNDA.n1021 GNDA.n98 1.70563
R17555 GNDA.n1027 GNDA.n98 1.70563
R17556 GNDA.n1033 GNDA.n98 1.70563
R17557 GNDA.n1091 GNDA.n1059 1.70563
R17558 GNDA.n1099 GNDA.n1059 1.70563
R17559 GNDA.n1107 GNDA.n1059 1.70563
R17560 GNDA.n1146 GNDA.n1059 1.70563
R17561 GNDA.n1163 GNDA.n1161 1.70563
R17562 GNDA.n1163 GNDA.n1160 1.70563
R17563 GNDA.n1163 GNDA.n1157 1.70563
R17564 GNDA.n1163 GNDA.n1156 1.70563
R17565 GNDA.n1163 GNDA.n1153 1.70563
R17566 GNDA.n1163 GNDA.n1152 1.70563
R17567 GNDA.n1163 GNDA.n1149 1.70563
R17568 GNDA.n1148 GNDA.n1147 1.70563
R17569 GNDA.n1147 GNDA.n1144 1.70563
R17570 GNDA.n1147 GNDA.n1142 1.70563
R17571 GNDA.n1147 GNDA.n1140 1.70563
R17572 GNDA.n1147 GNDA.n1138 1.70563
R17573 GNDA.n1147 GNDA.n1136 1.70563
R17574 GNDA.n1147 GNDA.n1134 1.70563
R17575 GNDA.n1147 GNDA.n1132 1.70563
R17576 GNDA.n1165 GNDA.n1075 1.70563
R17577 GNDA.n1053 GNDA.n1051 1.70563
R17578 GNDA.n1053 GNDA.n1050 1.70563
R17579 GNDA.n1053 GNDA.n1047 1.70563
R17580 GNDA.n1053 GNDA.n1046 1.70563
R17581 GNDA.n1053 GNDA.n1043 1.70563
R17582 GNDA.n1053 GNDA.n1042 1.70563
R17583 GNDA.n1053 GNDA.n1039 1.70563
R17584 GNDA.n1054 GNDA.n1053 1.70563
R17585 GNDA.n869 GNDA.n868 1.70563
R17586 GNDA.n869 GNDA.n864 1.70563
R17587 GNDA.n869 GNDA.n860 1.70563
R17588 GNDA.n901 GNDA.n869 1.70563
R17589 GNDA.n899 GNDA.n898 1.70563
R17590 GNDA.n899 GNDA.n896 1.70563
R17591 GNDA.n899 GNDA.n894 1.70563
R17592 GNDA.n899 GNDA.n892 1.70563
R17593 GNDA.n899 GNDA.n890 1.70563
R17594 GNDA.n899 GNDA.n888 1.70563
R17595 GNDA.n899 GNDA.n886 1.70563
R17596 GNDA.n900 GNDA.n899 1.70563
R17597 GNDA.n974 GNDA.n971 1.70556
R17598 GNDA.n974 GNDA.n967 1.70556
R17599 GNDA.n974 GNDA.n963 1.70556
R17600 GNDA.n994 GNDA.n98 1.70556
R17601 GNDA.n1000 GNDA.n98 1.70556
R17602 GNDA.n1006 GNDA.n98 1.70556
R17603 GNDA.n1012 GNDA.n98 1.70556
R17604 GNDA.n1018 GNDA.n98 1.70556
R17605 GNDA.n1024 GNDA.n98 1.70556
R17606 GNDA.n1030 GNDA.n98 1.70556
R17607 GNDA.n1095 GNDA.n1059 1.70556
R17608 GNDA.n1103 GNDA.n1059 1.70556
R17609 GNDA.n1111 GNDA.n1059 1.70556
R17610 GNDA.n1147 GNDA.n1145 1.70556
R17611 GNDA.n1147 GNDA.n1143 1.70556
R17612 GNDA.n1147 GNDA.n1141 1.70556
R17613 GNDA.n1147 GNDA.n1139 1.70556
R17614 GNDA.n1147 GNDA.n1137 1.70556
R17615 GNDA.n1147 GNDA.n1135 1.70556
R17616 GNDA.n1147 GNDA.n1133 1.70556
R17617 GNDA.n869 GNDA.n866 1.70556
R17618 GNDA.n869 GNDA.n862 1.70556
R17619 GNDA.n869 GNDA.n858 1.70556
R17620 GNDA.n899 GNDA.n897 1.70556
R17621 GNDA.n899 GNDA.n895 1.70556
R17622 GNDA.n899 GNDA.n893 1.70556
R17623 GNDA.n899 GNDA.n891 1.70556
R17624 GNDA.n899 GNDA.n889 1.70556
R17625 GNDA.n899 GNDA.n887 1.70556
R17626 GNDA.n899 GNDA.n885 1.70556
R17627 GNDA.n1514 GNDA.n1375 1.69433
R17628 GNDA.n1514 GNDA.n1372 1.69433
R17629 GNDA.n1514 GNDA.n1369 1.69433
R17630 GNDA.n1514 GNDA.n1366 1.69433
R17631 GNDA.n1514 GNDA.n1363 1.69433
R17632 GNDA.n1514 GNDA.n1360 1.69433
R17633 GNDA.n1514 GNDA.n1357 1.69433
R17634 GNDA.n1624 GNDA.n728 1.69433
R17635 GNDA.n1633 GNDA.n728 1.69433
R17636 GNDA.n1642 GNDA.n728 1.69433
R17637 GNDA.n1651 GNDA.n728 1.69433
R17638 GNDA.n1660 GNDA.n728 1.69433
R17639 GNDA.n1669 GNDA.n728 1.69433
R17640 GNDA.n1678 GNDA.n728 1.69433
R17641 GNDA.n1938 GNDA.n750 1.69433
R17642 GNDA.n1938 GNDA.n747 1.69433
R17643 GNDA.n1938 GNDA.n744 1.69433
R17644 GNDA.n1938 GNDA.n741 1.69433
R17645 GNDA.n1938 GNDA.n738 1.69433
R17646 GNDA.n1938 GNDA.n735 1.69433
R17647 GNDA.n1938 GNDA.n732 1.69433
R17648 GNDA.n2098 GNDA.n1959 1.69433
R17649 GNDA.n2098 GNDA.n1956 1.69433
R17650 GNDA.n2098 GNDA.n1953 1.69433
R17651 GNDA.n2098 GNDA.n1950 1.69433
R17652 GNDA.n2098 GNDA.n1947 1.69433
R17653 GNDA.n2098 GNDA.n1944 1.69433
R17654 GNDA.n2098 GNDA.n1941 1.69433
R17655 GNDA.n2211 GNDA.n665 1.69433
R17656 GNDA.n2220 GNDA.n665 1.69433
R17657 GNDA.n2229 GNDA.n665 1.69433
R17658 GNDA.n2238 GNDA.n665 1.69433
R17659 GNDA.n2247 GNDA.n665 1.69433
R17660 GNDA.n2256 GNDA.n665 1.69433
R17661 GNDA.n2265 GNDA.n665 1.69433
R17662 GNDA.n2561 GNDA.n2422 1.69433
R17663 GNDA.n2561 GNDA.n2419 1.69433
R17664 GNDA.n2561 GNDA.n2416 1.69433
R17665 GNDA.n2561 GNDA.n2413 1.69433
R17666 GNDA.n2561 GNDA.n2410 1.69433
R17667 GNDA.n2561 GNDA.n2407 1.69433
R17668 GNDA.n2561 GNDA.n2404 1.69433
R17669 GNDA.n2671 GNDA.n599 1.69433
R17670 GNDA.n2680 GNDA.n599 1.69433
R17671 GNDA.n2689 GNDA.n599 1.69433
R17672 GNDA.n2698 GNDA.n599 1.69433
R17673 GNDA.n2707 GNDA.n599 1.69433
R17674 GNDA.n2716 GNDA.n599 1.69433
R17675 GNDA.n2725 GNDA.n599 1.69433
R17676 GNDA.n2863 GNDA.n621 1.69433
R17677 GNDA.n2863 GNDA.n618 1.69433
R17678 GNDA.n2863 GNDA.n615 1.69433
R17679 GNDA.n2863 GNDA.n612 1.69433
R17680 GNDA.n2863 GNDA.n609 1.69433
R17681 GNDA.n2863 GNDA.n606 1.69433
R17682 GNDA.n2863 GNDA.n603 1.69433
R17683 GNDA.n2401 GNDA.n687 1.69433
R17684 GNDA.n2401 GNDA.n684 1.69433
R17685 GNDA.n2401 GNDA.n681 1.69433
R17686 GNDA.n2401 GNDA.n678 1.69433
R17687 GNDA.n2401 GNDA.n675 1.69433
R17688 GNDA.n2401 GNDA.n672 1.69433
R17689 GNDA.n2401 GNDA.n669 1.69433
R17690 GNDA.n3037 GNDA.n2885 1.69433
R17691 GNDA.n3037 GNDA.n2882 1.69433
R17692 GNDA.n3037 GNDA.n2879 1.69433
R17693 GNDA.n3037 GNDA.n2876 1.69433
R17694 GNDA.n3037 GNDA.n2873 1.69433
R17695 GNDA.n3037 GNDA.n2870 1.69433
R17696 GNDA.n3037 GNDA.n2867 1.69433
R17697 GNDA.n3197 GNDA.n3058 1.69433
R17698 GNDA.n3197 GNDA.n3055 1.69433
R17699 GNDA.n3197 GNDA.n3052 1.69433
R17700 GNDA.n3197 GNDA.n3049 1.69433
R17701 GNDA.n3197 GNDA.n3046 1.69433
R17702 GNDA.n3197 GNDA.n3043 1.69433
R17703 GNDA.n3197 GNDA.n3040 1.69433
R17704 GNDA.n3308 GNDA.n329 1.69433
R17705 GNDA.n3317 GNDA.n329 1.69433
R17706 GNDA.n3326 GNDA.n329 1.69433
R17707 GNDA.n3335 GNDA.n329 1.69433
R17708 GNDA.n3344 GNDA.n329 1.69433
R17709 GNDA.n3353 GNDA.n329 1.69433
R17710 GNDA.n3362 GNDA.n329 1.69433
R17711 GNDA.n5135 GNDA.n374 1.69433
R17712 GNDA.n5135 GNDA.n371 1.69433
R17713 GNDA.n5135 GNDA.n368 1.69433
R17714 GNDA.n5135 GNDA.n365 1.69433
R17715 GNDA.n5135 GNDA.n362 1.69433
R17716 GNDA.n5135 GNDA.n359 1.69433
R17717 GNDA.n5135 GNDA.n356 1.69433
R17718 GNDA.n505 GNDA.n377 1.69433
R17719 GNDA.n514 GNDA.n377 1.69433
R17720 GNDA.n523 GNDA.n377 1.69433
R17721 GNDA.n532 GNDA.n377 1.69433
R17722 GNDA.n541 GNDA.n377 1.69433
R17723 GNDA.n550 GNDA.n377 1.69433
R17724 GNDA.n559 GNDA.n377 1.69433
R17725 GNDA.n3611 GNDA.n3459 1.69433
R17726 GNDA.n3620 GNDA.n3459 1.69433
R17727 GNDA.n3629 GNDA.n3459 1.69433
R17728 GNDA.n3638 GNDA.n3459 1.69433
R17729 GNDA.n3647 GNDA.n3459 1.69433
R17730 GNDA.n3656 GNDA.n3459 1.69433
R17731 GNDA.n3665 GNDA.n3459 1.69433
R17732 GNDA.n3969 GNDA.n3825 1.69433
R17733 GNDA.n3969 GNDA.n3822 1.69433
R17734 GNDA.n3969 GNDA.n3819 1.69433
R17735 GNDA.n3969 GNDA.n3816 1.69433
R17736 GNDA.n3969 GNDA.n3813 1.69433
R17737 GNDA.n3969 GNDA.n3810 1.69433
R17738 GNDA.n3969 GNDA.n3807 1.69433
R17739 GNDA.n4135 GNDA.n3991 1.69433
R17740 GNDA.n4135 GNDA.n3988 1.69433
R17741 GNDA.n4135 GNDA.n3985 1.69433
R17742 GNDA.n4135 GNDA.n3982 1.69433
R17743 GNDA.n4135 GNDA.n3979 1.69433
R17744 GNDA.n4135 GNDA.n3976 1.69433
R17745 GNDA.n4135 GNDA.n3973 1.69433
R17746 GNDA.n3803 GNDA.n3481 1.69433
R17747 GNDA.n3803 GNDA.n3478 1.69433
R17748 GNDA.n3803 GNDA.n3475 1.69433
R17749 GNDA.n3803 GNDA.n3472 1.69433
R17750 GNDA.n3803 GNDA.n3469 1.69433
R17751 GNDA.n3803 GNDA.n3466 1.69433
R17752 GNDA.n3803 GNDA.n3463 1.69433
R17753 GNDA.n4301 GNDA.n4157 1.69433
R17754 GNDA.n4301 GNDA.n4154 1.69433
R17755 GNDA.n4301 GNDA.n4151 1.69433
R17756 GNDA.n4301 GNDA.n4148 1.69433
R17757 GNDA.n4301 GNDA.n4145 1.69433
R17758 GNDA.n4301 GNDA.n4142 1.69433
R17759 GNDA.n4301 GNDA.n4139 1.69433
R17760 GNDA.n4467 GNDA.n4323 1.69433
R17761 GNDA.n4467 GNDA.n4320 1.69433
R17762 GNDA.n4467 GNDA.n4317 1.69433
R17763 GNDA.n4467 GNDA.n4314 1.69433
R17764 GNDA.n4467 GNDA.n4311 1.69433
R17765 GNDA.n4467 GNDA.n4308 1.69433
R17766 GNDA.n4467 GNDA.n4305 1.69433
R17767 GNDA.n4633 GNDA.n4489 1.69433
R17768 GNDA.n4633 GNDA.n4486 1.69433
R17769 GNDA.n4633 GNDA.n4483 1.69433
R17770 GNDA.n4633 GNDA.n4480 1.69433
R17771 GNDA.n4633 GNDA.n4477 1.69433
R17772 GNDA.n4633 GNDA.n4474 1.69433
R17773 GNDA.n4633 GNDA.n4471 1.69433
R17774 GNDA.n4799 GNDA.n4655 1.69433
R17775 GNDA.n4799 GNDA.n4652 1.69433
R17776 GNDA.n4799 GNDA.n4649 1.69433
R17777 GNDA.n4799 GNDA.n4646 1.69433
R17778 GNDA.n4799 GNDA.n4643 1.69433
R17779 GNDA.n4799 GNDA.n4640 1.69433
R17780 GNDA.n4799 GNDA.n4637 1.69433
R17781 GNDA.n4959 GNDA.n4820 1.69433
R17782 GNDA.n4959 GNDA.n4817 1.69433
R17783 GNDA.n4959 GNDA.n4814 1.69433
R17784 GNDA.n4959 GNDA.n4811 1.69433
R17785 GNDA.n4959 GNDA.n4808 1.69433
R17786 GNDA.n4959 GNDA.n4805 1.69433
R17787 GNDA.n4959 GNDA.n4802 1.69433
R17788 GNDA.n5272 GNDA.n350 1.69433
R17789 GNDA.n5272 GNDA.n347 1.69433
R17790 GNDA.n5272 GNDA.n344 1.69433
R17791 GNDA.n5272 GNDA.n341 1.69433
R17792 GNDA.n5272 GNDA.n338 1.69433
R17793 GNDA.n5272 GNDA.n335 1.69433
R17794 GNDA.n5272 GNDA.n332 1.69433
R17795 GNDA.n7065 GNDA.n120 1.69433
R17796 GNDA.n7065 GNDA.n117 1.69433
R17797 GNDA.n7065 GNDA.n114 1.69433
R17798 GNDA.n7065 GNDA.n111 1.69433
R17799 GNDA.n7065 GNDA.n108 1.69433
R17800 GNDA.n7065 GNDA.n105 1.69433
R17801 GNDA.n7065 GNDA.n102 1.69433
R17802 GNDA.n7225 GNDA.n7087 1.69433
R17803 GNDA.n7225 GNDA.n7084 1.69433
R17804 GNDA.n7225 GNDA.n7081 1.69433
R17805 GNDA.n7225 GNDA.n7078 1.69433
R17806 GNDA.n7225 GNDA.n7075 1.69433
R17807 GNDA.n7225 GNDA.n7072 1.69433
R17808 GNDA.n7225 GNDA.n7069 1.69433
R17809 GNDA.n1354 GNDA.n1189 1.69337
R17810 GNDA.n1354 GNDA.n1188 1.69337
R17811 GNDA.n1354 GNDA.n1186 1.69337
R17812 GNDA.n1354 GNDA.n1185 1.69337
R17813 GNDA.n1354 GNDA.n1183 1.69337
R17814 GNDA.n1354 GNDA.n1182 1.69337
R17815 GNDA.n1354 GNDA.n1180 1.69337
R17816 GNDA.n1354 GNDA.n1179 1.69337
R17817 GNDA.n1354 GNDA.n1177 1.69337
R17818 GNDA.n1354 GNDA.n1176 1.69337
R17819 GNDA.n1354 GNDA.n1174 1.69337
R17820 GNDA.n1354 GNDA.n1173 1.69337
R17821 GNDA.n1354 GNDA.n1171 1.69337
R17822 GNDA.n1354 GNDA.n1170 1.69337
R17823 GNDA.n1354 GNDA.n1168 1.69337
R17824 GNDA.n1354 GNDA.n1167 1.69337
R17825 GNDA.n1514 GNDA.n1377 1.6924
R17826 GNDA.n1514 GNDA.n1376 1.6924
R17827 GNDA.n1514 GNDA.n1374 1.6924
R17828 GNDA.n1514 GNDA.n1373 1.6924
R17829 GNDA.n1514 GNDA.n1371 1.6924
R17830 GNDA.n1514 GNDA.n1370 1.6924
R17831 GNDA.n1514 GNDA.n1368 1.6924
R17832 GNDA.n1514 GNDA.n1367 1.6924
R17833 GNDA.n1514 GNDA.n1365 1.6924
R17834 GNDA.n1514 GNDA.n1364 1.6924
R17835 GNDA.n1514 GNDA.n1362 1.6924
R17836 GNDA.n1514 GNDA.n1361 1.6924
R17837 GNDA.n1514 GNDA.n1359 1.6924
R17838 GNDA.n1514 GNDA.n1358 1.6924
R17839 GNDA.n1514 GNDA.n1356 1.6924
R17840 GNDA.n1514 GNDA.n1355 1.6924
R17841 GNDA.n1618 GNDA.n728 1.6924
R17842 GNDA.n1621 GNDA.n728 1.6924
R17843 GNDA.n1627 GNDA.n728 1.6924
R17844 GNDA.n1630 GNDA.n728 1.6924
R17845 GNDA.n1636 GNDA.n728 1.6924
R17846 GNDA.n1639 GNDA.n728 1.6924
R17847 GNDA.n1645 GNDA.n728 1.6924
R17848 GNDA.n1648 GNDA.n728 1.6924
R17849 GNDA.n1654 GNDA.n728 1.6924
R17850 GNDA.n1657 GNDA.n728 1.6924
R17851 GNDA.n1663 GNDA.n728 1.6924
R17852 GNDA.n1666 GNDA.n728 1.6924
R17853 GNDA.n1672 GNDA.n728 1.6924
R17854 GNDA.n1675 GNDA.n728 1.6924
R17855 GNDA.n1681 GNDA.n728 1.6924
R17856 GNDA.n1684 GNDA.n728 1.6924
R17857 GNDA.n1938 GNDA.n752 1.6924
R17858 GNDA.n1938 GNDA.n751 1.6924
R17859 GNDA.n1938 GNDA.n749 1.6924
R17860 GNDA.n1938 GNDA.n748 1.6924
R17861 GNDA.n1938 GNDA.n746 1.6924
R17862 GNDA.n1938 GNDA.n745 1.6924
R17863 GNDA.n1938 GNDA.n743 1.6924
R17864 GNDA.n1938 GNDA.n742 1.6924
R17865 GNDA.n1938 GNDA.n740 1.6924
R17866 GNDA.n1938 GNDA.n739 1.6924
R17867 GNDA.n1938 GNDA.n737 1.6924
R17868 GNDA.n1938 GNDA.n736 1.6924
R17869 GNDA.n1938 GNDA.n734 1.6924
R17870 GNDA.n1938 GNDA.n733 1.6924
R17871 GNDA.n1938 GNDA.n731 1.6924
R17872 GNDA.n1938 GNDA.n730 1.6924
R17873 GNDA.n2098 GNDA.n1961 1.6924
R17874 GNDA.n2098 GNDA.n1960 1.6924
R17875 GNDA.n2098 GNDA.n1958 1.6924
R17876 GNDA.n2098 GNDA.n1957 1.6924
R17877 GNDA.n2098 GNDA.n1955 1.6924
R17878 GNDA.n2098 GNDA.n1954 1.6924
R17879 GNDA.n2098 GNDA.n1952 1.6924
R17880 GNDA.n2098 GNDA.n1951 1.6924
R17881 GNDA.n2098 GNDA.n1949 1.6924
R17882 GNDA.n2098 GNDA.n1948 1.6924
R17883 GNDA.n2098 GNDA.n1946 1.6924
R17884 GNDA.n2098 GNDA.n1945 1.6924
R17885 GNDA.n2098 GNDA.n1943 1.6924
R17886 GNDA.n2098 GNDA.n1942 1.6924
R17887 GNDA.n2098 GNDA.n1940 1.6924
R17888 GNDA.n2098 GNDA.n1939 1.6924
R17889 GNDA.n2205 GNDA.n665 1.6924
R17890 GNDA.n2208 GNDA.n665 1.6924
R17891 GNDA.n2214 GNDA.n665 1.6924
R17892 GNDA.n2217 GNDA.n665 1.6924
R17893 GNDA.n2223 GNDA.n665 1.6924
R17894 GNDA.n2226 GNDA.n665 1.6924
R17895 GNDA.n2232 GNDA.n665 1.6924
R17896 GNDA.n2235 GNDA.n665 1.6924
R17897 GNDA.n2241 GNDA.n665 1.6924
R17898 GNDA.n2244 GNDA.n665 1.6924
R17899 GNDA.n2250 GNDA.n665 1.6924
R17900 GNDA.n2253 GNDA.n665 1.6924
R17901 GNDA.n2259 GNDA.n665 1.6924
R17902 GNDA.n2262 GNDA.n665 1.6924
R17903 GNDA.n2268 GNDA.n665 1.6924
R17904 GNDA.n2271 GNDA.n665 1.6924
R17905 GNDA.n2561 GNDA.n2424 1.6924
R17906 GNDA.n2561 GNDA.n2423 1.6924
R17907 GNDA.n2561 GNDA.n2421 1.6924
R17908 GNDA.n2561 GNDA.n2420 1.6924
R17909 GNDA.n2561 GNDA.n2418 1.6924
R17910 GNDA.n2561 GNDA.n2417 1.6924
R17911 GNDA.n2561 GNDA.n2415 1.6924
R17912 GNDA.n2561 GNDA.n2414 1.6924
R17913 GNDA.n2561 GNDA.n2412 1.6924
R17914 GNDA.n2561 GNDA.n2411 1.6924
R17915 GNDA.n2561 GNDA.n2409 1.6924
R17916 GNDA.n2561 GNDA.n2408 1.6924
R17917 GNDA.n2561 GNDA.n2406 1.6924
R17918 GNDA.n2561 GNDA.n2405 1.6924
R17919 GNDA.n2561 GNDA.n2403 1.6924
R17920 GNDA.n2561 GNDA.n2402 1.6924
R17921 GNDA.n2665 GNDA.n599 1.6924
R17922 GNDA.n2668 GNDA.n599 1.6924
R17923 GNDA.n2674 GNDA.n599 1.6924
R17924 GNDA.n2677 GNDA.n599 1.6924
R17925 GNDA.n2683 GNDA.n599 1.6924
R17926 GNDA.n2686 GNDA.n599 1.6924
R17927 GNDA.n2692 GNDA.n599 1.6924
R17928 GNDA.n2695 GNDA.n599 1.6924
R17929 GNDA.n2701 GNDA.n599 1.6924
R17930 GNDA.n2704 GNDA.n599 1.6924
R17931 GNDA.n2710 GNDA.n599 1.6924
R17932 GNDA.n2713 GNDA.n599 1.6924
R17933 GNDA.n2719 GNDA.n599 1.6924
R17934 GNDA.n2722 GNDA.n599 1.6924
R17935 GNDA.n2728 GNDA.n599 1.6924
R17936 GNDA.n2731 GNDA.n599 1.6924
R17937 GNDA.n2863 GNDA.n623 1.6924
R17938 GNDA.n2863 GNDA.n622 1.6924
R17939 GNDA.n2863 GNDA.n620 1.6924
R17940 GNDA.n2863 GNDA.n619 1.6924
R17941 GNDA.n2863 GNDA.n617 1.6924
R17942 GNDA.n2863 GNDA.n616 1.6924
R17943 GNDA.n2863 GNDA.n614 1.6924
R17944 GNDA.n2863 GNDA.n613 1.6924
R17945 GNDA.n2863 GNDA.n611 1.6924
R17946 GNDA.n2863 GNDA.n610 1.6924
R17947 GNDA.n2863 GNDA.n608 1.6924
R17948 GNDA.n2863 GNDA.n607 1.6924
R17949 GNDA.n2863 GNDA.n605 1.6924
R17950 GNDA.n2863 GNDA.n604 1.6924
R17951 GNDA.n2863 GNDA.n602 1.6924
R17952 GNDA.n2863 GNDA.n601 1.6924
R17953 GNDA.n2401 GNDA.n689 1.6924
R17954 GNDA.n2401 GNDA.n688 1.6924
R17955 GNDA.n2401 GNDA.n686 1.6924
R17956 GNDA.n2401 GNDA.n685 1.6924
R17957 GNDA.n2401 GNDA.n683 1.6924
R17958 GNDA.n2401 GNDA.n682 1.6924
R17959 GNDA.n2401 GNDA.n680 1.6924
R17960 GNDA.n2401 GNDA.n679 1.6924
R17961 GNDA.n2401 GNDA.n677 1.6924
R17962 GNDA.n2401 GNDA.n676 1.6924
R17963 GNDA.n2401 GNDA.n674 1.6924
R17964 GNDA.n2401 GNDA.n673 1.6924
R17965 GNDA.n2401 GNDA.n671 1.6924
R17966 GNDA.n2401 GNDA.n670 1.6924
R17967 GNDA.n2401 GNDA.n668 1.6924
R17968 GNDA.n2401 GNDA.n667 1.6924
R17969 GNDA.n3037 GNDA.n2887 1.6924
R17970 GNDA.n3037 GNDA.n2886 1.6924
R17971 GNDA.n3037 GNDA.n2884 1.6924
R17972 GNDA.n3037 GNDA.n2883 1.6924
R17973 GNDA.n3037 GNDA.n2881 1.6924
R17974 GNDA.n3037 GNDA.n2880 1.6924
R17975 GNDA.n3037 GNDA.n2878 1.6924
R17976 GNDA.n3037 GNDA.n2877 1.6924
R17977 GNDA.n3037 GNDA.n2875 1.6924
R17978 GNDA.n3037 GNDA.n2874 1.6924
R17979 GNDA.n3037 GNDA.n2872 1.6924
R17980 GNDA.n3037 GNDA.n2871 1.6924
R17981 GNDA.n3037 GNDA.n2869 1.6924
R17982 GNDA.n3037 GNDA.n2868 1.6924
R17983 GNDA.n3037 GNDA.n2866 1.6924
R17984 GNDA.n3037 GNDA.n2865 1.6924
R17985 GNDA.n3197 GNDA.n3060 1.6924
R17986 GNDA.n3197 GNDA.n3059 1.6924
R17987 GNDA.n3197 GNDA.n3057 1.6924
R17988 GNDA.n3197 GNDA.n3056 1.6924
R17989 GNDA.n3197 GNDA.n3054 1.6924
R17990 GNDA.n3197 GNDA.n3053 1.6924
R17991 GNDA.n3197 GNDA.n3051 1.6924
R17992 GNDA.n3197 GNDA.n3050 1.6924
R17993 GNDA.n3197 GNDA.n3048 1.6924
R17994 GNDA.n3197 GNDA.n3047 1.6924
R17995 GNDA.n3197 GNDA.n3045 1.6924
R17996 GNDA.n3197 GNDA.n3044 1.6924
R17997 GNDA.n3197 GNDA.n3042 1.6924
R17998 GNDA.n3197 GNDA.n3041 1.6924
R17999 GNDA.n3197 GNDA.n3039 1.6924
R18000 GNDA.n3197 GNDA.n3038 1.6924
R18001 GNDA.n3302 GNDA.n329 1.6924
R18002 GNDA.n3305 GNDA.n329 1.6924
R18003 GNDA.n3311 GNDA.n329 1.6924
R18004 GNDA.n3314 GNDA.n329 1.6924
R18005 GNDA.n3320 GNDA.n329 1.6924
R18006 GNDA.n3323 GNDA.n329 1.6924
R18007 GNDA.n3329 GNDA.n329 1.6924
R18008 GNDA.n3332 GNDA.n329 1.6924
R18009 GNDA.n3338 GNDA.n329 1.6924
R18010 GNDA.n3341 GNDA.n329 1.6924
R18011 GNDA.n3347 GNDA.n329 1.6924
R18012 GNDA.n3350 GNDA.n329 1.6924
R18013 GNDA.n3356 GNDA.n329 1.6924
R18014 GNDA.n3359 GNDA.n329 1.6924
R18015 GNDA.n3365 GNDA.n329 1.6924
R18016 GNDA.n3368 GNDA.n329 1.6924
R18017 GNDA.n5135 GNDA.n376 1.6924
R18018 GNDA.n5135 GNDA.n375 1.6924
R18019 GNDA.n5135 GNDA.n373 1.6924
R18020 GNDA.n5135 GNDA.n372 1.6924
R18021 GNDA.n5135 GNDA.n370 1.6924
R18022 GNDA.n5135 GNDA.n369 1.6924
R18023 GNDA.n5135 GNDA.n367 1.6924
R18024 GNDA.n5135 GNDA.n366 1.6924
R18025 GNDA.n5135 GNDA.n364 1.6924
R18026 GNDA.n5135 GNDA.n363 1.6924
R18027 GNDA.n5135 GNDA.n361 1.6924
R18028 GNDA.n5135 GNDA.n360 1.6924
R18029 GNDA.n5135 GNDA.n358 1.6924
R18030 GNDA.n5135 GNDA.n357 1.6924
R18031 GNDA.n5135 GNDA.n355 1.6924
R18032 GNDA.n5135 GNDA.n354 1.6924
R18033 GNDA.n499 GNDA.n377 1.6924
R18034 GNDA.n502 GNDA.n377 1.6924
R18035 GNDA.n508 GNDA.n377 1.6924
R18036 GNDA.n511 GNDA.n377 1.6924
R18037 GNDA.n517 GNDA.n377 1.6924
R18038 GNDA.n520 GNDA.n377 1.6924
R18039 GNDA.n526 GNDA.n377 1.6924
R18040 GNDA.n529 GNDA.n377 1.6924
R18041 GNDA.n535 GNDA.n377 1.6924
R18042 GNDA.n538 GNDA.n377 1.6924
R18043 GNDA.n544 GNDA.n377 1.6924
R18044 GNDA.n547 GNDA.n377 1.6924
R18045 GNDA.n553 GNDA.n377 1.6924
R18046 GNDA.n556 GNDA.n377 1.6924
R18047 GNDA.n562 GNDA.n377 1.6924
R18048 GNDA.n565 GNDA.n377 1.6924
R18049 GNDA.n3605 GNDA.n3459 1.6924
R18050 GNDA.n3608 GNDA.n3459 1.6924
R18051 GNDA.n3614 GNDA.n3459 1.6924
R18052 GNDA.n3617 GNDA.n3459 1.6924
R18053 GNDA.n3623 GNDA.n3459 1.6924
R18054 GNDA.n3626 GNDA.n3459 1.6924
R18055 GNDA.n3632 GNDA.n3459 1.6924
R18056 GNDA.n3635 GNDA.n3459 1.6924
R18057 GNDA.n3641 GNDA.n3459 1.6924
R18058 GNDA.n3644 GNDA.n3459 1.6924
R18059 GNDA.n3650 GNDA.n3459 1.6924
R18060 GNDA.n3653 GNDA.n3459 1.6924
R18061 GNDA.n3659 GNDA.n3459 1.6924
R18062 GNDA.n3662 GNDA.n3459 1.6924
R18063 GNDA.n3668 GNDA.n3459 1.6924
R18064 GNDA.n3671 GNDA.n3459 1.6924
R18065 GNDA.n3969 GNDA.n3827 1.6924
R18066 GNDA.n3969 GNDA.n3826 1.6924
R18067 GNDA.n3969 GNDA.n3824 1.6924
R18068 GNDA.n3969 GNDA.n3823 1.6924
R18069 GNDA.n3969 GNDA.n3821 1.6924
R18070 GNDA.n3969 GNDA.n3820 1.6924
R18071 GNDA.n3969 GNDA.n3818 1.6924
R18072 GNDA.n3969 GNDA.n3817 1.6924
R18073 GNDA.n3969 GNDA.n3815 1.6924
R18074 GNDA.n3969 GNDA.n3814 1.6924
R18075 GNDA.n3969 GNDA.n3812 1.6924
R18076 GNDA.n3969 GNDA.n3811 1.6924
R18077 GNDA.n3969 GNDA.n3809 1.6924
R18078 GNDA.n3969 GNDA.n3808 1.6924
R18079 GNDA.n3969 GNDA.n3806 1.6924
R18080 GNDA.n3969 GNDA.n3805 1.6924
R18081 GNDA.n4135 GNDA.n3993 1.6924
R18082 GNDA.n4135 GNDA.n3992 1.6924
R18083 GNDA.n4135 GNDA.n3990 1.6924
R18084 GNDA.n4135 GNDA.n3989 1.6924
R18085 GNDA.n4135 GNDA.n3987 1.6924
R18086 GNDA.n4135 GNDA.n3986 1.6924
R18087 GNDA.n4135 GNDA.n3984 1.6924
R18088 GNDA.n4135 GNDA.n3983 1.6924
R18089 GNDA.n4135 GNDA.n3981 1.6924
R18090 GNDA.n4135 GNDA.n3980 1.6924
R18091 GNDA.n4135 GNDA.n3978 1.6924
R18092 GNDA.n4135 GNDA.n3977 1.6924
R18093 GNDA.n4135 GNDA.n3975 1.6924
R18094 GNDA.n4135 GNDA.n3974 1.6924
R18095 GNDA.n4135 GNDA.n3972 1.6924
R18096 GNDA.n4135 GNDA.n3971 1.6924
R18097 GNDA.n3803 GNDA.n3483 1.6924
R18098 GNDA.n3803 GNDA.n3482 1.6924
R18099 GNDA.n3803 GNDA.n3480 1.6924
R18100 GNDA.n3803 GNDA.n3479 1.6924
R18101 GNDA.n3803 GNDA.n3477 1.6924
R18102 GNDA.n3803 GNDA.n3476 1.6924
R18103 GNDA.n3803 GNDA.n3474 1.6924
R18104 GNDA.n3803 GNDA.n3473 1.6924
R18105 GNDA.n3803 GNDA.n3471 1.6924
R18106 GNDA.n3803 GNDA.n3470 1.6924
R18107 GNDA.n3803 GNDA.n3468 1.6924
R18108 GNDA.n3803 GNDA.n3467 1.6924
R18109 GNDA.n3803 GNDA.n3465 1.6924
R18110 GNDA.n3803 GNDA.n3464 1.6924
R18111 GNDA.n3803 GNDA.n3462 1.6924
R18112 GNDA.n3803 GNDA.n3461 1.6924
R18113 GNDA.n4301 GNDA.n4159 1.6924
R18114 GNDA.n4301 GNDA.n4158 1.6924
R18115 GNDA.n4301 GNDA.n4156 1.6924
R18116 GNDA.n4301 GNDA.n4155 1.6924
R18117 GNDA.n4301 GNDA.n4153 1.6924
R18118 GNDA.n4301 GNDA.n4152 1.6924
R18119 GNDA.n4301 GNDA.n4150 1.6924
R18120 GNDA.n4301 GNDA.n4149 1.6924
R18121 GNDA.n4301 GNDA.n4147 1.6924
R18122 GNDA.n4301 GNDA.n4146 1.6924
R18123 GNDA.n4301 GNDA.n4144 1.6924
R18124 GNDA.n4301 GNDA.n4143 1.6924
R18125 GNDA.n4301 GNDA.n4141 1.6924
R18126 GNDA.n4301 GNDA.n4140 1.6924
R18127 GNDA.n4301 GNDA.n4138 1.6924
R18128 GNDA.n4301 GNDA.n4137 1.6924
R18129 GNDA.n4467 GNDA.n4325 1.6924
R18130 GNDA.n4467 GNDA.n4324 1.6924
R18131 GNDA.n4467 GNDA.n4322 1.6924
R18132 GNDA.n4467 GNDA.n4321 1.6924
R18133 GNDA.n4467 GNDA.n4319 1.6924
R18134 GNDA.n4467 GNDA.n4318 1.6924
R18135 GNDA.n4467 GNDA.n4316 1.6924
R18136 GNDA.n4467 GNDA.n4315 1.6924
R18137 GNDA.n4467 GNDA.n4313 1.6924
R18138 GNDA.n4467 GNDA.n4312 1.6924
R18139 GNDA.n4467 GNDA.n4310 1.6924
R18140 GNDA.n4467 GNDA.n4309 1.6924
R18141 GNDA.n4467 GNDA.n4307 1.6924
R18142 GNDA.n4467 GNDA.n4306 1.6924
R18143 GNDA.n4467 GNDA.n4304 1.6924
R18144 GNDA.n4467 GNDA.n4303 1.6924
R18145 GNDA.n4633 GNDA.n4491 1.6924
R18146 GNDA.n4633 GNDA.n4490 1.6924
R18147 GNDA.n4633 GNDA.n4488 1.6924
R18148 GNDA.n4633 GNDA.n4487 1.6924
R18149 GNDA.n4633 GNDA.n4485 1.6924
R18150 GNDA.n4633 GNDA.n4484 1.6924
R18151 GNDA.n4633 GNDA.n4482 1.6924
R18152 GNDA.n4633 GNDA.n4481 1.6924
R18153 GNDA.n4633 GNDA.n4479 1.6924
R18154 GNDA.n4633 GNDA.n4478 1.6924
R18155 GNDA.n4633 GNDA.n4476 1.6924
R18156 GNDA.n4633 GNDA.n4475 1.6924
R18157 GNDA.n4633 GNDA.n4473 1.6924
R18158 GNDA.n4633 GNDA.n4472 1.6924
R18159 GNDA.n4633 GNDA.n4470 1.6924
R18160 GNDA.n4633 GNDA.n4469 1.6924
R18161 GNDA.n4799 GNDA.n4657 1.6924
R18162 GNDA.n4799 GNDA.n4656 1.6924
R18163 GNDA.n4799 GNDA.n4654 1.6924
R18164 GNDA.n4799 GNDA.n4653 1.6924
R18165 GNDA.n4799 GNDA.n4651 1.6924
R18166 GNDA.n4799 GNDA.n4650 1.6924
R18167 GNDA.n4799 GNDA.n4648 1.6924
R18168 GNDA.n4799 GNDA.n4647 1.6924
R18169 GNDA.n4799 GNDA.n4645 1.6924
R18170 GNDA.n4799 GNDA.n4644 1.6924
R18171 GNDA.n4799 GNDA.n4642 1.6924
R18172 GNDA.n4799 GNDA.n4641 1.6924
R18173 GNDA.n4799 GNDA.n4639 1.6924
R18174 GNDA.n4799 GNDA.n4638 1.6924
R18175 GNDA.n4799 GNDA.n4636 1.6924
R18176 GNDA.n4799 GNDA.n4635 1.6924
R18177 GNDA.n4959 GNDA.n4822 1.6924
R18178 GNDA.n4959 GNDA.n4821 1.6924
R18179 GNDA.n4959 GNDA.n4819 1.6924
R18180 GNDA.n4959 GNDA.n4818 1.6924
R18181 GNDA.n4959 GNDA.n4816 1.6924
R18182 GNDA.n4959 GNDA.n4815 1.6924
R18183 GNDA.n4959 GNDA.n4813 1.6924
R18184 GNDA.n4959 GNDA.n4812 1.6924
R18185 GNDA.n4959 GNDA.n4810 1.6924
R18186 GNDA.n4959 GNDA.n4809 1.6924
R18187 GNDA.n4959 GNDA.n4807 1.6924
R18188 GNDA.n4959 GNDA.n4806 1.6924
R18189 GNDA.n4959 GNDA.n4804 1.6924
R18190 GNDA.n4959 GNDA.n4803 1.6924
R18191 GNDA.n4959 GNDA.n4801 1.6924
R18192 GNDA.n4959 GNDA.n4800 1.6924
R18193 GNDA.n5272 GNDA.n352 1.6924
R18194 GNDA.n5272 GNDA.n351 1.6924
R18195 GNDA.n5272 GNDA.n349 1.6924
R18196 GNDA.n5272 GNDA.n348 1.6924
R18197 GNDA.n5272 GNDA.n346 1.6924
R18198 GNDA.n5272 GNDA.n345 1.6924
R18199 GNDA.n5272 GNDA.n343 1.6924
R18200 GNDA.n5272 GNDA.n342 1.6924
R18201 GNDA.n5272 GNDA.n340 1.6924
R18202 GNDA.n5272 GNDA.n339 1.6924
R18203 GNDA.n5272 GNDA.n337 1.6924
R18204 GNDA.n5272 GNDA.n336 1.6924
R18205 GNDA.n5272 GNDA.n334 1.6924
R18206 GNDA.n5272 GNDA.n333 1.6924
R18207 GNDA.n5272 GNDA.n331 1.6924
R18208 GNDA.n5272 GNDA.n330 1.6924
R18209 GNDA.n7065 GNDA.n122 1.6924
R18210 GNDA.n7065 GNDA.n121 1.6924
R18211 GNDA.n7065 GNDA.n119 1.6924
R18212 GNDA.n7065 GNDA.n118 1.6924
R18213 GNDA.n7065 GNDA.n116 1.6924
R18214 GNDA.n7065 GNDA.n115 1.6924
R18215 GNDA.n7065 GNDA.n113 1.6924
R18216 GNDA.n7065 GNDA.n112 1.6924
R18217 GNDA.n7065 GNDA.n110 1.6924
R18218 GNDA.n7065 GNDA.n109 1.6924
R18219 GNDA.n7065 GNDA.n107 1.6924
R18220 GNDA.n7065 GNDA.n106 1.6924
R18221 GNDA.n7065 GNDA.n104 1.6924
R18222 GNDA.n7065 GNDA.n103 1.6924
R18223 GNDA.n7065 GNDA.n101 1.6924
R18224 GNDA.n7065 GNDA.n100 1.6924
R18225 GNDA.n7225 GNDA.n7224 1.6924
R18226 GNDA.n7225 GNDA.n7088 1.6924
R18227 GNDA.n7225 GNDA.n7086 1.6924
R18228 GNDA.n7225 GNDA.n7085 1.6924
R18229 GNDA.n7225 GNDA.n7083 1.6924
R18230 GNDA.n7225 GNDA.n7082 1.6924
R18231 GNDA.n7225 GNDA.n7080 1.6924
R18232 GNDA.n7225 GNDA.n7079 1.6924
R18233 GNDA.n7225 GNDA.n7077 1.6924
R18234 GNDA.n7225 GNDA.n7076 1.6924
R18235 GNDA.n7225 GNDA.n7074 1.6924
R18236 GNDA.n7225 GNDA.n7073 1.6924
R18237 GNDA.n7225 GNDA.n7071 1.6924
R18238 GNDA.n7225 GNDA.n7070 1.6924
R18239 GNDA.n7225 GNDA.n7068 1.6924
R18240 GNDA.n7225 GNDA.n7067 1.6924
R18241 GNDA.n1354 GNDA.n1353 1.6924
R18242 GNDA.n1354 GNDA.n1187 1.6924
R18243 GNDA.n1354 GNDA.n1184 1.6924
R18244 GNDA.n1354 GNDA.n1181 1.6924
R18245 GNDA.n1354 GNDA.n1178 1.6924
R18246 GNDA.n1354 GNDA.n1175 1.6924
R18247 GNDA.n1354 GNDA.n1172 1.6924
R18248 GNDA.n1354 GNDA.n1169 1.6924
R18249 GNDA.n6777 GNDA.n6662 1.63592
R18250 GNDA.t46 GNDA.t145 1.57352
R18251 GNDA.n1775 GNDA.n1706 1.56997
R18252 GNDA.n1772 GNDA.n1707 1.56997
R18253 GNDA.n3431 GNDA.n3430 1.5005
R18254 GNDA.n1811 GNDA.n1810 1.5005
R18255 GNDA.n2281 GNDA.n715 1.5005
R18256 GNDA.n3679 GNDA.n3678 1.5005
R18257 GNDA.n6551 GNDA.n6548 1.47392
R18258 GNDA.n6574 GNDA.n5405 1.47392
R18259 GNDA.n5762 GNDA.n5639 1.47392
R18260 GNDA.n5882 GNDA.n5880 1.47392
R18261 GNDA.n7006 GNDA.n7005 1.47392
R18262 GNDA.n7392 GNDA.n7315 1.47392
R18263 GNDA.n5409 GNDA.t279 1.31483
R18264 GNDA.n3427 GNDA.n3425 1.07342
R18265 GNDA.n1805 GNDA.n1804 1.07342
R18266 GNDA.t126 GNDA.t34 1.06911
R18267 GNDA.n1776 GNDA.n1775 1.063
R18268 GNDA.n1772 GNDA.n1771 1.063
R18269 GNDA.t70 GNDA.t332 1.02079
R18270 GNDA.n7052 GNDA.n7051 1.01092
R18271 GNDA.n7234 GNDA.n7233 0.839515
R18272 GNDA.n6445 GNDA.n6345 0.8197
R18273 GNDA.n6444 GNDA.n6346 0.8197
R18274 GNDA.n6358 GNDA.n6355 0.8197
R18275 GNDA.n6361 GNDA.n6360 0.8197
R18276 GNDA.n6369 GNDA.n6368 0.8197
R18277 GNDA.n6372 GNDA.n6354 0.8197
R18278 GNDA.n6374 GNDA.n6373 0.8197
R18279 GNDA.n7479 GNDA.n56 0.8197
R18280 GNDA.n6540 GNDA.n6324 0.8197
R18281 GNDA.n6539 GNDA.n6325 0.8197
R18282 GNDA.n6459 GNDA.n6456 0.8197
R18283 GNDA.n6462 GNDA.n6461 0.8197
R18284 GNDA.n6472 GNDA.n6469 0.8197
R18285 GNDA.n6473 GNDA.n6455 0.8197
R18286 GNDA.n6477 GNDA.n6476 0.8197
R18287 GNDA.n6481 GNDA.n6480 0.8197
R18288 GNDA.n6974 GNDA.n6973 0.8197
R18289 GNDA.n6960 GNDA.n5345 0.8197
R18290 GNDA.n6967 GNDA.n6961 0.8197
R18291 GNDA.n6966 GNDA.n6963 0.8197
R18292 GNDA.n6979 GNDA.n5323 0.8197
R18293 GNDA.n6839 GNDA.n6838 0.8197
R18294 GNDA.n6846 GNDA.n6837 0.8197
R18295 GNDA.n6848 GNDA.n6847 0.8197
R18296 GNDA.n6819 GNDA.n6576 0.8197
R18297 GNDA.n6816 GNDA.n6815 0.8197
R18298 GNDA.n6797 GNDA.n6641 0.8197
R18299 GNDA.n6809 GNDA.n6798 0.8197
R18300 GNDA.n6802 GNDA.n6801 0.8197
R18301 GNDA.n6828 GNDA.n5399 0.8197
R18302 GNDA.n6830 GNDA.n6829 0.8197
R18303 GNDA.n6908 GNDA.n5395 0.8197
R18304 GNDA.n5743 GNDA.n5742 0.8197
R18305 GNDA.n5739 GNDA.n5738 0.8197
R18306 GNDA.n5735 GNDA.n5719 0.8197
R18307 GNDA.n5734 GNDA.n5731 0.8197
R18308 GNDA.n5727 GNDA.n5724 0.8197
R18309 GNDA.n5721 GNDA.n5643 0.8197
R18310 GNDA.n5749 GNDA.n5748 0.8197
R18311 GNDA.n5752 GNDA.n5642 0.8197
R18312 GNDA.n6062 GNDA.n5452 0.8197
R18313 GNDA.n6061 GNDA.n5454 0.8197
R18314 GNDA.n5506 GNDA.n5488 0.8197
R18315 GNDA.n5505 GNDA.n5503 0.8197
R18316 GNDA.n5499 GNDA.n5498 0.8197
R18317 GNDA.n5495 GNDA.n5491 0.8197
R18318 GNDA.n5494 GNDA.n5474 0.8197
R18319 GNDA.n6003 GNDA.n6002 0.8197
R18320 GNDA.n5993 GNDA.n5885 0.8197
R18321 GNDA.n5990 GNDA.n5989 0.8197
R18322 GNDA.n5986 GNDA.n5888 0.8197
R18323 GNDA.n5985 GNDA.n5889 0.8197
R18324 GNDA.n5920 GNDA.n5917 0.8197
R18325 GNDA.n5921 GNDA.n5911 0.8197
R18326 GNDA.n5925 GNDA.n5924 0.8197
R18327 GNDA.n5929 GNDA.n5928 0.8197
R18328 GNDA.n6740 GNDA.n6670 0.8197
R18329 GNDA.n6751 GNDA.n6750 0.8197
R18330 GNDA.n6668 GNDA.n6667 0.8197
R18331 GNDA.n6760 GNDA.n6757 0.8197
R18332 GNDA.n7021 GNDA.n7020 0.8197
R18333 GNDA.n294 GNDA.n293 0.8197
R18334 GNDA.n7029 GNDA.n290 0.8197
R18335 GNDA.n7028 GNDA.n291 0.8197
R18336 GNDA.n7486 GNDA.n7485 0.8197
R18337 GNDA.n32 GNDA.n23 0.8197
R18338 GNDA.n39 GNDA.n33 0.8197
R18339 GNDA.n38 GNDA.n35 0.8197
R18340 GNDA.n7491 GNDA.n1 0.8197
R18341 GNDA.n7376 GNDA.n7373 0.8197
R18342 GNDA.n7379 GNDA.n7378 0.8197
R18343 GNDA.n7382 GNDA.n7372 0.8197
R18344 GNDA.n3419 GNDA.n3418 0.786958
R18345 GNDA.n1799 GNDA.n1798 0.786958
R18346 GNDA.n5314 GNDA.n318 0.78175
R18347 GNDA.n3401 GNDA.n3398 0.78175
R18348 GNDA.n5277 GNDA.n5275 0.776542
R18349 GNDA.n4963 GNDA.n4962 0.776542
R18350 GNDA.n4682 GNDA.n3451 0.776542
R18351 GNDA.n4516 GNDA.n3446 0.776542
R18352 GNDA.n4350 GNDA.n3441 0.776542
R18353 GNDA.n4184 GNDA.n3436 0.776542
R18354 GNDA.n4018 GNDA.n584 0.776542
R18355 GNDA.n3852 GNDA.n579 0.776542
R18356 GNDA.n570 GNDA.n569 0.776542
R18357 GNDA.n5018 GNDA.n5017 0.776542
R18358 GNDA.n3373 GNDA.n3372 0.776542
R18359 GNDA.n3201 GNDA.n3200 0.776542
R18360 GNDA.n2920 GNDA.n2919 0.776542
R18361 GNDA.n2746 GNDA.n2745 0.776542
R18362 GNDA.n2736 GNDA.n2735 0.776542
R18363 GNDA.n2565 GNDA.n2564 0.776542
R18364 GNDA.n1821 GNDA.n1820 0.776542
R18365 GNDA.n1689 GNDA.n1688 0.776542
R18366 GNDA.n1518 GNDA.n1517 0.776542
R18367 GNDA.n1239 GNDA.n1238 0.776542
R18368 GNDA.n2102 GNDA.n2101 0.776542
R18369 GNDA.n3686 GNDA.n3685 0.77295
R18370 GNDA.n2276 GNDA.n2275 0.77295
R18371 GNDA.n3676 GNDA.n3675 0.755708
R18372 GNDA.n2284 GNDA.n2283 0.755708
R18373 GNDA.n3676 GNDA.n573 0.751
R18374 GNDA.n2283 GNDA.n2282 0.751
R18375 GNDA.n5315 GNDA.n317 0.729667
R18376 GNDA.n1726 GNDA.n318 0.729667
R18377 GNDA.n3398 GNDA.n590 0.729667
R18378 GNDA.n3429 GNDA.n3404 0.729667
R18379 GNDA.n6946 GNDA.n5355 0.71925
R18380 GNDA.n5315 GNDA.n5314 0.688
R18381 GNDA.n3404 GNDA.n3401 0.688
R18382 GNDA.n1743 GNDA.n1742 0.688
R18383 GNDA.n1756 GNDA.n1717 0.688
R18384 GNDA.n7059 GNDA.n7058 0.677583
R18385 GNDA.n6778 GNDA.n6777 0.65675
R18386 GNDA.n6365 GNDA 0.5637
R18387 GNDA.n6466 GNDA 0.5637
R18388 GNDA.n6962 GNDA 0.5637
R18389 GNDA.n6808 GNDA 0.5637
R18390 GNDA GNDA.n5720 0.5637
R18391 GNDA.n5502 GNDA 0.5637
R18392 GNDA GNDA.n5912 0.5637
R18393 GNDA.n6759 GNDA 0.5637
R18394 GNDA.n34 GNDA 0.5637
R18395 GNDA.n5304 GNDA.n5302 0.563
R18396 GNDA.n5302 GNDA.n5300 0.563
R18397 GNDA.n5300 GNDA.n5298 0.563
R18398 GNDA.n5298 GNDA.n5296 0.563
R18399 GNDA.n5296 GNDA.n5294 0.563
R18400 GNDA.n5294 GNDA.n5292 0.563
R18401 GNDA.n5292 GNDA.n5290 0.563
R18402 GNDA.n5290 GNDA.n5288 0.563
R18403 GNDA.n5288 GNDA.n5286 0.563
R18404 GNDA.n5286 GNDA.n5284 0.563
R18405 GNDA.n1788 GNDA.n1786 0.464042
R18406 GNDA.n1742 GNDA.n1717 0.396333
R18407 GNDA.n7235 GNDA.n7234 0.369818
R18408 GNDA.n1763 GNDA.n1761 0.34425
R18409 GNDA.n1785 GNDA.n1702 0.34425
R18410 GNDA.n1726 GNDA.n590 0.313
R18411 GNDA.n1743 GNDA.n1724 0.292167
R18412 GNDA.n1757 GNDA.n1756 0.292167
R18413 GNDA.n1230 GNDA.n1227 0.28175
R18414 GNDA.n1237 GNDA.n1232 0.28175
R18415 GNDA.n1520 GNDA.n789 0.28175
R18416 GNDA.n1691 GNDA.n1522 0.28175
R18417 GNDA.n2281 GNDA.n2280 0.28175
R18418 GNDA.n2738 GNDA.n2569 0.28175
R18419 GNDA.n2742 GNDA.n2740 0.28175
R18420 GNDA.n3203 GNDA.n594 0.28175
R18421 GNDA.n5014 GNDA.n323 0.28175
R18422 GNDA.n5010 GNDA.n5009 0.28175
R18423 GNDA.n3682 GNDA.n3679 0.28175
R18424 GNDA.n4994 GNDA.n4993 0.28175
R18425 GNDA.n4982 GNDA.n4981 0.28175
R18426 GNDA.n4978 GNDA.n4977 0.28175
R18427 GNDA.n4974 GNDA.n4973 0.28175
R18428 GNDA.n4970 GNDA.n4969 0.28175
R18429 GNDA.n2109 GNDA.n2106 0.271333
R18430 GNDA GNDA.n6364 0.2565
R18431 GNDA GNDA.n6465 0.2565
R18432 GNDA.n6980 GNDA 0.2565
R18433 GNDA.n6800 GNDA 0.2565
R18434 GNDA.n5728 GNDA 0.2565
R18435 GNDA.n5490 GNDA 0.2565
R18436 GNDA.n5915 GNDA 0.2565
R18437 GNDA GNDA.n6758 0.2565
R18438 GNDA GNDA.n0 0.2565
R18439 GNDA.n6571 GNDA.n5409 0.255468
R18440 GNDA.n2916 GNDA.n320 0.224458
R18441 GNDA.n5280 GNDA.n324 0.21925
R18442 GNDA.n3387 GNDA.n3386 0.208833
R18443 GNDA.n1729 GNDA.n1728 0.208833
R18444 GNDA.n2104 GNDA.n723 0.198417
R18445 GNDA.n2567 GNDA.n660 0.198417
R18446 GNDA.n3380 GNDA.n3379 0.198417
R18447 GNDA.n5006 GNDA.n5005 0.198417
R18448 GNDA.n4998 GNDA.n4997 0.188
R18449 GNDA.n6949 GNDA.n6948 0.188
R18450 GNDA.n6944 GNDA.n6943 0.188
R18451 GNDA.n1770 GNDA.n1766 0.172375
R18452 GNDA.n1782 GNDA.n1781 0.172375
R18453 GNDA.n7043 GNDA.n7042 0.15675
R18454 GNDA.n7039 GNDA.n7038 0.15675
R18455 GNDA.n7048 GNDA.n7047 0.151542
R18456 GNDA.n6660 GNDA.n93 0.147453
R18457 GNDA.n5159 GNDA.n327 0.146333
R18458 GNDA.n5164 GNDA.n5159 0.146333
R18459 GNDA.n5165 GNDA.n5164 0.146333
R18460 GNDA.n5175 GNDA.n5174 0.146333
R18461 GNDA.n5178 GNDA.n5175 0.146333
R18462 GNDA.n5178 GNDA.n5155 0.146333
R18463 GNDA.n5188 GNDA.n5153 0.146333
R18464 GNDA.n5194 GNDA.n5153 0.146333
R18465 GNDA.n5195 GNDA.n5194 0.146333
R18466 GNDA.n5205 GNDA.n5204 0.146333
R18467 GNDA.n5208 GNDA.n5205 0.146333
R18468 GNDA.n5208 GNDA.n5149 0.146333
R18469 GNDA.n5218 GNDA.n5147 0.146333
R18470 GNDA.n5224 GNDA.n5147 0.146333
R18471 GNDA.n5225 GNDA.n5224 0.146333
R18472 GNDA.n5235 GNDA.n5234 0.146333
R18473 GNDA.n5238 GNDA.n5235 0.146333
R18474 GNDA.n5238 GNDA.n5143 0.146333
R18475 GNDA.n5248 GNDA.n5141 0.146333
R18476 GNDA.n5254 GNDA.n5141 0.146333
R18477 GNDA.n5255 GNDA.n5254 0.146333
R18478 GNDA.n5265 GNDA.n5264 0.146333
R18479 GNDA.n5268 GNDA.n5265 0.146333
R18480 GNDA.n5268 GNDA.n5137 0.146333
R18481 GNDA.n4846 GNDA.n3457 0.146333
R18482 GNDA.n4851 GNDA.n4846 0.146333
R18483 GNDA.n4852 GNDA.n4851 0.146333
R18484 GNDA.n4862 GNDA.n4861 0.146333
R18485 GNDA.n4865 GNDA.n4862 0.146333
R18486 GNDA.n4865 GNDA.n4842 0.146333
R18487 GNDA.n4875 GNDA.n4840 0.146333
R18488 GNDA.n4881 GNDA.n4840 0.146333
R18489 GNDA.n4882 GNDA.n4881 0.146333
R18490 GNDA.n4892 GNDA.n4891 0.146333
R18491 GNDA.n4895 GNDA.n4892 0.146333
R18492 GNDA.n4895 GNDA.n4836 0.146333
R18493 GNDA.n4905 GNDA.n4834 0.146333
R18494 GNDA.n4911 GNDA.n4834 0.146333
R18495 GNDA.n4912 GNDA.n4911 0.146333
R18496 GNDA.n4922 GNDA.n4921 0.146333
R18497 GNDA.n4925 GNDA.n4922 0.146333
R18498 GNDA.n4925 GNDA.n4830 0.146333
R18499 GNDA.n4935 GNDA.n4828 0.146333
R18500 GNDA.n4941 GNDA.n4828 0.146333
R18501 GNDA.n4942 GNDA.n4941 0.146333
R18502 GNDA.n4952 GNDA.n4951 0.146333
R18503 GNDA.n4955 GNDA.n4952 0.146333
R18504 GNDA.n4955 GNDA.n4824 0.146333
R18505 GNDA.n4685 GNDA.n4681 0.146333
R18506 GNDA.n4691 GNDA.n4681 0.146333
R18507 GNDA.n4692 GNDA.n4691 0.146333
R18508 GNDA.n4702 GNDA.n4701 0.146333
R18509 GNDA.n4705 GNDA.n4702 0.146333
R18510 GNDA.n4705 GNDA.n4677 0.146333
R18511 GNDA.n4715 GNDA.n4675 0.146333
R18512 GNDA.n4721 GNDA.n4675 0.146333
R18513 GNDA.n4722 GNDA.n4721 0.146333
R18514 GNDA.n4732 GNDA.n4731 0.146333
R18515 GNDA.n4735 GNDA.n4732 0.146333
R18516 GNDA.n4735 GNDA.n4671 0.146333
R18517 GNDA.n4745 GNDA.n4669 0.146333
R18518 GNDA.n4751 GNDA.n4669 0.146333
R18519 GNDA.n4752 GNDA.n4751 0.146333
R18520 GNDA.n4762 GNDA.n4761 0.146333
R18521 GNDA.n4765 GNDA.n4762 0.146333
R18522 GNDA.n4765 GNDA.n4665 0.146333
R18523 GNDA.n4775 GNDA.n4663 0.146333
R18524 GNDA.n4781 GNDA.n4663 0.146333
R18525 GNDA.n4782 GNDA.n4781 0.146333
R18526 GNDA.n4792 GNDA.n4791 0.146333
R18527 GNDA.n4795 GNDA.n4792 0.146333
R18528 GNDA.n4795 GNDA.n4659 0.146333
R18529 GNDA.n4519 GNDA.n4515 0.146333
R18530 GNDA.n4525 GNDA.n4515 0.146333
R18531 GNDA.n4526 GNDA.n4525 0.146333
R18532 GNDA.n4536 GNDA.n4535 0.146333
R18533 GNDA.n4539 GNDA.n4536 0.146333
R18534 GNDA.n4539 GNDA.n4511 0.146333
R18535 GNDA.n4549 GNDA.n4509 0.146333
R18536 GNDA.n4555 GNDA.n4509 0.146333
R18537 GNDA.n4556 GNDA.n4555 0.146333
R18538 GNDA.n4566 GNDA.n4565 0.146333
R18539 GNDA.n4569 GNDA.n4566 0.146333
R18540 GNDA.n4569 GNDA.n4505 0.146333
R18541 GNDA.n4579 GNDA.n4503 0.146333
R18542 GNDA.n4585 GNDA.n4503 0.146333
R18543 GNDA.n4586 GNDA.n4585 0.146333
R18544 GNDA.n4596 GNDA.n4595 0.146333
R18545 GNDA.n4599 GNDA.n4596 0.146333
R18546 GNDA.n4599 GNDA.n4499 0.146333
R18547 GNDA.n4609 GNDA.n4497 0.146333
R18548 GNDA.n4615 GNDA.n4497 0.146333
R18549 GNDA.n4616 GNDA.n4615 0.146333
R18550 GNDA.n4626 GNDA.n4625 0.146333
R18551 GNDA.n4629 GNDA.n4626 0.146333
R18552 GNDA.n4629 GNDA.n4493 0.146333
R18553 GNDA.n4353 GNDA.n4349 0.146333
R18554 GNDA.n4359 GNDA.n4349 0.146333
R18555 GNDA.n4360 GNDA.n4359 0.146333
R18556 GNDA.n4370 GNDA.n4369 0.146333
R18557 GNDA.n4373 GNDA.n4370 0.146333
R18558 GNDA.n4373 GNDA.n4345 0.146333
R18559 GNDA.n4383 GNDA.n4343 0.146333
R18560 GNDA.n4389 GNDA.n4343 0.146333
R18561 GNDA.n4390 GNDA.n4389 0.146333
R18562 GNDA.n4400 GNDA.n4399 0.146333
R18563 GNDA.n4403 GNDA.n4400 0.146333
R18564 GNDA.n4403 GNDA.n4339 0.146333
R18565 GNDA.n4413 GNDA.n4337 0.146333
R18566 GNDA.n4419 GNDA.n4337 0.146333
R18567 GNDA.n4420 GNDA.n4419 0.146333
R18568 GNDA.n4430 GNDA.n4429 0.146333
R18569 GNDA.n4433 GNDA.n4430 0.146333
R18570 GNDA.n4433 GNDA.n4333 0.146333
R18571 GNDA.n4443 GNDA.n4331 0.146333
R18572 GNDA.n4449 GNDA.n4331 0.146333
R18573 GNDA.n4450 GNDA.n4449 0.146333
R18574 GNDA.n4460 GNDA.n4459 0.146333
R18575 GNDA.n4463 GNDA.n4460 0.146333
R18576 GNDA.n4463 GNDA.n4327 0.146333
R18577 GNDA.n4187 GNDA.n4183 0.146333
R18578 GNDA.n4193 GNDA.n4183 0.146333
R18579 GNDA.n4194 GNDA.n4193 0.146333
R18580 GNDA.n4204 GNDA.n4203 0.146333
R18581 GNDA.n4207 GNDA.n4204 0.146333
R18582 GNDA.n4207 GNDA.n4179 0.146333
R18583 GNDA.n4217 GNDA.n4177 0.146333
R18584 GNDA.n4223 GNDA.n4177 0.146333
R18585 GNDA.n4224 GNDA.n4223 0.146333
R18586 GNDA.n4234 GNDA.n4233 0.146333
R18587 GNDA.n4237 GNDA.n4234 0.146333
R18588 GNDA.n4237 GNDA.n4173 0.146333
R18589 GNDA.n4247 GNDA.n4171 0.146333
R18590 GNDA.n4253 GNDA.n4171 0.146333
R18591 GNDA.n4254 GNDA.n4253 0.146333
R18592 GNDA.n4264 GNDA.n4263 0.146333
R18593 GNDA.n4267 GNDA.n4264 0.146333
R18594 GNDA.n4267 GNDA.n4167 0.146333
R18595 GNDA.n4277 GNDA.n4165 0.146333
R18596 GNDA.n4283 GNDA.n4165 0.146333
R18597 GNDA.n4284 GNDA.n4283 0.146333
R18598 GNDA.n4294 GNDA.n4293 0.146333
R18599 GNDA.n4297 GNDA.n4294 0.146333
R18600 GNDA.n4297 GNDA.n4161 0.146333
R18601 GNDA.n3689 GNDA.n3507 0.146333
R18602 GNDA.n3695 GNDA.n3507 0.146333
R18603 GNDA.n3696 GNDA.n3695 0.146333
R18604 GNDA.n3706 GNDA.n3705 0.146333
R18605 GNDA.n3709 GNDA.n3706 0.146333
R18606 GNDA.n3709 GNDA.n3503 0.146333
R18607 GNDA.n3719 GNDA.n3501 0.146333
R18608 GNDA.n3725 GNDA.n3501 0.146333
R18609 GNDA.n3726 GNDA.n3725 0.146333
R18610 GNDA.n3736 GNDA.n3735 0.146333
R18611 GNDA.n3739 GNDA.n3736 0.146333
R18612 GNDA.n3739 GNDA.n3497 0.146333
R18613 GNDA.n3749 GNDA.n3495 0.146333
R18614 GNDA.n3755 GNDA.n3495 0.146333
R18615 GNDA.n3756 GNDA.n3755 0.146333
R18616 GNDA.n3766 GNDA.n3765 0.146333
R18617 GNDA.n3769 GNDA.n3766 0.146333
R18618 GNDA.n3769 GNDA.n3491 0.146333
R18619 GNDA.n3779 GNDA.n3489 0.146333
R18620 GNDA.n3785 GNDA.n3489 0.146333
R18621 GNDA.n3786 GNDA.n3785 0.146333
R18622 GNDA.n3796 GNDA.n3795 0.146333
R18623 GNDA.n3799 GNDA.n3796 0.146333
R18624 GNDA.n3799 GNDA.n3485 0.146333
R18625 GNDA.n4021 GNDA.n4017 0.146333
R18626 GNDA.n4027 GNDA.n4017 0.146333
R18627 GNDA.n4028 GNDA.n4027 0.146333
R18628 GNDA.n4038 GNDA.n4037 0.146333
R18629 GNDA.n4041 GNDA.n4038 0.146333
R18630 GNDA.n4041 GNDA.n4013 0.146333
R18631 GNDA.n4051 GNDA.n4011 0.146333
R18632 GNDA.n4057 GNDA.n4011 0.146333
R18633 GNDA.n4058 GNDA.n4057 0.146333
R18634 GNDA.n4068 GNDA.n4067 0.146333
R18635 GNDA.n4071 GNDA.n4068 0.146333
R18636 GNDA.n4071 GNDA.n4007 0.146333
R18637 GNDA.n4081 GNDA.n4005 0.146333
R18638 GNDA.n4087 GNDA.n4005 0.146333
R18639 GNDA.n4088 GNDA.n4087 0.146333
R18640 GNDA.n4098 GNDA.n4097 0.146333
R18641 GNDA.n4101 GNDA.n4098 0.146333
R18642 GNDA.n4101 GNDA.n4001 0.146333
R18643 GNDA.n4111 GNDA.n3999 0.146333
R18644 GNDA.n4117 GNDA.n3999 0.146333
R18645 GNDA.n4118 GNDA.n4117 0.146333
R18646 GNDA.n4128 GNDA.n4127 0.146333
R18647 GNDA.n4131 GNDA.n4128 0.146333
R18648 GNDA.n4131 GNDA.n3995 0.146333
R18649 GNDA.n3855 GNDA.n3851 0.146333
R18650 GNDA.n3861 GNDA.n3851 0.146333
R18651 GNDA.n3862 GNDA.n3861 0.146333
R18652 GNDA.n3872 GNDA.n3871 0.146333
R18653 GNDA.n3875 GNDA.n3872 0.146333
R18654 GNDA.n3875 GNDA.n3847 0.146333
R18655 GNDA.n3885 GNDA.n3845 0.146333
R18656 GNDA.n3891 GNDA.n3845 0.146333
R18657 GNDA.n3892 GNDA.n3891 0.146333
R18658 GNDA.n3902 GNDA.n3901 0.146333
R18659 GNDA.n3905 GNDA.n3902 0.146333
R18660 GNDA.n3905 GNDA.n3841 0.146333
R18661 GNDA.n3915 GNDA.n3839 0.146333
R18662 GNDA.n3921 GNDA.n3839 0.146333
R18663 GNDA.n3922 GNDA.n3921 0.146333
R18664 GNDA.n3932 GNDA.n3931 0.146333
R18665 GNDA.n3935 GNDA.n3932 0.146333
R18666 GNDA.n3935 GNDA.n3835 0.146333
R18667 GNDA.n3945 GNDA.n3833 0.146333
R18668 GNDA.n3951 GNDA.n3833 0.146333
R18669 GNDA.n3952 GNDA.n3951 0.146333
R18670 GNDA.n3962 GNDA.n3961 0.146333
R18671 GNDA.n3965 GNDA.n3962 0.146333
R18672 GNDA.n3965 GNDA.n3829 0.146333
R18673 GNDA.n3513 GNDA.n3512 0.146333
R18674 GNDA.n3514 GNDA.n3513 0.146333
R18675 GNDA.n3515 GNDA.n3514 0.146333
R18676 GNDA.n3519 GNDA.n3518 0.146333
R18677 GNDA.n3520 GNDA.n3519 0.146333
R18678 GNDA.n3521 GNDA.n3520 0.146333
R18679 GNDA.n3525 GNDA.n3524 0.146333
R18680 GNDA.n3526 GNDA.n3525 0.146333
R18681 GNDA.n3527 GNDA.n3526 0.146333
R18682 GNDA.n3531 GNDA.n3530 0.146333
R18683 GNDA.n3532 GNDA.n3531 0.146333
R18684 GNDA.n3533 GNDA.n3532 0.146333
R18685 GNDA.n3537 GNDA.n3536 0.146333
R18686 GNDA.n3538 GNDA.n3537 0.146333
R18687 GNDA.n3539 GNDA.n3538 0.146333
R18688 GNDA.n3543 GNDA.n3542 0.146333
R18689 GNDA.n3544 GNDA.n3543 0.146333
R18690 GNDA.n3545 GNDA.n3544 0.146333
R18691 GNDA.n3549 GNDA.n3548 0.146333
R18692 GNDA.n3550 GNDA.n3549 0.146333
R18693 GNDA.n3551 GNDA.n3550 0.146333
R18694 GNDA.n3555 GNDA.n3554 0.146333
R18695 GNDA.n3556 GNDA.n3555 0.146333
R18696 GNDA.n3557 GNDA.n3556 0.146333
R18697 GNDA.n407 GNDA.n406 0.146333
R18698 GNDA.n408 GNDA.n407 0.146333
R18699 GNDA.n409 GNDA.n408 0.146333
R18700 GNDA.n413 GNDA.n412 0.146333
R18701 GNDA.n414 GNDA.n413 0.146333
R18702 GNDA.n415 GNDA.n414 0.146333
R18703 GNDA.n419 GNDA.n418 0.146333
R18704 GNDA.n420 GNDA.n419 0.146333
R18705 GNDA.n421 GNDA.n420 0.146333
R18706 GNDA.n425 GNDA.n424 0.146333
R18707 GNDA.n426 GNDA.n425 0.146333
R18708 GNDA.n427 GNDA.n426 0.146333
R18709 GNDA.n431 GNDA.n430 0.146333
R18710 GNDA.n432 GNDA.n431 0.146333
R18711 GNDA.n433 GNDA.n432 0.146333
R18712 GNDA.n437 GNDA.n436 0.146333
R18713 GNDA.n438 GNDA.n437 0.146333
R18714 GNDA.n439 GNDA.n438 0.146333
R18715 GNDA.n443 GNDA.n442 0.146333
R18716 GNDA.n444 GNDA.n443 0.146333
R18717 GNDA.n445 GNDA.n444 0.146333
R18718 GNDA.n449 GNDA.n448 0.146333
R18719 GNDA.n450 GNDA.n449 0.146333
R18720 GNDA.n451 GNDA.n450 0.146333
R18721 GNDA.n5021 GNDA.n401 0.146333
R18722 GNDA.n5027 GNDA.n401 0.146333
R18723 GNDA.n5028 GNDA.n5027 0.146333
R18724 GNDA.n5038 GNDA.n5037 0.146333
R18725 GNDA.n5041 GNDA.n5038 0.146333
R18726 GNDA.n5041 GNDA.n397 0.146333
R18727 GNDA.n5051 GNDA.n395 0.146333
R18728 GNDA.n5057 GNDA.n395 0.146333
R18729 GNDA.n5058 GNDA.n5057 0.146333
R18730 GNDA.n5068 GNDA.n5067 0.146333
R18731 GNDA.n5071 GNDA.n5068 0.146333
R18732 GNDA.n5071 GNDA.n391 0.146333
R18733 GNDA.n5081 GNDA.n389 0.146333
R18734 GNDA.n5087 GNDA.n389 0.146333
R18735 GNDA.n5088 GNDA.n5087 0.146333
R18736 GNDA.n5098 GNDA.n5097 0.146333
R18737 GNDA.n5101 GNDA.n5098 0.146333
R18738 GNDA.n5101 GNDA.n385 0.146333
R18739 GNDA.n5111 GNDA.n383 0.146333
R18740 GNDA.n5117 GNDA.n383 0.146333
R18741 GNDA.n5118 GNDA.n5117 0.146333
R18742 GNDA.n5128 GNDA.n5127 0.146333
R18743 GNDA.n5131 GNDA.n5128 0.146333
R18744 GNDA.n5131 GNDA.n379 0.146333
R18745 GNDA.n3210 GNDA.n3209 0.146333
R18746 GNDA.n3211 GNDA.n3210 0.146333
R18747 GNDA.n3212 GNDA.n3211 0.146333
R18748 GNDA.n3216 GNDA.n3215 0.146333
R18749 GNDA.n3217 GNDA.n3216 0.146333
R18750 GNDA.n3218 GNDA.n3217 0.146333
R18751 GNDA.n3222 GNDA.n3221 0.146333
R18752 GNDA.n3223 GNDA.n3222 0.146333
R18753 GNDA.n3224 GNDA.n3223 0.146333
R18754 GNDA.n3228 GNDA.n3227 0.146333
R18755 GNDA.n3229 GNDA.n3228 0.146333
R18756 GNDA.n3230 GNDA.n3229 0.146333
R18757 GNDA.n3234 GNDA.n3233 0.146333
R18758 GNDA.n3235 GNDA.n3234 0.146333
R18759 GNDA.n3236 GNDA.n3235 0.146333
R18760 GNDA.n3240 GNDA.n3239 0.146333
R18761 GNDA.n3241 GNDA.n3240 0.146333
R18762 GNDA.n3242 GNDA.n3241 0.146333
R18763 GNDA.n3246 GNDA.n3245 0.146333
R18764 GNDA.n3247 GNDA.n3246 0.146333
R18765 GNDA.n3248 GNDA.n3247 0.146333
R18766 GNDA.n3252 GNDA.n3251 0.146333
R18767 GNDA.n3253 GNDA.n3252 0.146333
R18768 GNDA.n3254 GNDA.n3253 0.146333
R18769 GNDA.n3084 GNDA.n597 0.146333
R18770 GNDA.n3089 GNDA.n3084 0.146333
R18771 GNDA.n3090 GNDA.n3089 0.146333
R18772 GNDA.n3100 GNDA.n3099 0.146333
R18773 GNDA.n3103 GNDA.n3100 0.146333
R18774 GNDA.n3103 GNDA.n3080 0.146333
R18775 GNDA.n3113 GNDA.n3078 0.146333
R18776 GNDA.n3119 GNDA.n3078 0.146333
R18777 GNDA.n3120 GNDA.n3119 0.146333
R18778 GNDA.n3130 GNDA.n3129 0.146333
R18779 GNDA.n3133 GNDA.n3130 0.146333
R18780 GNDA.n3133 GNDA.n3074 0.146333
R18781 GNDA.n3143 GNDA.n3072 0.146333
R18782 GNDA.n3149 GNDA.n3072 0.146333
R18783 GNDA.n3150 GNDA.n3149 0.146333
R18784 GNDA.n3160 GNDA.n3159 0.146333
R18785 GNDA.n3163 GNDA.n3160 0.146333
R18786 GNDA.n3163 GNDA.n3068 0.146333
R18787 GNDA.n3173 GNDA.n3066 0.146333
R18788 GNDA.n3179 GNDA.n3066 0.146333
R18789 GNDA.n3180 GNDA.n3179 0.146333
R18790 GNDA.n3190 GNDA.n3189 0.146333
R18791 GNDA.n3193 GNDA.n3190 0.146333
R18792 GNDA.n3193 GNDA.n3062 0.146333
R18793 GNDA.n2923 GNDA.n2911 0.146333
R18794 GNDA.n2929 GNDA.n2911 0.146333
R18795 GNDA.n2930 GNDA.n2929 0.146333
R18796 GNDA.n2940 GNDA.n2939 0.146333
R18797 GNDA.n2943 GNDA.n2940 0.146333
R18798 GNDA.n2943 GNDA.n2907 0.146333
R18799 GNDA.n2953 GNDA.n2905 0.146333
R18800 GNDA.n2959 GNDA.n2905 0.146333
R18801 GNDA.n2960 GNDA.n2959 0.146333
R18802 GNDA.n2970 GNDA.n2969 0.146333
R18803 GNDA.n2973 GNDA.n2970 0.146333
R18804 GNDA.n2973 GNDA.n2901 0.146333
R18805 GNDA.n2983 GNDA.n2899 0.146333
R18806 GNDA.n2989 GNDA.n2899 0.146333
R18807 GNDA.n2990 GNDA.n2989 0.146333
R18808 GNDA.n3000 GNDA.n2999 0.146333
R18809 GNDA.n3003 GNDA.n3000 0.146333
R18810 GNDA.n3003 GNDA.n2895 0.146333
R18811 GNDA.n3013 GNDA.n2893 0.146333
R18812 GNDA.n3019 GNDA.n2893 0.146333
R18813 GNDA.n3020 GNDA.n3019 0.146333
R18814 GNDA.n3030 GNDA.n3029 0.146333
R18815 GNDA.n3033 GNDA.n3030 0.146333
R18816 GNDA.n3033 GNDA.n2889 0.146333
R18817 GNDA.n2287 GNDA.n713 0.146333
R18818 GNDA.n2293 GNDA.n713 0.146333
R18819 GNDA.n2294 GNDA.n2293 0.146333
R18820 GNDA.n2304 GNDA.n2303 0.146333
R18821 GNDA.n2307 GNDA.n2304 0.146333
R18822 GNDA.n2307 GNDA.n709 0.146333
R18823 GNDA.n2317 GNDA.n707 0.146333
R18824 GNDA.n2323 GNDA.n707 0.146333
R18825 GNDA.n2324 GNDA.n2323 0.146333
R18826 GNDA.n2334 GNDA.n2333 0.146333
R18827 GNDA.n2337 GNDA.n2334 0.146333
R18828 GNDA.n2337 GNDA.n703 0.146333
R18829 GNDA.n2347 GNDA.n701 0.146333
R18830 GNDA.n2353 GNDA.n701 0.146333
R18831 GNDA.n2354 GNDA.n2353 0.146333
R18832 GNDA.n2364 GNDA.n2363 0.146333
R18833 GNDA.n2367 GNDA.n2364 0.146333
R18834 GNDA.n2367 GNDA.n697 0.146333
R18835 GNDA.n2377 GNDA.n695 0.146333
R18836 GNDA.n2383 GNDA.n695 0.146333
R18837 GNDA.n2384 GNDA.n2383 0.146333
R18838 GNDA.n2394 GNDA.n2393 0.146333
R18839 GNDA.n2397 GNDA.n2394 0.146333
R18840 GNDA.n2397 GNDA.n691 0.146333
R18841 GNDA.n2749 GNDA.n647 0.146333
R18842 GNDA.n2755 GNDA.n647 0.146333
R18843 GNDA.n2756 GNDA.n2755 0.146333
R18844 GNDA.n2766 GNDA.n2765 0.146333
R18845 GNDA.n2769 GNDA.n2766 0.146333
R18846 GNDA.n2769 GNDA.n643 0.146333
R18847 GNDA.n2779 GNDA.n641 0.146333
R18848 GNDA.n2785 GNDA.n641 0.146333
R18849 GNDA.n2786 GNDA.n2785 0.146333
R18850 GNDA.n2796 GNDA.n2795 0.146333
R18851 GNDA.n2799 GNDA.n2796 0.146333
R18852 GNDA.n2799 GNDA.n637 0.146333
R18853 GNDA.n2809 GNDA.n635 0.146333
R18854 GNDA.n2815 GNDA.n635 0.146333
R18855 GNDA.n2816 GNDA.n2815 0.146333
R18856 GNDA.n2826 GNDA.n2825 0.146333
R18857 GNDA.n2829 GNDA.n2826 0.146333
R18858 GNDA.n2829 GNDA.n631 0.146333
R18859 GNDA.n2839 GNDA.n629 0.146333
R18860 GNDA.n2845 GNDA.n629 0.146333
R18861 GNDA.n2846 GNDA.n2845 0.146333
R18862 GNDA.n2856 GNDA.n2855 0.146333
R18863 GNDA.n2859 GNDA.n2856 0.146333
R18864 GNDA.n2859 GNDA.n625 0.146333
R18865 GNDA.n2573 GNDA.n2572 0.146333
R18866 GNDA.n2574 GNDA.n2573 0.146333
R18867 GNDA.n2575 GNDA.n2574 0.146333
R18868 GNDA.n2579 GNDA.n2578 0.146333
R18869 GNDA.n2580 GNDA.n2579 0.146333
R18870 GNDA.n2581 GNDA.n2580 0.146333
R18871 GNDA.n2585 GNDA.n2584 0.146333
R18872 GNDA.n2586 GNDA.n2585 0.146333
R18873 GNDA.n2587 GNDA.n2586 0.146333
R18874 GNDA.n2591 GNDA.n2590 0.146333
R18875 GNDA.n2592 GNDA.n2591 0.146333
R18876 GNDA.n2593 GNDA.n2592 0.146333
R18877 GNDA.n2597 GNDA.n2596 0.146333
R18878 GNDA.n2598 GNDA.n2597 0.146333
R18879 GNDA.n2599 GNDA.n2598 0.146333
R18880 GNDA.n2603 GNDA.n2602 0.146333
R18881 GNDA.n2604 GNDA.n2603 0.146333
R18882 GNDA.n2605 GNDA.n2604 0.146333
R18883 GNDA.n2609 GNDA.n2608 0.146333
R18884 GNDA.n2610 GNDA.n2609 0.146333
R18885 GNDA.n2611 GNDA.n2610 0.146333
R18886 GNDA.n2615 GNDA.n2614 0.146333
R18887 GNDA.n2616 GNDA.n2615 0.146333
R18888 GNDA.n2617 GNDA.n2616 0.146333
R18889 GNDA.n2448 GNDA.n663 0.146333
R18890 GNDA.n2453 GNDA.n2448 0.146333
R18891 GNDA.n2454 GNDA.n2453 0.146333
R18892 GNDA.n2464 GNDA.n2463 0.146333
R18893 GNDA.n2467 GNDA.n2464 0.146333
R18894 GNDA.n2467 GNDA.n2444 0.146333
R18895 GNDA.n2477 GNDA.n2442 0.146333
R18896 GNDA.n2483 GNDA.n2442 0.146333
R18897 GNDA.n2484 GNDA.n2483 0.146333
R18898 GNDA.n2494 GNDA.n2493 0.146333
R18899 GNDA.n2497 GNDA.n2494 0.146333
R18900 GNDA.n2497 GNDA.n2438 0.146333
R18901 GNDA.n2507 GNDA.n2436 0.146333
R18902 GNDA.n2513 GNDA.n2436 0.146333
R18903 GNDA.n2514 GNDA.n2513 0.146333
R18904 GNDA.n2524 GNDA.n2523 0.146333
R18905 GNDA.n2527 GNDA.n2524 0.146333
R18906 GNDA.n2527 GNDA.n2432 0.146333
R18907 GNDA.n2537 GNDA.n2430 0.146333
R18908 GNDA.n2543 GNDA.n2430 0.146333
R18909 GNDA.n2544 GNDA.n2543 0.146333
R18910 GNDA.n2554 GNDA.n2553 0.146333
R18911 GNDA.n2557 GNDA.n2554 0.146333
R18912 GNDA.n2557 GNDA.n2426 0.146333
R18913 GNDA.n2113 GNDA.n2112 0.146333
R18914 GNDA.n2114 GNDA.n2113 0.146333
R18915 GNDA.n2115 GNDA.n2114 0.146333
R18916 GNDA.n2119 GNDA.n2118 0.146333
R18917 GNDA.n2120 GNDA.n2119 0.146333
R18918 GNDA.n2121 GNDA.n2120 0.146333
R18919 GNDA.n2125 GNDA.n2124 0.146333
R18920 GNDA.n2126 GNDA.n2125 0.146333
R18921 GNDA.n2127 GNDA.n2126 0.146333
R18922 GNDA.n2131 GNDA.n2130 0.146333
R18923 GNDA.n2132 GNDA.n2131 0.146333
R18924 GNDA.n2133 GNDA.n2132 0.146333
R18925 GNDA.n2137 GNDA.n2136 0.146333
R18926 GNDA.n2138 GNDA.n2137 0.146333
R18927 GNDA.n2139 GNDA.n2138 0.146333
R18928 GNDA.n2143 GNDA.n2142 0.146333
R18929 GNDA.n2144 GNDA.n2143 0.146333
R18930 GNDA.n2145 GNDA.n2144 0.146333
R18931 GNDA.n2149 GNDA.n2148 0.146333
R18932 GNDA.n2150 GNDA.n2149 0.146333
R18933 GNDA.n2151 GNDA.n2150 0.146333
R18934 GNDA.n2155 GNDA.n2154 0.146333
R18935 GNDA.n2156 GNDA.n2155 0.146333
R18936 GNDA.n2157 GNDA.n2156 0.146333
R18937 GNDA.n1985 GNDA.n726 0.146333
R18938 GNDA.n1990 GNDA.n1985 0.146333
R18939 GNDA.n1991 GNDA.n1990 0.146333
R18940 GNDA.n2001 GNDA.n2000 0.146333
R18941 GNDA.n2004 GNDA.n2001 0.146333
R18942 GNDA.n2004 GNDA.n1981 0.146333
R18943 GNDA.n2014 GNDA.n1979 0.146333
R18944 GNDA.n2020 GNDA.n1979 0.146333
R18945 GNDA.n2021 GNDA.n2020 0.146333
R18946 GNDA.n2031 GNDA.n2030 0.146333
R18947 GNDA.n2034 GNDA.n2031 0.146333
R18948 GNDA.n2034 GNDA.n1975 0.146333
R18949 GNDA.n2044 GNDA.n1973 0.146333
R18950 GNDA.n2050 GNDA.n1973 0.146333
R18951 GNDA.n2051 GNDA.n2050 0.146333
R18952 GNDA.n2061 GNDA.n2060 0.146333
R18953 GNDA.n2064 GNDA.n2061 0.146333
R18954 GNDA.n2064 GNDA.n1969 0.146333
R18955 GNDA.n2074 GNDA.n1967 0.146333
R18956 GNDA.n2080 GNDA.n1967 0.146333
R18957 GNDA.n2081 GNDA.n2080 0.146333
R18958 GNDA.n2091 GNDA.n2090 0.146333
R18959 GNDA.n2094 GNDA.n2091 0.146333
R18960 GNDA.n2094 GNDA.n1963 0.146333
R18961 GNDA.n1824 GNDA.n776 0.146333
R18962 GNDA.n1830 GNDA.n776 0.146333
R18963 GNDA.n1831 GNDA.n1830 0.146333
R18964 GNDA.n1841 GNDA.n1840 0.146333
R18965 GNDA.n1844 GNDA.n1841 0.146333
R18966 GNDA.n1844 GNDA.n772 0.146333
R18967 GNDA.n1854 GNDA.n770 0.146333
R18968 GNDA.n1860 GNDA.n770 0.146333
R18969 GNDA.n1861 GNDA.n1860 0.146333
R18970 GNDA.n1871 GNDA.n1870 0.146333
R18971 GNDA.n1874 GNDA.n1871 0.146333
R18972 GNDA.n1874 GNDA.n766 0.146333
R18973 GNDA.n1884 GNDA.n764 0.146333
R18974 GNDA.n1890 GNDA.n764 0.146333
R18975 GNDA.n1891 GNDA.n1890 0.146333
R18976 GNDA.n1901 GNDA.n1900 0.146333
R18977 GNDA.n1904 GNDA.n1901 0.146333
R18978 GNDA.n1904 GNDA.n760 0.146333
R18979 GNDA.n1914 GNDA.n758 0.146333
R18980 GNDA.n1920 GNDA.n758 0.146333
R18981 GNDA.n1921 GNDA.n1920 0.146333
R18982 GNDA.n1931 GNDA.n1930 0.146333
R18983 GNDA.n1934 GNDA.n1931 0.146333
R18984 GNDA.n1934 GNDA.n754 0.146333
R18985 GNDA.n1526 GNDA.n1525 0.146333
R18986 GNDA.n1527 GNDA.n1526 0.146333
R18987 GNDA.n1528 GNDA.n1527 0.146333
R18988 GNDA.n1532 GNDA.n1531 0.146333
R18989 GNDA.n1533 GNDA.n1532 0.146333
R18990 GNDA.n1534 GNDA.n1533 0.146333
R18991 GNDA.n1538 GNDA.n1537 0.146333
R18992 GNDA.n1539 GNDA.n1538 0.146333
R18993 GNDA.n1540 GNDA.n1539 0.146333
R18994 GNDA.n1544 GNDA.n1543 0.146333
R18995 GNDA.n1545 GNDA.n1544 0.146333
R18996 GNDA.n1546 GNDA.n1545 0.146333
R18997 GNDA.n1550 GNDA.n1549 0.146333
R18998 GNDA.n1551 GNDA.n1550 0.146333
R18999 GNDA.n1552 GNDA.n1551 0.146333
R19000 GNDA.n1556 GNDA.n1555 0.146333
R19001 GNDA.n1557 GNDA.n1556 0.146333
R19002 GNDA.n1558 GNDA.n1557 0.146333
R19003 GNDA.n1562 GNDA.n1561 0.146333
R19004 GNDA.n1563 GNDA.n1562 0.146333
R19005 GNDA.n1564 GNDA.n1563 0.146333
R19006 GNDA.n1568 GNDA.n1567 0.146333
R19007 GNDA.n1569 GNDA.n1568 0.146333
R19008 GNDA.n1570 GNDA.n1569 0.146333
R19009 GNDA.n1401 GNDA.n792 0.146333
R19010 GNDA.n1406 GNDA.n1401 0.146333
R19011 GNDA.n1407 GNDA.n1406 0.146333
R19012 GNDA.n1417 GNDA.n1416 0.146333
R19013 GNDA.n1420 GNDA.n1417 0.146333
R19014 GNDA.n1420 GNDA.n1397 0.146333
R19015 GNDA.n1430 GNDA.n1395 0.146333
R19016 GNDA.n1436 GNDA.n1395 0.146333
R19017 GNDA.n1437 GNDA.n1436 0.146333
R19018 GNDA.n1447 GNDA.n1446 0.146333
R19019 GNDA.n1450 GNDA.n1447 0.146333
R19020 GNDA.n1450 GNDA.n1391 0.146333
R19021 GNDA.n1460 GNDA.n1389 0.146333
R19022 GNDA.n1466 GNDA.n1389 0.146333
R19023 GNDA.n1467 GNDA.n1466 0.146333
R19024 GNDA.n1477 GNDA.n1476 0.146333
R19025 GNDA.n1480 GNDA.n1477 0.146333
R19026 GNDA.n1480 GNDA.n1385 0.146333
R19027 GNDA.n1490 GNDA.n1383 0.146333
R19028 GNDA.n1496 GNDA.n1383 0.146333
R19029 GNDA.n1497 GNDA.n1496 0.146333
R19030 GNDA.n1507 GNDA.n1506 0.146333
R19031 GNDA.n1510 GNDA.n1507 0.146333
R19032 GNDA.n1510 GNDA.n1379 0.146333
R19033 GNDA.n1244 GNDA.n1241 0.146333
R19034 GNDA.n1247 GNDA.n1244 0.146333
R19035 GNDA.n1247 GNDA.n1213 0.146333
R19036 GNDA.n1257 GNDA.n1211 0.146333
R19037 GNDA.n1261 GNDA.n1211 0.146333
R19038 GNDA.n1264 GNDA.n1261 0.146333
R19039 GNDA.n1274 GNDA.n1271 0.146333
R19040 GNDA.n1277 GNDA.n1274 0.146333
R19041 GNDA.n1277 GNDA.n1207 0.146333
R19042 GNDA.n1287 GNDA.n1205 0.146333
R19043 GNDA.n1291 GNDA.n1205 0.146333
R19044 GNDA.n1294 GNDA.n1291 0.146333
R19045 GNDA.n1304 GNDA.n1301 0.146333
R19046 GNDA.n1307 GNDA.n1304 0.146333
R19047 GNDA.n1307 GNDA.n1201 0.146333
R19048 GNDA.n1317 GNDA.n1199 0.146333
R19049 GNDA.n1321 GNDA.n1199 0.146333
R19050 GNDA.n1324 GNDA.n1321 0.146333
R19051 GNDA.n1334 GNDA.n1331 0.146333
R19052 GNDA.n1337 GNDA.n1334 0.146333
R19053 GNDA.n1337 GNDA.n1195 0.146333
R19054 GNDA.n1346 GNDA.n1192 0.146333
R19055 GNDA.n1351 GNDA.n1192 0.146333
R19056 GNDA.n1351 GNDA.n1193 0.146333
R19057 GNDA.n7135 GNDA.n7134 0.146333
R19058 GNDA.n7138 GNDA.n7135 0.146333
R19059 GNDA.n7138 GNDA.n7128 0.146333
R19060 GNDA.n7146 GNDA.n7124 0.146333
R19061 GNDA.n7150 GNDA.n7124 0.146333
R19062 GNDA.n7151 GNDA.n7150 0.146333
R19063 GNDA.n7159 GNDA.n7158 0.146333
R19064 GNDA.n7162 GNDA.n7159 0.146333
R19065 GNDA.n7162 GNDA.n7116 0.146333
R19066 GNDA.n7170 GNDA.n7112 0.146333
R19067 GNDA.n7174 GNDA.n7112 0.146333
R19068 GNDA.n7175 GNDA.n7174 0.146333
R19069 GNDA.n7183 GNDA.n7182 0.146333
R19070 GNDA.n7186 GNDA.n7183 0.146333
R19071 GNDA.n7186 GNDA.n7104 0.146333
R19072 GNDA.n7194 GNDA.n7100 0.146333
R19073 GNDA.n7198 GNDA.n7100 0.146333
R19074 GNDA.n7199 GNDA.n7198 0.146333
R19075 GNDA.n7207 GNDA.n7206 0.146333
R19076 GNDA.n7210 GNDA.n7207 0.146333
R19077 GNDA.n7210 GNDA.n7092 0.146333
R19078 GNDA.n7218 GNDA.n7090 0.146333
R19079 GNDA.n7222 GNDA.n7090 0.146333
R19080 GNDA.n7222 GNDA.n96 0.146333
R19081 GNDA.n151 GNDA.n150 0.146333
R19082 GNDA.n151 GNDA.n145 0.146333
R19083 GNDA.n161 GNDA.n143 0.146333
R19084 GNDA.n169 GNDA.n143 0.146333
R19085 GNDA.n170 GNDA.n169 0.146333
R19086 GNDA.n180 GNDA.n179 0.146333
R19087 GNDA.n181 GNDA.n180 0.146333
R19088 GNDA.n181 GNDA.n139 0.146333
R19089 GNDA.n191 GNDA.n137 0.146333
R19090 GNDA.n199 GNDA.n137 0.146333
R19091 GNDA.n200 GNDA.n199 0.146333
R19092 GNDA.n210 GNDA.n209 0.146333
R19093 GNDA.n211 GNDA.n210 0.146333
R19094 GNDA.n211 GNDA.n133 0.146333
R19095 GNDA.n221 GNDA.n131 0.146333
R19096 GNDA.n229 GNDA.n131 0.146333
R19097 GNDA.n230 GNDA.n229 0.146333
R19098 GNDA.n240 GNDA.n239 0.146333
R19099 GNDA.n241 GNDA.n240 0.146333
R19100 GNDA.n241 GNDA.n127 0.146333
R19101 GNDA.n251 GNDA.n125 0.146333
R19102 GNDA.n259 GNDA.n125 0.146333
R19103 GNDA.n260 GNDA.n259 0.146333
R19104 GNDA.n148 GNDA.n146 0.146333
R19105 GNDA.n154 GNDA.n146 0.146333
R19106 GNDA.n155 GNDA.n154 0.146333
R19107 GNDA.n165 GNDA.n164 0.146333
R19108 GNDA.n168 GNDA.n165 0.146333
R19109 GNDA.n168 GNDA.n142 0.146333
R19110 GNDA.n178 GNDA.n140 0.146333
R19111 GNDA.n184 GNDA.n140 0.146333
R19112 GNDA.n185 GNDA.n184 0.146333
R19113 GNDA.n195 GNDA.n194 0.146333
R19114 GNDA.n198 GNDA.n195 0.146333
R19115 GNDA.n198 GNDA.n136 0.146333
R19116 GNDA.n208 GNDA.n134 0.146333
R19117 GNDA.n214 GNDA.n134 0.146333
R19118 GNDA.n215 GNDA.n214 0.146333
R19119 GNDA.n225 GNDA.n224 0.146333
R19120 GNDA.n228 GNDA.n225 0.146333
R19121 GNDA.n228 GNDA.n130 0.146333
R19122 GNDA.n238 GNDA.n128 0.146333
R19123 GNDA.n244 GNDA.n128 0.146333
R19124 GNDA.n245 GNDA.n244 0.146333
R19125 GNDA.n255 GNDA.n254 0.146333
R19126 GNDA.n258 GNDA.n255 0.146333
R19127 GNDA.n258 GNDA.n124 0.146333
R19128 GNDA.n5274 GNDA.n327 0.135917
R19129 GNDA.n5168 GNDA.n5165 0.135917
R19130 GNDA.n5174 GNDA.n5157 0.135917
R19131 GNDA.n5184 GNDA.n5155 0.135917
R19132 GNDA.n5188 GNDA.n5185 0.135917
R19133 GNDA.n5198 GNDA.n5195 0.135917
R19134 GNDA.n5204 GNDA.n5151 0.135917
R19135 GNDA.n5214 GNDA.n5149 0.135917
R19136 GNDA.n5218 GNDA.n5215 0.135917
R19137 GNDA.n5228 GNDA.n5225 0.135917
R19138 GNDA.n5234 GNDA.n5145 0.135917
R19139 GNDA.n5244 GNDA.n5143 0.135917
R19140 GNDA.n5248 GNDA.n5245 0.135917
R19141 GNDA.n5258 GNDA.n5255 0.135917
R19142 GNDA.n5264 GNDA.n5139 0.135917
R19143 GNDA.n4961 GNDA.n3457 0.135917
R19144 GNDA.n4855 GNDA.n4852 0.135917
R19145 GNDA.n4861 GNDA.n4844 0.135917
R19146 GNDA.n4871 GNDA.n4842 0.135917
R19147 GNDA.n4875 GNDA.n4872 0.135917
R19148 GNDA.n4885 GNDA.n4882 0.135917
R19149 GNDA.n4891 GNDA.n4838 0.135917
R19150 GNDA.n4901 GNDA.n4836 0.135917
R19151 GNDA.n4905 GNDA.n4902 0.135917
R19152 GNDA.n4915 GNDA.n4912 0.135917
R19153 GNDA.n4921 GNDA.n4832 0.135917
R19154 GNDA.n4931 GNDA.n4830 0.135917
R19155 GNDA.n4935 GNDA.n4932 0.135917
R19156 GNDA.n4945 GNDA.n4942 0.135917
R19157 GNDA.n4951 GNDA.n4826 0.135917
R19158 GNDA.n4685 GNDA.n4683 0.135917
R19159 GNDA.n4695 GNDA.n4692 0.135917
R19160 GNDA.n4701 GNDA.n4679 0.135917
R19161 GNDA.n4711 GNDA.n4677 0.135917
R19162 GNDA.n4715 GNDA.n4712 0.135917
R19163 GNDA.n4725 GNDA.n4722 0.135917
R19164 GNDA.n4731 GNDA.n4673 0.135917
R19165 GNDA.n4741 GNDA.n4671 0.135917
R19166 GNDA.n4745 GNDA.n4742 0.135917
R19167 GNDA.n4755 GNDA.n4752 0.135917
R19168 GNDA.n4761 GNDA.n4667 0.135917
R19169 GNDA.n4771 GNDA.n4665 0.135917
R19170 GNDA.n4775 GNDA.n4772 0.135917
R19171 GNDA.n4785 GNDA.n4782 0.135917
R19172 GNDA.n4791 GNDA.n4661 0.135917
R19173 GNDA.n4519 GNDA.n4517 0.135917
R19174 GNDA.n4529 GNDA.n4526 0.135917
R19175 GNDA.n4535 GNDA.n4513 0.135917
R19176 GNDA.n4545 GNDA.n4511 0.135917
R19177 GNDA.n4549 GNDA.n4546 0.135917
R19178 GNDA.n4559 GNDA.n4556 0.135917
R19179 GNDA.n4565 GNDA.n4507 0.135917
R19180 GNDA.n4575 GNDA.n4505 0.135917
R19181 GNDA.n4579 GNDA.n4576 0.135917
R19182 GNDA.n4589 GNDA.n4586 0.135917
R19183 GNDA.n4595 GNDA.n4501 0.135917
R19184 GNDA.n4605 GNDA.n4499 0.135917
R19185 GNDA.n4609 GNDA.n4606 0.135917
R19186 GNDA.n4619 GNDA.n4616 0.135917
R19187 GNDA.n4625 GNDA.n4495 0.135917
R19188 GNDA.n4353 GNDA.n4351 0.135917
R19189 GNDA.n4363 GNDA.n4360 0.135917
R19190 GNDA.n4369 GNDA.n4347 0.135917
R19191 GNDA.n4379 GNDA.n4345 0.135917
R19192 GNDA.n4383 GNDA.n4380 0.135917
R19193 GNDA.n4393 GNDA.n4390 0.135917
R19194 GNDA.n4399 GNDA.n4341 0.135917
R19195 GNDA.n4409 GNDA.n4339 0.135917
R19196 GNDA.n4413 GNDA.n4410 0.135917
R19197 GNDA.n4423 GNDA.n4420 0.135917
R19198 GNDA.n4429 GNDA.n4335 0.135917
R19199 GNDA.n4439 GNDA.n4333 0.135917
R19200 GNDA.n4443 GNDA.n4440 0.135917
R19201 GNDA.n4453 GNDA.n4450 0.135917
R19202 GNDA.n4459 GNDA.n4329 0.135917
R19203 GNDA.n4187 GNDA.n4185 0.135917
R19204 GNDA.n4197 GNDA.n4194 0.135917
R19205 GNDA.n4203 GNDA.n4181 0.135917
R19206 GNDA.n4213 GNDA.n4179 0.135917
R19207 GNDA.n4217 GNDA.n4214 0.135917
R19208 GNDA.n4227 GNDA.n4224 0.135917
R19209 GNDA.n4233 GNDA.n4175 0.135917
R19210 GNDA.n4243 GNDA.n4173 0.135917
R19211 GNDA.n4247 GNDA.n4244 0.135917
R19212 GNDA.n4257 GNDA.n4254 0.135917
R19213 GNDA.n4263 GNDA.n4169 0.135917
R19214 GNDA.n4273 GNDA.n4167 0.135917
R19215 GNDA.n4277 GNDA.n4274 0.135917
R19216 GNDA.n4287 GNDA.n4284 0.135917
R19217 GNDA.n4293 GNDA.n4163 0.135917
R19218 GNDA.n3689 GNDA.n3687 0.135917
R19219 GNDA.n3699 GNDA.n3696 0.135917
R19220 GNDA.n3705 GNDA.n3505 0.135917
R19221 GNDA.n3715 GNDA.n3503 0.135917
R19222 GNDA.n3719 GNDA.n3716 0.135917
R19223 GNDA.n3729 GNDA.n3726 0.135917
R19224 GNDA.n3735 GNDA.n3499 0.135917
R19225 GNDA.n3745 GNDA.n3497 0.135917
R19226 GNDA.n3749 GNDA.n3746 0.135917
R19227 GNDA.n3759 GNDA.n3756 0.135917
R19228 GNDA.n3765 GNDA.n3493 0.135917
R19229 GNDA.n3775 GNDA.n3491 0.135917
R19230 GNDA.n3779 GNDA.n3776 0.135917
R19231 GNDA.n3789 GNDA.n3786 0.135917
R19232 GNDA.n3795 GNDA.n3487 0.135917
R19233 GNDA.n4021 GNDA.n4019 0.135917
R19234 GNDA.n4031 GNDA.n4028 0.135917
R19235 GNDA.n4037 GNDA.n4015 0.135917
R19236 GNDA.n4047 GNDA.n4013 0.135917
R19237 GNDA.n4051 GNDA.n4048 0.135917
R19238 GNDA.n4061 GNDA.n4058 0.135917
R19239 GNDA.n4067 GNDA.n4009 0.135917
R19240 GNDA.n4077 GNDA.n4007 0.135917
R19241 GNDA.n4081 GNDA.n4078 0.135917
R19242 GNDA.n4091 GNDA.n4088 0.135917
R19243 GNDA.n4097 GNDA.n4003 0.135917
R19244 GNDA.n4107 GNDA.n4001 0.135917
R19245 GNDA.n4111 GNDA.n4108 0.135917
R19246 GNDA.n4121 GNDA.n4118 0.135917
R19247 GNDA.n4127 GNDA.n3997 0.135917
R19248 GNDA.n3855 GNDA.n3853 0.135917
R19249 GNDA.n3865 GNDA.n3862 0.135917
R19250 GNDA.n3871 GNDA.n3849 0.135917
R19251 GNDA.n3881 GNDA.n3847 0.135917
R19252 GNDA.n3885 GNDA.n3882 0.135917
R19253 GNDA.n3895 GNDA.n3892 0.135917
R19254 GNDA.n3901 GNDA.n3843 0.135917
R19255 GNDA.n3911 GNDA.n3841 0.135917
R19256 GNDA.n3915 GNDA.n3912 0.135917
R19257 GNDA.n3925 GNDA.n3922 0.135917
R19258 GNDA.n3931 GNDA.n3837 0.135917
R19259 GNDA.n3941 GNDA.n3835 0.135917
R19260 GNDA.n3945 GNDA.n3942 0.135917
R19261 GNDA.n3955 GNDA.n3952 0.135917
R19262 GNDA.n3961 GNDA.n3831 0.135917
R19263 GNDA.n3674 GNDA.n3512 0.135917
R19264 GNDA.n3516 GNDA.n3515 0.135917
R19265 GNDA.n3518 GNDA.n3517 0.135917
R19266 GNDA.n3522 GNDA.n3521 0.135917
R19267 GNDA.n3524 GNDA.n3523 0.135917
R19268 GNDA.n3528 GNDA.n3527 0.135917
R19269 GNDA.n3530 GNDA.n3529 0.135917
R19270 GNDA.n3534 GNDA.n3533 0.135917
R19271 GNDA.n3536 GNDA.n3535 0.135917
R19272 GNDA.n3540 GNDA.n3539 0.135917
R19273 GNDA.n3542 GNDA.n3541 0.135917
R19274 GNDA.n3546 GNDA.n3545 0.135917
R19275 GNDA.n3548 GNDA.n3547 0.135917
R19276 GNDA.n3552 GNDA.n3551 0.135917
R19277 GNDA.n3554 GNDA.n3553 0.135917
R19278 GNDA.n568 GNDA.n406 0.135917
R19279 GNDA.n410 GNDA.n409 0.135917
R19280 GNDA.n412 GNDA.n411 0.135917
R19281 GNDA.n416 GNDA.n415 0.135917
R19282 GNDA.n418 GNDA.n417 0.135917
R19283 GNDA.n422 GNDA.n421 0.135917
R19284 GNDA.n424 GNDA.n423 0.135917
R19285 GNDA.n428 GNDA.n427 0.135917
R19286 GNDA.n430 GNDA.n429 0.135917
R19287 GNDA.n434 GNDA.n433 0.135917
R19288 GNDA.n436 GNDA.n435 0.135917
R19289 GNDA.n440 GNDA.n439 0.135917
R19290 GNDA.n442 GNDA.n441 0.135917
R19291 GNDA.n446 GNDA.n445 0.135917
R19292 GNDA.n448 GNDA.n447 0.135917
R19293 GNDA.n5021 GNDA.n5019 0.135917
R19294 GNDA.n5031 GNDA.n5028 0.135917
R19295 GNDA.n5037 GNDA.n399 0.135917
R19296 GNDA.n5047 GNDA.n397 0.135917
R19297 GNDA.n5051 GNDA.n5048 0.135917
R19298 GNDA.n5061 GNDA.n5058 0.135917
R19299 GNDA.n5067 GNDA.n393 0.135917
R19300 GNDA.n5077 GNDA.n391 0.135917
R19301 GNDA.n5081 GNDA.n5078 0.135917
R19302 GNDA.n5091 GNDA.n5088 0.135917
R19303 GNDA.n5097 GNDA.n387 0.135917
R19304 GNDA.n5107 GNDA.n385 0.135917
R19305 GNDA.n5111 GNDA.n5108 0.135917
R19306 GNDA.n5121 GNDA.n5118 0.135917
R19307 GNDA.n5127 GNDA.n381 0.135917
R19308 GNDA.n3371 GNDA.n3209 0.135917
R19309 GNDA.n3213 GNDA.n3212 0.135917
R19310 GNDA.n3215 GNDA.n3214 0.135917
R19311 GNDA.n3219 GNDA.n3218 0.135917
R19312 GNDA.n3221 GNDA.n3220 0.135917
R19313 GNDA.n3225 GNDA.n3224 0.135917
R19314 GNDA.n3227 GNDA.n3226 0.135917
R19315 GNDA.n3231 GNDA.n3230 0.135917
R19316 GNDA.n3233 GNDA.n3232 0.135917
R19317 GNDA.n3237 GNDA.n3236 0.135917
R19318 GNDA.n3239 GNDA.n3238 0.135917
R19319 GNDA.n3243 GNDA.n3242 0.135917
R19320 GNDA.n3245 GNDA.n3244 0.135917
R19321 GNDA.n3249 GNDA.n3248 0.135917
R19322 GNDA.n3251 GNDA.n3250 0.135917
R19323 GNDA.n3199 GNDA.n597 0.135917
R19324 GNDA.n3093 GNDA.n3090 0.135917
R19325 GNDA.n3099 GNDA.n3082 0.135917
R19326 GNDA.n3109 GNDA.n3080 0.135917
R19327 GNDA.n3113 GNDA.n3110 0.135917
R19328 GNDA.n3123 GNDA.n3120 0.135917
R19329 GNDA.n3129 GNDA.n3076 0.135917
R19330 GNDA.n3139 GNDA.n3074 0.135917
R19331 GNDA.n3143 GNDA.n3140 0.135917
R19332 GNDA.n3153 GNDA.n3150 0.135917
R19333 GNDA.n3159 GNDA.n3070 0.135917
R19334 GNDA.n3169 GNDA.n3068 0.135917
R19335 GNDA.n3173 GNDA.n3170 0.135917
R19336 GNDA.n3183 GNDA.n3180 0.135917
R19337 GNDA.n3189 GNDA.n3064 0.135917
R19338 GNDA.n2923 GNDA.n2921 0.135917
R19339 GNDA.n2933 GNDA.n2930 0.135917
R19340 GNDA.n2939 GNDA.n2909 0.135917
R19341 GNDA.n2949 GNDA.n2907 0.135917
R19342 GNDA.n2953 GNDA.n2950 0.135917
R19343 GNDA.n2963 GNDA.n2960 0.135917
R19344 GNDA.n2969 GNDA.n2903 0.135917
R19345 GNDA.n2979 GNDA.n2901 0.135917
R19346 GNDA.n2983 GNDA.n2980 0.135917
R19347 GNDA.n2993 GNDA.n2990 0.135917
R19348 GNDA.n2999 GNDA.n2897 0.135917
R19349 GNDA.n3009 GNDA.n2895 0.135917
R19350 GNDA.n3013 GNDA.n3010 0.135917
R19351 GNDA.n3023 GNDA.n3020 0.135917
R19352 GNDA.n3029 GNDA.n2891 0.135917
R19353 GNDA.n2287 GNDA.n2285 0.135917
R19354 GNDA.n2297 GNDA.n2294 0.135917
R19355 GNDA.n2303 GNDA.n711 0.135917
R19356 GNDA.n2313 GNDA.n709 0.135917
R19357 GNDA.n2317 GNDA.n2314 0.135917
R19358 GNDA.n2327 GNDA.n2324 0.135917
R19359 GNDA.n2333 GNDA.n705 0.135917
R19360 GNDA.n2343 GNDA.n703 0.135917
R19361 GNDA.n2347 GNDA.n2344 0.135917
R19362 GNDA.n2357 GNDA.n2354 0.135917
R19363 GNDA.n2363 GNDA.n699 0.135917
R19364 GNDA.n2373 GNDA.n697 0.135917
R19365 GNDA.n2377 GNDA.n2374 0.135917
R19366 GNDA.n2387 GNDA.n2384 0.135917
R19367 GNDA.n2393 GNDA.n693 0.135917
R19368 GNDA.n2749 GNDA.n2747 0.135917
R19369 GNDA.n2759 GNDA.n2756 0.135917
R19370 GNDA.n2765 GNDA.n645 0.135917
R19371 GNDA.n2775 GNDA.n643 0.135917
R19372 GNDA.n2779 GNDA.n2776 0.135917
R19373 GNDA.n2789 GNDA.n2786 0.135917
R19374 GNDA.n2795 GNDA.n639 0.135917
R19375 GNDA.n2805 GNDA.n637 0.135917
R19376 GNDA.n2809 GNDA.n2806 0.135917
R19377 GNDA.n2819 GNDA.n2816 0.135917
R19378 GNDA.n2825 GNDA.n633 0.135917
R19379 GNDA.n2835 GNDA.n631 0.135917
R19380 GNDA.n2839 GNDA.n2836 0.135917
R19381 GNDA.n2849 GNDA.n2846 0.135917
R19382 GNDA.n2855 GNDA.n627 0.135917
R19383 GNDA.n2734 GNDA.n2572 0.135917
R19384 GNDA.n2576 GNDA.n2575 0.135917
R19385 GNDA.n2578 GNDA.n2577 0.135917
R19386 GNDA.n2582 GNDA.n2581 0.135917
R19387 GNDA.n2584 GNDA.n2583 0.135917
R19388 GNDA.n2588 GNDA.n2587 0.135917
R19389 GNDA.n2590 GNDA.n2589 0.135917
R19390 GNDA.n2594 GNDA.n2593 0.135917
R19391 GNDA.n2596 GNDA.n2595 0.135917
R19392 GNDA.n2600 GNDA.n2599 0.135917
R19393 GNDA.n2602 GNDA.n2601 0.135917
R19394 GNDA.n2606 GNDA.n2605 0.135917
R19395 GNDA.n2608 GNDA.n2607 0.135917
R19396 GNDA.n2612 GNDA.n2611 0.135917
R19397 GNDA.n2614 GNDA.n2613 0.135917
R19398 GNDA.n2563 GNDA.n663 0.135917
R19399 GNDA.n2457 GNDA.n2454 0.135917
R19400 GNDA.n2463 GNDA.n2446 0.135917
R19401 GNDA.n2473 GNDA.n2444 0.135917
R19402 GNDA.n2477 GNDA.n2474 0.135917
R19403 GNDA.n2487 GNDA.n2484 0.135917
R19404 GNDA.n2493 GNDA.n2440 0.135917
R19405 GNDA.n2503 GNDA.n2438 0.135917
R19406 GNDA.n2507 GNDA.n2504 0.135917
R19407 GNDA.n2517 GNDA.n2514 0.135917
R19408 GNDA.n2523 GNDA.n2434 0.135917
R19409 GNDA.n2533 GNDA.n2432 0.135917
R19410 GNDA.n2537 GNDA.n2534 0.135917
R19411 GNDA.n2547 GNDA.n2544 0.135917
R19412 GNDA.n2553 GNDA.n2428 0.135917
R19413 GNDA.n2274 GNDA.n2112 0.135917
R19414 GNDA.n2116 GNDA.n2115 0.135917
R19415 GNDA.n2118 GNDA.n2117 0.135917
R19416 GNDA.n2122 GNDA.n2121 0.135917
R19417 GNDA.n2124 GNDA.n2123 0.135917
R19418 GNDA.n2128 GNDA.n2127 0.135917
R19419 GNDA.n2130 GNDA.n2129 0.135917
R19420 GNDA.n2134 GNDA.n2133 0.135917
R19421 GNDA.n2136 GNDA.n2135 0.135917
R19422 GNDA.n2140 GNDA.n2139 0.135917
R19423 GNDA.n2142 GNDA.n2141 0.135917
R19424 GNDA.n2146 GNDA.n2145 0.135917
R19425 GNDA.n2148 GNDA.n2147 0.135917
R19426 GNDA.n2152 GNDA.n2151 0.135917
R19427 GNDA.n2154 GNDA.n2153 0.135917
R19428 GNDA.n2100 GNDA.n726 0.135917
R19429 GNDA.n1994 GNDA.n1991 0.135917
R19430 GNDA.n2000 GNDA.n1983 0.135917
R19431 GNDA.n2010 GNDA.n1981 0.135917
R19432 GNDA.n2014 GNDA.n2011 0.135917
R19433 GNDA.n2024 GNDA.n2021 0.135917
R19434 GNDA.n2030 GNDA.n1977 0.135917
R19435 GNDA.n2040 GNDA.n1975 0.135917
R19436 GNDA.n2044 GNDA.n2041 0.135917
R19437 GNDA.n2054 GNDA.n2051 0.135917
R19438 GNDA.n2060 GNDA.n1971 0.135917
R19439 GNDA.n2070 GNDA.n1969 0.135917
R19440 GNDA.n2074 GNDA.n2071 0.135917
R19441 GNDA.n2084 GNDA.n2081 0.135917
R19442 GNDA.n2090 GNDA.n1965 0.135917
R19443 GNDA.n1824 GNDA.n1822 0.135917
R19444 GNDA.n1834 GNDA.n1831 0.135917
R19445 GNDA.n1840 GNDA.n774 0.135917
R19446 GNDA.n1850 GNDA.n772 0.135917
R19447 GNDA.n1854 GNDA.n1851 0.135917
R19448 GNDA.n1864 GNDA.n1861 0.135917
R19449 GNDA.n1870 GNDA.n768 0.135917
R19450 GNDA.n1880 GNDA.n766 0.135917
R19451 GNDA.n1884 GNDA.n1881 0.135917
R19452 GNDA.n1894 GNDA.n1891 0.135917
R19453 GNDA.n1900 GNDA.n762 0.135917
R19454 GNDA.n1910 GNDA.n760 0.135917
R19455 GNDA.n1914 GNDA.n1911 0.135917
R19456 GNDA.n1924 GNDA.n1921 0.135917
R19457 GNDA.n1930 GNDA.n756 0.135917
R19458 GNDA.n1687 GNDA.n1525 0.135917
R19459 GNDA.n1529 GNDA.n1528 0.135917
R19460 GNDA.n1531 GNDA.n1530 0.135917
R19461 GNDA.n1535 GNDA.n1534 0.135917
R19462 GNDA.n1537 GNDA.n1536 0.135917
R19463 GNDA.n1541 GNDA.n1540 0.135917
R19464 GNDA.n1543 GNDA.n1542 0.135917
R19465 GNDA.n1547 GNDA.n1546 0.135917
R19466 GNDA.n1549 GNDA.n1548 0.135917
R19467 GNDA.n1553 GNDA.n1552 0.135917
R19468 GNDA.n1555 GNDA.n1554 0.135917
R19469 GNDA.n1559 GNDA.n1558 0.135917
R19470 GNDA.n1561 GNDA.n1560 0.135917
R19471 GNDA.n1565 GNDA.n1564 0.135917
R19472 GNDA.n1567 GNDA.n1566 0.135917
R19473 GNDA.n1516 GNDA.n792 0.135917
R19474 GNDA.n1410 GNDA.n1407 0.135917
R19475 GNDA.n1416 GNDA.n1399 0.135917
R19476 GNDA.n1426 GNDA.n1397 0.135917
R19477 GNDA.n1430 GNDA.n1427 0.135917
R19478 GNDA.n1440 GNDA.n1437 0.135917
R19479 GNDA.n1446 GNDA.n1393 0.135917
R19480 GNDA.n1456 GNDA.n1391 0.135917
R19481 GNDA.n1460 GNDA.n1457 0.135917
R19482 GNDA.n1470 GNDA.n1467 0.135917
R19483 GNDA.n1476 GNDA.n1387 0.135917
R19484 GNDA.n1486 GNDA.n1385 0.135917
R19485 GNDA.n1490 GNDA.n1487 0.135917
R19486 GNDA.n1500 GNDA.n1497 0.135917
R19487 GNDA.n1506 GNDA.n1381 0.135917
R19488 GNDA.n1241 GNDA.n1215 0.135917
R19489 GNDA.n1251 GNDA.n1213 0.135917
R19490 GNDA.n1257 GNDA.n1254 0.135917
R19491 GNDA.n1267 GNDA.n1264 0.135917
R19492 GNDA.n1271 GNDA.n1209 0.135917
R19493 GNDA.n1281 GNDA.n1207 0.135917
R19494 GNDA.n1287 GNDA.n1284 0.135917
R19495 GNDA.n1297 GNDA.n1294 0.135917
R19496 GNDA.n1301 GNDA.n1203 0.135917
R19497 GNDA.n1311 GNDA.n1201 0.135917
R19498 GNDA.n1317 GNDA.n1314 0.135917
R19499 GNDA.n1327 GNDA.n1324 0.135917
R19500 GNDA.n1331 GNDA.n1197 0.135917
R19501 GNDA.n1341 GNDA.n1195 0.135917
R19502 GNDA.n1346 GNDA.n1344 0.135917
R19503 GNDA.n7142 GNDA.n7128 0.135917
R19504 GNDA.n7146 GNDA.n7143 0.135917
R19505 GNDA.n7154 GNDA.n7151 0.135917
R19506 GNDA.n7158 GNDA.n7120 0.135917
R19507 GNDA.n7166 GNDA.n7116 0.135917
R19508 GNDA.n7170 GNDA.n7167 0.135917
R19509 GNDA.n7178 GNDA.n7175 0.135917
R19510 GNDA.n7182 GNDA.n7108 0.135917
R19511 GNDA.n7190 GNDA.n7104 0.135917
R19512 GNDA.n7194 GNDA.n7191 0.135917
R19513 GNDA.n7202 GNDA.n7199 0.135917
R19514 GNDA.n7206 GNDA.n7096 0.135917
R19515 GNDA.n7214 GNDA.n7092 0.135917
R19516 GNDA.n7218 GNDA.n7215 0.135917
R19517 GNDA.n7227 GNDA.n96 0.135917
R19518 GNDA.n159 GNDA.n145 0.135917
R19519 GNDA.n161 GNDA.n160 0.135917
R19520 GNDA.n171 GNDA.n170 0.135917
R19521 GNDA.n179 GNDA.n141 0.135917
R19522 GNDA.n189 GNDA.n139 0.135917
R19523 GNDA.n191 GNDA.n190 0.135917
R19524 GNDA.n201 GNDA.n200 0.135917
R19525 GNDA.n209 GNDA.n135 0.135917
R19526 GNDA.n219 GNDA.n133 0.135917
R19527 GNDA.n221 GNDA.n220 0.135917
R19528 GNDA.n231 GNDA.n230 0.135917
R19529 GNDA.n239 GNDA.n129 0.135917
R19530 GNDA.n249 GNDA.n127 0.135917
R19531 GNDA.n251 GNDA.n250 0.135917
R19532 GNDA.n7062 GNDA.n260 0.135917
R19533 GNDA.n158 GNDA.n155 0.135917
R19534 GNDA.n164 GNDA.n144 0.135917
R19535 GNDA.n174 GNDA.n142 0.135917
R19536 GNDA.n178 GNDA.n175 0.135917
R19537 GNDA.n188 GNDA.n185 0.135917
R19538 GNDA.n194 GNDA.n138 0.135917
R19539 GNDA.n204 GNDA.n136 0.135917
R19540 GNDA.n208 GNDA.n205 0.135917
R19541 GNDA.n218 GNDA.n215 0.135917
R19542 GNDA.n224 GNDA.n132 0.135917
R19543 GNDA.n234 GNDA.n130 0.135917
R19544 GNDA.n238 GNDA.n235 0.135917
R19545 GNDA.n248 GNDA.n245 0.135917
R19546 GNDA.n254 GNDA.n126 0.135917
R19547 GNDA.n7063 GNDA.n124 0.135917
R19548 GNDA.n5168 GNDA.n5157 0.1255
R19549 GNDA.n5185 GNDA.n5184 0.1255
R19550 GNDA.n5198 GNDA.n5151 0.1255
R19551 GNDA.n5215 GNDA.n5214 0.1255
R19552 GNDA.n5228 GNDA.n5145 0.1255
R19553 GNDA.n5245 GNDA.n5244 0.1255
R19554 GNDA.n5258 GNDA.n5139 0.1255
R19555 GNDA.n4855 GNDA.n4844 0.1255
R19556 GNDA.n4872 GNDA.n4871 0.1255
R19557 GNDA.n4885 GNDA.n4838 0.1255
R19558 GNDA.n4902 GNDA.n4901 0.1255
R19559 GNDA.n4915 GNDA.n4832 0.1255
R19560 GNDA.n4932 GNDA.n4931 0.1255
R19561 GNDA.n4945 GNDA.n4826 0.1255
R19562 GNDA.n4695 GNDA.n4679 0.1255
R19563 GNDA.n4712 GNDA.n4711 0.1255
R19564 GNDA.n4725 GNDA.n4673 0.1255
R19565 GNDA.n4742 GNDA.n4741 0.1255
R19566 GNDA.n4755 GNDA.n4667 0.1255
R19567 GNDA.n4772 GNDA.n4771 0.1255
R19568 GNDA.n4785 GNDA.n4661 0.1255
R19569 GNDA.n4529 GNDA.n4513 0.1255
R19570 GNDA.n4546 GNDA.n4545 0.1255
R19571 GNDA.n4559 GNDA.n4507 0.1255
R19572 GNDA.n4576 GNDA.n4575 0.1255
R19573 GNDA.n4589 GNDA.n4501 0.1255
R19574 GNDA.n4606 GNDA.n4605 0.1255
R19575 GNDA.n4619 GNDA.n4495 0.1255
R19576 GNDA.n4363 GNDA.n4347 0.1255
R19577 GNDA.n4380 GNDA.n4379 0.1255
R19578 GNDA.n4393 GNDA.n4341 0.1255
R19579 GNDA.n4410 GNDA.n4409 0.1255
R19580 GNDA.n4423 GNDA.n4335 0.1255
R19581 GNDA.n4440 GNDA.n4439 0.1255
R19582 GNDA.n4453 GNDA.n4329 0.1255
R19583 GNDA.n4197 GNDA.n4181 0.1255
R19584 GNDA.n4214 GNDA.n4213 0.1255
R19585 GNDA.n4227 GNDA.n4175 0.1255
R19586 GNDA.n4244 GNDA.n4243 0.1255
R19587 GNDA.n4257 GNDA.n4169 0.1255
R19588 GNDA.n4274 GNDA.n4273 0.1255
R19589 GNDA.n4287 GNDA.n4163 0.1255
R19590 GNDA.n3699 GNDA.n3505 0.1255
R19591 GNDA.n3716 GNDA.n3715 0.1255
R19592 GNDA.n3729 GNDA.n3499 0.1255
R19593 GNDA.n3746 GNDA.n3745 0.1255
R19594 GNDA.n3759 GNDA.n3493 0.1255
R19595 GNDA.n3776 GNDA.n3775 0.1255
R19596 GNDA.n3789 GNDA.n3487 0.1255
R19597 GNDA.n4031 GNDA.n4015 0.1255
R19598 GNDA.n4048 GNDA.n4047 0.1255
R19599 GNDA.n4061 GNDA.n4009 0.1255
R19600 GNDA.n4078 GNDA.n4077 0.1255
R19601 GNDA.n4091 GNDA.n4003 0.1255
R19602 GNDA.n4108 GNDA.n4107 0.1255
R19603 GNDA.n4121 GNDA.n3997 0.1255
R19604 GNDA.n3865 GNDA.n3849 0.1255
R19605 GNDA.n3882 GNDA.n3881 0.1255
R19606 GNDA.n3895 GNDA.n3843 0.1255
R19607 GNDA.n3912 GNDA.n3911 0.1255
R19608 GNDA.n3925 GNDA.n3837 0.1255
R19609 GNDA.n3942 GNDA.n3941 0.1255
R19610 GNDA.n3955 GNDA.n3831 0.1255
R19611 GNDA.n3517 GNDA.n3516 0.1255
R19612 GNDA.n3523 GNDA.n3522 0.1255
R19613 GNDA.n3529 GNDA.n3528 0.1255
R19614 GNDA.n3535 GNDA.n3534 0.1255
R19615 GNDA.n3541 GNDA.n3540 0.1255
R19616 GNDA.n3547 GNDA.n3546 0.1255
R19617 GNDA.n3553 GNDA.n3552 0.1255
R19618 GNDA.n411 GNDA.n410 0.1255
R19619 GNDA.n417 GNDA.n416 0.1255
R19620 GNDA.n423 GNDA.n422 0.1255
R19621 GNDA.n429 GNDA.n428 0.1255
R19622 GNDA.n435 GNDA.n434 0.1255
R19623 GNDA.n441 GNDA.n440 0.1255
R19624 GNDA.n447 GNDA.n446 0.1255
R19625 GNDA.n5031 GNDA.n399 0.1255
R19626 GNDA.n5048 GNDA.n5047 0.1255
R19627 GNDA.n5061 GNDA.n393 0.1255
R19628 GNDA.n5078 GNDA.n5077 0.1255
R19629 GNDA.n5091 GNDA.n387 0.1255
R19630 GNDA.n5108 GNDA.n5107 0.1255
R19631 GNDA.n5121 GNDA.n381 0.1255
R19632 GNDA.n3214 GNDA.n3213 0.1255
R19633 GNDA.n3220 GNDA.n3219 0.1255
R19634 GNDA.n3226 GNDA.n3225 0.1255
R19635 GNDA.n3232 GNDA.n3231 0.1255
R19636 GNDA.n3238 GNDA.n3237 0.1255
R19637 GNDA.n3244 GNDA.n3243 0.1255
R19638 GNDA.n3250 GNDA.n3249 0.1255
R19639 GNDA.n3093 GNDA.n3082 0.1255
R19640 GNDA.n3110 GNDA.n3109 0.1255
R19641 GNDA.n3123 GNDA.n3076 0.1255
R19642 GNDA.n3140 GNDA.n3139 0.1255
R19643 GNDA.n3153 GNDA.n3070 0.1255
R19644 GNDA.n3170 GNDA.n3169 0.1255
R19645 GNDA.n3183 GNDA.n3064 0.1255
R19646 GNDA.n2933 GNDA.n2909 0.1255
R19647 GNDA.n2950 GNDA.n2949 0.1255
R19648 GNDA.n2963 GNDA.n2903 0.1255
R19649 GNDA.n2980 GNDA.n2979 0.1255
R19650 GNDA.n2993 GNDA.n2897 0.1255
R19651 GNDA.n3010 GNDA.n3009 0.1255
R19652 GNDA.n3023 GNDA.n2891 0.1255
R19653 GNDA.n2297 GNDA.n711 0.1255
R19654 GNDA.n2314 GNDA.n2313 0.1255
R19655 GNDA.n2327 GNDA.n705 0.1255
R19656 GNDA.n2344 GNDA.n2343 0.1255
R19657 GNDA.n2357 GNDA.n699 0.1255
R19658 GNDA.n2374 GNDA.n2373 0.1255
R19659 GNDA.n2387 GNDA.n693 0.1255
R19660 GNDA.n2759 GNDA.n645 0.1255
R19661 GNDA.n2776 GNDA.n2775 0.1255
R19662 GNDA.n2789 GNDA.n639 0.1255
R19663 GNDA.n2806 GNDA.n2805 0.1255
R19664 GNDA.n2819 GNDA.n633 0.1255
R19665 GNDA.n2836 GNDA.n2835 0.1255
R19666 GNDA.n2849 GNDA.n627 0.1255
R19667 GNDA.n2577 GNDA.n2576 0.1255
R19668 GNDA.n2583 GNDA.n2582 0.1255
R19669 GNDA.n2589 GNDA.n2588 0.1255
R19670 GNDA.n2595 GNDA.n2594 0.1255
R19671 GNDA.n2601 GNDA.n2600 0.1255
R19672 GNDA.n2607 GNDA.n2606 0.1255
R19673 GNDA.n2613 GNDA.n2612 0.1255
R19674 GNDA.n2457 GNDA.n2446 0.1255
R19675 GNDA.n2474 GNDA.n2473 0.1255
R19676 GNDA.n2487 GNDA.n2440 0.1255
R19677 GNDA.n2504 GNDA.n2503 0.1255
R19678 GNDA.n2517 GNDA.n2434 0.1255
R19679 GNDA.n2534 GNDA.n2533 0.1255
R19680 GNDA.n2547 GNDA.n2428 0.1255
R19681 GNDA.n2117 GNDA.n2116 0.1255
R19682 GNDA.n2123 GNDA.n2122 0.1255
R19683 GNDA.n2129 GNDA.n2128 0.1255
R19684 GNDA.n2135 GNDA.n2134 0.1255
R19685 GNDA.n2141 GNDA.n2140 0.1255
R19686 GNDA.n2147 GNDA.n2146 0.1255
R19687 GNDA.n2153 GNDA.n2152 0.1255
R19688 GNDA.n1994 GNDA.n1983 0.1255
R19689 GNDA.n2011 GNDA.n2010 0.1255
R19690 GNDA.n2024 GNDA.n1977 0.1255
R19691 GNDA.n2041 GNDA.n2040 0.1255
R19692 GNDA.n2054 GNDA.n1971 0.1255
R19693 GNDA.n2071 GNDA.n2070 0.1255
R19694 GNDA.n2084 GNDA.n1965 0.1255
R19695 GNDA.n1834 GNDA.n774 0.1255
R19696 GNDA.n1851 GNDA.n1850 0.1255
R19697 GNDA.n1864 GNDA.n768 0.1255
R19698 GNDA.n1881 GNDA.n1880 0.1255
R19699 GNDA.n1894 GNDA.n762 0.1255
R19700 GNDA.n1911 GNDA.n1910 0.1255
R19701 GNDA.n1924 GNDA.n756 0.1255
R19702 GNDA.n1530 GNDA.n1529 0.1255
R19703 GNDA.n1536 GNDA.n1535 0.1255
R19704 GNDA.n1542 GNDA.n1541 0.1255
R19705 GNDA.n1548 GNDA.n1547 0.1255
R19706 GNDA.n1554 GNDA.n1553 0.1255
R19707 GNDA.n1560 GNDA.n1559 0.1255
R19708 GNDA.n1566 GNDA.n1565 0.1255
R19709 GNDA.n1410 GNDA.n1399 0.1255
R19710 GNDA.n1427 GNDA.n1426 0.1255
R19711 GNDA.n1440 GNDA.n1393 0.1255
R19712 GNDA.n1457 GNDA.n1456 0.1255
R19713 GNDA.n1470 GNDA.n1387 0.1255
R19714 GNDA.n1487 GNDA.n1486 0.1255
R19715 GNDA.n1500 GNDA.n1381 0.1255
R19716 GNDA.n1254 GNDA.n1251 0.1255
R19717 GNDA.n1267 GNDA.n1209 0.1255
R19718 GNDA.n1284 GNDA.n1281 0.1255
R19719 GNDA.n1297 GNDA.n1203 0.1255
R19720 GNDA.n1314 GNDA.n1311 0.1255
R19721 GNDA.n1327 GNDA.n1197 0.1255
R19722 GNDA.n1344 GNDA.n1341 0.1255
R19723 GNDA.n1817 GNDA.n1815 0.1255
R19724 GNDA.n4990 GNDA.n4989 0.1255
R19725 GNDA.n6942 GNDA.n5359 0.1255
R19726 GNDA.n6951 GNDA.n6950 0.1255
R19727 GNDA.n7143 GNDA.n7142 0.1255
R19728 GNDA.n7154 GNDA.n7120 0.1255
R19729 GNDA.n7167 GNDA.n7166 0.1255
R19730 GNDA.n7178 GNDA.n7108 0.1255
R19731 GNDA.n7191 GNDA.n7190 0.1255
R19732 GNDA.n7202 GNDA.n7096 0.1255
R19733 GNDA.n7215 GNDA.n7214 0.1255
R19734 GNDA.n160 GNDA.n159 0.1255
R19735 GNDA.n171 GNDA.n141 0.1255
R19736 GNDA.n190 GNDA.n189 0.1255
R19737 GNDA.n201 GNDA.n135 0.1255
R19738 GNDA.n220 GNDA.n219 0.1255
R19739 GNDA.n231 GNDA.n129 0.1255
R19740 GNDA.n250 GNDA.n249 0.1255
R19741 GNDA.n158 GNDA.n144 0.1255
R19742 GNDA.n175 GNDA.n174 0.1255
R19743 GNDA.n188 GNDA.n138 0.1255
R19744 GNDA.n205 GNDA.n204 0.1255
R19745 GNDA.n218 GNDA.n132 0.1255
R19746 GNDA.n235 GNDA.n234 0.1255
R19747 GNDA.n248 GNDA.n126 0.1255
R19748 GNDA.n1053 GNDA.n1038 0.120864
R19749 GNDA.n1059 GNDA.n1058 0.115944
R19750 GNDA.n3412 GNDA.n3410 0.115083
R19751 GNDA.n3414 GNDA.n3412 0.115083
R19752 GNDA.n3416 GNDA.n3414 0.115083
R19753 GNDA.n3418 GNDA.n3416 0.115083
R19754 GNDA.n1775 GNDA.n1774 0.115083
R19755 GNDA.n1774 GNDA.n1772 0.115083
R19756 GNDA.n1798 GNDA.n1796 0.115083
R19757 GNDA.n1796 GNDA.n1794 0.115083
R19758 GNDA.n1794 GNDA.n1792 0.115083
R19759 GNDA.n1792 GNDA.n1790 0.115083
R19760 GNDA.n1790 GNDA.n1788 0.115083
R19761 GNDA.n7051 GNDA.n7050 0.115083
R19762 GNDA.n7050 GNDA.n7049 0.115083
R19763 GNDA.n7047 GNDA.n7046 0.115083
R19764 GNDA.n7046 GNDA.n7045 0.115083
R19765 GNDA.n7045 GNDA.n7044 0.115083
R19766 GNDA.n7044 GNDA.n7043 0.115083
R19767 GNDA.n7042 GNDA.n7041 0.115083
R19768 GNDA.n7041 GNDA.n7040 0.115083
R19769 GNDA.n7040 GNDA.n7039 0.115083
R19770 GNDA.n7038 GNDA.n7037 0.115083
R19771 GNDA.n7037 GNDA.n7036 0.115083
R19772 GNDA.n7036 GNDA.n7035 0.115083
R19773 GNDA.n2282 GNDA.n660 0.105167
R19774 GNDA.n5005 GNDA.n573 0.105167
R19775 GNDA.n2278 GNDA.n2109 0.09425
R19776 GNDA.n4998 GNDA.n576 0.09425
R19777 GNDA.n7065 GNDA.n98 0.0925906
R19778 GNDA.n3380 GNDA.n3205 0.0838333
R19779 GNDA.n5160 GNDA.n326 0.0734167
R19780 GNDA.n5161 GNDA.n5160 0.0734167
R19781 GNDA.n5161 GNDA.n5158 0.0734167
R19782 GNDA.n5171 GNDA.n5156 0.0734167
R19783 GNDA.n5179 GNDA.n5156 0.0734167
R19784 GNDA.n5180 GNDA.n5179 0.0734167
R19785 GNDA.n5190 GNDA.n5189 0.0734167
R19786 GNDA.n5191 GNDA.n5190 0.0734167
R19787 GNDA.n5191 GNDA.n5152 0.0734167
R19788 GNDA.n5201 GNDA.n5150 0.0734167
R19789 GNDA.n5209 GNDA.n5150 0.0734167
R19790 GNDA.n5210 GNDA.n5209 0.0734167
R19791 GNDA.n5220 GNDA.n5219 0.0734167
R19792 GNDA.n5221 GNDA.n5220 0.0734167
R19793 GNDA.n5221 GNDA.n5146 0.0734167
R19794 GNDA.n5231 GNDA.n5144 0.0734167
R19795 GNDA.n5239 GNDA.n5144 0.0734167
R19796 GNDA.n5240 GNDA.n5239 0.0734167
R19797 GNDA.n5250 GNDA.n5249 0.0734167
R19798 GNDA.n5251 GNDA.n5250 0.0734167
R19799 GNDA.n5251 GNDA.n5140 0.0734167
R19800 GNDA.n5261 GNDA.n5138 0.0734167
R19801 GNDA.n5269 GNDA.n5138 0.0734167
R19802 GNDA.n4847 GNDA.n3456 0.0734167
R19803 GNDA.n4848 GNDA.n4847 0.0734167
R19804 GNDA.n4848 GNDA.n4845 0.0734167
R19805 GNDA.n4858 GNDA.n4843 0.0734167
R19806 GNDA.n4866 GNDA.n4843 0.0734167
R19807 GNDA.n4867 GNDA.n4866 0.0734167
R19808 GNDA.n4877 GNDA.n4876 0.0734167
R19809 GNDA.n4878 GNDA.n4877 0.0734167
R19810 GNDA.n4878 GNDA.n4839 0.0734167
R19811 GNDA.n4888 GNDA.n4837 0.0734167
R19812 GNDA.n4896 GNDA.n4837 0.0734167
R19813 GNDA.n4897 GNDA.n4896 0.0734167
R19814 GNDA.n4907 GNDA.n4906 0.0734167
R19815 GNDA.n4908 GNDA.n4907 0.0734167
R19816 GNDA.n4908 GNDA.n4833 0.0734167
R19817 GNDA.n4918 GNDA.n4831 0.0734167
R19818 GNDA.n4926 GNDA.n4831 0.0734167
R19819 GNDA.n4927 GNDA.n4926 0.0734167
R19820 GNDA.n4937 GNDA.n4936 0.0734167
R19821 GNDA.n4938 GNDA.n4937 0.0734167
R19822 GNDA.n4938 GNDA.n4827 0.0734167
R19823 GNDA.n4948 GNDA.n4825 0.0734167
R19824 GNDA.n4956 GNDA.n4825 0.0734167
R19825 GNDA.n4687 GNDA.n4686 0.0734167
R19826 GNDA.n4688 GNDA.n4687 0.0734167
R19827 GNDA.n4688 GNDA.n4680 0.0734167
R19828 GNDA.n4698 GNDA.n4678 0.0734167
R19829 GNDA.n4706 GNDA.n4678 0.0734167
R19830 GNDA.n4707 GNDA.n4706 0.0734167
R19831 GNDA.n4717 GNDA.n4716 0.0734167
R19832 GNDA.n4718 GNDA.n4717 0.0734167
R19833 GNDA.n4718 GNDA.n4674 0.0734167
R19834 GNDA.n4728 GNDA.n4672 0.0734167
R19835 GNDA.n4736 GNDA.n4672 0.0734167
R19836 GNDA.n4737 GNDA.n4736 0.0734167
R19837 GNDA.n4747 GNDA.n4746 0.0734167
R19838 GNDA.n4748 GNDA.n4747 0.0734167
R19839 GNDA.n4748 GNDA.n4668 0.0734167
R19840 GNDA.n4758 GNDA.n4666 0.0734167
R19841 GNDA.n4766 GNDA.n4666 0.0734167
R19842 GNDA.n4767 GNDA.n4766 0.0734167
R19843 GNDA.n4777 GNDA.n4776 0.0734167
R19844 GNDA.n4778 GNDA.n4777 0.0734167
R19845 GNDA.n4778 GNDA.n4662 0.0734167
R19846 GNDA.n4788 GNDA.n4660 0.0734167
R19847 GNDA.n4796 GNDA.n4660 0.0734167
R19848 GNDA.n4521 GNDA.n4520 0.0734167
R19849 GNDA.n4522 GNDA.n4521 0.0734167
R19850 GNDA.n4522 GNDA.n4514 0.0734167
R19851 GNDA.n4532 GNDA.n4512 0.0734167
R19852 GNDA.n4540 GNDA.n4512 0.0734167
R19853 GNDA.n4541 GNDA.n4540 0.0734167
R19854 GNDA.n4551 GNDA.n4550 0.0734167
R19855 GNDA.n4552 GNDA.n4551 0.0734167
R19856 GNDA.n4552 GNDA.n4508 0.0734167
R19857 GNDA.n4562 GNDA.n4506 0.0734167
R19858 GNDA.n4570 GNDA.n4506 0.0734167
R19859 GNDA.n4571 GNDA.n4570 0.0734167
R19860 GNDA.n4581 GNDA.n4580 0.0734167
R19861 GNDA.n4582 GNDA.n4581 0.0734167
R19862 GNDA.n4582 GNDA.n4502 0.0734167
R19863 GNDA.n4592 GNDA.n4500 0.0734167
R19864 GNDA.n4600 GNDA.n4500 0.0734167
R19865 GNDA.n4601 GNDA.n4600 0.0734167
R19866 GNDA.n4611 GNDA.n4610 0.0734167
R19867 GNDA.n4612 GNDA.n4611 0.0734167
R19868 GNDA.n4612 GNDA.n4496 0.0734167
R19869 GNDA.n4622 GNDA.n4494 0.0734167
R19870 GNDA.n4630 GNDA.n4494 0.0734167
R19871 GNDA.n4355 GNDA.n4354 0.0734167
R19872 GNDA.n4356 GNDA.n4355 0.0734167
R19873 GNDA.n4356 GNDA.n4348 0.0734167
R19874 GNDA.n4366 GNDA.n4346 0.0734167
R19875 GNDA.n4374 GNDA.n4346 0.0734167
R19876 GNDA.n4375 GNDA.n4374 0.0734167
R19877 GNDA.n4385 GNDA.n4384 0.0734167
R19878 GNDA.n4386 GNDA.n4385 0.0734167
R19879 GNDA.n4386 GNDA.n4342 0.0734167
R19880 GNDA.n4396 GNDA.n4340 0.0734167
R19881 GNDA.n4404 GNDA.n4340 0.0734167
R19882 GNDA.n4405 GNDA.n4404 0.0734167
R19883 GNDA.n4415 GNDA.n4414 0.0734167
R19884 GNDA.n4416 GNDA.n4415 0.0734167
R19885 GNDA.n4416 GNDA.n4336 0.0734167
R19886 GNDA.n4426 GNDA.n4334 0.0734167
R19887 GNDA.n4434 GNDA.n4334 0.0734167
R19888 GNDA.n4435 GNDA.n4434 0.0734167
R19889 GNDA.n4445 GNDA.n4444 0.0734167
R19890 GNDA.n4446 GNDA.n4445 0.0734167
R19891 GNDA.n4446 GNDA.n4330 0.0734167
R19892 GNDA.n4456 GNDA.n4328 0.0734167
R19893 GNDA.n4464 GNDA.n4328 0.0734167
R19894 GNDA.n4189 GNDA.n4188 0.0734167
R19895 GNDA.n4190 GNDA.n4189 0.0734167
R19896 GNDA.n4190 GNDA.n4182 0.0734167
R19897 GNDA.n4200 GNDA.n4180 0.0734167
R19898 GNDA.n4208 GNDA.n4180 0.0734167
R19899 GNDA.n4209 GNDA.n4208 0.0734167
R19900 GNDA.n4219 GNDA.n4218 0.0734167
R19901 GNDA.n4220 GNDA.n4219 0.0734167
R19902 GNDA.n4220 GNDA.n4176 0.0734167
R19903 GNDA.n4230 GNDA.n4174 0.0734167
R19904 GNDA.n4238 GNDA.n4174 0.0734167
R19905 GNDA.n4239 GNDA.n4238 0.0734167
R19906 GNDA.n4249 GNDA.n4248 0.0734167
R19907 GNDA.n4250 GNDA.n4249 0.0734167
R19908 GNDA.n4250 GNDA.n4170 0.0734167
R19909 GNDA.n4260 GNDA.n4168 0.0734167
R19910 GNDA.n4268 GNDA.n4168 0.0734167
R19911 GNDA.n4269 GNDA.n4268 0.0734167
R19912 GNDA.n4279 GNDA.n4278 0.0734167
R19913 GNDA.n4280 GNDA.n4279 0.0734167
R19914 GNDA.n4280 GNDA.n4164 0.0734167
R19915 GNDA.n4290 GNDA.n4162 0.0734167
R19916 GNDA.n4298 GNDA.n4162 0.0734167
R19917 GNDA.n3691 GNDA.n3690 0.0734167
R19918 GNDA.n3692 GNDA.n3691 0.0734167
R19919 GNDA.n3692 GNDA.n3506 0.0734167
R19920 GNDA.n3702 GNDA.n3504 0.0734167
R19921 GNDA.n3710 GNDA.n3504 0.0734167
R19922 GNDA.n3711 GNDA.n3710 0.0734167
R19923 GNDA.n3721 GNDA.n3720 0.0734167
R19924 GNDA.n3722 GNDA.n3721 0.0734167
R19925 GNDA.n3722 GNDA.n3500 0.0734167
R19926 GNDA.n3732 GNDA.n3498 0.0734167
R19927 GNDA.n3740 GNDA.n3498 0.0734167
R19928 GNDA.n3741 GNDA.n3740 0.0734167
R19929 GNDA.n3751 GNDA.n3750 0.0734167
R19930 GNDA.n3752 GNDA.n3751 0.0734167
R19931 GNDA.n3752 GNDA.n3494 0.0734167
R19932 GNDA.n3762 GNDA.n3492 0.0734167
R19933 GNDA.n3770 GNDA.n3492 0.0734167
R19934 GNDA.n3771 GNDA.n3770 0.0734167
R19935 GNDA.n3781 GNDA.n3780 0.0734167
R19936 GNDA.n3782 GNDA.n3781 0.0734167
R19937 GNDA.n3782 GNDA.n3488 0.0734167
R19938 GNDA.n3792 GNDA.n3486 0.0734167
R19939 GNDA.n3800 GNDA.n3486 0.0734167
R19940 GNDA.n4023 GNDA.n4022 0.0734167
R19941 GNDA.n4024 GNDA.n4023 0.0734167
R19942 GNDA.n4024 GNDA.n4016 0.0734167
R19943 GNDA.n4034 GNDA.n4014 0.0734167
R19944 GNDA.n4042 GNDA.n4014 0.0734167
R19945 GNDA.n4043 GNDA.n4042 0.0734167
R19946 GNDA.n4053 GNDA.n4052 0.0734167
R19947 GNDA.n4054 GNDA.n4053 0.0734167
R19948 GNDA.n4054 GNDA.n4010 0.0734167
R19949 GNDA.n4064 GNDA.n4008 0.0734167
R19950 GNDA.n4072 GNDA.n4008 0.0734167
R19951 GNDA.n4073 GNDA.n4072 0.0734167
R19952 GNDA.n4083 GNDA.n4082 0.0734167
R19953 GNDA.n4084 GNDA.n4083 0.0734167
R19954 GNDA.n4084 GNDA.n4004 0.0734167
R19955 GNDA.n4094 GNDA.n4002 0.0734167
R19956 GNDA.n4102 GNDA.n4002 0.0734167
R19957 GNDA.n4103 GNDA.n4102 0.0734167
R19958 GNDA.n4113 GNDA.n4112 0.0734167
R19959 GNDA.n4114 GNDA.n4113 0.0734167
R19960 GNDA.n4114 GNDA.n3998 0.0734167
R19961 GNDA.n4124 GNDA.n3996 0.0734167
R19962 GNDA.n4132 GNDA.n3996 0.0734167
R19963 GNDA.n3857 GNDA.n3856 0.0734167
R19964 GNDA.n3858 GNDA.n3857 0.0734167
R19965 GNDA.n3858 GNDA.n3850 0.0734167
R19966 GNDA.n3868 GNDA.n3848 0.0734167
R19967 GNDA.n3876 GNDA.n3848 0.0734167
R19968 GNDA.n3877 GNDA.n3876 0.0734167
R19969 GNDA.n3887 GNDA.n3886 0.0734167
R19970 GNDA.n3888 GNDA.n3887 0.0734167
R19971 GNDA.n3888 GNDA.n3844 0.0734167
R19972 GNDA.n3898 GNDA.n3842 0.0734167
R19973 GNDA.n3906 GNDA.n3842 0.0734167
R19974 GNDA.n3907 GNDA.n3906 0.0734167
R19975 GNDA.n3917 GNDA.n3916 0.0734167
R19976 GNDA.n3918 GNDA.n3917 0.0734167
R19977 GNDA.n3918 GNDA.n3838 0.0734167
R19978 GNDA.n3928 GNDA.n3836 0.0734167
R19979 GNDA.n3936 GNDA.n3836 0.0734167
R19980 GNDA.n3937 GNDA.n3936 0.0734167
R19981 GNDA.n3947 GNDA.n3946 0.0734167
R19982 GNDA.n3948 GNDA.n3947 0.0734167
R19983 GNDA.n3948 GNDA.n3832 0.0734167
R19984 GNDA.n3958 GNDA.n3830 0.0734167
R19985 GNDA.n3966 GNDA.n3830 0.0734167
R19986 GNDA.n3558 GNDA.n3511 0.0734167
R19987 GNDA.n3559 GNDA.n3558 0.0734167
R19988 GNDA.n3560 GNDA.n3559 0.0734167
R19989 GNDA.n3564 GNDA.n3563 0.0734167
R19990 GNDA.n3565 GNDA.n3564 0.0734167
R19991 GNDA.n3566 GNDA.n3565 0.0734167
R19992 GNDA.n3570 GNDA.n3569 0.0734167
R19993 GNDA.n3571 GNDA.n3570 0.0734167
R19994 GNDA.n3572 GNDA.n3571 0.0734167
R19995 GNDA.n3576 GNDA.n3575 0.0734167
R19996 GNDA.n3577 GNDA.n3576 0.0734167
R19997 GNDA.n3578 GNDA.n3577 0.0734167
R19998 GNDA.n3582 GNDA.n3581 0.0734167
R19999 GNDA.n3583 GNDA.n3582 0.0734167
R20000 GNDA.n3584 GNDA.n3583 0.0734167
R20001 GNDA.n3588 GNDA.n3587 0.0734167
R20002 GNDA.n3589 GNDA.n3588 0.0734167
R20003 GNDA.n3590 GNDA.n3589 0.0734167
R20004 GNDA.n3594 GNDA.n3593 0.0734167
R20005 GNDA.n3595 GNDA.n3594 0.0734167
R20006 GNDA.n3596 GNDA.n3595 0.0734167
R20007 GNDA.n3600 GNDA.n3599 0.0734167
R20008 GNDA.n3601 GNDA.n3600 0.0734167
R20009 GNDA.n452 GNDA.n405 0.0734167
R20010 GNDA.n453 GNDA.n452 0.0734167
R20011 GNDA.n454 GNDA.n453 0.0734167
R20012 GNDA.n458 GNDA.n457 0.0734167
R20013 GNDA.n459 GNDA.n458 0.0734167
R20014 GNDA.n460 GNDA.n459 0.0734167
R20015 GNDA.n464 GNDA.n463 0.0734167
R20016 GNDA.n465 GNDA.n464 0.0734167
R20017 GNDA.n466 GNDA.n465 0.0734167
R20018 GNDA.n470 GNDA.n469 0.0734167
R20019 GNDA.n471 GNDA.n470 0.0734167
R20020 GNDA.n472 GNDA.n471 0.0734167
R20021 GNDA.n476 GNDA.n475 0.0734167
R20022 GNDA.n477 GNDA.n476 0.0734167
R20023 GNDA.n478 GNDA.n477 0.0734167
R20024 GNDA.n482 GNDA.n481 0.0734167
R20025 GNDA.n483 GNDA.n482 0.0734167
R20026 GNDA.n484 GNDA.n483 0.0734167
R20027 GNDA.n488 GNDA.n487 0.0734167
R20028 GNDA.n489 GNDA.n488 0.0734167
R20029 GNDA.n490 GNDA.n489 0.0734167
R20030 GNDA.n494 GNDA.n493 0.0734167
R20031 GNDA.n495 GNDA.n494 0.0734167
R20032 GNDA.n5023 GNDA.n5022 0.0734167
R20033 GNDA.n5024 GNDA.n5023 0.0734167
R20034 GNDA.n5024 GNDA.n400 0.0734167
R20035 GNDA.n5034 GNDA.n398 0.0734167
R20036 GNDA.n5042 GNDA.n398 0.0734167
R20037 GNDA.n5043 GNDA.n5042 0.0734167
R20038 GNDA.n5053 GNDA.n5052 0.0734167
R20039 GNDA.n5054 GNDA.n5053 0.0734167
R20040 GNDA.n5054 GNDA.n394 0.0734167
R20041 GNDA.n5064 GNDA.n392 0.0734167
R20042 GNDA.n5072 GNDA.n392 0.0734167
R20043 GNDA.n5073 GNDA.n5072 0.0734167
R20044 GNDA.n5083 GNDA.n5082 0.0734167
R20045 GNDA.n5084 GNDA.n5083 0.0734167
R20046 GNDA.n5084 GNDA.n388 0.0734167
R20047 GNDA.n5094 GNDA.n386 0.0734167
R20048 GNDA.n5102 GNDA.n386 0.0734167
R20049 GNDA.n5103 GNDA.n5102 0.0734167
R20050 GNDA.n5113 GNDA.n5112 0.0734167
R20051 GNDA.n5114 GNDA.n5113 0.0734167
R20052 GNDA.n5114 GNDA.n382 0.0734167
R20053 GNDA.n5124 GNDA.n380 0.0734167
R20054 GNDA.n5132 GNDA.n380 0.0734167
R20055 GNDA.n3255 GNDA.n3208 0.0734167
R20056 GNDA.n3256 GNDA.n3255 0.0734167
R20057 GNDA.n3257 GNDA.n3256 0.0734167
R20058 GNDA.n3261 GNDA.n3260 0.0734167
R20059 GNDA.n3262 GNDA.n3261 0.0734167
R20060 GNDA.n3263 GNDA.n3262 0.0734167
R20061 GNDA.n3267 GNDA.n3266 0.0734167
R20062 GNDA.n3268 GNDA.n3267 0.0734167
R20063 GNDA.n3269 GNDA.n3268 0.0734167
R20064 GNDA.n3273 GNDA.n3272 0.0734167
R20065 GNDA.n3274 GNDA.n3273 0.0734167
R20066 GNDA.n3275 GNDA.n3274 0.0734167
R20067 GNDA.n3279 GNDA.n3278 0.0734167
R20068 GNDA.n3280 GNDA.n3279 0.0734167
R20069 GNDA.n3281 GNDA.n3280 0.0734167
R20070 GNDA.n3285 GNDA.n3284 0.0734167
R20071 GNDA.n3286 GNDA.n3285 0.0734167
R20072 GNDA.n3287 GNDA.n3286 0.0734167
R20073 GNDA.n3291 GNDA.n3290 0.0734167
R20074 GNDA.n3292 GNDA.n3291 0.0734167
R20075 GNDA.n3293 GNDA.n3292 0.0734167
R20076 GNDA.n3297 GNDA.n3296 0.0734167
R20077 GNDA.n3298 GNDA.n3297 0.0734167
R20078 GNDA.n3085 GNDA.n596 0.0734167
R20079 GNDA.n3086 GNDA.n3085 0.0734167
R20080 GNDA.n3086 GNDA.n3083 0.0734167
R20081 GNDA.n3096 GNDA.n3081 0.0734167
R20082 GNDA.n3104 GNDA.n3081 0.0734167
R20083 GNDA.n3105 GNDA.n3104 0.0734167
R20084 GNDA.n3115 GNDA.n3114 0.0734167
R20085 GNDA.n3116 GNDA.n3115 0.0734167
R20086 GNDA.n3116 GNDA.n3077 0.0734167
R20087 GNDA.n3126 GNDA.n3075 0.0734167
R20088 GNDA.n3134 GNDA.n3075 0.0734167
R20089 GNDA.n3135 GNDA.n3134 0.0734167
R20090 GNDA.n3145 GNDA.n3144 0.0734167
R20091 GNDA.n3146 GNDA.n3145 0.0734167
R20092 GNDA.n3146 GNDA.n3071 0.0734167
R20093 GNDA.n3156 GNDA.n3069 0.0734167
R20094 GNDA.n3164 GNDA.n3069 0.0734167
R20095 GNDA.n3165 GNDA.n3164 0.0734167
R20096 GNDA.n3175 GNDA.n3174 0.0734167
R20097 GNDA.n3176 GNDA.n3175 0.0734167
R20098 GNDA.n3176 GNDA.n3065 0.0734167
R20099 GNDA.n3186 GNDA.n3063 0.0734167
R20100 GNDA.n3194 GNDA.n3063 0.0734167
R20101 GNDA.n2925 GNDA.n2924 0.0734167
R20102 GNDA.n2926 GNDA.n2925 0.0734167
R20103 GNDA.n2926 GNDA.n2910 0.0734167
R20104 GNDA.n2936 GNDA.n2908 0.0734167
R20105 GNDA.n2944 GNDA.n2908 0.0734167
R20106 GNDA.n2945 GNDA.n2944 0.0734167
R20107 GNDA.n2955 GNDA.n2954 0.0734167
R20108 GNDA.n2956 GNDA.n2955 0.0734167
R20109 GNDA.n2956 GNDA.n2904 0.0734167
R20110 GNDA.n2966 GNDA.n2902 0.0734167
R20111 GNDA.n2974 GNDA.n2902 0.0734167
R20112 GNDA.n2975 GNDA.n2974 0.0734167
R20113 GNDA.n2985 GNDA.n2984 0.0734167
R20114 GNDA.n2986 GNDA.n2985 0.0734167
R20115 GNDA.n2986 GNDA.n2898 0.0734167
R20116 GNDA.n2996 GNDA.n2896 0.0734167
R20117 GNDA.n3004 GNDA.n2896 0.0734167
R20118 GNDA.n3005 GNDA.n3004 0.0734167
R20119 GNDA.n3015 GNDA.n3014 0.0734167
R20120 GNDA.n3016 GNDA.n3015 0.0734167
R20121 GNDA.n3016 GNDA.n2892 0.0734167
R20122 GNDA.n3026 GNDA.n2890 0.0734167
R20123 GNDA.n3034 GNDA.n2890 0.0734167
R20124 GNDA.n2289 GNDA.n2288 0.0734167
R20125 GNDA.n2290 GNDA.n2289 0.0734167
R20126 GNDA.n2290 GNDA.n712 0.0734167
R20127 GNDA.n2300 GNDA.n710 0.0734167
R20128 GNDA.n2308 GNDA.n710 0.0734167
R20129 GNDA.n2309 GNDA.n2308 0.0734167
R20130 GNDA.n2319 GNDA.n2318 0.0734167
R20131 GNDA.n2320 GNDA.n2319 0.0734167
R20132 GNDA.n2320 GNDA.n706 0.0734167
R20133 GNDA.n2330 GNDA.n704 0.0734167
R20134 GNDA.n2338 GNDA.n704 0.0734167
R20135 GNDA.n2339 GNDA.n2338 0.0734167
R20136 GNDA.n2349 GNDA.n2348 0.0734167
R20137 GNDA.n2350 GNDA.n2349 0.0734167
R20138 GNDA.n2350 GNDA.n700 0.0734167
R20139 GNDA.n2360 GNDA.n698 0.0734167
R20140 GNDA.n2368 GNDA.n698 0.0734167
R20141 GNDA.n2369 GNDA.n2368 0.0734167
R20142 GNDA.n2379 GNDA.n2378 0.0734167
R20143 GNDA.n2380 GNDA.n2379 0.0734167
R20144 GNDA.n2380 GNDA.n694 0.0734167
R20145 GNDA.n2390 GNDA.n692 0.0734167
R20146 GNDA.n2398 GNDA.n692 0.0734167
R20147 GNDA.n2751 GNDA.n2750 0.0734167
R20148 GNDA.n2752 GNDA.n2751 0.0734167
R20149 GNDA.n2752 GNDA.n646 0.0734167
R20150 GNDA.n2762 GNDA.n644 0.0734167
R20151 GNDA.n2770 GNDA.n644 0.0734167
R20152 GNDA.n2771 GNDA.n2770 0.0734167
R20153 GNDA.n2781 GNDA.n2780 0.0734167
R20154 GNDA.n2782 GNDA.n2781 0.0734167
R20155 GNDA.n2782 GNDA.n640 0.0734167
R20156 GNDA.n2792 GNDA.n638 0.0734167
R20157 GNDA.n2800 GNDA.n638 0.0734167
R20158 GNDA.n2801 GNDA.n2800 0.0734167
R20159 GNDA.n2811 GNDA.n2810 0.0734167
R20160 GNDA.n2812 GNDA.n2811 0.0734167
R20161 GNDA.n2812 GNDA.n634 0.0734167
R20162 GNDA.n2822 GNDA.n632 0.0734167
R20163 GNDA.n2830 GNDA.n632 0.0734167
R20164 GNDA.n2831 GNDA.n2830 0.0734167
R20165 GNDA.n2841 GNDA.n2840 0.0734167
R20166 GNDA.n2842 GNDA.n2841 0.0734167
R20167 GNDA.n2842 GNDA.n628 0.0734167
R20168 GNDA.n2852 GNDA.n626 0.0734167
R20169 GNDA.n2860 GNDA.n626 0.0734167
R20170 GNDA.n2618 GNDA.n2571 0.0734167
R20171 GNDA.n2619 GNDA.n2618 0.0734167
R20172 GNDA.n2620 GNDA.n2619 0.0734167
R20173 GNDA.n2624 GNDA.n2623 0.0734167
R20174 GNDA.n2625 GNDA.n2624 0.0734167
R20175 GNDA.n2626 GNDA.n2625 0.0734167
R20176 GNDA.n2630 GNDA.n2629 0.0734167
R20177 GNDA.n2631 GNDA.n2630 0.0734167
R20178 GNDA.n2632 GNDA.n2631 0.0734167
R20179 GNDA.n2636 GNDA.n2635 0.0734167
R20180 GNDA.n2637 GNDA.n2636 0.0734167
R20181 GNDA.n2638 GNDA.n2637 0.0734167
R20182 GNDA.n2642 GNDA.n2641 0.0734167
R20183 GNDA.n2643 GNDA.n2642 0.0734167
R20184 GNDA.n2644 GNDA.n2643 0.0734167
R20185 GNDA.n2648 GNDA.n2647 0.0734167
R20186 GNDA.n2649 GNDA.n2648 0.0734167
R20187 GNDA.n2650 GNDA.n2649 0.0734167
R20188 GNDA.n2654 GNDA.n2653 0.0734167
R20189 GNDA.n2655 GNDA.n2654 0.0734167
R20190 GNDA.n2656 GNDA.n2655 0.0734167
R20191 GNDA.n2660 GNDA.n2659 0.0734167
R20192 GNDA.n2661 GNDA.n2660 0.0734167
R20193 GNDA.n2449 GNDA.n662 0.0734167
R20194 GNDA.n2450 GNDA.n2449 0.0734167
R20195 GNDA.n2450 GNDA.n2447 0.0734167
R20196 GNDA.n2460 GNDA.n2445 0.0734167
R20197 GNDA.n2468 GNDA.n2445 0.0734167
R20198 GNDA.n2469 GNDA.n2468 0.0734167
R20199 GNDA.n2479 GNDA.n2478 0.0734167
R20200 GNDA.n2480 GNDA.n2479 0.0734167
R20201 GNDA.n2480 GNDA.n2441 0.0734167
R20202 GNDA.n2490 GNDA.n2439 0.0734167
R20203 GNDA.n2498 GNDA.n2439 0.0734167
R20204 GNDA.n2499 GNDA.n2498 0.0734167
R20205 GNDA.n2509 GNDA.n2508 0.0734167
R20206 GNDA.n2510 GNDA.n2509 0.0734167
R20207 GNDA.n2510 GNDA.n2435 0.0734167
R20208 GNDA.n2520 GNDA.n2433 0.0734167
R20209 GNDA.n2528 GNDA.n2433 0.0734167
R20210 GNDA.n2529 GNDA.n2528 0.0734167
R20211 GNDA.n2539 GNDA.n2538 0.0734167
R20212 GNDA.n2540 GNDA.n2539 0.0734167
R20213 GNDA.n2540 GNDA.n2429 0.0734167
R20214 GNDA.n2550 GNDA.n2427 0.0734167
R20215 GNDA.n2558 GNDA.n2427 0.0734167
R20216 GNDA.n2158 GNDA.n2111 0.0734167
R20217 GNDA.n2159 GNDA.n2158 0.0734167
R20218 GNDA.n2160 GNDA.n2159 0.0734167
R20219 GNDA.n2164 GNDA.n2163 0.0734167
R20220 GNDA.n2165 GNDA.n2164 0.0734167
R20221 GNDA.n2166 GNDA.n2165 0.0734167
R20222 GNDA.n2170 GNDA.n2169 0.0734167
R20223 GNDA.n2171 GNDA.n2170 0.0734167
R20224 GNDA.n2172 GNDA.n2171 0.0734167
R20225 GNDA.n2176 GNDA.n2175 0.0734167
R20226 GNDA.n2177 GNDA.n2176 0.0734167
R20227 GNDA.n2178 GNDA.n2177 0.0734167
R20228 GNDA.n2182 GNDA.n2181 0.0734167
R20229 GNDA.n2183 GNDA.n2182 0.0734167
R20230 GNDA.n2184 GNDA.n2183 0.0734167
R20231 GNDA.n2188 GNDA.n2187 0.0734167
R20232 GNDA.n2189 GNDA.n2188 0.0734167
R20233 GNDA.n2190 GNDA.n2189 0.0734167
R20234 GNDA.n2194 GNDA.n2193 0.0734167
R20235 GNDA.n2195 GNDA.n2194 0.0734167
R20236 GNDA.n2196 GNDA.n2195 0.0734167
R20237 GNDA.n2200 GNDA.n2199 0.0734167
R20238 GNDA.n2201 GNDA.n2200 0.0734167
R20239 GNDA.n1986 GNDA.n725 0.0734167
R20240 GNDA.n1987 GNDA.n1986 0.0734167
R20241 GNDA.n1987 GNDA.n1984 0.0734167
R20242 GNDA.n1997 GNDA.n1982 0.0734167
R20243 GNDA.n2005 GNDA.n1982 0.0734167
R20244 GNDA.n2006 GNDA.n2005 0.0734167
R20245 GNDA.n2016 GNDA.n2015 0.0734167
R20246 GNDA.n2017 GNDA.n2016 0.0734167
R20247 GNDA.n2017 GNDA.n1978 0.0734167
R20248 GNDA.n2027 GNDA.n1976 0.0734167
R20249 GNDA.n2035 GNDA.n1976 0.0734167
R20250 GNDA.n2036 GNDA.n2035 0.0734167
R20251 GNDA.n2046 GNDA.n2045 0.0734167
R20252 GNDA.n2047 GNDA.n2046 0.0734167
R20253 GNDA.n2047 GNDA.n1972 0.0734167
R20254 GNDA.n2057 GNDA.n1970 0.0734167
R20255 GNDA.n2065 GNDA.n1970 0.0734167
R20256 GNDA.n2066 GNDA.n2065 0.0734167
R20257 GNDA.n2076 GNDA.n2075 0.0734167
R20258 GNDA.n2077 GNDA.n2076 0.0734167
R20259 GNDA.n2077 GNDA.n1966 0.0734167
R20260 GNDA.n2087 GNDA.n1964 0.0734167
R20261 GNDA.n2095 GNDA.n1964 0.0734167
R20262 GNDA.n1826 GNDA.n1825 0.0734167
R20263 GNDA.n1827 GNDA.n1826 0.0734167
R20264 GNDA.n1827 GNDA.n775 0.0734167
R20265 GNDA.n1837 GNDA.n773 0.0734167
R20266 GNDA.n1845 GNDA.n773 0.0734167
R20267 GNDA.n1846 GNDA.n1845 0.0734167
R20268 GNDA.n1856 GNDA.n1855 0.0734167
R20269 GNDA.n1857 GNDA.n1856 0.0734167
R20270 GNDA.n1857 GNDA.n769 0.0734167
R20271 GNDA.n1867 GNDA.n767 0.0734167
R20272 GNDA.n1875 GNDA.n767 0.0734167
R20273 GNDA.n1876 GNDA.n1875 0.0734167
R20274 GNDA.n1886 GNDA.n1885 0.0734167
R20275 GNDA.n1887 GNDA.n1886 0.0734167
R20276 GNDA.n1887 GNDA.n763 0.0734167
R20277 GNDA.n1897 GNDA.n761 0.0734167
R20278 GNDA.n1905 GNDA.n761 0.0734167
R20279 GNDA.n1906 GNDA.n1905 0.0734167
R20280 GNDA.n1916 GNDA.n1915 0.0734167
R20281 GNDA.n1917 GNDA.n1916 0.0734167
R20282 GNDA.n1917 GNDA.n757 0.0734167
R20283 GNDA.n1927 GNDA.n755 0.0734167
R20284 GNDA.n1935 GNDA.n755 0.0734167
R20285 GNDA.n1571 GNDA.n1524 0.0734167
R20286 GNDA.n1572 GNDA.n1571 0.0734167
R20287 GNDA.n1573 GNDA.n1572 0.0734167
R20288 GNDA.n1577 GNDA.n1576 0.0734167
R20289 GNDA.n1578 GNDA.n1577 0.0734167
R20290 GNDA.n1579 GNDA.n1578 0.0734167
R20291 GNDA.n1583 GNDA.n1582 0.0734167
R20292 GNDA.n1584 GNDA.n1583 0.0734167
R20293 GNDA.n1585 GNDA.n1584 0.0734167
R20294 GNDA.n1589 GNDA.n1588 0.0734167
R20295 GNDA.n1590 GNDA.n1589 0.0734167
R20296 GNDA.n1591 GNDA.n1590 0.0734167
R20297 GNDA.n1595 GNDA.n1594 0.0734167
R20298 GNDA.n1596 GNDA.n1595 0.0734167
R20299 GNDA.n1597 GNDA.n1596 0.0734167
R20300 GNDA.n1601 GNDA.n1600 0.0734167
R20301 GNDA.n1602 GNDA.n1601 0.0734167
R20302 GNDA.n1603 GNDA.n1602 0.0734167
R20303 GNDA.n1607 GNDA.n1606 0.0734167
R20304 GNDA.n1608 GNDA.n1607 0.0734167
R20305 GNDA.n1609 GNDA.n1608 0.0734167
R20306 GNDA.n1613 GNDA.n1612 0.0734167
R20307 GNDA.n1614 GNDA.n1613 0.0734167
R20308 GNDA.n1402 GNDA.n791 0.0734167
R20309 GNDA.n1403 GNDA.n1402 0.0734167
R20310 GNDA.n1403 GNDA.n1400 0.0734167
R20311 GNDA.n1413 GNDA.n1398 0.0734167
R20312 GNDA.n1421 GNDA.n1398 0.0734167
R20313 GNDA.n1422 GNDA.n1421 0.0734167
R20314 GNDA.n1432 GNDA.n1431 0.0734167
R20315 GNDA.n1433 GNDA.n1432 0.0734167
R20316 GNDA.n1433 GNDA.n1394 0.0734167
R20317 GNDA.n1443 GNDA.n1392 0.0734167
R20318 GNDA.n1451 GNDA.n1392 0.0734167
R20319 GNDA.n1452 GNDA.n1451 0.0734167
R20320 GNDA.n1462 GNDA.n1461 0.0734167
R20321 GNDA.n1463 GNDA.n1462 0.0734167
R20322 GNDA.n1463 GNDA.n1388 0.0734167
R20323 GNDA.n1473 GNDA.n1386 0.0734167
R20324 GNDA.n1481 GNDA.n1386 0.0734167
R20325 GNDA.n1482 GNDA.n1481 0.0734167
R20326 GNDA.n1492 GNDA.n1491 0.0734167
R20327 GNDA.n1493 GNDA.n1492 0.0734167
R20328 GNDA.n1493 GNDA.n1382 0.0734167
R20329 GNDA.n1503 GNDA.n1380 0.0734167
R20330 GNDA.n1511 GNDA.n1380 0.0734167
R20331 GNDA.n1240 GNDA.n1214 0.0734167
R20332 GNDA.n1248 GNDA.n1214 0.0734167
R20333 GNDA.n1249 GNDA.n1248 0.0734167
R20334 GNDA.n1259 GNDA.n1258 0.0734167
R20335 GNDA.n1260 GNDA.n1259 0.0734167
R20336 GNDA.n1260 GNDA.n1210 0.0734167
R20337 GNDA.n1270 GNDA.n1208 0.0734167
R20338 GNDA.n1278 GNDA.n1208 0.0734167
R20339 GNDA.n1279 GNDA.n1278 0.0734167
R20340 GNDA.n1289 GNDA.n1288 0.0734167
R20341 GNDA.n1290 GNDA.n1289 0.0734167
R20342 GNDA.n1290 GNDA.n1204 0.0734167
R20343 GNDA.n1300 GNDA.n1202 0.0734167
R20344 GNDA.n1308 GNDA.n1202 0.0734167
R20345 GNDA.n1309 GNDA.n1308 0.0734167
R20346 GNDA.n1319 GNDA.n1318 0.0734167
R20347 GNDA.n1320 GNDA.n1319 0.0734167
R20348 GNDA.n1320 GNDA.n1198 0.0734167
R20349 GNDA.n1330 GNDA.n1196 0.0734167
R20350 GNDA.n1338 GNDA.n1196 0.0734167
R20351 GNDA.n1339 GNDA.n1338 0.0734167
R20352 GNDA.n1348 GNDA.n1347 0.0734167
R20353 GNDA.n1350 GNDA.n1348 0.0734167
R20354 GNDA.n1813 GNDA.n1693 0.0734167
R20355 GNDA.n4986 GNDA.n4985 0.0734167
R20356 GNDA.n7139 GNDA.n7131 0.0734167
R20357 GNDA.n7140 GNDA.n7139 0.0734167
R20358 GNDA.n7148 GNDA.n7147 0.0734167
R20359 GNDA.n7149 GNDA.n7148 0.0734167
R20360 GNDA.n7149 GNDA.n7123 0.0734167
R20361 GNDA.n7157 GNDA.n7119 0.0734167
R20362 GNDA.n7163 GNDA.n7119 0.0734167
R20363 GNDA.n7164 GNDA.n7163 0.0734167
R20364 GNDA.n7172 GNDA.n7171 0.0734167
R20365 GNDA.n7173 GNDA.n7172 0.0734167
R20366 GNDA.n7173 GNDA.n7111 0.0734167
R20367 GNDA.n7181 GNDA.n7107 0.0734167
R20368 GNDA.n7187 GNDA.n7107 0.0734167
R20369 GNDA.n7188 GNDA.n7187 0.0734167
R20370 GNDA.n7196 GNDA.n7195 0.0734167
R20371 GNDA.n7197 GNDA.n7196 0.0734167
R20372 GNDA.n7197 GNDA.n7099 0.0734167
R20373 GNDA.n7205 GNDA.n7095 0.0734167
R20374 GNDA.n7211 GNDA.n7095 0.0734167
R20375 GNDA.n7212 GNDA.n7211 0.0734167
R20376 GNDA.n7220 GNDA.n7219 0.0734167
R20377 GNDA.n7221 GNDA.n7220 0.0734167
R20378 GNDA.n7221 GNDA.n95 0.0734167
R20379 GNDA.n1354 GNDA.n1166 0.0682094
R20380 GNDA.n5275 GNDA.n326 0.0682083
R20381 GNDA.n5169 GNDA.n5158 0.0682083
R20382 GNDA.n5171 GNDA.n5170 0.0682083
R20383 GNDA.n5181 GNDA.n5180 0.0682083
R20384 GNDA.n5189 GNDA.n5154 0.0682083
R20385 GNDA.n5199 GNDA.n5152 0.0682083
R20386 GNDA.n5201 GNDA.n5200 0.0682083
R20387 GNDA.n5211 GNDA.n5210 0.0682083
R20388 GNDA.n5219 GNDA.n5148 0.0682083
R20389 GNDA.n5229 GNDA.n5146 0.0682083
R20390 GNDA.n5231 GNDA.n5230 0.0682083
R20391 GNDA.n5241 GNDA.n5240 0.0682083
R20392 GNDA.n5249 GNDA.n5142 0.0682083
R20393 GNDA.n5259 GNDA.n5140 0.0682083
R20394 GNDA.n5261 GNDA.n5260 0.0682083
R20395 GNDA.n4962 GNDA.n3456 0.0682083
R20396 GNDA.n4856 GNDA.n4845 0.0682083
R20397 GNDA.n4858 GNDA.n4857 0.0682083
R20398 GNDA.n4868 GNDA.n4867 0.0682083
R20399 GNDA.n4876 GNDA.n4841 0.0682083
R20400 GNDA.n4886 GNDA.n4839 0.0682083
R20401 GNDA.n4888 GNDA.n4887 0.0682083
R20402 GNDA.n4898 GNDA.n4897 0.0682083
R20403 GNDA.n4906 GNDA.n4835 0.0682083
R20404 GNDA.n4916 GNDA.n4833 0.0682083
R20405 GNDA.n4918 GNDA.n4917 0.0682083
R20406 GNDA.n4928 GNDA.n4927 0.0682083
R20407 GNDA.n4936 GNDA.n4829 0.0682083
R20408 GNDA.n4946 GNDA.n4827 0.0682083
R20409 GNDA.n4948 GNDA.n4947 0.0682083
R20410 GNDA.n4686 GNDA.n4682 0.0682083
R20411 GNDA.n4696 GNDA.n4680 0.0682083
R20412 GNDA.n4698 GNDA.n4697 0.0682083
R20413 GNDA.n4708 GNDA.n4707 0.0682083
R20414 GNDA.n4716 GNDA.n4676 0.0682083
R20415 GNDA.n4726 GNDA.n4674 0.0682083
R20416 GNDA.n4728 GNDA.n4727 0.0682083
R20417 GNDA.n4738 GNDA.n4737 0.0682083
R20418 GNDA.n4746 GNDA.n4670 0.0682083
R20419 GNDA.n4756 GNDA.n4668 0.0682083
R20420 GNDA.n4758 GNDA.n4757 0.0682083
R20421 GNDA.n4768 GNDA.n4767 0.0682083
R20422 GNDA.n4776 GNDA.n4664 0.0682083
R20423 GNDA.n4786 GNDA.n4662 0.0682083
R20424 GNDA.n4788 GNDA.n4787 0.0682083
R20425 GNDA.n4520 GNDA.n4516 0.0682083
R20426 GNDA.n4530 GNDA.n4514 0.0682083
R20427 GNDA.n4532 GNDA.n4531 0.0682083
R20428 GNDA.n4542 GNDA.n4541 0.0682083
R20429 GNDA.n4550 GNDA.n4510 0.0682083
R20430 GNDA.n4560 GNDA.n4508 0.0682083
R20431 GNDA.n4562 GNDA.n4561 0.0682083
R20432 GNDA.n4572 GNDA.n4571 0.0682083
R20433 GNDA.n4580 GNDA.n4504 0.0682083
R20434 GNDA.n4590 GNDA.n4502 0.0682083
R20435 GNDA.n4592 GNDA.n4591 0.0682083
R20436 GNDA.n4602 GNDA.n4601 0.0682083
R20437 GNDA.n4610 GNDA.n4498 0.0682083
R20438 GNDA.n4620 GNDA.n4496 0.0682083
R20439 GNDA.n4622 GNDA.n4621 0.0682083
R20440 GNDA.n4354 GNDA.n4350 0.0682083
R20441 GNDA.n4364 GNDA.n4348 0.0682083
R20442 GNDA.n4366 GNDA.n4365 0.0682083
R20443 GNDA.n4376 GNDA.n4375 0.0682083
R20444 GNDA.n4384 GNDA.n4344 0.0682083
R20445 GNDA.n4394 GNDA.n4342 0.0682083
R20446 GNDA.n4396 GNDA.n4395 0.0682083
R20447 GNDA.n4406 GNDA.n4405 0.0682083
R20448 GNDA.n4414 GNDA.n4338 0.0682083
R20449 GNDA.n4424 GNDA.n4336 0.0682083
R20450 GNDA.n4426 GNDA.n4425 0.0682083
R20451 GNDA.n4436 GNDA.n4435 0.0682083
R20452 GNDA.n4444 GNDA.n4332 0.0682083
R20453 GNDA.n4454 GNDA.n4330 0.0682083
R20454 GNDA.n4456 GNDA.n4455 0.0682083
R20455 GNDA.n4188 GNDA.n4184 0.0682083
R20456 GNDA.n4198 GNDA.n4182 0.0682083
R20457 GNDA.n4200 GNDA.n4199 0.0682083
R20458 GNDA.n4210 GNDA.n4209 0.0682083
R20459 GNDA.n4218 GNDA.n4178 0.0682083
R20460 GNDA.n4228 GNDA.n4176 0.0682083
R20461 GNDA.n4230 GNDA.n4229 0.0682083
R20462 GNDA.n4240 GNDA.n4239 0.0682083
R20463 GNDA.n4248 GNDA.n4172 0.0682083
R20464 GNDA.n4258 GNDA.n4170 0.0682083
R20465 GNDA.n4260 GNDA.n4259 0.0682083
R20466 GNDA.n4270 GNDA.n4269 0.0682083
R20467 GNDA.n4278 GNDA.n4166 0.0682083
R20468 GNDA.n4288 GNDA.n4164 0.0682083
R20469 GNDA.n4290 GNDA.n4289 0.0682083
R20470 GNDA.n3690 GNDA.n3686 0.0682083
R20471 GNDA.n3700 GNDA.n3506 0.0682083
R20472 GNDA.n3702 GNDA.n3701 0.0682083
R20473 GNDA.n3712 GNDA.n3711 0.0682083
R20474 GNDA.n3720 GNDA.n3502 0.0682083
R20475 GNDA.n3730 GNDA.n3500 0.0682083
R20476 GNDA.n3732 GNDA.n3731 0.0682083
R20477 GNDA.n3742 GNDA.n3741 0.0682083
R20478 GNDA.n3750 GNDA.n3496 0.0682083
R20479 GNDA.n3760 GNDA.n3494 0.0682083
R20480 GNDA.n3762 GNDA.n3761 0.0682083
R20481 GNDA.n3772 GNDA.n3771 0.0682083
R20482 GNDA.n3780 GNDA.n3490 0.0682083
R20483 GNDA.n3790 GNDA.n3488 0.0682083
R20484 GNDA.n3792 GNDA.n3791 0.0682083
R20485 GNDA.n4022 GNDA.n4018 0.0682083
R20486 GNDA.n4032 GNDA.n4016 0.0682083
R20487 GNDA.n4034 GNDA.n4033 0.0682083
R20488 GNDA.n4044 GNDA.n4043 0.0682083
R20489 GNDA.n4052 GNDA.n4012 0.0682083
R20490 GNDA.n4062 GNDA.n4010 0.0682083
R20491 GNDA.n4064 GNDA.n4063 0.0682083
R20492 GNDA.n4074 GNDA.n4073 0.0682083
R20493 GNDA.n4082 GNDA.n4006 0.0682083
R20494 GNDA.n4092 GNDA.n4004 0.0682083
R20495 GNDA.n4094 GNDA.n4093 0.0682083
R20496 GNDA.n4104 GNDA.n4103 0.0682083
R20497 GNDA.n4112 GNDA.n4000 0.0682083
R20498 GNDA.n4122 GNDA.n3998 0.0682083
R20499 GNDA.n4124 GNDA.n4123 0.0682083
R20500 GNDA.n3856 GNDA.n3852 0.0682083
R20501 GNDA.n3866 GNDA.n3850 0.0682083
R20502 GNDA.n3868 GNDA.n3867 0.0682083
R20503 GNDA.n3878 GNDA.n3877 0.0682083
R20504 GNDA.n3886 GNDA.n3846 0.0682083
R20505 GNDA.n3896 GNDA.n3844 0.0682083
R20506 GNDA.n3898 GNDA.n3897 0.0682083
R20507 GNDA.n3908 GNDA.n3907 0.0682083
R20508 GNDA.n3916 GNDA.n3840 0.0682083
R20509 GNDA.n3926 GNDA.n3838 0.0682083
R20510 GNDA.n3928 GNDA.n3927 0.0682083
R20511 GNDA.n3938 GNDA.n3937 0.0682083
R20512 GNDA.n3946 GNDA.n3834 0.0682083
R20513 GNDA.n3956 GNDA.n3832 0.0682083
R20514 GNDA.n3958 GNDA.n3957 0.0682083
R20515 GNDA.n3675 GNDA.n3511 0.0682083
R20516 GNDA.n3561 GNDA.n3560 0.0682083
R20517 GNDA.n3563 GNDA.n3562 0.0682083
R20518 GNDA.n3567 GNDA.n3566 0.0682083
R20519 GNDA.n3569 GNDA.n3568 0.0682083
R20520 GNDA.n3573 GNDA.n3572 0.0682083
R20521 GNDA.n3575 GNDA.n3574 0.0682083
R20522 GNDA.n3579 GNDA.n3578 0.0682083
R20523 GNDA.n3581 GNDA.n3580 0.0682083
R20524 GNDA.n3585 GNDA.n3584 0.0682083
R20525 GNDA.n3587 GNDA.n3586 0.0682083
R20526 GNDA.n3591 GNDA.n3590 0.0682083
R20527 GNDA.n3593 GNDA.n3592 0.0682083
R20528 GNDA.n3597 GNDA.n3596 0.0682083
R20529 GNDA.n3599 GNDA.n3598 0.0682083
R20530 GNDA.n569 GNDA.n405 0.0682083
R20531 GNDA.n455 GNDA.n454 0.0682083
R20532 GNDA.n457 GNDA.n456 0.0682083
R20533 GNDA.n461 GNDA.n460 0.0682083
R20534 GNDA.n463 GNDA.n462 0.0682083
R20535 GNDA.n467 GNDA.n466 0.0682083
R20536 GNDA.n469 GNDA.n468 0.0682083
R20537 GNDA.n473 GNDA.n472 0.0682083
R20538 GNDA.n475 GNDA.n474 0.0682083
R20539 GNDA.n479 GNDA.n478 0.0682083
R20540 GNDA.n481 GNDA.n480 0.0682083
R20541 GNDA.n485 GNDA.n484 0.0682083
R20542 GNDA.n487 GNDA.n486 0.0682083
R20543 GNDA.n491 GNDA.n490 0.0682083
R20544 GNDA.n493 GNDA.n492 0.0682083
R20545 GNDA.n5022 GNDA.n5018 0.0682083
R20546 GNDA.n5032 GNDA.n400 0.0682083
R20547 GNDA.n5034 GNDA.n5033 0.0682083
R20548 GNDA.n5044 GNDA.n5043 0.0682083
R20549 GNDA.n5052 GNDA.n396 0.0682083
R20550 GNDA.n5062 GNDA.n394 0.0682083
R20551 GNDA.n5064 GNDA.n5063 0.0682083
R20552 GNDA.n5074 GNDA.n5073 0.0682083
R20553 GNDA.n5082 GNDA.n390 0.0682083
R20554 GNDA.n5092 GNDA.n388 0.0682083
R20555 GNDA.n5094 GNDA.n5093 0.0682083
R20556 GNDA.n5104 GNDA.n5103 0.0682083
R20557 GNDA.n5112 GNDA.n384 0.0682083
R20558 GNDA.n5122 GNDA.n382 0.0682083
R20559 GNDA.n5124 GNDA.n5123 0.0682083
R20560 GNDA.n3372 GNDA.n3208 0.0682083
R20561 GNDA.n3258 GNDA.n3257 0.0682083
R20562 GNDA.n3260 GNDA.n3259 0.0682083
R20563 GNDA.n3264 GNDA.n3263 0.0682083
R20564 GNDA.n3266 GNDA.n3265 0.0682083
R20565 GNDA.n3270 GNDA.n3269 0.0682083
R20566 GNDA.n3272 GNDA.n3271 0.0682083
R20567 GNDA.n3276 GNDA.n3275 0.0682083
R20568 GNDA.n3278 GNDA.n3277 0.0682083
R20569 GNDA.n3282 GNDA.n3281 0.0682083
R20570 GNDA.n3284 GNDA.n3283 0.0682083
R20571 GNDA.n3288 GNDA.n3287 0.0682083
R20572 GNDA.n3290 GNDA.n3289 0.0682083
R20573 GNDA.n3294 GNDA.n3293 0.0682083
R20574 GNDA.n3296 GNDA.n3295 0.0682083
R20575 GNDA.n3200 GNDA.n596 0.0682083
R20576 GNDA.n3094 GNDA.n3083 0.0682083
R20577 GNDA.n3096 GNDA.n3095 0.0682083
R20578 GNDA.n3106 GNDA.n3105 0.0682083
R20579 GNDA.n3114 GNDA.n3079 0.0682083
R20580 GNDA.n3124 GNDA.n3077 0.0682083
R20581 GNDA.n3126 GNDA.n3125 0.0682083
R20582 GNDA.n3136 GNDA.n3135 0.0682083
R20583 GNDA.n3144 GNDA.n3073 0.0682083
R20584 GNDA.n3154 GNDA.n3071 0.0682083
R20585 GNDA.n3156 GNDA.n3155 0.0682083
R20586 GNDA.n3166 GNDA.n3165 0.0682083
R20587 GNDA.n3174 GNDA.n3067 0.0682083
R20588 GNDA.n3184 GNDA.n3065 0.0682083
R20589 GNDA.n3186 GNDA.n3185 0.0682083
R20590 GNDA.n2924 GNDA.n2920 0.0682083
R20591 GNDA.n2934 GNDA.n2910 0.0682083
R20592 GNDA.n2936 GNDA.n2935 0.0682083
R20593 GNDA.n2946 GNDA.n2945 0.0682083
R20594 GNDA.n2954 GNDA.n2906 0.0682083
R20595 GNDA.n2964 GNDA.n2904 0.0682083
R20596 GNDA.n2966 GNDA.n2965 0.0682083
R20597 GNDA.n2976 GNDA.n2975 0.0682083
R20598 GNDA.n2984 GNDA.n2900 0.0682083
R20599 GNDA.n2994 GNDA.n2898 0.0682083
R20600 GNDA.n2996 GNDA.n2995 0.0682083
R20601 GNDA.n3006 GNDA.n3005 0.0682083
R20602 GNDA.n3014 GNDA.n2894 0.0682083
R20603 GNDA.n3024 GNDA.n2892 0.0682083
R20604 GNDA.n3026 GNDA.n3025 0.0682083
R20605 GNDA.n2288 GNDA.n2284 0.0682083
R20606 GNDA.n2298 GNDA.n712 0.0682083
R20607 GNDA.n2300 GNDA.n2299 0.0682083
R20608 GNDA.n2310 GNDA.n2309 0.0682083
R20609 GNDA.n2318 GNDA.n708 0.0682083
R20610 GNDA.n2328 GNDA.n706 0.0682083
R20611 GNDA.n2330 GNDA.n2329 0.0682083
R20612 GNDA.n2340 GNDA.n2339 0.0682083
R20613 GNDA.n2348 GNDA.n702 0.0682083
R20614 GNDA.n2358 GNDA.n700 0.0682083
R20615 GNDA.n2360 GNDA.n2359 0.0682083
R20616 GNDA.n2370 GNDA.n2369 0.0682083
R20617 GNDA.n2378 GNDA.n696 0.0682083
R20618 GNDA.n2388 GNDA.n694 0.0682083
R20619 GNDA.n2390 GNDA.n2389 0.0682083
R20620 GNDA.n2750 GNDA.n2746 0.0682083
R20621 GNDA.n2760 GNDA.n646 0.0682083
R20622 GNDA.n2762 GNDA.n2761 0.0682083
R20623 GNDA.n2772 GNDA.n2771 0.0682083
R20624 GNDA.n2780 GNDA.n642 0.0682083
R20625 GNDA.n2790 GNDA.n640 0.0682083
R20626 GNDA.n2792 GNDA.n2791 0.0682083
R20627 GNDA.n2802 GNDA.n2801 0.0682083
R20628 GNDA.n2810 GNDA.n636 0.0682083
R20629 GNDA.n2820 GNDA.n634 0.0682083
R20630 GNDA.n2822 GNDA.n2821 0.0682083
R20631 GNDA.n2832 GNDA.n2831 0.0682083
R20632 GNDA.n2840 GNDA.n630 0.0682083
R20633 GNDA.n2850 GNDA.n628 0.0682083
R20634 GNDA.n2852 GNDA.n2851 0.0682083
R20635 GNDA.n2735 GNDA.n2571 0.0682083
R20636 GNDA.n2621 GNDA.n2620 0.0682083
R20637 GNDA.n2623 GNDA.n2622 0.0682083
R20638 GNDA.n2627 GNDA.n2626 0.0682083
R20639 GNDA.n2629 GNDA.n2628 0.0682083
R20640 GNDA.n2633 GNDA.n2632 0.0682083
R20641 GNDA.n2635 GNDA.n2634 0.0682083
R20642 GNDA.n2639 GNDA.n2638 0.0682083
R20643 GNDA.n2641 GNDA.n2640 0.0682083
R20644 GNDA.n2645 GNDA.n2644 0.0682083
R20645 GNDA.n2647 GNDA.n2646 0.0682083
R20646 GNDA.n2651 GNDA.n2650 0.0682083
R20647 GNDA.n2653 GNDA.n2652 0.0682083
R20648 GNDA.n2657 GNDA.n2656 0.0682083
R20649 GNDA.n2659 GNDA.n2658 0.0682083
R20650 GNDA.n2564 GNDA.n662 0.0682083
R20651 GNDA.n2458 GNDA.n2447 0.0682083
R20652 GNDA.n2460 GNDA.n2459 0.0682083
R20653 GNDA.n2470 GNDA.n2469 0.0682083
R20654 GNDA.n2478 GNDA.n2443 0.0682083
R20655 GNDA.n2488 GNDA.n2441 0.0682083
R20656 GNDA.n2490 GNDA.n2489 0.0682083
R20657 GNDA.n2500 GNDA.n2499 0.0682083
R20658 GNDA.n2508 GNDA.n2437 0.0682083
R20659 GNDA.n2518 GNDA.n2435 0.0682083
R20660 GNDA.n2520 GNDA.n2519 0.0682083
R20661 GNDA.n2530 GNDA.n2529 0.0682083
R20662 GNDA.n2538 GNDA.n2431 0.0682083
R20663 GNDA.n2548 GNDA.n2429 0.0682083
R20664 GNDA.n2550 GNDA.n2549 0.0682083
R20665 GNDA.n2275 GNDA.n2111 0.0682083
R20666 GNDA.n2161 GNDA.n2160 0.0682083
R20667 GNDA.n2163 GNDA.n2162 0.0682083
R20668 GNDA.n2167 GNDA.n2166 0.0682083
R20669 GNDA.n2169 GNDA.n2168 0.0682083
R20670 GNDA.n2173 GNDA.n2172 0.0682083
R20671 GNDA.n2175 GNDA.n2174 0.0682083
R20672 GNDA.n2179 GNDA.n2178 0.0682083
R20673 GNDA.n2181 GNDA.n2180 0.0682083
R20674 GNDA.n2185 GNDA.n2184 0.0682083
R20675 GNDA.n2187 GNDA.n2186 0.0682083
R20676 GNDA.n2191 GNDA.n2190 0.0682083
R20677 GNDA.n2193 GNDA.n2192 0.0682083
R20678 GNDA.n2197 GNDA.n2196 0.0682083
R20679 GNDA.n2199 GNDA.n2198 0.0682083
R20680 GNDA.n2101 GNDA.n725 0.0682083
R20681 GNDA.n1995 GNDA.n1984 0.0682083
R20682 GNDA.n1997 GNDA.n1996 0.0682083
R20683 GNDA.n2007 GNDA.n2006 0.0682083
R20684 GNDA.n2015 GNDA.n1980 0.0682083
R20685 GNDA.n2025 GNDA.n1978 0.0682083
R20686 GNDA.n2027 GNDA.n2026 0.0682083
R20687 GNDA.n2037 GNDA.n2036 0.0682083
R20688 GNDA.n2045 GNDA.n1974 0.0682083
R20689 GNDA.n2055 GNDA.n1972 0.0682083
R20690 GNDA.n2057 GNDA.n2056 0.0682083
R20691 GNDA.n2067 GNDA.n2066 0.0682083
R20692 GNDA.n2075 GNDA.n1968 0.0682083
R20693 GNDA.n2085 GNDA.n1966 0.0682083
R20694 GNDA.n2087 GNDA.n2086 0.0682083
R20695 GNDA.n1825 GNDA.n1821 0.0682083
R20696 GNDA.n1835 GNDA.n775 0.0682083
R20697 GNDA.n1837 GNDA.n1836 0.0682083
R20698 GNDA.n1847 GNDA.n1846 0.0682083
R20699 GNDA.n1855 GNDA.n771 0.0682083
R20700 GNDA.n1865 GNDA.n769 0.0682083
R20701 GNDA.n1867 GNDA.n1866 0.0682083
R20702 GNDA.n1877 GNDA.n1876 0.0682083
R20703 GNDA.n1885 GNDA.n765 0.0682083
R20704 GNDA.n1895 GNDA.n763 0.0682083
R20705 GNDA.n1897 GNDA.n1896 0.0682083
R20706 GNDA.n1907 GNDA.n1906 0.0682083
R20707 GNDA.n1915 GNDA.n759 0.0682083
R20708 GNDA.n1925 GNDA.n757 0.0682083
R20709 GNDA.n1927 GNDA.n1926 0.0682083
R20710 GNDA.n1688 GNDA.n1524 0.0682083
R20711 GNDA.n1574 GNDA.n1573 0.0682083
R20712 GNDA.n1576 GNDA.n1575 0.0682083
R20713 GNDA.n1580 GNDA.n1579 0.0682083
R20714 GNDA.n1582 GNDA.n1581 0.0682083
R20715 GNDA.n1586 GNDA.n1585 0.0682083
R20716 GNDA.n1588 GNDA.n1587 0.0682083
R20717 GNDA.n1592 GNDA.n1591 0.0682083
R20718 GNDA.n1594 GNDA.n1593 0.0682083
R20719 GNDA.n1598 GNDA.n1597 0.0682083
R20720 GNDA.n1600 GNDA.n1599 0.0682083
R20721 GNDA.n1604 GNDA.n1603 0.0682083
R20722 GNDA.n1606 GNDA.n1605 0.0682083
R20723 GNDA.n1610 GNDA.n1609 0.0682083
R20724 GNDA.n1612 GNDA.n1611 0.0682083
R20725 GNDA.n1517 GNDA.n791 0.0682083
R20726 GNDA.n1411 GNDA.n1400 0.0682083
R20727 GNDA.n1413 GNDA.n1412 0.0682083
R20728 GNDA.n1423 GNDA.n1422 0.0682083
R20729 GNDA.n1431 GNDA.n1396 0.0682083
R20730 GNDA.n1441 GNDA.n1394 0.0682083
R20731 GNDA.n1443 GNDA.n1442 0.0682083
R20732 GNDA.n1453 GNDA.n1452 0.0682083
R20733 GNDA.n1461 GNDA.n1390 0.0682083
R20734 GNDA.n1471 GNDA.n1388 0.0682083
R20735 GNDA.n1473 GNDA.n1472 0.0682083
R20736 GNDA.n1483 GNDA.n1482 0.0682083
R20737 GNDA.n1491 GNDA.n1384 0.0682083
R20738 GNDA.n1501 GNDA.n1382 0.0682083
R20739 GNDA.n1503 GNDA.n1502 0.0682083
R20740 GNDA.n1240 GNDA.n1239 0.0682083
R20741 GNDA.n1250 GNDA.n1249 0.0682083
R20742 GNDA.n1258 GNDA.n1212 0.0682083
R20743 GNDA.n1268 GNDA.n1210 0.0682083
R20744 GNDA.n1270 GNDA.n1269 0.0682083
R20745 GNDA.n1280 GNDA.n1279 0.0682083
R20746 GNDA.n1288 GNDA.n1206 0.0682083
R20747 GNDA.n1298 GNDA.n1204 0.0682083
R20748 GNDA.n1300 GNDA.n1299 0.0682083
R20749 GNDA.n1310 GNDA.n1309 0.0682083
R20750 GNDA.n1318 GNDA.n1200 0.0682083
R20751 GNDA.n1328 GNDA.n1198 0.0682083
R20752 GNDA.n1330 GNDA.n1329 0.0682083
R20753 GNDA.n1340 GNDA.n1339 0.0682083
R20754 GNDA.n1347 GNDA.n1194 0.0682083
R20755 GNDA.n7141 GNDA.n7140 0.0682083
R20756 GNDA.n7147 GNDA.n7127 0.0682083
R20757 GNDA.n7155 GNDA.n7123 0.0682083
R20758 GNDA.n7157 GNDA.n7156 0.0682083
R20759 GNDA.n7165 GNDA.n7164 0.0682083
R20760 GNDA.n7171 GNDA.n7115 0.0682083
R20761 GNDA.n7179 GNDA.n7111 0.0682083
R20762 GNDA.n7181 GNDA.n7180 0.0682083
R20763 GNDA.n7189 GNDA.n7188 0.0682083
R20764 GNDA.n7195 GNDA.n7103 0.0682083
R20765 GNDA.n7203 GNDA.n7099 0.0682083
R20766 GNDA.n7205 GNDA.n7204 0.0682083
R20767 GNDA.n7213 GNDA.n7212 0.0682083
R20768 GNDA.n7219 GNDA.n7091 0.0682083
R20769 GNDA.n7228 GNDA.n95 0.0682083
R20770 GNDA.n7134 GNDA.n7132 0.0672139
R20771 GNDA.n5270 GNDA.n5137 0.0672139
R20772 GNDA.n4957 GNDA.n4824 0.0672139
R20773 GNDA.n4797 GNDA.n4659 0.0672139
R20774 GNDA.n4631 GNDA.n4493 0.0672139
R20775 GNDA.n4465 GNDA.n4327 0.0672139
R20776 GNDA.n4299 GNDA.n4161 0.0672139
R20777 GNDA.n3801 GNDA.n3485 0.0672139
R20778 GNDA.n4133 GNDA.n3995 0.0672139
R20779 GNDA.n3967 GNDA.n3829 0.0672139
R20780 GNDA.n3602 GNDA.n3557 0.0672139
R20781 GNDA.n496 GNDA.n451 0.0672139
R20782 GNDA.n5133 GNDA.n379 0.0672139
R20783 GNDA.n3299 GNDA.n3254 0.0672139
R20784 GNDA.n3195 GNDA.n3062 0.0672139
R20785 GNDA.n3035 GNDA.n2889 0.0672139
R20786 GNDA.n2399 GNDA.n691 0.0672139
R20787 GNDA.n2861 GNDA.n625 0.0672139
R20788 GNDA.n2662 GNDA.n2617 0.0672139
R20789 GNDA.n2559 GNDA.n2426 0.0672139
R20790 GNDA.n2202 GNDA.n2157 0.0672139
R20791 GNDA.n2096 GNDA.n1963 0.0672139
R20792 GNDA.n1936 GNDA.n754 0.0672139
R20793 GNDA.n1615 GNDA.n1570 0.0672139
R20794 GNDA.n1512 GNDA.n1379 0.0672139
R20795 GNDA.n1349 GNDA.n1193 0.0672139
R20796 GNDA.n149 GNDA.n148 0.0667303
R20797 GNDA.n7225 GNDA.n7065 0.0661531
R20798 GNDA.n5170 GNDA.n5169 0.063
R20799 GNDA.n5181 GNDA.n5154 0.063
R20800 GNDA.n5200 GNDA.n5199 0.063
R20801 GNDA.n5211 GNDA.n5148 0.063
R20802 GNDA.n5230 GNDA.n5229 0.063
R20803 GNDA.n5241 GNDA.n5142 0.063
R20804 GNDA.n5260 GNDA.n5259 0.063
R20805 GNDA.n4857 GNDA.n4856 0.063
R20806 GNDA.n4868 GNDA.n4841 0.063
R20807 GNDA.n4887 GNDA.n4886 0.063
R20808 GNDA.n4898 GNDA.n4835 0.063
R20809 GNDA.n4917 GNDA.n4916 0.063
R20810 GNDA.n4928 GNDA.n4829 0.063
R20811 GNDA.n4947 GNDA.n4946 0.063
R20812 GNDA.n4697 GNDA.n4696 0.063
R20813 GNDA.n4708 GNDA.n4676 0.063
R20814 GNDA.n4727 GNDA.n4726 0.063
R20815 GNDA.n4738 GNDA.n4670 0.063
R20816 GNDA.n4757 GNDA.n4756 0.063
R20817 GNDA.n4768 GNDA.n4664 0.063
R20818 GNDA.n4787 GNDA.n4786 0.063
R20819 GNDA.n4531 GNDA.n4530 0.063
R20820 GNDA.n4542 GNDA.n4510 0.063
R20821 GNDA.n4561 GNDA.n4560 0.063
R20822 GNDA.n4572 GNDA.n4504 0.063
R20823 GNDA.n4591 GNDA.n4590 0.063
R20824 GNDA.n4602 GNDA.n4498 0.063
R20825 GNDA.n4621 GNDA.n4620 0.063
R20826 GNDA.n4365 GNDA.n4364 0.063
R20827 GNDA.n4376 GNDA.n4344 0.063
R20828 GNDA.n4395 GNDA.n4394 0.063
R20829 GNDA.n4406 GNDA.n4338 0.063
R20830 GNDA.n4425 GNDA.n4424 0.063
R20831 GNDA.n4436 GNDA.n4332 0.063
R20832 GNDA.n4455 GNDA.n4454 0.063
R20833 GNDA.n4199 GNDA.n4198 0.063
R20834 GNDA.n4210 GNDA.n4178 0.063
R20835 GNDA.n4229 GNDA.n4228 0.063
R20836 GNDA.n4240 GNDA.n4172 0.063
R20837 GNDA.n4259 GNDA.n4258 0.063
R20838 GNDA.n4270 GNDA.n4166 0.063
R20839 GNDA.n4289 GNDA.n4288 0.063
R20840 GNDA.n3701 GNDA.n3700 0.063
R20841 GNDA.n3712 GNDA.n3502 0.063
R20842 GNDA.n3731 GNDA.n3730 0.063
R20843 GNDA.n3742 GNDA.n3496 0.063
R20844 GNDA.n3761 GNDA.n3760 0.063
R20845 GNDA.n3772 GNDA.n3490 0.063
R20846 GNDA.n3791 GNDA.n3790 0.063
R20847 GNDA.n4033 GNDA.n4032 0.063
R20848 GNDA.n4044 GNDA.n4012 0.063
R20849 GNDA.n4063 GNDA.n4062 0.063
R20850 GNDA.n4074 GNDA.n4006 0.063
R20851 GNDA.n4093 GNDA.n4092 0.063
R20852 GNDA.n4104 GNDA.n4000 0.063
R20853 GNDA.n4123 GNDA.n4122 0.063
R20854 GNDA.n3867 GNDA.n3866 0.063
R20855 GNDA.n3878 GNDA.n3846 0.063
R20856 GNDA.n3897 GNDA.n3896 0.063
R20857 GNDA.n3908 GNDA.n3840 0.063
R20858 GNDA.n3927 GNDA.n3926 0.063
R20859 GNDA.n3938 GNDA.n3834 0.063
R20860 GNDA.n3957 GNDA.n3956 0.063
R20861 GNDA.n3562 GNDA.n3561 0.063
R20862 GNDA.n3568 GNDA.n3567 0.063
R20863 GNDA.n3574 GNDA.n3573 0.063
R20864 GNDA.n3580 GNDA.n3579 0.063
R20865 GNDA.n3586 GNDA.n3585 0.063
R20866 GNDA.n3592 GNDA.n3591 0.063
R20867 GNDA.n3598 GNDA.n3597 0.063
R20868 GNDA.n456 GNDA.n455 0.063
R20869 GNDA.n462 GNDA.n461 0.063
R20870 GNDA.n468 GNDA.n467 0.063
R20871 GNDA.n474 GNDA.n473 0.063
R20872 GNDA.n480 GNDA.n479 0.063
R20873 GNDA.n486 GNDA.n485 0.063
R20874 GNDA.n492 GNDA.n491 0.063
R20875 GNDA.n5033 GNDA.n5032 0.063
R20876 GNDA.n5044 GNDA.n396 0.063
R20877 GNDA.n5063 GNDA.n5062 0.063
R20878 GNDA.n5074 GNDA.n390 0.063
R20879 GNDA.n5093 GNDA.n5092 0.063
R20880 GNDA.n5104 GNDA.n384 0.063
R20881 GNDA.n5123 GNDA.n5122 0.063
R20882 GNDA.n3259 GNDA.n3258 0.063
R20883 GNDA.n3265 GNDA.n3264 0.063
R20884 GNDA.n3271 GNDA.n3270 0.063
R20885 GNDA.n3277 GNDA.n3276 0.063
R20886 GNDA.n3283 GNDA.n3282 0.063
R20887 GNDA.n3289 GNDA.n3288 0.063
R20888 GNDA.n3295 GNDA.n3294 0.063
R20889 GNDA.n3095 GNDA.n3094 0.063
R20890 GNDA.n3106 GNDA.n3079 0.063
R20891 GNDA.n3125 GNDA.n3124 0.063
R20892 GNDA.n3136 GNDA.n3073 0.063
R20893 GNDA.n3155 GNDA.n3154 0.063
R20894 GNDA.n3166 GNDA.n3067 0.063
R20895 GNDA.n3185 GNDA.n3184 0.063
R20896 GNDA.n2935 GNDA.n2934 0.063
R20897 GNDA.n2946 GNDA.n2906 0.063
R20898 GNDA.n2965 GNDA.n2964 0.063
R20899 GNDA.n2976 GNDA.n2900 0.063
R20900 GNDA.n2995 GNDA.n2994 0.063
R20901 GNDA.n3006 GNDA.n2894 0.063
R20902 GNDA.n3025 GNDA.n3024 0.063
R20903 GNDA.n2299 GNDA.n2298 0.063
R20904 GNDA.n2310 GNDA.n708 0.063
R20905 GNDA.n2329 GNDA.n2328 0.063
R20906 GNDA.n2340 GNDA.n702 0.063
R20907 GNDA.n2359 GNDA.n2358 0.063
R20908 GNDA.n2370 GNDA.n696 0.063
R20909 GNDA.n2389 GNDA.n2388 0.063
R20910 GNDA.n2761 GNDA.n2760 0.063
R20911 GNDA.n2772 GNDA.n642 0.063
R20912 GNDA.n2791 GNDA.n2790 0.063
R20913 GNDA.n2802 GNDA.n636 0.063
R20914 GNDA.n2821 GNDA.n2820 0.063
R20915 GNDA.n2832 GNDA.n630 0.063
R20916 GNDA.n2851 GNDA.n2850 0.063
R20917 GNDA.n2622 GNDA.n2621 0.063
R20918 GNDA.n2628 GNDA.n2627 0.063
R20919 GNDA.n2634 GNDA.n2633 0.063
R20920 GNDA.n2640 GNDA.n2639 0.063
R20921 GNDA.n2646 GNDA.n2645 0.063
R20922 GNDA.n2652 GNDA.n2651 0.063
R20923 GNDA.n2658 GNDA.n2657 0.063
R20924 GNDA.n2459 GNDA.n2458 0.063
R20925 GNDA.n2470 GNDA.n2443 0.063
R20926 GNDA.n2489 GNDA.n2488 0.063
R20927 GNDA.n2500 GNDA.n2437 0.063
R20928 GNDA.n2519 GNDA.n2518 0.063
R20929 GNDA.n2530 GNDA.n2431 0.063
R20930 GNDA.n2549 GNDA.n2548 0.063
R20931 GNDA.n2162 GNDA.n2161 0.063
R20932 GNDA.n2168 GNDA.n2167 0.063
R20933 GNDA.n2174 GNDA.n2173 0.063
R20934 GNDA.n2180 GNDA.n2179 0.063
R20935 GNDA.n2186 GNDA.n2185 0.063
R20936 GNDA.n2192 GNDA.n2191 0.063
R20937 GNDA.n2198 GNDA.n2197 0.063
R20938 GNDA.n1996 GNDA.n1995 0.063
R20939 GNDA.n2007 GNDA.n1980 0.063
R20940 GNDA.n2026 GNDA.n2025 0.063
R20941 GNDA.n2037 GNDA.n1974 0.063
R20942 GNDA.n2056 GNDA.n2055 0.063
R20943 GNDA.n2067 GNDA.n1968 0.063
R20944 GNDA.n2086 GNDA.n2085 0.063
R20945 GNDA.n1836 GNDA.n1835 0.063
R20946 GNDA.n1847 GNDA.n771 0.063
R20947 GNDA.n1866 GNDA.n1865 0.063
R20948 GNDA.n1877 GNDA.n765 0.063
R20949 GNDA.n1896 GNDA.n1895 0.063
R20950 GNDA.n1907 GNDA.n759 0.063
R20951 GNDA.n1926 GNDA.n1925 0.063
R20952 GNDA.n1575 GNDA.n1574 0.063
R20953 GNDA.n1581 GNDA.n1580 0.063
R20954 GNDA.n1587 GNDA.n1586 0.063
R20955 GNDA.n1593 GNDA.n1592 0.063
R20956 GNDA.n1599 GNDA.n1598 0.063
R20957 GNDA.n1605 GNDA.n1604 0.063
R20958 GNDA.n1611 GNDA.n1610 0.063
R20959 GNDA.n1412 GNDA.n1411 0.063
R20960 GNDA.n1423 GNDA.n1396 0.063
R20961 GNDA.n1442 GNDA.n1441 0.063
R20962 GNDA.n1453 GNDA.n1390 0.063
R20963 GNDA.n1472 GNDA.n1471 0.063
R20964 GNDA.n1483 GNDA.n1384 0.063
R20965 GNDA.n1502 GNDA.n1501 0.063
R20966 GNDA.n1250 GNDA.n1212 0.063
R20967 GNDA.n1269 GNDA.n1268 0.063
R20968 GNDA.n1280 GNDA.n1206 0.063
R20969 GNDA.n1299 GNDA.n1298 0.063
R20970 GNDA.n1310 GNDA.n1200 0.063
R20971 GNDA.n1329 GNDA.n1328 0.063
R20972 GNDA.n1340 GNDA.n1194 0.063
R20973 GNDA.n3376 GNDA.n324 0.063
R20974 GNDA.n7141 GNDA.n7127 0.063
R20975 GNDA.n7156 GNDA.n7155 0.063
R20976 GNDA.n7165 GNDA.n7115 0.063
R20977 GNDA.n7180 GNDA.n7179 0.063
R20978 GNDA.n7189 GNDA.n7103 0.063
R20979 GNDA.n7204 GNDA.n7203 0.063
R20980 GNDA.n7213 GNDA.n7091 0.063
R20981 GNDA.n7049 GNDA.n7048 0.063
R20982 GNDA.n2282 GNDA.n2281 0.0629369
R20983 GNDA.n3679 GNDA.n573 0.0629369
R20984 GNDA.n5359 GNDA.n5358 0.0626438
R20985 GNDA.n6951 GNDA.n5351 0.0626438
R20986 GNDA.n649 GNDA.n320 0.0577917
R20987 GNDA.n5163 GNDA.n5162 0.0553333
R20988 GNDA.n5177 GNDA.n5176 0.0553333
R20989 GNDA.n5193 GNDA.n5192 0.0553333
R20990 GNDA.n5207 GNDA.n5206 0.0553333
R20991 GNDA.n5223 GNDA.n5222 0.0553333
R20992 GNDA.n5237 GNDA.n5236 0.0553333
R20993 GNDA.n5253 GNDA.n5252 0.0553333
R20994 GNDA.n5267 GNDA.n5266 0.0553333
R20995 GNDA.n4850 GNDA.n4849 0.0553333
R20996 GNDA.n4864 GNDA.n4863 0.0553333
R20997 GNDA.n4880 GNDA.n4879 0.0553333
R20998 GNDA.n4894 GNDA.n4893 0.0553333
R20999 GNDA.n4910 GNDA.n4909 0.0553333
R21000 GNDA.n4924 GNDA.n4923 0.0553333
R21001 GNDA.n4940 GNDA.n4939 0.0553333
R21002 GNDA.n4954 GNDA.n4953 0.0553333
R21003 GNDA.n4690 GNDA.n4689 0.0553333
R21004 GNDA.n4704 GNDA.n4703 0.0553333
R21005 GNDA.n4720 GNDA.n4719 0.0553333
R21006 GNDA.n4734 GNDA.n4733 0.0553333
R21007 GNDA.n4750 GNDA.n4749 0.0553333
R21008 GNDA.n4764 GNDA.n4763 0.0553333
R21009 GNDA.n4780 GNDA.n4779 0.0553333
R21010 GNDA.n4794 GNDA.n4793 0.0553333
R21011 GNDA.n4524 GNDA.n4523 0.0553333
R21012 GNDA.n4538 GNDA.n4537 0.0553333
R21013 GNDA.n4554 GNDA.n4553 0.0553333
R21014 GNDA.n4568 GNDA.n4567 0.0553333
R21015 GNDA.n4584 GNDA.n4583 0.0553333
R21016 GNDA.n4598 GNDA.n4597 0.0553333
R21017 GNDA.n4614 GNDA.n4613 0.0553333
R21018 GNDA.n4628 GNDA.n4627 0.0553333
R21019 GNDA.n4358 GNDA.n4357 0.0553333
R21020 GNDA.n4372 GNDA.n4371 0.0553333
R21021 GNDA.n4388 GNDA.n4387 0.0553333
R21022 GNDA.n4402 GNDA.n4401 0.0553333
R21023 GNDA.n4418 GNDA.n4417 0.0553333
R21024 GNDA.n4432 GNDA.n4431 0.0553333
R21025 GNDA.n4448 GNDA.n4447 0.0553333
R21026 GNDA.n4462 GNDA.n4461 0.0553333
R21027 GNDA.n4192 GNDA.n4191 0.0553333
R21028 GNDA.n4206 GNDA.n4205 0.0553333
R21029 GNDA.n4222 GNDA.n4221 0.0553333
R21030 GNDA.n4236 GNDA.n4235 0.0553333
R21031 GNDA.n4252 GNDA.n4251 0.0553333
R21032 GNDA.n4266 GNDA.n4265 0.0553333
R21033 GNDA.n4282 GNDA.n4281 0.0553333
R21034 GNDA.n4296 GNDA.n4295 0.0553333
R21035 GNDA.n3694 GNDA.n3693 0.0553333
R21036 GNDA.n3708 GNDA.n3707 0.0553333
R21037 GNDA.n3724 GNDA.n3723 0.0553333
R21038 GNDA.n3738 GNDA.n3737 0.0553333
R21039 GNDA.n3754 GNDA.n3753 0.0553333
R21040 GNDA.n3768 GNDA.n3767 0.0553333
R21041 GNDA.n3784 GNDA.n3783 0.0553333
R21042 GNDA.n3798 GNDA.n3797 0.0553333
R21043 GNDA.n4026 GNDA.n4025 0.0553333
R21044 GNDA.n4040 GNDA.n4039 0.0553333
R21045 GNDA.n4056 GNDA.n4055 0.0553333
R21046 GNDA.n4070 GNDA.n4069 0.0553333
R21047 GNDA.n4086 GNDA.n4085 0.0553333
R21048 GNDA.n4100 GNDA.n4099 0.0553333
R21049 GNDA.n4116 GNDA.n4115 0.0553333
R21050 GNDA.n4130 GNDA.n4129 0.0553333
R21051 GNDA.n3860 GNDA.n3859 0.0553333
R21052 GNDA.n3874 GNDA.n3873 0.0553333
R21053 GNDA.n3890 GNDA.n3889 0.0553333
R21054 GNDA.n3904 GNDA.n3903 0.0553333
R21055 GNDA.n3920 GNDA.n3919 0.0553333
R21056 GNDA.n3934 GNDA.n3933 0.0553333
R21057 GNDA.n3950 GNDA.n3949 0.0553333
R21058 GNDA.n3964 GNDA.n3963 0.0553333
R21059 GNDA.n3670 GNDA.n3669 0.0553333
R21060 GNDA.n3661 GNDA.n3660 0.0553333
R21061 GNDA.n3652 GNDA.n3651 0.0553333
R21062 GNDA.n3643 GNDA.n3642 0.0553333
R21063 GNDA.n3634 GNDA.n3633 0.0553333
R21064 GNDA.n3625 GNDA.n3624 0.0553333
R21065 GNDA.n3616 GNDA.n3615 0.0553333
R21066 GNDA.n3607 GNDA.n3606 0.0553333
R21067 GNDA.n564 GNDA.n563 0.0553333
R21068 GNDA.n555 GNDA.n554 0.0553333
R21069 GNDA.n546 GNDA.n545 0.0553333
R21070 GNDA.n537 GNDA.n536 0.0553333
R21071 GNDA.n528 GNDA.n527 0.0553333
R21072 GNDA.n519 GNDA.n518 0.0553333
R21073 GNDA.n510 GNDA.n509 0.0553333
R21074 GNDA.n501 GNDA.n500 0.0553333
R21075 GNDA.n5026 GNDA.n5025 0.0553333
R21076 GNDA.n5040 GNDA.n5039 0.0553333
R21077 GNDA.n5056 GNDA.n5055 0.0553333
R21078 GNDA.n5070 GNDA.n5069 0.0553333
R21079 GNDA.n5086 GNDA.n5085 0.0553333
R21080 GNDA.n5100 GNDA.n5099 0.0553333
R21081 GNDA.n5116 GNDA.n5115 0.0553333
R21082 GNDA.n5130 GNDA.n5129 0.0553333
R21083 GNDA.n3367 GNDA.n3366 0.0553333
R21084 GNDA.n3358 GNDA.n3357 0.0553333
R21085 GNDA.n3349 GNDA.n3348 0.0553333
R21086 GNDA.n3340 GNDA.n3339 0.0553333
R21087 GNDA.n3331 GNDA.n3330 0.0553333
R21088 GNDA.n3322 GNDA.n3321 0.0553333
R21089 GNDA.n3313 GNDA.n3312 0.0553333
R21090 GNDA.n3304 GNDA.n3303 0.0553333
R21091 GNDA.n3088 GNDA.n3087 0.0553333
R21092 GNDA.n3102 GNDA.n3101 0.0553333
R21093 GNDA.n3118 GNDA.n3117 0.0553333
R21094 GNDA.n3132 GNDA.n3131 0.0553333
R21095 GNDA.n3148 GNDA.n3147 0.0553333
R21096 GNDA.n3162 GNDA.n3161 0.0553333
R21097 GNDA.n3178 GNDA.n3177 0.0553333
R21098 GNDA.n3192 GNDA.n3191 0.0553333
R21099 GNDA.n2928 GNDA.n2927 0.0553333
R21100 GNDA.n2942 GNDA.n2941 0.0553333
R21101 GNDA.n2958 GNDA.n2957 0.0553333
R21102 GNDA.n2972 GNDA.n2971 0.0553333
R21103 GNDA.n2988 GNDA.n2987 0.0553333
R21104 GNDA.n3002 GNDA.n3001 0.0553333
R21105 GNDA.n3018 GNDA.n3017 0.0553333
R21106 GNDA.n3032 GNDA.n3031 0.0553333
R21107 GNDA.n2292 GNDA.n2291 0.0553333
R21108 GNDA.n2306 GNDA.n2305 0.0553333
R21109 GNDA.n2322 GNDA.n2321 0.0553333
R21110 GNDA.n2336 GNDA.n2335 0.0553333
R21111 GNDA.n2352 GNDA.n2351 0.0553333
R21112 GNDA.n2366 GNDA.n2365 0.0553333
R21113 GNDA.n2382 GNDA.n2381 0.0553333
R21114 GNDA.n2396 GNDA.n2395 0.0553333
R21115 GNDA.n2754 GNDA.n2753 0.0553333
R21116 GNDA.n2768 GNDA.n2767 0.0553333
R21117 GNDA.n2784 GNDA.n2783 0.0553333
R21118 GNDA.n2798 GNDA.n2797 0.0553333
R21119 GNDA.n2814 GNDA.n2813 0.0553333
R21120 GNDA.n2828 GNDA.n2827 0.0553333
R21121 GNDA.n2844 GNDA.n2843 0.0553333
R21122 GNDA.n2858 GNDA.n2857 0.0553333
R21123 GNDA.n2730 GNDA.n2729 0.0553333
R21124 GNDA.n2721 GNDA.n2720 0.0553333
R21125 GNDA.n2712 GNDA.n2711 0.0553333
R21126 GNDA.n2703 GNDA.n2702 0.0553333
R21127 GNDA.n2694 GNDA.n2693 0.0553333
R21128 GNDA.n2685 GNDA.n2684 0.0553333
R21129 GNDA.n2676 GNDA.n2675 0.0553333
R21130 GNDA.n2667 GNDA.n2666 0.0553333
R21131 GNDA.n2452 GNDA.n2451 0.0553333
R21132 GNDA.n2466 GNDA.n2465 0.0553333
R21133 GNDA.n2482 GNDA.n2481 0.0553333
R21134 GNDA.n2496 GNDA.n2495 0.0553333
R21135 GNDA.n2512 GNDA.n2511 0.0553333
R21136 GNDA.n2526 GNDA.n2525 0.0553333
R21137 GNDA.n2542 GNDA.n2541 0.0553333
R21138 GNDA.n2556 GNDA.n2555 0.0553333
R21139 GNDA.n2270 GNDA.n2269 0.0553333
R21140 GNDA.n2261 GNDA.n2260 0.0553333
R21141 GNDA.n2252 GNDA.n2251 0.0553333
R21142 GNDA.n2243 GNDA.n2242 0.0553333
R21143 GNDA.n2234 GNDA.n2233 0.0553333
R21144 GNDA.n2225 GNDA.n2224 0.0553333
R21145 GNDA.n2216 GNDA.n2215 0.0553333
R21146 GNDA.n2207 GNDA.n2206 0.0553333
R21147 GNDA.n1989 GNDA.n1988 0.0553333
R21148 GNDA.n2003 GNDA.n2002 0.0553333
R21149 GNDA.n2019 GNDA.n2018 0.0553333
R21150 GNDA.n2033 GNDA.n2032 0.0553333
R21151 GNDA.n2049 GNDA.n2048 0.0553333
R21152 GNDA.n2063 GNDA.n2062 0.0553333
R21153 GNDA.n2079 GNDA.n2078 0.0553333
R21154 GNDA.n2093 GNDA.n2092 0.0553333
R21155 GNDA.n1829 GNDA.n1828 0.0553333
R21156 GNDA.n1843 GNDA.n1842 0.0553333
R21157 GNDA.n1859 GNDA.n1858 0.0553333
R21158 GNDA.n1873 GNDA.n1872 0.0553333
R21159 GNDA.n1889 GNDA.n1888 0.0553333
R21160 GNDA.n1903 GNDA.n1902 0.0553333
R21161 GNDA.n1919 GNDA.n1918 0.0553333
R21162 GNDA.n1933 GNDA.n1932 0.0553333
R21163 GNDA.n1683 GNDA.n1682 0.0553333
R21164 GNDA.n1674 GNDA.n1673 0.0553333
R21165 GNDA.n1665 GNDA.n1664 0.0553333
R21166 GNDA.n1656 GNDA.n1655 0.0553333
R21167 GNDA.n1647 GNDA.n1646 0.0553333
R21168 GNDA.n1638 GNDA.n1637 0.0553333
R21169 GNDA.n1629 GNDA.n1628 0.0553333
R21170 GNDA.n1620 GNDA.n1619 0.0553333
R21171 GNDA.n1405 GNDA.n1404 0.0553333
R21172 GNDA.n1419 GNDA.n1418 0.0553333
R21173 GNDA.n1435 GNDA.n1434 0.0553333
R21174 GNDA.n1449 GNDA.n1448 0.0553333
R21175 GNDA.n1465 GNDA.n1464 0.0553333
R21176 GNDA.n1479 GNDA.n1478 0.0553333
R21177 GNDA.n1495 GNDA.n1494 0.0553333
R21178 GNDA.n1509 GNDA.n1508 0.0553333
R21179 GNDA.n1243 GNDA.n1242 0.0553333
R21180 GNDA.n1246 GNDA.n1245 0.0553333
R21181 GNDA.n1256 GNDA.n1255 0.0553333
R21182 GNDA.n1263 GNDA.n1262 0.0553333
R21183 GNDA.n1273 GNDA.n1272 0.0553333
R21184 GNDA.n1276 GNDA.n1275 0.0553333
R21185 GNDA.n1286 GNDA.n1285 0.0553333
R21186 GNDA.n1293 GNDA.n1292 0.0553333
R21187 GNDA.n1303 GNDA.n1302 0.0553333
R21188 GNDA.n1306 GNDA.n1305 0.0553333
R21189 GNDA.n1316 GNDA.n1315 0.0553333
R21190 GNDA.n1323 GNDA.n1322 0.0553333
R21191 GNDA.n1333 GNDA.n1332 0.0553333
R21192 GNDA.n1336 GNDA.n1335 0.0553333
R21193 GNDA.n1345 GNDA.n1190 0.0553333
R21194 GNDA.n1352 GNDA.n1191 0.0553333
R21195 GNDA.n7137 GNDA.n7136 0.0553333
R21196 GNDA.n7126 GNDA.n7125 0.0553333
R21197 GNDA.n7161 GNDA.n7160 0.0553333
R21198 GNDA.n7114 GNDA.n7113 0.0553333
R21199 GNDA.n7185 GNDA.n7184 0.0553333
R21200 GNDA.n7102 GNDA.n7101 0.0553333
R21201 GNDA.n7209 GNDA.n7208 0.0553333
R21202 GNDA.n7223 GNDA.n7089 0.0553333
R21203 GNDA.n153 GNDA.n152 0.0553333
R21204 GNDA.n167 GNDA.n166 0.0553333
R21205 GNDA.n183 GNDA.n182 0.0553333
R21206 GNDA.n197 GNDA.n196 0.0553333
R21207 GNDA.n213 GNDA.n212 0.0553333
R21208 GNDA.n227 GNDA.n226 0.0553333
R21209 GNDA.n243 GNDA.n242 0.0553333
R21210 GNDA.n257 GNDA.n256 0.0553333
R21211 GNDA.n6364 GNDA 0.0517
R21212 GNDA.n6465 GNDA 0.0517
R21213 GNDA.n6980 GNDA 0.0517
R21214 GNDA GNDA.n6800 0.0517
R21215 GNDA.n5728 GNDA 0.0517
R21216 GNDA GNDA.n5490 0.0517
R21217 GNDA GNDA.n5915 0.0517
R21218 GNDA.n6758 GNDA 0.0517
R21219 GNDA GNDA.n0 0.0517
R21220 GNDA.n5273 GNDA.n328 0.0514167
R21221 GNDA.n5167 GNDA.n5166 0.0514167
R21222 GNDA.n5173 GNDA.n5172 0.0514167
R21223 GNDA.n5183 GNDA.n5182 0.0514167
R21224 GNDA.n5187 GNDA.n5186 0.0514167
R21225 GNDA.n5197 GNDA.n5196 0.0514167
R21226 GNDA.n5203 GNDA.n5202 0.0514167
R21227 GNDA.n5213 GNDA.n5212 0.0514167
R21228 GNDA.n5217 GNDA.n5216 0.0514167
R21229 GNDA.n5227 GNDA.n5226 0.0514167
R21230 GNDA.n5233 GNDA.n5232 0.0514167
R21231 GNDA.n5243 GNDA.n5242 0.0514167
R21232 GNDA.n5247 GNDA.n5246 0.0514167
R21233 GNDA.n5257 GNDA.n5256 0.0514167
R21234 GNDA.n5263 GNDA.n5262 0.0514167
R21235 GNDA.n5271 GNDA.n5136 0.0514167
R21236 GNDA.n4960 GNDA.n3458 0.0514167
R21237 GNDA.n4854 GNDA.n4853 0.0514167
R21238 GNDA.n4860 GNDA.n4859 0.0514167
R21239 GNDA.n4870 GNDA.n4869 0.0514167
R21240 GNDA.n4874 GNDA.n4873 0.0514167
R21241 GNDA.n4884 GNDA.n4883 0.0514167
R21242 GNDA.n4890 GNDA.n4889 0.0514167
R21243 GNDA.n4900 GNDA.n4899 0.0514167
R21244 GNDA.n4904 GNDA.n4903 0.0514167
R21245 GNDA.n4914 GNDA.n4913 0.0514167
R21246 GNDA.n4920 GNDA.n4919 0.0514167
R21247 GNDA.n4930 GNDA.n4929 0.0514167
R21248 GNDA.n4934 GNDA.n4933 0.0514167
R21249 GNDA.n4944 GNDA.n4943 0.0514167
R21250 GNDA.n4950 GNDA.n4949 0.0514167
R21251 GNDA.n4958 GNDA.n4823 0.0514167
R21252 GNDA.n4684 GNDA.n4634 0.0514167
R21253 GNDA.n4694 GNDA.n4693 0.0514167
R21254 GNDA.n4700 GNDA.n4699 0.0514167
R21255 GNDA.n4710 GNDA.n4709 0.0514167
R21256 GNDA.n4714 GNDA.n4713 0.0514167
R21257 GNDA.n4724 GNDA.n4723 0.0514167
R21258 GNDA.n4730 GNDA.n4729 0.0514167
R21259 GNDA.n4740 GNDA.n4739 0.0514167
R21260 GNDA.n4744 GNDA.n4743 0.0514167
R21261 GNDA.n4754 GNDA.n4753 0.0514167
R21262 GNDA.n4760 GNDA.n4759 0.0514167
R21263 GNDA.n4770 GNDA.n4769 0.0514167
R21264 GNDA.n4774 GNDA.n4773 0.0514167
R21265 GNDA.n4784 GNDA.n4783 0.0514167
R21266 GNDA.n4790 GNDA.n4789 0.0514167
R21267 GNDA.n4798 GNDA.n4658 0.0514167
R21268 GNDA.n4518 GNDA.n4468 0.0514167
R21269 GNDA.n4528 GNDA.n4527 0.0514167
R21270 GNDA.n4534 GNDA.n4533 0.0514167
R21271 GNDA.n4544 GNDA.n4543 0.0514167
R21272 GNDA.n4548 GNDA.n4547 0.0514167
R21273 GNDA.n4558 GNDA.n4557 0.0514167
R21274 GNDA.n4564 GNDA.n4563 0.0514167
R21275 GNDA.n4574 GNDA.n4573 0.0514167
R21276 GNDA.n4578 GNDA.n4577 0.0514167
R21277 GNDA.n4588 GNDA.n4587 0.0514167
R21278 GNDA.n4594 GNDA.n4593 0.0514167
R21279 GNDA.n4604 GNDA.n4603 0.0514167
R21280 GNDA.n4608 GNDA.n4607 0.0514167
R21281 GNDA.n4618 GNDA.n4617 0.0514167
R21282 GNDA.n4624 GNDA.n4623 0.0514167
R21283 GNDA.n4632 GNDA.n4492 0.0514167
R21284 GNDA.n4352 GNDA.n4302 0.0514167
R21285 GNDA.n4362 GNDA.n4361 0.0514167
R21286 GNDA.n4368 GNDA.n4367 0.0514167
R21287 GNDA.n4378 GNDA.n4377 0.0514167
R21288 GNDA.n4382 GNDA.n4381 0.0514167
R21289 GNDA.n4392 GNDA.n4391 0.0514167
R21290 GNDA.n4398 GNDA.n4397 0.0514167
R21291 GNDA.n4408 GNDA.n4407 0.0514167
R21292 GNDA.n4412 GNDA.n4411 0.0514167
R21293 GNDA.n4422 GNDA.n4421 0.0514167
R21294 GNDA.n4428 GNDA.n4427 0.0514167
R21295 GNDA.n4438 GNDA.n4437 0.0514167
R21296 GNDA.n4442 GNDA.n4441 0.0514167
R21297 GNDA.n4452 GNDA.n4451 0.0514167
R21298 GNDA.n4458 GNDA.n4457 0.0514167
R21299 GNDA.n4466 GNDA.n4326 0.0514167
R21300 GNDA.n4186 GNDA.n4136 0.0514167
R21301 GNDA.n4196 GNDA.n4195 0.0514167
R21302 GNDA.n4202 GNDA.n4201 0.0514167
R21303 GNDA.n4212 GNDA.n4211 0.0514167
R21304 GNDA.n4216 GNDA.n4215 0.0514167
R21305 GNDA.n4226 GNDA.n4225 0.0514167
R21306 GNDA.n4232 GNDA.n4231 0.0514167
R21307 GNDA.n4242 GNDA.n4241 0.0514167
R21308 GNDA.n4246 GNDA.n4245 0.0514167
R21309 GNDA.n4256 GNDA.n4255 0.0514167
R21310 GNDA.n4262 GNDA.n4261 0.0514167
R21311 GNDA.n4272 GNDA.n4271 0.0514167
R21312 GNDA.n4276 GNDA.n4275 0.0514167
R21313 GNDA.n4286 GNDA.n4285 0.0514167
R21314 GNDA.n4292 GNDA.n4291 0.0514167
R21315 GNDA.n4300 GNDA.n4160 0.0514167
R21316 GNDA.n3688 GNDA.n3460 0.0514167
R21317 GNDA.n3698 GNDA.n3697 0.0514167
R21318 GNDA.n3704 GNDA.n3703 0.0514167
R21319 GNDA.n3714 GNDA.n3713 0.0514167
R21320 GNDA.n3718 GNDA.n3717 0.0514167
R21321 GNDA.n3728 GNDA.n3727 0.0514167
R21322 GNDA.n3734 GNDA.n3733 0.0514167
R21323 GNDA.n3744 GNDA.n3743 0.0514167
R21324 GNDA.n3748 GNDA.n3747 0.0514167
R21325 GNDA.n3758 GNDA.n3757 0.0514167
R21326 GNDA.n3764 GNDA.n3763 0.0514167
R21327 GNDA.n3774 GNDA.n3773 0.0514167
R21328 GNDA.n3778 GNDA.n3777 0.0514167
R21329 GNDA.n3788 GNDA.n3787 0.0514167
R21330 GNDA.n3794 GNDA.n3793 0.0514167
R21331 GNDA.n3802 GNDA.n3484 0.0514167
R21332 GNDA.n4020 GNDA.n3970 0.0514167
R21333 GNDA.n4030 GNDA.n4029 0.0514167
R21334 GNDA.n4036 GNDA.n4035 0.0514167
R21335 GNDA.n4046 GNDA.n4045 0.0514167
R21336 GNDA.n4050 GNDA.n4049 0.0514167
R21337 GNDA.n4060 GNDA.n4059 0.0514167
R21338 GNDA.n4066 GNDA.n4065 0.0514167
R21339 GNDA.n4076 GNDA.n4075 0.0514167
R21340 GNDA.n4080 GNDA.n4079 0.0514167
R21341 GNDA.n4090 GNDA.n4089 0.0514167
R21342 GNDA.n4096 GNDA.n4095 0.0514167
R21343 GNDA.n4106 GNDA.n4105 0.0514167
R21344 GNDA.n4110 GNDA.n4109 0.0514167
R21345 GNDA.n4120 GNDA.n4119 0.0514167
R21346 GNDA.n4126 GNDA.n4125 0.0514167
R21347 GNDA.n4134 GNDA.n3994 0.0514167
R21348 GNDA.n3854 GNDA.n3804 0.0514167
R21349 GNDA.n3864 GNDA.n3863 0.0514167
R21350 GNDA.n3870 GNDA.n3869 0.0514167
R21351 GNDA.n3880 GNDA.n3879 0.0514167
R21352 GNDA.n3884 GNDA.n3883 0.0514167
R21353 GNDA.n3894 GNDA.n3893 0.0514167
R21354 GNDA.n3900 GNDA.n3899 0.0514167
R21355 GNDA.n3910 GNDA.n3909 0.0514167
R21356 GNDA.n3914 GNDA.n3913 0.0514167
R21357 GNDA.n3924 GNDA.n3923 0.0514167
R21358 GNDA.n3930 GNDA.n3929 0.0514167
R21359 GNDA.n3940 GNDA.n3939 0.0514167
R21360 GNDA.n3944 GNDA.n3943 0.0514167
R21361 GNDA.n3954 GNDA.n3953 0.0514167
R21362 GNDA.n3960 GNDA.n3959 0.0514167
R21363 GNDA.n3968 GNDA.n3828 0.0514167
R21364 GNDA.n3673 GNDA.n3672 0.0514167
R21365 GNDA.n3667 GNDA.n3666 0.0514167
R21366 GNDA.n3664 GNDA.n3663 0.0514167
R21367 GNDA.n3658 GNDA.n3657 0.0514167
R21368 GNDA.n3655 GNDA.n3654 0.0514167
R21369 GNDA.n3649 GNDA.n3648 0.0514167
R21370 GNDA.n3646 GNDA.n3645 0.0514167
R21371 GNDA.n3640 GNDA.n3639 0.0514167
R21372 GNDA.n3637 GNDA.n3636 0.0514167
R21373 GNDA.n3631 GNDA.n3630 0.0514167
R21374 GNDA.n3628 GNDA.n3627 0.0514167
R21375 GNDA.n3622 GNDA.n3621 0.0514167
R21376 GNDA.n3619 GNDA.n3618 0.0514167
R21377 GNDA.n3613 GNDA.n3612 0.0514167
R21378 GNDA.n3610 GNDA.n3609 0.0514167
R21379 GNDA.n3604 GNDA.n3603 0.0514167
R21380 GNDA.n567 GNDA.n566 0.0514167
R21381 GNDA.n561 GNDA.n560 0.0514167
R21382 GNDA.n558 GNDA.n557 0.0514167
R21383 GNDA.n552 GNDA.n551 0.0514167
R21384 GNDA.n549 GNDA.n548 0.0514167
R21385 GNDA.n543 GNDA.n542 0.0514167
R21386 GNDA.n540 GNDA.n539 0.0514167
R21387 GNDA.n534 GNDA.n533 0.0514167
R21388 GNDA.n531 GNDA.n530 0.0514167
R21389 GNDA.n525 GNDA.n524 0.0514167
R21390 GNDA.n522 GNDA.n521 0.0514167
R21391 GNDA.n516 GNDA.n515 0.0514167
R21392 GNDA.n513 GNDA.n512 0.0514167
R21393 GNDA.n507 GNDA.n506 0.0514167
R21394 GNDA.n504 GNDA.n503 0.0514167
R21395 GNDA.n498 GNDA.n497 0.0514167
R21396 GNDA.n5020 GNDA.n353 0.0514167
R21397 GNDA.n5030 GNDA.n5029 0.0514167
R21398 GNDA.n5036 GNDA.n5035 0.0514167
R21399 GNDA.n5046 GNDA.n5045 0.0514167
R21400 GNDA.n5050 GNDA.n5049 0.0514167
R21401 GNDA.n5060 GNDA.n5059 0.0514167
R21402 GNDA.n5066 GNDA.n5065 0.0514167
R21403 GNDA.n5076 GNDA.n5075 0.0514167
R21404 GNDA.n5080 GNDA.n5079 0.0514167
R21405 GNDA.n5090 GNDA.n5089 0.0514167
R21406 GNDA.n5096 GNDA.n5095 0.0514167
R21407 GNDA.n5106 GNDA.n5105 0.0514167
R21408 GNDA.n5110 GNDA.n5109 0.0514167
R21409 GNDA.n5120 GNDA.n5119 0.0514167
R21410 GNDA.n5126 GNDA.n5125 0.0514167
R21411 GNDA.n5134 GNDA.n378 0.0514167
R21412 GNDA.n3370 GNDA.n3369 0.0514167
R21413 GNDA.n3364 GNDA.n3363 0.0514167
R21414 GNDA.n3361 GNDA.n3360 0.0514167
R21415 GNDA.n3355 GNDA.n3354 0.0514167
R21416 GNDA.n3352 GNDA.n3351 0.0514167
R21417 GNDA.n3346 GNDA.n3345 0.0514167
R21418 GNDA.n3343 GNDA.n3342 0.0514167
R21419 GNDA.n3337 GNDA.n3336 0.0514167
R21420 GNDA.n3334 GNDA.n3333 0.0514167
R21421 GNDA.n3328 GNDA.n3327 0.0514167
R21422 GNDA.n3325 GNDA.n3324 0.0514167
R21423 GNDA.n3319 GNDA.n3318 0.0514167
R21424 GNDA.n3316 GNDA.n3315 0.0514167
R21425 GNDA.n3310 GNDA.n3309 0.0514167
R21426 GNDA.n3307 GNDA.n3306 0.0514167
R21427 GNDA.n3301 GNDA.n3300 0.0514167
R21428 GNDA.n3198 GNDA.n598 0.0514167
R21429 GNDA.n3092 GNDA.n3091 0.0514167
R21430 GNDA.n3098 GNDA.n3097 0.0514167
R21431 GNDA.n3108 GNDA.n3107 0.0514167
R21432 GNDA.n3112 GNDA.n3111 0.0514167
R21433 GNDA.n3122 GNDA.n3121 0.0514167
R21434 GNDA.n3128 GNDA.n3127 0.0514167
R21435 GNDA.n3138 GNDA.n3137 0.0514167
R21436 GNDA.n3142 GNDA.n3141 0.0514167
R21437 GNDA.n3152 GNDA.n3151 0.0514167
R21438 GNDA.n3158 GNDA.n3157 0.0514167
R21439 GNDA.n3168 GNDA.n3167 0.0514167
R21440 GNDA.n3172 GNDA.n3171 0.0514167
R21441 GNDA.n3182 GNDA.n3181 0.0514167
R21442 GNDA.n3188 GNDA.n3187 0.0514167
R21443 GNDA.n3196 GNDA.n3061 0.0514167
R21444 GNDA.n2922 GNDA.n2864 0.0514167
R21445 GNDA.n2932 GNDA.n2931 0.0514167
R21446 GNDA.n2938 GNDA.n2937 0.0514167
R21447 GNDA.n2948 GNDA.n2947 0.0514167
R21448 GNDA.n2952 GNDA.n2951 0.0514167
R21449 GNDA.n2962 GNDA.n2961 0.0514167
R21450 GNDA.n2968 GNDA.n2967 0.0514167
R21451 GNDA.n2978 GNDA.n2977 0.0514167
R21452 GNDA.n2982 GNDA.n2981 0.0514167
R21453 GNDA.n2992 GNDA.n2991 0.0514167
R21454 GNDA.n2998 GNDA.n2997 0.0514167
R21455 GNDA.n3008 GNDA.n3007 0.0514167
R21456 GNDA.n3012 GNDA.n3011 0.0514167
R21457 GNDA.n3022 GNDA.n3021 0.0514167
R21458 GNDA.n3028 GNDA.n3027 0.0514167
R21459 GNDA.n3036 GNDA.n2888 0.0514167
R21460 GNDA.n2286 GNDA.n666 0.0514167
R21461 GNDA.n2296 GNDA.n2295 0.0514167
R21462 GNDA.n2302 GNDA.n2301 0.0514167
R21463 GNDA.n2312 GNDA.n2311 0.0514167
R21464 GNDA.n2316 GNDA.n2315 0.0514167
R21465 GNDA.n2326 GNDA.n2325 0.0514167
R21466 GNDA.n2332 GNDA.n2331 0.0514167
R21467 GNDA.n2342 GNDA.n2341 0.0514167
R21468 GNDA.n2346 GNDA.n2345 0.0514167
R21469 GNDA.n2356 GNDA.n2355 0.0514167
R21470 GNDA.n2362 GNDA.n2361 0.0514167
R21471 GNDA.n2372 GNDA.n2371 0.0514167
R21472 GNDA.n2376 GNDA.n2375 0.0514167
R21473 GNDA.n2386 GNDA.n2385 0.0514167
R21474 GNDA.n2392 GNDA.n2391 0.0514167
R21475 GNDA.n2400 GNDA.n690 0.0514167
R21476 GNDA.n2748 GNDA.n600 0.0514167
R21477 GNDA.n2758 GNDA.n2757 0.0514167
R21478 GNDA.n2764 GNDA.n2763 0.0514167
R21479 GNDA.n2774 GNDA.n2773 0.0514167
R21480 GNDA.n2778 GNDA.n2777 0.0514167
R21481 GNDA.n2788 GNDA.n2787 0.0514167
R21482 GNDA.n2794 GNDA.n2793 0.0514167
R21483 GNDA.n2804 GNDA.n2803 0.0514167
R21484 GNDA.n2808 GNDA.n2807 0.0514167
R21485 GNDA.n2818 GNDA.n2817 0.0514167
R21486 GNDA.n2824 GNDA.n2823 0.0514167
R21487 GNDA.n2834 GNDA.n2833 0.0514167
R21488 GNDA.n2838 GNDA.n2837 0.0514167
R21489 GNDA.n2848 GNDA.n2847 0.0514167
R21490 GNDA.n2854 GNDA.n2853 0.0514167
R21491 GNDA.n2862 GNDA.n624 0.0514167
R21492 GNDA.n2733 GNDA.n2732 0.0514167
R21493 GNDA.n2727 GNDA.n2726 0.0514167
R21494 GNDA.n2724 GNDA.n2723 0.0514167
R21495 GNDA.n2718 GNDA.n2717 0.0514167
R21496 GNDA.n2715 GNDA.n2714 0.0514167
R21497 GNDA.n2709 GNDA.n2708 0.0514167
R21498 GNDA.n2706 GNDA.n2705 0.0514167
R21499 GNDA.n2700 GNDA.n2699 0.0514167
R21500 GNDA.n2697 GNDA.n2696 0.0514167
R21501 GNDA.n2691 GNDA.n2690 0.0514167
R21502 GNDA.n2688 GNDA.n2687 0.0514167
R21503 GNDA.n2682 GNDA.n2681 0.0514167
R21504 GNDA.n2679 GNDA.n2678 0.0514167
R21505 GNDA.n2673 GNDA.n2672 0.0514167
R21506 GNDA.n2670 GNDA.n2669 0.0514167
R21507 GNDA.n2664 GNDA.n2663 0.0514167
R21508 GNDA.n2562 GNDA.n664 0.0514167
R21509 GNDA.n2456 GNDA.n2455 0.0514167
R21510 GNDA.n2462 GNDA.n2461 0.0514167
R21511 GNDA.n2472 GNDA.n2471 0.0514167
R21512 GNDA.n2476 GNDA.n2475 0.0514167
R21513 GNDA.n2486 GNDA.n2485 0.0514167
R21514 GNDA.n2492 GNDA.n2491 0.0514167
R21515 GNDA.n2502 GNDA.n2501 0.0514167
R21516 GNDA.n2506 GNDA.n2505 0.0514167
R21517 GNDA.n2516 GNDA.n2515 0.0514167
R21518 GNDA.n2522 GNDA.n2521 0.0514167
R21519 GNDA.n2532 GNDA.n2531 0.0514167
R21520 GNDA.n2536 GNDA.n2535 0.0514167
R21521 GNDA.n2546 GNDA.n2545 0.0514167
R21522 GNDA.n2552 GNDA.n2551 0.0514167
R21523 GNDA.n2560 GNDA.n2425 0.0514167
R21524 GNDA.n2273 GNDA.n2272 0.0514167
R21525 GNDA.n2267 GNDA.n2266 0.0514167
R21526 GNDA.n2264 GNDA.n2263 0.0514167
R21527 GNDA.n2258 GNDA.n2257 0.0514167
R21528 GNDA.n2255 GNDA.n2254 0.0514167
R21529 GNDA.n2249 GNDA.n2248 0.0514167
R21530 GNDA.n2246 GNDA.n2245 0.0514167
R21531 GNDA.n2240 GNDA.n2239 0.0514167
R21532 GNDA.n2237 GNDA.n2236 0.0514167
R21533 GNDA.n2231 GNDA.n2230 0.0514167
R21534 GNDA.n2228 GNDA.n2227 0.0514167
R21535 GNDA.n2222 GNDA.n2221 0.0514167
R21536 GNDA.n2219 GNDA.n2218 0.0514167
R21537 GNDA.n2213 GNDA.n2212 0.0514167
R21538 GNDA.n2210 GNDA.n2209 0.0514167
R21539 GNDA.n2204 GNDA.n2203 0.0514167
R21540 GNDA.n2099 GNDA.n727 0.0514167
R21541 GNDA.n1993 GNDA.n1992 0.0514167
R21542 GNDA.n1999 GNDA.n1998 0.0514167
R21543 GNDA.n2009 GNDA.n2008 0.0514167
R21544 GNDA.n2013 GNDA.n2012 0.0514167
R21545 GNDA.n2023 GNDA.n2022 0.0514167
R21546 GNDA.n2029 GNDA.n2028 0.0514167
R21547 GNDA.n2039 GNDA.n2038 0.0514167
R21548 GNDA.n2043 GNDA.n2042 0.0514167
R21549 GNDA.n2053 GNDA.n2052 0.0514167
R21550 GNDA.n2059 GNDA.n2058 0.0514167
R21551 GNDA.n2069 GNDA.n2068 0.0514167
R21552 GNDA.n2073 GNDA.n2072 0.0514167
R21553 GNDA.n2083 GNDA.n2082 0.0514167
R21554 GNDA.n2089 GNDA.n2088 0.0514167
R21555 GNDA.n2097 GNDA.n1962 0.0514167
R21556 GNDA.n1823 GNDA.n729 0.0514167
R21557 GNDA.n1833 GNDA.n1832 0.0514167
R21558 GNDA.n1839 GNDA.n1838 0.0514167
R21559 GNDA.n1849 GNDA.n1848 0.0514167
R21560 GNDA.n1853 GNDA.n1852 0.0514167
R21561 GNDA.n1863 GNDA.n1862 0.0514167
R21562 GNDA.n1869 GNDA.n1868 0.0514167
R21563 GNDA.n1879 GNDA.n1878 0.0514167
R21564 GNDA.n1883 GNDA.n1882 0.0514167
R21565 GNDA.n1893 GNDA.n1892 0.0514167
R21566 GNDA.n1899 GNDA.n1898 0.0514167
R21567 GNDA.n1909 GNDA.n1908 0.0514167
R21568 GNDA.n1913 GNDA.n1912 0.0514167
R21569 GNDA.n1923 GNDA.n1922 0.0514167
R21570 GNDA.n1929 GNDA.n1928 0.0514167
R21571 GNDA.n1937 GNDA.n753 0.0514167
R21572 GNDA.n1686 GNDA.n1685 0.0514167
R21573 GNDA.n1680 GNDA.n1679 0.0514167
R21574 GNDA.n1677 GNDA.n1676 0.0514167
R21575 GNDA.n1671 GNDA.n1670 0.0514167
R21576 GNDA.n1668 GNDA.n1667 0.0514167
R21577 GNDA.n1662 GNDA.n1661 0.0514167
R21578 GNDA.n1659 GNDA.n1658 0.0514167
R21579 GNDA.n1653 GNDA.n1652 0.0514167
R21580 GNDA.n1650 GNDA.n1649 0.0514167
R21581 GNDA.n1644 GNDA.n1643 0.0514167
R21582 GNDA.n1641 GNDA.n1640 0.0514167
R21583 GNDA.n1635 GNDA.n1634 0.0514167
R21584 GNDA.n1632 GNDA.n1631 0.0514167
R21585 GNDA.n1626 GNDA.n1625 0.0514167
R21586 GNDA.n1623 GNDA.n1622 0.0514167
R21587 GNDA.n1617 GNDA.n1616 0.0514167
R21588 GNDA.n1515 GNDA.n793 0.0514167
R21589 GNDA.n1409 GNDA.n1408 0.0514167
R21590 GNDA.n1415 GNDA.n1414 0.0514167
R21591 GNDA.n1425 GNDA.n1424 0.0514167
R21592 GNDA.n1429 GNDA.n1428 0.0514167
R21593 GNDA.n1439 GNDA.n1438 0.0514167
R21594 GNDA.n1445 GNDA.n1444 0.0514167
R21595 GNDA.n1455 GNDA.n1454 0.0514167
R21596 GNDA.n1459 GNDA.n1458 0.0514167
R21597 GNDA.n1469 GNDA.n1468 0.0514167
R21598 GNDA.n1475 GNDA.n1474 0.0514167
R21599 GNDA.n1485 GNDA.n1484 0.0514167
R21600 GNDA.n1489 GNDA.n1488 0.0514167
R21601 GNDA.n1499 GNDA.n1498 0.0514167
R21602 GNDA.n1505 GNDA.n1504 0.0514167
R21603 GNDA.n1513 GNDA.n1378 0.0514167
R21604 GNDA.n7133 GNDA.n7066 0.0514167
R21605 GNDA.n7130 GNDA.n7129 0.0514167
R21606 GNDA.n7145 GNDA.n7144 0.0514167
R21607 GNDA.n7153 GNDA.n7152 0.0514167
R21608 GNDA.n7122 GNDA.n7121 0.0514167
R21609 GNDA.n7118 GNDA.n7117 0.0514167
R21610 GNDA.n7169 GNDA.n7168 0.0514167
R21611 GNDA.n7177 GNDA.n7176 0.0514167
R21612 GNDA.n7110 GNDA.n7109 0.0514167
R21613 GNDA.n7106 GNDA.n7105 0.0514167
R21614 GNDA.n7193 GNDA.n7192 0.0514167
R21615 GNDA.n7201 GNDA.n7200 0.0514167
R21616 GNDA.n7098 GNDA.n7097 0.0514167
R21617 GNDA.n7094 GNDA.n7093 0.0514167
R21618 GNDA.n7217 GNDA.n7216 0.0514167
R21619 GNDA.n7226 GNDA.n97 0.0514167
R21620 GNDA.n147 GNDA.n99 0.0514167
R21621 GNDA.n157 GNDA.n156 0.0514167
R21622 GNDA.n163 GNDA.n162 0.0514167
R21623 GNDA.n173 GNDA.n172 0.0514167
R21624 GNDA.n177 GNDA.n176 0.0514167
R21625 GNDA.n187 GNDA.n186 0.0514167
R21626 GNDA.n193 GNDA.n192 0.0514167
R21627 GNDA.n203 GNDA.n202 0.0514167
R21628 GNDA.n207 GNDA.n206 0.0514167
R21629 GNDA.n217 GNDA.n216 0.0514167
R21630 GNDA.n223 GNDA.n222 0.0514167
R21631 GNDA.n233 GNDA.n232 0.0514167
R21632 GNDA.n237 GNDA.n236 0.0514167
R21633 GNDA.n247 GNDA.n246 0.0514167
R21634 GNDA.n253 GNDA.n252 0.0514167
R21635 GNDA.n7064 GNDA.n123 0.0514167
R21636 GNDA.n1253 GNDA.n1252 0.0475
R21637 GNDA.n1266 GNDA.n1265 0.0475
R21638 GNDA.n1283 GNDA.n1282 0.0475
R21639 GNDA.n1296 GNDA.n1295 0.0475
R21640 GNDA.n1313 GNDA.n1312 0.0475
R21641 GNDA.n1326 GNDA.n1325 0.0475
R21642 GNDA.n1343 GNDA.n1342 0.0475
R21643 GNDA.n3406 GNDA.n589 0.0421667
R21644 GNDA.n1724 GNDA.n1718 0.0421667
R21645 GNDA.n1769 GNDA.n1767 0.0421667
R21646 GNDA.n1784 GNDA.n1703 0.0421667
R21647 GNDA.n3678 GNDA.n3676 0.0421667
R21648 GNDA.n2283 GNDA.n715 0.0421667
R21649 GNDA.n1227 GNDA.n1220 0.0421667
R21650 GNDA.n1232 GNDA.n1217 0.0421667
R21651 GNDA.n1234 GNDA.n789 0.0421667
R21652 GNDA.n1522 GNDA.n786 0.0421667
R21653 GNDA.n1693 GNDA.n783 0.0421667
R21654 GNDA.n1815 GNDA.n780 0.0421667
R21655 GNDA.n778 GNDA.n723 0.0421667
R21656 GNDA.n2106 GNDA.n720 0.0421667
R21657 GNDA.n2280 GNDA.n716 0.0421667
R21658 GNDA.n2569 GNDA.n655 0.0421667
R21659 GNDA.n2740 GNDA.n652 0.0421667
R21660 GNDA.n650 GNDA.n649 0.0421667
R21661 GNDA.n2913 GNDA.n594 0.0421667
R21662 GNDA.n3205 GNDA.n591 0.0421667
R21663 GNDA.n3377 GNDA.n3376 0.0421667
R21664 GNDA.n5278 GNDA.n323 0.0421667
R21665 GNDA.n5011 GNDA.n5010 0.0421667
R21666 GNDA.n5007 GNDA.n5006 0.0421667
R21667 GNDA.n3509 GNDA.n576 0.0421667
R21668 GNDA.n4995 GNDA.n4994 0.0421667
R21669 GNDA.n4991 GNDA.n4990 0.0421667
R21670 GNDA.n4987 GNDA.n4986 0.0421667
R21671 GNDA.n4983 GNDA.n4982 0.0421667
R21672 GNDA.n4979 GNDA.n4978 0.0421667
R21673 GNDA.n4975 GNDA.n4974 0.0421667
R21674 GNDA.n4971 GNDA.n4970 0.0421667
R21675 GNDA.n4967 GNDA.n4966 0.0421667
R21676 GNDA.n6778 GNDA.n6654 0.0421667
R21677 GNDA.n7231 GNDA.n94 0.0421667
R21678 GNDA.n1057 GNDA 0.0414781
R21679 GNDA.n5162 GNDA.n330 0.028198
R21680 GNDA.n5166 GNDA.n331 0.028198
R21681 GNDA.n5176 GNDA.n333 0.028198
R21682 GNDA.n5182 GNDA.n334 0.028198
R21683 GNDA.n5192 GNDA.n336 0.028198
R21684 GNDA.n5196 GNDA.n337 0.028198
R21685 GNDA.n5206 GNDA.n339 0.028198
R21686 GNDA.n5212 GNDA.n340 0.028198
R21687 GNDA.n5222 GNDA.n342 0.028198
R21688 GNDA.n5226 GNDA.n343 0.028198
R21689 GNDA.n5236 GNDA.n345 0.028198
R21690 GNDA.n5242 GNDA.n346 0.028198
R21691 GNDA.n5252 GNDA.n348 0.028198
R21692 GNDA.n5256 GNDA.n349 0.028198
R21693 GNDA.n5266 GNDA.n351 0.028198
R21694 GNDA.n5136 GNDA.n352 0.028198
R21695 GNDA.n4849 GNDA.n4800 0.028198
R21696 GNDA.n4853 GNDA.n4801 0.028198
R21697 GNDA.n4863 GNDA.n4803 0.028198
R21698 GNDA.n4869 GNDA.n4804 0.028198
R21699 GNDA.n4879 GNDA.n4806 0.028198
R21700 GNDA.n4883 GNDA.n4807 0.028198
R21701 GNDA.n4893 GNDA.n4809 0.028198
R21702 GNDA.n4899 GNDA.n4810 0.028198
R21703 GNDA.n4909 GNDA.n4812 0.028198
R21704 GNDA.n4913 GNDA.n4813 0.028198
R21705 GNDA.n4923 GNDA.n4815 0.028198
R21706 GNDA.n4929 GNDA.n4816 0.028198
R21707 GNDA.n4939 GNDA.n4818 0.028198
R21708 GNDA.n4943 GNDA.n4819 0.028198
R21709 GNDA.n4953 GNDA.n4821 0.028198
R21710 GNDA.n4823 GNDA.n4822 0.028198
R21711 GNDA.n4689 GNDA.n4635 0.028198
R21712 GNDA.n4693 GNDA.n4636 0.028198
R21713 GNDA.n4703 GNDA.n4638 0.028198
R21714 GNDA.n4709 GNDA.n4639 0.028198
R21715 GNDA.n4719 GNDA.n4641 0.028198
R21716 GNDA.n4723 GNDA.n4642 0.028198
R21717 GNDA.n4733 GNDA.n4644 0.028198
R21718 GNDA.n4739 GNDA.n4645 0.028198
R21719 GNDA.n4749 GNDA.n4647 0.028198
R21720 GNDA.n4753 GNDA.n4648 0.028198
R21721 GNDA.n4763 GNDA.n4650 0.028198
R21722 GNDA.n4769 GNDA.n4651 0.028198
R21723 GNDA.n4779 GNDA.n4653 0.028198
R21724 GNDA.n4783 GNDA.n4654 0.028198
R21725 GNDA.n4793 GNDA.n4656 0.028198
R21726 GNDA.n4658 GNDA.n4657 0.028198
R21727 GNDA.n4523 GNDA.n4469 0.028198
R21728 GNDA.n4527 GNDA.n4470 0.028198
R21729 GNDA.n4537 GNDA.n4472 0.028198
R21730 GNDA.n4543 GNDA.n4473 0.028198
R21731 GNDA.n4553 GNDA.n4475 0.028198
R21732 GNDA.n4557 GNDA.n4476 0.028198
R21733 GNDA.n4567 GNDA.n4478 0.028198
R21734 GNDA.n4573 GNDA.n4479 0.028198
R21735 GNDA.n4583 GNDA.n4481 0.028198
R21736 GNDA.n4587 GNDA.n4482 0.028198
R21737 GNDA.n4597 GNDA.n4484 0.028198
R21738 GNDA.n4603 GNDA.n4485 0.028198
R21739 GNDA.n4613 GNDA.n4487 0.028198
R21740 GNDA.n4617 GNDA.n4488 0.028198
R21741 GNDA.n4627 GNDA.n4490 0.028198
R21742 GNDA.n4492 GNDA.n4491 0.028198
R21743 GNDA.n4357 GNDA.n4303 0.028198
R21744 GNDA.n4361 GNDA.n4304 0.028198
R21745 GNDA.n4371 GNDA.n4306 0.028198
R21746 GNDA.n4377 GNDA.n4307 0.028198
R21747 GNDA.n4387 GNDA.n4309 0.028198
R21748 GNDA.n4391 GNDA.n4310 0.028198
R21749 GNDA.n4401 GNDA.n4312 0.028198
R21750 GNDA.n4407 GNDA.n4313 0.028198
R21751 GNDA.n4417 GNDA.n4315 0.028198
R21752 GNDA.n4421 GNDA.n4316 0.028198
R21753 GNDA.n4431 GNDA.n4318 0.028198
R21754 GNDA.n4437 GNDA.n4319 0.028198
R21755 GNDA.n4447 GNDA.n4321 0.028198
R21756 GNDA.n4451 GNDA.n4322 0.028198
R21757 GNDA.n4461 GNDA.n4324 0.028198
R21758 GNDA.n4326 GNDA.n4325 0.028198
R21759 GNDA.n4191 GNDA.n4137 0.028198
R21760 GNDA.n4195 GNDA.n4138 0.028198
R21761 GNDA.n4205 GNDA.n4140 0.028198
R21762 GNDA.n4211 GNDA.n4141 0.028198
R21763 GNDA.n4221 GNDA.n4143 0.028198
R21764 GNDA.n4225 GNDA.n4144 0.028198
R21765 GNDA.n4235 GNDA.n4146 0.028198
R21766 GNDA.n4241 GNDA.n4147 0.028198
R21767 GNDA.n4251 GNDA.n4149 0.028198
R21768 GNDA.n4255 GNDA.n4150 0.028198
R21769 GNDA.n4265 GNDA.n4152 0.028198
R21770 GNDA.n4271 GNDA.n4153 0.028198
R21771 GNDA.n4281 GNDA.n4155 0.028198
R21772 GNDA.n4285 GNDA.n4156 0.028198
R21773 GNDA.n4295 GNDA.n4158 0.028198
R21774 GNDA.n4160 GNDA.n4159 0.028198
R21775 GNDA.n3693 GNDA.n3461 0.028198
R21776 GNDA.n3697 GNDA.n3462 0.028198
R21777 GNDA.n3707 GNDA.n3464 0.028198
R21778 GNDA.n3713 GNDA.n3465 0.028198
R21779 GNDA.n3723 GNDA.n3467 0.028198
R21780 GNDA.n3727 GNDA.n3468 0.028198
R21781 GNDA.n3737 GNDA.n3470 0.028198
R21782 GNDA.n3743 GNDA.n3471 0.028198
R21783 GNDA.n3753 GNDA.n3473 0.028198
R21784 GNDA.n3757 GNDA.n3474 0.028198
R21785 GNDA.n3767 GNDA.n3476 0.028198
R21786 GNDA.n3773 GNDA.n3477 0.028198
R21787 GNDA.n3783 GNDA.n3479 0.028198
R21788 GNDA.n3787 GNDA.n3480 0.028198
R21789 GNDA.n3797 GNDA.n3482 0.028198
R21790 GNDA.n3484 GNDA.n3483 0.028198
R21791 GNDA.n4025 GNDA.n3971 0.028198
R21792 GNDA.n4029 GNDA.n3972 0.028198
R21793 GNDA.n4039 GNDA.n3974 0.028198
R21794 GNDA.n4045 GNDA.n3975 0.028198
R21795 GNDA.n4055 GNDA.n3977 0.028198
R21796 GNDA.n4059 GNDA.n3978 0.028198
R21797 GNDA.n4069 GNDA.n3980 0.028198
R21798 GNDA.n4075 GNDA.n3981 0.028198
R21799 GNDA.n4085 GNDA.n3983 0.028198
R21800 GNDA.n4089 GNDA.n3984 0.028198
R21801 GNDA.n4099 GNDA.n3986 0.028198
R21802 GNDA.n4105 GNDA.n3987 0.028198
R21803 GNDA.n4115 GNDA.n3989 0.028198
R21804 GNDA.n4119 GNDA.n3990 0.028198
R21805 GNDA.n4129 GNDA.n3992 0.028198
R21806 GNDA.n3994 GNDA.n3993 0.028198
R21807 GNDA.n3859 GNDA.n3805 0.028198
R21808 GNDA.n3863 GNDA.n3806 0.028198
R21809 GNDA.n3873 GNDA.n3808 0.028198
R21810 GNDA.n3879 GNDA.n3809 0.028198
R21811 GNDA.n3889 GNDA.n3811 0.028198
R21812 GNDA.n3893 GNDA.n3812 0.028198
R21813 GNDA.n3903 GNDA.n3814 0.028198
R21814 GNDA.n3909 GNDA.n3815 0.028198
R21815 GNDA.n3919 GNDA.n3817 0.028198
R21816 GNDA.n3923 GNDA.n3818 0.028198
R21817 GNDA.n3933 GNDA.n3820 0.028198
R21818 GNDA.n3939 GNDA.n3821 0.028198
R21819 GNDA.n3949 GNDA.n3823 0.028198
R21820 GNDA.n3953 GNDA.n3824 0.028198
R21821 GNDA.n3963 GNDA.n3826 0.028198
R21822 GNDA.n3828 GNDA.n3827 0.028198
R21823 GNDA.n3671 GNDA.n3670 0.028198
R21824 GNDA.n3668 GNDA.n3667 0.028198
R21825 GNDA.n3662 GNDA.n3661 0.028198
R21826 GNDA.n3659 GNDA.n3658 0.028198
R21827 GNDA.n3653 GNDA.n3652 0.028198
R21828 GNDA.n3650 GNDA.n3649 0.028198
R21829 GNDA.n3644 GNDA.n3643 0.028198
R21830 GNDA.n3641 GNDA.n3640 0.028198
R21831 GNDA.n3635 GNDA.n3634 0.028198
R21832 GNDA.n3632 GNDA.n3631 0.028198
R21833 GNDA.n3626 GNDA.n3625 0.028198
R21834 GNDA.n3623 GNDA.n3622 0.028198
R21835 GNDA.n3617 GNDA.n3616 0.028198
R21836 GNDA.n3614 GNDA.n3613 0.028198
R21837 GNDA.n3608 GNDA.n3607 0.028198
R21838 GNDA.n3605 GNDA.n3604 0.028198
R21839 GNDA.n565 GNDA.n564 0.028198
R21840 GNDA.n562 GNDA.n561 0.028198
R21841 GNDA.n556 GNDA.n555 0.028198
R21842 GNDA.n553 GNDA.n552 0.028198
R21843 GNDA.n547 GNDA.n546 0.028198
R21844 GNDA.n544 GNDA.n543 0.028198
R21845 GNDA.n538 GNDA.n537 0.028198
R21846 GNDA.n535 GNDA.n534 0.028198
R21847 GNDA.n529 GNDA.n528 0.028198
R21848 GNDA.n526 GNDA.n525 0.028198
R21849 GNDA.n520 GNDA.n519 0.028198
R21850 GNDA.n517 GNDA.n516 0.028198
R21851 GNDA.n511 GNDA.n510 0.028198
R21852 GNDA.n508 GNDA.n507 0.028198
R21853 GNDA.n502 GNDA.n501 0.028198
R21854 GNDA.n499 GNDA.n498 0.028198
R21855 GNDA.n5025 GNDA.n354 0.028198
R21856 GNDA.n5029 GNDA.n355 0.028198
R21857 GNDA.n5039 GNDA.n357 0.028198
R21858 GNDA.n5045 GNDA.n358 0.028198
R21859 GNDA.n5055 GNDA.n360 0.028198
R21860 GNDA.n5059 GNDA.n361 0.028198
R21861 GNDA.n5069 GNDA.n363 0.028198
R21862 GNDA.n5075 GNDA.n364 0.028198
R21863 GNDA.n5085 GNDA.n366 0.028198
R21864 GNDA.n5089 GNDA.n367 0.028198
R21865 GNDA.n5099 GNDA.n369 0.028198
R21866 GNDA.n5105 GNDA.n370 0.028198
R21867 GNDA.n5115 GNDA.n372 0.028198
R21868 GNDA.n5119 GNDA.n373 0.028198
R21869 GNDA.n5129 GNDA.n375 0.028198
R21870 GNDA.n378 GNDA.n376 0.028198
R21871 GNDA.n3368 GNDA.n3367 0.028198
R21872 GNDA.n3365 GNDA.n3364 0.028198
R21873 GNDA.n3359 GNDA.n3358 0.028198
R21874 GNDA.n3356 GNDA.n3355 0.028198
R21875 GNDA.n3350 GNDA.n3349 0.028198
R21876 GNDA.n3347 GNDA.n3346 0.028198
R21877 GNDA.n3341 GNDA.n3340 0.028198
R21878 GNDA.n3338 GNDA.n3337 0.028198
R21879 GNDA.n3332 GNDA.n3331 0.028198
R21880 GNDA.n3329 GNDA.n3328 0.028198
R21881 GNDA.n3323 GNDA.n3322 0.028198
R21882 GNDA.n3320 GNDA.n3319 0.028198
R21883 GNDA.n3314 GNDA.n3313 0.028198
R21884 GNDA.n3311 GNDA.n3310 0.028198
R21885 GNDA.n3305 GNDA.n3304 0.028198
R21886 GNDA.n3302 GNDA.n3301 0.028198
R21887 GNDA.n3087 GNDA.n3038 0.028198
R21888 GNDA.n3091 GNDA.n3039 0.028198
R21889 GNDA.n3101 GNDA.n3041 0.028198
R21890 GNDA.n3107 GNDA.n3042 0.028198
R21891 GNDA.n3117 GNDA.n3044 0.028198
R21892 GNDA.n3121 GNDA.n3045 0.028198
R21893 GNDA.n3131 GNDA.n3047 0.028198
R21894 GNDA.n3137 GNDA.n3048 0.028198
R21895 GNDA.n3147 GNDA.n3050 0.028198
R21896 GNDA.n3151 GNDA.n3051 0.028198
R21897 GNDA.n3161 GNDA.n3053 0.028198
R21898 GNDA.n3167 GNDA.n3054 0.028198
R21899 GNDA.n3177 GNDA.n3056 0.028198
R21900 GNDA.n3181 GNDA.n3057 0.028198
R21901 GNDA.n3191 GNDA.n3059 0.028198
R21902 GNDA.n3061 GNDA.n3060 0.028198
R21903 GNDA.n2927 GNDA.n2865 0.028198
R21904 GNDA.n2931 GNDA.n2866 0.028198
R21905 GNDA.n2941 GNDA.n2868 0.028198
R21906 GNDA.n2947 GNDA.n2869 0.028198
R21907 GNDA.n2957 GNDA.n2871 0.028198
R21908 GNDA.n2961 GNDA.n2872 0.028198
R21909 GNDA.n2971 GNDA.n2874 0.028198
R21910 GNDA.n2977 GNDA.n2875 0.028198
R21911 GNDA.n2987 GNDA.n2877 0.028198
R21912 GNDA.n2991 GNDA.n2878 0.028198
R21913 GNDA.n3001 GNDA.n2880 0.028198
R21914 GNDA.n3007 GNDA.n2881 0.028198
R21915 GNDA.n3017 GNDA.n2883 0.028198
R21916 GNDA.n3021 GNDA.n2884 0.028198
R21917 GNDA.n3031 GNDA.n2886 0.028198
R21918 GNDA.n2888 GNDA.n2887 0.028198
R21919 GNDA.n2291 GNDA.n667 0.028198
R21920 GNDA.n2295 GNDA.n668 0.028198
R21921 GNDA.n2305 GNDA.n670 0.028198
R21922 GNDA.n2311 GNDA.n671 0.028198
R21923 GNDA.n2321 GNDA.n673 0.028198
R21924 GNDA.n2325 GNDA.n674 0.028198
R21925 GNDA.n2335 GNDA.n676 0.028198
R21926 GNDA.n2341 GNDA.n677 0.028198
R21927 GNDA.n2351 GNDA.n679 0.028198
R21928 GNDA.n2355 GNDA.n680 0.028198
R21929 GNDA.n2365 GNDA.n682 0.028198
R21930 GNDA.n2371 GNDA.n683 0.028198
R21931 GNDA.n2381 GNDA.n685 0.028198
R21932 GNDA.n2385 GNDA.n686 0.028198
R21933 GNDA.n2395 GNDA.n688 0.028198
R21934 GNDA.n690 GNDA.n689 0.028198
R21935 GNDA.n2753 GNDA.n601 0.028198
R21936 GNDA.n2757 GNDA.n602 0.028198
R21937 GNDA.n2767 GNDA.n604 0.028198
R21938 GNDA.n2773 GNDA.n605 0.028198
R21939 GNDA.n2783 GNDA.n607 0.028198
R21940 GNDA.n2787 GNDA.n608 0.028198
R21941 GNDA.n2797 GNDA.n610 0.028198
R21942 GNDA.n2803 GNDA.n611 0.028198
R21943 GNDA.n2813 GNDA.n613 0.028198
R21944 GNDA.n2817 GNDA.n614 0.028198
R21945 GNDA.n2827 GNDA.n616 0.028198
R21946 GNDA.n2833 GNDA.n617 0.028198
R21947 GNDA.n2843 GNDA.n619 0.028198
R21948 GNDA.n2847 GNDA.n620 0.028198
R21949 GNDA.n2857 GNDA.n622 0.028198
R21950 GNDA.n624 GNDA.n623 0.028198
R21951 GNDA.n2731 GNDA.n2730 0.028198
R21952 GNDA.n2728 GNDA.n2727 0.028198
R21953 GNDA.n2722 GNDA.n2721 0.028198
R21954 GNDA.n2719 GNDA.n2718 0.028198
R21955 GNDA.n2713 GNDA.n2712 0.028198
R21956 GNDA.n2710 GNDA.n2709 0.028198
R21957 GNDA.n2704 GNDA.n2703 0.028198
R21958 GNDA.n2701 GNDA.n2700 0.028198
R21959 GNDA.n2695 GNDA.n2694 0.028198
R21960 GNDA.n2692 GNDA.n2691 0.028198
R21961 GNDA.n2686 GNDA.n2685 0.028198
R21962 GNDA.n2683 GNDA.n2682 0.028198
R21963 GNDA.n2677 GNDA.n2676 0.028198
R21964 GNDA.n2674 GNDA.n2673 0.028198
R21965 GNDA.n2668 GNDA.n2667 0.028198
R21966 GNDA.n2665 GNDA.n2664 0.028198
R21967 GNDA.n2451 GNDA.n2402 0.028198
R21968 GNDA.n2455 GNDA.n2403 0.028198
R21969 GNDA.n2465 GNDA.n2405 0.028198
R21970 GNDA.n2471 GNDA.n2406 0.028198
R21971 GNDA.n2481 GNDA.n2408 0.028198
R21972 GNDA.n2485 GNDA.n2409 0.028198
R21973 GNDA.n2495 GNDA.n2411 0.028198
R21974 GNDA.n2501 GNDA.n2412 0.028198
R21975 GNDA.n2511 GNDA.n2414 0.028198
R21976 GNDA.n2515 GNDA.n2415 0.028198
R21977 GNDA.n2525 GNDA.n2417 0.028198
R21978 GNDA.n2531 GNDA.n2418 0.028198
R21979 GNDA.n2541 GNDA.n2420 0.028198
R21980 GNDA.n2545 GNDA.n2421 0.028198
R21981 GNDA.n2555 GNDA.n2423 0.028198
R21982 GNDA.n2425 GNDA.n2424 0.028198
R21983 GNDA.n2271 GNDA.n2270 0.028198
R21984 GNDA.n2268 GNDA.n2267 0.028198
R21985 GNDA.n2262 GNDA.n2261 0.028198
R21986 GNDA.n2259 GNDA.n2258 0.028198
R21987 GNDA.n2253 GNDA.n2252 0.028198
R21988 GNDA.n2250 GNDA.n2249 0.028198
R21989 GNDA.n2244 GNDA.n2243 0.028198
R21990 GNDA.n2241 GNDA.n2240 0.028198
R21991 GNDA.n2235 GNDA.n2234 0.028198
R21992 GNDA.n2232 GNDA.n2231 0.028198
R21993 GNDA.n2226 GNDA.n2225 0.028198
R21994 GNDA.n2223 GNDA.n2222 0.028198
R21995 GNDA.n2217 GNDA.n2216 0.028198
R21996 GNDA.n2214 GNDA.n2213 0.028198
R21997 GNDA.n2208 GNDA.n2207 0.028198
R21998 GNDA.n2205 GNDA.n2204 0.028198
R21999 GNDA.n1988 GNDA.n1939 0.028198
R22000 GNDA.n1992 GNDA.n1940 0.028198
R22001 GNDA.n2002 GNDA.n1942 0.028198
R22002 GNDA.n2008 GNDA.n1943 0.028198
R22003 GNDA.n2018 GNDA.n1945 0.028198
R22004 GNDA.n2022 GNDA.n1946 0.028198
R22005 GNDA.n2032 GNDA.n1948 0.028198
R22006 GNDA.n2038 GNDA.n1949 0.028198
R22007 GNDA.n2048 GNDA.n1951 0.028198
R22008 GNDA.n2052 GNDA.n1952 0.028198
R22009 GNDA.n2062 GNDA.n1954 0.028198
R22010 GNDA.n2068 GNDA.n1955 0.028198
R22011 GNDA.n2078 GNDA.n1957 0.028198
R22012 GNDA.n2082 GNDA.n1958 0.028198
R22013 GNDA.n2092 GNDA.n1960 0.028198
R22014 GNDA.n1962 GNDA.n1961 0.028198
R22015 GNDA.n1828 GNDA.n730 0.028198
R22016 GNDA.n1832 GNDA.n731 0.028198
R22017 GNDA.n1842 GNDA.n733 0.028198
R22018 GNDA.n1848 GNDA.n734 0.028198
R22019 GNDA.n1858 GNDA.n736 0.028198
R22020 GNDA.n1862 GNDA.n737 0.028198
R22021 GNDA.n1872 GNDA.n739 0.028198
R22022 GNDA.n1878 GNDA.n740 0.028198
R22023 GNDA.n1888 GNDA.n742 0.028198
R22024 GNDA.n1892 GNDA.n743 0.028198
R22025 GNDA.n1902 GNDA.n745 0.028198
R22026 GNDA.n1908 GNDA.n746 0.028198
R22027 GNDA.n1918 GNDA.n748 0.028198
R22028 GNDA.n1922 GNDA.n749 0.028198
R22029 GNDA.n1932 GNDA.n751 0.028198
R22030 GNDA.n753 GNDA.n752 0.028198
R22031 GNDA.n1684 GNDA.n1683 0.028198
R22032 GNDA.n1681 GNDA.n1680 0.028198
R22033 GNDA.n1675 GNDA.n1674 0.028198
R22034 GNDA.n1672 GNDA.n1671 0.028198
R22035 GNDA.n1666 GNDA.n1665 0.028198
R22036 GNDA.n1663 GNDA.n1662 0.028198
R22037 GNDA.n1657 GNDA.n1656 0.028198
R22038 GNDA.n1654 GNDA.n1653 0.028198
R22039 GNDA.n1648 GNDA.n1647 0.028198
R22040 GNDA.n1645 GNDA.n1644 0.028198
R22041 GNDA.n1639 GNDA.n1638 0.028198
R22042 GNDA.n1636 GNDA.n1635 0.028198
R22043 GNDA.n1630 GNDA.n1629 0.028198
R22044 GNDA.n1627 GNDA.n1626 0.028198
R22045 GNDA.n1621 GNDA.n1620 0.028198
R22046 GNDA.n1618 GNDA.n1617 0.028198
R22047 GNDA.n1404 GNDA.n1355 0.028198
R22048 GNDA.n1408 GNDA.n1356 0.028198
R22049 GNDA.n1418 GNDA.n1358 0.028198
R22050 GNDA.n1424 GNDA.n1359 0.028198
R22051 GNDA.n1434 GNDA.n1361 0.028198
R22052 GNDA.n1438 GNDA.n1362 0.028198
R22053 GNDA.n1448 GNDA.n1364 0.028198
R22054 GNDA.n1454 GNDA.n1365 0.028198
R22055 GNDA.n1464 GNDA.n1367 0.028198
R22056 GNDA.n1468 GNDA.n1368 0.028198
R22057 GNDA.n1478 GNDA.n1370 0.028198
R22058 GNDA.n1484 GNDA.n1371 0.028198
R22059 GNDA.n1494 GNDA.n1373 0.028198
R22060 GNDA.n1498 GNDA.n1374 0.028198
R22061 GNDA.n1508 GNDA.n1376 0.028198
R22062 GNDA.n1378 GNDA.n1377 0.028198
R22063 GNDA.n1509 GNDA.n1377 0.028198
R22064 GNDA.n1505 GNDA.n1376 0.028198
R22065 GNDA.n1495 GNDA.n1374 0.028198
R22066 GNDA.n1489 GNDA.n1373 0.028198
R22067 GNDA.n1479 GNDA.n1371 0.028198
R22068 GNDA.n1475 GNDA.n1370 0.028198
R22069 GNDA.n1465 GNDA.n1368 0.028198
R22070 GNDA.n1459 GNDA.n1367 0.028198
R22071 GNDA.n1449 GNDA.n1365 0.028198
R22072 GNDA.n1445 GNDA.n1364 0.028198
R22073 GNDA.n1435 GNDA.n1362 0.028198
R22074 GNDA.n1429 GNDA.n1361 0.028198
R22075 GNDA.n1419 GNDA.n1359 0.028198
R22076 GNDA.n1415 GNDA.n1358 0.028198
R22077 GNDA.n1405 GNDA.n1356 0.028198
R22078 GNDA.n1355 GNDA.n793 0.028198
R22079 GNDA.n1619 GNDA.n1618 0.028198
R22080 GNDA.n1622 GNDA.n1621 0.028198
R22081 GNDA.n1628 GNDA.n1627 0.028198
R22082 GNDA.n1631 GNDA.n1630 0.028198
R22083 GNDA.n1637 GNDA.n1636 0.028198
R22084 GNDA.n1640 GNDA.n1639 0.028198
R22085 GNDA.n1646 GNDA.n1645 0.028198
R22086 GNDA.n1649 GNDA.n1648 0.028198
R22087 GNDA.n1655 GNDA.n1654 0.028198
R22088 GNDA.n1658 GNDA.n1657 0.028198
R22089 GNDA.n1664 GNDA.n1663 0.028198
R22090 GNDA.n1667 GNDA.n1666 0.028198
R22091 GNDA.n1673 GNDA.n1672 0.028198
R22092 GNDA.n1676 GNDA.n1675 0.028198
R22093 GNDA.n1682 GNDA.n1681 0.028198
R22094 GNDA.n1685 GNDA.n1684 0.028198
R22095 GNDA.n1933 GNDA.n752 0.028198
R22096 GNDA.n1929 GNDA.n751 0.028198
R22097 GNDA.n1919 GNDA.n749 0.028198
R22098 GNDA.n1913 GNDA.n748 0.028198
R22099 GNDA.n1903 GNDA.n746 0.028198
R22100 GNDA.n1899 GNDA.n745 0.028198
R22101 GNDA.n1889 GNDA.n743 0.028198
R22102 GNDA.n1883 GNDA.n742 0.028198
R22103 GNDA.n1873 GNDA.n740 0.028198
R22104 GNDA.n1869 GNDA.n739 0.028198
R22105 GNDA.n1859 GNDA.n737 0.028198
R22106 GNDA.n1853 GNDA.n736 0.028198
R22107 GNDA.n1843 GNDA.n734 0.028198
R22108 GNDA.n1839 GNDA.n733 0.028198
R22109 GNDA.n1829 GNDA.n731 0.028198
R22110 GNDA.n1823 GNDA.n730 0.028198
R22111 GNDA.n2093 GNDA.n1961 0.028198
R22112 GNDA.n2089 GNDA.n1960 0.028198
R22113 GNDA.n2079 GNDA.n1958 0.028198
R22114 GNDA.n2073 GNDA.n1957 0.028198
R22115 GNDA.n2063 GNDA.n1955 0.028198
R22116 GNDA.n2059 GNDA.n1954 0.028198
R22117 GNDA.n2049 GNDA.n1952 0.028198
R22118 GNDA.n2043 GNDA.n1951 0.028198
R22119 GNDA.n2033 GNDA.n1949 0.028198
R22120 GNDA.n2029 GNDA.n1948 0.028198
R22121 GNDA.n2019 GNDA.n1946 0.028198
R22122 GNDA.n2013 GNDA.n1945 0.028198
R22123 GNDA.n2003 GNDA.n1943 0.028198
R22124 GNDA.n1999 GNDA.n1942 0.028198
R22125 GNDA.n1989 GNDA.n1940 0.028198
R22126 GNDA.n1939 GNDA.n727 0.028198
R22127 GNDA.n2206 GNDA.n2205 0.028198
R22128 GNDA.n2209 GNDA.n2208 0.028198
R22129 GNDA.n2215 GNDA.n2214 0.028198
R22130 GNDA.n2218 GNDA.n2217 0.028198
R22131 GNDA.n2224 GNDA.n2223 0.028198
R22132 GNDA.n2227 GNDA.n2226 0.028198
R22133 GNDA.n2233 GNDA.n2232 0.028198
R22134 GNDA.n2236 GNDA.n2235 0.028198
R22135 GNDA.n2242 GNDA.n2241 0.028198
R22136 GNDA.n2245 GNDA.n2244 0.028198
R22137 GNDA.n2251 GNDA.n2250 0.028198
R22138 GNDA.n2254 GNDA.n2253 0.028198
R22139 GNDA.n2260 GNDA.n2259 0.028198
R22140 GNDA.n2263 GNDA.n2262 0.028198
R22141 GNDA.n2269 GNDA.n2268 0.028198
R22142 GNDA.n2272 GNDA.n2271 0.028198
R22143 GNDA.n2556 GNDA.n2424 0.028198
R22144 GNDA.n2552 GNDA.n2423 0.028198
R22145 GNDA.n2542 GNDA.n2421 0.028198
R22146 GNDA.n2536 GNDA.n2420 0.028198
R22147 GNDA.n2526 GNDA.n2418 0.028198
R22148 GNDA.n2522 GNDA.n2417 0.028198
R22149 GNDA.n2512 GNDA.n2415 0.028198
R22150 GNDA.n2506 GNDA.n2414 0.028198
R22151 GNDA.n2496 GNDA.n2412 0.028198
R22152 GNDA.n2492 GNDA.n2411 0.028198
R22153 GNDA.n2482 GNDA.n2409 0.028198
R22154 GNDA.n2476 GNDA.n2408 0.028198
R22155 GNDA.n2466 GNDA.n2406 0.028198
R22156 GNDA.n2462 GNDA.n2405 0.028198
R22157 GNDA.n2452 GNDA.n2403 0.028198
R22158 GNDA.n2402 GNDA.n664 0.028198
R22159 GNDA.n2666 GNDA.n2665 0.028198
R22160 GNDA.n2669 GNDA.n2668 0.028198
R22161 GNDA.n2675 GNDA.n2674 0.028198
R22162 GNDA.n2678 GNDA.n2677 0.028198
R22163 GNDA.n2684 GNDA.n2683 0.028198
R22164 GNDA.n2687 GNDA.n2686 0.028198
R22165 GNDA.n2693 GNDA.n2692 0.028198
R22166 GNDA.n2696 GNDA.n2695 0.028198
R22167 GNDA.n2702 GNDA.n2701 0.028198
R22168 GNDA.n2705 GNDA.n2704 0.028198
R22169 GNDA.n2711 GNDA.n2710 0.028198
R22170 GNDA.n2714 GNDA.n2713 0.028198
R22171 GNDA.n2720 GNDA.n2719 0.028198
R22172 GNDA.n2723 GNDA.n2722 0.028198
R22173 GNDA.n2729 GNDA.n2728 0.028198
R22174 GNDA.n2732 GNDA.n2731 0.028198
R22175 GNDA.n2858 GNDA.n623 0.028198
R22176 GNDA.n2854 GNDA.n622 0.028198
R22177 GNDA.n2844 GNDA.n620 0.028198
R22178 GNDA.n2838 GNDA.n619 0.028198
R22179 GNDA.n2828 GNDA.n617 0.028198
R22180 GNDA.n2824 GNDA.n616 0.028198
R22181 GNDA.n2814 GNDA.n614 0.028198
R22182 GNDA.n2808 GNDA.n613 0.028198
R22183 GNDA.n2798 GNDA.n611 0.028198
R22184 GNDA.n2794 GNDA.n610 0.028198
R22185 GNDA.n2784 GNDA.n608 0.028198
R22186 GNDA.n2778 GNDA.n607 0.028198
R22187 GNDA.n2768 GNDA.n605 0.028198
R22188 GNDA.n2764 GNDA.n604 0.028198
R22189 GNDA.n2754 GNDA.n602 0.028198
R22190 GNDA.n2748 GNDA.n601 0.028198
R22191 GNDA.n2396 GNDA.n689 0.028198
R22192 GNDA.n2392 GNDA.n688 0.028198
R22193 GNDA.n2382 GNDA.n686 0.028198
R22194 GNDA.n2376 GNDA.n685 0.028198
R22195 GNDA.n2366 GNDA.n683 0.028198
R22196 GNDA.n2362 GNDA.n682 0.028198
R22197 GNDA.n2352 GNDA.n680 0.028198
R22198 GNDA.n2346 GNDA.n679 0.028198
R22199 GNDA.n2336 GNDA.n677 0.028198
R22200 GNDA.n2332 GNDA.n676 0.028198
R22201 GNDA.n2322 GNDA.n674 0.028198
R22202 GNDA.n2316 GNDA.n673 0.028198
R22203 GNDA.n2306 GNDA.n671 0.028198
R22204 GNDA.n2302 GNDA.n670 0.028198
R22205 GNDA.n2292 GNDA.n668 0.028198
R22206 GNDA.n2286 GNDA.n667 0.028198
R22207 GNDA.n3032 GNDA.n2887 0.028198
R22208 GNDA.n3028 GNDA.n2886 0.028198
R22209 GNDA.n3018 GNDA.n2884 0.028198
R22210 GNDA.n3012 GNDA.n2883 0.028198
R22211 GNDA.n3002 GNDA.n2881 0.028198
R22212 GNDA.n2998 GNDA.n2880 0.028198
R22213 GNDA.n2988 GNDA.n2878 0.028198
R22214 GNDA.n2982 GNDA.n2877 0.028198
R22215 GNDA.n2972 GNDA.n2875 0.028198
R22216 GNDA.n2968 GNDA.n2874 0.028198
R22217 GNDA.n2958 GNDA.n2872 0.028198
R22218 GNDA.n2952 GNDA.n2871 0.028198
R22219 GNDA.n2942 GNDA.n2869 0.028198
R22220 GNDA.n2938 GNDA.n2868 0.028198
R22221 GNDA.n2928 GNDA.n2866 0.028198
R22222 GNDA.n2922 GNDA.n2865 0.028198
R22223 GNDA.n3192 GNDA.n3060 0.028198
R22224 GNDA.n3188 GNDA.n3059 0.028198
R22225 GNDA.n3178 GNDA.n3057 0.028198
R22226 GNDA.n3172 GNDA.n3056 0.028198
R22227 GNDA.n3162 GNDA.n3054 0.028198
R22228 GNDA.n3158 GNDA.n3053 0.028198
R22229 GNDA.n3148 GNDA.n3051 0.028198
R22230 GNDA.n3142 GNDA.n3050 0.028198
R22231 GNDA.n3132 GNDA.n3048 0.028198
R22232 GNDA.n3128 GNDA.n3047 0.028198
R22233 GNDA.n3118 GNDA.n3045 0.028198
R22234 GNDA.n3112 GNDA.n3044 0.028198
R22235 GNDA.n3102 GNDA.n3042 0.028198
R22236 GNDA.n3098 GNDA.n3041 0.028198
R22237 GNDA.n3088 GNDA.n3039 0.028198
R22238 GNDA.n3038 GNDA.n598 0.028198
R22239 GNDA.n3303 GNDA.n3302 0.028198
R22240 GNDA.n3306 GNDA.n3305 0.028198
R22241 GNDA.n3312 GNDA.n3311 0.028198
R22242 GNDA.n3315 GNDA.n3314 0.028198
R22243 GNDA.n3321 GNDA.n3320 0.028198
R22244 GNDA.n3324 GNDA.n3323 0.028198
R22245 GNDA.n3330 GNDA.n3329 0.028198
R22246 GNDA.n3333 GNDA.n3332 0.028198
R22247 GNDA.n3339 GNDA.n3338 0.028198
R22248 GNDA.n3342 GNDA.n3341 0.028198
R22249 GNDA.n3348 GNDA.n3347 0.028198
R22250 GNDA.n3351 GNDA.n3350 0.028198
R22251 GNDA.n3357 GNDA.n3356 0.028198
R22252 GNDA.n3360 GNDA.n3359 0.028198
R22253 GNDA.n3366 GNDA.n3365 0.028198
R22254 GNDA.n3369 GNDA.n3368 0.028198
R22255 GNDA.n5130 GNDA.n376 0.028198
R22256 GNDA.n5126 GNDA.n375 0.028198
R22257 GNDA.n5116 GNDA.n373 0.028198
R22258 GNDA.n5110 GNDA.n372 0.028198
R22259 GNDA.n5100 GNDA.n370 0.028198
R22260 GNDA.n5096 GNDA.n369 0.028198
R22261 GNDA.n5086 GNDA.n367 0.028198
R22262 GNDA.n5080 GNDA.n366 0.028198
R22263 GNDA.n5070 GNDA.n364 0.028198
R22264 GNDA.n5066 GNDA.n363 0.028198
R22265 GNDA.n5056 GNDA.n361 0.028198
R22266 GNDA.n5050 GNDA.n360 0.028198
R22267 GNDA.n5040 GNDA.n358 0.028198
R22268 GNDA.n5036 GNDA.n357 0.028198
R22269 GNDA.n5026 GNDA.n355 0.028198
R22270 GNDA.n5020 GNDA.n354 0.028198
R22271 GNDA.n500 GNDA.n499 0.028198
R22272 GNDA.n503 GNDA.n502 0.028198
R22273 GNDA.n509 GNDA.n508 0.028198
R22274 GNDA.n512 GNDA.n511 0.028198
R22275 GNDA.n518 GNDA.n517 0.028198
R22276 GNDA.n521 GNDA.n520 0.028198
R22277 GNDA.n527 GNDA.n526 0.028198
R22278 GNDA.n530 GNDA.n529 0.028198
R22279 GNDA.n536 GNDA.n535 0.028198
R22280 GNDA.n539 GNDA.n538 0.028198
R22281 GNDA.n545 GNDA.n544 0.028198
R22282 GNDA.n548 GNDA.n547 0.028198
R22283 GNDA.n554 GNDA.n553 0.028198
R22284 GNDA.n557 GNDA.n556 0.028198
R22285 GNDA.n563 GNDA.n562 0.028198
R22286 GNDA.n566 GNDA.n565 0.028198
R22287 GNDA.n3606 GNDA.n3605 0.028198
R22288 GNDA.n3609 GNDA.n3608 0.028198
R22289 GNDA.n3615 GNDA.n3614 0.028198
R22290 GNDA.n3618 GNDA.n3617 0.028198
R22291 GNDA.n3624 GNDA.n3623 0.028198
R22292 GNDA.n3627 GNDA.n3626 0.028198
R22293 GNDA.n3633 GNDA.n3632 0.028198
R22294 GNDA.n3636 GNDA.n3635 0.028198
R22295 GNDA.n3642 GNDA.n3641 0.028198
R22296 GNDA.n3645 GNDA.n3644 0.028198
R22297 GNDA.n3651 GNDA.n3650 0.028198
R22298 GNDA.n3654 GNDA.n3653 0.028198
R22299 GNDA.n3660 GNDA.n3659 0.028198
R22300 GNDA.n3663 GNDA.n3662 0.028198
R22301 GNDA.n3669 GNDA.n3668 0.028198
R22302 GNDA.n3672 GNDA.n3671 0.028198
R22303 GNDA.n3964 GNDA.n3827 0.028198
R22304 GNDA.n3960 GNDA.n3826 0.028198
R22305 GNDA.n3950 GNDA.n3824 0.028198
R22306 GNDA.n3944 GNDA.n3823 0.028198
R22307 GNDA.n3934 GNDA.n3821 0.028198
R22308 GNDA.n3930 GNDA.n3820 0.028198
R22309 GNDA.n3920 GNDA.n3818 0.028198
R22310 GNDA.n3914 GNDA.n3817 0.028198
R22311 GNDA.n3904 GNDA.n3815 0.028198
R22312 GNDA.n3900 GNDA.n3814 0.028198
R22313 GNDA.n3890 GNDA.n3812 0.028198
R22314 GNDA.n3884 GNDA.n3811 0.028198
R22315 GNDA.n3874 GNDA.n3809 0.028198
R22316 GNDA.n3870 GNDA.n3808 0.028198
R22317 GNDA.n3860 GNDA.n3806 0.028198
R22318 GNDA.n3854 GNDA.n3805 0.028198
R22319 GNDA.n4130 GNDA.n3993 0.028198
R22320 GNDA.n4126 GNDA.n3992 0.028198
R22321 GNDA.n4116 GNDA.n3990 0.028198
R22322 GNDA.n4110 GNDA.n3989 0.028198
R22323 GNDA.n4100 GNDA.n3987 0.028198
R22324 GNDA.n4096 GNDA.n3986 0.028198
R22325 GNDA.n4086 GNDA.n3984 0.028198
R22326 GNDA.n4080 GNDA.n3983 0.028198
R22327 GNDA.n4070 GNDA.n3981 0.028198
R22328 GNDA.n4066 GNDA.n3980 0.028198
R22329 GNDA.n4056 GNDA.n3978 0.028198
R22330 GNDA.n4050 GNDA.n3977 0.028198
R22331 GNDA.n4040 GNDA.n3975 0.028198
R22332 GNDA.n4036 GNDA.n3974 0.028198
R22333 GNDA.n4026 GNDA.n3972 0.028198
R22334 GNDA.n4020 GNDA.n3971 0.028198
R22335 GNDA.n3798 GNDA.n3483 0.028198
R22336 GNDA.n3794 GNDA.n3482 0.028198
R22337 GNDA.n3784 GNDA.n3480 0.028198
R22338 GNDA.n3778 GNDA.n3479 0.028198
R22339 GNDA.n3768 GNDA.n3477 0.028198
R22340 GNDA.n3764 GNDA.n3476 0.028198
R22341 GNDA.n3754 GNDA.n3474 0.028198
R22342 GNDA.n3748 GNDA.n3473 0.028198
R22343 GNDA.n3738 GNDA.n3471 0.028198
R22344 GNDA.n3734 GNDA.n3470 0.028198
R22345 GNDA.n3724 GNDA.n3468 0.028198
R22346 GNDA.n3718 GNDA.n3467 0.028198
R22347 GNDA.n3708 GNDA.n3465 0.028198
R22348 GNDA.n3704 GNDA.n3464 0.028198
R22349 GNDA.n3694 GNDA.n3462 0.028198
R22350 GNDA.n3688 GNDA.n3461 0.028198
R22351 GNDA.n4296 GNDA.n4159 0.028198
R22352 GNDA.n4292 GNDA.n4158 0.028198
R22353 GNDA.n4282 GNDA.n4156 0.028198
R22354 GNDA.n4276 GNDA.n4155 0.028198
R22355 GNDA.n4266 GNDA.n4153 0.028198
R22356 GNDA.n4262 GNDA.n4152 0.028198
R22357 GNDA.n4252 GNDA.n4150 0.028198
R22358 GNDA.n4246 GNDA.n4149 0.028198
R22359 GNDA.n4236 GNDA.n4147 0.028198
R22360 GNDA.n4232 GNDA.n4146 0.028198
R22361 GNDA.n4222 GNDA.n4144 0.028198
R22362 GNDA.n4216 GNDA.n4143 0.028198
R22363 GNDA.n4206 GNDA.n4141 0.028198
R22364 GNDA.n4202 GNDA.n4140 0.028198
R22365 GNDA.n4192 GNDA.n4138 0.028198
R22366 GNDA.n4186 GNDA.n4137 0.028198
R22367 GNDA.n4462 GNDA.n4325 0.028198
R22368 GNDA.n4458 GNDA.n4324 0.028198
R22369 GNDA.n4448 GNDA.n4322 0.028198
R22370 GNDA.n4442 GNDA.n4321 0.028198
R22371 GNDA.n4432 GNDA.n4319 0.028198
R22372 GNDA.n4428 GNDA.n4318 0.028198
R22373 GNDA.n4418 GNDA.n4316 0.028198
R22374 GNDA.n4412 GNDA.n4315 0.028198
R22375 GNDA.n4402 GNDA.n4313 0.028198
R22376 GNDA.n4398 GNDA.n4312 0.028198
R22377 GNDA.n4388 GNDA.n4310 0.028198
R22378 GNDA.n4382 GNDA.n4309 0.028198
R22379 GNDA.n4372 GNDA.n4307 0.028198
R22380 GNDA.n4368 GNDA.n4306 0.028198
R22381 GNDA.n4358 GNDA.n4304 0.028198
R22382 GNDA.n4352 GNDA.n4303 0.028198
R22383 GNDA.n4628 GNDA.n4491 0.028198
R22384 GNDA.n4624 GNDA.n4490 0.028198
R22385 GNDA.n4614 GNDA.n4488 0.028198
R22386 GNDA.n4608 GNDA.n4487 0.028198
R22387 GNDA.n4598 GNDA.n4485 0.028198
R22388 GNDA.n4594 GNDA.n4484 0.028198
R22389 GNDA.n4584 GNDA.n4482 0.028198
R22390 GNDA.n4578 GNDA.n4481 0.028198
R22391 GNDA.n4568 GNDA.n4479 0.028198
R22392 GNDA.n4564 GNDA.n4478 0.028198
R22393 GNDA.n4554 GNDA.n4476 0.028198
R22394 GNDA.n4548 GNDA.n4475 0.028198
R22395 GNDA.n4538 GNDA.n4473 0.028198
R22396 GNDA.n4534 GNDA.n4472 0.028198
R22397 GNDA.n4524 GNDA.n4470 0.028198
R22398 GNDA.n4518 GNDA.n4469 0.028198
R22399 GNDA.n4794 GNDA.n4657 0.028198
R22400 GNDA.n4790 GNDA.n4656 0.028198
R22401 GNDA.n4780 GNDA.n4654 0.028198
R22402 GNDA.n4774 GNDA.n4653 0.028198
R22403 GNDA.n4764 GNDA.n4651 0.028198
R22404 GNDA.n4760 GNDA.n4650 0.028198
R22405 GNDA.n4750 GNDA.n4648 0.028198
R22406 GNDA.n4744 GNDA.n4647 0.028198
R22407 GNDA.n4734 GNDA.n4645 0.028198
R22408 GNDA.n4730 GNDA.n4644 0.028198
R22409 GNDA.n4720 GNDA.n4642 0.028198
R22410 GNDA.n4714 GNDA.n4641 0.028198
R22411 GNDA.n4704 GNDA.n4639 0.028198
R22412 GNDA.n4700 GNDA.n4638 0.028198
R22413 GNDA.n4690 GNDA.n4636 0.028198
R22414 GNDA.n4684 GNDA.n4635 0.028198
R22415 GNDA.n4954 GNDA.n4822 0.028198
R22416 GNDA.n4950 GNDA.n4821 0.028198
R22417 GNDA.n4940 GNDA.n4819 0.028198
R22418 GNDA.n4934 GNDA.n4818 0.028198
R22419 GNDA.n4924 GNDA.n4816 0.028198
R22420 GNDA.n4920 GNDA.n4815 0.028198
R22421 GNDA.n4910 GNDA.n4813 0.028198
R22422 GNDA.n4904 GNDA.n4812 0.028198
R22423 GNDA.n4894 GNDA.n4810 0.028198
R22424 GNDA.n4890 GNDA.n4809 0.028198
R22425 GNDA.n4880 GNDA.n4807 0.028198
R22426 GNDA.n4874 GNDA.n4806 0.028198
R22427 GNDA.n4864 GNDA.n4804 0.028198
R22428 GNDA.n4860 GNDA.n4803 0.028198
R22429 GNDA.n4850 GNDA.n4801 0.028198
R22430 GNDA.n4800 GNDA.n3458 0.028198
R22431 GNDA.n5267 GNDA.n352 0.028198
R22432 GNDA.n5263 GNDA.n351 0.028198
R22433 GNDA.n5253 GNDA.n349 0.028198
R22434 GNDA.n5247 GNDA.n348 0.028198
R22435 GNDA.n5237 GNDA.n346 0.028198
R22436 GNDA.n5233 GNDA.n345 0.028198
R22437 GNDA.n5223 GNDA.n343 0.028198
R22438 GNDA.n5217 GNDA.n342 0.028198
R22439 GNDA.n5207 GNDA.n340 0.028198
R22440 GNDA.n5203 GNDA.n339 0.028198
R22441 GNDA.n5193 GNDA.n337 0.028198
R22442 GNDA.n5187 GNDA.n336 0.028198
R22443 GNDA.n5177 GNDA.n334 0.028198
R22444 GNDA.n5173 GNDA.n333 0.028198
R22445 GNDA.n5163 GNDA.n331 0.028198
R22446 GNDA.n330 GNDA.n328 0.028198
R22447 GNDA.n7136 GNDA.n7067 0.028198
R22448 GNDA.n7129 GNDA.n7068 0.028198
R22449 GNDA.n7125 GNDA.n7070 0.028198
R22450 GNDA.n7152 GNDA.n7071 0.028198
R22451 GNDA.n7160 GNDA.n7073 0.028198
R22452 GNDA.n7117 GNDA.n7074 0.028198
R22453 GNDA.n7113 GNDA.n7076 0.028198
R22454 GNDA.n7176 GNDA.n7077 0.028198
R22455 GNDA.n7184 GNDA.n7079 0.028198
R22456 GNDA.n7105 GNDA.n7080 0.028198
R22457 GNDA.n7101 GNDA.n7082 0.028198
R22458 GNDA.n7200 GNDA.n7083 0.028198
R22459 GNDA.n7208 GNDA.n7085 0.028198
R22460 GNDA.n7093 GNDA.n7086 0.028198
R22461 GNDA.n7089 GNDA.n7088 0.028198
R22462 GNDA.n7224 GNDA.n97 0.028198
R22463 GNDA.n152 GNDA.n100 0.028198
R22464 GNDA.n156 GNDA.n101 0.028198
R22465 GNDA.n166 GNDA.n103 0.028198
R22466 GNDA.n172 GNDA.n104 0.028198
R22467 GNDA.n182 GNDA.n106 0.028198
R22468 GNDA.n186 GNDA.n107 0.028198
R22469 GNDA.n196 GNDA.n109 0.028198
R22470 GNDA.n202 GNDA.n110 0.028198
R22471 GNDA.n212 GNDA.n112 0.028198
R22472 GNDA.n216 GNDA.n113 0.028198
R22473 GNDA.n226 GNDA.n115 0.028198
R22474 GNDA.n232 GNDA.n116 0.028198
R22475 GNDA.n242 GNDA.n118 0.028198
R22476 GNDA.n246 GNDA.n119 0.028198
R22477 GNDA.n256 GNDA.n121 0.028198
R22478 GNDA.n123 GNDA.n122 0.028198
R22479 GNDA.n257 GNDA.n122 0.028198
R22480 GNDA.n253 GNDA.n121 0.028198
R22481 GNDA.n243 GNDA.n119 0.028198
R22482 GNDA.n237 GNDA.n118 0.028198
R22483 GNDA.n227 GNDA.n116 0.028198
R22484 GNDA.n223 GNDA.n115 0.028198
R22485 GNDA.n213 GNDA.n113 0.028198
R22486 GNDA.n207 GNDA.n112 0.028198
R22487 GNDA.n197 GNDA.n110 0.028198
R22488 GNDA.n193 GNDA.n109 0.028198
R22489 GNDA.n183 GNDA.n107 0.028198
R22490 GNDA.n177 GNDA.n106 0.028198
R22491 GNDA.n167 GNDA.n104 0.028198
R22492 GNDA.n163 GNDA.n103 0.028198
R22493 GNDA.n153 GNDA.n101 0.028198
R22494 GNDA.n147 GNDA.n100 0.028198
R22495 GNDA.n7224 GNDA.n7223 0.028198
R22496 GNDA.n7217 GNDA.n7088 0.028198
R22497 GNDA.n7209 GNDA.n7086 0.028198
R22498 GNDA.n7098 GNDA.n7085 0.028198
R22499 GNDA.n7102 GNDA.n7083 0.028198
R22500 GNDA.n7193 GNDA.n7082 0.028198
R22501 GNDA.n7185 GNDA.n7080 0.028198
R22502 GNDA.n7110 GNDA.n7079 0.028198
R22503 GNDA.n7114 GNDA.n7077 0.028198
R22504 GNDA.n7169 GNDA.n7076 0.028198
R22505 GNDA.n7161 GNDA.n7074 0.028198
R22506 GNDA.n7122 GNDA.n7073 0.028198
R22507 GNDA.n7126 GNDA.n7071 0.028198
R22508 GNDA.n7145 GNDA.n7070 0.028198
R22509 GNDA.n7137 GNDA.n7068 0.028198
R22510 GNDA.n7133 GNDA.n7067 0.028198
R22511 GNDA.n1243 GNDA.n1169 0.028198
R22512 GNDA.n1255 GNDA.n1172 0.028198
R22513 GNDA.n1273 GNDA.n1175 0.028198
R22514 GNDA.n1285 GNDA.n1178 0.028198
R22515 GNDA.n1303 GNDA.n1181 0.028198
R22516 GNDA.n1315 GNDA.n1184 0.028198
R22517 GNDA.n1333 GNDA.n1187 0.028198
R22518 GNDA.n1353 GNDA.n1190 0.028198
R22519 GNDA.n1353 GNDA.n1352 0.028198
R22520 GNDA.n1336 GNDA.n1187 0.028198
R22521 GNDA.n1322 GNDA.n1184 0.028198
R22522 GNDA.n1306 GNDA.n1181 0.028198
R22523 GNDA.n1292 GNDA.n1178 0.028198
R22524 GNDA.n1276 GNDA.n1175 0.028198
R22525 GNDA.n1262 GNDA.n1172 0.028198
R22526 GNDA.n1246 GNDA.n1169 0.028198
R22527 GNDA.n1245 GNDA.n1170 0.0262697
R22528 GNDA.n1253 GNDA.n1171 0.0262697
R22529 GNDA.n1263 GNDA.n1173 0.0262697
R22530 GNDA.n1265 GNDA.n1174 0.0262697
R22531 GNDA.n1275 GNDA.n1176 0.0262697
R22532 GNDA.n1283 GNDA.n1177 0.0262697
R22533 GNDA.n1293 GNDA.n1179 0.0262697
R22534 GNDA.n1295 GNDA.n1180 0.0262697
R22535 GNDA.n1305 GNDA.n1182 0.0262697
R22536 GNDA.n1313 GNDA.n1183 0.0262697
R22537 GNDA.n1323 GNDA.n1185 0.0262697
R22538 GNDA.n1325 GNDA.n1186 0.0262697
R22539 GNDA.n1335 GNDA.n1188 0.0262697
R22540 GNDA.n1343 GNDA.n1189 0.0262697
R22541 GNDA.n1191 GNDA.n1167 0.0262697
R22542 GNDA.n1345 GNDA.n1189 0.0262697
R22543 GNDA.n1342 GNDA.n1188 0.0262697
R22544 GNDA.n1332 GNDA.n1186 0.0262697
R22545 GNDA.n1326 GNDA.n1185 0.0262697
R22546 GNDA.n1316 GNDA.n1183 0.0262697
R22547 GNDA.n1312 GNDA.n1182 0.0262697
R22548 GNDA.n1302 GNDA.n1180 0.0262697
R22549 GNDA.n1296 GNDA.n1179 0.0262697
R22550 GNDA.n1286 GNDA.n1177 0.0262697
R22551 GNDA.n1282 GNDA.n1176 0.0262697
R22552 GNDA.n1272 GNDA.n1174 0.0262697
R22553 GNDA.n1266 GNDA.n1173 0.0262697
R22554 GNDA.n1256 GNDA.n1171 0.0262697
R22555 GNDA.n1252 GNDA.n1170 0.0262697
R22556 GNDA.n1242 GNDA.n1168 0.0262697
R22557 GNDA.n5172 GNDA.n332 0.0243392
R22558 GNDA.n5186 GNDA.n335 0.0243392
R22559 GNDA.n5202 GNDA.n338 0.0243392
R22560 GNDA.n5216 GNDA.n341 0.0243392
R22561 GNDA.n5232 GNDA.n344 0.0243392
R22562 GNDA.n5246 GNDA.n347 0.0243392
R22563 GNDA.n5262 GNDA.n350 0.0243392
R22564 GNDA.n4859 GNDA.n4802 0.0243392
R22565 GNDA.n4873 GNDA.n4805 0.0243392
R22566 GNDA.n4889 GNDA.n4808 0.0243392
R22567 GNDA.n4903 GNDA.n4811 0.0243392
R22568 GNDA.n4919 GNDA.n4814 0.0243392
R22569 GNDA.n4933 GNDA.n4817 0.0243392
R22570 GNDA.n4949 GNDA.n4820 0.0243392
R22571 GNDA.n4699 GNDA.n4637 0.0243392
R22572 GNDA.n4713 GNDA.n4640 0.0243392
R22573 GNDA.n4729 GNDA.n4643 0.0243392
R22574 GNDA.n4743 GNDA.n4646 0.0243392
R22575 GNDA.n4759 GNDA.n4649 0.0243392
R22576 GNDA.n4773 GNDA.n4652 0.0243392
R22577 GNDA.n4789 GNDA.n4655 0.0243392
R22578 GNDA.n4533 GNDA.n4471 0.0243392
R22579 GNDA.n4547 GNDA.n4474 0.0243392
R22580 GNDA.n4563 GNDA.n4477 0.0243392
R22581 GNDA.n4577 GNDA.n4480 0.0243392
R22582 GNDA.n4593 GNDA.n4483 0.0243392
R22583 GNDA.n4607 GNDA.n4486 0.0243392
R22584 GNDA.n4623 GNDA.n4489 0.0243392
R22585 GNDA.n4367 GNDA.n4305 0.0243392
R22586 GNDA.n4381 GNDA.n4308 0.0243392
R22587 GNDA.n4397 GNDA.n4311 0.0243392
R22588 GNDA.n4411 GNDA.n4314 0.0243392
R22589 GNDA.n4427 GNDA.n4317 0.0243392
R22590 GNDA.n4441 GNDA.n4320 0.0243392
R22591 GNDA.n4457 GNDA.n4323 0.0243392
R22592 GNDA.n4201 GNDA.n4139 0.0243392
R22593 GNDA.n4215 GNDA.n4142 0.0243392
R22594 GNDA.n4231 GNDA.n4145 0.0243392
R22595 GNDA.n4245 GNDA.n4148 0.0243392
R22596 GNDA.n4261 GNDA.n4151 0.0243392
R22597 GNDA.n4275 GNDA.n4154 0.0243392
R22598 GNDA.n4291 GNDA.n4157 0.0243392
R22599 GNDA.n3703 GNDA.n3463 0.0243392
R22600 GNDA.n3717 GNDA.n3466 0.0243392
R22601 GNDA.n3733 GNDA.n3469 0.0243392
R22602 GNDA.n3747 GNDA.n3472 0.0243392
R22603 GNDA.n3763 GNDA.n3475 0.0243392
R22604 GNDA.n3777 GNDA.n3478 0.0243392
R22605 GNDA.n3793 GNDA.n3481 0.0243392
R22606 GNDA.n4035 GNDA.n3973 0.0243392
R22607 GNDA.n4049 GNDA.n3976 0.0243392
R22608 GNDA.n4065 GNDA.n3979 0.0243392
R22609 GNDA.n4079 GNDA.n3982 0.0243392
R22610 GNDA.n4095 GNDA.n3985 0.0243392
R22611 GNDA.n4109 GNDA.n3988 0.0243392
R22612 GNDA.n4125 GNDA.n3991 0.0243392
R22613 GNDA.n3869 GNDA.n3807 0.0243392
R22614 GNDA.n3883 GNDA.n3810 0.0243392
R22615 GNDA.n3899 GNDA.n3813 0.0243392
R22616 GNDA.n3913 GNDA.n3816 0.0243392
R22617 GNDA.n3929 GNDA.n3819 0.0243392
R22618 GNDA.n3943 GNDA.n3822 0.0243392
R22619 GNDA.n3959 GNDA.n3825 0.0243392
R22620 GNDA.n3665 GNDA.n3664 0.0243392
R22621 GNDA.n3656 GNDA.n3655 0.0243392
R22622 GNDA.n3647 GNDA.n3646 0.0243392
R22623 GNDA.n3638 GNDA.n3637 0.0243392
R22624 GNDA.n3629 GNDA.n3628 0.0243392
R22625 GNDA.n3620 GNDA.n3619 0.0243392
R22626 GNDA.n3611 GNDA.n3610 0.0243392
R22627 GNDA.n559 GNDA.n558 0.0243392
R22628 GNDA.n550 GNDA.n549 0.0243392
R22629 GNDA.n541 GNDA.n540 0.0243392
R22630 GNDA.n532 GNDA.n531 0.0243392
R22631 GNDA.n523 GNDA.n522 0.0243392
R22632 GNDA.n514 GNDA.n513 0.0243392
R22633 GNDA.n505 GNDA.n504 0.0243392
R22634 GNDA.n5035 GNDA.n356 0.0243392
R22635 GNDA.n5049 GNDA.n359 0.0243392
R22636 GNDA.n5065 GNDA.n362 0.0243392
R22637 GNDA.n5079 GNDA.n365 0.0243392
R22638 GNDA.n5095 GNDA.n368 0.0243392
R22639 GNDA.n5109 GNDA.n371 0.0243392
R22640 GNDA.n5125 GNDA.n374 0.0243392
R22641 GNDA.n3362 GNDA.n3361 0.0243392
R22642 GNDA.n3353 GNDA.n3352 0.0243392
R22643 GNDA.n3344 GNDA.n3343 0.0243392
R22644 GNDA.n3335 GNDA.n3334 0.0243392
R22645 GNDA.n3326 GNDA.n3325 0.0243392
R22646 GNDA.n3317 GNDA.n3316 0.0243392
R22647 GNDA.n3308 GNDA.n3307 0.0243392
R22648 GNDA.n3097 GNDA.n3040 0.0243392
R22649 GNDA.n3111 GNDA.n3043 0.0243392
R22650 GNDA.n3127 GNDA.n3046 0.0243392
R22651 GNDA.n3141 GNDA.n3049 0.0243392
R22652 GNDA.n3157 GNDA.n3052 0.0243392
R22653 GNDA.n3171 GNDA.n3055 0.0243392
R22654 GNDA.n3187 GNDA.n3058 0.0243392
R22655 GNDA.n2937 GNDA.n2867 0.0243392
R22656 GNDA.n2951 GNDA.n2870 0.0243392
R22657 GNDA.n2967 GNDA.n2873 0.0243392
R22658 GNDA.n2981 GNDA.n2876 0.0243392
R22659 GNDA.n2997 GNDA.n2879 0.0243392
R22660 GNDA.n3011 GNDA.n2882 0.0243392
R22661 GNDA.n3027 GNDA.n2885 0.0243392
R22662 GNDA.n2301 GNDA.n669 0.0243392
R22663 GNDA.n2315 GNDA.n672 0.0243392
R22664 GNDA.n2331 GNDA.n675 0.0243392
R22665 GNDA.n2345 GNDA.n678 0.0243392
R22666 GNDA.n2361 GNDA.n681 0.0243392
R22667 GNDA.n2375 GNDA.n684 0.0243392
R22668 GNDA.n2391 GNDA.n687 0.0243392
R22669 GNDA.n2763 GNDA.n603 0.0243392
R22670 GNDA.n2777 GNDA.n606 0.0243392
R22671 GNDA.n2793 GNDA.n609 0.0243392
R22672 GNDA.n2807 GNDA.n612 0.0243392
R22673 GNDA.n2823 GNDA.n615 0.0243392
R22674 GNDA.n2837 GNDA.n618 0.0243392
R22675 GNDA.n2853 GNDA.n621 0.0243392
R22676 GNDA.n2725 GNDA.n2724 0.0243392
R22677 GNDA.n2716 GNDA.n2715 0.0243392
R22678 GNDA.n2707 GNDA.n2706 0.0243392
R22679 GNDA.n2698 GNDA.n2697 0.0243392
R22680 GNDA.n2689 GNDA.n2688 0.0243392
R22681 GNDA.n2680 GNDA.n2679 0.0243392
R22682 GNDA.n2671 GNDA.n2670 0.0243392
R22683 GNDA.n2461 GNDA.n2404 0.0243392
R22684 GNDA.n2475 GNDA.n2407 0.0243392
R22685 GNDA.n2491 GNDA.n2410 0.0243392
R22686 GNDA.n2505 GNDA.n2413 0.0243392
R22687 GNDA.n2521 GNDA.n2416 0.0243392
R22688 GNDA.n2535 GNDA.n2419 0.0243392
R22689 GNDA.n2551 GNDA.n2422 0.0243392
R22690 GNDA.n2265 GNDA.n2264 0.0243392
R22691 GNDA.n2256 GNDA.n2255 0.0243392
R22692 GNDA.n2247 GNDA.n2246 0.0243392
R22693 GNDA.n2238 GNDA.n2237 0.0243392
R22694 GNDA.n2229 GNDA.n2228 0.0243392
R22695 GNDA.n2220 GNDA.n2219 0.0243392
R22696 GNDA.n2211 GNDA.n2210 0.0243392
R22697 GNDA.n1998 GNDA.n1941 0.0243392
R22698 GNDA.n2012 GNDA.n1944 0.0243392
R22699 GNDA.n2028 GNDA.n1947 0.0243392
R22700 GNDA.n2042 GNDA.n1950 0.0243392
R22701 GNDA.n2058 GNDA.n1953 0.0243392
R22702 GNDA.n2072 GNDA.n1956 0.0243392
R22703 GNDA.n2088 GNDA.n1959 0.0243392
R22704 GNDA.n1838 GNDA.n732 0.0243392
R22705 GNDA.n1852 GNDA.n735 0.0243392
R22706 GNDA.n1868 GNDA.n738 0.0243392
R22707 GNDA.n1882 GNDA.n741 0.0243392
R22708 GNDA.n1898 GNDA.n744 0.0243392
R22709 GNDA.n1912 GNDA.n747 0.0243392
R22710 GNDA.n1928 GNDA.n750 0.0243392
R22711 GNDA.n1678 GNDA.n1677 0.0243392
R22712 GNDA.n1669 GNDA.n1668 0.0243392
R22713 GNDA.n1660 GNDA.n1659 0.0243392
R22714 GNDA.n1651 GNDA.n1650 0.0243392
R22715 GNDA.n1642 GNDA.n1641 0.0243392
R22716 GNDA.n1633 GNDA.n1632 0.0243392
R22717 GNDA.n1624 GNDA.n1623 0.0243392
R22718 GNDA.n1414 GNDA.n1357 0.0243392
R22719 GNDA.n1428 GNDA.n1360 0.0243392
R22720 GNDA.n1444 GNDA.n1363 0.0243392
R22721 GNDA.n1458 GNDA.n1366 0.0243392
R22722 GNDA.n1474 GNDA.n1369 0.0243392
R22723 GNDA.n1488 GNDA.n1372 0.0243392
R22724 GNDA.n1504 GNDA.n1375 0.0243392
R22725 GNDA.n1499 GNDA.n1375 0.0243392
R22726 GNDA.n1485 GNDA.n1372 0.0243392
R22727 GNDA.n1469 GNDA.n1369 0.0243392
R22728 GNDA.n1455 GNDA.n1366 0.0243392
R22729 GNDA.n1439 GNDA.n1363 0.0243392
R22730 GNDA.n1425 GNDA.n1360 0.0243392
R22731 GNDA.n1409 GNDA.n1357 0.0243392
R22732 GNDA.n1625 GNDA.n1624 0.0243392
R22733 GNDA.n1634 GNDA.n1633 0.0243392
R22734 GNDA.n1643 GNDA.n1642 0.0243392
R22735 GNDA.n1652 GNDA.n1651 0.0243392
R22736 GNDA.n1661 GNDA.n1660 0.0243392
R22737 GNDA.n1670 GNDA.n1669 0.0243392
R22738 GNDA.n1679 GNDA.n1678 0.0243392
R22739 GNDA.n1923 GNDA.n750 0.0243392
R22740 GNDA.n1909 GNDA.n747 0.0243392
R22741 GNDA.n1893 GNDA.n744 0.0243392
R22742 GNDA.n1879 GNDA.n741 0.0243392
R22743 GNDA.n1863 GNDA.n738 0.0243392
R22744 GNDA.n1849 GNDA.n735 0.0243392
R22745 GNDA.n1833 GNDA.n732 0.0243392
R22746 GNDA.n2083 GNDA.n1959 0.0243392
R22747 GNDA.n2069 GNDA.n1956 0.0243392
R22748 GNDA.n2053 GNDA.n1953 0.0243392
R22749 GNDA.n2039 GNDA.n1950 0.0243392
R22750 GNDA.n2023 GNDA.n1947 0.0243392
R22751 GNDA.n2009 GNDA.n1944 0.0243392
R22752 GNDA.n1993 GNDA.n1941 0.0243392
R22753 GNDA.n2212 GNDA.n2211 0.0243392
R22754 GNDA.n2221 GNDA.n2220 0.0243392
R22755 GNDA.n2230 GNDA.n2229 0.0243392
R22756 GNDA.n2239 GNDA.n2238 0.0243392
R22757 GNDA.n2248 GNDA.n2247 0.0243392
R22758 GNDA.n2257 GNDA.n2256 0.0243392
R22759 GNDA.n2266 GNDA.n2265 0.0243392
R22760 GNDA.n2546 GNDA.n2422 0.0243392
R22761 GNDA.n2532 GNDA.n2419 0.0243392
R22762 GNDA.n2516 GNDA.n2416 0.0243392
R22763 GNDA.n2502 GNDA.n2413 0.0243392
R22764 GNDA.n2486 GNDA.n2410 0.0243392
R22765 GNDA.n2472 GNDA.n2407 0.0243392
R22766 GNDA.n2456 GNDA.n2404 0.0243392
R22767 GNDA.n2672 GNDA.n2671 0.0243392
R22768 GNDA.n2681 GNDA.n2680 0.0243392
R22769 GNDA.n2690 GNDA.n2689 0.0243392
R22770 GNDA.n2699 GNDA.n2698 0.0243392
R22771 GNDA.n2708 GNDA.n2707 0.0243392
R22772 GNDA.n2717 GNDA.n2716 0.0243392
R22773 GNDA.n2726 GNDA.n2725 0.0243392
R22774 GNDA.n2848 GNDA.n621 0.0243392
R22775 GNDA.n2834 GNDA.n618 0.0243392
R22776 GNDA.n2818 GNDA.n615 0.0243392
R22777 GNDA.n2804 GNDA.n612 0.0243392
R22778 GNDA.n2788 GNDA.n609 0.0243392
R22779 GNDA.n2774 GNDA.n606 0.0243392
R22780 GNDA.n2758 GNDA.n603 0.0243392
R22781 GNDA.n2386 GNDA.n687 0.0243392
R22782 GNDA.n2372 GNDA.n684 0.0243392
R22783 GNDA.n2356 GNDA.n681 0.0243392
R22784 GNDA.n2342 GNDA.n678 0.0243392
R22785 GNDA.n2326 GNDA.n675 0.0243392
R22786 GNDA.n2312 GNDA.n672 0.0243392
R22787 GNDA.n2296 GNDA.n669 0.0243392
R22788 GNDA.n3022 GNDA.n2885 0.0243392
R22789 GNDA.n3008 GNDA.n2882 0.0243392
R22790 GNDA.n2992 GNDA.n2879 0.0243392
R22791 GNDA.n2978 GNDA.n2876 0.0243392
R22792 GNDA.n2962 GNDA.n2873 0.0243392
R22793 GNDA.n2948 GNDA.n2870 0.0243392
R22794 GNDA.n2932 GNDA.n2867 0.0243392
R22795 GNDA.n3182 GNDA.n3058 0.0243392
R22796 GNDA.n3168 GNDA.n3055 0.0243392
R22797 GNDA.n3152 GNDA.n3052 0.0243392
R22798 GNDA.n3138 GNDA.n3049 0.0243392
R22799 GNDA.n3122 GNDA.n3046 0.0243392
R22800 GNDA.n3108 GNDA.n3043 0.0243392
R22801 GNDA.n3092 GNDA.n3040 0.0243392
R22802 GNDA.n3309 GNDA.n3308 0.0243392
R22803 GNDA.n3318 GNDA.n3317 0.0243392
R22804 GNDA.n3327 GNDA.n3326 0.0243392
R22805 GNDA.n3336 GNDA.n3335 0.0243392
R22806 GNDA.n3345 GNDA.n3344 0.0243392
R22807 GNDA.n3354 GNDA.n3353 0.0243392
R22808 GNDA.n3363 GNDA.n3362 0.0243392
R22809 GNDA.n5120 GNDA.n374 0.0243392
R22810 GNDA.n5106 GNDA.n371 0.0243392
R22811 GNDA.n5090 GNDA.n368 0.0243392
R22812 GNDA.n5076 GNDA.n365 0.0243392
R22813 GNDA.n5060 GNDA.n362 0.0243392
R22814 GNDA.n5046 GNDA.n359 0.0243392
R22815 GNDA.n5030 GNDA.n356 0.0243392
R22816 GNDA.n506 GNDA.n505 0.0243392
R22817 GNDA.n515 GNDA.n514 0.0243392
R22818 GNDA.n524 GNDA.n523 0.0243392
R22819 GNDA.n533 GNDA.n532 0.0243392
R22820 GNDA.n542 GNDA.n541 0.0243392
R22821 GNDA.n551 GNDA.n550 0.0243392
R22822 GNDA.n560 GNDA.n559 0.0243392
R22823 GNDA.n3612 GNDA.n3611 0.0243392
R22824 GNDA.n3621 GNDA.n3620 0.0243392
R22825 GNDA.n3630 GNDA.n3629 0.0243392
R22826 GNDA.n3639 GNDA.n3638 0.0243392
R22827 GNDA.n3648 GNDA.n3647 0.0243392
R22828 GNDA.n3657 GNDA.n3656 0.0243392
R22829 GNDA.n3666 GNDA.n3665 0.0243392
R22830 GNDA.n3954 GNDA.n3825 0.0243392
R22831 GNDA.n3940 GNDA.n3822 0.0243392
R22832 GNDA.n3924 GNDA.n3819 0.0243392
R22833 GNDA.n3910 GNDA.n3816 0.0243392
R22834 GNDA.n3894 GNDA.n3813 0.0243392
R22835 GNDA.n3880 GNDA.n3810 0.0243392
R22836 GNDA.n3864 GNDA.n3807 0.0243392
R22837 GNDA.n4120 GNDA.n3991 0.0243392
R22838 GNDA.n4106 GNDA.n3988 0.0243392
R22839 GNDA.n4090 GNDA.n3985 0.0243392
R22840 GNDA.n4076 GNDA.n3982 0.0243392
R22841 GNDA.n4060 GNDA.n3979 0.0243392
R22842 GNDA.n4046 GNDA.n3976 0.0243392
R22843 GNDA.n4030 GNDA.n3973 0.0243392
R22844 GNDA.n3788 GNDA.n3481 0.0243392
R22845 GNDA.n3774 GNDA.n3478 0.0243392
R22846 GNDA.n3758 GNDA.n3475 0.0243392
R22847 GNDA.n3744 GNDA.n3472 0.0243392
R22848 GNDA.n3728 GNDA.n3469 0.0243392
R22849 GNDA.n3714 GNDA.n3466 0.0243392
R22850 GNDA.n3698 GNDA.n3463 0.0243392
R22851 GNDA.n4286 GNDA.n4157 0.0243392
R22852 GNDA.n4272 GNDA.n4154 0.0243392
R22853 GNDA.n4256 GNDA.n4151 0.0243392
R22854 GNDA.n4242 GNDA.n4148 0.0243392
R22855 GNDA.n4226 GNDA.n4145 0.0243392
R22856 GNDA.n4212 GNDA.n4142 0.0243392
R22857 GNDA.n4196 GNDA.n4139 0.0243392
R22858 GNDA.n4452 GNDA.n4323 0.0243392
R22859 GNDA.n4438 GNDA.n4320 0.0243392
R22860 GNDA.n4422 GNDA.n4317 0.0243392
R22861 GNDA.n4408 GNDA.n4314 0.0243392
R22862 GNDA.n4392 GNDA.n4311 0.0243392
R22863 GNDA.n4378 GNDA.n4308 0.0243392
R22864 GNDA.n4362 GNDA.n4305 0.0243392
R22865 GNDA.n4618 GNDA.n4489 0.0243392
R22866 GNDA.n4604 GNDA.n4486 0.0243392
R22867 GNDA.n4588 GNDA.n4483 0.0243392
R22868 GNDA.n4574 GNDA.n4480 0.0243392
R22869 GNDA.n4558 GNDA.n4477 0.0243392
R22870 GNDA.n4544 GNDA.n4474 0.0243392
R22871 GNDA.n4528 GNDA.n4471 0.0243392
R22872 GNDA.n4784 GNDA.n4655 0.0243392
R22873 GNDA.n4770 GNDA.n4652 0.0243392
R22874 GNDA.n4754 GNDA.n4649 0.0243392
R22875 GNDA.n4740 GNDA.n4646 0.0243392
R22876 GNDA.n4724 GNDA.n4643 0.0243392
R22877 GNDA.n4710 GNDA.n4640 0.0243392
R22878 GNDA.n4694 GNDA.n4637 0.0243392
R22879 GNDA.n4944 GNDA.n4820 0.0243392
R22880 GNDA.n4930 GNDA.n4817 0.0243392
R22881 GNDA.n4914 GNDA.n4814 0.0243392
R22882 GNDA.n4900 GNDA.n4811 0.0243392
R22883 GNDA.n4884 GNDA.n4808 0.0243392
R22884 GNDA.n4870 GNDA.n4805 0.0243392
R22885 GNDA.n4854 GNDA.n4802 0.0243392
R22886 GNDA.n5257 GNDA.n350 0.0243392
R22887 GNDA.n5243 GNDA.n347 0.0243392
R22888 GNDA.n5227 GNDA.n344 0.0243392
R22889 GNDA.n5213 GNDA.n341 0.0243392
R22890 GNDA.n5197 GNDA.n338 0.0243392
R22891 GNDA.n5183 GNDA.n335 0.0243392
R22892 GNDA.n5167 GNDA.n332 0.0243392
R22893 GNDA.n7144 GNDA.n7069 0.0243392
R22894 GNDA.n7121 GNDA.n7072 0.0243392
R22895 GNDA.n7168 GNDA.n7075 0.0243392
R22896 GNDA.n7109 GNDA.n7078 0.0243392
R22897 GNDA.n7192 GNDA.n7081 0.0243392
R22898 GNDA.n7097 GNDA.n7084 0.0243392
R22899 GNDA.n7216 GNDA.n7087 0.0243392
R22900 GNDA.n162 GNDA.n102 0.0243392
R22901 GNDA.n176 GNDA.n105 0.0243392
R22902 GNDA.n192 GNDA.n108 0.0243392
R22903 GNDA.n206 GNDA.n111 0.0243392
R22904 GNDA.n222 GNDA.n114 0.0243392
R22905 GNDA.n236 GNDA.n117 0.0243392
R22906 GNDA.n252 GNDA.n120 0.0243392
R22907 GNDA.n247 GNDA.n120 0.0243392
R22908 GNDA.n233 GNDA.n117 0.0243392
R22909 GNDA.n217 GNDA.n114 0.0243392
R22910 GNDA.n203 GNDA.n111 0.0243392
R22911 GNDA.n187 GNDA.n108 0.0243392
R22912 GNDA.n173 GNDA.n105 0.0243392
R22913 GNDA.n157 GNDA.n102 0.0243392
R22914 GNDA.n7094 GNDA.n7087 0.0243392
R22915 GNDA.n7201 GNDA.n7084 0.0243392
R22916 GNDA.n7106 GNDA.n7081 0.0243392
R22917 GNDA.n7177 GNDA.n7078 0.0243392
R22918 GNDA.n7118 GNDA.n7075 0.0243392
R22919 GNDA.n7153 GNDA.n7072 0.0243392
R22920 GNDA.n7130 GNDA.n7069 0.0243392
R22921 GNDA.n3424 GNDA.n3423 0.0217373
R22922 GNDA.n3427 GNDA.n3426 0.0217373
R22923 GNDA.n3430 GNDA.n588 0.0217373
R22924 GNDA.n3433 GNDA.n587 0.0217373
R22925 GNDA.n3432 GNDA.n587 0.0217373
R22926 GNDA.n3422 GNDA.n3407 0.0217373
R22927 GNDA.n3425 GNDA.n3424 0.0217373
R22928 GNDA.n1695 GNDA.n317 0.0217373
R22929 GNDA.n3426 GNDA.n3405 0.0217373
R22930 GNDA.n3405 GNDA.n588 0.0217373
R22931 GNDA.n1719 GNDA.n1718 0.0217373
R22932 GNDA.n1770 GNDA.n1710 0.0217373
R22933 GNDA.n1762 GNDA.n1712 0.0217373
R22934 GNDA.n1758 GNDA.n1715 0.0217373
R22935 GNDA.n1764 GNDA.n1713 0.0217373
R22936 GNDA.n1763 GNDA.n1762 0.0217373
R22937 GNDA.n1759 GNDA.n1716 0.0217373
R22938 GNDA.n1776 GNDA.n1704 0.0217373
R22939 GNDA.n1768 GNDA.n1708 0.0217373
R22940 GNDA.n1710 GNDA.n1708 0.0217373
R22941 GNDA.n1780 GNDA.n1779 0.0217373
R22942 GNDA.n1783 GNDA.n1782 0.0217373
R22943 GNDA.n1785 GNDA.n1701 0.0217373
R22944 GNDA.n1722 GNDA.n1720 0.0217373
R22945 GNDA.n1723 GNDA.n1722 0.0217373
R22946 GNDA.n1778 GNDA.n1704 0.0217373
R22947 GNDA.n1781 GNDA.n1780 0.0217373
R22948 GNDA.n1720 GNDA.n1702 0.0217373
R22949 GNDA.n1721 GNDA.n1719 0.0217373
R22950 GNDA.n1799 GNDA.n1697 0.0217373
R22951 GNDA.n1783 GNDA.n1699 0.0217373
R22952 GNDA.n1701 GNDA.n1699 0.0217373
R22953 GNDA.n1803 GNDA.n1802 0.0217373
R22954 GNDA.n1809 GNDA.n1808 0.0217373
R22955 GNDA.n1811 GNDA.n781 0.0217373
R22956 GNDA.n1814 GNDA.n782 0.0217373
R22957 GNDA.n1801 GNDA.n1697 0.0217373
R22958 GNDA.n1804 GNDA.n1803 0.0217373
R22959 GNDA.n1807 GNDA.n1695 0.0217373
R22960 GNDA.n1810 GNDA.n1809 0.0217373
R22961 GNDA.n325 GNDA.n322 0.0217373
R22962 GNDA.n5276 GNDA.n325 0.0217373
R22963 GNDA.n4964 GNDA.n3454 0.0217373
R22964 GNDA.n4965 GNDA.n3454 0.0217373
R22965 GNDA.n3452 GNDA.n3449 0.0217373
R22966 GNDA.n3453 GNDA.n3449 0.0217373
R22967 GNDA.n3447 GNDA.n3444 0.0217373
R22968 GNDA.n3448 GNDA.n3444 0.0217373
R22969 GNDA.n3442 GNDA.n3439 0.0217373
R22970 GNDA.n3443 GNDA.n3439 0.0217373
R22971 GNDA.n3437 GNDA.n3434 0.0217373
R22972 GNDA.n3438 GNDA.n3434 0.0217373
R22973 GNDA.n585 GNDA.n582 0.0217373
R22974 GNDA.n586 GNDA.n582 0.0217373
R22975 GNDA.n580 GNDA.n577 0.0217373
R22976 GNDA.n581 GNDA.n577 0.0217373
R22977 GNDA.n571 GNDA.n403 0.0217373
R22978 GNDA.n572 GNDA.n403 0.0217373
R22979 GNDA.n5015 GNDA.n5012 0.0217373
R22980 GNDA.n5016 GNDA.n5015 0.0217373
R22981 GNDA.n3374 GNDA.n3206 0.0217373
R22982 GNDA.n3375 GNDA.n3206 0.0217373
R22983 GNDA.n595 GNDA.n593 0.0217373
R22984 GNDA.n595 GNDA.n592 0.0217373
R22985 GNDA.n2917 GNDA.n2914 0.0217373
R22986 GNDA.n2918 GNDA.n2917 0.0217373
R22987 GNDA.n2743 GNDA.n651 0.0217373
R22988 GNDA.n2744 GNDA.n2743 0.0217373
R22989 GNDA.n2570 GNDA.n654 0.0217373
R22990 GNDA.n2570 GNDA.n653 0.0217373
R22991 GNDA.n661 GNDA.n657 0.0217373
R22992 GNDA.n661 GNDA.n656 0.0217373
R22993 GNDA.n724 GNDA.n722 0.0217373
R22994 GNDA.n724 GNDA.n721 0.0217373
R22995 GNDA.n1818 GNDA.n779 0.0217373
R22996 GNDA.n1819 GNDA.n1818 0.0217373
R22997 GNDA.n1523 GNDA.n785 0.0217373
R22998 GNDA.n1523 GNDA.n784 0.0217373
R22999 GNDA.n790 GNDA.n788 0.0217373
R23000 GNDA.n790 GNDA.n787 0.0217373
R23001 GNDA.n1238 GNDA.n1216 0.0217373
R23002 GNDA.n1231 GNDA.n1219 0.0217373
R23003 GNDA.n1226 GNDA.n1222 0.0217373
R23004 GNDA.n1519 GNDA.n786 0.0217373
R23005 GNDA.n1690 GNDA.n783 0.0217373
R23006 GNDA.n778 GNDA.n777 0.0217373
R23007 GNDA.n2103 GNDA.n720 0.0217373
R23008 GNDA.n2277 GNDA.n716 0.0217373
R23009 GNDA.n2566 GNDA.n655 0.0217373
R23010 GNDA.n2737 GNDA.n652 0.0217373
R23011 GNDA.n650 GNDA.n648 0.0217373
R23012 GNDA.n2913 GNDA.n2912 0.0217373
R23013 GNDA.n3202 GNDA.n591 0.0217373
R23014 GNDA.n3378 GNDA.n3377 0.0217373
R23015 GNDA.n5279 GNDA.n5278 0.0217373
R23016 GNDA.n5011 GNDA.n402 0.0217373
R23017 GNDA.n5008 GNDA.n5007 0.0217373
R23018 GNDA.n3509 GNDA.n3508 0.0217373
R23019 GNDA.n4996 GNDA.n4995 0.0217373
R23020 GNDA.n4992 GNDA.n4991 0.0217373
R23021 GNDA.n4988 GNDA.n4987 0.0217373
R23022 GNDA.n4984 GNDA.n4983 0.0217373
R23023 GNDA.n4980 GNDA.n4979 0.0217373
R23024 GNDA.n4976 GNDA.n4975 0.0217373
R23025 GNDA.n4972 GNDA.n4971 0.0217373
R23026 GNDA.n4968 GNDA.n4967 0.0217373
R23027 GNDA.n1223 GNDA.n1221 0.0217373
R23028 GNDA.n1223 GNDA.n1222 0.0217373
R23029 GNDA.n1228 GNDA.n1218 0.0217373
R23030 GNDA.n1228 GNDA.n1219 0.0217373
R23031 GNDA.n1235 GNDA.n1233 0.0217373
R23032 GNDA.n1233 GNDA.n1216 0.0217373
R23033 GNDA.n1521 GNDA.n788 0.0217373
R23034 GNDA.n1518 GNDA.n787 0.0217373
R23035 GNDA.n1520 GNDA.n1519 0.0217373
R23036 GNDA.n1692 GNDA.n785 0.0217373
R23037 GNDA.n1689 GNDA.n784 0.0217373
R23038 GNDA.n1691 GNDA.n1690 0.0217373
R23039 GNDA.n1816 GNDA.n779 0.0217373
R23040 GNDA.n1820 GNDA.n1819 0.0217373
R23041 GNDA.n1817 GNDA.n777 0.0217373
R23042 GNDA.n2105 GNDA.n722 0.0217373
R23043 GNDA.n2102 GNDA.n721 0.0217373
R23044 GNDA.n2104 GNDA.n2103 0.0217373
R23045 GNDA.n2278 GNDA.n2277 0.0217373
R23046 GNDA.n2568 GNDA.n657 0.0217373
R23047 GNDA.n2565 GNDA.n656 0.0217373
R23048 GNDA.n2567 GNDA.n2566 0.0217373
R23049 GNDA.n2739 GNDA.n654 0.0217373
R23050 GNDA.n2736 GNDA.n653 0.0217373
R23051 GNDA.n2738 GNDA.n2737 0.0217373
R23052 GNDA.n2741 GNDA.n651 0.0217373
R23053 GNDA.n2745 GNDA.n2744 0.0217373
R23054 GNDA.n2742 GNDA.n648 0.0217373
R23055 GNDA.n2915 GNDA.n2914 0.0217373
R23056 GNDA.n2919 GNDA.n2918 0.0217373
R23057 GNDA.n2916 GNDA.n2912 0.0217373
R23058 GNDA.n3204 GNDA.n593 0.0217373
R23059 GNDA.n3201 GNDA.n592 0.0217373
R23060 GNDA.n3203 GNDA.n3202 0.0217373
R23061 GNDA.n3374 GNDA.n3207 0.0217373
R23062 GNDA.n3375 GNDA.n3373 0.0217373
R23063 GNDA.n3379 GNDA.n3378 0.0217373
R23064 GNDA.n5013 GNDA.n5012 0.0217373
R23065 GNDA.n5017 GNDA.n5016 0.0217373
R23066 GNDA.n5014 GNDA.n402 0.0217373
R23067 GNDA.n571 GNDA.n404 0.0217373
R23068 GNDA.n572 GNDA.n570 0.0217373
R23069 GNDA.n5009 GNDA.n5008 0.0217373
R23070 GNDA.n580 GNDA.n578 0.0217373
R23071 GNDA.n581 GNDA.n579 0.0217373
R23072 GNDA.n4997 GNDA.n4996 0.0217373
R23073 GNDA.n585 GNDA.n583 0.0217373
R23074 GNDA.n586 GNDA.n584 0.0217373
R23075 GNDA.n4993 GNDA.n4992 0.0217373
R23076 GNDA.n3682 GNDA.n3508 0.0217373
R23077 GNDA.n3437 GNDA.n3435 0.0217373
R23078 GNDA.n3438 GNDA.n3436 0.0217373
R23079 GNDA.n4985 GNDA.n4984 0.0217373
R23080 GNDA.n3442 GNDA.n3440 0.0217373
R23081 GNDA.n3443 GNDA.n3441 0.0217373
R23082 GNDA.n4981 GNDA.n4980 0.0217373
R23083 GNDA.n3447 GNDA.n3445 0.0217373
R23084 GNDA.n3448 GNDA.n3446 0.0217373
R23085 GNDA.n4977 GNDA.n4976 0.0217373
R23086 GNDA.n3452 GNDA.n3450 0.0217373
R23087 GNDA.n3453 GNDA.n3451 0.0217373
R23088 GNDA.n4973 GNDA.n4972 0.0217373
R23089 GNDA.n4964 GNDA.n3455 0.0217373
R23090 GNDA.n4965 GNDA.n4963 0.0217373
R23091 GNDA.n4969 GNDA.n4968 0.0217373
R23092 GNDA.n1694 GNDA.n781 0.0217373
R23093 GNDA.n1694 GNDA.n782 0.0217373
R23094 GNDA.n3433 GNDA.n3431 0.0217373
R23095 GNDA.n4989 GNDA.n4988 0.0217373
R23096 GNDA.n5281 GNDA.n322 0.0217373
R23097 GNDA.n5277 GNDA.n5276 0.0217373
R23098 GNDA.n5280 GNDA.n5279 0.0217373
R23099 GNDA.n6944 GNDA.n5357 0.0217373
R23100 GNDA.n6653 GNDA.n5355 0.0217373
R23101 GNDA.n5356 GNDA.n5353 0.0217373
R23102 GNDA.n5357 GNDA.n5354 0.0217373
R23103 GNDA.n6779 GNDA.n6652 0.0217373
R23104 GNDA.n6653 GNDA.n6652 0.0217373
R23105 GNDA.n7230 GNDA.n7229 0.0217373
R23106 GNDA.n7232 GNDA.n92 0.0217373
R23107 GNDA.n6657 GNDA.n6655 0.0217373
R23108 GNDA.n6658 GNDA.n6656 0.0217373
R23109 GNDA.n7230 GNDA.n90 0.0217373
R23110 GNDA.n92 GNDA.n90 0.0217373
R23111 GNDA.n7052 GNDA.n268 0.0217373
R23112 GNDA.n7059 GNDA.n7057 0.0217373
R23113 GNDA.n7055 GNDA.n262 0.0217373
R23114 GNDA.n267 GNDA.n265 0.0217373
R23115 GNDA.n7057 GNDA.n263 0.0217373
R23116 GNDA.n7056 GNDA.n7055 0.0217373
R23117 GNDA.n268 GNDA.n266 0.0217373
R23118 GNDA.n3422 GNDA.n3421 0.0217373
R23119 GNDA.n3423 GNDA.n3420 0.0217373
R23120 GNDA.n3421 GNDA.n3419 0.0217373
R23121 GNDA.n1807 GNDA.n1696 0.0217373
R23122 GNDA.n3429 GNDA.n3428 0.0217373
R23123 GNDA.n3428 GNDA.n3406 0.0217373
R23124 GNDA.n1716 GNDA.n1714 0.0217373
R23125 GNDA.n1713 GNDA.n1711 0.0217373
R23126 GNDA.n1765 GNDA.n1712 0.0217373
R23127 GNDA.n1760 GNDA.n1715 0.0217373
R23128 GNDA.n1766 GNDA.n1765 0.0217373
R23129 GNDA.n1761 GNDA.n1760 0.0217373
R23130 GNDA.n1757 GNDA.n1714 0.0217373
R23131 GNDA.n1778 GNDA.n1705 0.0217373
R23132 GNDA.n1771 GNDA.n1709 0.0217373
R23133 GNDA.n1767 GNDA.n1709 0.0217373
R23134 GNDA.n1779 GNDA.n1777 0.0217373
R23135 GNDA.n1801 GNDA.n1698 0.0217373
R23136 GNDA.n1786 GNDA.n1700 0.0217373
R23137 GNDA.n1703 GNDA.n1700 0.0217373
R23138 GNDA.n1802 GNDA.n1800 0.0217373
R23139 GNDA.n1808 GNDA.n1806 0.0217373
R23140 GNDA.n1806 GNDA.n1805 0.0217373
R23141 GNDA.n1225 GNDA.n1224 0.0217373
R23142 GNDA.n1230 GNDA.n1229 0.0217373
R23143 GNDA.n1237 GNDA.n1236 0.0217373
R23144 GNDA.n1813 GNDA.n1812 0.0217373
R23145 GNDA.n1224 GNDA.n1220 0.0217373
R23146 GNDA.n1229 GNDA.n1217 0.0217373
R23147 GNDA.n1236 GNDA.n1234 0.0217373
R23148 GNDA.n1812 GNDA.n780 0.0217373
R23149 GNDA.n6947 GNDA.n5354 0.0217373
R23150 GNDA.n6945 GNDA.n5356 0.0217373
R23151 GNDA.n6946 GNDA.n6945 0.0217373
R23152 GNDA.n6948 GNDA.n6947 0.0217373
R23153 GNDA.n6781 GNDA.n6780 0.0217373
R23154 GNDA.n6661 GNDA.n6656 0.0217373
R23155 GNDA.n6780 GNDA.n6654 0.0217373
R23156 GNDA.n6659 GNDA.n6657 0.0217373
R23157 GNDA.n6660 GNDA.n6659 0.0217373
R23158 GNDA.n6662 GNDA.n6661 0.0217373
R23159 GNDA.n7233 GNDA.n91 0.0217373
R23160 GNDA.n94 GNDA.n91 0.0217373
R23161 GNDA.n266 GNDA.n264 0.0217373
R23162 GNDA.n263 GNDA.n261 0.0217373
R23163 GNDA.n7060 GNDA.n262 0.0217373
R23164 GNDA.n7053 GNDA.n265 0.0217373
R23165 GNDA.n7061 GNDA.n7060 0.0217373
R23166 GNDA.n7054 GNDA.n7053 0.0217373
R23167 GNDA.n3683 GNDA.n3510 0.0181756
R23168 GNDA.n3684 GNDA.n3683 0.0181756
R23169 GNDA.n2110 GNDA.n719 0.0181756
R23170 GNDA.n2110 GNDA.n717 0.0181756
R23171 GNDA.n2279 GNDA.n719 0.0181756
R23172 GNDA.n2276 GNDA.n717 0.0181756
R23173 GNDA.n3681 GNDA.n3510 0.0181756
R23174 GNDA.n3685 GNDA.n3684 0.0181756
R23175 GNDA.n1514 GNDA.n1354 0.00564062
R23176 GNDA.n1514 GNDA.n728 0.00564062
R23177 GNDA.n1938 GNDA.n728 0.00564062
R23178 GNDA.n2098 GNDA.n1938 0.00564062
R23179 GNDA.n2098 GNDA.n665 0.00564062
R23180 GNDA.n2401 GNDA.n665 0.00564062
R23181 GNDA.n2561 GNDA.n2401 0.00564062
R23182 GNDA.n2561 GNDA.n599 0.00564062
R23183 GNDA.n2863 GNDA.n599 0.00564062
R23184 GNDA.n3037 GNDA.n2863 0.00564062
R23185 GNDA.n3197 GNDA.n3037 0.00564062
R23186 GNDA.n3197 GNDA.n329 0.00564062
R23187 GNDA.n5272 GNDA.n329 0.00564062
R23188 GNDA.n5272 GNDA.n5135 0.00564062
R23189 GNDA.n5135 GNDA.n377 0.00564062
R23190 GNDA.n3459 GNDA.n377 0.00564062
R23191 GNDA.n3803 GNDA.n3459 0.00564062
R23192 GNDA.n3969 GNDA.n3803 0.00564062
R23193 GNDA.n4135 GNDA.n3969 0.00564062
R23194 GNDA.n4301 GNDA.n4135 0.00564062
R23195 GNDA.n4467 GNDA.n4301 0.00564062
R23196 GNDA.n4633 GNDA.n4467 0.00564062
R23197 GNDA.n4799 GNDA.n4633 0.00564062
R23198 GNDA.n4959 GNDA.n4799 0.00564062
R23199 GNDA.n1164 GNDA.n1130 0.00189531
R23200 GNDA.n1162 GNDA.n1130 0.00189531
R23201 GNDA.n1037 GNDA.n975 0.00189531
R23202 GNDA.n975 GNDA.n945 0.00189531
R23203 GNDA.n1111 GNDA.n1077 0.00188102
R23204 GNDA.n1103 GNDA.n1081 0.00188102
R23205 GNDA.n1095 GNDA.n1085 0.00188102
R23206 GNDA.n963 GNDA.n919 0.00188102
R23207 GNDA.n967 GNDA.n923 0.00188102
R23208 GNDA.n971 GNDA.n927 0.00188102
R23209 GNDA.n994 GNDA.n959 0.00188102
R23210 GNDA.n1000 GNDA.n957 0.00188102
R23211 GNDA.n1006 GNDA.n955 0.00188102
R23212 GNDA.n1012 GNDA.n953 0.00188102
R23213 GNDA.n1018 GNDA.n951 0.00188102
R23214 GNDA.n1024 GNDA.n949 0.00188102
R23215 GNDA.n1030 GNDA.n947 0.00188102
R23216 GNDA.n897 GNDA.n853 0.00188102
R23217 GNDA.n895 GNDA.n851 0.00188102
R23218 GNDA.n893 GNDA.n849 0.00188102
R23219 GNDA.n891 GNDA.n847 0.00188102
R23220 GNDA.n889 GNDA.n845 0.00188102
R23221 GNDA.n887 GNDA.n843 0.00188102
R23222 GNDA.n885 GNDA.n841 0.00188102
R23223 GNDA.n1145 GNDA.n808 0.00188102
R23224 GNDA.n1143 GNDA.n806 0.00188102
R23225 GNDA.n1141 GNDA.n804 0.00188102
R23226 GNDA.n1139 GNDA.n802 0.00188102
R23227 GNDA.n1137 GNDA.n800 0.00188102
R23228 GNDA.n1135 GNDA.n798 0.00188102
R23229 GNDA.n1133 GNDA.n796 0.00188102
R23230 GNDA.n971 GNDA.n934 0.00188102
R23231 GNDA.n967 GNDA.n938 0.00188102
R23232 GNDA.n963 GNDA.n942 0.00188102
R23233 GNDA.n995 GNDA.n994 0.00188102
R23234 GNDA.n1001 GNDA.n1000 0.00188102
R23235 GNDA.n1007 GNDA.n1006 0.00188102
R23236 GNDA.n1013 GNDA.n1012 0.00188102
R23237 GNDA.n1019 GNDA.n1018 0.00188102
R23238 GNDA.n1025 GNDA.n1024 0.00188102
R23239 GNDA.n1031 GNDA.n1030 0.00188102
R23240 GNDA.n1096 GNDA.n1095 0.00188102
R23241 GNDA.n1104 GNDA.n1103 0.00188102
R23242 GNDA.n1112 GNDA.n1111 0.00188102
R23243 GNDA.n1145 GNDA.n1060 0.00188102
R23244 GNDA.n1143 GNDA.n1062 0.00188102
R23245 GNDA.n1141 GNDA.n1064 0.00188102
R23246 GNDA.n1139 GNDA.n1066 0.00188102
R23247 GNDA.n1137 GNDA.n1068 0.00188102
R23248 GNDA.n1135 GNDA.n1070 0.00188102
R23249 GNDA.n1133 GNDA.n1072 0.00188102
R23250 GNDA.n858 GNDA.n812 0.00188102
R23251 GNDA.n862 GNDA.n816 0.00188102
R23252 GNDA.n866 GNDA.n820 0.00188102
R23253 GNDA.n866 GNDA.n828 0.00188102
R23254 GNDA.n862 GNDA.n832 0.00188102
R23255 GNDA.n858 GNDA.n836 0.00188102
R23256 GNDA.n897 GNDA.n871 0.00188102
R23257 GNDA.n895 GNDA.n873 0.00188102
R23258 GNDA.n893 GNDA.n875 0.00188102
R23259 GNDA.n891 GNDA.n877 0.00188102
R23260 GNDA.n889 GNDA.n879 0.00188102
R23261 GNDA.n887 GNDA.n881 0.00188102
R23262 GNDA.n885 GNDA.n883 0.00188102
R23263 GNDA.n1147 GNDA.n1075 0.00173422
R23264 GNDA.n1147 GNDA.n1146 0.00173422
R23265 GNDA.n1149 GNDA.n1076 0.00173422
R23266 GNDA.n1152 GNDA.n1079 0.00173422
R23267 GNDA.n1107 GNDA.n1079 0.00173422
R23268 GNDA.n1153 GNDA.n1080 0.00173422
R23269 GNDA.n1156 GNDA.n1083 0.00173422
R23270 GNDA.n1099 GNDA.n1083 0.00173422
R23271 GNDA.n1157 GNDA.n1084 0.00173422
R23272 GNDA.n1160 GNDA.n1087 0.00173422
R23273 GNDA.n1091 GNDA.n1087 0.00173422
R23274 GNDA.n1161 GNDA.n1088 0.00173422
R23275 GNDA.n977 GNDA.n917 0.00173422
R23276 GNDA.n961 GNDA.n917 0.00173422
R23277 GNDA.n978 GNDA.n918 0.00173422
R23278 GNDA.n981 GNDA.n921 0.00173422
R23279 GNDA.n965 GNDA.n921 0.00173422
R23280 GNDA.n982 GNDA.n922 0.00173422
R23281 GNDA.n985 GNDA.n925 0.00173422
R23282 GNDA.n969 GNDA.n925 0.00173422
R23283 GNDA.n986 GNDA.n926 0.00173422
R23284 GNDA.n989 GNDA.n929 0.00173422
R23285 GNDA.n973 GNDA.n929 0.00173422
R23286 GNDA.n990 GNDA.n930 0.00173422
R23287 GNDA.n991 GNDA.n960 0.00173422
R23288 GNDA.n997 GNDA.n958 0.00173422
R23289 GNDA.n1003 GNDA.n956 0.00173422
R23290 GNDA.n1009 GNDA.n954 0.00173422
R23291 GNDA.n1015 GNDA.n952 0.00173422
R23292 GNDA.n1021 GNDA.n950 0.00173422
R23293 GNDA.n1027 GNDA.n948 0.00173422
R23294 GNDA.n1033 GNDA.n946 0.00173422
R23295 GNDA.n898 GNDA.n855 0.00173422
R23296 GNDA.n896 GNDA.n852 0.00173422
R23297 GNDA.n894 GNDA.n850 0.00173422
R23298 GNDA.n892 GNDA.n848 0.00173422
R23299 GNDA.n890 GNDA.n846 0.00173422
R23300 GNDA.n888 GNDA.n844 0.00173422
R23301 GNDA.n886 GNDA.n842 0.00173422
R23302 GNDA.n900 GNDA.n840 0.00173422
R23303 GNDA.n1148 GNDA.n809 0.00173422
R23304 GNDA.n1144 GNDA.n807 0.00173422
R23305 GNDA.n1142 GNDA.n805 0.00173422
R23306 GNDA.n1140 GNDA.n803 0.00173422
R23307 GNDA.n1138 GNDA.n801 0.00173422
R23308 GNDA.n1136 GNDA.n799 0.00173422
R23309 GNDA.n1134 GNDA.n797 0.00173422
R23310 GNDA.n1132 GNDA.n795 0.00173422
R23311 GNDA.n973 GNDA.n932 0.00173422
R23312 GNDA.n969 GNDA.n936 0.00173422
R23313 GNDA.n965 GNDA.n940 0.00173422
R23314 GNDA.n961 GNDA.n944 0.00173422
R23315 GNDA.n992 GNDA.n991 0.00173422
R23316 GNDA.n990 GNDA.n932 0.00173422
R23317 GNDA.n989 GNDA.n933 0.00173422
R23318 GNDA.n986 GNDA.n936 0.00173422
R23319 GNDA.n985 GNDA.n937 0.00173422
R23320 GNDA.n982 GNDA.n940 0.00173422
R23321 GNDA.n981 GNDA.n941 0.00173422
R23322 GNDA.n978 GNDA.n944 0.00173422
R23323 GNDA.n977 GNDA.n945 0.00173422
R23324 GNDA.n998 GNDA.n997 0.00173422
R23325 GNDA.n1004 GNDA.n1003 0.00173422
R23326 GNDA.n1010 GNDA.n1009 0.00173422
R23327 GNDA.n1016 GNDA.n1015 0.00173422
R23328 GNDA.n1022 GNDA.n1021 0.00173422
R23329 GNDA.n1028 GNDA.n1027 0.00173422
R23330 GNDA.n1036 GNDA.n1033 0.00173422
R23331 GNDA.n1092 GNDA.n1091 0.00173422
R23332 GNDA.n1100 GNDA.n1099 0.00173422
R23333 GNDA.n1108 GNDA.n1107 0.00173422
R23334 GNDA.n1146 GNDA.n1115 0.00173422
R23335 GNDA.n1161 GNDA.n1092 0.00173422
R23336 GNDA.n1160 GNDA.n1094 0.00173422
R23337 GNDA.n1157 GNDA.n1100 0.00173422
R23338 GNDA.n1156 GNDA.n1102 0.00173422
R23339 GNDA.n1153 GNDA.n1108 0.00173422
R23340 GNDA.n1152 GNDA.n1110 0.00173422
R23341 GNDA.n1149 GNDA.n1115 0.00173422
R23342 GNDA.n1163 GNDA.n1148 0.00173422
R23343 GNDA.n1144 GNDA.n1061 0.00173422
R23344 GNDA.n1142 GNDA.n1063 0.00173422
R23345 GNDA.n1140 GNDA.n1065 0.00173422
R23346 GNDA.n1138 GNDA.n1067 0.00173422
R23347 GNDA.n1136 GNDA.n1069 0.00173422
R23348 GNDA.n1134 GNDA.n1071 0.00173422
R23349 GNDA.n1132 GNDA.n1073 0.00173422
R23350 GNDA.n1162 GNDA.n1075 0.00173422
R23351 GNDA.n1055 GNDA.n1054 0.00173422
R23352 GNDA.n915 GNDA.n901 0.00173422
R23353 GNDA.n1039 GNDA.n838 0.00173422
R23354 GNDA.n1042 GNDA.n835 0.00173422
R23355 GNDA.n860 GNDA.n814 0.00173422
R23356 GNDA.n1043 GNDA.n834 0.00173422
R23357 GNDA.n1046 GNDA.n831 0.00173422
R23358 GNDA.n864 GNDA.n818 0.00173422
R23359 GNDA.n1047 GNDA.n830 0.00173422
R23360 GNDA.n1050 GNDA.n827 0.00173422
R23361 GNDA.n868 GNDA.n822 0.00173422
R23362 GNDA.n1051 GNDA.n826 0.00173422
R23363 GNDA.n1051 GNDA.n823 0.00173422
R23364 GNDA.n1050 GNDA.n822 0.00173422
R23365 GNDA.n1047 GNDA.n819 0.00173422
R23366 GNDA.n1046 GNDA.n818 0.00173422
R23367 GNDA.n1043 GNDA.n815 0.00173422
R23368 GNDA.n1042 GNDA.n814 0.00173422
R23369 GNDA.n1039 GNDA.n811 0.00173422
R23370 GNDA.n1054 GNDA.n915 0.00173422
R23371 GNDA.n868 GNDA.n826 0.00173422
R23372 GNDA.n864 GNDA.n830 0.00173422
R23373 GNDA.n860 GNDA.n834 0.00173422
R23374 GNDA.n901 GNDA.n838 0.00173422
R23375 GNDA.n898 GNDA.n869 0.00173422
R23376 GNDA.n896 GNDA.n872 0.00173422
R23377 GNDA.n894 GNDA.n874 0.00173422
R23378 GNDA.n892 GNDA.n876 0.00173422
R23379 GNDA.n890 GNDA.n878 0.00173422
R23380 GNDA.n888 GNDA.n880 0.00173422
R23381 GNDA.n886 GNDA.n882 0.00173422
R23382 GNDA.n1056 GNDA.n900 0.00173422
R23383 GNDA.n1113 GNDA.n1076 0.00169751
R23384 GNDA.n1150 GNDA.n1077 0.00169751
R23385 GNDA.n1151 GNDA.n1078 0.00169751
R23386 GNDA.n1109 GNDA.n1078 0.00169751
R23387 GNDA.n1105 GNDA.n1080 0.00169751
R23388 GNDA.n1154 GNDA.n1081 0.00169751
R23389 GNDA.n1155 GNDA.n1082 0.00169751
R23390 GNDA.n1101 GNDA.n1082 0.00169751
R23391 GNDA.n1097 GNDA.n1084 0.00169751
R23392 GNDA.n1158 GNDA.n1085 0.00169751
R23393 GNDA.n1159 GNDA.n1086 0.00169751
R23394 GNDA.n1093 GNDA.n1086 0.00169751
R23395 GNDA.n1089 GNDA.n1088 0.00169751
R23396 GNDA.n1166 GNDA.n794 0.00169751
R23397 GNDA.n962 GNDA.n918 0.00169751
R23398 GNDA.n979 GNDA.n919 0.00169751
R23399 GNDA.n980 GNDA.n920 0.00169751
R23400 GNDA.n964 GNDA.n920 0.00169751
R23401 GNDA.n966 GNDA.n922 0.00169751
R23402 GNDA.n983 GNDA.n923 0.00169751
R23403 GNDA.n984 GNDA.n924 0.00169751
R23404 GNDA.n968 GNDA.n924 0.00169751
R23405 GNDA.n970 GNDA.n926 0.00169751
R23406 GNDA.n987 GNDA.n927 0.00169751
R23407 GNDA.n988 GNDA.n928 0.00169751
R23408 GNDA.n972 GNDA.n928 0.00169751
R23409 GNDA.n1034 GNDA.n930 0.00169751
R23410 GNDA.n931 GNDA.n98 0.00169751
R23411 GNDA.n1035 GNDA.n1034 0.00169751
R23412 GNDA.n972 GNDA.n933 0.00169751
R23413 GNDA.n970 GNDA.n935 0.00169751
R23414 GNDA.n968 GNDA.n937 0.00169751
R23415 GNDA.n966 GNDA.n939 0.00169751
R23416 GNDA.n964 GNDA.n941 0.00169751
R23417 GNDA.n962 GNDA.n943 0.00169751
R23418 GNDA.n988 GNDA.n934 0.00169751
R23419 GNDA.n987 GNDA.n935 0.00169751
R23420 GNDA.n984 GNDA.n938 0.00169751
R23421 GNDA.n983 GNDA.n939 0.00169751
R23422 GNDA.n980 GNDA.n942 0.00169751
R23423 GNDA.n979 GNDA.n943 0.00169751
R23424 GNDA.n1035 GNDA.n931 0.00169751
R23425 GNDA.n1090 GNDA.n1089 0.00169751
R23426 GNDA.n1094 GNDA.n1093 0.00169751
R23427 GNDA.n1098 GNDA.n1097 0.00169751
R23428 GNDA.n1102 GNDA.n1101 0.00169751
R23429 GNDA.n1106 GNDA.n1105 0.00169751
R23430 GNDA.n1110 GNDA.n1109 0.00169751
R23431 GNDA.n1114 GNDA.n1113 0.00169751
R23432 GNDA.n1090 GNDA.n794 0.00169751
R23433 GNDA.n1159 GNDA.n1096 0.00169751
R23434 GNDA.n1158 GNDA.n1098 0.00169751
R23435 GNDA.n1155 GNDA.n1104 0.00169751
R23436 GNDA.n1154 GNDA.n1106 0.00169751
R23437 GNDA.n1151 GNDA.n1112 0.00169751
R23438 GNDA.n1150 GNDA.n1114 0.00169751
R23439 GNDA.n1057 GNDA.n856 0.00169751
R23440 GNDA.n1055 GNDA.n839 0.00169751
R23441 GNDA.n857 GNDA.n811 0.00169751
R23442 GNDA.n1040 GNDA.n837 0.00169751
R23443 GNDA.n1041 GNDA.n836 0.00169751
R23444 GNDA.n859 GNDA.n813 0.00169751
R23445 GNDA.n861 GNDA.n815 0.00169751
R23446 GNDA.n1044 GNDA.n833 0.00169751
R23447 GNDA.n1045 GNDA.n832 0.00169751
R23448 GNDA.n863 GNDA.n817 0.00169751
R23449 GNDA.n865 GNDA.n819 0.00169751
R23450 GNDA.n1048 GNDA.n829 0.00169751
R23451 GNDA.n1049 GNDA.n828 0.00169751
R23452 GNDA.n867 GNDA.n821 0.00169751
R23453 GNDA.n854 GNDA.n823 0.00169751
R23454 GNDA.n870 GNDA.n824 0.00169751
R23455 GNDA.n1049 GNDA.n821 0.00169751
R23456 GNDA.n1048 GNDA.n820 0.00169751
R23457 GNDA.n1045 GNDA.n817 0.00169751
R23458 GNDA.n1044 GNDA.n816 0.00169751
R23459 GNDA.n1041 GNDA.n813 0.00169751
R23460 GNDA.n1040 GNDA.n812 0.00169751
R23461 GNDA.n899 GNDA.n856 0.00169751
R23462 GNDA.n867 GNDA.n827 0.00169751
R23463 GNDA.n865 GNDA.n829 0.00169751
R23464 GNDA.n863 GNDA.n831 0.00169751
R23465 GNDA.n861 GNDA.n833 0.00169751
R23466 GNDA.n859 GNDA.n835 0.00169751
R23467 GNDA.n857 GNDA.n837 0.00169751
R23468 GNDA.n854 GNDA.n825 0.00169751
R23469 GNDA.n870 GNDA.n825 0.00169751
R23470 GNDA.n899 GNDA.n839 0.00169751
R23471 GNDA.n992 GNDA.n976 0.00166081
R23472 GNDA.n995 GNDA.n993 0.00166081
R23473 GNDA.n998 GNDA.n996 0.00166081
R23474 GNDA.n1001 GNDA.n999 0.00166081
R23475 GNDA.n1004 GNDA.n1002 0.00166081
R23476 GNDA.n1007 GNDA.n1005 0.00166081
R23477 GNDA.n1010 GNDA.n1008 0.00166081
R23478 GNDA.n1013 GNDA.n1011 0.00166081
R23479 GNDA.n1016 GNDA.n1014 0.00166081
R23480 GNDA.n1019 GNDA.n1017 0.00166081
R23481 GNDA.n1022 GNDA.n1020 0.00166081
R23482 GNDA.n1025 GNDA.n1023 0.00166081
R23483 GNDA.n1028 GNDA.n1026 0.00166081
R23484 GNDA.n1031 GNDA.n1029 0.00166081
R23485 GNDA.n1036 GNDA.n1032 0.00166081
R23486 GNDA.n1038 GNDA.n916 0.00166081
R23487 GNDA.n1052 GNDA.n869 0.00166081
R23488 GNDA.n902 GNDA.n871 0.00166081
R23489 GNDA.n903 GNDA.n872 0.00166081
R23490 GNDA.n904 GNDA.n873 0.00166081
R23491 GNDA.n905 GNDA.n874 0.00166081
R23492 GNDA.n906 GNDA.n875 0.00166081
R23493 GNDA.n907 GNDA.n876 0.00166081
R23494 GNDA.n908 GNDA.n877 0.00166081
R23495 GNDA.n909 GNDA.n878 0.00166081
R23496 GNDA.n910 GNDA.n879 0.00166081
R23497 GNDA.n911 GNDA.n880 0.00166081
R23498 GNDA.n912 GNDA.n881 0.00166081
R23499 GNDA.n913 GNDA.n882 0.00166081
R23500 GNDA.n914 GNDA.n883 0.00166081
R23501 GNDA.n1056 GNDA.n884 0.00166081
R23502 GNDA.n1058 GNDA.n810 0.00166081
R23503 GNDA.n1163 GNDA.n1131 0.00166081
R23504 GNDA.n1116 GNDA.n1060 0.00166081
R23505 GNDA.n1117 GNDA.n1061 0.00166081
R23506 GNDA.n1118 GNDA.n1062 0.00166081
R23507 GNDA.n1119 GNDA.n1063 0.00166081
R23508 GNDA.n1120 GNDA.n1064 0.00166081
R23509 GNDA.n1121 GNDA.n1065 0.00166081
R23510 GNDA.n1122 GNDA.n1066 0.00166081
R23511 GNDA.n1123 GNDA.n1067 0.00166081
R23512 GNDA.n1124 GNDA.n1068 0.00166081
R23513 GNDA.n1125 GNDA.n1069 0.00166081
R23514 GNDA.n1126 GNDA.n1070 0.00166081
R23515 GNDA.n1127 GNDA.n1071 0.00166081
R23516 GNDA.n1128 GNDA.n1072 0.00166081
R23517 GNDA.n1129 GNDA.n1073 0.00166081
R23518 GNDA.n1165 GNDA.n1074 0.00166081
R23519 GNDA.n976 GNDA.n974 0.00166081
R23520 GNDA.n993 GNDA.n960 0.00166081
R23521 GNDA.n996 GNDA.n959 0.00166081
R23522 GNDA.n999 GNDA.n958 0.00166081
R23523 GNDA.n1002 GNDA.n957 0.00166081
R23524 GNDA.n1005 GNDA.n956 0.00166081
R23525 GNDA.n1008 GNDA.n955 0.00166081
R23526 GNDA.n1011 GNDA.n954 0.00166081
R23527 GNDA.n1014 GNDA.n953 0.00166081
R23528 GNDA.n1017 GNDA.n952 0.00166081
R23529 GNDA.n1020 GNDA.n951 0.00166081
R23530 GNDA.n1023 GNDA.n950 0.00166081
R23531 GNDA.n1026 GNDA.n949 0.00166081
R23532 GNDA.n1029 GNDA.n948 0.00166081
R23533 GNDA.n1032 GNDA.n947 0.00166081
R23534 GNDA.n946 GNDA.n916 0.00166081
R23535 GNDA.n1131 GNDA.n1059 0.00166081
R23536 GNDA.n1116 GNDA.n809 0.00166081
R23537 GNDA.n1117 GNDA.n808 0.00166081
R23538 GNDA.n1118 GNDA.n807 0.00166081
R23539 GNDA.n1119 GNDA.n806 0.00166081
R23540 GNDA.n1120 GNDA.n805 0.00166081
R23541 GNDA.n1121 GNDA.n804 0.00166081
R23542 GNDA.n1122 GNDA.n803 0.00166081
R23543 GNDA.n1123 GNDA.n802 0.00166081
R23544 GNDA.n1124 GNDA.n801 0.00166081
R23545 GNDA.n1125 GNDA.n800 0.00166081
R23546 GNDA.n1126 GNDA.n799 0.00166081
R23547 GNDA.n1127 GNDA.n798 0.00166081
R23548 GNDA.n1128 GNDA.n797 0.00166081
R23549 GNDA.n1129 GNDA.n796 0.00166081
R23550 GNDA.n1074 GNDA.n795 0.00166081
R23551 GNDA.n1053 GNDA.n1052 0.00166081
R23552 GNDA.n902 GNDA.n855 0.00166081
R23553 GNDA.n903 GNDA.n853 0.00166081
R23554 GNDA.n904 GNDA.n852 0.00166081
R23555 GNDA.n905 GNDA.n851 0.00166081
R23556 GNDA.n906 GNDA.n850 0.00166081
R23557 GNDA.n907 GNDA.n849 0.00166081
R23558 GNDA.n908 GNDA.n848 0.00166081
R23559 GNDA.n909 GNDA.n847 0.00166081
R23560 GNDA.n910 GNDA.n846 0.00166081
R23561 GNDA.n911 GNDA.n845 0.00166081
R23562 GNDA.n912 GNDA.n844 0.00166081
R23563 GNDA.n913 GNDA.n843 0.00166081
R23564 GNDA.n914 GNDA.n842 0.00166081
R23565 GNDA.n884 GNDA.n841 0.00166081
R23566 GNDA.n840 GNDA.n810 0.00166081
R23567 VIN+.n0 VIN+.t8 1097.62
R23568 VIN+ VIN+.n9 433.019
R23569 VIN+.n9 VIN+.t4 273.134
R23570 VIN+.n0 VIN+.t6 273.134
R23571 VIN+.n8 VIN+.t0 273.134
R23572 VIN+.n7 VIN+.t3 273.134
R23573 VIN+.n6 VIN+.t10 273.134
R23574 VIN+.n5 VIN+.t2 273.134
R23575 VIN+.n4 VIN+.t7 273.134
R23576 VIN+.n3 VIN+.t5 273.134
R23577 VIN+.n2 VIN+.t9 273.134
R23578 VIN+.n1 VIN+.t1 273.134
R23579 VIN+.n1 VIN+.n0 176.733
R23580 VIN+.n2 VIN+.n1 176.733
R23581 VIN+.n3 VIN+.n2 176.733
R23582 VIN+.n4 VIN+.n3 176.733
R23583 VIN+.n5 VIN+.n4 176.733
R23584 VIN+.n6 VIN+.n5 176.733
R23585 VIN+.n7 VIN+.n6 176.733
R23586 VIN+.n8 VIN+.n7 176.733
R23587 VIN+.n9 VIN+.n8 176.733
R23588 two_stage_opamp_dummy_magic_25_0.V_source.n17 two_stage_opamp_dummy_magic_25_0.V_source.t11 82.6422
R23589 two_stage_opamp_dummy_magic_25_0.V_source.n32 two_stage_opamp_dummy_magic_25_0.V_source.n31 49.3505
R23590 two_stage_opamp_dummy_magic_25_0.V_source.n30 two_stage_opamp_dummy_magic_25_0.V_source.n29 49.3505
R23591 two_stage_opamp_dummy_magic_25_0.V_source.n22 two_stage_opamp_dummy_magic_25_0.V_source.n21 49.3505
R23592 two_stage_opamp_dummy_magic_25_0.V_source.n38 two_stage_opamp_dummy_magic_25_0.V_source.n37 49.3505
R23593 two_stage_opamp_dummy_magic_25_0.V_source.n35 two_stage_opamp_dummy_magic_25_0.V_source.n34 49.3505
R23594 two_stage_opamp_dummy_magic_25_0.V_source.n47 two_stage_opamp_dummy_magic_25_0.V_source.n46 49.3505
R23595 two_stage_opamp_dummy_magic_25_0.V_source.n43 two_stage_opamp_dummy_magic_25_0.V_source.n42 49.3505
R23596 two_stage_opamp_dummy_magic_25_0.V_source.n41 two_stage_opamp_dummy_magic_25_0.V_source.n40 49.3505
R23597 two_stage_opamp_dummy_magic_25_0.V_source.n26 two_stage_opamp_dummy_magic_25_0.V_source.n25 49.3505
R23598 two_stage_opamp_dummy_magic_25_0.V_source.n24 two_stage_opamp_dummy_magic_25_0.V_source.n23 49.3505
R23599 two_stage_opamp_dummy_magic_25_0.V_source.n9 two_stage_opamp_dummy_magic_25_0.V_source.n49 32.3838
R23600 two_stage_opamp_dummy_magic_25_0.V_source.n51 two_stage_opamp_dummy_magic_25_0.V_source.n50 32.3838
R23601 two_stage_opamp_dummy_magic_25_0.V_source.n4 two_stage_opamp_dummy_magic_25_0.V_source.n12 32.3838
R23602 two_stage_opamp_dummy_magic_25_0.V_source.n16 two_stage_opamp_dummy_magic_25_0.V_source.n15 32.3838
R23603 two_stage_opamp_dummy_magic_25_0.V_source.n14 two_stage_opamp_dummy_magic_25_0.V_source.n13 32.3838
R23604 two_stage_opamp_dummy_magic_25_0.V_source.n19 two_stage_opamp_dummy_magic_25_0.V_source.n18 32.3838
R23605 two_stage_opamp_dummy_magic_25_0.V_source.n55 two_stage_opamp_dummy_magic_25_0.V_source.n54 32.3838
R23606 two_stage_opamp_dummy_magic_25_0.V_source.n57 two_stage_opamp_dummy_magic_25_0.V_source.n56 32.3838
R23607 two_stage_opamp_dummy_magic_25_0.V_source.n59 two_stage_opamp_dummy_magic_25_0.V_source.n58 32.3838
R23608 two_stage_opamp_dummy_magic_25_0.V_source.n53 two_stage_opamp_dummy_magic_25_0.V_source.n52 32.3838
R23609 two_stage_opamp_dummy_magic_25_0.V_source.n31 two_stage_opamp_dummy_magic_25_0.V_source.t9 16.0005
R23610 two_stage_opamp_dummy_magic_25_0.V_source.n31 two_stage_opamp_dummy_magic_25_0.V_source.t32 16.0005
R23611 two_stage_opamp_dummy_magic_25_0.V_source.n29 two_stage_opamp_dummy_magic_25_0.V_source.t2 16.0005
R23612 two_stage_opamp_dummy_magic_25_0.V_source.n29 two_stage_opamp_dummy_magic_25_0.V_source.t38 16.0005
R23613 two_stage_opamp_dummy_magic_25_0.V_source.n21 two_stage_opamp_dummy_magic_25_0.V_source.t29 16.0005
R23614 two_stage_opamp_dummy_magic_25_0.V_source.n21 two_stage_opamp_dummy_magic_25_0.V_source.t1 16.0005
R23615 two_stage_opamp_dummy_magic_25_0.V_source.n37 two_stage_opamp_dummy_magic_25_0.V_source.t16 16.0005
R23616 two_stage_opamp_dummy_magic_25_0.V_source.n37 two_stage_opamp_dummy_magic_25_0.V_source.t18 16.0005
R23617 two_stage_opamp_dummy_magic_25_0.V_source.n34 two_stage_opamp_dummy_magic_25_0.V_source.t17 16.0005
R23618 two_stage_opamp_dummy_magic_25_0.V_source.n34 two_stage_opamp_dummy_magic_25_0.V_source.t12 16.0005
R23619 two_stage_opamp_dummy_magic_25_0.V_source.n46 two_stage_opamp_dummy_magic_25_0.V_source.t20 16.0005
R23620 two_stage_opamp_dummy_magic_25_0.V_source.n46 two_stage_opamp_dummy_magic_25_0.V_source.t19 16.0005
R23621 two_stage_opamp_dummy_magic_25_0.V_source.n42 two_stage_opamp_dummy_magic_25_0.V_source.t15 16.0005
R23622 two_stage_opamp_dummy_magic_25_0.V_source.n42 two_stage_opamp_dummy_magic_25_0.V_source.t21 16.0005
R23623 two_stage_opamp_dummy_magic_25_0.V_source.n40 two_stage_opamp_dummy_magic_25_0.V_source.t13 16.0005
R23624 two_stage_opamp_dummy_magic_25_0.V_source.n40 two_stage_opamp_dummy_magic_25_0.V_source.t14 16.0005
R23625 two_stage_opamp_dummy_magic_25_0.V_source.n25 two_stage_opamp_dummy_magic_25_0.V_source.t27 16.0005
R23626 two_stage_opamp_dummy_magic_25_0.V_source.n25 two_stage_opamp_dummy_magic_25_0.V_source.t28 16.0005
R23627 two_stage_opamp_dummy_magic_25_0.V_source.n23 two_stage_opamp_dummy_magic_25_0.V_source.t26 16.0005
R23628 two_stage_opamp_dummy_magic_25_0.V_source.n23 two_stage_opamp_dummy_magic_25_0.V_source.t0 16.0005
R23629 two_stage_opamp_dummy_magic_25_0.V_source.n49 two_stage_opamp_dummy_magic_25_0.V_source.t33 9.6005
R23630 two_stage_opamp_dummy_magic_25_0.V_source.n49 two_stage_opamp_dummy_magic_25_0.V_source.t40 9.6005
R23631 two_stage_opamp_dummy_magic_25_0.V_source.n50 two_stage_opamp_dummy_magic_25_0.V_source.t22 9.6005
R23632 two_stage_opamp_dummy_magic_25_0.V_source.n50 two_stage_opamp_dummy_magic_25_0.V_source.t39 9.6005
R23633 two_stage_opamp_dummy_magic_25_0.V_source.n12 two_stage_opamp_dummy_magic_25_0.V_source.t24 9.6005
R23634 two_stage_opamp_dummy_magic_25_0.V_source.n12 two_stage_opamp_dummy_magic_25_0.V_source.t5 9.6005
R23635 two_stage_opamp_dummy_magic_25_0.V_source.n15 two_stage_opamp_dummy_magic_25_0.V_source.t31 9.6005
R23636 two_stage_opamp_dummy_magic_25_0.V_source.n15 two_stage_opamp_dummy_magic_25_0.V_source.t37 9.6005
R23637 two_stage_opamp_dummy_magic_25_0.V_source.n13 two_stage_opamp_dummy_magic_25_0.V_source.t7 9.6005
R23638 two_stage_opamp_dummy_magic_25_0.V_source.n13 two_stage_opamp_dummy_magic_25_0.V_source.t35 9.6005
R23639 two_stage_opamp_dummy_magic_25_0.V_source.n18 two_stage_opamp_dummy_magic_25_0.V_source.t8 9.6005
R23640 two_stage_opamp_dummy_magic_25_0.V_source.n18 two_stage_opamp_dummy_magic_25_0.V_source.t6 9.6005
R23641 two_stage_opamp_dummy_magic_25_0.V_source.n54 two_stage_opamp_dummy_magic_25_0.V_source.t34 9.6005
R23642 two_stage_opamp_dummy_magic_25_0.V_source.n54 two_stage_opamp_dummy_magic_25_0.V_source.t36 9.6005
R23643 two_stage_opamp_dummy_magic_25_0.V_source.n56 two_stage_opamp_dummy_magic_25_0.V_source.t10 9.6005
R23644 two_stage_opamp_dummy_magic_25_0.V_source.n56 two_stage_opamp_dummy_magic_25_0.V_source.t25 9.6005
R23645 two_stage_opamp_dummy_magic_25_0.V_source.n58 two_stage_opamp_dummy_magic_25_0.V_source.t4 9.6005
R23646 two_stage_opamp_dummy_magic_25_0.V_source.n58 two_stage_opamp_dummy_magic_25_0.V_source.t30 9.6005
R23647 two_stage_opamp_dummy_magic_25_0.V_source.n52 two_stage_opamp_dummy_magic_25_0.V_source.t3 9.6005
R23648 two_stage_opamp_dummy_magic_25_0.V_source.n52 two_stage_opamp_dummy_magic_25_0.V_source.t23 9.6005
R23649 two_stage_opamp_dummy_magic_25_0.V_source.n61 two_stage_opamp_dummy_magic_25_0.V_source.n4 5.85227
R23650 two_stage_opamp_dummy_magic_25_0.V_source.n51 two_stage_opamp_dummy_magic_25_0.V_source.n8 5.71925
R23651 two_stage_opamp_dummy_magic_25_0.V_source.n5 two_stage_opamp_dummy_magic_25_0.V_source.n4 5.71925
R23652 two_stage_opamp_dummy_magic_25_0.V_source.n41 two_stage_opamp_dummy_magic_25_0.V_source.n2 5.51092
R23653 two_stage_opamp_dummy_magic_25_0.V_source.n1 two_stage_opamp_dummy_magic_25_0.V_source.n22 5.51092
R23654 two_stage_opamp_dummy_magic_25_0.V_source.n44 two_stage_opamp_dummy_magic_25_0.V_source.n41 5.45883
R23655 two_stage_opamp_dummy_magic_25_0.V_source.n22 two_stage_opamp_dummy_magic_25_0.V_source.n20 5.45883
R23656 two_stage_opamp_dummy_magic_25_0.V_source.n8 two_stage_opamp_dummy_magic_25_0.V_source.n9 5.3755
R23657 two_stage_opamp_dummy_magic_25_0.V_source.n5 two_stage_opamp_dummy_magic_25_0.V_source.n14 5.3755
R23658 two_stage_opamp_dummy_magic_25_0.V_source.n7 two_stage_opamp_dummy_magic_25_0.V_source.n19 5.3755
R23659 two_stage_opamp_dummy_magic_25_0.V_source.n6 two_stage_opamp_dummy_magic_25_0.V_source.n55 5.3755
R23660 two_stage_opamp_dummy_magic_25_0.V_source.n6 two_stage_opamp_dummy_magic_25_0.V_source.n57 5.3755
R23661 two_stage_opamp_dummy_magic_25_0.V_source.n59 two_stage_opamp_dummy_magic_25_0.V_source.n7 5.3755
R23662 two_stage_opamp_dummy_magic_25_0.V_source.n53 two_stage_opamp_dummy_magic_25_0.V_source.n8 5.3755
R23663 two_stage_opamp_dummy_magic_25_0.V_source.n55 two_stage_opamp_dummy_magic_25_0.V_source.n3 5.188
R23664 two_stage_opamp_dummy_magic_25_0.V_source.n57 two_stage_opamp_dummy_magic_25_0.V_source.n3 5.188
R23665 two_stage_opamp_dummy_magic_25_0.V_source.n60 two_stage_opamp_dummy_magic_25_0.V_source.n59 5.188
R23666 two_stage_opamp_dummy_magic_25_0.V_source.n2 two_stage_opamp_dummy_magic_25_0.V_source.n47 5.16717
R23667 two_stage_opamp_dummy_magic_25_0.V_source.n43 two_stage_opamp_dummy_magic_25_0.V_source.n2 5.16717
R23668 two_stage_opamp_dummy_magic_25_0.V_source.n26 two_stage_opamp_dummy_magic_25_0.V_source.n1 5.16717
R23669 two_stage_opamp_dummy_magic_25_0.V_source.n1 two_stage_opamp_dummy_magic_25_0.V_source.n24 5.16717
R23670 two_stage_opamp_dummy_magic_25_0.V_source.n39 two_stage_opamp_dummy_magic_25_0.V_source.n38 4.89633
R23671 two_stage_opamp_dummy_magic_25_0.V_source.n47 two_stage_opamp_dummy_magic_25_0.V_source.n45 4.89633
R23672 two_stage_opamp_dummy_magic_25_0.V_source.n44 two_stage_opamp_dummy_magic_25_0.V_source.n43 4.89633
R23673 two_stage_opamp_dummy_magic_25_0.V_source.n33 two_stage_opamp_dummy_magic_25_0.V_source.n32 4.89633
R23674 two_stage_opamp_dummy_magic_25_0.V_source.n36 two_stage_opamp_dummy_magic_25_0.V_source.n35 4.89633
R23675 two_stage_opamp_dummy_magic_25_0.V_source.n27 two_stage_opamp_dummy_magic_25_0.V_source.n26 4.89633
R23676 two_stage_opamp_dummy_magic_25_0.V_source.n24 two_stage_opamp_dummy_magic_25_0.V_source.n20 4.89633
R23677 two_stage_opamp_dummy_magic_25_0.V_source.n30 two_stage_opamp_dummy_magic_25_0.V_source.n28 4.89633
R23678 two_stage_opamp_dummy_magic_25_0.V_source.n5 two_stage_opamp_dummy_magic_25_0.V_source.n17 4.5005
R23679 two_stage_opamp_dummy_magic_25_0.V_source.n36 two_stage_opamp_dummy_magic_25_0.V_source.n33 3.6255
R23680 two_stage_opamp_dummy_magic_25_0.V_source.n48 two_stage_opamp_dummy_magic_25_0.V_source.n0 2.2076
R23681 two_stage_opamp_dummy_magic_25_0.V_source.n11 two_stage_opamp_dummy_magic_25_0.V_source.n48 2.16822
R23682 two_stage_opamp_dummy_magic_25_0.V_source.n0 two_stage_opamp_dummy_magic_25_0.V_source.n10 2.16822
R23683 two_stage_opamp_dummy_magic_25_0.V_source.n3 two_stage_opamp_dummy_magic_25_0.V_source.n11 2.02255
R23684 two_stage_opamp_dummy_magic_25_0.V_source.n10 two_stage_opamp_dummy_magic_25_0.V_source.n61 1.36007
R23685 two_stage_opamp_dummy_magic_25_0.V_source.n7 two_stage_opamp_dummy_magic_25_0.V_source.n5 1.03175
R23686 two_stage_opamp_dummy_magic_25_0.V_source.n17 two_stage_opamp_dummy_magic_25_0.V_source.n16 0.8755
R23687 two_stage_opamp_dummy_magic_25_0.V_source.n38 two_stage_opamp_dummy_magic_25_0.V_source.n11 0.871494
R23688 two_stage_opamp_dummy_magic_25_0.V_source.n32 two_stage_opamp_dummy_magic_25_0.V_source.n10 0.871494
R23689 two_stage_opamp_dummy_magic_25_0.V_source.n48 two_stage_opamp_dummy_magic_25_0.V_source.n2 0.854052
R23690 two_stage_opamp_dummy_magic_25_0.V_source.n1 two_stage_opamp_dummy_magic_25_0.V_source.n0 0.854052
R23691 two_stage_opamp_dummy_magic_25_0.V_source.n6 two_stage_opamp_dummy_magic_25_0.V_source.n8 0.688
R23692 two_stage_opamp_dummy_magic_25_0.V_source.n7 two_stage_opamp_dummy_magic_25_0.V_source.n6 0.688
R23693 two_stage_opamp_dummy_magic_25_0.V_source.n60 two_stage_opamp_dummy_magic_25_0.V_source.n3 0.688
R23694 two_stage_opamp_dummy_magic_25_0.V_source.n61 two_stage_opamp_dummy_magic_25_0.V_source.n60 0.664374
R23695 two_stage_opamp_dummy_magic_25_0.V_source.n11 two_stage_opamp_dummy_magic_25_0.V_source.n9 0.6255
R23696 two_stage_opamp_dummy_magic_25_0.V_source.n11 two_stage_opamp_dummy_magic_25_0.V_source.n51 0.6255
R23697 two_stage_opamp_dummy_magic_25_0.V_source.n19 two_stage_opamp_dummy_magic_25_0.V_source.n10 0.6255
R23698 two_stage_opamp_dummy_magic_25_0.V_source.n14 two_stage_opamp_dummy_magic_25_0.V_source.n10 0.6255
R23699 two_stage_opamp_dummy_magic_25_0.V_source.n16 two_stage_opamp_dummy_magic_25_0.V_source.n10 0.6255
R23700 two_stage_opamp_dummy_magic_25_0.V_source.n11 two_stage_opamp_dummy_magic_25_0.V_source.n53 0.6255
R23701 two_stage_opamp_dummy_magic_25_0.V_source.n35 two_stage_opamp_dummy_magic_25_0.V_source.n11 0.604667
R23702 two_stage_opamp_dummy_magic_25_0.V_source.n10 two_stage_opamp_dummy_magic_25_0.V_source.n30 0.604667
R23703 two_stage_opamp_dummy_magic_25_0.V_source.n45 two_stage_opamp_dummy_magic_25_0.V_source.n44 0.563
R23704 two_stage_opamp_dummy_magic_25_0.V_source.n45 two_stage_opamp_dummy_magic_25_0.V_source.n39 0.563
R23705 two_stage_opamp_dummy_magic_25_0.V_source.n39 two_stage_opamp_dummy_magic_25_0.V_source.n36 0.563
R23706 two_stage_opamp_dummy_magic_25_0.V_source.n33 two_stage_opamp_dummy_magic_25_0.V_source.n28 0.563
R23707 two_stage_opamp_dummy_magic_25_0.V_source.n27 two_stage_opamp_dummy_magic_25_0.V_source.n20 0.563
R23708 two_stage_opamp_dummy_magic_25_0.V_source.n28 two_stage_opamp_dummy_magic_25_0.V_source.n27 0.563
R23709 two_stage_opamp_dummy_magic_25_0.VD2.n15 two_stage_opamp_dummy_magic_25_0.VD2.n14 49.3505
R23710 two_stage_opamp_dummy_magic_25_0.VD2.n18 two_stage_opamp_dummy_magic_25_0.VD2.n17 49.3505
R23711 two_stage_opamp_dummy_magic_25_0.VD2.n4 two_stage_opamp_dummy_magic_25_0.VD2.n3 49.3505
R23712 two_stage_opamp_dummy_magic_25_0.VD2.n43 two_stage_opamp_dummy_magic_25_0.VD2.n42 49.3505
R23713 two_stage_opamp_dummy_magic_25_0.VD2.n9 two_stage_opamp_dummy_magic_25_0.VD2.n8 49.3505
R23714 two_stage_opamp_dummy_magic_25_0.VD2.n12 two_stage_opamp_dummy_magic_25_0.VD2.n11 49.3505
R23715 two_stage_opamp_dummy_magic_25_0.VD2.n25 two_stage_opamp_dummy_magic_25_0.VD2.n24 49.3505
R23716 two_stage_opamp_dummy_magic_25_0.VD2.n28 two_stage_opamp_dummy_magic_25_0.VD2.n27 49.3505
R23717 two_stage_opamp_dummy_magic_25_0.VD2.n32 two_stage_opamp_dummy_magic_25_0.VD2.n31 49.3505
R23718 two_stage_opamp_dummy_magic_25_0.VD2.n7 two_stage_opamp_dummy_magic_25_0.VD2.n6 49.3505
R23719 two_stage_opamp_dummy_magic_25_0.VD2.n39 two_stage_opamp_dummy_magic_25_0.VD2.n38 49.3505
R23720 two_stage_opamp_dummy_magic_25_0.VD2.n14 two_stage_opamp_dummy_magic_25_0.VD2.t17 16.0005
R23721 two_stage_opamp_dummy_magic_25_0.VD2.n14 two_stage_opamp_dummy_magic_25_0.VD2.t10 16.0005
R23722 two_stage_opamp_dummy_magic_25_0.VD2.n17 two_stage_opamp_dummy_magic_25_0.VD2.t15 16.0005
R23723 two_stage_opamp_dummy_magic_25_0.VD2.n17 two_stage_opamp_dummy_magic_25_0.VD2.t8 16.0005
R23724 two_stage_opamp_dummy_magic_25_0.VD2.n3 two_stage_opamp_dummy_magic_25_0.VD2.t11 16.0005
R23725 two_stage_opamp_dummy_magic_25_0.VD2.n3 two_stage_opamp_dummy_magic_25_0.VD2.t9 16.0005
R23726 two_stage_opamp_dummy_magic_25_0.VD2.n42 two_stage_opamp_dummy_magic_25_0.VD2.t14 16.0005
R23727 two_stage_opamp_dummy_magic_25_0.VD2.n42 two_stage_opamp_dummy_magic_25_0.VD2.t7 16.0005
R23728 two_stage_opamp_dummy_magic_25_0.VD2.n8 two_stage_opamp_dummy_magic_25_0.VD2.t1 16.0005
R23729 two_stage_opamp_dummy_magic_25_0.VD2.n8 two_stage_opamp_dummy_magic_25_0.VD2.t3 16.0005
R23730 two_stage_opamp_dummy_magic_25_0.VD2.n11 two_stage_opamp_dummy_magic_25_0.VD2.t19 16.0005
R23731 two_stage_opamp_dummy_magic_25_0.VD2.n11 two_stage_opamp_dummy_magic_25_0.VD2.t5 16.0005
R23732 two_stage_opamp_dummy_magic_25_0.VD2.n24 two_stage_opamp_dummy_magic_25_0.VD2.t6 16.0005
R23733 two_stage_opamp_dummy_magic_25_0.VD2.n24 two_stage_opamp_dummy_magic_25_0.VD2.t0 16.0005
R23734 two_stage_opamp_dummy_magic_25_0.VD2.n27 two_stage_opamp_dummy_magic_25_0.VD2.t21 16.0005
R23735 two_stage_opamp_dummy_magic_25_0.VD2.n27 two_stage_opamp_dummy_magic_25_0.VD2.t4 16.0005
R23736 two_stage_opamp_dummy_magic_25_0.VD2.n31 two_stage_opamp_dummy_magic_25_0.VD2.t2 16.0005
R23737 two_stage_opamp_dummy_magic_25_0.VD2.n31 two_stage_opamp_dummy_magic_25_0.VD2.t20 16.0005
R23738 two_stage_opamp_dummy_magic_25_0.VD2.n6 two_stage_opamp_dummy_magic_25_0.VD2.t12 16.0005
R23739 two_stage_opamp_dummy_magic_25_0.VD2.n6 two_stage_opamp_dummy_magic_25_0.VD2.t18 16.0005
R23740 two_stage_opamp_dummy_magic_25_0.VD2.n38 two_stage_opamp_dummy_magic_25_0.VD2.t13 16.0005
R23741 two_stage_opamp_dummy_magic_25_0.VD2.n38 two_stage_opamp_dummy_magic_25_0.VD2.t16 16.0005
R23742 two_stage_opamp_dummy_magic_25_0.VD2.n23 two_stage_opamp_dummy_magic_25_0.VD2.n13 6.2505
R23743 two_stage_opamp_dummy_magic_25_0.VD2.n33 two_stage_opamp_dummy_magic_25_0.VD2.n2 6.2505
R23744 two_stage_opamp_dummy_magic_25_0.VD2.n21 two_stage_opamp_dummy_magic_25_0.VD2.n20 6.2505
R23745 two_stage_opamp_dummy_magic_25_0.VD2.n36 two_stage_opamp_dummy_magic_25_0.VD2.n35 6.2505
R23746 two_stage_opamp_dummy_magic_25_0.VD2.n26 two_stage_opamp_dummy_magic_25_0.VD2.n12 5.6255
R23747 two_stage_opamp_dummy_magic_25_0.VD2.n30 two_stage_opamp_dummy_magic_25_0.VD2.n9 5.6255
R23748 two_stage_opamp_dummy_magic_25_0.VD2.n40 two_stage_opamp_dummy_magic_25_0.VD2.n7 5.438
R23749 two_stage_opamp_dummy_magic_25_0.VD2.n16 two_stage_opamp_dummy_magic_25_0.VD2.n15 5.438
R23750 two_stage_opamp_dummy_magic_25_0.VD2.n36 two_stage_opamp_dummy_magic_25_0.VD2.n7 5.31821
R23751 two_stage_opamp_dummy_magic_25_0.VD2.n20 two_stage_opamp_dummy_magic_25_0.VD2.n15 5.31821
R23752 two_stage_opamp_dummy_magic_25_0.VD2.n19 two_stage_opamp_dummy_magic_25_0.VD2.n18 5.08383
R23753 two_stage_opamp_dummy_magic_25_0.VD2.n4 two_stage_opamp_dummy_magic_25_0.VD2.n1 5.08383
R23754 two_stage_opamp_dummy_magic_25_0.VD2.n44 two_stage_opamp_dummy_magic_25_0.VD2.n43 5.08383
R23755 two_stage_opamp_dummy_magic_25_0.VD2.n39 two_stage_opamp_dummy_magic_25_0.VD2.n37 5.08383
R23756 two_stage_opamp_dummy_magic_25_0.VD2.n26 two_stage_opamp_dummy_magic_25_0.VD2.n25 5.063
R23757 two_stage_opamp_dummy_magic_25_0.VD2.n29 two_stage_opamp_dummy_magic_25_0.VD2.n28 5.063
R23758 two_stage_opamp_dummy_magic_25_0.VD2.n32 two_stage_opamp_dummy_magic_25_0.VD2.n30 5.063
R23759 two_stage_opamp_dummy_magic_25_0.VD2.n35 two_stage_opamp_dummy_magic_25_0.VD2.n34 5.063
R23760 two_stage_opamp_dummy_magic_25_0.VD2.n22 two_stage_opamp_dummy_magic_25_0.VD2.n21 5.063
R23761 two_stage_opamp_dummy_magic_25_0.VD2.n18 two_stage_opamp_dummy_magic_25_0.VD2.n16 4.8755
R23762 two_stage_opamp_dummy_magic_25_0.VD2.n5 two_stage_opamp_dummy_magic_25_0.VD2.n4 4.8755
R23763 two_stage_opamp_dummy_magic_25_0.VD2.n43 two_stage_opamp_dummy_magic_25_0.VD2.n41 4.8755
R23764 two_stage_opamp_dummy_magic_25_0.VD2.n40 two_stage_opamp_dummy_magic_25_0.VD2.n39 4.8755
R23765 two_stage_opamp_dummy_magic_25_0.VD2 two_stage_opamp_dummy_magic_25_0.VD2.n45 4.60467
R23766 two_stage_opamp_dummy_magic_25_0.VD2.n34 two_stage_opamp_dummy_magic_25_0.VD2.n33 4.5005
R23767 two_stage_opamp_dummy_magic_25_0.VD2.n10 two_stage_opamp_dummy_magic_25_0.VD2.n0 4.5005
R23768 two_stage_opamp_dummy_magic_25_0.VD2.n23 two_stage_opamp_dummy_magic_25_0.VD2.n22 4.5005
R23769 two_stage_opamp_dummy_magic_25_0.VD2 two_stage_opamp_dummy_magic_25_0.VD2.n0 1.64633
R23770 two_stage_opamp_dummy_magic_25_0.VD2.n34 two_stage_opamp_dummy_magic_25_0.VD2.n10 0.563
R23771 two_stage_opamp_dummy_magic_25_0.VD2.n22 two_stage_opamp_dummy_magic_25_0.VD2.n10 0.563
R23772 two_stage_opamp_dummy_magic_25_0.VD2.n29 two_stage_opamp_dummy_magic_25_0.VD2.n26 0.563
R23773 two_stage_opamp_dummy_magic_25_0.VD2.n30 two_stage_opamp_dummy_magic_25_0.VD2.n29 0.563
R23774 two_stage_opamp_dummy_magic_25_0.VD2.n16 two_stage_opamp_dummy_magic_25_0.VD2.n5 0.563
R23775 two_stage_opamp_dummy_magic_25_0.VD2.n41 two_stage_opamp_dummy_magic_25_0.VD2.n5 0.563
R23776 two_stage_opamp_dummy_magic_25_0.VD2.n41 two_stage_opamp_dummy_magic_25_0.VD2.n40 0.563
R23777 two_stage_opamp_dummy_magic_25_0.VD2.n25 two_stage_opamp_dummy_magic_25_0.VD2.n23 0.3755
R23778 two_stage_opamp_dummy_magic_25_0.VD2.n28 two_stage_opamp_dummy_magic_25_0.VD2.n0 0.3755
R23779 two_stage_opamp_dummy_magic_25_0.VD2.n33 two_stage_opamp_dummy_magic_25_0.VD2.n32 0.3755
R23780 two_stage_opamp_dummy_magic_25_0.VD2.n21 two_stage_opamp_dummy_magic_25_0.VD2.n12 0.3755
R23781 two_stage_opamp_dummy_magic_25_0.VD2.n35 two_stage_opamp_dummy_magic_25_0.VD2.n9 0.3755
R23782 two_stage_opamp_dummy_magic_25_0.VD2.n37 two_stage_opamp_dummy_magic_25_0.VD2.n36 0.234875
R23783 two_stage_opamp_dummy_magic_25_0.VD2.n37 two_stage_opamp_dummy_magic_25_0.VD2.n2 0.234875
R23784 two_stage_opamp_dummy_magic_25_0.VD2.n44 two_stage_opamp_dummy_magic_25_0.VD2.n2 0.234875
R23785 two_stage_opamp_dummy_magic_25_0.VD2.n45 two_stage_opamp_dummy_magic_25_0.VD2.n44 0.234875
R23786 two_stage_opamp_dummy_magic_25_0.VD2.n45 two_stage_opamp_dummy_magic_25_0.VD2.n1 0.234875
R23787 two_stage_opamp_dummy_magic_25_0.VD2.n13 two_stage_opamp_dummy_magic_25_0.VD2.n1 0.234875
R23788 two_stage_opamp_dummy_magic_25_0.VD2.n19 two_stage_opamp_dummy_magic_25_0.VD2.n13 0.234875
R23789 two_stage_opamp_dummy_magic_25_0.VD2.n20 two_stage_opamp_dummy_magic_25_0.VD2.n19 0.234875
R23790 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.n15 325.473
R23791 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.n8 325.473
R23792 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.n3 325.473
R23793 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t15 310.488
R23794 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t14 310.488
R23795 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t13 310.488
R23796 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.t10 184.097
R23797 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.t0 184.097
R23798 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.t2 184.097
R23799 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.n12 167.094
R23800 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.n5 167.094
R23801 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.n0 167.094
R23802 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.n7 152
R23803 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.n2 152
R23804 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n14 152
R23805 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t17 120.501
R23806 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.t4 120.501
R23807 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t18 120.501
R23808 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.t8 120.501
R23809 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t16 120.501
R23810 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.t6 120.501
R23811 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.t12 106.933
R23812 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.n13 40.7027
R23813 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.n6 40.7027
R23814 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.n1 40.7027
R23815 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.t9 39.4005
R23816 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.t1 39.4005
R23817 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.t7 39.4005
R23818 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.t3 39.4005
R23819 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.t5 39.4005
R23820 bgr_11_0.V_mir2.t11 bgr_11_0.V_mir2.n16 39.4005
R23821 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n4 15.9255
R23822 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n11 15.9255
R23823 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.n9 9.3005
R23824 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n10 4.5005
R23825 two_stage_opamp_dummy_magic_25_0.Vb1.n8 two_stage_opamp_dummy_magic_25_0.Vb1.t6 449.868
R23826 two_stage_opamp_dummy_magic_25_0.Vb1.n7 two_stage_opamp_dummy_magic_25_0.Vb1.t4 449.868
R23827 two_stage_opamp_dummy_magic_25_0.Vb1.n14 two_stage_opamp_dummy_magic_25_0.Vb1.t20 449.868
R23828 two_stage_opamp_dummy_magic_25_0.Vb1.n33 two_stage_opamp_dummy_magic_25_0.Vb1.n32 435.659
R23829 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.Vb1.n22 433.519
R23830 two_stage_opamp_dummy_magic_25_0.Vb1.n23 two_stage_opamp_dummy_magic_25_0.Vb1 433.519
R23831 two_stage_opamp_dummy_magic_25_0.Vb1.n8 two_stage_opamp_dummy_magic_25_0.Vb1.t0 273.134
R23832 two_stage_opamp_dummy_magic_25_0.Vb1.n7 two_stage_opamp_dummy_magic_25_0.Vb1.t2 273.134
R23833 two_stage_opamp_dummy_magic_25_0.Vb1.n32 two_stage_opamp_dummy_magic_25_0.Vb1.t14 273.134
R23834 two_stage_opamp_dummy_magic_25_0.Vb1.n23 two_stage_opamp_dummy_magic_25_0.Vb1.t21 273.134
R23835 two_stage_opamp_dummy_magic_25_0.Vb1.n22 two_stage_opamp_dummy_magic_25_0.Vb1.t19 273.134
R23836 two_stage_opamp_dummy_magic_25_0.Vb1.n21 two_stage_opamp_dummy_magic_25_0.Vb1.t29 273.134
R23837 two_stage_opamp_dummy_magic_25_0.Vb1.n20 two_stage_opamp_dummy_magic_25_0.Vb1.t18 273.134
R23838 two_stage_opamp_dummy_magic_25_0.Vb1.n19 two_stage_opamp_dummy_magic_25_0.Vb1.t27 273.134
R23839 two_stage_opamp_dummy_magic_25_0.Vb1.n18 two_stage_opamp_dummy_magic_25_0.Vb1.t15 273.134
R23840 two_stage_opamp_dummy_magic_25_0.Vb1.n17 two_stage_opamp_dummy_magic_25_0.Vb1.t28 273.134
R23841 two_stage_opamp_dummy_magic_25_0.Vb1.n16 two_stage_opamp_dummy_magic_25_0.Vb1.t16 273.134
R23842 two_stage_opamp_dummy_magic_25_0.Vb1.n15 two_stage_opamp_dummy_magic_25_0.Vb1.t26 273.134
R23843 two_stage_opamp_dummy_magic_25_0.Vb1.n14 two_stage_opamp_dummy_magic_25_0.Vb1.t13 273.134
R23844 two_stage_opamp_dummy_magic_25_0.Vb1.n31 two_stage_opamp_dummy_magic_25_0.Vb1.t25 273.134
R23845 two_stage_opamp_dummy_magic_25_0.Vb1.n30 two_stage_opamp_dummy_magic_25_0.Vb1.t32 273.134
R23846 two_stage_opamp_dummy_magic_25_0.Vb1.n29 two_stage_opamp_dummy_magic_25_0.Vb1.t24 273.134
R23847 two_stage_opamp_dummy_magic_25_0.Vb1.n28 two_stage_opamp_dummy_magic_25_0.Vb1.t31 273.134
R23848 two_stage_opamp_dummy_magic_25_0.Vb1.n27 two_stage_opamp_dummy_magic_25_0.Vb1.t22 273.134
R23849 two_stage_opamp_dummy_magic_25_0.Vb1.n26 two_stage_opamp_dummy_magic_25_0.Vb1.t17 273.134
R23850 two_stage_opamp_dummy_magic_25_0.Vb1.n25 two_stage_opamp_dummy_magic_25_0.Vb1.t23 273.134
R23851 two_stage_opamp_dummy_magic_25_0.Vb1.n24 two_stage_opamp_dummy_magic_25_0.Vb1.t30 273.134
R23852 two_stage_opamp_dummy_magic_25_0.Vb1.n15 two_stage_opamp_dummy_magic_25_0.Vb1.n14 176.733
R23853 two_stage_opamp_dummy_magic_25_0.Vb1.n16 two_stage_opamp_dummy_magic_25_0.Vb1.n15 176.733
R23854 two_stage_opamp_dummy_magic_25_0.Vb1.n17 two_stage_opamp_dummy_magic_25_0.Vb1.n16 176.733
R23855 two_stage_opamp_dummy_magic_25_0.Vb1.n18 two_stage_opamp_dummy_magic_25_0.Vb1.n17 176.733
R23856 two_stage_opamp_dummy_magic_25_0.Vb1.n19 two_stage_opamp_dummy_magic_25_0.Vb1.n18 176.733
R23857 two_stage_opamp_dummy_magic_25_0.Vb1.n20 two_stage_opamp_dummy_magic_25_0.Vb1.n19 176.733
R23858 two_stage_opamp_dummy_magic_25_0.Vb1.n21 two_stage_opamp_dummy_magic_25_0.Vb1.n20 176.733
R23859 two_stage_opamp_dummy_magic_25_0.Vb1.n22 two_stage_opamp_dummy_magic_25_0.Vb1.n21 176.733
R23860 two_stage_opamp_dummy_magic_25_0.Vb1.n24 two_stage_opamp_dummy_magic_25_0.Vb1.n23 176.733
R23861 two_stage_opamp_dummy_magic_25_0.Vb1.n25 two_stage_opamp_dummy_magic_25_0.Vb1.n24 176.733
R23862 two_stage_opamp_dummy_magic_25_0.Vb1.n26 two_stage_opamp_dummy_magic_25_0.Vb1.n25 176.733
R23863 two_stage_opamp_dummy_magic_25_0.Vb1.n27 two_stage_opamp_dummy_magic_25_0.Vb1.n26 176.733
R23864 two_stage_opamp_dummy_magic_25_0.Vb1.n28 two_stage_opamp_dummy_magic_25_0.Vb1.n27 176.733
R23865 two_stage_opamp_dummy_magic_25_0.Vb1.n29 two_stage_opamp_dummy_magic_25_0.Vb1.n28 176.733
R23866 two_stage_opamp_dummy_magic_25_0.Vb1.n30 two_stage_opamp_dummy_magic_25_0.Vb1.n29 176.733
R23867 two_stage_opamp_dummy_magic_25_0.Vb1.n31 two_stage_opamp_dummy_magic_25_0.Vb1.n30 176.733
R23868 two_stage_opamp_dummy_magic_25_0.Vb1.n32 two_stage_opamp_dummy_magic_25_0.Vb1.n31 176.733
R23869 two_stage_opamp_dummy_magic_25_0.Vb1.n3 two_stage_opamp_dummy_magic_25_0.Vb1.t12 166.847
R23870 two_stage_opamp_dummy_magic_25_0.Vb1.t12 two_stage_opamp_dummy_magic_25_0.Vb1.n5 166.847
R23871 two_stage_opamp_dummy_magic_25_0.Vb1.n0 two_stage_opamp_dummy_magic_25_0.Vb1.n9 161.3
R23872 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.Vb1.n6 151.863
R23873 two_stage_opamp_dummy_magic_25_0.Vb1.n0 two_stage_opamp_dummy_magic_25_0.Vb1.n12 49.3505
R23874 two_stage_opamp_dummy_magic_25_0.Vb1.n11 two_stage_opamp_dummy_magic_25_0.Vb1.n10 49.3505
R23875 two_stage_opamp_dummy_magic_25_0.Vb1.n9 two_stage_opamp_dummy_magic_25_0.Vb1.n8 45.5227
R23876 two_stage_opamp_dummy_magic_25_0.Vb1.n9 two_stage_opamp_dummy_magic_25_0.Vb1.n7 45.5227
R23877 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.Vb1.n33 36.6255
R23878 two_stage_opamp_dummy_magic_25_0.Vb1.n6 two_stage_opamp_dummy_magic_25_0.Vb1.t11 19.7005
R23879 two_stage_opamp_dummy_magic_25_0.Vb1.n6 two_stage_opamp_dummy_magic_25_0.Vb1.t8 19.7005
R23880 two_stage_opamp_dummy_magic_25_0.Vb1.n12 two_stage_opamp_dummy_magic_25_0.Vb1.t3 16.0005
R23881 two_stage_opamp_dummy_magic_25_0.Vb1.n12 two_stage_opamp_dummy_magic_25_0.Vb1.t1 16.0005
R23882 two_stage_opamp_dummy_magic_25_0.Vb1.n10 two_stage_opamp_dummy_magic_25_0.Vb1.t9 16.0005
R23883 two_stage_opamp_dummy_magic_25_0.Vb1.n10 two_stage_opamp_dummy_magic_25_0.Vb1.t5 16.0005
R23884 two_stage_opamp_dummy_magic_25_0.Vb1.n13 two_stage_opamp_dummy_magic_25_0.Vb1.t7 16.0005
R23885 two_stage_opamp_dummy_magic_25_0.Vb1.n13 two_stage_opamp_dummy_magic_25_0.Vb1.t10 16.0005
R23886 two_stage_opamp_dummy_magic_25_0.Vb1.n1 two_stage_opamp_dummy_magic_25_0.Vb1.n0 4.938
R23887 two_stage_opamp_dummy_magic_25_0.Vb1.n13 two_stage_opamp_dummy_magic_25_0.Vb1.n2 51.6321
R23888 two_stage_opamp_dummy_magic_25_0.Vb1.n11 two_stage_opamp_dummy_magic_25_0.Vb1.n5 4.938
R23889 two_stage_opamp_dummy_magic_25_0.Vb1.n3 two_stage_opamp_dummy_magic_25_0.Vb1.n11 4.938
R23890 two_stage_opamp_dummy_magic_25_0.Vb1.n0 two_stage_opamp_dummy_magic_25_0.Vb1.n4 4.938
R23891 two_stage_opamp_dummy_magic_25_0.Vb1.n1 two_stage_opamp_dummy_magic_25_0.Vb1.n2 0.376365
R23892 two_stage_opamp_dummy_magic_25_0.Vb1.n33 two_stage_opamp_dummy_magic_25_0.Vb1.n1 4.90706
R23893 two_stage_opamp_dummy_magic_25_0.Vb1.n2 two_stage_opamp_dummy_magic_25_0.Vb1.n4 0.376365
R23894 two_stage_opamp_dummy_magic_25_0.Vb1.n1 two_stage_opamp_dummy_magic_25_0.Vb1.n5 0.688
R23895 two_stage_opamp_dummy_magic_25_0.Vb1.n4 two_stage_opamp_dummy_magic_25_0.Vb1.n3 0.688
R23896 two_stage_opamp_dummy_magic_25_0.Vb1_2.n1 two_stage_opamp_dummy_magic_25_0.Vb1_2.t4 65.3505
R23897 two_stage_opamp_dummy_magic_25_0.Vb1_2.n3 two_stage_opamp_dummy_magic_25_0.Vb1_2.n2 49.3505
R23898 two_stage_opamp_dummy_magic_25_0.Vb1_2.n6 two_stage_opamp_dummy_magic_25_0.Vb1_2.n5 49.3505
R23899 two_stage_opamp_dummy_magic_25_0.Vb1_2.n2 two_stage_opamp_dummy_magic_25_0.Vb1_2.t2 16.0005
R23900 two_stage_opamp_dummy_magic_25_0.Vb1_2.n2 two_stage_opamp_dummy_magic_25_0.Vb1_2.t0 16.0005
R23901 two_stage_opamp_dummy_magic_25_0.Vb1_2.t3 two_stage_opamp_dummy_magic_25_0.Vb1_2.n6 16.0005
R23902 two_stage_opamp_dummy_magic_25_0.Vb1_2.n6 two_stage_opamp_dummy_magic_25_0.Vb1_2.t1 16.0005
R23903 two_stage_opamp_dummy_magic_25_0.Vb1_2.n1 two_stage_opamp_dummy_magic_25_0.Vb1_2.n0 6.41717
R23904 two_stage_opamp_dummy_magic_25_0.Vb1_2.n4 two_stage_opamp_dummy_magic_25_0.Vb1_2.n1 5.85467
R23905 two_stage_opamp_dummy_magic_25_0.Vb1_2.n3 two_stage_opamp_dummy_magic_25_0.Vb1_2.n0 5.72967
R23906 two_stage_opamp_dummy_magic_25_0.Vb1_2.n4 two_stage_opamp_dummy_magic_25_0.Vb1_2.n3 5.51092
R23907 two_stage_opamp_dummy_magic_25_0.Vb1_2.n5 two_stage_opamp_dummy_magic_25_0.Vb1_2.n0 5.16717
R23908 two_stage_opamp_dummy_magic_25_0.Vb1_2.n5 two_stage_opamp_dummy_magic_25_0.Vb1_2.n4 5.16717
R23909 two_stage_opamp_dummy_magic_25_0.Y.n74 two_stage_opamp_dummy_magic_25_0.Y.t48 1172.87
R23910 two_stage_opamp_dummy_magic_25_0.Y.n70 two_stage_opamp_dummy_magic_25_0.Y.t39 1172.87
R23911 two_stage_opamp_dummy_magic_25_0.Y.n74 two_stage_opamp_dummy_magic_25_0.Y.t40 996.134
R23912 two_stage_opamp_dummy_magic_25_0.Y.n75 two_stage_opamp_dummy_magic_25_0.Y.t28 996.134
R23913 two_stage_opamp_dummy_magic_25_0.Y.n76 two_stage_opamp_dummy_magic_25_0.Y.t44 996.134
R23914 two_stage_opamp_dummy_magic_25_0.Y.n77 two_stage_opamp_dummy_magic_25_0.Y.t30 996.134
R23915 two_stage_opamp_dummy_magic_25_0.Y.n73 two_stage_opamp_dummy_magic_25_0.Y.t47 996.134
R23916 two_stage_opamp_dummy_magic_25_0.Y.n72 two_stage_opamp_dummy_magic_25_0.Y.t52 996.134
R23917 two_stage_opamp_dummy_magic_25_0.Y.n71 two_stage_opamp_dummy_magic_25_0.Y.t35 996.134
R23918 two_stage_opamp_dummy_magic_25_0.Y.n70 two_stage_opamp_dummy_magic_25_0.Y.t25 996.134
R23919 two_stage_opamp_dummy_magic_25_0.Y.n46 two_stage_opamp_dummy_magic_25_0.Y.t43 690.867
R23920 two_stage_opamp_dummy_magic_25_0.Y.n39 two_stage_opamp_dummy_magic_25_0.Y.t33 690.867
R23921 two_stage_opamp_dummy_magic_25_0.Y.n55 two_stage_opamp_dummy_magic_25_0.Y.t46 530.201
R23922 two_stage_opamp_dummy_magic_25_0.Y.n48 two_stage_opamp_dummy_magic_25_0.Y.t36 530.201
R23923 two_stage_opamp_dummy_magic_25_0.Y.n46 two_stage_opamp_dummy_magic_25_0.Y.t34 514.134
R23924 two_stage_opamp_dummy_magic_25_0.Y.n39 two_stage_opamp_dummy_magic_25_0.Y.t51 514.134
R23925 two_stage_opamp_dummy_magic_25_0.Y.n40 two_stage_opamp_dummy_magic_25_0.Y.t31 514.134
R23926 two_stage_opamp_dummy_magic_25_0.Y.n41 two_stage_opamp_dummy_magic_25_0.Y.t49 514.134
R23927 two_stage_opamp_dummy_magic_25_0.Y.n42 two_stage_opamp_dummy_magic_25_0.Y.t42 514.134
R23928 two_stage_opamp_dummy_magic_25_0.Y.n43 two_stage_opamp_dummy_magic_25_0.Y.t27 514.134
R23929 two_stage_opamp_dummy_magic_25_0.Y.n44 two_stage_opamp_dummy_magic_25_0.Y.t38 514.134
R23930 two_stage_opamp_dummy_magic_25_0.Y.n45 two_stage_opamp_dummy_magic_25_0.Y.t54 514.134
R23931 two_stage_opamp_dummy_magic_25_0.Y.n55 two_stage_opamp_dummy_magic_25_0.Y.t37 353.467
R23932 two_stage_opamp_dummy_magic_25_0.Y.n54 two_stage_opamp_dummy_magic_25_0.Y.t26 353.467
R23933 two_stage_opamp_dummy_magic_25_0.Y.n53 two_stage_opamp_dummy_magic_25_0.Y.t41 353.467
R23934 two_stage_opamp_dummy_magic_25_0.Y.n52 two_stage_opamp_dummy_magic_25_0.Y.t29 353.467
R23935 two_stage_opamp_dummy_magic_25_0.Y.n51 two_stage_opamp_dummy_magic_25_0.Y.t45 353.467
R23936 two_stage_opamp_dummy_magic_25_0.Y.n50 two_stage_opamp_dummy_magic_25_0.Y.t50 353.467
R23937 two_stage_opamp_dummy_magic_25_0.Y.n49 two_stage_opamp_dummy_magic_25_0.Y.t32 353.467
R23938 two_stage_opamp_dummy_magic_25_0.Y.n48 two_stage_opamp_dummy_magic_25_0.Y.t53 353.467
R23939 two_stage_opamp_dummy_magic_25_0.Y.n73 two_stage_opamp_dummy_magic_25_0.Y.n72 176.733
R23940 two_stage_opamp_dummy_magic_25_0.Y.n72 two_stage_opamp_dummy_magic_25_0.Y.n71 176.733
R23941 two_stage_opamp_dummy_magic_25_0.Y.n71 two_stage_opamp_dummy_magic_25_0.Y.n70 176.733
R23942 two_stage_opamp_dummy_magic_25_0.Y.n75 two_stage_opamp_dummy_magic_25_0.Y.n74 176.733
R23943 two_stage_opamp_dummy_magic_25_0.Y.n76 two_stage_opamp_dummy_magic_25_0.Y.n75 176.733
R23944 two_stage_opamp_dummy_magic_25_0.Y.n77 two_stage_opamp_dummy_magic_25_0.Y.n76 176.733
R23945 two_stage_opamp_dummy_magic_25_0.Y.n54 two_stage_opamp_dummy_magic_25_0.Y.n53 176.733
R23946 two_stage_opamp_dummy_magic_25_0.Y.n53 two_stage_opamp_dummy_magic_25_0.Y.n52 176.733
R23947 two_stage_opamp_dummy_magic_25_0.Y.n52 two_stage_opamp_dummy_magic_25_0.Y.n51 176.733
R23948 two_stage_opamp_dummy_magic_25_0.Y.n51 two_stage_opamp_dummy_magic_25_0.Y.n50 176.733
R23949 two_stage_opamp_dummy_magic_25_0.Y.n50 two_stage_opamp_dummy_magic_25_0.Y.n49 176.733
R23950 two_stage_opamp_dummy_magic_25_0.Y.n49 two_stage_opamp_dummy_magic_25_0.Y.n48 176.733
R23951 two_stage_opamp_dummy_magic_25_0.Y.n45 two_stage_opamp_dummy_magic_25_0.Y.n44 176.733
R23952 two_stage_opamp_dummy_magic_25_0.Y.n44 two_stage_opamp_dummy_magic_25_0.Y.n43 176.733
R23953 two_stage_opamp_dummy_magic_25_0.Y.n43 two_stage_opamp_dummy_magic_25_0.Y.n42 176.733
R23954 two_stage_opamp_dummy_magic_25_0.Y.n42 two_stage_opamp_dummy_magic_25_0.Y.n41 176.733
R23955 two_stage_opamp_dummy_magic_25_0.Y.n41 two_stage_opamp_dummy_magic_25_0.Y.n40 176.733
R23956 two_stage_opamp_dummy_magic_25_0.Y.n40 two_stage_opamp_dummy_magic_25_0.Y.n39 176.733
R23957 two_stage_opamp_dummy_magic_25_0.Y.n57 two_stage_opamp_dummy_magic_25_0.Y.n56 165.472
R23958 two_stage_opamp_dummy_magic_25_0.Y.n57 two_stage_opamp_dummy_magic_25_0.Y.n47 165.472
R23959 two_stage_opamp_dummy_magic_25_0.Y.n80 two_stage_opamp_dummy_magic_25_0.Y.n79 152
R23960 two_stage_opamp_dummy_magic_25_0.Y.n81 two_stage_opamp_dummy_magic_25_0.Y.n80 131.571
R23961 two_stage_opamp_dummy_magic_25_0.Y.n80 two_stage_opamp_dummy_magic_25_0.Y.n78 124.517
R23962 two_stage_opamp_dummy_magic_25_0.Y.n147 two_stage_opamp_dummy_magic_25_0.Y.n57 74.5372
R23963 two_stage_opamp_dummy_magic_25_0.Y.n107 two_stage_opamp_dummy_magic_25_0.Y.n106 66.0338
R23964 two_stage_opamp_dummy_magic_25_0.Y.n98 two_stage_opamp_dummy_magic_25_0.Y.n97 66.0338
R23965 two_stage_opamp_dummy_magic_25_0.Y.n96 two_stage_opamp_dummy_magic_25_0.Y.n95 66.0338
R23966 two_stage_opamp_dummy_magic_25_0.Y.n101 two_stage_opamp_dummy_magic_25_0.Y.n100 66.0338
R23967 two_stage_opamp_dummy_magic_25_0.Y.n104 two_stage_opamp_dummy_magic_25_0.Y.n103 66.0338
R23968 two_stage_opamp_dummy_magic_25_0.Y.n110 two_stage_opamp_dummy_magic_25_0.Y.n109 66.0338
R23969 two_stage_opamp_dummy_magic_25_0.Y.n7 two_stage_opamp_dummy_magic_25_0.Y.n6 49.3505
R23970 two_stage_opamp_dummy_magic_25_0.Y.n11 two_stage_opamp_dummy_magic_25_0.Y.n10 49.3505
R23971 two_stage_opamp_dummy_magic_25_0.Y.n20 two_stage_opamp_dummy_magic_25_0.Y.n19 49.3505
R23972 two_stage_opamp_dummy_magic_25_0.Y.n30 two_stage_opamp_dummy_magic_25_0.Y.n29 49.3505
R23973 two_stage_opamp_dummy_magic_25_0.Y.n26 two_stage_opamp_dummy_magic_25_0.Y.n25 49.3505
R23974 two_stage_opamp_dummy_magic_25_0.Y.n23 two_stage_opamp_dummy_magic_25_0.Y.n22 49.3505
R23975 two_stage_opamp_dummy_magic_25_0.Y.n64 two_stage_opamp_dummy_magic_25_0.Y.t20 41.0384
R23976 two_stage_opamp_dummy_magic_25_0.Y.n78 two_stage_opamp_dummy_magic_25_0.Y.n73 40.1672
R23977 two_stage_opamp_dummy_magic_25_0.Y.n78 two_stage_opamp_dummy_magic_25_0.Y.n77 40.1672
R23978 two_stage_opamp_dummy_magic_25_0.Y.n56 two_stage_opamp_dummy_magic_25_0.Y.n54 40.1672
R23979 two_stage_opamp_dummy_magic_25_0.Y.n56 two_stage_opamp_dummy_magic_25_0.Y.n55 40.1672
R23980 two_stage_opamp_dummy_magic_25_0.Y.n47 two_stage_opamp_dummy_magic_25_0.Y.n45 40.1672
R23981 two_stage_opamp_dummy_magic_25_0.Y.n47 two_stage_opamp_dummy_magic_25_0.Y.n46 40.1672
R23982 two_stage_opamp_dummy_magic_25_0.Y.n82 two_stage_opamp_dummy_magic_25_0.Y.n81 16.3217
R23983 two_stage_opamp_dummy_magic_25_0.Y.n6 two_stage_opamp_dummy_magic_25_0.Y.t9 16.0005
R23984 two_stage_opamp_dummy_magic_25_0.Y.n6 two_stage_opamp_dummy_magic_25_0.Y.t22 16.0005
R23985 two_stage_opamp_dummy_magic_25_0.Y.n10 two_stage_opamp_dummy_magic_25_0.Y.t21 16.0005
R23986 two_stage_opamp_dummy_magic_25_0.Y.n10 two_stage_opamp_dummy_magic_25_0.Y.t7 16.0005
R23987 two_stage_opamp_dummy_magic_25_0.Y.n19 two_stage_opamp_dummy_magic_25_0.Y.t2 16.0005
R23988 two_stage_opamp_dummy_magic_25_0.Y.n19 two_stage_opamp_dummy_magic_25_0.Y.t5 16.0005
R23989 two_stage_opamp_dummy_magic_25_0.Y.n29 two_stage_opamp_dummy_magic_25_0.Y.t8 16.0005
R23990 two_stage_opamp_dummy_magic_25_0.Y.n29 two_stage_opamp_dummy_magic_25_0.Y.t6 16.0005
R23991 two_stage_opamp_dummy_magic_25_0.Y.n25 two_stage_opamp_dummy_magic_25_0.Y.t1 16.0005
R23992 two_stage_opamp_dummy_magic_25_0.Y.n25 two_stage_opamp_dummy_magic_25_0.Y.t4 16.0005
R23993 two_stage_opamp_dummy_magic_25_0.Y.n22 two_stage_opamp_dummy_magic_25_0.Y.t0 16.0005
R23994 two_stage_opamp_dummy_magic_25_0.Y.n22 two_stage_opamp_dummy_magic_25_0.Y.t3 16.0005
R23995 two_stage_opamp_dummy_magic_25_0.Y.n79 two_stage_opamp_dummy_magic_25_0.Y.n69 12.8005
R23996 two_stage_opamp_dummy_magic_25_0.Y.n106 two_stage_opamp_dummy_magic_25_0.Y.t16 11.2576
R23997 two_stage_opamp_dummy_magic_25_0.Y.n106 two_stage_opamp_dummy_magic_25_0.Y.t24 11.2576
R23998 two_stage_opamp_dummy_magic_25_0.Y.n97 two_stage_opamp_dummy_magic_25_0.Y.t23 11.2576
R23999 two_stage_opamp_dummy_magic_25_0.Y.n97 two_stage_opamp_dummy_magic_25_0.Y.t12 11.2576
R24000 two_stage_opamp_dummy_magic_25_0.Y.n95 two_stage_opamp_dummy_magic_25_0.Y.t14 11.2576
R24001 two_stage_opamp_dummy_magic_25_0.Y.n95 two_stage_opamp_dummy_magic_25_0.Y.t17 11.2576
R24002 two_stage_opamp_dummy_magic_25_0.Y.n100 two_stage_opamp_dummy_magic_25_0.Y.t19 11.2576
R24003 two_stage_opamp_dummy_magic_25_0.Y.n100 two_stage_opamp_dummy_magic_25_0.Y.t10 11.2576
R24004 two_stage_opamp_dummy_magic_25_0.Y.n103 two_stage_opamp_dummy_magic_25_0.Y.t11 11.2576
R24005 two_stage_opamp_dummy_magic_25_0.Y.n103 two_stage_opamp_dummy_magic_25_0.Y.t13 11.2576
R24006 two_stage_opamp_dummy_magic_25_0.Y.n109 two_stage_opamp_dummy_magic_25_0.Y.t15 11.2576
R24007 two_stage_opamp_dummy_magic_25_0.Y.n109 two_stage_opamp_dummy_magic_25_0.Y.t18 11.2576
R24008 two_stage_opamp_dummy_magic_25_0.Y.n79 two_stage_opamp_dummy_magic_25_0.Y.n67 9.36264
R24009 two_stage_opamp_dummy_magic_25_0.Y.n69 two_stage_opamp_dummy_magic_25_0.Y.n68 9.3005
R24010 two_stage_opamp_dummy_magic_25_0.Y.n99 two_stage_opamp_dummy_magic_25_0.Y.n98 5.91717
R24011 two_stage_opamp_dummy_magic_25_0.Y.n108 two_stage_opamp_dummy_magic_25_0.Y.n107 5.91717
R24012 two_stage_opamp_dummy_magic_25_0.Y.n21 two_stage_opamp_dummy_magic_25_0.Y.n11 5.6255
R24013 two_stage_opamp_dummy_magic_25_0.Y.n24 two_stage_opamp_dummy_magic_25_0.Y.n7 5.6255
R24014 two_stage_opamp_dummy_magic_25_0.Y.n81 two_stage_opamp_dummy_magic_25_0.Y.n69 5.33141
R24015 two_stage_opamp_dummy_magic_25_0.Y.n99 two_stage_opamp_dummy_magic_25_0.Y.n96 5.29217
R24016 two_stage_opamp_dummy_magic_25_0.Y.n102 two_stage_opamp_dummy_magic_25_0.Y.n101 5.29217
R24017 two_stage_opamp_dummy_magic_25_0.Y.n105 two_stage_opamp_dummy_magic_25_0.Y.n104 5.29217
R24018 two_stage_opamp_dummy_magic_25_0.Y.n110 two_stage_opamp_dummy_magic_25_0.Y.n108 5.29217
R24019 two_stage_opamp_dummy_magic_25_0.Y.n112 two_stage_opamp_dummy_magic_25_0.Y.n86 5.1255
R24020 two_stage_opamp_dummy_magic_25_0.Y.n115 two_stage_opamp_dummy_magic_25_0.Y.n94 5.1255
R24021 two_stage_opamp_dummy_magic_25_0.Y.n21 two_stage_opamp_dummy_magic_25_0.Y.n20 5.063
R24022 two_stage_opamp_dummy_magic_25_0.Y.n30 two_stage_opamp_dummy_magic_25_0.Y.n28 5.063
R24023 two_stage_opamp_dummy_magic_25_0.Y.n27 two_stage_opamp_dummy_magic_25_0.Y.n26 5.063
R24024 two_stage_opamp_dummy_magic_25_0.Y.n24 two_stage_opamp_dummy_magic_25_0.Y.n23 5.063
R24025 two_stage_opamp_dummy_magic_25_0.Y.n35 two_stage_opamp_dummy_magic_25_0.Y.n34 5.063
R24026 two_stage_opamp_dummy_magic_25_0.Y.n12 two_stage_opamp_dummy_magic_25_0.Y.n8 5.063
R24027 two_stage_opamp_dummy_magic_25_0.Y.n112 two_stage_opamp_dummy_magic_25_0.Y.n111 4.5005
R24028 two_stage_opamp_dummy_magic_25_0.Y.n113 two_stage_opamp_dummy_magic_25_0.Y.n89 4.5005
R24029 two_stage_opamp_dummy_magic_25_0.Y.n114 two_stage_opamp_dummy_magic_25_0.Y.n92 4.5005
R24030 two_stage_opamp_dummy_magic_25_0.Y.n116 two_stage_opamp_dummy_magic_25_0.Y.n115 4.5005
R24031 two_stage_opamp_dummy_magic_25_0.Y.n141 two_stage_opamp_dummy_magic_25_0.Y.n140 4.5005
R24032 two_stage_opamp_dummy_magic_25_0.Y.n34 two_stage_opamp_dummy_magic_25_0.Y.n5 4.5005
R24033 two_stage_opamp_dummy_magic_25_0.Y.n33 two_stage_opamp_dummy_magic_25_0.Y.n1 4.5005
R24034 two_stage_opamp_dummy_magic_25_0.Y.n32 two_stage_opamp_dummy_magic_25_0.Y.n31 4.5005
R24035 two_stage_opamp_dummy_magic_25_0.Y.n18 two_stage_opamp_dummy_magic_25_0.Y.n8 4.5005
R24036 two_stage_opamp_dummy_magic_25_0.Y.n148 two_stage_opamp_dummy_magic_25_0.Y.n36 4.5005
R24037 two_stage_opamp_dummy_magic_25_0.Y.n147 two_stage_opamp_dummy_magic_25_0.Y.n146 4.5005
R24038 two_stage_opamp_dummy_magic_25_0.Y.n148 two_stage_opamp_dummy_magic_25_0.Y.n147 4.5005
R24039 two_stage_opamp_dummy_magic_25_0.Y.n83 two_stage_opamp_dummy_magic_25_0.Y.n82 4.5005
R24040 two_stage_opamp_dummy_magic_25_0.Y.n61 two_stage_opamp_dummy_magic_25_0.Y.n60 4.5005
R24041 two_stage_opamp_dummy_magic_25_0.Y.n62 two_stage_opamp_dummy_magic_25_0.Y.n59 2.26187
R24042 two_stage_opamp_dummy_magic_25_0.Y.n138 two_stage_opamp_dummy_magic_25_0.Y.n84 2.26187
R24043 two_stage_opamp_dummy_magic_25_0.Y.n139 two_stage_opamp_dummy_magic_25_0.Y.n138 2.26187
R24044 two_stage_opamp_dummy_magic_25_0.Y.n63 two_stage_opamp_dummy_magic_25_0.Y.n62 2.26187
R24045 two_stage_opamp_dummy_magic_25_0.Y.n142 two_stage_opamp_dummy_magic_25_0.Y.n137 2.24063
R24046 two_stage_opamp_dummy_magic_25_0.Y.n143 two_stage_opamp_dummy_magic_25_0.Y.n84 2.24063
R24047 two_stage_opamp_dummy_magic_25_0.Y.n146 two_stage_opamp_dummy_magic_25_0.Y.n145 2.24063
R24048 two_stage_opamp_dummy_magic_25_0.Y.n58 two_stage_opamp_dummy_magic_25_0.Y.n38 2.24063
R24049 two_stage_opamp_dummy_magic_25_0.Y.n66 two_stage_opamp_dummy_magic_25_0.Y.n59 2.24063
R24050 two_stage_opamp_dummy_magic_25_0.Y.n144 two_stage_opamp_dummy_magic_25_0.Y.n37 2.24063
R24051 two_stage_opamp_dummy_magic_25_0.Y.n65 two_stage_opamp_dummy_magic_25_0.Y.n64 2.24063
R24052 two_stage_opamp_dummy_magic_25_0.Y.n83 two_stage_opamp_dummy_magic_25_0.Y.n67 2.22018
R24053 two_stage_opamp_dummy_magic_25_0.Y.n136 two_stage_opamp_dummy_magic_25_0.Y.n135 1.5005
R24054 two_stage_opamp_dummy_magic_25_0.Y.n134 two_stage_opamp_dummy_magic_25_0.Y.n85 1.5005
R24055 two_stage_opamp_dummy_magic_25_0.Y.n133 two_stage_opamp_dummy_magic_25_0.Y.n132 1.5005
R24056 two_stage_opamp_dummy_magic_25_0.Y.n131 two_stage_opamp_dummy_magic_25_0.Y.n87 1.5005
R24057 two_stage_opamp_dummy_magic_25_0.Y.n130 two_stage_opamp_dummy_magic_25_0.Y.n129 1.5005
R24058 two_stage_opamp_dummy_magic_25_0.Y.n128 two_stage_opamp_dummy_magic_25_0.Y.n88 1.5005
R24059 two_stage_opamp_dummy_magic_25_0.Y.n127 two_stage_opamp_dummy_magic_25_0.Y.n126 1.5005
R24060 two_stage_opamp_dummy_magic_25_0.Y.n125 two_stage_opamp_dummy_magic_25_0.Y.n90 1.5005
R24061 two_stage_opamp_dummy_magic_25_0.Y.n124 two_stage_opamp_dummy_magic_25_0.Y.n123 1.5005
R24062 two_stage_opamp_dummy_magic_25_0.Y.n122 two_stage_opamp_dummy_magic_25_0.Y.n91 1.5005
R24063 two_stage_opamp_dummy_magic_25_0.Y.n121 two_stage_opamp_dummy_magic_25_0.Y.n120 1.5005
R24064 two_stage_opamp_dummy_magic_25_0.Y.n119 two_stage_opamp_dummy_magic_25_0.Y.n93 1.5005
R24065 two_stage_opamp_dummy_magic_25_0.Y.n150 two_stage_opamp_dummy_magic_25_0.Y.n149 1.5005
R24066 two_stage_opamp_dummy_magic_25_0.Y.n151 two_stage_opamp_dummy_magic_25_0.Y.n4 1.5005
R24067 two_stage_opamp_dummy_magic_25_0.Y.n153 two_stage_opamp_dummy_magic_25_0.Y.n152 1.5005
R24068 two_stage_opamp_dummy_magic_25_0.Y.n154 two_stage_opamp_dummy_magic_25_0.Y.n2 1.5005
R24069 two_stage_opamp_dummy_magic_25_0.Y.n156 two_stage_opamp_dummy_magic_25_0.Y.n155 1.5005
R24070 two_stage_opamp_dummy_magic_25_0.Y.n3 two_stage_opamp_dummy_magic_25_0.Y.n0 1.5005
R24071 two_stage_opamp_dummy_magic_25_0.Y.n14 two_stage_opamp_dummy_magic_25_0.Y.n9 1.5005
R24072 two_stage_opamp_dummy_magic_25_0.Y.n16 two_stage_opamp_dummy_magic_25_0.Y.n15 1.5005
R24073 two_stage_opamp_dummy_magic_25_0.Y.n13 two_stage_opamp_dummy_magic_25_0.Y.n12 1.43397
R24074 two_stage_opamp_dummy_magic_25_0.Y.n18 two_stage_opamp_dummy_magic_25_0.Y.n17 1.3755
R24075 two_stage_opamp_dummy_magic_25_0.Y.n31 two_stage_opamp_dummy_magic_25_0.Y.n9 1.3755
R24076 two_stage_opamp_dummy_magic_25_0.Y.n156 two_stage_opamp_dummy_magic_25_0.Y.n1 1.3755
R24077 two_stage_opamp_dummy_magic_25_0.Y.n152 two_stage_opamp_dummy_magic_25_0.Y.n5 1.3755
R24078 two_stage_opamp_dummy_magic_25_0.Y.n150 two_stage_opamp_dummy_magic_25_0.Y.n35 1.3755
R24079 two_stage_opamp_dummy_magic_25_0.Y.n144 two_stage_opamp_dummy_magic_25_0.Y.n143 0.979667
R24080 two_stage_opamp_dummy_magic_25_0.Y.n116 two_stage_opamp_dummy_magic_25_0.Y.n96 0.792167
R24081 two_stage_opamp_dummy_magic_25_0.Y.n101 two_stage_opamp_dummy_magic_25_0.Y.n92 0.792167
R24082 two_stage_opamp_dummy_magic_25_0.Y.n104 two_stage_opamp_dummy_magic_25_0.Y.n89 0.792167
R24083 two_stage_opamp_dummy_magic_25_0.Y.n111 two_stage_opamp_dummy_magic_25_0.Y.n110 0.792167
R24084 two_stage_opamp_dummy_magic_25_0.Y.n98 two_stage_opamp_dummy_magic_25_0.Y.n94 0.792167
R24085 two_stage_opamp_dummy_magic_25_0.Y.n107 two_stage_opamp_dummy_magic_25_0.Y.n86 0.792167
R24086 two_stage_opamp_dummy_magic_25_0.Y.n83 two_stage_opamp_dummy_magic_25_0.Y.n66 0.682792
R24087 two_stage_opamp_dummy_magic_25_0.Y.n149 two_stage_opamp_dummy_magic_25_0.Y.n148 0.630708
R24088 two_stage_opamp_dummy_magic_25_0.Y.n113 two_stage_opamp_dummy_magic_25_0.Y.n112 0.6255
R24089 two_stage_opamp_dummy_magic_25_0.Y.n114 two_stage_opamp_dummy_magic_25_0.Y.n113 0.6255
R24090 two_stage_opamp_dummy_magic_25_0.Y.n115 two_stage_opamp_dummy_magic_25_0.Y.n114 0.6255
R24091 two_stage_opamp_dummy_magic_25_0.Y.n102 two_stage_opamp_dummy_magic_25_0.Y.n99 0.6255
R24092 two_stage_opamp_dummy_magic_25_0.Y.n105 two_stage_opamp_dummy_magic_25_0.Y.n102 0.6255
R24093 two_stage_opamp_dummy_magic_25_0.Y.n108 two_stage_opamp_dummy_magic_25_0.Y.n105 0.6255
R24094 two_stage_opamp_dummy_magic_25_0.Y.n137 two_stage_opamp_dummy_magic_25_0.Y.n136 0.609875
R24095 two_stage_opamp_dummy_magic_25_0.Y.n15 two_stage_opamp_dummy_magic_25_0.Y.n13 0.564601
R24096 two_stage_opamp_dummy_magic_25_0.Y.n34 two_stage_opamp_dummy_magic_25_0.Y.n33 0.563
R24097 two_stage_opamp_dummy_magic_25_0.Y.n33 two_stage_opamp_dummy_magic_25_0.Y.n32 0.563
R24098 two_stage_opamp_dummy_magic_25_0.Y.n32 two_stage_opamp_dummy_magic_25_0.Y.n8 0.563
R24099 two_stage_opamp_dummy_magic_25_0.Y.n28 two_stage_opamp_dummy_magic_25_0.Y.n21 0.563
R24100 two_stage_opamp_dummy_magic_25_0.Y.n28 two_stage_opamp_dummy_magic_25_0.Y.n27 0.563
R24101 two_stage_opamp_dummy_magic_25_0.Y.n27 two_stage_opamp_dummy_magic_25_0.Y.n24 0.563
R24102 two_stage_opamp_dummy_magic_25_0.Y.n118 two_stage_opamp_dummy_magic_25_0.Y.n94 0.533638
R24103 two_stage_opamp_dummy_magic_25_0.Y.n117 two_stage_opamp_dummy_magic_25_0.Y.n116 0.46925
R24104 two_stage_opamp_dummy_magic_25_0.Y.n122 two_stage_opamp_dummy_magic_25_0.Y.n92 0.46925
R24105 two_stage_opamp_dummy_magic_25_0.Y.n127 two_stage_opamp_dummy_magic_25_0.Y.n89 0.46925
R24106 two_stage_opamp_dummy_magic_25_0.Y.n111 two_stage_opamp_dummy_magic_25_0.Y.n87 0.46925
R24107 two_stage_opamp_dummy_magic_25_0.Y.n135 two_stage_opamp_dummy_magic_25_0.Y.n86 0.46925
R24108 two_stage_opamp_dummy_magic_25_0.Y.n146 two_stage_opamp_dummy_magic_25_0.Y.n83 0.46925
R24109 two_stage_opamp_dummy_magic_25_0.Y.n119 two_stage_opamp_dummy_magic_25_0.Y.n118 0.427973
R24110 two_stage_opamp_dummy_magic_25_0.Y.n20 two_stage_opamp_dummy_magic_25_0.Y.n18 0.3755
R24111 two_stage_opamp_dummy_magic_25_0.Y.n31 two_stage_opamp_dummy_magic_25_0.Y.n30 0.3755
R24112 two_stage_opamp_dummy_magic_25_0.Y.n26 two_stage_opamp_dummy_magic_25_0.Y.n1 0.3755
R24113 two_stage_opamp_dummy_magic_25_0.Y.n23 two_stage_opamp_dummy_magic_25_0.Y.n5 0.3755
R24114 two_stage_opamp_dummy_magic_25_0.Y.n12 two_stage_opamp_dummy_magic_25_0.Y.n11 0.3755
R24115 two_stage_opamp_dummy_magic_25_0.Y.n35 two_stage_opamp_dummy_magic_25_0.Y.n7 0.3755
R24116 two_stage_opamp_dummy_magic_25_0.Y.n82 two_stage_opamp_dummy_magic_25_0.Y.n68 0.1255
R24117 two_stage_opamp_dummy_magic_25_0.Y.n68 two_stage_opamp_dummy_magic_25_0.Y.n67 0.0626438
R24118 two_stage_opamp_dummy_magic_25_0.Y.n118 two_stage_opamp_dummy_magic_25_0.Y.n117 0.0587394
R24119 two_stage_opamp_dummy_magic_25_0.Y.n17 two_stage_opamp_dummy_magic_25_0.Y.n16 0.0577917
R24120 two_stage_opamp_dummy_magic_25_0.Y.n16 two_stage_opamp_dummy_magic_25_0.Y.n9 0.0577917
R24121 two_stage_opamp_dummy_magic_25_0.Y.n9 two_stage_opamp_dummy_magic_25_0.Y.n0 0.0577917
R24122 two_stage_opamp_dummy_magic_25_0.Y.n156 two_stage_opamp_dummy_magic_25_0.Y.n2 0.0577917
R24123 two_stage_opamp_dummy_magic_25_0.Y.n152 two_stage_opamp_dummy_magic_25_0.Y.n2 0.0577917
R24124 two_stage_opamp_dummy_magic_25_0.Y.n152 two_stage_opamp_dummy_magic_25_0.Y.n151 0.0577917
R24125 two_stage_opamp_dummy_magic_25_0.Y.n151 two_stage_opamp_dummy_magic_25_0.Y.n150 0.0577917
R24126 two_stage_opamp_dummy_magic_25_0.Y.n15 two_stage_opamp_dummy_magic_25_0.Y.n14 0.0577917
R24127 two_stage_opamp_dummy_magic_25_0.Y.n14 two_stage_opamp_dummy_magic_25_0.Y.n3 0.0577917
R24128 two_stage_opamp_dummy_magic_25_0.Y.n155 two_stage_opamp_dummy_magic_25_0.Y.n3 0.0577917
R24129 two_stage_opamp_dummy_magic_25_0.Y.n155 two_stage_opamp_dummy_magic_25_0.Y.n154 0.0577917
R24130 two_stage_opamp_dummy_magic_25_0.Y.n154 two_stage_opamp_dummy_magic_25_0.Y.n153 0.0577917
R24131 two_stage_opamp_dummy_magic_25_0.Y.n153 two_stage_opamp_dummy_magic_25_0.Y.n4 0.0577917
R24132 two_stage_opamp_dummy_magic_25_0.Y.n149 two_stage_opamp_dummy_magic_25_0.Y.n4 0.0577917
R24133 two_stage_opamp_dummy_magic_25_0.Y.n17 two_stage_opamp_dummy_magic_25_0.Y.n13 0.054517
R24134 two_stage_opamp_dummy_magic_25_0.Y.n117 two_stage_opamp_dummy_magic_25_0.Y.n93 0.0421667
R24135 two_stage_opamp_dummy_magic_25_0.Y.n121 two_stage_opamp_dummy_magic_25_0.Y.n93 0.0421667
R24136 two_stage_opamp_dummy_magic_25_0.Y.n122 two_stage_opamp_dummy_magic_25_0.Y.n121 0.0421667
R24137 two_stage_opamp_dummy_magic_25_0.Y.n123 two_stage_opamp_dummy_magic_25_0.Y.n122 0.0421667
R24138 two_stage_opamp_dummy_magic_25_0.Y.n123 two_stage_opamp_dummy_magic_25_0.Y.n90 0.0421667
R24139 two_stage_opamp_dummy_magic_25_0.Y.n127 two_stage_opamp_dummy_magic_25_0.Y.n90 0.0421667
R24140 two_stage_opamp_dummy_magic_25_0.Y.n128 two_stage_opamp_dummy_magic_25_0.Y.n127 0.0421667
R24141 two_stage_opamp_dummy_magic_25_0.Y.n129 two_stage_opamp_dummy_magic_25_0.Y.n128 0.0421667
R24142 two_stage_opamp_dummy_magic_25_0.Y.n129 two_stage_opamp_dummy_magic_25_0.Y.n87 0.0421667
R24143 two_stage_opamp_dummy_magic_25_0.Y.n133 two_stage_opamp_dummy_magic_25_0.Y.n87 0.0421667
R24144 two_stage_opamp_dummy_magic_25_0.Y.n134 two_stage_opamp_dummy_magic_25_0.Y.n133 0.0421667
R24145 two_stage_opamp_dummy_magic_25_0.Y.n135 two_stage_opamp_dummy_magic_25_0.Y.n134 0.0421667
R24146 two_stage_opamp_dummy_magic_25_0.Y.n120 two_stage_opamp_dummy_magic_25_0.Y.n119 0.0421667
R24147 two_stage_opamp_dummy_magic_25_0.Y.n120 two_stage_opamp_dummy_magic_25_0.Y.n91 0.0421667
R24148 two_stage_opamp_dummy_magic_25_0.Y.n124 two_stage_opamp_dummy_magic_25_0.Y.n91 0.0421667
R24149 two_stage_opamp_dummy_magic_25_0.Y.n125 two_stage_opamp_dummy_magic_25_0.Y.n124 0.0421667
R24150 two_stage_opamp_dummy_magic_25_0.Y.n126 two_stage_opamp_dummy_magic_25_0.Y.n125 0.0421667
R24151 two_stage_opamp_dummy_magic_25_0.Y.n126 two_stage_opamp_dummy_magic_25_0.Y.n88 0.0421667
R24152 two_stage_opamp_dummy_magic_25_0.Y.n130 two_stage_opamp_dummy_magic_25_0.Y.n88 0.0421667
R24153 two_stage_opamp_dummy_magic_25_0.Y.n131 two_stage_opamp_dummy_magic_25_0.Y.n130 0.0421667
R24154 two_stage_opamp_dummy_magic_25_0.Y.n132 two_stage_opamp_dummy_magic_25_0.Y.n131 0.0421667
R24155 two_stage_opamp_dummy_magic_25_0.Y.n132 two_stage_opamp_dummy_magic_25_0.Y.n85 0.0421667
R24156 two_stage_opamp_dummy_magic_25_0.Y.n136 two_stage_opamp_dummy_magic_25_0.Y.n85 0.0421667
R24157 two_stage_opamp_dummy_magic_25_0.Y.n146 two_stage_opamp_dummy_magic_25_0.Y.n58 0.0421667
R24158 two_stage_opamp_dummy_magic_25_0.Y two_stage_opamp_dummy_magic_25_0.Y.n0 0.0369583
R24159 two_stage_opamp_dummy_magic_25_0.Y.n142 two_stage_opamp_dummy_magic_25_0.Y.n141 0.0217373
R24160 two_stage_opamp_dummy_magic_25_0.Y.n145 two_stage_opamp_dummy_magic_25_0.Y.n144 0.0217373
R24161 two_stage_opamp_dummy_magic_25_0.Y.n147 two_stage_opamp_dummy_magic_25_0.Y.n38 0.0217373
R24162 two_stage_opamp_dummy_magic_25_0.Y.n140 two_stage_opamp_dummy_magic_25_0.Y.n84 0.0217373
R24163 two_stage_opamp_dummy_magic_25_0.Y.n143 two_stage_opamp_dummy_magic_25_0.Y.n142 0.0217373
R24164 two_stage_opamp_dummy_magic_25_0.Y.n145 two_stage_opamp_dummy_magic_25_0.Y.n36 0.0217373
R24165 two_stage_opamp_dummy_magic_25_0.Y.n38 two_stage_opamp_dummy_magic_25_0.Y.n36 0.0217373
R24166 two_stage_opamp_dummy_magic_25_0.Y.n61 two_stage_opamp_dummy_magic_25_0.Y.n59 0.0217373
R24167 two_stage_opamp_dummy_magic_25_0.Y.n62 two_stage_opamp_dummy_magic_25_0.Y.n60 0.0217373
R24168 two_stage_opamp_dummy_magic_25_0.Y.n140 two_stage_opamp_dummy_magic_25_0.Y.n139 0.0217373
R24169 two_stage_opamp_dummy_magic_25_0.Y.n141 two_stage_opamp_dummy_magic_25_0.Y.n138 0.0217373
R24170 two_stage_opamp_dummy_magic_25_0.Y.n139 two_stage_opamp_dummy_magic_25_0.Y.n137 0.0217373
R24171 two_stage_opamp_dummy_magic_25_0.Y.n148 two_stage_opamp_dummy_magic_25_0.Y.n37 0.0217373
R24172 two_stage_opamp_dummy_magic_25_0.Y.n65 two_stage_opamp_dummy_magic_25_0.Y.n60 0.0217373
R24173 two_stage_opamp_dummy_magic_25_0.Y.n58 two_stage_opamp_dummy_magic_25_0.Y.n37 0.0217373
R24174 two_stage_opamp_dummy_magic_25_0.Y.n63 two_stage_opamp_dummy_magic_25_0.Y.n61 0.0217373
R24175 two_stage_opamp_dummy_magic_25_0.Y.n64 two_stage_opamp_dummy_magic_25_0.Y.n63 0.0217373
R24176 two_stage_opamp_dummy_magic_25_0.Y.n66 two_stage_opamp_dummy_magic_25_0.Y.n65 0.0217373
R24177 two_stage_opamp_dummy_magic_25_0.Y two_stage_opamp_dummy_magic_25_0.Y.n156 0.0213333
R24178 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 344.178
R24179 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 339.272
R24180 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 339.272
R24181 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 339.272
R24182 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 334.772
R24183 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 334.772
R24184 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t20 310.682
R24185 bgr_11_0.V_TOP bgr_11_0.V_TOP.t41 310.541
R24186 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.t16 310.401
R24187 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.t29 310.401
R24188 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.t34 310.401
R24189 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t45 310.401
R24190 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t43 310.401
R24191 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t19 310.401
R24192 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t31 310.401
R24193 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t46 310.401
R24194 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t22 310.401
R24195 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t32 310.401
R24196 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t42 310.401
R24197 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t21 310.401
R24198 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t37 305.901
R24199 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t47 305.901
R24200 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.t1 108.424
R24201 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t7 99.005
R24202 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t0 39.4005
R24203 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t10 39.4005
R24204 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t2 39.4005
R24205 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t12 39.4005
R24206 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t4 39.4005
R24207 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t5 39.4005
R24208 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t9 39.4005
R24209 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t6 39.4005
R24210 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t3 39.4005
R24211 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t8 39.4005
R24212 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t11 39.4005
R24213 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t13 39.4005
R24214 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 29.0745
R24215 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 16.0376
R24216 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 4.90675
R24217 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t38 4.8295
R24218 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t27 4.8295
R24219 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t30 4.8295
R24220 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t15 4.8295
R24221 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t18 4.8295
R24222 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t40 4.8295
R24223 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t28 4.8295
R24224 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t49 4.8295
R24225 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t39 4.8295
R24226 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t44 4.5005
R24227 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t36 4.5005
R24228 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t35 4.5005
R24229 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t26 4.5005
R24230 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t25 4.5005
R24231 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t14 4.5005
R24232 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t33 4.5005
R24233 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t24 4.5005
R24234 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t17 4.5005
R24235 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t23 4.5005
R24236 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t48 4.5005
R24237 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 4.5005
R24238 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n0 4.5005
R24239 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 4.5005
R24240 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R24241 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 1.563
R24242 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 1.188
R24243 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 1.1255
R24244 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 1.1255
R24245 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n29 1.1255
R24246 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R24247 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R24248 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R24249 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R24250 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.n17 0.3295
R24251 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 0.3295
R24252 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R24253 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R24254 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n13 0.2825
R24255 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.2825
R24256 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 0.28175
R24257 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 0.28175
R24258 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 0.28175
R24259 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 0.28175
R24260 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n5 0.28175
R24261 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 0.28175
R24262 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 0.28175
R24263 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 0.28175
R24264 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 0.28175
R24265 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.n39 0.28175
R24266 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.n40 0.28175
R24267 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.n41 0.28175
R24268 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n0 0.141125
R24269 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n0 0.141125
R24270 bgr_11_0.V_TOP bgr_11_0.V_TOP.n42 0.141125
R24271 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n7 0.141125
R24272 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 0.141125
R24273 a_6470_28110.t0 a_6470_28110.t1 178.133
R24274 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n0 345.264
R24275 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n1 344.7
R24276 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n3 292.5
R24277 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t11 121.931
R24278 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n7 118.861
R24279 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n9 118.861
R24280 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n13 118.861
R24281 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n16 118.861
R24282 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n19 118.861
R24283 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n22 75.438
R24284 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n2 52.763
R24285 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n4 51.8547
R24286 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t13 39.4005
R24287 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t15 39.4005
R24288 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t16 39.4005
R24289 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t0 39.4005
R24290 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t14 39.4005
R24291 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t12 39.4005
R24292 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t3 19.7005
R24293 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t6 19.7005
R24294 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t10 19.7005
R24295 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t5 19.7005
R24296 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t9 19.7005
R24297 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t4 19.7005
R24298 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t2 19.7005
R24299 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t8 19.7005
R24300 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t1 19.7005
R24301 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t7 19.7005
R24302 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n21 5.90675
R24303 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n8 5.60467
R24304 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n18 5.54217
R24305 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n6 5.54217
R24306 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n10 5.04217
R24307 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n12 5.04217
R24308 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n5 5.04217
R24309 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n20 5.04217
R24310 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n6 4.97967
R24311 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n14 4.97967
R24312 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n17 4.97967
R24313 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n15 0.563
R24314 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n6 0.563
R24315 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n11 0.563
R24316 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n5 0.563
R24317 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n5 0.563
R24318 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t18 369.534
R24319 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t20 369.534
R24320 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t22 369.534
R24321 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t19 369.534
R24322 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t12 369.534
R24323 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t10 369.534
R24324 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t0 369.534
R24325 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n1 359.836
R24326 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t6 249.034
R24327 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t17 192.8
R24328 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t5 192.8
R24329 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t11 192.8
R24330 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t8 192.8
R24331 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t14 192.8
R24332 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t7 192.8
R24333 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t9 192.8
R24334 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t16 192.8
R24335 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t15 192.8
R24336 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t21 192.8
R24337 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t13 192.8
R24338 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R24339 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R24340 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.n11 176.733
R24341 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 176.733
R24342 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n6 167.843
R24343 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n9 166.343
R24344 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 166.343
R24345 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n18 166.343
R24346 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n0 141.752
R24347 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 56.2338
R24348 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n2 56.2338
R24349 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 56.2338
R24350 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R24351 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n14 56.2338
R24352 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n13 56.2338
R24353 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.n17 56.2338
R24354 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t4 39.4005
R24355 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t3 39.4005
R24356 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t2 24.0005
R24357 bgr_11_0.NFET_GATE_10uA.t1 bgr_11_0.NFET_GATE_10uA.n19 24.0005
R24358 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n16 2.01612
R24359 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n10 1.5005
R24360 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t13 119.785
R24361 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n0 107.121
R24362 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n1 97.4332
R24363 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n20 69.8443
R24364 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n2 38.8443
R24365 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n5 24.288
R24366 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n7 24.288
R24367 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n11 24.288
R24368 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n14 24.288
R24369 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n17 24.288
R24370 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t14 24.0005
R24371 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t0 24.0005
R24372 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t2 24.0005
R24373 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t1 24.0005
R24374 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t6 8.0005
R24375 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t9 8.0005
R24376 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t3 8.0005
R24377 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t8 8.0005
R24378 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t12 8.0005
R24379 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t7 8.0005
R24380 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t5 8.0005
R24381 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t11 8.0005
R24382 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t4 8.0005
R24383 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t10 8.0005
R24384 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n16 5.7505
R24385 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n4 5.7505
R24386 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n6 5.7505
R24387 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n19 5.6255
R24388 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n8 5.188
R24389 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n4 5.188
R24390 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n10 5.188
R24391 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n12 5.188
R24392 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n3 5.188
R24393 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n15 5.188
R24394 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n18 5.188
R24395 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n13 0.563
R24396 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n4 0.563
R24397 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n9 0.563
R24398 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n3 0.563
R24399 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n3 0.563
R24400 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t21 758.64
R24401 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n0 510.991
R24402 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n25 509.226
R24403 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t25 369.534
R24404 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t24 369.534
R24405 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t17 369.534
R24406 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t22 369.534
R24407 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t20 369.534
R24408 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t19 369.534
R24409 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n11 339.272
R24410 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 339.272
R24411 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n7 339.272
R24412 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.n5 339.272
R24413 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t15 249.034
R24414 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t23 249.034
R24415 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t16 192.8
R24416 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t10 192.8
R24417 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t26 192.8
R24418 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t11 192.8
R24419 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t18 192.8
R24420 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t28 192.8
R24421 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t14 192.8
R24422 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t13 192.8
R24423 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t12 192.8
R24424 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t27 192.8
R24425 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R24426 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R24427 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.n22 176.733
R24428 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R24429 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n17 166.541
R24430 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n3 166.343
R24431 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.t9 118.65
R24432 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t6 105.516
R24433 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 56.2338
R24434 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n15 56.2338
R24435 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n2 56.2338
R24436 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R24437 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n21 56.2338
R24438 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 56.2338
R24439 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t0 39.4005
R24440 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R24441 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R24442 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t2 39.4005
R24443 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R24444 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t1 39.4005
R24445 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R24446 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t3 39.4005
R24447 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n14 10.5429
R24448 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 6.15675
R24449 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n18 2.29514
R24450 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n4 2.28175
R24451 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.n13 1.3755
R24452 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n6 1.1255
R24453 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 1.1255
R24454 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n10 1.1255
R24455 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.n15 325.473
R24456 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 325.473
R24457 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 325.473
R24458 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t14 310.488
R24459 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t18 310.488
R24460 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t13 310.488
R24461 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.t5 184.097
R24462 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t3 184.097
R24463 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t7 184.097
R24464 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 167.094
R24465 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R24466 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R24467 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 152
R24468 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 152
R24469 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 152
R24470 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t16 120.501
R24471 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t11 120.501
R24472 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t17 120.501
R24473 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t9 120.501
R24474 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t15 120.501
R24475 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t1 120.501
R24476 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t0 106.933
R24477 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 40.7027
R24478 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R24479 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R24480 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t4 39.4005
R24481 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t10 39.4005
R24482 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t8 39.4005
R24483 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t2 39.4005
R24484 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.t6 39.4005
R24485 bgr_11_0.V_mir1.t12 bgr_11_0.V_mir1.n16 39.4005
R24486 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 15.9255
R24487 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n4 15.9255
R24488 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n11 9.3005
R24489 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.n10 4.5005
R24490 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t20 354.854
R24491 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t7 346.8
R24492 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.n6 339.522
R24493 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n15 339.522
R24494 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.n10 335.022
R24495 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t32 184.097
R24496 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t25 184.097
R24497 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t8 184.097
R24498 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t17 184.097
R24499 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 166.05
R24500 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n13 166.05
R24501 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t0 106.558
R24502 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.n4 53.7134
R24503 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t3 39.4005
R24504 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t5 39.4005
R24505 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t2 39.4005
R24506 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t1 39.4005
R24507 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t4 39.4005
R24508 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t6 39.4005
R24509 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t10 4.8295
R24510 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t28 4.8295
R24511 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t30 4.8295
R24512 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t19 4.8295
R24513 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t23 4.8295
R24514 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t12 4.8295
R24515 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t29 4.8295
R24516 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t16 4.8295
R24517 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t21 4.8295
R24518 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.n11 4.5005
R24519 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t31 4.5005
R24520 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t9 4.5005
R24521 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t24 4.5005
R24522 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t27 4.5005
R24523 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t14 4.5005
R24524 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R24525 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t22 4.5005
R24526 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t26 4.5005
R24527 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t13 4.5005
R24528 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t15 4.5005
R24529 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t11 4.5005
R24530 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n14 1.3755
R24531 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.n9 1.3755
R24532 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.n5 1.188
R24533 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n2 0.8935
R24534 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n0 0.8935
R24535 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n3 0.6585
R24536 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.6585
R24537 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n12 0.6255
R24538 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n7 0.6255
R24539 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n16 0.438
R24540 two_stage_opamp_dummy_magic_25_0.V_err_gate.n2 two_stage_opamp_dummy_magic_25_0.V_err_gate.t8 479.322
R24541 two_stage_opamp_dummy_magic_25_0.V_err_gate.n2 two_stage_opamp_dummy_magic_25_0.V_err_gate.t6 479.322
R24542 two_stage_opamp_dummy_magic_25_0.V_err_gate.n6 two_stage_opamp_dummy_magic_25_0.V_err_gate.t7 479.322
R24543 two_stage_opamp_dummy_magic_25_0.V_err_gate.n6 two_stage_opamp_dummy_magic_25_0.V_err_gate.t9 479.322
R24544 two_stage_opamp_dummy_magic_25_0.V_err_gate.n3 two_stage_opamp_dummy_magic_25_0.V_err_gate.n1 178.625
R24545 two_stage_opamp_dummy_magic_25_0.V_err_gate.n5 two_stage_opamp_dummy_magic_25_0.V_err_gate.n4 177.987
R24546 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.V_err_gate.n0 169.452
R24547 two_stage_opamp_dummy_magic_25_0.V_err_gate.n3 two_stage_opamp_dummy_magic_25_0.V_err_gate.n2 165.8
R24548 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.V_err_gate.n6 165.8
R24549 two_stage_opamp_dummy_magic_25_0.V_err_gate.n0 two_stage_opamp_dummy_magic_25_0.V_err_gate.t0 24.0005
R24550 two_stage_opamp_dummy_magic_25_0.V_err_gate.n0 two_stage_opamp_dummy_magic_25_0.V_err_gate.t1 24.0005
R24551 two_stage_opamp_dummy_magic_25_0.V_err_gate.n4 two_stage_opamp_dummy_magic_25_0.V_err_gate.t3 15.7605
R24552 two_stage_opamp_dummy_magic_25_0.V_err_gate.n4 two_stage_opamp_dummy_magic_25_0.V_err_gate.t5 15.7605
R24553 two_stage_opamp_dummy_magic_25_0.V_err_gate.n1 two_stage_opamp_dummy_magic_25_0.V_err_gate.t2 15.7605
R24554 two_stage_opamp_dummy_magic_25_0.V_err_gate.n1 two_stage_opamp_dummy_magic_25_0.V_err_gate.t4 15.7605
R24555 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.V_err_gate.n5 1.76612
R24556 two_stage_opamp_dummy_magic_25_0.V_err_gate.n5 two_stage_opamp_dummy_magic_25_0.V_err_gate.n3 0.641125
R24557 two_stage_opamp_dummy_magic_25_0.V_tot.n2 two_stage_opamp_dummy_magic_25_0.V_tot.t5 648.343
R24558 two_stage_opamp_dummy_magic_25_0.V_tot.n1 two_stage_opamp_dummy_magic_25_0.V_tot.t4 648.343
R24559 two_stage_opamp_dummy_magic_25_0.V_tot.n3 two_stage_opamp_dummy_magic_25_0.V_tot.t1 117.591
R24560 two_stage_opamp_dummy_magic_25_0.V_tot.n0 two_stage_opamp_dummy_magic_25_0.V_tot.t3 117.591
R24561 two_stage_opamp_dummy_magic_25_0.V_tot.n0 two_stage_opamp_dummy_magic_25_0.V_tot.t2 108.424
R24562 two_stage_opamp_dummy_magic_25_0.V_tot.t0 two_stage_opamp_dummy_magic_25_0.V_tot.n3 108.424
R24563 two_stage_opamp_dummy_magic_25_0.V_tot.n1 two_stage_opamp_dummy_magic_25_0.V_tot.n0 43.0496
R24564 two_stage_opamp_dummy_magic_25_0.V_tot.n3 two_stage_opamp_dummy_magic_25_0.V_tot.n2 43.0496
R24565 two_stage_opamp_dummy_magic_25_0.V_tot.n2 two_stage_opamp_dummy_magic_25_0.V_tot.n1 1.563
R24566 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t5 573.044
R24567 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t3 433.8
R24568 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n0 184.643
R24569 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n1 163.978
R24570 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n2 33.0088
R24571 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t0 15.7605
R24572 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t2 15.7605
R24573 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t4 9.6005
R24574 two_stage_opamp_dummy_magic_25_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_25_0.err_amp_mir.n3 9.6005
R24575 two_stage_opamp_dummy_magic_25_0.V_err_p.n1 two_stage_opamp_dummy_magic_25_0.V_err_p.n0 365.07
R24576 two_stage_opamp_dummy_magic_25_0.V_err_p.n0 two_stage_opamp_dummy_magic_25_0.V_err_p.t3 15.7605
R24577 two_stage_opamp_dummy_magic_25_0.V_err_p.n0 two_stage_opamp_dummy_magic_25_0.V_err_p.t0 15.7605
R24578 two_stage_opamp_dummy_magic_25_0.V_err_p.t1 two_stage_opamp_dummy_magic_25_0.V_err_p.n1 15.7605
R24579 two_stage_opamp_dummy_magic_25_0.V_err_p.n1 two_stage_opamp_dummy_magic_25_0.V_err_p.t2 15.7605
R24580 two_stage_opamp_dummy_magic_25_0.VD1.n15 two_stage_opamp_dummy_magic_25_0.VD1.n14 49.3505
R24581 two_stage_opamp_dummy_magic_25_0.VD1.n7 two_stage_opamp_dummy_magic_25_0.VD1.n6 49.3505
R24582 two_stage_opamp_dummy_magic_25_0.VD1.n39 two_stage_opamp_dummy_magic_25_0.VD1.n38 49.3505
R24583 two_stage_opamp_dummy_magic_25_0.VD1.n43 two_stage_opamp_dummy_magic_25_0.VD1.n42 49.3505
R24584 two_stage_opamp_dummy_magic_25_0.VD1.n4 two_stage_opamp_dummy_magic_25_0.VD1.n3 49.3505
R24585 two_stage_opamp_dummy_magic_25_0.VD1.n25 two_stage_opamp_dummy_magic_25_0.VD1.n24 49.3505
R24586 two_stage_opamp_dummy_magic_25_0.VD1.n9 two_stage_opamp_dummy_magic_25_0.VD1.n8 49.3505
R24587 two_stage_opamp_dummy_magic_25_0.VD1.n32 two_stage_opamp_dummy_magic_25_0.VD1.n31 49.3505
R24588 two_stage_opamp_dummy_magic_25_0.VD1.n28 two_stage_opamp_dummy_magic_25_0.VD1.n27 49.3505
R24589 two_stage_opamp_dummy_magic_25_0.VD1.n18 two_stage_opamp_dummy_magic_25_0.VD1.n17 49.3505
R24590 two_stage_opamp_dummy_magic_25_0.VD1.n12 two_stage_opamp_dummy_magic_25_0.VD1.n11 49.3505
R24591 two_stage_opamp_dummy_magic_25_0.VD1.n14 two_stage_opamp_dummy_magic_25_0.VD1.t15 16.0005
R24592 two_stage_opamp_dummy_magic_25_0.VD1.n14 two_stage_opamp_dummy_magic_25_0.VD1.t19 16.0005
R24593 two_stage_opamp_dummy_magic_25_0.VD1.n6 two_stage_opamp_dummy_magic_25_0.VD1.t20 16.0005
R24594 two_stage_opamp_dummy_magic_25_0.VD1.n6 two_stage_opamp_dummy_magic_25_0.VD1.t14 16.0005
R24595 two_stage_opamp_dummy_magic_25_0.VD1.n38 two_stage_opamp_dummy_magic_25_0.VD1.t21 16.0005
R24596 two_stage_opamp_dummy_magic_25_0.VD1.n38 two_stage_opamp_dummy_magic_25_0.VD1.t13 16.0005
R24597 two_stage_opamp_dummy_magic_25_0.VD1.n42 two_stage_opamp_dummy_magic_25_0.VD1.t18 16.0005
R24598 two_stage_opamp_dummy_magic_25_0.VD1.n42 two_stage_opamp_dummy_magic_25_0.VD1.t12 16.0005
R24599 two_stage_opamp_dummy_magic_25_0.VD1.n3 two_stage_opamp_dummy_magic_25_0.VD1.t10 16.0005
R24600 two_stage_opamp_dummy_magic_25_0.VD1.n3 two_stage_opamp_dummy_magic_25_0.VD1.t17 16.0005
R24601 two_stage_opamp_dummy_magic_25_0.VD1.n24 two_stage_opamp_dummy_magic_25_0.VD1.t3 16.0005
R24602 two_stage_opamp_dummy_magic_25_0.VD1.n24 two_stage_opamp_dummy_magic_25_0.VD1.t7 16.0005
R24603 two_stage_opamp_dummy_magic_25_0.VD1.n8 two_stage_opamp_dummy_magic_25_0.VD1.t0 16.0005
R24604 two_stage_opamp_dummy_magic_25_0.VD1.n8 two_stage_opamp_dummy_magic_25_0.VD1.t5 16.0005
R24605 two_stage_opamp_dummy_magic_25_0.VD1.n31 two_stage_opamp_dummy_magic_25_0.VD1.t2 16.0005
R24606 two_stage_opamp_dummy_magic_25_0.VD1.n31 two_stage_opamp_dummy_magic_25_0.VD1.t6 16.0005
R24607 two_stage_opamp_dummy_magic_25_0.VD1.n27 two_stage_opamp_dummy_magic_25_0.VD1.t1 16.0005
R24608 two_stage_opamp_dummy_magic_25_0.VD1.n27 two_stage_opamp_dummy_magic_25_0.VD1.t8 16.0005
R24609 two_stage_opamp_dummy_magic_25_0.VD1.n17 two_stage_opamp_dummy_magic_25_0.VD1.t11 16.0005
R24610 two_stage_opamp_dummy_magic_25_0.VD1.n17 two_stage_opamp_dummy_magic_25_0.VD1.t16 16.0005
R24611 two_stage_opamp_dummy_magic_25_0.VD1.n11 two_stage_opamp_dummy_magic_25_0.VD1.t4 16.0005
R24612 two_stage_opamp_dummy_magic_25_0.VD1.n11 two_stage_opamp_dummy_magic_25_0.VD1.t9 16.0005
R24613 two_stage_opamp_dummy_magic_25_0.VD1.n33 two_stage_opamp_dummy_magic_25_0.VD1.n2 6.2505
R24614 two_stage_opamp_dummy_magic_25_0.VD1.n36 two_stage_opamp_dummy_magic_25_0.VD1.n35 6.2505
R24615 two_stage_opamp_dummy_magic_25_0.VD1.n23 two_stage_opamp_dummy_magic_25_0.VD1.n13 6.2505
R24616 two_stage_opamp_dummy_magic_25_0.VD1.n21 two_stage_opamp_dummy_magic_25_0.VD1.n20 6.2505
R24617 two_stage_opamp_dummy_magic_25_0.VD1.n30 two_stage_opamp_dummy_magic_25_0.VD1.n9 5.6255
R24618 two_stage_opamp_dummy_magic_25_0.VD1.n26 two_stage_opamp_dummy_magic_25_0.VD1.n12 5.6255
R24619 two_stage_opamp_dummy_magic_25_0.VD1.n40 two_stage_opamp_dummy_magic_25_0.VD1.n7 5.438
R24620 two_stage_opamp_dummy_magic_25_0.VD1.n16 two_stage_opamp_dummy_magic_25_0.VD1.n15 5.438
R24621 two_stage_opamp_dummy_magic_25_0.VD1.n36 two_stage_opamp_dummy_magic_25_0.VD1.n7 5.31821
R24622 two_stage_opamp_dummy_magic_25_0.VD1.n20 two_stage_opamp_dummy_magic_25_0.VD1.n15 5.31821
R24623 two_stage_opamp_dummy_magic_25_0.VD1.n39 two_stage_opamp_dummy_magic_25_0.VD1.n37 5.08383
R24624 two_stage_opamp_dummy_magic_25_0.VD1.n44 two_stage_opamp_dummy_magic_25_0.VD1.n43 5.08383
R24625 two_stage_opamp_dummy_magic_25_0.VD1.n4 two_stage_opamp_dummy_magic_25_0.VD1.n1 5.08383
R24626 two_stage_opamp_dummy_magic_25_0.VD1.n19 two_stage_opamp_dummy_magic_25_0.VD1.n18 5.08383
R24627 two_stage_opamp_dummy_magic_25_0.VD1.n32 two_stage_opamp_dummy_magic_25_0.VD1.n30 5.063
R24628 two_stage_opamp_dummy_magic_25_0.VD1.n29 two_stage_opamp_dummy_magic_25_0.VD1.n28 5.063
R24629 two_stage_opamp_dummy_magic_25_0.VD1.n22 two_stage_opamp_dummy_magic_25_0.VD1.n21 5.063
R24630 two_stage_opamp_dummy_magic_25_0.VD1.n35 two_stage_opamp_dummy_magic_25_0.VD1.n34 5.063
R24631 two_stage_opamp_dummy_magic_25_0.VD1.n26 two_stage_opamp_dummy_magic_25_0.VD1.n25 5.063
R24632 two_stage_opamp_dummy_magic_25_0.VD1.n40 two_stage_opamp_dummy_magic_25_0.VD1.n39 4.8755
R24633 two_stage_opamp_dummy_magic_25_0.VD1.n43 two_stage_opamp_dummy_magic_25_0.VD1.n41 4.8755
R24634 two_stage_opamp_dummy_magic_25_0.VD1.n5 two_stage_opamp_dummy_magic_25_0.VD1.n4 4.8755
R24635 two_stage_opamp_dummy_magic_25_0.VD1.n18 two_stage_opamp_dummy_magic_25_0.VD1.n16 4.8755
R24636 two_stage_opamp_dummy_magic_25_0.VD1 two_stage_opamp_dummy_magic_25_0.VD1.n45 4.60467
R24637 two_stage_opamp_dummy_magic_25_0.VD1.n10 two_stage_opamp_dummy_magic_25_0.VD1.n0 4.5005
R24638 two_stage_opamp_dummy_magic_25_0.VD1.n34 two_stage_opamp_dummy_magic_25_0.VD1.n33 4.5005
R24639 two_stage_opamp_dummy_magic_25_0.VD1.n23 two_stage_opamp_dummy_magic_25_0.VD1.n22 4.5005
R24640 two_stage_opamp_dummy_magic_25_0.VD1 two_stage_opamp_dummy_magic_25_0.VD1.n0 1.64633
R24641 two_stage_opamp_dummy_magic_25_0.VD1.n22 two_stage_opamp_dummy_magic_25_0.VD1.n10 0.563
R24642 two_stage_opamp_dummy_magic_25_0.VD1.n34 two_stage_opamp_dummy_magic_25_0.VD1.n10 0.563
R24643 two_stage_opamp_dummy_magic_25_0.VD1.n30 two_stage_opamp_dummy_magic_25_0.VD1.n29 0.563
R24644 two_stage_opamp_dummy_magic_25_0.VD1.n29 two_stage_opamp_dummy_magic_25_0.VD1.n26 0.563
R24645 two_stage_opamp_dummy_magic_25_0.VD1.n41 two_stage_opamp_dummy_magic_25_0.VD1.n40 0.563
R24646 two_stage_opamp_dummy_magic_25_0.VD1.n41 two_stage_opamp_dummy_magic_25_0.VD1.n5 0.563
R24647 two_stage_opamp_dummy_magic_25_0.VD1.n16 two_stage_opamp_dummy_magic_25_0.VD1.n5 0.563
R24648 two_stage_opamp_dummy_magic_25_0.VD1.n33 two_stage_opamp_dummy_magic_25_0.VD1.n32 0.3755
R24649 two_stage_opamp_dummy_magic_25_0.VD1.n28 two_stage_opamp_dummy_magic_25_0.VD1.n0 0.3755
R24650 two_stage_opamp_dummy_magic_25_0.VD1.n35 two_stage_opamp_dummy_magic_25_0.VD1.n9 0.3755
R24651 two_stage_opamp_dummy_magic_25_0.VD1.n25 two_stage_opamp_dummy_magic_25_0.VD1.n23 0.3755
R24652 two_stage_opamp_dummy_magic_25_0.VD1.n21 two_stage_opamp_dummy_magic_25_0.VD1.n12 0.3755
R24653 two_stage_opamp_dummy_magic_25_0.VD1.n20 two_stage_opamp_dummy_magic_25_0.VD1.n19 0.234875
R24654 two_stage_opamp_dummy_magic_25_0.VD1.n19 two_stage_opamp_dummy_magic_25_0.VD1.n13 0.234875
R24655 two_stage_opamp_dummy_magic_25_0.VD1.n13 two_stage_opamp_dummy_magic_25_0.VD1.n1 0.234875
R24656 two_stage_opamp_dummy_magic_25_0.VD1.n45 two_stage_opamp_dummy_magic_25_0.VD1.n1 0.234875
R24657 two_stage_opamp_dummy_magic_25_0.VD1.n45 two_stage_opamp_dummy_magic_25_0.VD1.n44 0.234875
R24658 two_stage_opamp_dummy_magic_25_0.VD1.n44 two_stage_opamp_dummy_magic_25_0.VD1.n2 0.234875
R24659 two_stage_opamp_dummy_magic_25_0.VD1.n37 two_stage_opamp_dummy_magic_25_0.VD1.n2 0.234875
R24660 two_stage_opamp_dummy_magic_25_0.VD1.n37 two_stage_opamp_dummy_magic_25_0.VD1.n36 0.234875
R24661 a_12070_29568.t0 a_12070_29568.t1 178.133
R24662 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t3 536.909
R24663 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 370.586
R24664 bgr_11_0.V_CUR_REF_REG.t0 bgr_11_0.V_CUR_REF_REG.n1 152.224
R24665 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t1 39.4005
R24666 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R24667 bgr_11_0.1st_Vout_2.n15 bgr_11_0.1st_Vout_2.t19 355.293
R24668 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t20 346.8
R24669 bgr_11_0.1st_Vout_2.n16 bgr_11_0.1st_Vout_2.n15 339.522
R24670 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n6 339.522
R24671 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.n10 335.022
R24672 bgr_11_0.1st_Vout_2.n13 bgr_11_0.1st_Vout_2.t26 184.097
R24673 bgr_11_0.1st_Vout_2.n13 bgr_11_0.1st_Vout_2.t12 184.097
R24674 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t31 184.097
R24675 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t15 184.097
R24676 bgr_11_0.1st_Vout_2.n14 bgr_11_0.1st_Vout_2.n13 166.05
R24677 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n8 166.05
R24678 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t6 106.558
R24679 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.n4 53.6509
R24680 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t4 39.4005
R24681 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t0 39.4005
R24682 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t3 39.4005
R24683 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t1 39.4005
R24684 bgr_11_0.1st_Vout_2.t5 bgr_11_0.1st_Vout_2.n16 39.4005
R24685 bgr_11_0.1st_Vout_2.n16 bgr_11_0.1st_Vout_2.t2 39.4005
R24686 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t18 4.8295
R24687 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t25 4.8295
R24688 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t10 4.8295
R24689 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t17 4.8295
R24690 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t29 4.8295
R24691 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t8 4.8295
R24692 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t9 4.8295
R24693 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t14 4.8295
R24694 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t7 4.8295
R24695 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t11 4.5005
R24696 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t32 4.5005
R24697 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t30 4.5005
R24698 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t24 4.5005
R24699 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t23 4.5005
R24700 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t16 4.5005
R24701 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t28 4.5005
R24702 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t22 4.5005
R24703 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t27 4.5005
R24704 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t21 4.5005
R24705 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.t13 4.5005
R24706 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n11 4.5005
R24707 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n9 1.3755
R24708 bgr_11_0.1st_Vout_2.n15 bgr_11_0.1st_Vout_2.n14 1.3755
R24709 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n5 1.188
R24710 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n2 0.8935
R24711 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n0 0.8935
R24712 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n3 0.6585
R24713 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n1 0.6585
R24714 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n7 0.6255
R24715 bgr_11_0.1st_Vout_2.n14 bgr_11_0.1st_Vout_2.n12 0.6255
R24716 bgr_11_0.cap_res2.t20 bgr_11_0.cap_res2.t14 121.245
R24717 bgr_11_0.cap_res2.t9 bgr_11_0.cap_res2.t4 0.1603
R24718 bgr_11_0.cap_res2.t3 bgr_11_0.cap_res2.t17 0.1603
R24719 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.t2 0.1603
R24720 bgr_11_0.cap_res2.t1 bgr_11_0.cap_res2.t16 0.1603
R24721 bgr_11_0.cap_res2.t15 bgr_11_0.cap_res2.t10 0.1603
R24722 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t0 0.159278
R24723 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t6 0.159278
R24724 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t12 0.159278
R24725 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t8 0.159278
R24726 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t19 0.1368
R24727 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t9 0.1368
R24728 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t13 0.1368
R24729 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t3 0.1368
R24730 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t18 0.1368
R24731 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t7 0.1368
R24732 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t11 0.1368
R24733 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t1 0.1368
R24734 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t5 0.1368
R24735 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t15 0.1368
R24736 bgr_11_0.cap_res2.t0 bgr_11_0.cap_res2.n0 0.00152174
R24737 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.n1 0.00152174
R24738 bgr_11_0.cap_res2.t12 bgr_11_0.cap_res2.n2 0.00152174
R24739 bgr_11_0.cap_res2.t8 bgr_11_0.cap_res2.n3 0.00152174
R24740 bgr_11_0.cap_res2.t14 bgr_11_0.cap_res2.n4 0.00152174
R24741 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n0 344.837
R24742 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n1 344.274
R24743 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n3 292.5
R24744 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t0 121.785
R24745 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n7 118.861
R24746 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n9 118.861
R24747 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n13 118.861
R24748 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n16 118.861
R24749 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n19 118.861
R24750 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n22 77.4067
R24751 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n2 52.3363
R24752 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n4 52.2813
R24753 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t16 39.4005
R24754 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t13 39.4005
R24755 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t11 39.4005
R24756 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t14 39.4005
R24757 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t12 39.4005
R24758 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t15 39.4005
R24759 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t9 19.7005
R24760 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t4 19.7005
R24761 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t10 19.7005
R24762 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t5 19.7005
R24763 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t2 19.7005
R24764 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t6 19.7005
R24765 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t1 19.7005
R24766 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t8 19.7005
R24767 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t3 19.7005
R24768 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t7 19.7005
R24769 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n21 5.90675
R24770 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n8 5.60467
R24771 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n18 5.54217
R24772 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n6 5.54217
R24773 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n10 5.04217
R24774 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n12 5.04217
R24775 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n5 5.04217
R24776 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n20 5.04217
R24777 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n6 4.97967
R24778 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n14 4.97967
R24779 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n17 4.97967
R24780 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n15 0.563
R24781 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n6 0.563
R24782 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n11 0.563
R24783 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n5 0.563
R24784 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n5 0.563
R24785 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t14 119.785
R24786 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n0 107.121
R24787 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n1 97.4332
R24788 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n20 65.8443
R24789 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n2 30.2474
R24790 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n5 24.288
R24791 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n7 24.288
R24792 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n11 24.288
R24793 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n14 24.288
R24794 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n17 24.288
R24795 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t2 24.0005
R24796 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t13 24.0005
R24797 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t0 24.0005
R24798 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t1 24.0005
R24799 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t12 8.0005
R24800 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t7 8.0005
R24801 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t3 8.0005
R24802 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t8 8.0005
R24803 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t5 8.0005
R24804 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t9 8.0005
R24805 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t4 8.0005
R24806 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t11 8.0005
R24807 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t6 8.0005
R24808 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t10 8.0005
R24809 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n16 5.7505
R24810 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n4 5.7505
R24811 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n6 5.7505
R24812 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n19 5.6255
R24813 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n8 5.188
R24814 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n4 5.188
R24815 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n10 5.188
R24816 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n12 5.188
R24817 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n3 5.188
R24818 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n15 5.188
R24819 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n18 5.188
R24820 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n13 0.563
R24821 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n4 0.563
R24822 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n9 0.563
R24823 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n3 0.563
R24824 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n3 0.563
R24825 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R24826 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R24827 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 167.332
R24828 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t5 130.001
R24829 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 111.796
R24830 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 105.171
R24831 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t4 81.7074
R24832 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.8552
R24833 bgr_11_0.START_UP bgr_11_0.START_UP.n5 14.4693
R24834 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t2 13.1338
R24835 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t0 13.1338
R24836 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t1 13.1338
R24837 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t3 13.1338
R24838 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R24839 VIN-.n0 VIN-.t7 1097.62
R24840 VIN- VIN-.n9 433.019
R24841 VIN-.n9 VIN-.t10 273.134
R24842 VIN-.n0 VIN-.t9 273.134
R24843 VIN-.n1 VIN-.t3 273.134
R24844 VIN-.n2 VIN-.t8 273.134
R24845 VIN-.n3 VIN-.t1 273.134
R24846 VIN-.n4 VIN-.t5 273.134
R24847 VIN-.n5 VIN-.t2 273.134
R24848 VIN-.n6 VIN-.t6 273.134
R24849 VIN-.n7 VIN-.t0 273.134
R24850 VIN-.n8 VIN-.t4 273.134
R24851 VIN-.n9 VIN-.n8 176.733
R24852 VIN-.n8 VIN-.n7 176.733
R24853 VIN-.n7 VIN-.n6 176.733
R24854 VIN-.n6 VIN-.n5 176.733
R24855 VIN-.n5 VIN-.n4 176.733
R24856 VIN-.n4 VIN-.n3 176.733
R24857 VIN-.n3 VIN-.n2 176.733
R24858 VIN-.n2 VIN-.n1 176.733
R24859 VIN-.n1 VIN-.n0 176.733
R24860 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t14 610.534
R24861 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t24 610.534
R24862 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t22 433.8
R24863 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t27 433.8
R24864 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t16 433.8
R24865 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t25 433.8
R24866 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t12 433.8
R24867 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t20 433.8
R24868 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t30 433.8
R24869 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t18 433.8
R24870 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t15 433.8
R24871 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t17 433.8
R24872 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t26 433.8
R24873 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t13 433.8
R24874 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t21 433.8
R24875 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t31 433.8
R24876 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t19 433.8
R24877 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t29 433.8
R24878 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t23 433.8
R24879 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t28 433.8
R24880 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n27 287.264
R24881 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n23 287.264
R24882 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n24 287.264
R24883 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n30 287.264
R24884 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n10 176.733
R24885 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n9 176.733
R24886 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n8 176.733
R24887 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n7 176.733
R24888 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n6 176.733
R24889 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n5 176.733
R24890 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n4 176.733
R24891 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n3 176.733
R24892 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n13 176.733
R24893 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n14 176.733
R24894 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n15 176.733
R24895 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n16 176.733
R24896 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n17 176.733
R24897 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n18 176.733
R24898 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n20 176.733
R24899 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate.n12 161.863
R24900 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate.n22 161.863
R24901 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n31 62.6961
R24902 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n2 62.6953
R24903 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n0 62.6953
R24904 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n2 52.5725
R24905 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n29 52.5725
R24906 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n28 52.01
R24907 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n25 52.01
R24908 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate.n32 50.4989
R24909 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate.n33 50.4989
R24910 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_25_0.V_tail_gate 46.7517
R24911 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n11 45.5227
R24912 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n19 45.5227
R24913 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n21 45.5227
R24914 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n12 45.5227
R24915 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t7 39.4005
R24916 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t4 39.4005
R24917 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t3 39.4005
R24918 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t8 39.4005
R24919 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t9 39.4005
R24920 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t5 39.4005
R24921 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t10 39.4005
R24922 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t6 39.4005
R24923 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t0 16.0005
R24924 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t1 16.0005
R24925 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t2 16.0005
R24926 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t11 16.0005
R24927 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate.n1 15.9442
R24928 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate.n0 7.03346
R24929 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n26 0.563
R24930 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n1 0.340713
R24931 a_5700_29568.t0 a_5700_29568.t1 178.133
R24932 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t7 651.405
R24933 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t9 648.03
R24934 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t8 540.458
R24935 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t0 125.486
R24936 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n2 109.829
R24937 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n5 105.454
R24938 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n3 105.454
R24939 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n7 69.813
R24940 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t3 13.1338
R24941 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t1 13.1338
R24942 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t4 13.1338
R24943 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t5 13.1338
R24944 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t2 13.1338
R24945 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t6 13.1338
R24946 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n6 10.0317
R24947 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n4 4.3755
R24948 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n1 2.84425
R24949 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n0 1.53175
R24950 bgr_11_0.cap_res1.t0 bgr_11_0.cap_res1.t16 121.245
R24951 bgr_11_0.cap_res1.t14 bgr_11_0.cap_res1.t18 0.1603
R24952 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.t13 0.1603
R24953 bgr_11_0.cap_res1.t12 bgr_11_0.cap_res1.t17 0.1603
R24954 bgr_11_0.cap_res1.t5 bgr_11_0.cap_res1.t11 0.1603
R24955 bgr_11_0.cap_res1.t20 bgr_11_0.cap_res1.t4 0.1603
R24956 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t1 0.159278
R24957 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t7 0.159278
R24958 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t15 0.159278
R24959 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t9 0.159278
R24960 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t14 0.1368
R24961 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t10 0.1368
R24962 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t6 0.1368
R24963 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t3 0.1368
R24964 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t12 0.1368
R24965 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t8 0.1368
R24966 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t5 0.1368
R24967 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t2 0.1368
R24968 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t20 0.1368
R24969 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t19 0.1368
R24970 bgr_11_0.cap_res1.t1 bgr_11_0.cap_res1.n0 0.00152174
R24971 bgr_11_0.cap_res1.t7 bgr_11_0.cap_res1.n1 0.00152174
R24972 bgr_11_0.cap_res1.t15 bgr_11_0.cap_res1.n2 0.00152174
R24973 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.n3 0.00152174
R24974 bgr_11_0.cap_res1.t16 bgr_11_0.cap_res1.n4 0.00152174
R24975 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t8 525.38
R24976 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t7 525.38
R24977 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t6 525.38
R24978 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t5 525.38
R24979 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n4 491.151
R24980 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n1 491.151
R24981 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t4 281.168
R24982 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t9 281.168
R24983 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t2 281.168
R24984 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t3 281.168
R24985 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n3 244.214
R24986 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n0 244.214
R24987 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t1 118.129
R24988 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n5 118.129
R24989 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n2 23.3755
R24990 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t8 539.797
R24991 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 351.865
R24992 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n17 141.667
R24993 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.t5 117.817
R24994 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n3 109.204
R24995 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n4 104.829
R24996 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n18 84.0884
R24997 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 83.5719
R24998 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n0 83.5719
R24999 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n1 83.5719
R25000 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t0 65.0299
R25001 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t7 39.4005
R25002 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t6 39.4005
R25003 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 26.074
R25004 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n15 26.074
R25005 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n16 26.074
R25006 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 24.3755
R25007 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 17.188
R25008 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t3 13.1338
R25009 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t4 13.1338
R25010 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t1 13.1338
R25011 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t2 13.1338
R25012 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 11.0943
R25013 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n5 3.8755
R25014 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n19 1.56836
R25015 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n11 1.56363
R25016 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n20 1.5505
R25017 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n2 1.5505
R25018 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n1 1.14402
R25019 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n0 0.885803
R25020 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 0.77514
R25021 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R25022 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n1 0.701365
R25023 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n10 0.530034
R25024 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.t0 0.290206
R25025 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n21 0.203382
R25026 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n2 0.0183571
R25027 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n2 0.00817857
R25028 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 201.124
R25029 bgr_11_0.V_p_2.t0 bgr_11_0.V_p_2.n0 9.6005
R25030 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t1 9.6005
R25031 two_stage_opamp_dummy_magic_25_0.Vb2_2.n2 two_stage_opamp_dummy_magic_25_0.Vb2_2.t6 661.375
R25032 two_stage_opamp_dummy_magic_25_0.Vb2_2.n4 two_stage_opamp_dummy_magic_25_0.Vb2_2.t3 661.375
R25033 two_stage_opamp_dummy_magic_25_0.Vb2_2.t7 two_stage_opamp_dummy_magic_25_0.Vb2_2.n0 213.131
R25034 two_stage_opamp_dummy_magic_25_0.Vb2_2.n3 two_stage_opamp_dummy_magic_25_0.Vb2_2.t4 213.131
R25035 two_stage_opamp_dummy_magic_25_0.Vb2_2.n6 two_stage_opamp_dummy_magic_25_0.Vb2_2.n1 155.123
R25036 two_stage_opamp_dummy_magic_25_0.Vb2_2.t0 two_stage_opamp_dummy_magic_25_0.Vb2_2.t7 146.155
R25037 two_stage_opamp_dummy_magic_25_0.Vb2_2.t4 two_stage_opamp_dummy_magic_25_0.Vb2_2.t0 146.155
R25038 two_stage_opamp_dummy_magic_25_0.Vb2_2.t8 two_stage_opamp_dummy_magic_25_0.Vb2_2.n0 76.2576
R25039 two_stage_opamp_dummy_magic_25_0.Vb2_2.n3 two_stage_opamp_dummy_magic_25_0.Vb2_2.t5 76.2576
R25040 two_stage_opamp_dummy_magic_25_0.Vb2_2.n7 two_stage_opamp_dummy_magic_25_0.Vb2_2.n6 66.4336
R25041 two_stage_opamp_dummy_magic_25_0.Vb2_2.n1 two_stage_opamp_dummy_magic_25_0.Vb2_2.t9 21.8894
R25042 two_stage_opamp_dummy_magic_25_0.Vb2_2.n1 two_stage_opamp_dummy_magic_25_0.Vb2_2.t2 21.8894
R25043 two_stage_opamp_dummy_magic_25_0.Vb2_2.t8 two_stage_opamp_dummy_magic_25_0.Vb2_2.n7 11.2576
R25044 two_stage_opamp_dummy_magic_25_0.Vb2_2.n7 two_stage_opamp_dummy_magic_25_0.Vb2_2.t1 11.2576
R25045 two_stage_opamp_dummy_magic_25_0.Vb2_2.n5 two_stage_opamp_dummy_magic_25_0.Vb2_2.n4 5.1255
R25046 two_stage_opamp_dummy_magic_25_0.Vb2_2.n6 two_stage_opamp_dummy_magic_25_0.Vb2_2.n5 4.92976
R25047 two_stage_opamp_dummy_magic_25_0.Vb2_2.n5 two_stage_opamp_dummy_magic_25_0.Vb2_2.n2 4.7505
R25048 two_stage_opamp_dummy_magic_25_0.Vb2_2.n4 two_stage_opamp_dummy_magic_25_0.Vb2_2.n3 1.888
R25049 two_stage_opamp_dummy_magic_25_0.Vb2_2.n2 two_stage_opamp_dummy_magic_25_0.Vb2_2.n0 1.888
R25050 two_stage_opamp_dummy_magic_25_0.V_p_mir.n0 two_stage_opamp_dummy_magic_25_0.V_p_mir.t3 16.0005
R25051 two_stage_opamp_dummy_magic_25_0.V_p_mir.n0 two_stage_opamp_dummy_magic_25_0.V_p_mir.t2 16.0005
R25052 two_stage_opamp_dummy_magic_25_0.V_p_mir.n1 two_stage_opamp_dummy_magic_25_0.V_p_mir.t0 9.6005
R25053 two_stage_opamp_dummy_magic_25_0.V_p_mir.t1 two_stage_opamp_dummy_magic_25_0.V_p_mir.n1 9.6005
R25054 two_stage_opamp_dummy_magic_25_0.V_p_mir.n1 two_stage_opamp_dummy_magic_25_0.V_p_mir.n0 89.8428
R25055 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 529.879
R25056 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t0 148.653
R25057 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t1 125.418
R25058 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n1 106.609
R25059 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 104.484
R25060 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n0 24.6434
R25061 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 18.2193
R25062 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t3 13.1338
R25063 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t2 13.1338
R25064 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t5 13.1338
R25065 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t4 13.1338
R25066 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 6.53175
R25067 two_stage_opamp_dummy_magic_25_0.V_err_mir_p two_stage_opamp_dummy_magic_25_0.V_err_mir_p.n1 187.316
R25068 two_stage_opamp_dummy_magic_25_0.V_err_mir_p two_stage_opamp_dummy_magic_25_0.V_err_mir_p.n0 177.754
R25069 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t0 15.7605
R25070 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t3 15.7605
R25071 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t2 15.7605
R25072 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_25_0.V_err_mir_p.t1 15.7605
R25073 a_6350_29718.t0 a_6350_29718.t1 178.133
R25074 a_13840_3288.t0 a_13840_3288.t1 294.339
R25075 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R25076 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t3 661.375
R25077 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t0 661.375
R25078 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n6 213.131
R25079 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t4 213.131
R25080 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t1 146.155
R25081 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t7 146.155
R25082 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t2 76.2576
R25083 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n7 76.2576
R25084 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n1 72.5885
R25085 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n2 66.4444
R25086 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t8 11.2576
R25087 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t5 11.2576
R25088 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t9 11.2576
R25089 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.t10 11.2576
R25090 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n4 5.1255
R25091 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n3 4.91892
R25092 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n0 4.7505
R25093 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n5 1.888
R25094 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_25_0.Vb2_Vb3.n0 1.888
R25095 a_3690_3288.t0 a_3690_3288.t1 294.339
R25096 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 172.969
R25097 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R25098 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R25099 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R25100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R25101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R25102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R25103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R25104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R25105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R25106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R25107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R25108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R25109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R25110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R25111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R25112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R25113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R25114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R25115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R25116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R25117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R25118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R25119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R25120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R25121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R25122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R25123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R25124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R25125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R25126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R25127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R25128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R25129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R25130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R25131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R25132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R25133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R25134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 65.0299
R25135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R25136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R25137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R25138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R25139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R25140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R25141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R25142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R25143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R25144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R25145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R25146 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R25147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R25148 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R25149 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R25150 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25151 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25152 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R25153 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25154 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25155 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25156 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R25157 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25158 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25159 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25160 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25161 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R25162 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R25163 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25164 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25165 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25166 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R25167 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25168 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25169 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25170 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R25171 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25172 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25173 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25174 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R25175 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R25176 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R25177 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25178 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25179 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25180 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R25181 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25182 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25183 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25184 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R25185 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25186 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25187 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25188 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25189 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25190 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25191 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25192 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25193 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25194 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25195 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25196 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25197 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R25198 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R25199 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25200 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25201 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25202 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25203 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R25204 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R25205 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R25206 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R25207 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R25208 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R25209 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R25210 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R25211 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R25212 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R25213 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R25214 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R25215 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R25216 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R25217 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R25218 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R25219 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R25220 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R25221 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R25222 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R25223 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R25224 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R25225 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R25226 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R25227 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R25228 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R25229 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R25230 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R25231 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R25232 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R25233 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R25234 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R25235 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R25236 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R25237 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R25238 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R25239 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R25240 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R25241 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R25242 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R25243 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R25244 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R25245 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R25246 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R25247 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R25248 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R25249 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R25250 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R25251 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R25252 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R25253 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R25254 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R25255 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R25256 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R25257 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R25258 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R25259 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R25260 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R25261 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R25262 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R25263 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R25264 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R25265 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R25266 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R25267 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R25268 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R25269 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R25270 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R25271 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R25272 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R25273 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R25274 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R25275 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R25276 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R25277 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R25278 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R25279 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R25280 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R25281 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R25282 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R25283 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R25284 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R25285 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R25286 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R25287 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R25288 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R25289 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R25290 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R25291 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R25292 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R25293 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R25294 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R25295 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R25296 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R25297 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R25298 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R25299 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R25300 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R25301 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R25302 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R25303 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R25304 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R25305 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 0.290206
R25306 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R25307 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R25308 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R25309 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R25310 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R25311 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R25312 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25313 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25314 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25315 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R25316 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25317 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R25318 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R25319 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R25320 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R25321 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R25322 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R25323 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R25324 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R25325 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R25326 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R25327 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R25328 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R25329 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R25330 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R25331 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R25332 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R25333 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R25334 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R25335 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R25336 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R25337 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R25338 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R25339 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R25340 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R25341 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R25342 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R25343 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R25344 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R25345 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R25346 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R25347 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R25348 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R25349 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R25350 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R25351 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R25352 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R25353 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R25354 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R25355 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R25356 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R25357 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R25358 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R25359 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R25360 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R25361 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R25362 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R25363 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R25364 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R25365 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R25366 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R25367 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R25368 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R25369 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R25370 a_13960_3288.t0 a_13960_3288.t1 169.905
R25371 a_11420_29718.t0 a_11420_29718.t1 178.133
R25372 a_11950_28360.t0 a_11950_28360.t1 178.133
R25373 two_stage_opamp_dummy_magic_25_0.err_amp_out.n1 two_stage_opamp_dummy_magic_25_0.err_amp_out.t4 1025.2
R25374 two_stage_opamp_dummy_magic_25_0.err_amp_out.n1 two_stage_opamp_dummy_magic_25_0.err_amp_out.n0 179.382
R25375 two_stage_opamp_dummy_magic_25_0.err_amp_out.n2 two_stage_opamp_dummy_magic_25_0.err_amp_out.n1 39.3422
R25376 two_stage_opamp_dummy_magic_25_0.err_amp_out.n0 two_stage_opamp_dummy_magic_25_0.err_amp_out.t2 15.7605
R25377 two_stage_opamp_dummy_magic_25_0.err_amp_out.n0 two_stage_opamp_dummy_magic_25_0.err_amp_out.t1 15.7605
R25378 two_stage_opamp_dummy_magic_25_0.err_amp_out.t0 two_stage_opamp_dummy_magic_25_0.err_amp_out.n2 9.6005
R25379 two_stage_opamp_dummy_magic_25_0.err_amp_out.n2 two_stage_opamp_dummy_magic_25_0.err_amp_out.t3 9.6005
R25380 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t2 99.603
R25381 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t1 9.6005
R25382 bgr_11_0.V_p_1.t0 bgr_11_0.V_p_1.n0 9.6005
R25383 a_11300_28110.t0 a_11300_28110.t1 178.133
R25384 a_13940_n584.t0 a_13940_n584.t1 169.905
R25385 a_5820_28304.t0 a_5820_28304.t1 178.133
R25386 a_3830_n584.t0 a_3830_n584.t1 169.905
R25387 a_3810_3288.t0 a_3810_3288.t1 169.905
C0 two_stage_opamp_dummy_magic_25_0.V_tail_gate VOUT- 1.28602f
C1 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_25_0.V_tail_gate 0.582261f
C2 bgr_11_0.Vin+ bgr_11_0.START_UP 0.170149f
C3 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.V_err_mir_p 0.047104f
C4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.058662f
C5 bgr_11_0.START_UP_NFET1 VDDA 0.187957f
C6 VDDA VOUT- 15.3137f
C7 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_25_0.V_err_gate 0.104624f
C8 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.VD1 0.329453f
C9 bgr_11_0.PFET_GATE_10uA VDDA 9.53048f
C10 two_stage_opamp_dummy_magic_25_0.V_tail_gate VIN+ 0.059812f
C11 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.VD2 0.357127f
C12 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.cap_res_X 0.15916f
C13 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.Vb1 3.27161f
C14 two_stage_opamp_dummy_magic_25_0.Y two_stage_opamp_dummy_magic_25_0.V_err_mir_p 0.013108f
C15 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref bgr_11_0.Vin+ 0.228924f
C16 bgr_11_0.V_TOP bgr_11_0.START_UP 1.37397f
C17 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.cap_res_Y 0.218019f
C18 VOUT+ VOUT- 0.118487f
C19 two_stage_opamp_dummy_magic_25_0.V_tail_gate VIN- 0.057394f
C20 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.X 0.40038f
C21 two_stage_opamp_dummy_magic_25_0.V_err_gate bgr_11_0.START_UP 0.683079f
C22 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.Y 0.875295f
C23 two_stage_opamp_dummy_magic_25_0.V_err_mir_p VDDA 0.684276f
C24 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.010685f
C25 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref bgr_11_0.V_TOP 0.891713f
C26 bgr_11_0.1st_Vout_1 VDDA 1.54682f
C27 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.V_tail_gate 0.640804f
C28 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.01235f
C29 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_25_0.V_tail_gate 0.014649f
C30 two_stage_opamp_dummy_magic_25_0.cap_res_Y two_stage_opamp_dummy_magic_25_0.cap_res_X 0.345243f
C31 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.V_err_gate 0.742191f
C32 two_stage_opamp_dummy_magic_25_0.Vb1 VDDA 11.6536f
C33 bgr_11_0.Vin+ VDDA 1.74802f
C34 two_stage_opamp_dummy_magic_25_0.X two_stage_opamp_dummy_magic_25_0.cap_res_X 0.056362f
C35 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref bgr_11_0.START_UP 1.39042f
C36 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.X 0.202531f
C37 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_25_0.V_tail_gate 0.028081f
C38 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.Y 0.013749f
C39 two_stage_opamp_dummy_magic_25_0.Vb1 VOUT+ 0.110607f
C40 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.cap_res_X 2.08159f
C41 bgr_11_0.V_TOP VDDA 15.802401f
C42 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.V_tail_gate 0.169248f
C43 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C44 two_stage_opamp_dummy_magic_25_0.cap_res_X VDDA 7.87029f
C45 VIN+ VIN- 0.075694f
C46 two_stage_opamp_dummy_magic_25_0.V_err_gate VDDA 2.94416f
C47 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.cap_res_Y 0.157188f
C48 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_25_0.Vb1 0.091831f
C49 two_stage_opamp_dummy_magic_25_0.X two_stage_opamp_dummy_magic_25_0.VD1 6.06356f
C50 two_stage_opamp_dummy_magic_25_0.Y two_stage_opamp_dummy_magic_25_0.VD2 6.06356f
C51 two_stage_opamp_dummy_magic_25_0.cap_res_X VOUT+ 0.011897f
C52 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.Y 0.143814f
C53 bgr_11_0.START_UP VDDA 2.33963f
C54 two_stage_opamp_dummy_magic_25_0.Vb1 VIN+ 0.020966f
C55 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.VD1 0.015556f
C56 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.VD2 0.016071f
C57 two_stage_opamp_dummy_magic_25_0.Y two_stage_opamp_dummy_magic_25_0.cap_res_Y 0.056362f
C58 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref two_stage_opamp_dummy_magic_25_0.V_tail_gate 0.130473f
C59 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.177962f
C60 two_stage_opamp_dummy_magic_25_0.Y two_stage_opamp_dummy_magic_25_0.X 0.081053f
C61 two_stage_opamp_dummy_magic_25_0.cap_res_X VOUT- 50.9226f
C62 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.cap_res_Y 2.08159f
C63 two_stage_opamp_dummy_magic_25_0.Vb1 VIN- 0.015071f
C64 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref VDDA 6.18351f
C65 two_stage_opamp_dummy_magic_25_0.V_err_gate VOUT- 0.019632f
C66 bgr_11_0.Vin+ bgr_11_0.1st_Vout_1 0.147603f
C67 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.X 0.030556f
C68 two_stage_opamp_dummy_magic_25_0.cap_res_Y VDDA 7.87058f
C69 two_stage_opamp_dummy_magic_25_0.V_tail_gate two_stage_opamp_dummy_magic_25_0.Y 0.030556f
C70 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C71 two_stage_opamp_dummy_magic_25_0.X VDDA 8.62924f
C72 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref VOUT+ 0.020461f
C73 two_stage_opamp_dummy_magic_25_0.Y VDDA 8.69539f
C74 bgr_11_0.V_TOP bgr_11_0.1st_Vout_1 2.56012f
C75 two_stage_opamp_dummy_magic_25_0.cap_res_Y VOUT+ 50.9212f
C76 two_stage_opamp_dummy_magic_25_0.V_tail_gate VDDA 7.94882f
C77 two_stage_opamp_dummy_magic_25_0.V_err_gate two_stage_opamp_dummy_magic_25_0.V_err_mir_p 0.429395f
C78 two_stage_opamp_dummy_magic_25_0.Y VOUT+ 3.89591f
C79 two_stage_opamp_dummy_magic_25_0.V_err_gate bgr_11_0.1st_Vout_1 0.043022f
C80 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_25_0.V_err_amp_ref 0.643757f
C81 bgr_11_0.Vin+ bgr_11_0.V_TOP 1.90298f
C82 two_stage_opamp_dummy_magic_25_0.cap_res_Y VOUT- 0.011897f
C83 two_stage_opamp_dummy_magic_25_0.Vb1 two_stage_opamp_dummy_magic_25_0.cap_res_X 0.05001f
C84 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.24327f
C85 two_stage_opamp_dummy_magic_25_0.V_tail_gate VOUT+ 1.28602f
C86 two_stage_opamp_dummy_magic_25_0.VD2 VIN+ 0.533286f
C87 two_stage_opamp_dummy_magic_25_0.X VOUT- 3.89591f
C88 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.045039f
C89 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_25_0.V_err_gate 0.067034f
C90 VDDA VOUT+ 15.306099f
C91 two_stage_opamp_dummy_magic_25_0.VD1 VIN- 0.533286f
C92 VIN- GNDA 1.838f
C93 VIN+ GNDA 1.83367f
C94 VOUT- GNDA 26.046717f
C95 VOUT+ GNDA 25.908194f
C96 VDDA GNDA 0.261144p
C97 two_stage_opamp_dummy_magic_25_0.VD1 GNDA 3.177854f
C98 two_stage_opamp_dummy_magic_25_0.VD2 GNDA 3.163774f
C99 two_stage_opamp_dummy_magic_25_0.cap_res_X GNDA 41.644634f
C100 two_stage_opamp_dummy_magic_25_0.V_err_mir_p GNDA 0.106697f
C101 two_stage_opamp_dummy_magic_25_0.cap_res_Y GNDA 41.564934f
C102 two_stage_opamp_dummy_magic_25_0.X GNDA 12.164685f
C103 two_stage_opamp_dummy_magic_25_0.Y GNDA 11.827178f
C104 two_stage_opamp_dummy_magic_25_0.V_tail_gate GNDA 38.94952f
C105 two_stage_opamp_dummy_magic_25_0.Vb1 GNDA 15.744164f
C106 bgr_11_0.1st_Vout_1 GNDA 7.409633f
C107 bgr_11_0.START_UP GNDA 6.548946f
C108 bgr_11_0.START_UP_NFET1 GNDA 5.23986f
C109 two_stage_opamp_dummy_magic_25_0.V_err_gate GNDA 11.64701f
C110 bgr_11_0.V_TOP GNDA 11.27345f
C111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.2176f
C112 bgr_11_0.Vin+ GNDA 4.633147f
C113 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref GNDA 9.387731f
C114 bgr_11_0.PFET_GATE_10uA GNDA 8.581967f
C115 two_stage_opamp_dummy_magic_25_0.err_amp_out.t3 GNDA 0.036496f
C116 two_stage_opamp_dummy_magic_25_0.err_amp_out.t4 GNDA 0.08233f
C117 two_stage_opamp_dummy_magic_25_0.err_amp_out.t2 GNDA 0.036496f
C118 two_stage_opamp_dummy_magic_25_0.err_amp_out.t1 GNDA 0.036496f
C119 two_stage_opamp_dummy_magic_25_0.err_amp_out.n0 GNDA 0.114419f
C120 two_stage_opamp_dummy_magic_25_0.err_amp_out.n1 GNDA 1.7352f
C121 two_stage_opamp_dummy_magic_25_0.err_amp_out.n2 GNDA 0.122064f
C122 two_stage_opamp_dummy_magic_25_0.err_amp_out.t0 GNDA 0.036496f
C123 bgr_11_0.Vin+.t1 GNDA 0.217964f
C124 bgr_11_0.Vin+.t0 GNDA 0.09447f
C125 bgr_11_0.Vin+.n0 GNDA 1.43218f
C126 bgr_11_0.Vin+.t5 GNDA 0.03247f
C127 bgr_11_0.Vin+.t4 GNDA 0.03247f
C128 bgr_11_0.Vin+.n1 GNDA 0.082826f
C129 bgr_11_0.Vin+.t3 GNDA 0.03247f
C130 bgr_11_0.Vin+.t2 GNDA 0.03247f
C131 bgr_11_0.Vin+.n2 GNDA 0.077621f
C132 bgr_11_0.Vin+.n3 GNDA 0.774879f
C133 bgr_11_0.Vin+.n4 GNDA 0.620062f
C134 bgr_11_0.Vin+.t6 GNDA 0.051901f
C135 bgr_11_0.Vin-.n0 GNDA 0.075564f
C136 bgr_11_0.Vin-.n1 GNDA 0.084904f
C137 bgr_11_0.Vin-.n2 GNDA 0.122462f
C138 bgr_11_0.Vin-.t0 GNDA 0.283423f
C139 bgr_11_0.Vin-.t1 GNDA 0.029362f
C140 bgr_11_0.Vin-.t2 GNDA 0.029362f
C141 bgr_11_0.Vin-.n3 GNDA 0.082506f
C142 bgr_11_0.Vin-.t3 GNDA 0.029362f
C143 bgr_11_0.Vin-.t4 GNDA 0.029362f
C144 bgr_11_0.Vin-.n4 GNDA 0.071244f
C145 bgr_11_0.Vin-.n5 GNDA 0.60965f
C146 bgr_11_0.Vin-.n6 GNDA 0.030323f
C147 bgr_11_0.Vin-.n7 GNDA 0.405894f
C148 bgr_11_0.Vin-.t8 GNDA 0.047558f
C149 bgr_11_0.Vin-.n8 GNDA 0.580314f
C150 bgr_11_0.Vin-.t5 GNDA 0.123953f
C151 bgr_11_0.Vin-.n9 GNDA 0.699939f
C152 bgr_11_0.Vin-.n10 GNDA 1.30859f
C153 bgr_11_0.Vin-.n11 GNDA 0.510732f
C154 bgr_11_0.Vin-.n12 GNDA 0.076413f
C155 bgr_11_0.Vin-.n13 GNDA 0.129472f
C156 bgr_11_0.Vin-.n14 GNDA 0.075704f
C157 bgr_11_0.Vin-.n15 GNDA 0.149744f
C158 bgr_11_0.Vin-.n16 GNDA 0.149744f
C159 bgr_11_0.Vin-.n17 GNDA -0.292f
C160 bgr_11_0.Vin-.n18 GNDA 0.482615f
C161 bgr_11_0.Vin-.n19 GNDA 0.231364f
C162 bgr_11_0.Vin-.n20 GNDA 0.437116f
C163 bgr_11_0.Vin-.n21 GNDA 0.041603f
C164 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.04415f
C165 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t1 GNDA 0.155439f
C166 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t2 GNDA 0.385095f
C167 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t5 GNDA 0.457048f
C168 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t3 GNDA 0.385095f
C169 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t6 GNDA 0.457048f
C170 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n0 GNDA 0.241409f
C171 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n1 GNDA 0.271017f
C172 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n2 GNDA 0.847851f
C173 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t4 GNDA 0.385095f
C174 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t9 GNDA 0.385095f
C175 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t7 GNDA 0.457048f
C176 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n3 GNDA 0.241409f
C177 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t8 GNDA 0.457048f
C178 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n4 GNDA 0.271017f
C179 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.n5 GNDA 0.847851f
C180 two_stage_opamp_dummy_magic_25_0.V_b_2nd_stage.t0 GNDA 0.155439f
C181 bgr_11_0.cap_res1.t10 GNDA 0.331712f
C182 bgr_11_0.cap_res1.t18 GNDA 0.349187f
C183 bgr_11_0.cap_res1.t14 GNDA 0.350452f
C184 bgr_11_0.cap_res1.t3 GNDA 0.331712f
C185 bgr_11_0.cap_res1.t13 GNDA 0.349187f
C186 bgr_11_0.cap_res1.t6 GNDA 0.350452f
C187 bgr_11_0.cap_res1.t8 GNDA 0.331712f
C188 bgr_11_0.cap_res1.t17 GNDA 0.349187f
C189 bgr_11_0.cap_res1.t12 GNDA 0.350452f
C190 bgr_11_0.cap_res1.t2 GNDA 0.331712f
C191 bgr_11_0.cap_res1.t11 GNDA 0.349187f
C192 bgr_11_0.cap_res1.t5 GNDA 0.350452f
C193 bgr_11_0.cap_res1.t19 GNDA 0.331712f
C194 bgr_11_0.cap_res1.t4 GNDA 0.349187f
C195 bgr_11_0.cap_res1.t20 GNDA 0.350452f
C196 bgr_11_0.cap_res1.n0 GNDA 0.23406f
C197 bgr_11_0.cap_res1.t1 GNDA 0.186395f
C198 bgr_11_0.cap_res1.n1 GNDA 0.253961f
C199 bgr_11_0.cap_res1.t7 GNDA 0.186395f
C200 bgr_11_0.cap_res1.n2 GNDA 0.253961f
C201 bgr_11_0.cap_res1.t15 GNDA 0.186395f
C202 bgr_11_0.cap_res1.n3 GNDA 0.253961f
C203 bgr_11_0.cap_res1.t9 GNDA 0.186395f
C204 bgr_11_0.cap_res1.n4 GNDA 0.253961f
C205 bgr_11_0.cap_res1.t16 GNDA 0.363549f
C206 bgr_11_0.cap_res1.t0 GNDA 0.08421f
C207 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t7 GNDA 0.082848f
C208 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t9 GNDA 0.081431f
C209 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n0 GNDA 0.599299f
C210 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t0 GNDA 0.377424f
C211 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t8 GNDA 0.117755f
C212 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n1 GNDA 2.02279f
C213 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t2 GNDA 0.072086f
C214 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t6 GNDA 0.072086f
C215 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n2 GNDA 0.209012f
C216 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t4 GNDA 0.072086f
C217 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t5 GNDA 0.072086f
C218 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n3 GNDA 0.179801f
C219 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n4 GNDA 1.60076f
C220 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t3 GNDA 0.072086f
C221 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.t1 GNDA 0.072086f
C222 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n5 GNDA 0.179801f
C223 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n6 GNDA 1.05162f
C224 two_stage_opamp_dummy_magic_25_0.V_err_amp_ref.n7 GNDA 2.64979f
C225 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n0 GNDA 5.38141f
C226 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n1 GNDA 4.56768f
C227 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n2 GNDA 0.111227f
C228 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t15 GNDA 0.01395f
C229 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t18 GNDA 0.01395f
C230 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t30 GNDA 0.01395f
C231 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t20 GNDA 0.01395f
C232 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t12 GNDA 0.01395f
C233 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t25 GNDA 0.01395f
C234 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t16 GNDA 0.01395f
C235 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t27 GNDA 0.01395f
C236 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t22 GNDA 0.01395f
C237 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t14 GNDA 0.016282f
C238 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n3 GNDA 0.015351f
C239 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t17 GNDA 0.01395f
C240 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t26 GNDA 0.01395f
C241 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t13 GNDA 0.01395f
C242 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t21 GNDA 0.01395f
C243 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t31 GNDA 0.01395f
C244 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t19 GNDA 0.01395f
C245 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t29 GNDA 0.01395f
C246 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t24 GNDA 0.016282f
C247 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n13 GNDA 0.015351f
C248 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t28 GNDA 0.01395f
C249 two_stage_opamp_dummy_magic_25_0.V_tail_gate.t23 GNDA 0.01395f
C250 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n23 GNDA 0.010479f
C251 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n24 GNDA 0.010479f
C252 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n25 GNDA 0.110924f
C253 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n26 GNDA 0.059996f
C254 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n27 GNDA 0.010479f
C255 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n28 GNDA 0.019028f
C256 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n29 GNDA 0.059996f
C257 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n30 GNDA 0.010479f
C258 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n31 GNDA 0.111233f
C259 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n32 GNDA 0.018776f
C260 two_stage_opamp_dummy_magic_25_0.V_tail_gate.n33 GNDA 0.018776f
C261 bgr_11_0.START_UP.t4 GNDA 1.6772f
C262 bgr_11_0.START_UP.t5 GNDA 0.044089f
C263 bgr_11_0.START_UP.n0 GNDA 1.12266f
C264 bgr_11_0.START_UP.t1 GNDA 0.042075f
C265 bgr_11_0.START_UP.t3 GNDA 0.042075f
C266 bgr_11_0.START_UP.n1 GNDA 0.131329f
C267 bgr_11_0.START_UP.t2 GNDA 0.042075f
C268 bgr_11_0.START_UP.t0 GNDA 0.042075f
C269 bgr_11_0.START_UP.n2 GNDA 0.103645f
C270 bgr_11_0.START_UP.n3 GNDA 0.998514f
C271 bgr_11_0.START_UP.t6 GNDA 0.015811f
C272 bgr_11_0.START_UP.t7 GNDA 0.015811f
C273 bgr_11_0.START_UP.n4 GNDA 0.04536f
C274 bgr_11_0.START_UP.n5 GNDA 0.446231f
C275 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t2 GNDA 0.030692f
C276 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t13 GNDA 0.030692f
C277 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n0 GNDA 0.096522f
C278 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t0 GNDA 0.030692f
C279 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t1 GNDA 0.030692f
C280 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n1 GNDA 0.065837f
C281 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n2 GNDA 2.85633f
C282 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t14 GNDA 0.376143f
C283 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n3 GNDA 0.106757f
C284 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n4 GNDA 0.183688f
C285 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t12 GNDA 0.092077f
C286 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t7 GNDA 0.092077f
C287 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n5 GNDA 0.196934f
C288 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n6 GNDA 0.616009f
C289 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t3 GNDA 0.092077f
C290 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t8 GNDA 0.092077f
C291 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n7 GNDA 0.196934f
C292 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n8 GNDA 0.599325f
C293 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n9 GNDA 0.183688f
C294 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n10 GNDA 0.106757f
C295 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t5 GNDA 0.092077f
C296 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t9 GNDA 0.092077f
C297 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n11 GNDA 0.196934f
C298 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n12 GNDA 0.599325f
C299 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n13 GNDA 0.106757f
C300 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t4 GNDA 0.092077f
C301 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t11 GNDA 0.092077f
C302 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n14 GNDA 0.196934f
C303 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n15 GNDA 0.599325f
C304 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n16 GNDA 0.183688f
C305 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t6 GNDA 0.092077f
C306 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.t10 GNDA 0.092077f
C307 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n17 GNDA 0.196934f
C308 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n18 GNDA 0.607667f
C309 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n19 GNDA 0.212952f
C310 two_stage_opamp_dummy_magic_25_0.V_CMFB_S2.n20 GNDA 3.20423f
C311 bgr_11_0.V_CMFB_S2 GNDA 5.96679f
C312 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t12 GNDA 0.020331f
C313 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t15 GNDA 0.020331f
C314 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n0 GNDA 0.050962f
C315 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t11 GNDA 0.020331f
C316 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t14 GNDA 0.020331f
C317 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n1 GNDA 0.050693f
C318 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n2 GNDA 0.450559f
C319 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t16 GNDA 0.020331f
C320 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t13 GNDA 0.020331f
C321 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n3 GNDA 0.040661f
C322 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n4 GNDA 0.076236f
C323 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t0 GNDA 0.256696f
C324 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n5 GNDA 0.064224f
C325 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n6 GNDA 0.1136f
C326 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t9 GNDA 0.040661f
C327 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t4 GNDA 0.040661f
C328 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n7 GNDA 0.083136f
C329 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n8 GNDA 0.279251f
C330 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t10 GNDA 0.040661f
C331 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t5 GNDA 0.040661f
C332 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n9 GNDA 0.083136f
C333 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n10 GNDA 0.268921f
C334 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n11 GNDA 0.109199f
C335 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n12 GNDA 0.064224f
C336 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t2 GNDA 0.040661f
C337 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t6 GNDA 0.040661f
C338 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n13 GNDA 0.083136f
C339 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n14 GNDA 0.268921f
C340 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n15 GNDA 0.066572f
C341 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t1 GNDA 0.040661f
C342 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t8 GNDA 0.040661f
C343 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n16 GNDA 0.083136f
C344 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n17 GNDA 0.268921f
C345 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n18 GNDA 0.1136f
C346 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t3 GNDA 0.040661f
C347 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.t7 GNDA 0.040661f
C348 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n19 GNDA 0.083136f
C349 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n20 GNDA 0.274233f
C350 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n21 GNDA 0.148209f
C351 two_stage_opamp_dummy_magic_25_0.V_CMFB_S1.n22 GNDA 2.42166f
C352 bgr_11_0.V_CMFB_S1 GNDA 2.36838f
C353 bgr_11_0.cap_res2.t4 GNDA 0.353782f
C354 bgr_11_0.cap_res2.t9 GNDA 0.355064f
C355 bgr_11_0.cap_res2.t19 GNDA 0.336077f
C356 bgr_11_0.cap_res2.t17 GNDA 0.353782f
C357 bgr_11_0.cap_res2.t3 GNDA 0.355064f
C358 bgr_11_0.cap_res2.t13 GNDA 0.336077f
C359 bgr_11_0.cap_res2.t2 GNDA 0.353782f
C360 bgr_11_0.cap_res2.t7 GNDA 0.355064f
C361 bgr_11_0.cap_res2.t18 GNDA 0.336077f
C362 bgr_11_0.cap_res2.t16 GNDA 0.353782f
C363 bgr_11_0.cap_res2.t1 GNDA 0.355064f
C364 bgr_11_0.cap_res2.t11 GNDA 0.336077f
C365 bgr_11_0.cap_res2.t10 GNDA 0.353782f
C366 bgr_11_0.cap_res2.t15 GNDA 0.355064f
C367 bgr_11_0.cap_res2.t5 GNDA 0.336077f
C368 bgr_11_0.cap_res2.n0 GNDA 0.23714f
C369 bgr_11_0.cap_res2.t0 GNDA 0.188847f
C370 bgr_11_0.cap_res2.n1 GNDA 0.257303f
C371 bgr_11_0.cap_res2.t6 GNDA 0.188847f
C372 bgr_11_0.cap_res2.n2 GNDA 0.257303f
C373 bgr_11_0.cap_res2.t12 GNDA 0.188847f
C374 bgr_11_0.cap_res2.n3 GNDA 0.257303f
C375 bgr_11_0.cap_res2.t8 GNDA 0.188847f
C376 bgr_11_0.cap_res2.n4 GNDA 0.257303f
C377 bgr_11_0.cap_res2.t14 GNDA 0.368333f
C378 bgr_11_0.cap_res2.t20 GNDA 0.085318f
C379 bgr_11_0.1st_Vout_2.n0 GNDA 0.558332f
C380 bgr_11_0.1st_Vout_2.n1 GNDA 0.24492f
C381 bgr_11_0.1st_Vout_2.n2 GNDA 1.00873f
C382 bgr_11_0.1st_Vout_2.n3 GNDA 1.10006f
C383 bgr_11_0.1st_Vout_2.t19 GNDA 0.021918f
C384 bgr_11_0.1st_Vout_2.t27 GNDA 0.365297f
C385 bgr_11_0.1st_Vout_2.t18 GNDA 0.371519f
C386 bgr_11_0.1st_Vout_2.t11 GNDA 0.365297f
C387 bgr_11_0.1st_Vout_2.t32 GNDA 0.365297f
C388 bgr_11_0.1st_Vout_2.t25 GNDA 0.371519f
C389 bgr_11_0.1st_Vout_2.t10 GNDA 0.371519f
C390 bgr_11_0.1st_Vout_2.t30 GNDA 0.365297f
C391 bgr_11_0.1st_Vout_2.t24 GNDA 0.365297f
C392 bgr_11_0.1st_Vout_2.t17 GNDA 0.371519f
C393 bgr_11_0.1st_Vout_2.t29 GNDA 0.371519f
C394 bgr_11_0.1st_Vout_2.t23 GNDA 0.365297f
C395 bgr_11_0.1st_Vout_2.t16 GNDA 0.365297f
C396 bgr_11_0.1st_Vout_2.t8 GNDA 0.371519f
C397 bgr_11_0.1st_Vout_2.t9 GNDA 0.371519f
C398 bgr_11_0.1st_Vout_2.t28 GNDA 0.365297f
C399 bgr_11_0.1st_Vout_2.t22 GNDA 0.365297f
C400 bgr_11_0.1st_Vout_2.t14 GNDA 0.371519f
C401 bgr_11_0.1st_Vout_2.t7 GNDA 0.371519f
C402 bgr_11_0.1st_Vout_2.t13 GNDA 0.365297f
C403 bgr_11_0.1st_Vout_2.t21 GNDA 0.365297f
C404 bgr_11_0.1st_Vout_2.n4 GNDA 0.755526f
C405 bgr_11_0.1st_Vout_2.t20 GNDA 0.023864f
C406 bgr_11_0.1st_Vout_2.n5 GNDA 0.732025f
C407 bgr_11_0.1st_Vout_2.n6 GNDA 0.023021f
C408 bgr_11_0.1st_Vout_2.n7 GNDA 0.108486f
C409 bgr_11_0.1st_Vout_2.t15 GNDA 0.013912f
C410 bgr_11_0.1st_Vout_2.t31 GNDA 0.013912f
C411 bgr_11_0.1st_Vout_2.n8 GNDA 0.030949f
C412 bgr_11_0.1st_Vout_2.n9 GNDA 0.085519f
C413 bgr_11_0.1st_Vout_2.t6 GNDA 0.124099f
C414 bgr_11_0.1st_Vout_2.n10 GNDA 0.022067f
C415 bgr_11_0.1st_Vout_2.n11 GNDA 0.133286f
C416 bgr_11_0.1st_Vout_2.n12 GNDA 0.040183f
C417 bgr_11_0.1st_Vout_2.t12 GNDA 0.013912f
C418 bgr_11_0.1st_Vout_2.t26 GNDA 0.013912f
C419 bgr_11_0.1st_Vout_2.n13 GNDA 0.030949f
C420 bgr_11_0.1st_Vout_2.n14 GNDA 0.085519f
C421 bgr_11_0.1st_Vout_2.n15 GNDA 0.175152f
C422 bgr_11_0.1st_Vout_2.n16 GNDA 0.023021f
C423 bgr_11_0.V_CUR_REF_REG.t1 GNDA 0.011797f
C424 bgr_11_0.V_CUR_REF_REG.t2 GNDA 0.011797f
C425 bgr_11_0.V_CUR_REF_REG.n0 GNDA 0.081855f
C426 bgr_11_0.V_CUR_REF_REG.t3 GNDA 0.059852f
C427 bgr_11_0.V_CUR_REF_REG.n1 GNDA 2.5866f
C428 bgr_11_0.V_CUR_REF_REG.t0 GNDA 0.348101f
C429 two_stage_opamp_dummy_magic_25_0.VD1.n0 GNDA 0.259344f
C430 two_stage_opamp_dummy_magic_25_0.VD1.n1 GNDA 0.073525f
C431 two_stage_opamp_dummy_magic_25_0.VD1.n2 GNDA 0.119354f
C432 two_stage_opamp_dummy_magic_25_0.VD1.t10 GNDA 0.048999f
C433 two_stage_opamp_dummy_magic_25_0.VD1.t17 GNDA 0.048999f
C434 two_stage_opamp_dummy_magic_25_0.VD1.n3 GNDA 0.106617f
C435 two_stage_opamp_dummy_magic_25_0.VD1.n4 GNDA 0.410788f
C436 two_stage_opamp_dummy_magic_25_0.VD1.n5 GNDA 0.104207f
C437 two_stage_opamp_dummy_magic_25_0.VD1.t20 GNDA 0.048999f
C438 two_stage_opamp_dummy_magic_25_0.VD1.t14 GNDA 0.048999f
C439 two_stage_opamp_dummy_magic_25_0.VD1.n6 GNDA 0.106617f
C440 two_stage_opamp_dummy_magic_25_0.VD1.n7 GNDA 0.422242f
C441 two_stage_opamp_dummy_magic_25_0.VD1.t0 GNDA 0.048999f
C442 two_stage_opamp_dummy_magic_25_0.VD1.t5 GNDA 0.048999f
C443 two_stage_opamp_dummy_magic_25_0.VD1.n8 GNDA 0.106617f
C444 two_stage_opamp_dummy_magic_25_0.VD1.n9 GNDA 0.340702f
C445 two_stage_opamp_dummy_magic_25_0.VD1.n10 GNDA 0.097999f
C446 two_stage_opamp_dummy_magic_25_0.VD1.t4 GNDA 0.048999f
C447 two_stage_opamp_dummy_magic_25_0.VD1.t9 GNDA 0.048999f
C448 two_stage_opamp_dummy_magic_25_0.VD1.n11 GNDA 0.106617f
C449 two_stage_opamp_dummy_magic_25_0.VD1.n12 GNDA 0.340702f
C450 two_stage_opamp_dummy_magic_25_0.VD1.n13 GNDA 0.119354f
C451 two_stage_opamp_dummy_magic_25_0.VD1.t15 GNDA 0.048999f
C452 two_stage_opamp_dummy_magic_25_0.VD1.t19 GNDA 0.048999f
C453 two_stage_opamp_dummy_magic_25_0.VD1.n14 GNDA 0.106617f
C454 two_stage_opamp_dummy_magic_25_0.VD1.n15 GNDA 0.422242f
C455 two_stage_opamp_dummy_magic_25_0.VD1.n16 GNDA 0.177134f
C456 two_stage_opamp_dummy_magic_25_0.VD1.t11 GNDA 0.048999f
C457 two_stage_opamp_dummy_magic_25_0.VD1.t16 GNDA 0.048999f
C458 two_stage_opamp_dummy_magic_25_0.VD1.n17 GNDA 0.106617f
C459 two_stage_opamp_dummy_magic_25_0.VD1.n18 GNDA 0.410788f
C460 two_stage_opamp_dummy_magic_25_0.VD1.n19 GNDA 0.073525f
C461 two_stage_opamp_dummy_magic_25_0.VD1.n20 GNDA 0.185267f
C462 two_stage_opamp_dummy_magic_25_0.VD1.n21 GNDA 0.442387f
C463 two_stage_opamp_dummy_magic_25_0.VD1.n22 GNDA 0.164783f
C464 two_stage_opamp_dummy_magic_25_0.VD1.n23 GNDA 0.434039f
C465 two_stage_opamp_dummy_magic_25_0.VD1.t3 GNDA 0.048999f
C466 two_stage_opamp_dummy_magic_25_0.VD1.t7 GNDA 0.048999f
C467 two_stage_opamp_dummy_magic_25_0.VD1.n24 GNDA 0.106617f
C468 two_stage_opamp_dummy_magic_25_0.VD1.n25 GNDA 0.332043f
C469 two_stage_opamp_dummy_magic_25_0.VD1.n26 GNDA 0.187379f
C470 two_stage_opamp_dummy_magic_25_0.VD1.t1 GNDA 0.048999f
C471 two_stage_opamp_dummy_magic_25_0.VD1.t8 GNDA 0.048999f
C472 two_stage_opamp_dummy_magic_25_0.VD1.n27 GNDA 0.106617f
C473 two_stage_opamp_dummy_magic_25_0.VD1.n28 GNDA 0.332043f
C474 two_stage_opamp_dummy_magic_25_0.VD1.n29 GNDA 0.109452f
C475 two_stage_opamp_dummy_magic_25_0.VD1.n30 GNDA 0.187379f
C476 two_stage_opamp_dummy_magic_25_0.VD1.t2 GNDA 0.048999f
C477 two_stage_opamp_dummy_magic_25_0.VD1.t6 GNDA 0.048999f
C478 two_stage_opamp_dummy_magic_25_0.VD1.n31 GNDA 0.106617f
C479 two_stage_opamp_dummy_magic_25_0.VD1.n32 GNDA 0.332043f
C480 two_stage_opamp_dummy_magic_25_0.VD1.n33 GNDA 0.434039f
C481 two_stage_opamp_dummy_magic_25_0.VD1.n34 GNDA 0.164783f
C482 two_stage_opamp_dummy_magic_25_0.VD1.n35 GNDA 0.442387f
C483 two_stage_opamp_dummy_magic_25_0.VD1.n36 GNDA 0.185267f
C484 two_stage_opamp_dummy_magic_25_0.VD1.n37 GNDA 0.073525f
C485 two_stage_opamp_dummy_magic_25_0.VD1.t21 GNDA 0.048999f
C486 two_stage_opamp_dummy_magic_25_0.VD1.t13 GNDA 0.048999f
C487 two_stage_opamp_dummy_magic_25_0.VD1.n38 GNDA 0.106617f
C488 two_stage_opamp_dummy_magic_25_0.VD1.n39 GNDA 0.410788f
C489 two_stage_opamp_dummy_magic_25_0.VD1.n40 GNDA 0.177134f
C490 two_stage_opamp_dummy_magic_25_0.VD1.n41 GNDA 0.104207f
C491 two_stage_opamp_dummy_magic_25_0.VD1.t18 GNDA 0.048999f
C492 two_stage_opamp_dummy_magic_25_0.VD1.t12 GNDA 0.048999f
C493 two_stage_opamp_dummy_magic_25_0.VD1.n42 GNDA 0.106617f
C494 two_stage_opamp_dummy_magic_25_0.VD1.n43 GNDA 0.410788f
C495 two_stage_opamp_dummy_magic_25_0.VD1.n44 GNDA 0.073525f
C496 two_stage_opamp_dummy_magic_25_0.VD1.n45 GNDA 0.056907f
C497 two_stage_opamp_dummy_magic_25_0.V_tot.t1 GNDA 0.204389f
C498 two_stage_opamp_dummy_magic_25_0.V_tot.t3 GNDA 0.204389f
C499 two_stage_opamp_dummy_magic_25_0.V_tot.t2 GNDA 0.191871f
C500 two_stage_opamp_dummy_magic_25_0.V_tot.n0 GNDA 1.15943f
C501 two_stage_opamp_dummy_magic_25_0.V_tot.t4 GNDA 0.058137f
C502 two_stage_opamp_dummy_magic_25_0.V_tot.n1 GNDA 1.08618f
C503 two_stage_opamp_dummy_magic_25_0.V_tot.t5 GNDA 0.058137f
C504 two_stage_opamp_dummy_magic_25_0.V_tot.n2 GNDA 1.08618f
C505 two_stage_opamp_dummy_magic_25_0.V_tot.n3 GNDA 1.15943f
C506 two_stage_opamp_dummy_magic_25_0.V_tot.t0 GNDA 0.191871f
C507 two_stage_opamp_dummy_magic_25_0.V_err_gate.t0 GNDA 0.019597f
C508 two_stage_opamp_dummy_magic_25_0.V_err_gate.t1 GNDA 0.019597f
C509 two_stage_opamp_dummy_magic_25_0.V_err_gate.n0 GNDA 0.231028f
C510 two_stage_opamp_dummy_magic_25_0.V_err_gate.t2 GNDA 0.048991f
C511 two_stage_opamp_dummy_magic_25_0.V_err_gate.t4 GNDA 0.048991f
C512 two_stage_opamp_dummy_magic_25_0.V_err_gate.n1 GNDA 0.150096f
C513 two_stage_opamp_dummy_magic_25_0.V_err_gate.t6 GNDA 0.054707f
C514 two_stage_opamp_dummy_magic_25_0.V_err_gate.t8 GNDA 0.054707f
C515 two_stage_opamp_dummy_magic_25_0.V_err_gate.n2 GNDA 0.082174f
C516 two_stage_opamp_dummy_magic_25_0.V_err_gate.n3 GNDA 0.303282f
C517 two_stage_opamp_dummy_magic_25_0.V_err_gate.t3 GNDA 0.048991f
C518 two_stage_opamp_dummy_magic_25_0.V_err_gate.t5 GNDA 0.048991f
C519 two_stage_opamp_dummy_magic_25_0.V_err_gate.n4 GNDA 0.149445f
C520 two_stage_opamp_dummy_magic_25_0.V_err_gate.n5 GNDA 0.232053f
C521 two_stage_opamp_dummy_magic_25_0.V_err_gate.t9 GNDA 0.054707f
C522 two_stage_opamp_dummy_magic_25_0.V_err_gate.t7 GNDA 0.054707f
C523 two_stage_opamp_dummy_magic_25_0.V_err_gate.n6 GNDA 0.082174f
C524 bgr_11_0.1st_Vout_1.n0 GNDA 0.444858f
C525 bgr_11_0.1st_Vout_1.n1 GNDA 0.195143f
C526 bgr_11_0.1st_Vout_1.n2 GNDA 0.803718f
C527 bgr_11_0.1st_Vout_1.n3 GNDA 0.749146f
C528 bgr_11_0.1st_Vout_1.n4 GNDA 0.730009f
C529 bgr_11_0.1st_Vout_1.t10 GNDA 0.296012f
C530 bgr_11_0.1st_Vout_1.t31 GNDA 0.291054f
C531 bgr_11_0.1st_Vout_1.t28 GNDA 0.296012f
C532 bgr_11_0.1st_Vout_1.t9 GNDA 0.291054f
C533 bgr_11_0.1st_Vout_1.t30 GNDA 0.296012f
C534 bgr_11_0.1st_Vout_1.t24 GNDA 0.291054f
C535 bgr_11_0.1st_Vout_1.t19 GNDA 0.296012f
C536 bgr_11_0.1st_Vout_1.t27 GNDA 0.291054f
C537 bgr_11_0.1st_Vout_1.t23 GNDA 0.296012f
C538 bgr_11_0.1st_Vout_1.t14 GNDA 0.291054f
C539 bgr_11_0.1st_Vout_1.t12 GNDA 0.296012f
C540 bgr_11_0.1st_Vout_1.t18 GNDA 0.291054f
C541 bgr_11_0.1st_Vout_1.t29 GNDA 0.296012f
C542 bgr_11_0.1st_Vout_1.t22 GNDA 0.291054f
C543 bgr_11_0.1st_Vout_1.t16 GNDA 0.296012f
C544 bgr_11_0.1st_Vout_1.t26 GNDA 0.291054f
C545 bgr_11_0.1st_Vout_1.t21 GNDA 0.296012f
C546 bgr_11_0.1st_Vout_1.t13 GNDA 0.291054f
C547 bgr_11_0.1st_Vout_1.t15 GNDA 0.291054f
C548 bgr_11_0.1st_Vout_1.t11 GNDA 0.291054f
C549 bgr_11_0.1st_Vout_1.t7 GNDA 0.019014f
C550 bgr_11_0.1st_Vout_1.n5 GNDA 0.584006f
C551 bgr_11_0.1st_Vout_1.n6 GNDA 0.018342f
C552 bgr_11_0.1st_Vout_1.n7 GNDA 0.086437f
C553 bgr_11_0.1st_Vout_1.t25 GNDA 0.011085f
C554 bgr_11_0.1st_Vout_1.t32 GNDA 0.011085f
C555 bgr_11_0.1st_Vout_1.n8 GNDA 0.024659f
C556 bgr_11_0.1st_Vout_1.n9 GNDA 0.068138f
C557 bgr_11_0.1st_Vout_1.t0 GNDA 0.098878f
C558 bgr_11_0.1st_Vout_1.n10 GNDA 0.017582f
C559 bgr_11_0.1st_Vout_1.n11 GNDA 0.106197f
C560 bgr_11_0.1st_Vout_1.n12 GNDA 0.032016f
C561 bgr_11_0.1st_Vout_1.t17 GNDA 0.011085f
C562 bgr_11_0.1st_Vout_1.t8 GNDA 0.011085f
C563 bgr_11_0.1st_Vout_1.n13 GNDA 0.024659f
C564 bgr_11_0.1st_Vout_1.n14 GNDA 0.068138f
C565 bgr_11_0.1st_Vout_1.n15 GNDA 0.018342f
C566 bgr_11_0.1st_Vout_1.n16 GNDA 0.086437f
C567 bgr_11_0.1st_Vout_1.t20 GNDA 0.017398f
C568 bgr_11_0.PFET_GATE_10uA.t23 GNDA 0.023201f
C569 bgr_11_0.PFET_GATE_10uA.t15 GNDA 0.023201f
C570 bgr_11_0.PFET_GATE_10uA.n0 GNDA 0.081236f
C571 bgr_11_0.PFET_GATE_10uA.t27 GNDA 0.019989f
C572 bgr_11_0.PFET_GATE_10uA.t19 GNDA 0.029549f
C573 bgr_11_0.PFET_GATE_10uA.n1 GNDA 0.03256f
C574 bgr_11_0.PFET_GATE_10uA.t12 GNDA 0.019989f
C575 bgr_11_0.PFET_GATE_10uA.t20 GNDA 0.029549f
C576 bgr_11_0.PFET_GATE_10uA.n2 GNDA 0.03256f
C577 bgr_11_0.PFET_GATE_10uA.n3 GNDA 0.031895f
C578 bgr_11_0.PFET_GATE_10uA.n4 GNDA 1.01606f
C579 bgr_11_0.PFET_GATE_10uA.t9 GNDA 0.346712f
C580 bgr_11_0.PFET_GATE_10uA.t6 GNDA 0.305144f
C581 bgr_11_0.PFET_GATE_10uA.t7 GNDA 0.020502f
C582 bgr_11_0.PFET_GATE_10uA.t3 GNDA 0.020502f
C583 bgr_11_0.PFET_GATE_10uA.n5 GNDA 0.051047f
C584 bgr_11_0.PFET_GATE_10uA.n6 GNDA 0.838031f
C585 bgr_11_0.PFET_GATE_10uA.t5 GNDA 0.020502f
C586 bgr_11_0.PFET_GATE_10uA.t1 GNDA 0.020502f
C587 bgr_11_0.PFET_GATE_10uA.n7 GNDA 0.051047f
C588 bgr_11_0.PFET_GATE_10uA.n8 GNDA 0.414341f
C589 bgr_11_0.PFET_GATE_10uA.t4 GNDA 0.020502f
C590 bgr_11_0.PFET_GATE_10uA.t2 GNDA 0.020502f
C591 bgr_11_0.PFET_GATE_10uA.n9 GNDA 0.051047f
C592 bgr_11_0.PFET_GATE_10uA.n10 GNDA 0.414341f
C593 bgr_11_0.PFET_GATE_10uA.t0 GNDA 0.020502f
C594 bgr_11_0.PFET_GATE_10uA.t8 GNDA 0.020502f
C595 bgr_11_0.PFET_GATE_10uA.n11 GNDA 0.051047f
C596 bgr_11_0.PFET_GATE_10uA.n12 GNDA 0.654887f
C597 bgr_11_0.PFET_GATE_10uA.n13 GNDA 2.81264f
C598 bgr_11_0.PFET_GATE_10uA.t21 GNDA 0.072894f
C599 bgr_11_0.PFET_GATE_10uA.n14 GNDA 1.57977f
C600 bgr_11_0.PFET_GATE_10uA.t10 GNDA 0.019989f
C601 bgr_11_0.PFET_GATE_10uA.t24 GNDA 0.029549f
C602 bgr_11_0.PFET_GATE_10uA.n15 GNDA 0.03256f
C603 bgr_11_0.PFET_GATE_10uA.t16 GNDA 0.019989f
C604 bgr_11_0.PFET_GATE_10uA.t25 GNDA 0.029549f
C605 bgr_11_0.PFET_GATE_10uA.n16 GNDA 0.03256f
C606 bgr_11_0.PFET_GATE_10uA.n17 GNDA 0.031303f
C607 bgr_11_0.PFET_GATE_10uA.n18 GNDA 1.25111f
C608 bgr_11_0.PFET_GATE_10uA.t28 GNDA 0.019989f
C609 bgr_11_0.PFET_GATE_10uA.t14 GNDA 0.019989f
C610 bgr_11_0.PFET_GATE_10uA.t13 GNDA 0.019989f
C611 bgr_11_0.PFET_GATE_10uA.t22 GNDA 0.029549f
C612 bgr_11_0.PFET_GATE_10uA.n19 GNDA 0.036569f
C613 bgr_11_0.PFET_GATE_10uA.n20 GNDA 0.02614f
C614 bgr_11_0.PFET_GATE_10uA.n21 GNDA 0.020374f
C615 bgr_11_0.PFET_GATE_10uA.t18 GNDA 0.019989f
C616 bgr_11_0.PFET_GATE_10uA.t11 GNDA 0.019989f
C617 bgr_11_0.PFET_GATE_10uA.t26 GNDA 0.019989f
C618 bgr_11_0.PFET_GATE_10uA.t17 GNDA 0.029549f
C619 bgr_11_0.PFET_GATE_10uA.n22 GNDA 0.036569f
C620 bgr_11_0.PFET_GATE_10uA.n23 GNDA 0.02614f
C621 bgr_11_0.PFET_GATE_10uA.n24 GNDA 0.020374f
C622 bgr_11_0.PFET_GATE_10uA.n25 GNDA 0.057999f
C623 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t14 GNDA 0.028461f
C624 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t0 GNDA 0.028461f
C625 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n0 GNDA 0.089504f
C626 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t2 GNDA 0.028461f
C627 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t1 GNDA 0.028461f
C628 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n1 GNDA 0.061051f
C629 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n2 GNDA 1.86327f
C630 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t13 GNDA 0.348794f
C631 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n3 GNDA 0.098995f
C632 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n4 GNDA 0.170332f
C633 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t6 GNDA 0.085382f
C634 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t9 GNDA 0.085382f
C635 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n5 GNDA 0.182615f
C636 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n6 GNDA 0.571221f
C637 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t3 GNDA 0.085382f
C638 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t8 GNDA 0.085382f
C639 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n7 GNDA 0.182615f
C640 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n8 GNDA 0.55575f
C641 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n9 GNDA 0.170332f
C642 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n10 GNDA 0.098995f
C643 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t12 GNDA 0.085382f
C644 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t7 GNDA 0.085382f
C645 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n11 GNDA 0.182615f
C646 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n12 GNDA 0.55575f
C647 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n13 GNDA 0.098995f
C648 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t5 GNDA 0.085382f
C649 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t11 GNDA 0.085382f
C650 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n14 GNDA 0.182615f
C651 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n15 GNDA 0.55575f
C652 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n16 GNDA 0.170332f
C653 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t4 GNDA 0.085382f
C654 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.t10 GNDA 0.085382f
C655 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n17 GNDA 0.182615f
C656 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n18 GNDA 0.563485f
C657 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n19 GNDA 0.197469f
C658 two_stage_opamp_dummy_magic_25_0.V_CMFB_S4.n20 GNDA 3.03697f
C659 bgr_11_0.V_CMFB_S4 GNDA 4.512259f
C660 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t14 GNDA 0.020674f
C661 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t12 GNDA 0.020674f
C662 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n0 GNDA 0.051844f
C663 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t16 GNDA 0.020674f
C664 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t0 GNDA 0.020674f
C665 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n1 GNDA 0.051571f
C666 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n2 GNDA 0.458445f
C667 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t13 GNDA 0.020674f
C668 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t15 GNDA 0.020674f
C669 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n3 GNDA 0.041347f
C670 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n4 GNDA 0.077494f
C671 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t11 GNDA 0.260751f
C672 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n5 GNDA 0.065308f
C673 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n6 GNDA 0.115516f
C674 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t3 GNDA 0.041347f
C675 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t6 GNDA 0.041347f
C676 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n7 GNDA 0.084538f
C677 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n8 GNDA 0.283962f
C678 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t10 GNDA 0.041347f
C679 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t5 GNDA 0.041347f
C680 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n9 GNDA 0.084538f
C681 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n10 GNDA 0.273457f
C682 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n11 GNDA 0.111041f
C683 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n12 GNDA 0.065308f
C684 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t9 GNDA 0.041347f
C685 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t4 GNDA 0.041347f
C686 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n13 GNDA 0.084538f
C687 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n14 GNDA 0.273457f
C688 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n15 GNDA 0.067695f
C689 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t2 GNDA 0.041347f
C690 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t8 GNDA 0.041347f
C691 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n16 GNDA 0.084538f
C692 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n17 GNDA 0.273457f
C693 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n18 GNDA 0.115516f
C694 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t1 GNDA 0.041347f
C695 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.t7 GNDA 0.041347f
C696 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n19 GNDA 0.084538f
C697 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n20 GNDA 0.278859f
C698 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n21 GNDA 0.150709f
C699 two_stage_opamp_dummy_magic_25_0.V_CMFB_S3.n22 GNDA 2.4891f
C700 bgr_11_0.V_CMFB_S3 GNDA 2.63496f
C701 bgr_11_0.V_TOP.n0 GNDA 0.016534f
C702 bgr_11_0.V_TOP.t47 GNDA 0.126443f
C703 bgr_11_0.V_TOP.t20 GNDA 0.127563f
C704 bgr_11_0.V_TOP.t21 GNDA 0.127246f
C705 bgr_11_0.V_TOP.n1 GNDA 0.166356f
C706 bgr_11_0.V_TOP.t42 GNDA 0.127246f
C707 bgr_11_0.V_TOP.n2 GNDA 0.087699f
C708 bgr_11_0.V_TOP.t32 GNDA 0.127246f
C709 bgr_11_0.V_TOP.n3 GNDA 0.087699f
C710 bgr_11_0.V_TOP.t22 GNDA 0.127246f
C711 bgr_11_0.V_TOP.n4 GNDA 0.087699f
C712 bgr_11_0.V_TOP.t46 GNDA 0.127246f
C713 bgr_11_0.V_TOP.n5 GNDA 0.087699f
C714 bgr_11_0.V_TOP.n6 GNDA 0.024801f
C715 bgr_11_0.V_TOP.n7 GNDA 0.056353f
C716 bgr_11_0.V_TOP.t7 GNDA 0.125958f
C717 bgr_11_0.V_TOP.t17 GNDA 0.367429f
C718 bgr_11_0.V_TOP.t38 GNDA 0.373687f
C719 bgr_11_0.V_TOP.t44 GNDA 0.367429f
C720 bgr_11_0.V_TOP.n8 GNDA 0.246349f
C721 bgr_11_0.V_TOP.t36 GNDA 0.367429f
C722 bgr_11_0.V_TOP.t27 GNDA 0.373687f
C723 bgr_11_0.V_TOP.n9 GNDA 0.315242f
C724 bgr_11_0.V_TOP.t30 GNDA 0.373687f
C725 bgr_11_0.V_TOP.t35 GNDA 0.367429f
C726 bgr_11_0.V_TOP.n10 GNDA 0.246349f
C727 bgr_11_0.V_TOP.t26 GNDA 0.367429f
C728 bgr_11_0.V_TOP.t15 GNDA 0.373687f
C729 bgr_11_0.V_TOP.n11 GNDA 0.384135f
C730 bgr_11_0.V_TOP.t18 GNDA 0.373687f
C731 bgr_11_0.V_TOP.t25 GNDA 0.367429f
C732 bgr_11_0.V_TOP.n12 GNDA 0.246349f
C733 bgr_11_0.V_TOP.t14 GNDA 0.367429f
C734 bgr_11_0.V_TOP.t40 GNDA 0.373687f
C735 bgr_11_0.V_TOP.n13 GNDA 0.384135f
C736 bgr_11_0.V_TOP.t28 GNDA 0.373687f
C737 bgr_11_0.V_TOP.t33 GNDA 0.367429f
C738 bgr_11_0.V_TOP.n14 GNDA 0.246349f
C739 bgr_11_0.V_TOP.t24 GNDA 0.367429f
C740 bgr_11_0.V_TOP.t49 GNDA 0.373687f
C741 bgr_11_0.V_TOP.n15 GNDA 0.384135f
C742 bgr_11_0.V_TOP.t39 GNDA 0.373687f
C743 bgr_11_0.V_TOP.t48 GNDA 0.367429f
C744 bgr_11_0.V_TOP.n16 GNDA 0.315242f
C745 bgr_11_0.V_TOP.t23 GNDA 0.367429f
C746 bgr_11_0.V_TOP.n17 GNDA 0.16075f
C747 bgr_11_0.V_TOP.n18 GNDA 0.811818f
C748 bgr_11_0.V_TOP.t1 GNDA 0.10339f
C749 bgr_11_0.V_TOP.n19 GNDA 1.36541f
C750 bgr_11_0.V_TOP.n20 GNDA 0.022154f
C751 bgr_11_0.V_TOP.n21 GNDA 0.022154f
C752 bgr_11_0.V_TOP.n22 GNDA 0.024486f
C753 bgr_11_0.V_TOP.n23 GNDA 0.252815f
C754 bgr_11_0.V_TOP.n24 GNDA 0.138596f
C755 bgr_11_0.V_TOP.n25 GNDA 0.620324f
C756 bgr_11_0.V_TOP.n26 GNDA 0.022871f
C757 bgr_11_0.V_TOP.n27 GNDA 0.185644f
C758 bgr_11_0.V_TOP.n28 GNDA 0.022871f
C759 bgr_11_0.V_TOP.n29 GNDA 0.185644f
C760 bgr_11_0.V_TOP.n30 GNDA 0.022871f
C761 bgr_11_0.V_TOP.n31 GNDA 0.172036f
C762 bgr_11_0.V_TOP.n32 GNDA 0.347396f
C763 bgr_11_0.V_TOP.n33 GNDA 0.086346f
C764 bgr_11_0.V_TOP.t37 GNDA 0.126443f
C765 bgr_11_0.V_TOP.n34 GNDA 0.056353f
C766 bgr_11_0.V_TOP.n35 GNDA 0.024801f
C767 bgr_11_0.V_TOP.t31 GNDA 0.127246f
C768 bgr_11_0.V_TOP.n36 GNDA 0.087699f
C769 bgr_11_0.V_TOP.t19 GNDA 0.127246f
C770 bgr_11_0.V_TOP.n37 GNDA 0.087699f
C771 bgr_11_0.V_TOP.t43 GNDA 0.127246f
C772 bgr_11_0.V_TOP.n38 GNDA 0.087699f
C773 bgr_11_0.V_TOP.t45 GNDA 0.127246f
C774 bgr_11_0.V_TOP.n39 GNDA 0.087699f
C775 bgr_11_0.V_TOP.t34 GNDA 0.127246f
C776 bgr_11_0.V_TOP.n40 GNDA 0.087699f
C777 bgr_11_0.V_TOP.t29 GNDA 0.127246f
C778 bgr_11_0.V_TOP.n41 GNDA 0.087699f
C779 bgr_11_0.V_TOP.t16 GNDA 0.127246f
C780 bgr_11_0.V_TOP.n42 GNDA 0.079432f
C781 bgr_11_0.V_TOP.t41 GNDA 0.127278f
C782 two_stage_opamp_dummy_magic_25_0.Y.n0 GNDA 0.083909f
C783 two_stage_opamp_dummy_magic_25_0.Y.n1 GNDA 0.162703f
C784 two_stage_opamp_dummy_magic_25_0.Y.n2 GNDA 0.102555f
C785 two_stage_opamp_dummy_magic_25_0.Y.n3 GNDA 0.102555f
C786 two_stage_opamp_dummy_magic_25_0.Y.n4 GNDA 0.102555f
C787 two_stage_opamp_dummy_magic_25_0.Y.n5 GNDA 0.162703f
C788 two_stage_opamp_dummy_magic_25_0.Y.t9 GNDA 0.023308f
C789 two_stage_opamp_dummy_magic_25_0.Y.t22 GNDA 0.023308f
C790 two_stage_opamp_dummy_magic_25_0.Y.n6 GNDA 0.050716f
C791 two_stage_opamp_dummy_magic_25_0.Y.n7 GNDA 0.162065f
C792 two_stage_opamp_dummy_magic_25_0.Y.n8 GNDA 0.078384f
C793 two_stage_opamp_dummy_magic_25_0.Y.n9 GNDA 0.239296f
C794 two_stage_opamp_dummy_magic_25_0.Y.t21 GNDA 0.023308f
C795 two_stage_opamp_dummy_magic_25_0.Y.t7 GNDA 0.023308f
C796 two_stage_opamp_dummy_magic_25_0.Y.n10 GNDA 0.050716f
C797 two_stage_opamp_dummy_magic_25_0.Y.n11 GNDA 0.162065f
C798 two_stage_opamp_dummy_magic_25_0.Y.n12 GNDA 0.177677f
C799 two_stage_opamp_dummy_magic_25_0.Y.n13 GNDA 0.327848f
C800 two_stage_opamp_dummy_magic_25_0.Y.n14 GNDA 0.102555f
C801 two_stage_opamp_dummy_magic_25_0.Y.n15 GNDA 0.351511f
C802 two_stage_opamp_dummy_magic_25_0.Y.n16 GNDA 0.102555f
C803 two_stage_opamp_dummy_magic_25_0.Y.n17 GNDA 0.273038f
C804 two_stage_opamp_dummy_magic_25_0.Y.n18 GNDA 0.162703f
C805 two_stage_opamp_dummy_magic_25_0.Y.t2 GNDA 0.023308f
C806 two_stage_opamp_dummy_magic_25_0.Y.t5 GNDA 0.023308f
C807 two_stage_opamp_dummy_magic_25_0.Y.n19 GNDA 0.050716f
C808 two_stage_opamp_dummy_magic_25_0.Y.n20 GNDA 0.157947f
C809 two_stage_opamp_dummy_magic_25_0.Y.n21 GNDA 0.089133f
C810 two_stage_opamp_dummy_magic_25_0.Y.t0 GNDA 0.023308f
C811 two_stage_opamp_dummy_magic_25_0.Y.t3 GNDA 0.023308f
C812 two_stage_opamp_dummy_magic_25_0.Y.n22 GNDA 0.050716f
C813 two_stage_opamp_dummy_magic_25_0.Y.n23 GNDA 0.157947f
C814 two_stage_opamp_dummy_magic_25_0.Y.n24 GNDA 0.089133f
C815 two_stage_opamp_dummy_magic_25_0.Y.t1 GNDA 0.023308f
C816 two_stage_opamp_dummy_magic_25_0.Y.t4 GNDA 0.023308f
C817 two_stage_opamp_dummy_magic_25_0.Y.n25 GNDA 0.050716f
C818 two_stage_opamp_dummy_magic_25_0.Y.n26 GNDA 0.157947f
C819 two_stage_opamp_dummy_magic_25_0.Y.n27 GNDA 0.052064f
C820 two_stage_opamp_dummy_magic_25_0.Y.n28 GNDA 0.052064f
C821 two_stage_opamp_dummy_magic_25_0.Y.t8 GNDA 0.023308f
C822 two_stage_opamp_dummy_magic_25_0.Y.t6 GNDA 0.023308f
C823 two_stage_opamp_dummy_magic_25_0.Y.n29 GNDA 0.050716f
C824 two_stage_opamp_dummy_magic_25_0.Y.n30 GNDA 0.157947f
C825 two_stage_opamp_dummy_magic_25_0.Y.n31 GNDA 0.162703f
C826 two_stage_opamp_dummy_magic_25_0.Y.n32 GNDA 0.046616f
C827 two_stage_opamp_dummy_magic_25_0.Y.n33 GNDA 0.046616f
C828 two_stage_opamp_dummy_magic_25_0.Y.n34 GNDA 0.078384f
C829 two_stage_opamp_dummy_magic_25_0.Y.n35 GNDA 0.166674f
C830 two_stage_opamp_dummy_magic_25_0.Y.n36 GNDA 0.074586f
C831 two_stage_opamp_dummy_magic_25_0.Y.t54 GNDA 0.050112f
C832 two_stage_opamp_dummy_magic_25_0.Y.t38 GNDA 0.050112f
C833 two_stage_opamp_dummy_magic_25_0.Y.t27 GNDA 0.050112f
C834 two_stage_opamp_dummy_magic_25_0.Y.t42 GNDA 0.050112f
C835 two_stage_opamp_dummy_magic_25_0.Y.t49 GNDA 0.050112f
C836 two_stage_opamp_dummy_magic_25_0.Y.t31 GNDA 0.050112f
C837 two_stage_opamp_dummy_magic_25_0.Y.t51 GNDA 0.050112f
C838 two_stage_opamp_dummy_magic_25_0.Y.t33 GNDA 0.056969f
C839 two_stage_opamp_dummy_magic_25_0.Y.n39 GNDA 0.051413f
C840 two_stage_opamp_dummy_magic_25_0.Y.n40 GNDA 0.031466f
C841 two_stage_opamp_dummy_magic_25_0.Y.n41 GNDA 0.031466f
C842 two_stage_opamp_dummy_magic_25_0.Y.n42 GNDA 0.031466f
C843 two_stage_opamp_dummy_magic_25_0.Y.n43 GNDA 0.031466f
C844 two_stage_opamp_dummy_magic_25_0.Y.n44 GNDA 0.031466f
C845 two_stage_opamp_dummy_magic_25_0.Y.n45 GNDA 0.026513f
C846 two_stage_opamp_dummy_magic_25_0.Y.t34 GNDA 0.050112f
C847 two_stage_opamp_dummy_magic_25_0.Y.t43 GNDA 0.056969f
C848 two_stage_opamp_dummy_magic_25_0.Y.n46 GNDA 0.04646f
C849 two_stage_opamp_dummy_magic_25_0.Y.n47 GNDA 0.012874f
C850 two_stage_opamp_dummy_magic_25_0.Y.t26 GNDA 0.032631f
C851 two_stage_opamp_dummy_magic_25_0.Y.t41 GNDA 0.032631f
C852 two_stage_opamp_dummy_magic_25_0.Y.t29 GNDA 0.032631f
C853 two_stage_opamp_dummy_magic_25_0.Y.t45 GNDA 0.032631f
C854 two_stage_opamp_dummy_magic_25_0.Y.t50 GNDA 0.032631f
C855 two_stage_opamp_dummy_magic_25_0.Y.t32 GNDA 0.032631f
C856 two_stage_opamp_dummy_magic_25_0.Y.t53 GNDA 0.032631f
C857 two_stage_opamp_dummy_magic_25_0.Y.t36 GNDA 0.039624f
C858 two_stage_opamp_dummy_magic_25_0.Y.n48 GNDA 0.039624f
C859 two_stage_opamp_dummy_magic_25_0.Y.n49 GNDA 0.025639f
C860 two_stage_opamp_dummy_magic_25_0.Y.n50 GNDA 0.025639f
C861 two_stage_opamp_dummy_magic_25_0.Y.n51 GNDA 0.025639f
C862 two_stage_opamp_dummy_magic_25_0.Y.n52 GNDA 0.025639f
C863 two_stage_opamp_dummy_magic_25_0.Y.n53 GNDA 0.025639f
C864 two_stage_opamp_dummy_magic_25_0.Y.n54 GNDA 0.020686f
C865 two_stage_opamp_dummy_magic_25_0.Y.t37 GNDA 0.032631f
C866 two_stage_opamp_dummy_magic_25_0.Y.t46 GNDA 0.039624f
C867 two_stage_opamp_dummy_magic_25_0.Y.n55 GNDA 0.034671f
C868 two_stage_opamp_dummy_magic_25_0.Y.n56 GNDA 0.012874f
C869 two_stage_opamp_dummy_magic_25_0.Y.n57 GNDA 0.080313f
C870 two_stage_opamp_dummy_magic_25_0.Y.n58 GNDA 0.074586f
C871 two_stage_opamp_dummy_magic_25_0.Y.n59 GNDA 0.073885f
C872 two_stage_opamp_dummy_magic_25_0.Y.n60 GNDA 0.074586f
C873 two_stage_opamp_dummy_magic_25_0.Y.t20 GNDA 0.644946f
C874 two_stage_opamp_dummy_magic_25_0.Y.n61 GNDA 0.074586f
C875 two_stage_opamp_dummy_magic_25_0.Y.n62 GNDA 0.074586f
C876 two_stage_opamp_dummy_magic_25_0.Y.n64 GNDA 0.692003f
C877 two_stage_opamp_dummy_magic_25_0.Y.n66 GNDA 0.647964f
C878 two_stage_opamp_dummy_magic_25_0.Y.n67 GNDA 0.024697f
C879 two_stage_opamp_dummy_magic_25_0.Y.n68 GNDA 0.024862f
C880 two_stage_opamp_dummy_magic_25_0.Y.n69 GNDA 0.024862f
C881 two_stage_opamp_dummy_magic_25_0.Y.t47 GNDA 0.102555f
C882 two_stage_opamp_dummy_magic_25_0.Y.t52 GNDA 0.102555f
C883 two_stage_opamp_dummy_magic_25_0.Y.t35 GNDA 0.102555f
C884 two_stage_opamp_dummy_magic_25_0.Y.t25 GNDA 0.102555f
C885 two_stage_opamp_dummy_magic_25_0.Y.t39 GNDA 0.109229f
C886 two_stage_opamp_dummy_magic_25_0.Y.n70 GNDA 0.086559f
C887 two_stage_opamp_dummy_magic_25_0.Y.n71 GNDA 0.048947f
C888 two_stage_opamp_dummy_magic_25_0.Y.n72 GNDA 0.048947f
C889 two_stage_opamp_dummy_magic_25_0.Y.n73 GNDA 0.043994f
C890 two_stage_opamp_dummy_magic_25_0.Y.t30 GNDA 0.102555f
C891 two_stage_opamp_dummy_magic_25_0.Y.t44 GNDA 0.102555f
C892 two_stage_opamp_dummy_magic_25_0.Y.t28 GNDA 0.102555f
C893 two_stage_opamp_dummy_magic_25_0.Y.t40 GNDA 0.102555f
C894 two_stage_opamp_dummy_magic_25_0.Y.t48 GNDA 0.109229f
C895 two_stage_opamp_dummy_magic_25_0.Y.n74 GNDA 0.086559f
C896 two_stage_opamp_dummy_magic_25_0.Y.n75 GNDA 0.048947f
C897 two_stage_opamp_dummy_magic_25_0.Y.n76 GNDA 0.048947f
C898 two_stage_opamp_dummy_magic_25_0.Y.n77 GNDA 0.043994f
C899 two_stage_opamp_dummy_magic_25_0.Y.n78 GNDA 0.010564f
C900 two_stage_opamp_dummy_magic_25_0.Y.n79 GNDA 0.025027f
C901 two_stage_opamp_dummy_magic_25_0.Y.n80 GNDA 0.058911f
C902 two_stage_opamp_dummy_magic_25_0.Y.n81 GNDA 0.0336f
C903 two_stage_opamp_dummy_magic_25_0.Y.n82 GNDA 0.038132f
C904 two_stage_opamp_dummy_magic_25_0.Y.n83 GNDA 1.03022f
C905 two_stage_opamp_dummy_magic_25_0.Y.n84 GNDA 0.073885f
C906 two_stage_opamp_dummy_magic_25_0.Y.n85 GNDA 0.074586f
C907 two_stage_opamp_dummy_magic_25_0.Y.n86 GNDA 0.100673f
C908 two_stage_opamp_dummy_magic_25_0.Y.n87 GNDA 0.121202f
C909 two_stage_opamp_dummy_magic_25_0.Y.n88 GNDA 0.074586f
C910 two_stage_opamp_dummy_magic_25_0.Y.n89 GNDA 0.096125f
C911 two_stage_opamp_dummy_magic_25_0.Y.n90 GNDA 0.074586f
C912 two_stage_opamp_dummy_magic_25_0.Y.n91 GNDA 0.074586f
C913 two_stage_opamp_dummy_magic_25_0.Y.n92 GNDA 0.096125f
C914 two_stage_opamp_dummy_magic_25_0.Y.n93 GNDA 0.074586f
C915 two_stage_opamp_dummy_magic_25_0.Y.n94 GNDA 0.122901f
C916 two_stage_opamp_dummy_magic_25_0.Y.t14 GNDA 0.054385f
C917 two_stage_opamp_dummy_magic_25_0.Y.t17 GNDA 0.054385f
C918 two_stage_opamp_dummy_magic_25_0.Y.n95 GNDA 0.111251f
C919 two_stage_opamp_dummy_magic_25_0.Y.n96 GNDA 0.297688f
C920 two_stage_opamp_dummy_magic_25_0.Y.t23 GNDA 0.054385f
C921 two_stage_opamp_dummy_magic_25_0.Y.t12 GNDA 0.054385f
C922 two_stage_opamp_dummy_magic_25_0.Y.n97 GNDA 0.111251f
C923 two_stage_opamp_dummy_magic_25_0.Y.n98 GNDA 0.302606f
C924 two_stage_opamp_dummy_magic_25_0.Y.n99 GNDA 0.100632f
C925 two_stage_opamp_dummy_magic_25_0.Y.t19 GNDA 0.054385f
C926 two_stage_opamp_dummy_magic_25_0.Y.t10 GNDA 0.054385f
C927 two_stage_opamp_dummy_magic_25_0.Y.n100 GNDA 0.111251f
C928 two_stage_opamp_dummy_magic_25_0.Y.n101 GNDA 0.297688f
C929 two_stage_opamp_dummy_magic_25_0.Y.n102 GNDA 0.058991f
C930 two_stage_opamp_dummy_magic_25_0.Y.t11 GNDA 0.054385f
C931 two_stage_opamp_dummy_magic_25_0.Y.t13 GNDA 0.054385f
C932 two_stage_opamp_dummy_magic_25_0.Y.n103 GNDA 0.111251f
C933 two_stage_opamp_dummy_magic_25_0.Y.n104 GNDA 0.297688f
C934 two_stage_opamp_dummy_magic_25_0.Y.n105 GNDA 0.058991f
C935 two_stage_opamp_dummy_magic_25_0.Y.t16 GNDA 0.054385f
C936 two_stage_opamp_dummy_magic_25_0.Y.t24 GNDA 0.054385f
C937 two_stage_opamp_dummy_magic_25_0.Y.n106 GNDA 0.111251f
C938 two_stage_opamp_dummy_magic_25_0.Y.n107 GNDA 0.302606f
C939 two_stage_opamp_dummy_magic_25_0.Y.n108 GNDA 0.100632f
C940 two_stage_opamp_dummy_magic_25_0.Y.t15 GNDA 0.054385f
C941 two_stage_opamp_dummy_magic_25_0.Y.t18 GNDA 0.054385f
C942 two_stage_opamp_dummy_magic_25_0.Y.n109 GNDA 0.111251f
C943 two_stage_opamp_dummy_magic_25_0.Y.n110 GNDA 0.297688f
C944 two_stage_opamp_dummy_magic_25_0.Y.n111 GNDA 0.096125f
C945 two_stage_opamp_dummy_magic_25_0.Y.n112 GNDA 0.082469f
C946 two_stage_opamp_dummy_magic_25_0.Y.n113 GNDA 0.049724f
C947 two_stage_opamp_dummy_magic_25_0.Y.n114 GNDA 0.049724f
C948 two_stage_opamp_dummy_magic_25_0.Y.n115 GNDA 0.082469f
C949 two_stage_opamp_dummy_magic_25_0.Y.n116 GNDA 0.096125f
C950 two_stage_opamp_dummy_magic_25_0.Y.n117 GNDA 0.170057f
C951 two_stage_opamp_dummy_magic_25_0.Y.n118 GNDA 0.251893f
C952 two_stage_opamp_dummy_magic_25_0.Y.n119 GNDA 0.320326f
C953 two_stage_opamp_dummy_magic_25_0.Y.n120 GNDA 0.074586f
C954 two_stage_opamp_dummy_magic_25_0.Y.n121 GNDA 0.074586f
C955 two_stage_opamp_dummy_magic_25_0.Y.n122 GNDA 0.121202f
C956 two_stage_opamp_dummy_magic_25_0.Y.n123 GNDA 0.074586f
C957 two_stage_opamp_dummy_magic_25_0.Y.n124 GNDA 0.074586f
C958 two_stage_opamp_dummy_magic_25_0.Y.n125 GNDA 0.074586f
C959 two_stage_opamp_dummy_magic_25_0.Y.n126 GNDA 0.074586f
C960 two_stage_opamp_dummy_magic_25_0.Y.n127 GNDA 0.121202f
C961 two_stage_opamp_dummy_magic_25_0.Y.n128 GNDA 0.074586f
C962 two_stage_opamp_dummy_magic_25_0.Y.n129 GNDA 0.074586f
C963 two_stage_opamp_dummy_magic_25_0.Y.n130 GNDA 0.074586f
C964 two_stage_opamp_dummy_magic_25_0.Y.n131 GNDA 0.074586f
C965 two_stage_opamp_dummy_magic_25_0.Y.n132 GNDA 0.074586f
C966 two_stage_opamp_dummy_magic_25_0.Y.n133 GNDA 0.074586f
C967 two_stage_opamp_dummy_magic_25_0.Y.n134 GNDA 0.074586f
C968 two_stage_opamp_dummy_magic_25_0.Y.n135 GNDA 0.121202f
C969 two_stage_opamp_dummy_magic_25_0.Y.n136 GNDA 0.582701f
C970 two_stage_opamp_dummy_magic_25_0.Y.n137 GNDA 0.582701f
C971 two_stage_opamp_dummy_magic_25_0.Y.n138 GNDA 0.074586f
C972 two_stage_opamp_dummy_magic_25_0.Y.n140 GNDA 0.074586f
C973 two_stage_opamp_dummy_magic_25_0.Y.n141 GNDA 0.074586f
C974 two_stage_opamp_dummy_magic_25_0.Y.n143 GNDA 0.913675f
C975 two_stage_opamp_dummy_magic_25_0.Y.n144 GNDA 0.913675f
C976 two_stage_opamp_dummy_magic_25_0.Y.n146 GNDA 0.456838f
C977 two_stage_opamp_dummy_magic_25_0.Y.n147 GNDA 2.20415f
C978 two_stage_opamp_dummy_magic_25_0.Y.n148 GNDA 0.601348f
C979 two_stage_opamp_dummy_magic_25_0.Y.n149 GNDA 0.615332f
C980 two_stage_opamp_dummy_magic_25_0.Y.n150 GNDA 0.225311f
C981 two_stage_opamp_dummy_magic_25_0.Y.n151 GNDA 0.102555f
C982 two_stage_opamp_dummy_magic_25_0.Y.n152 GNDA 0.239296f
C983 two_stage_opamp_dummy_magic_25_0.Y.n153 GNDA 0.102555f
C984 two_stage_opamp_dummy_magic_25_0.Y.n154 GNDA 0.102555f
C985 two_stage_opamp_dummy_magic_25_0.Y.n155 GNDA 0.102555f
C986 two_stage_opamp_dummy_magic_25_0.Y.n156 GNDA 0.206665f
C987 two_stage_opamp_dummy_magic_25_0.Vb1_2.t1 GNDA 0.046205f
C988 two_stage_opamp_dummy_magic_25_0.Vb1_2.n0 GNDA 0.312531f
C989 two_stage_opamp_dummy_magic_25_0.Vb1_2.t4 GNDA 0.157018f
C990 two_stage_opamp_dummy_magic_25_0.Vb1_2.n1 GNDA 0.539239f
C991 two_stage_opamp_dummy_magic_25_0.Vb1_2.t2 GNDA 0.046205f
C992 two_stage_opamp_dummy_magic_25_0.Vb1_2.t0 GNDA 0.046205f
C993 two_stage_opamp_dummy_magic_25_0.Vb1_2.n2 GNDA 0.100536f
C994 two_stage_opamp_dummy_magic_25_0.Vb1_2.n3 GNDA 0.474689f
C995 two_stage_opamp_dummy_magic_25_0.Vb1_2.n4 GNDA 0.470919f
C996 two_stage_opamp_dummy_magic_25_0.Vb1_2.n5 GNDA 0.459714f
C997 two_stage_opamp_dummy_magic_25_0.Vb1_2.n6 GNDA 0.100536f
C998 two_stage_opamp_dummy_magic_25_0.Vb1_2.t3 GNDA 0.046205f
C999 two_stage_opamp_dummy_magic_25_0.Vb1.n0 GNDA 0.259977f
C1000 two_stage_opamp_dummy_magic_25_0.Vb1.n1 GNDA 4.25266f
C1001 two_stage_opamp_dummy_magic_25_0.Vb1.n2 GNDA 0.217042f
C1002 two_stage_opamp_dummy_magic_25_0.Vb1.n3 GNDA 0.369053f
C1003 two_stage_opamp_dummy_magic_25_0.Vb1.n4 GNDA 0.177764f
C1004 two_stage_opamp_dummy_magic_25_0.Vb1.n5 GNDA 0.369053f
C1005 two_stage_opamp_dummy_magic_25_0.Vb1.t11 GNDA 0.037665f
C1006 two_stage_opamp_dummy_magic_25_0.Vb1.t8 GNDA 0.037665f
C1007 two_stage_opamp_dummy_magic_25_0.Vb1.n6 GNDA 0.085691f
C1008 two_stage_opamp_dummy_magic_25_0.Vb1.t2 GNDA 0.028955f
C1009 two_stage_opamp_dummy_magic_25_0.Vb1.t4 GNDA 0.037556f
C1010 two_stage_opamp_dummy_magic_25_0.Vb1.n7 GNDA 0.038612f
C1011 two_stage_opamp_dummy_magic_25_0.Vb1.t0 GNDA 0.028955f
C1012 two_stage_opamp_dummy_magic_25_0.Vb1.t6 GNDA 0.037556f
C1013 two_stage_opamp_dummy_magic_25_0.Vb1.n8 GNDA 0.038612f
C1014 two_stage_opamp_dummy_magic_25_0.Vb1.n9 GNDA 0.028781f
C1015 two_stage_opamp_dummy_magic_25_0.Vb1.t12 GNDA 1.08636f
C1016 two_stage_opamp_dummy_magic_25_0.Vb1.t9 GNDA 0.028249f
C1017 two_stage_opamp_dummy_magic_25_0.Vb1.t5 GNDA 0.028249f
C1018 two_stage_opamp_dummy_magic_25_0.Vb1.n10 GNDA 0.061466f
C1019 two_stage_opamp_dummy_magic_25_0.Vb1.n11 GNDA 0.227076f
C1020 two_stage_opamp_dummy_magic_25_0.Vb1.t3 GNDA 0.028249f
C1021 two_stage_opamp_dummy_magic_25_0.Vb1.t1 GNDA 0.028249f
C1022 two_stage_opamp_dummy_magic_25_0.Vb1.n12 GNDA 0.061466f
C1023 two_stage_opamp_dummy_magic_25_0.Vb1.t7 GNDA 0.028249f
C1024 two_stage_opamp_dummy_magic_25_0.Vb1.t10 GNDA 0.028249f
C1025 two_stage_opamp_dummy_magic_25_0.Vb1.n13 GNDA 0.0715f
C1026 two_stage_opamp_dummy_magic_25_0.Vb1.t14 GNDA 0.028955f
C1027 two_stage_opamp_dummy_magic_25_0.Vb1.t25 GNDA 0.028955f
C1028 two_stage_opamp_dummy_magic_25_0.Vb1.t32 GNDA 0.028955f
C1029 two_stage_opamp_dummy_magic_25_0.Vb1.t24 GNDA 0.028955f
C1030 two_stage_opamp_dummy_magic_25_0.Vb1.t31 GNDA 0.028955f
C1031 two_stage_opamp_dummy_magic_25_0.Vb1.t22 GNDA 0.028955f
C1032 two_stage_opamp_dummy_magic_25_0.Vb1.t17 GNDA 0.028955f
C1033 two_stage_opamp_dummy_magic_25_0.Vb1.t23 GNDA 0.028955f
C1034 two_stage_opamp_dummy_magic_25_0.Vb1.t30 GNDA 0.028955f
C1035 two_stage_opamp_dummy_magic_25_0.Vb1.t19 GNDA 0.028955f
C1036 two_stage_opamp_dummy_magic_25_0.Vb1.t29 GNDA 0.028955f
C1037 two_stage_opamp_dummy_magic_25_0.Vb1.t18 GNDA 0.028955f
C1038 two_stage_opamp_dummy_magic_25_0.Vb1.t27 GNDA 0.028955f
C1039 two_stage_opamp_dummy_magic_25_0.Vb1.t15 GNDA 0.028955f
C1040 two_stage_opamp_dummy_magic_25_0.Vb1.t28 GNDA 0.028955f
C1041 two_stage_opamp_dummy_magic_25_0.Vb1.t16 GNDA 0.028955f
C1042 two_stage_opamp_dummy_magic_25_0.Vb1.t26 GNDA 0.028955f
C1043 two_stage_opamp_dummy_magic_25_0.Vb1.t13 GNDA 0.028955f
C1044 two_stage_opamp_dummy_magic_25_0.Vb1.t20 GNDA 0.037556f
C1045 two_stage_opamp_dummy_magic_25_0.Vb1.n14 GNDA 0.040835f
C1046 two_stage_opamp_dummy_magic_25_0.Vb1.n15 GNDA 0.027542f
C1047 two_stage_opamp_dummy_magic_25_0.Vb1.n16 GNDA 0.027542f
C1048 two_stage_opamp_dummy_magic_25_0.Vb1.n17 GNDA 0.027542f
C1049 two_stage_opamp_dummy_magic_25_0.Vb1.n18 GNDA 0.027542f
C1050 two_stage_opamp_dummy_magic_25_0.Vb1.n19 GNDA 0.027542f
C1051 two_stage_opamp_dummy_magic_25_0.Vb1.n20 GNDA 0.027542f
C1052 two_stage_opamp_dummy_magic_25_0.Vb1.n21 GNDA 0.027542f
C1053 two_stage_opamp_dummy_magic_25_0.Vb1.n22 GNDA 0.049428f
C1054 two_stage_opamp_dummy_magic_25_0.Vb1.t21 GNDA 0.028955f
C1055 two_stage_opamp_dummy_magic_25_0.Vb1.n23 GNDA 0.049428f
C1056 two_stage_opamp_dummy_magic_25_0.Vb1.n24 GNDA 0.027542f
C1057 two_stage_opamp_dummy_magic_25_0.Vb1.n25 GNDA 0.027542f
C1058 two_stage_opamp_dummy_magic_25_0.Vb1.n26 GNDA 0.027542f
C1059 two_stage_opamp_dummy_magic_25_0.Vb1.n27 GNDA 0.027542f
C1060 two_stage_opamp_dummy_magic_25_0.Vb1.n28 GNDA 0.027542f
C1061 two_stage_opamp_dummy_magic_25_0.Vb1.n29 GNDA 0.027542f
C1062 two_stage_opamp_dummy_magic_25_0.Vb1.n30 GNDA 0.027542f
C1063 two_stage_opamp_dummy_magic_25_0.Vb1.n31 GNDA 0.027542f
C1064 two_stage_opamp_dummy_magic_25_0.Vb1.n32 GNDA 0.050581f
C1065 two_stage_opamp_dummy_magic_25_0.Vb1.n33 GNDA 5.63417f
C1066 two_stage_opamp_dummy_magic_25_0.VD2.n0 GNDA 0.259344f
C1067 two_stage_opamp_dummy_magic_25_0.VD2.n1 GNDA 0.073525f
C1068 two_stage_opamp_dummy_magic_25_0.VD2.n2 GNDA 0.119354f
C1069 two_stage_opamp_dummy_magic_25_0.VD2.t11 GNDA 0.048999f
C1070 two_stage_opamp_dummy_magic_25_0.VD2.t9 GNDA 0.048999f
C1071 two_stage_opamp_dummy_magic_25_0.VD2.n3 GNDA 0.106617f
C1072 two_stage_opamp_dummy_magic_25_0.VD2.n4 GNDA 0.410788f
C1073 two_stage_opamp_dummy_magic_25_0.VD2.n5 GNDA 0.104207f
C1074 two_stage_opamp_dummy_magic_25_0.VD2.t12 GNDA 0.048999f
C1075 two_stage_opamp_dummy_magic_25_0.VD2.t18 GNDA 0.048999f
C1076 two_stage_opamp_dummy_magic_25_0.VD2.n6 GNDA 0.106617f
C1077 two_stage_opamp_dummy_magic_25_0.VD2.n7 GNDA 0.422242f
C1078 two_stage_opamp_dummy_magic_25_0.VD2.t1 GNDA 0.048999f
C1079 two_stage_opamp_dummy_magic_25_0.VD2.t3 GNDA 0.048999f
C1080 two_stage_opamp_dummy_magic_25_0.VD2.n8 GNDA 0.106617f
C1081 two_stage_opamp_dummy_magic_25_0.VD2.n9 GNDA 0.340702f
C1082 two_stage_opamp_dummy_magic_25_0.VD2.n10 GNDA 0.097999f
C1083 two_stage_opamp_dummy_magic_25_0.VD2.t19 GNDA 0.048999f
C1084 two_stage_opamp_dummy_magic_25_0.VD2.t5 GNDA 0.048999f
C1085 two_stage_opamp_dummy_magic_25_0.VD2.n11 GNDA 0.106617f
C1086 two_stage_opamp_dummy_magic_25_0.VD2.n12 GNDA 0.340702f
C1087 two_stage_opamp_dummy_magic_25_0.VD2.n13 GNDA 0.119354f
C1088 two_stage_opamp_dummy_magic_25_0.VD2.t17 GNDA 0.048999f
C1089 two_stage_opamp_dummy_magic_25_0.VD2.t10 GNDA 0.048999f
C1090 two_stage_opamp_dummy_magic_25_0.VD2.n14 GNDA 0.106617f
C1091 two_stage_opamp_dummy_magic_25_0.VD2.n15 GNDA 0.422242f
C1092 two_stage_opamp_dummy_magic_25_0.VD2.n16 GNDA 0.177134f
C1093 two_stage_opamp_dummy_magic_25_0.VD2.t15 GNDA 0.048999f
C1094 two_stage_opamp_dummy_magic_25_0.VD2.t8 GNDA 0.048999f
C1095 two_stage_opamp_dummy_magic_25_0.VD2.n17 GNDA 0.106617f
C1096 two_stage_opamp_dummy_magic_25_0.VD2.n18 GNDA 0.410788f
C1097 two_stage_opamp_dummy_magic_25_0.VD2.n19 GNDA 0.073525f
C1098 two_stage_opamp_dummy_magic_25_0.VD2.n20 GNDA 0.185267f
C1099 two_stage_opamp_dummy_magic_25_0.VD2.n21 GNDA 0.442387f
C1100 two_stage_opamp_dummy_magic_25_0.VD2.n22 GNDA 0.164783f
C1101 two_stage_opamp_dummy_magic_25_0.VD2.n23 GNDA 0.434039f
C1102 two_stage_opamp_dummy_magic_25_0.VD2.t6 GNDA 0.048999f
C1103 two_stage_opamp_dummy_magic_25_0.VD2.t0 GNDA 0.048999f
C1104 two_stage_opamp_dummy_magic_25_0.VD2.n24 GNDA 0.106617f
C1105 two_stage_opamp_dummy_magic_25_0.VD2.n25 GNDA 0.332043f
C1106 two_stage_opamp_dummy_magic_25_0.VD2.n26 GNDA 0.187379f
C1107 two_stage_opamp_dummy_magic_25_0.VD2.t21 GNDA 0.048999f
C1108 two_stage_opamp_dummy_magic_25_0.VD2.t4 GNDA 0.048999f
C1109 two_stage_opamp_dummy_magic_25_0.VD2.n27 GNDA 0.106617f
C1110 two_stage_opamp_dummy_magic_25_0.VD2.n28 GNDA 0.332043f
C1111 two_stage_opamp_dummy_magic_25_0.VD2.n29 GNDA 0.109452f
C1112 two_stage_opamp_dummy_magic_25_0.VD2.n30 GNDA 0.187379f
C1113 two_stage_opamp_dummy_magic_25_0.VD2.t2 GNDA 0.048999f
C1114 two_stage_opamp_dummy_magic_25_0.VD2.t20 GNDA 0.048999f
C1115 two_stage_opamp_dummy_magic_25_0.VD2.n31 GNDA 0.106617f
C1116 two_stage_opamp_dummy_magic_25_0.VD2.n32 GNDA 0.332043f
C1117 two_stage_opamp_dummy_magic_25_0.VD2.n33 GNDA 0.434039f
C1118 two_stage_opamp_dummy_magic_25_0.VD2.n34 GNDA 0.164783f
C1119 two_stage_opamp_dummy_magic_25_0.VD2.n35 GNDA 0.442387f
C1120 two_stage_opamp_dummy_magic_25_0.VD2.n36 GNDA 0.185267f
C1121 two_stage_opamp_dummy_magic_25_0.VD2.n37 GNDA 0.073525f
C1122 two_stage_opamp_dummy_magic_25_0.VD2.t13 GNDA 0.048999f
C1123 two_stage_opamp_dummy_magic_25_0.VD2.t16 GNDA 0.048999f
C1124 two_stage_opamp_dummy_magic_25_0.VD2.n38 GNDA 0.106617f
C1125 two_stage_opamp_dummy_magic_25_0.VD2.n39 GNDA 0.410788f
C1126 two_stage_opamp_dummy_magic_25_0.VD2.n40 GNDA 0.177134f
C1127 two_stage_opamp_dummy_magic_25_0.VD2.n41 GNDA 0.104207f
C1128 two_stage_opamp_dummy_magic_25_0.VD2.t14 GNDA 0.048999f
C1129 two_stage_opamp_dummy_magic_25_0.VD2.t7 GNDA 0.048999f
C1130 two_stage_opamp_dummy_magic_25_0.VD2.n42 GNDA 0.106617f
C1131 two_stage_opamp_dummy_magic_25_0.VD2.n43 GNDA 0.410788f
C1132 two_stage_opamp_dummy_magic_25_0.VD2.n44 GNDA 0.073525f
C1133 two_stage_opamp_dummy_magic_25_0.VD2.n45 GNDA 0.056907f
C1134 two_stage_opamp_dummy_magic_25_0.V_source.n0 GNDA 0.232841f
C1135 two_stage_opamp_dummy_magic_25_0.V_source.n1 GNDA 0.195116f
C1136 two_stage_opamp_dummy_magic_25_0.V_source.n2 GNDA 0.195116f
C1137 two_stage_opamp_dummy_magic_25_0.V_source.n3 GNDA 0.252385f
C1138 two_stage_opamp_dummy_magic_25_0.V_source.n4 GNDA 0.273514f
C1139 two_stage_opamp_dummy_magic_25_0.V_source.n5 GNDA 0.175967f
C1140 two_stage_opamp_dummy_magic_25_0.V_source.n6 GNDA 0.138292f
C1141 two_stage_opamp_dummy_magic_25_0.V_source.n7 GNDA 0.138292f
C1142 two_stage_opamp_dummy_magic_25_0.V_source.n8 GNDA 0.185434f
C1143 two_stage_opamp_dummy_magic_25_0.V_source.n9 GNDA 0.215081f
C1144 two_stage_opamp_dummy_magic_25_0.V_source.n10 GNDA 2.10776f
C1145 two_stage_opamp_dummy_magic_25_0.V_source.n11 GNDA 2.14775f
C1146 two_stage_opamp_dummy_magic_25_0.V_source.t24 GNDA 0.033909f
C1147 two_stage_opamp_dummy_magic_25_0.V_source.t5 GNDA 0.033909f
C1148 two_stage_opamp_dummy_magic_25_0.V_source.n12 GNDA 0.072491f
C1149 two_stage_opamp_dummy_magic_25_0.V_source.t7 GNDA 0.033909f
C1150 two_stage_opamp_dummy_magic_25_0.V_source.t35 GNDA 0.033909f
C1151 two_stage_opamp_dummy_magic_25_0.V_source.n13 GNDA 0.072491f
C1152 two_stage_opamp_dummy_magic_25_0.V_source.n14 GNDA 0.215081f
C1153 two_stage_opamp_dummy_magic_25_0.V_source.t31 GNDA 0.033909f
C1154 two_stage_opamp_dummy_magic_25_0.V_source.t37 GNDA 0.033909f
C1155 two_stage_opamp_dummy_magic_25_0.V_source.n15 GNDA 0.072491f
C1156 two_stage_opamp_dummy_magic_25_0.V_source.n16 GNDA 0.166395f
C1157 two_stage_opamp_dummy_magic_25_0.V_source.t11 GNDA 0.075228f
C1158 two_stage_opamp_dummy_magic_25_0.V_source.n17 GNDA 0.31862f
C1159 two_stage_opamp_dummy_magic_25_0.V_source.t8 GNDA 0.033909f
C1160 two_stage_opamp_dummy_magic_25_0.V_source.t6 GNDA 0.033909f
C1161 two_stage_opamp_dummy_magic_25_0.V_source.n18 GNDA 0.072491f
C1162 two_stage_opamp_dummy_magic_25_0.V_source.n19 GNDA 0.215081f
C1163 two_stage_opamp_dummy_magic_25_0.V_source.n20 GNDA 0.07397f
C1164 two_stage_opamp_dummy_magic_25_0.V_source.t29 GNDA 0.020345f
C1165 two_stage_opamp_dummy_magic_25_0.V_source.t1 GNDA 0.020345f
C1166 two_stage_opamp_dummy_magic_25_0.V_source.n21 GNDA 0.044269f
C1167 two_stage_opamp_dummy_magic_25_0.V_source.n22 GNDA 0.185793f
C1168 two_stage_opamp_dummy_magic_25_0.V_source.t26 GNDA 0.020345f
C1169 two_stage_opamp_dummy_magic_25_0.V_source.t0 GNDA 0.020345f
C1170 two_stage_opamp_dummy_magic_25_0.V_source.n23 GNDA 0.044269f
C1171 two_stage_opamp_dummy_magic_25_0.V_source.n24 GNDA 0.179367f
C1172 two_stage_opamp_dummy_magic_25_0.V_source.t27 GNDA 0.020345f
C1173 two_stage_opamp_dummy_magic_25_0.V_source.t28 GNDA 0.020345f
C1174 two_stage_opamp_dummy_magic_25_0.V_source.n25 GNDA 0.044269f
C1175 two_stage_opamp_dummy_magic_25_0.V_source.n26 GNDA 0.179367f
C1176 two_stage_opamp_dummy_magic_25_0.V_source.n27 GNDA 0.043484f
C1177 two_stage_opamp_dummy_magic_25_0.V_source.n28 GNDA 0.043484f
C1178 two_stage_opamp_dummy_magic_25_0.V_source.t2 GNDA 0.020345f
C1179 two_stage_opamp_dummy_magic_25_0.V_source.t38 GNDA 0.020345f
C1180 two_stage_opamp_dummy_magic_25_0.V_source.n29 GNDA 0.044269f
C1181 two_stage_opamp_dummy_magic_25_0.V_source.n30 GNDA 0.134349f
C1182 two_stage_opamp_dummy_magic_25_0.V_source.t9 GNDA 0.020345f
C1183 two_stage_opamp_dummy_magic_25_0.V_source.t32 GNDA 0.020345f
C1184 two_stage_opamp_dummy_magic_25_0.V_source.n31 GNDA 0.044269f
C1185 two_stage_opamp_dummy_magic_25_0.V_source.n32 GNDA 0.134349f
C1186 two_stage_opamp_dummy_magic_25_0.V_source.n33 GNDA 0.109945f
C1187 two_stage_opamp_dummy_magic_25_0.V_source.t17 GNDA 0.020345f
C1188 two_stage_opamp_dummy_magic_25_0.V_source.t12 GNDA 0.020345f
C1189 two_stage_opamp_dummy_magic_25_0.V_source.n34 GNDA 0.044269f
C1190 two_stage_opamp_dummy_magic_25_0.V_source.n35 GNDA 0.134349f
C1191 two_stage_opamp_dummy_magic_25_0.V_source.n36 GNDA 0.109945f
C1192 two_stage_opamp_dummy_magic_25_0.V_source.t16 GNDA 0.020345f
C1193 two_stage_opamp_dummy_magic_25_0.V_source.t18 GNDA 0.020345f
C1194 two_stage_opamp_dummy_magic_25_0.V_source.n37 GNDA 0.044269f
C1195 two_stage_opamp_dummy_magic_25_0.V_source.n38 GNDA 0.134349f
C1196 two_stage_opamp_dummy_magic_25_0.V_source.n39 GNDA 0.043484f
C1197 two_stage_opamp_dummy_magic_25_0.V_source.t13 GNDA 0.020345f
C1198 two_stage_opamp_dummy_magic_25_0.V_source.t14 GNDA 0.020345f
C1199 two_stage_opamp_dummy_magic_25_0.V_source.n40 GNDA 0.044269f
C1200 two_stage_opamp_dummy_magic_25_0.V_source.n41 GNDA 0.185793f
C1201 two_stage_opamp_dummy_magic_25_0.V_source.t15 GNDA 0.020345f
C1202 two_stage_opamp_dummy_magic_25_0.V_source.t21 GNDA 0.020345f
C1203 two_stage_opamp_dummy_magic_25_0.V_source.n42 GNDA 0.044269f
C1204 two_stage_opamp_dummy_magic_25_0.V_source.n43 GNDA 0.179367f
C1205 two_stage_opamp_dummy_magic_25_0.V_source.n44 GNDA 0.07397f
C1206 two_stage_opamp_dummy_magic_25_0.V_source.n45 GNDA 0.043484f
C1207 two_stage_opamp_dummy_magic_25_0.V_source.t20 GNDA 0.020345f
C1208 two_stage_opamp_dummy_magic_25_0.V_source.t19 GNDA 0.020345f
C1209 two_stage_opamp_dummy_magic_25_0.V_source.n46 GNDA 0.044269f
C1210 two_stage_opamp_dummy_magic_25_0.V_source.n47 GNDA 0.179367f
C1211 two_stage_opamp_dummy_magic_25_0.V_source.n48 GNDA 0.232841f
C1212 two_stage_opamp_dummy_magic_25_0.V_source.t33 GNDA 0.033909f
C1213 two_stage_opamp_dummy_magic_25_0.V_source.t40 GNDA 0.033909f
C1214 two_stage_opamp_dummy_magic_25_0.V_source.n49 GNDA 0.072491f
C1215 two_stage_opamp_dummy_magic_25_0.V_source.t22 GNDA 0.033909f
C1216 two_stage_opamp_dummy_magic_25_0.V_source.t39 GNDA 0.033909f
C1217 two_stage_opamp_dummy_magic_25_0.V_source.n50 GNDA 0.072491f
C1218 two_stage_opamp_dummy_magic_25_0.V_source.n51 GNDA 0.218096f
C1219 two_stage_opamp_dummy_magic_25_0.V_source.t3 GNDA 0.033909f
C1220 two_stage_opamp_dummy_magic_25_0.V_source.t23 GNDA 0.033909f
C1221 two_stage_opamp_dummy_magic_25_0.V_source.n52 GNDA 0.072491f
C1222 two_stage_opamp_dummy_magic_25_0.V_source.n53 GNDA 0.215081f
C1223 two_stage_opamp_dummy_magic_25_0.V_source.t34 GNDA 0.033909f
C1224 two_stage_opamp_dummy_magic_25_0.V_source.t36 GNDA 0.033909f
C1225 two_stage_opamp_dummy_magic_25_0.V_source.n54 GNDA 0.072491f
C1226 two_stage_opamp_dummy_magic_25_0.V_source.n55 GNDA 0.260813f
C1227 two_stage_opamp_dummy_magic_25_0.V_source.t10 GNDA 0.033909f
C1228 two_stage_opamp_dummy_magic_25_0.V_source.t25 GNDA 0.033909f
C1229 two_stage_opamp_dummy_magic_25_0.V_source.n56 GNDA 0.072491f
C1230 two_stage_opamp_dummy_magic_25_0.V_source.n57 GNDA 0.260813f
C1231 two_stage_opamp_dummy_magic_25_0.V_source.t4 GNDA 0.033909f
C1232 two_stage_opamp_dummy_magic_25_0.V_source.t30 GNDA 0.033909f
C1233 two_stage_opamp_dummy_magic_25_0.V_source.n58 GNDA 0.072491f
C1234 two_stage_opamp_dummy_magic_25_0.V_source.n59 GNDA 0.260813f
C1235 two_stage_opamp_dummy_magic_25_0.V_source.n60 GNDA 0.104318f
C1236 two_stage_opamp_dummy_magic_25_0.V_source.n61 GNDA 0.178378f
C1237 two_stage_opamp_dummy_magic_25_0.X.n0 GNDA 0.069662f
C1238 two_stage_opamp_dummy_magic_25_0.X.n1 GNDA 0.102171f
C1239 two_stage_opamp_dummy_magic_25_0.X.n2 GNDA 0.2384f
C1240 two_stage_opamp_dummy_magic_25_0.X.n3 GNDA 0.162094f
C1241 two_stage_opamp_dummy_magic_25_0.X.n4 GNDA 0.272015f
C1242 two_stage_opamp_dummy_magic_25_0.X.t24 GNDA 0.023221f
C1243 two_stage_opamp_dummy_magic_25_0.X.t1 GNDA 0.023221f
C1244 two_stage_opamp_dummy_magic_25_0.X.n5 GNDA 0.050526f
C1245 two_stage_opamp_dummy_magic_25_0.X.n6 GNDA 0.161458f
C1246 two_stage_opamp_dummy_magic_25_0.X.n7 GNDA 0.046442f
C1247 two_stage_opamp_dummy_magic_25_0.X.n8 GNDA 0.088799f
C1248 two_stage_opamp_dummy_magic_25_0.X.t2 GNDA 0.023221f
C1249 two_stage_opamp_dummy_magic_25_0.X.t21 GNDA 0.023221f
C1250 two_stage_opamp_dummy_magic_25_0.X.n9 GNDA 0.050526f
C1251 two_stage_opamp_dummy_magic_25_0.X.n10 GNDA 0.161458f
C1252 two_stage_opamp_dummy_magic_25_0.X.n11 GNDA 0.16605f
C1253 two_stage_opamp_dummy_magic_25_0.X.n12 GNDA 0.102171f
C1254 two_stage_opamp_dummy_magic_25_0.X.n13 GNDA 0.102171f
C1255 two_stage_opamp_dummy_magic_25_0.X.n14 GNDA 0.074306f
C1256 two_stage_opamp_dummy_magic_25_0.X.t28 GNDA 0.049925f
C1257 two_stage_opamp_dummy_magic_25_0.X.t43 GNDA 0.056756f
C1258 two_stage_opamp_dummy_magic_25_0.X.n17 GNDA 0.046286f
C1259 two_stage_opamp_dummy_magic_25_0.X.t40 GNDA 0.049925f
C1260 two_stage_opamp_dummy_magic_25_0.X.t54 GNDA 0.049925f
C1261 two_stage_opamp_dummy_magic_25_0.X.t36 GNDA 0.049925f
C1262 two_stage_opamp_dummy_magic_25_0.X.t49 GNDA 0.049925f
C1263 two_stage_opamp_dummy_magic_25_0.X.t32 GNDA 0.049925f
C1264 two_stage_opamp_dummy_magic_25_0.X.t50 GNDA 0.049925f
C1265 two_stage_opamp_dummy_magic_25_0.X.t33 GNDA 0.049925f
C1266 two_stage_opamp_dummy_magic_25_0.X.t47 GNDA 0.056756f
C1267 two_stage_opamp_dummy_magic_25_0.X.n18 GNDA 0.051221f
C1268 two_stage_opamp_dummy_magic_25_0.X.n19 GNDA 0.031348f
C1269 two_stage_opamp_dummy_magic_25_0.X.n20 GNDA 0.031348f
C1270 two_stage_opamp_dummy_magic_25_0.X.n21 GNDA 0.031348f
C1271 two_stage_opamp_dummy_magic_25_0.X.n22 GNDA 0.031348f
C1272 two_stage_opamp_dummy_magic_25_0.X.n23 GNDA 0.031348f
C1273 two_stage_opamp_dummy_magic_25_0.X.n24 GNDA 0.026414f
C1274 two_stage_opamp_dummy_magic_25_0.X.n25 GNDA 0.012826f
C1275 two_stage_opamp_dummy_magic_25_0.X.t30 GNDA 0.032509f
C1276 two_stage_opamp_dummy_magic_25_0.X.t45 GNDA 0.039475f
C1277 two_stage_opamp_dummy_magic_25_0.X.n26 GNDA 0.034541f
C1278 two_stage_opamp_dummy_magic_25_0.X.t42 GNDA 0.032509f
C1279 two_stage_opamp_dummy_magic_25_0.X.t27 GNDA 0.032509f
C1280 two_stage_opamp_dummy_magic_25_0.X.t39 GNDA 0.032509f
C1281 two_stage_opamp_dummy_magic_25_0.X.t52 GNDA 0.032509f
C1282 two_stage_opamp_dummy_magic_25_0.X.t34 GNDA 0.032509f
C1283 two_stage_opamp_dummy_magic_25_0.X.t53 GNDA 0.032509f
C1284 two_stage_opamp_dummy_magic_25_0.X.t35 GNDA 0.032509f
C1285 two_stage_opamp_dummy_magic_25_0.X.t48 GNDA 0.039475f
C1286 two_stage_opamp_dummy_magic_25_0.X.n27 GNDA 0.039475f
C1287 two_stage_opamp_dummy_magic_25_0.X.n28 GNDA 0.025543f
C1288 two_stage_opamp_dummy_magic_25_0.X.n29 GNDA 0.025543f
C1289 two_stage_opamp_dummy_magic_25_0.X.n30 GNDA 0.025543f
C1290 two_stage_opamp_dummy_magic_25_0.X.n31 GNDA 0.025543f
C1291 two_stage_opamp_dummy_magic_25_0.X.n32 GNDA 0.025543f
C1292 two_stage_opamp_dummy_magic_25_0.X.n33 GNDA 0.020608f
C1293 two_stage_opamp_dummy_magic_25_0.X.n34 GNDA 0.012826f
C1294 two_stage_opamp_dummy_magic_25_0.X.n35 GNDA 0.080006f
C1295 two_stage_opamp_dummy_magic_25_0.X.n37 GNDA 0.074306f
C1296 two_stage_opamp_dummy_magic_25_0.X.t23 GNDA 0.642531f
C1297 two_stage_opamp_dummy_magic_25_0.X.n38 GNDA 0.074306f
C1298 two_stage_opamp_dummy_magic_25_0.X.n39 GNDA 0.074306f
C1299 two_stage_opamp_dummy_magic_25_0.X.n40 GNDA 0.073609f
C1300 two_stage_opamp_dummy_magic_25_0.X.n41 GNDA 0.689412f
C1301 two_stage_opamp_dummy_magic_25_0.X.n43 GNDA 0.645537f
C1302 two_stage_opamp_dummy_magic_25_0.X.n44 GNDA 0.024604f
C1303 two_stage_opamp_dummy_magic_25_0.X.n45 GNDA 0.024769f
C1304 two_stage_opamp_dummy_magic_25_0.X.n46 GNDA 0.024769f
C1305 two_stage_opamp_dummy_magic_25_0.X.t41 GNDA 0.102171f
C1306 two_stage_opamp_dummy_magic_25_0.X.t29 GNDA 0.102171f
C1307 two_stage_opamp_dummy_magic_25_0.X.t44 GNDA 0.102171f
C1308 two_stage_opamp_dummy_magic_25_0.X.t31 GNDA 0.102171f
C1309 two_stage_opamp_dummy_magic_25_0.X.t46 GNDA 0.108819f
C1310 two_stage_opamp_dummy_magic_25_0.X.n47 GNDA 0.086235f
C1311 two_stage_opamp_dummy_magic_25_0.X.n48 GNDA 0.048764f
C1312 two_stage_opamp_dummy_magic_25_0.X.n49 GNDA 0.048764f
C1313 two_stage_opamp_dummy_magic_25_0.X.n50 GNDA 0.043829f
C1314 two_stage_opamp_dummy_magic_25_0.X.t25 GNDA 0.102171f
C1315 two_stage_opamp_dummy_magic_25_0.X.t37 GNDA 0.102171f
C1316 two_stage_opamp_dummy_magic_25_0.X.t26 GNDA 0.102171f
C1317 two_stage_opamp_dummy_magic_25_0.X.t38 GNDA 0.102171f
C1318 two_stage_opamp_dummy_magic_25_0.X.t51 GNDA 0.108819f
C1319 two_stage_opamp_dummy_magic_25_0.X.n51 GNDA 0.086235f
C1320 two_stage_opamp_dummy_magic_25_0.X.n52 GNDA 0.048764f
C1321 two_stage_opamp_dummy_magic_25_0.X.n53 GNDA 0.048764f
C1322 two_stage_opamp_dummy_magic_25_0.X.n54 GNDA 0.043829f
C1323 two_stage_opamp_dummy_magic_25_0.X.n55 GNDA 0.010524f
C1324 two_stage_opamp_dummy_magic_25_0.X.n56 GNDA 0.024933f
C1325 two_stage_opamp_dummy_magic_25_0.X.n57 GNDA 0.058691f
C1326 two_stage_opamp_dummy_magic_25_0.X.n58 GNDA 0.033474f
C1327 two_stage_opamp_dummy_magic_25_0.X.n59 GNDA 0.037989f
C1328 two_stage_opamp_dummy_magic_25_0.X.n60 GNDA 1.02636f
C1329 two_stage_opamp_dummy_magic_25_0.X.n61 GNDA 0.074306f
C1330 two_stage_opamp_dummy_magic_25_0.X.n63 GNDA 0.074306f
C1331 two_stage_opamp_dummy_magic_25_0.X.n64 GNDA 0.074306f
C1332 two_stage_opamp_dummy_magic_25_0.X.n65 GNDA 0.100296f
C1333 two_stage_opamp_dummy_magic_25_0.X.n66 GNDA 0.120748f
C1334 two_stage_opamp_dummy_magic_25_0.X.n67 GNDA 0.074306f
C1335 two_stage_opamp_dummy_magic_25_0.X.n68 GNDA 0.095765f
C1336 two_stage_opamp_dummy_magic_25_0.X.n69 GNDA 0.074306f
C1337 two_stage_opamp_dummy_magic_25_0.X.n70 GNDA 0.074306f
C1338 two_stage_opamp_dummy_magic_25_0.X.n71 GNDA 0.095765f
C1339 two_stage_opamp_dummy_magic_25_0.X.n72 GNDA 0.074306f
C1340 two_stage_opamp_dummy_magic_25_0.X.n73 GNDA 0.122441f
C1341 two_stage_opamp_dummy_magic_25_0.X.t9 GNDA 0.054182f
C1342 two_stage_opamp_dummy_magic_25_0.X.t11 GNDA 0.054182f
C1343 two_stage_opamp_dummy_magic_25_0.X.n74 GNDA 0.110834f
C1344 two_stage_opamp_dummy_magic_25_0.X.n75 GNDA 0.296573f
C1345 two_stage_opamp_dummy_magic_25_0.X.t4 GNDA 0.054182f
C1346 two_stage_opamp_dummy_magic_25_0.X.t12 GNDA 0.054182f
C1347 two_stage_opamp_dummy_magic_25_0.X.n76 GNDA 0.110834f
C1348 two_stage_opamp_dummy_magic_25_0.X.n77 GNDA 0.301473f
C1349 two_stage_opamp_dummy_magic_25_0.X.t14 GNDA 0.054182f
C1350 two_stage_opamp_dummy_magic_25_0.X.t3 GNDA 0.054182f
C1351 two_stage_opamp_dummy_magic_25_0.X.n78 GNDA 0.110834f
C1352 two_stage_opamp_dummy_magic_25_0.X.n79 GNDA 0.301473f
C1353 two_stage_opamp_dummy_magic_25_0.X.n80 GNDA 0.100255f
C1354 two_stage_opamp_dummy_magic_25_0.X.t8 GNDA 0.054182f
C1355 two_stage_opamp_dummy_magic_25_0.X.t10 GNDA 0.054182f
C1356 two_stage_opamp_dummy_magic_25_0.X.n81 GNDA 0.110834f
C1357 two_stage_opamp_dummy_magic_25_0.X.n82 GNDA 0.296573f
C1358 two_stage_opamp_dummy_magic_25_0.X.n83 GNDA 0.05877f
C1359 two_stage_opamp_dummy_magic_25_0.X.t6 GNDA 0.054182f
C1360 two_stage_opamp_dummy_magic_25_0.X.t7 GNDA 0.054182f
C1361 two_stage_opamp_dummy_magic_25_0.X.n84 GNDA 0.110834f
C1362 two_stage_opamp_dummy_magic_25_0.X.n85 GNDA 0.296573f
C1363 two_stage_opamp_dummy_magic_25_0.X.n86 GNDA 0.05877f
C1364 two_stage_opamp_dummy_magic_25_0.X.n87 GNDA 0.100255f
C1365 two_stage_opamp_dummy_magic_25_0.X.t15 GNDA 0.054182f
C1366 two_stage_opamp_dummy_magic_25_0.X.t13 GNDA 0.054182f
C1367 two_stage_opamp_dummy_magic_25_0.X.n88 GNDA 0.110834f
C1368 two_stage_opamp_dummy_magic_25_0.X.n89 GNDA 0.296573f
C1369 two_stage_opamp_dummy_magic_25_0.X.n90 GNDA 0.095765f
C1370 two_stage_opamp_dummy_magic_25_0.X.n91 GNDA 0.08216f
C1371 two_stage_opamp_dummy_magic_25_0.X.n92 GNDA 0.049538f
C1372 two_stage_opamp_dummy_magic_25_0.X.n93 GNDA 0.049538f
C1373 two_stage_opamp_dummy_magic_25_0.X.n94 GNDA 0.08216f
C1374 two_stage_opamp_dummy_magic_25_0.X.n95 GNDA 0.095765f
C1375 two_stage_opamp_dummy_magic_25_0.X.n96 GNDA 0.16942f
C1376 two_stage_opamp_dummy_magic_25_0.X.n97 GNDA 0.25095f
C1377 two_stage_opamp_dummy_magic_25_0.X.n98 GNDA 0.319127f
C1378 two_stage_opamp_dummy_magic_25_0.X.n99 GNDA 0.074306f
C1379 two_stage_opamp_dummy_magic_25_0.X.n100 GNDA 0.074306f
C1380 two_stage_opamp_dummy_magic_25_0.X.n101 GNDA 0.120748f
C1381 two_stage_opamp_dummy_magic_25_0.X.n102 GNDA 0.074306f
C1382 two_stage_opamp_dummy_magic_25_0.X.n103 GNDA 0.074306f
C1383 two_stage_opamp_dummy_magic_25_0.X.n104 GNDA 0.074306f
C1384 two_stage_opamp_dummy_magic_25_0.X.n105 GNDA 0.074306f
C1385 two_stage_opamp_dummy_magic_25_0.X.n106 GNDA 0.120748f
C1386 two_stage_opamp_dummy_magic_25_0.X.n107 GNDA 0.074306f
C1387 two_stage_opamp_dummy_magic_25_0.X.n108 GNDA 0.074306f
C1388 two_stage_opamp_dummy_magic_25_0.X.n109 GNDA 0.074306f
C1389 two_stage_opamp_dummy_magic_25_0.X.n110 GNDA 0.074306f
C1390 two_stage_opamp_dummy_magic_25_0.X.n111 GNDA 0.074306f
C1391 two_stage_opamp_dummy_magic_25_0.X.n112 GNDA 0.074306f
C1392 two_stage_opamp_dummy_magic_25_0.X.n113 GNDA 0.074306f
C1393 two_stage_opamp_dummy_magic_25_0.X.n114 GNDA 0.120748f
C1394 two_stage_opamp_dummy_magic_25_0.X.n115 GNDA 0.580519f
C1395 two_stage_opamp_dummy_magic_25_0.X.n116 GNDA 0.580519f
C1396 two_stage_opamp_dummy_magic_25_0.X.n117 GNDA 0.073609f
C1397 two_stage_opamp_dummy_magic_25_0.X.n118 GNDA 0.074306f
C1398 two_stage_opamp_dummy_magic_25_0.X.n119 GNDA 0.074306f
C1399 two_stage_opamp_dummy_magic_25_0.X.n121 GNDA 0.910253f
C1400 two_stage_opamp_dummy_magic_25_0.X.n122 GNDA 0.910253f
C1401 two_stage_opamp_dummy_magic_25_0.X.n124 GNDA 0.455127f
C1402 two_stage_opamp_dummy_magic_25_0.X.n125 GNDA 2.1959f
C1403 two_stage_opamp_dummy_magic_25_0.X.n126 GNDA 0.599095f
C1404 two_stage_opamp_dummy_magic_25_0.X.n127 GNDA 0.224467f
C1405 two_stage_opamp_dummy_magic_25_0.X.n128 GNDA 0.613028f
C1406 two_stage_opamp_dummy_magic_25_0.X.n129 GNDA 0.102171f
C1407 two_stage_opamp_dummy_magic_25_0.X.n130 GNDA 0.102171f
C1408 two_stage_opamp_dummy_magic_25_0.X.n131 GNDA 0.102171f
C1409 two_stage_opamp_dummy_magic_25_0.X.n132 GNDA 0.2384f
C1410 two_stage_opamp_dummy_magic_25_0.X.t18 GNDA 0.023221f
C1411 two_stage_opamp_dummy_magic_25_0.X.t0 GNDA 0.023221f
C1412 two_stage_opamp_dummy_magic_25_0.X.n133 GNDA 0.050526f
C1413 two_stage_opamp_dummy_magic_25_0.X.n134 GNDA 0.157355f
C1414 two_stage_opamp_dummy_magic_25_0.X.n135 GNDA 0.162094f
C1415 two_stage_opamp_dummy_magic_25_0.X.n136 GNDA 0.078091f
C1416 two_stage_opamp_dummy_magic_25_0.X.n137 GNDA 0.046442f
C1417 two_stage_opamp_dummy_magic_25_0.X.n138 GNDA 0.162094f
C1418 two_stage_opamp_dummy_magic_25_0.X.t22 GNDA 0.023221f
C1419 two_stage_opamp_dummy_magic_25_0.X.t16 GNDA 0.023221f
C1420 two_stage_opamp_dummy_magic_25_0.X.n139 GNDA 0.050526f
C1421 two_stage_opamp_dummy_magic_25_0.X.n140 GNDA 0.157355f
C1422 two_stage_opamp_dummy_magic_25_0.X.n141 GNDA 0.051869f
C1423 two_stage_opamp_dummy_magic_25_0.X.t19 GNDA 0.023221f
C1424 two_stage_opamp_dummy_magic_25_0.X.t17 GNDA 0.023221f
C1425 two_stage_opamp_dummy_magic_25_0.X.n142 GNDA 0.050526f
C1426 two_stage_opamp_dummy_magic_25_0.X.n143 GNDA 0.157355f
C1427 two_stage_opamp_dummy_magic_25_0.X.n144 GNDA 0.051869f
C1428 two_stage_opamp_dummy_magic_25_0.X.n145 GNDA 0.088799f
C1429 two_stage_opamp_dummy_magic_25_0.X.t20 GNDA 0.023221f
C1430 two_stage_opamp_dummy_magic_25_0.X.t5 GNDA 0.023221f
C1431 two_stage_opamp_dummy_magic_25_0.X.n146 GNDA 0.050526f
C1432 two_stage_opamp_dummy_magic_25_0.X.n147 GNDA 0.157355f
C1433 two_stage_opamp_dummy_magic_25_0.X.n148 GNDA 0.162094f
C1434 two_stage_opamp_dummy_magic_25_0.X.n149 GNDA 0.078091f
C1435 two_stage_opamp_dummy_magic_25_0.X.n150 GNDA 0.177011f
C1436 two_stage_opamp_dummy_magic_25_0.X.n151 GNDA 0.32662f
C1437 two_stage_opamp_dummy_magic_25_0.X.n152 GNDA 0.350195f
C1438 two_stage_opamp_dummy_magic_25_0.X.n153 GNDA 0.102171f
C1439 two_stage_opamp_dummy_magic_25_0.X.n154 GNDA 0.2384f
C1440 two_stage_opamp_dummy_magic_25_0.X.n155 GNDA 0.102171f
C1441 two_stage_opamp_dummy_magic_25_0.X.n156 GNDA 0.083595f
C1442 two_stage_opamp_dummy_magic_25_0.Vb2.t7 GNDA 0.063923f
C1443 two_stage_opamp_dummy_magic_25_0.Vb2.t8 GNDA 0.018264f
C1444 two_stage_opamp_dummy_magic_25_0.Vb2.t5 GNDA 0.018264f
C1445 two_stage_opamp_dummy_magic_25_0.Vb2.n0 GNDA 0.061236f
C1446 two_stage_opamp_dummy_magic_25_0.Vb2.t1 GNDA 0.018264f
C1447 two_stage_opamp_dummy_magic_25_0.Vb2.t0 GNDA 0.018264f
C1448 two_stage_opamp_dummy_magic_25_0.Vb2.n1 GNDA 0.059556f
C1449 two_stage_opamp_dummy_magic_25_0.Vb2.n2 GNDA 0.54401f
C1450 two_stage_opamp_dummy_magic_25_0.Vb2.t10 GNDA 0.018264f
C1451 two_stage_opamp_dummy_magic_25_0.Vb2.t9 GNDA 0.018264f
C1452 two_stage_opamp_dummy_magic_25_0.Vb2.n3 GNDA 0.059556f
C1453 two_stage_opamp_dummy_magic_25_0.Vb2.n4 GNDA 0.356858f
C1454 two_stage_opamp_dummy_magic_25_0.Vb2.t6 GNDA 0.018264f
C1455 two_stage_opamp_dummy_magic_25_0.Vb2.t2 GNDA 0.018264f
C1456 two_stage_opamp_dummy_magic_25_0.Vb2.n5 GNDA 0.059556f
C1457 two_stage_opamp_dummy_magic_25_0.Vb2.n6 GNDA 2.3034f
C1458 two_stage_opamp_dummy_magic_25_0.Vb2.t22 GNDA 0.117487f
C1459 two_stage_opamp_dummy_magic_25_0.Vb2.n7 GNDA 2.10471f
C1460 two_stage_opamp_dummy_magic_25_0.Vb2.t25 GNDA 0.090406f
C1461 two_stage_opamp_dummy_magic_25_0.Vb2.t19 GNDA 0.090406f
C1462 two_stage_opamp_dummy_magic_25_0.Vb2.t23 GNDA 0.090406f
C1463 two_stage_opamp_dummy_magic_25_0.Vb2.t17 GNDA 0.090406f
C1464 two_stage_opamp_dummy_magic_25_0.Vb2.t12 GNDA 0.104328f
C1465 two_stage_opamp_dummy_magic_25_0.Vb2.n8 GNDA 0.084703f
C1466 two_stage_opamp_dummy_magic_25_0.Vb2.n9 GNDA 0.052052f
C1467 two_stage_opamp_dummy_magic_25_0.Vb2.n10 GNDA 0.052052f
C1468 two_stage_opamp_dummy_magic_25_0.Vb2.n11 GNDA 0.045639f
C1469 two_stage_opamp_dummy_magic_25_0.Vb2.t29 GNDA 0.090406f
C1470 two_stage_opamp_dummy_magic_25_0.Vb2.t32 GNDA 0.090406f
C1471 two_stage_opamp_dummy_magic_25_0.Vb2.t13 GNDA 0.090406f
C1472 two_stage_opamp_dummy_magic_25_0.Vb2.t11 GNDA 0.090406f
C1473 two_stage_opamp_dummy_magic_25_0.Vb2.t15 GNDA 0.104328f
C1474 two_stage_opamp_dummy_magic_25_0.Vb2.n12 GNDA 0.084703f
C1475 two_stage_opamp_dummy_magic_25_0.Vb2.n13 GNDA 0.052052f
C1476 two_stage_opamp_dummy_magic_25_0.Vb2.n14 GNDA 0.052052f
C1477 two_stage_opamp_dummy_magic_25_0.Vb2.n15 GNDA 0.045639f
C1478 two_stage_opamp_dummy_magic_25_0.Vb2.n16 GNDA 0.033825f
C1479 two_stage_opamp_dummy_magic_25_0.Vb2.t28 GNDA 0.090406f
C1480 two_stage_opamp_dummy_magic_25_0.Vb2.t26 GNDA 0.090406f
C1481 two_stage_opamp_dummy_magic_25_0.Vb2.t21 GNDA 0.090406f
C1482 two_stage_opamp_dummy_magic_25_0.Vb2.t16 GNDA 0.090406f
C1483 two_stage_opamp_dummy_magic_25_0.Vb2.t20 GNDA 0.104328f
C1484 two_stage_opamp_dummy_magic_25_0.Vb2.n17 GNDA 0.084703f
C1485 two_stage_opamp_dummy_magic_25_0.Vb2.n18 GNDA 0.052052f
C1486 two_stage_opamp_dummy_magic_25_0.Vb2.n19 GNDA 0.052052f
C1487 two_stage_opamp_dummy_magic_25_0.Vb2.n20 GNDA 0.045639f
C1488 two_stage_opamp_dummy_magic_25_0.Vb2.t30 GNDA 0.090406f
C1489 two_stage_opamp_dummy_magic_25_0.Vb2.t14 GNDA 0.090406f
C1490 two_stage_opamp_dummy_magic_25_0.Vb2.t18 GNDA 0.090406f
C1491 two_stage_opamp_dummy_magic_25_0.Vb2.t24 GNDA 0.090406f
C1492 two_stage_opamp_dummy_magic_25_0.Vb2.t27 GNDA 0.104328f
C1493 two_stage_opamp_dummy_magic_25_0.Vb2.n21 GNDA 0.084703f
C1494 two_stage_opamp_dummy_magic_25_0.Vb2.n22 GNDA 0.052052f
C1495 two_stage_opamp_dummy_magic_25_0.Vb2.n23 GNDA 0.052052f
C1496 two_stage_opamp_dummy_magic_25_0.Vb2.n24 GNDA 0.045639f
C1497 two_stage_opamp_dummy_magic_25_0.Vb2.n25 GNDA 0.033328f
C1498 two_stage_opamp_dummy_magic_25_0.Vb2.n26 GNDA 0.762106f
C1499 two_stage_opamp_dummy_magic_25_0.Vb2.n27 GNDA 0.374426f
C1500 two_stage_opamp_dummy_magic_25_0.Vb2.t31 GNDA 0.071661f
C1501 two_stage_opamp_dummy_magic_25_0.Vb2.n28 GNDA 0.27511f
C1502 two_stage_opamp_dummy_magic_25_0.Vb2.t3 GNDA 0.119327f
C1503 two_stage_opamp_dummy_magic_25_0.Vb2.n29 GNDA 0.552559f
C1504 two_stage_opamp_dummy_magic_25_0.Vb2.n30 GNDA 0.135746f
C1505 two_stage_opamp_dummy_magic_25_0.Vb2.t4 GNDA 0.063923f
C1506 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t43 GNDA 0.412258f
C1507 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t85 GNDA 0.434383f
C1508 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t61 GNDA 0.413752f
C1509 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t66 GNDA 0.412258f
C1510 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t100 GNDA 0.221432f
C1511 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n0 GNDA 0.255706f
C1512 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t89 GNDA 0.412258f
C1513 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t102 GNDA 0.434383f
C1514 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t1 GNDA 0.221432f
C1515 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n1 GNDA 0.235076f
C1516 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t131 GNDA 0.412258f
C1517 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t6 GNDA 0.434383f
C1518 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t36 GNDA 0.221432f
C1519 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n2 GNDA 0.235076f
C1520 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t34 GNDA 0.412258f
C1521 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t128 GNDA 0.434383f
C1522 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t17 GNDA 0.221432f
C1523 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n3 GNDA 0.235076f
C1524 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t13 GNDA 0.412258f
C1525 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t80 GNDA 0.413752f
C1526 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t33 GNDA 0.412258f
C1527 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t74 GNDA 0.413752f
C1528 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t124 GNDA 0.412258f
C1529 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t40 GNDA 0.413752f
C1530 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t18 GNDA 0.412258f
C1531 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t47 GNDA 0.413752f
C1532 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t130 GNDA 0.412258f
C1533 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t76 GNDA 0.413752f
C1534 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t51 GNDA 0.412258f
C1535 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t91 GNDA 0.413752f
C1536 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t25 GNDA 0.412258f
C1537 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t120 GNDA 0.413752f
C1538 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t24 GNDA 0.412258f
C1539 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t53 GNDA 0.413752f
C1540 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t136 GNDA 0.412258f
C1541 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t81 GNDA 0.413752f
C1542 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t59 GNDA 0.412258f
C1543 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t96 GNDA 0.413752f
C1544 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t31 GNDA 0.412258f
C1545 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t126 GNDA 0.413752f
C1546 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t98 GNDA 0.412258f
C1547 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t138 GNDA 0.413752f
C1548 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t67 GNDA 0.412258f
C1549 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t22 GNDA 0.413752f
C1550 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t65 GNDA 0.412258f
C1551 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t99 GNDA 0.413752f
C1552 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t32 GNDA 0.412258f
C1553 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t132 GNDA 0.413752f
C1554 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t108 GNDA 0.412258f
C1555 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t5 GNDA 0.413752f
C1556 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t75 GNDA 0.412258f
C1557 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t29 GNDA 0.413752f
C1558 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t8 GNDA 0.412258f
C1559 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t39 GNDA 0.413752f
C1560 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t118 GNDA 0.412258f
C1561 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t62 GNDA 0.413752f
C1562 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t41 GNDA 0.412258f
C1563 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t83 GNDA 0.413752f
C1564 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t14 GNDA 0.412258f
C1565 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t103 GNDA 0.413752f
C1566 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t12 GNDA 0.412258f
C1567 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t42 GNDA 0.413752f
C1568 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t125 GNDA 0.412258f
C1569 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t70 GNDA 0.413752f
C1570 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t46 GNDA 0.412258f
C1571 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t86 GNDA 0.413752f
C1572 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t20 GNDA 0.412258f
C1573 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t113 GNDA 0.413752f
C1574 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t90 GNDA 0.412258f
C1575 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t134 GNDA 0.413752f
C1576 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t56 GNDA 0.412258f
C1577 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t10 GNDA 0.413752f
C1578 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t52 GNDA 0.412258f
C1579 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t92 GNDA 0.413752f
C1580 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t26 GNDA 0.412258f
C1581 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t121 GNDA 0.413752f
C1582 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t116 GNDA 0.412258f
C1583 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t60 GNDA 0.413752f
C1584 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t109 GNDA 0.412258f
C1585 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t44 GNDA 0.413752f
C1586 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t106 GNDA 0.412258f
C1587 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t3 GNDA 0.413752f
C1588 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t73 GNDA 0.412258f
C1589 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t27 GNDA 0.413752f
C1590 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t2 GNDA 0.412258f
C1591 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t35 GNDA 0.413752f
C1592 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t110 GNDA 0.412258f
C1593 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t57 GNDA 0.413752f
C1594 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t45 GNDA 0.412258f
C1595 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t88 GNDA 0.432471f
C1596 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t87 GNDA 0.412258f
C1597 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t135 GNDA 0.221432f
C1598 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n4 GNDA 0.236987f
C1599 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t63 GNDA 0.412258f
C1600 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t104 GNDA 0.221432f
C1601 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n5 GNDA 0.235076f
C1602 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t101 GNDA 0.412258f
C1603 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t7 GNDA 0.221432f
C1604 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n6 GNDA 0.235076f
C1605 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t4 GNDA 0.412258f
C1606 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t38 GNDA 0.221432f
C1607 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n7 GNDA 0.235076f
C1608 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t37 GNDA 0.412258f
C1609 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t79 GNDA 0.221432f
C1610 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n8 GNDA 0.235076f
C1611 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t19 GNDA 0.412258f
C1612 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t55 GNDA 0.221432f
C1613 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n9 GNDA 0.235076f
C1614 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t50 GNDA 0.412258f
C1615 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t95 GNDA 0.221432f
C1616 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n10 GNDA 0.235076f
C1617 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t94 GNDA 0.412258f
C1618 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t137 GNDA 0.221432f
C1619 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n11 GNDA 0.235076f
C1620 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t72 GNDA 0.412258f
C1621 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t115 GNDA 0.221432f
C1622 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n12 GNDA 0.235076f
C1623 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t112 GNDA 0.412258f
C1624 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t9 GNDA 0.221432f
C1625 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n13 GNDA 0.235076f
C1626 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t48 GNDA 0.412258f
C1627 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t129 GNDA 0.413752f
C1628 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t15 GNDA 0.412258f
C1629 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t84 GNDA 0.413752f
C1630 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t119 GNDA 0.199307f
C1631 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n14 GNDA 0.257077f
C1632 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t16 GNDA 0.220062f
C1633 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n15 GNDA 0.279201f
C1634 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t58 GNDA 0.220062f
C1635 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n16 GNDA 0.299832f
C1636 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t28 GNDA 0.220062f
C1637 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n17 GNDA 0.299832f
C1638 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t97 GNDA 0.220062f
C1639 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n18 GNDA 0.299832f
C1640 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t123 GNDA 0.220062f
C1641 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n19 GNDA 0.299832f
C1642 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t11 GNDA 0.220062f
C1643 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n20 GNDA 0.299832f
C1644 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t114 GNDA 0.220062f
C1645 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n21 GNDA 0.299832f
C1646 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t71 GNDA 0.220062f
C1647 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n22 GNDA 0.299832f
C1648 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t107 GNDA 0.220062f
C1649 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n23 GNDA 0.299832f
C1650 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t64 GNDA 0.220062f
C1651 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n24 GNDA 0.299832f
C1652 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t30 GNDA 0.220062f
C1653 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n25 GNDA 0.299832f
C1654 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t133 GNDA 0.220062f
C1655 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n26 GNDA 0.299832f
C1656 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t23 GNDA 0.220062f
C1657 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n27 GNDA 0.299832f
C1658 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t127 GNDA 0.220062f
C1659 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n28 GNDA 0.299832f
C1660 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t82 GNDA 0.220062f
C1661 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n29 GNDA 0.299832f
C1662 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t122 GNDA 0.220062f
C1663 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n30 GNDA 0.299832f
C1664 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t77 GNDA 0.220062f
C1665 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n31 GNDA 0.299832f
C1666 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t78 GNDA 0.220062f
C1667 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n32 GNDA 0.299832f
C1668 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t117 GNDA 0.220062f
C1669 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n33 GNDA 0.276337f
C1670 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t111 GNDA 0.413752f
C1671 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t68 GNDA 0.413752f
C1672 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t105 GNDA 0.412258f
C1673 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t54 GNDA 0.434383f
C1674 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t93 GNDA 0.221432f
C1675 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n34 GNDA 0.255706f
C1676 two_stage_opamp_dummy_magic_25_0.cap_res_Y.n35 GNDA 0.235076f
C1677 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t49 GNDA 0.221432f
C1678 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t21 GNDA 0.434383f
C1679 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t69 GNDA 0.590705f
C1680 two_stage_opamp_dummy_magic_25_0.cap_res_Y.t0 GNDA 0.355571f
C1681 VOUT+.n0 GNDA 0.036192f
C1682 VOUT+.t12 GNDA 0.05278f
C1683 VOUT+.t9 GNDA 0.05278f
C1684 VOUT+.n1 GNDA 0.113404f
C1685 VOUT+.n2 GNDA 0.272735f
C1686 VOUT+.n3 GNDA 0.036192f
C1687 VOUT+.n4 GNDA 0.23372f
C1688 VOUT+.t4 GNDA 0.05278f
C1689 VOUT+.t3 GNDA 0.05278f
C1690 VOUT+.n5 GNDA 0.113404f
C1691 VOUT+.n6 GNDA 0.282262f
C1692 VOUT+.n7 GNDA 0.161339f
C1693 VOUT+.t0 GNDA 0.05278f
C1694 VOUT+.t10 GNDA 0.05278f
C1695 VOUT+.n8 GNDA 0.113404f
C1696 VOUT+.n9 GNDA 0.268146f
C1697 VOUT+.n10 GNDA 0.12306f
C1698 VOUT+.n11 GNDA 0.036192f
C1699 VOUT+.n12 GNDA 0.186755f
C1700 VOUT+.n13 GNDA 0.036192f
C1701 VOUT+.n14 GNDA 0.036192f
C1702 VOUT+.n15 GNDA 0.036192f
C1703 VOUT+.n16 GNDA 0.036192f
C1704 VOUT+.n17 GNDA 0.077474f
C1705 VOUT+.n18 GNDA 0.183223f
C1706 VOUT+.t1 GNDA 0.086088f
C1707 VOUT+.n19 GNDA 0.263015f
C1708 VOUT+.n20 GNDA 0.0754f
C1709 VOUT+.n23 GNDA 0.038454f
C1710 VOUT+.n25 GNDA 0.038454f
C1711 VOUT+.n28 GNDA 0.05655f
C1712 VOUT+.n29 GNDA 0.09425f
C1713 VOUT+.n30 GNDA 0.059913f
C1714 VOUT+.n31 GNDA 0.05655f
C1715 VOUT+.n33 GNDA 0.038454f
C1716 VOUT+.n34 GNDA 0.035853f
C1717 VOUT+.n35 GNDA 0.038454f
C1718 VOUT+.n36 GNDA 0.049764f
C1719 VOUT+.n37 GNDA 0.071798f
C1720 VOUT+.n38 GNDA 0.069871f
C1721 VOUT+.n39 GNDA 0.049764f
C1722 VOUT+.n40 GNDA 0.049764f
C1723 VOUT+.n41 GNDA 0.069871f
C1724 VOUT+.n42 GNDA 0.069871f
C1725 VOUT+.n43 GNDA 0.049764f
C1726 VOUT+.n44 GNDA 0.079669f
C1727 VOUT+.t14 GNDA 0.04524f
C1728 VOUT+.t18 GNDA 0.04524f
C1729 VOUT+.n45 GNDA 0.092697f
C1730 VOUT+.n46 GNDA 0.239278f
C1731 VOUT+.t5 GNDA 0.04524f
C1732 VOUT+.t15 GNDA 0.04524f
C1733 VOUT+.n47 GNDA 0.092697f
C1734 VOUT+.n48 GNDA 0.239278f
C1735 VOUT+.t11 GNDA 0.04524f
C1736 VOUT+.t17 GNDA 0.04524f
C1737 VOUT+.n49 GNDA 0.092697f
C1738 VOUT+.n50 GNDA 0.236867f
C1739 VOUT+.n51 GNDA 0.057528f
C1740 VOUT+.t16 GNDA 0.04524f
C1741 VOUT+.t8 GNDA 0.04524f
C1742 VOUT+.n52 GNDA 0.092697f
C1743 VOUT+.n53 GNDA 0.236867f
C1744 VOUT+.n54 GNDA 0.032609f
C1745 VOUT+.t13 GNDA 0.04524f
C1746 VOUT+.t2 GNDA 0.04524f
C1747 VOUT+.n55 GNDA 0.092697f
C1748 VOUT+.n56 GNDA 0.236867f
C1749 VOUT+.n57 GNDA 0.032609f
C1750 VOUT+.n58 GNDA 0.057528f
C1751 VOUT+.t7 GNDA 0.04524f
C1752 VOUT+.t6 GNDA 0.04524f
C1753 VOUT+.n59 GNDA 0.092697f
C1754 VOUT+.n60 GNDA 0.236867f
C1755 VOUT+.n61 GNDA 0.038035f
C1756 VOUT+.n62 GNDA 0.02262f
C1757 VOUT+.n63 GNDA 0.02262f
C1758 VOUT+.n64 GNDA 0.038035f
C1759 VOUT+.n65 GNDA 0.069871f
C1760 VOUT+.n66 GNDA 0.097805f
C1761 VOUT+.n67 GNDA 0.12187f
C1762 VOUT+.n68 GNDA 0.170568f
C1763 VOUT+.n69 GNDA 0.049764f
C1764 VOUT+.n70 GNDA 0.081432f
C1765 VOUT+.n71 GNDA 0.049764f
C1766 VOUT+.n72 GNDA 0.081432f
C1767 VOUT+.n73 GNDA 0.049764f
C1768 VOUT+.n74 GNDA 0.049764f
C1769 VOUT+.n75 GNDA 0.049764f
C1770 VOUT+.n76 GNDA 0.081432f
C1771 VOUT+.n77 GNDA 0.049764f
C1772 VOUT+.n78 GNDA 0.074646f
C1773 VOUT+.n79 GNDA 0.239773f
C1774 VOUT+.n81 GNDA 0.0754f
C1775 VOUT+.n82 GNDA 0.038454f
C1776 VOUT+.n84 GNDA 0.038454f
C1777 VOUT+.n87 GNDA 0.0754f
C1778 VOUT+.n88 GNDA 0.232987f
C1779 VOUT+.n89 GNDA 0.537227f
C1780 VOUT+.n92 GNDA 0.05655f
C1781 VOUT+.n93 GNDA 0.05655f
C1782 VOUT+.n94 GNDA 0.05655f
C1783 VOUT+.n95 GNDA 0.05655f
C1784 VOUT+.n96 GNDA 0.165871f
C1785 VOUT+.n97 GNDA 0.05655f
C1786 VOUT+.t38 GNDA 0.301601f
C1787 VOUT+.t142 GNDA 0.306738f
C1788 VOUT+.t73 GNDA 0.301601f
C1789 VOUT+.n98 GNDA 0.202214f
C1790 VOUT+.n99 GNDA 0.13195f
C1791 VOUT+.t45 GNDA 0.306095f
C1792 VOUT+.t85 GNDA 0.306095f
C1793 VOUT+.t63 GNDA 0.306095f
C1794 VOUT+.t107 GNDA 0.306095f
C1795 VOUT+.t138 GNDA 0.306095f
C1796 VOUT+.t120 GNDA 0.306095f
C1797 VOUT+.t153 GNDA 0.306095f
C1798 VOUT+.t56 GNDA 0.306095f
C1799 VOUT+.t94 GNDA 0.306095f
C1800 VOUT+.t70 GNDA 0.306095f
C1801 VOUT+.t112 GNDA 0.306095f
C1802 VOUT+.t69 GNDA 0.301601f
C1803 VOUT+.n100 GNDA 0.202857f
C1804 VOUT+.t22 GNDA 0.301601f
C1805 VOUT+.n101 GNDA 0.259407f
C1806 VOUT+.t53 GNDA 0.301601f
C1807 VOUT+.n102 GNDA 0.259407f
C1808 VOUT+.t150 GNDA 0.301601f
C1809 VOUT+.n103 GNDA 0.259407f
C1810 VOUT+.t119 GNDA 0.301601f
C1811 VOUT+.n104 GNDA 0.259407f
C1812 VOUT+.t78 GNDA 0.301601f
C1813 VOUT+.n105 GNDA 0.259407f
C1814 VOUT+.t102 GNDA 0.301601f
C1815 VOUT+.n106 GNDA 0.259407f
C1816 VOUT+.t62 GNDA 0.301601f
C1817 VOUT+.n107 GNDA 0.259407f
C1818 VOUT+.t20 GNDA 0.301601f
C1819 VOUT+.n108 GNDA 0.259407f
C1820 VOUT+.t42 GNDA 0.301601f
C1821 VOUT+.n109 GNDA 0.259407f
C1822 VOUT+.t148 GNDA 0.301601f
C1823 VOUT+.n110 GNDA 0.259407f
C1824 VOUT+.t141 GNDA 0.301601f
C1825 VOUT+.t109 GNDA 0.306738f
C1826 VOUT+.t28 GNDA 0.301601f
C1827 VOUT+.n111 GNDA 0.202214f
C1828 VOUT+.n112 GNDA 0.245051f
C1829 VOUT+.t155 GNDA 0.306738f
C1830 VOUT+.t122 GNDA 0.301601f
C1831 VOUT+.n113 GNDA 0.202214f
C1832 VOUT+.t99 GNDA 0.301601f
C1833 VOUT+.t47 GNDA 0.306738f
C1834 VOUT+.t100 GNDA 0.301601f
C1835 VOUT+.n114 GNDA 0.202214f
C1836 VOUT+.n115 GNDA 0.245051f
C1837 VOUT+.t51 GNDA 0.306738f
C1838 VOUT+.t154 GNDA 0.301601f
C1839 VOUT+.n116 GNDA 0.202214f
C1840 VOUT+.t129 GNDA 0.301601f
C1841 VOUT+.t84 GNDA 0.306738f
C1842 VOUT+.t130 GNDA 0.301601f
C1843 VOUT+.n117 GNDA 0.202214f
C1844 VOUT+.n118 GNDA 0.245051f
C1845 VOUT+.t41 GNDA 0.306738f
C1846 VOUT+.t97 GNDA 0.301601f
C1847 VOUT+.n119 GNDA 0.202214f
C1848 VOUT+.t60 GNDA 0.301601f
C1849 VOUT+.t48 GNDA 0.306738f
C1850 VOUT+.t113 GNDA 0.301601f
C1851 VOUT+.n120 GNDA 0.202214f
C1852 VOUT+.n121 GNDA 0.245051f
C1853 VOUT+.t105 GNDA 0.306738f
C1854 VOUT+.t65 GNDA 0.301601f
C1855 VOUT+.n122 GNDA 0.202214f
C1856 VOUT+.t34 GNDA 0.301601f
C1857 VOUT+.t131 GNDA 0.306738f
C1858 VOUT+.t36 GNDA 0.301601f
C1859 VOUT+.n123 GNDA 0.202214f
C1860 VOUT+.n124 GNDA 0.245051f
C1861 VOUT+.t67 GNDA 0.306738f
C1862 VOUT+.t23 GNDA 0.301601f
C1863 VOUT+.n125 GNDA 0.202214f
C1864 VOUT+.t146 GNDA 0.301601f
C1865 VOUT+.t101 GNDA 0.306738f
C1866 VOUT+.t147 GNDA 0.301601f
C1867 VOUT+.n126 GNDA 0.202214f
C1868 VOUT+.n127 GNDA 0.245051f
C1869 VOUT+.t111 GNDA 0.306738f
C1870 VOUT+.t71 GNDA 0.301601f
C1871 VOUT+.n128 GNDA 0.202214f
C1872 VOUT+.t43 GNDA 0.301601f
C1873 VOUT+.t137 GNDA 0.306738f
C1874 VOUT+.t44 GNDA 0.301601f
C1875 VOUT+.n129 GNDA 0.202214f
C1876 VOUT+.n130 GNDA 0.245051f
C1877 VOUT+.t52 GNDA 0.306738f
C1878 VOUT+.t103 GNDA 0.301601f
C1879 VOUT+.n131 GNDA 0.197501f
C1880 VOUT+.t88 GNDA 0.306738f
C1881 VOUT+.t136 GNDA 0.301601f
C1882 VOUT+.n132 GNDA 0.197501f
C1883 VOUT+.t123 GNDA 0.306738f
C1884 VOUT+.t29 GNDA 0.301601f
C1885 VOUT+.n133 GNDA 0.197501f
C1886 VOUT+.t26 GNDA 0.306738f
C1887 VOUT+.t151 GNDA 0.301601f
C1888 VOUT+.n134 GNDA 0.197501f
C1889 VOUT+.t68 GNDA 0.306738f
C1890 VOUT+.t55 GNDA 0.301601f
C1891 VOUT+.n135 GNDA 0.199386f
C1892 VOUT+.t91 GNDA 0.306347f
C1893 VOUT+.t114 GNDA 0.306738f
C1894 VOUT+.t72 GNDA 0.301601f
C1895 VOUT+.n136 GNDA 0.202214f
C1896 VOUT+.t96 GNDA 0.301601f
C1897 VOUT+.n137 GNDA 0.13195f
C1898 VOUT+.t57 GNDA 0.301601f
C1899 VOUT+.n138 GNDA 0.262925f
C1900 VOUT+.t156 GNDA 0.301601f
C1901 VOUT+.n139 GNDA 0.195098f
C1902 VOUT+.t121 GNDA 0.301601f
C1903 VOUT+.n140 GNDA 0.193213f
C1904 VOUT+.t140 GNDA 0.301601f
C1905 VOUT+.n141 GNDA 0.193213f
C1906 VOUT+.t108 GNDA 0.301601f
C1907 VOUT+.n142 GNDA 0.193213f
C1908 VOUT+.t64 GNDA 0.301601f
C1909 VOUT+.n143 GNDA 0.193213f
C1910 VOUT+.t89 GNDA 0.301601f
C1911 VOUT+.n144 GNDA 0.13195f
C1912 VOUT+.t46 GNDA 0.301601f
C1913 VOUT+.n145 GNDA 0.13195f
C1914 VOUT+.t40 GNDA 0.301601f
C1915 VOUT+.t144 GNDA 0.306738f
C1916 VOUT+.t77 GNDA 0.301601f
C1917 VOUT+.n146 GNDA 0.202214f
C1918 VOUT+.n147 GNDA 0.188501f
C1919 VOUT+.t124 GNDA 0.306738f
C1920 VOUT+.t83 GNDA 0.301601f
C1921 VOUT+.n148 GNDA 0.202214f
C1922 VOUT+.t79 GNDA 0.301601f
C1923 VOUT+.t33 GNDA 0.306738f
C1924 VOUT+.t117 GNDA 0.301601f
C1925 VOUT+.n149 GNDA 0.202214f
C1926 VOUT+.n150 GNDA 0.245051f
C1927 VOUT+.t139 GNDA 0.306738f
C1928 VOUT+.t110 GNDA 0.301601f
C1929 VOUT+.n151 GNDA 0.202214f
C1930 VOUT+.t80 GNDA 0.301601f
C1931 VOUT+.t27 GNDA 0.306738f
C1932 VOUT+.t81 GNDA 0.301601f
C1933 VOUT+.n152 GNDA 0.202214f
C1934 VOUT+.n153 GNDA 0.245051f
C1935 VOUT+.t106 GNDA 0.306738f
C1936 VOUT+.t66 GNDA 0.301601f
C1937 VOUT+.n154 GNDA 0.202214f
C1938 VOUT+.t35 GNDA 0.301601f
C1939 VOUT+.t132 GNDA 0.306738f
C1940 VOUT+.t37 GNDA 0.301601f
C1941 VOUT+.n155 GNDA 0.202214f
C1942 VOUT+.n156 GNDA 0.245051f
C1943 VOUT+.t133 GNDA 0.306738f
C1944 VOUT+.t104 GNDA 0.301601f
C1945 VOUT+.n157 GNDA 0.202214f
C1946 VOUT+.t75 GNDA 0.301601f
C1947 VOUT+.t21 GNDA 0.306738f
C1948 VOUT+.t76 GNDA 0.301601f
C1949 VOUT+.n158 GNDA 0.202214f
C1950 VOUT+.n159 GNDA 0.245051f
C1951 VOUT+.t98 GNDA 0.306738f
C1952 VOUT+.t61 GNDA 0.301601f
C1953 VOUT+.n160 GNDA 0.202214f
C1954 VOUT+.t30 GNDA 0.301601f
C1955 VOUT+.t126 GNDA 0.306738f
C1956 VOUT+.t31 GNDA 0.301601f
C1957 VOUT+.n161 GNDA 0.202214f
C1958 VOUT+.n162 GNDA 0.245051f
C1959 VOUT+.t59 GNDA 0.306738f
C1960 VOUT+.t19 GNDA 0.301601f
C1961 VOUT+.n163 GNDA 0.202214f
C1962 VOUT+.t134 GNDA 0.301601f
C1963 VOUT+.t90 GNDA 0.306738f
C1964 VOUT+.t135 GNDA 0.301601f
C1965 VOUT+.n164 GNDA 0.202214f
C1966 VOUT+.n165 GNDA 0.245051f
C1967 VOUT+.t92 GNDA 0.306738f
C1968 VOUT+.t58 GNDA 0.301601f
C1969 VOUT+.n166 GNDA 0.202214f
C1970 VOUT+.t24 GNDA 0.301601f
C1971 VOUT+.t125 GNDA 0.306738f
C1972 VOUT+.t25 GNDA 0.301601f
C1973 VOUT+.n167 GNDA 0.202214f
C1974 VOUT+.n168 GNDA 0.245051f
C1975 VOUT+.t49 GNDA 0.306738f
C1976 VOUT+.t152 GNDA 0.301601f
C1977 VOUT+.n169 GNDA 0.202214f
C1978 VOUT+.t127 GNDA 0.301601f
C1979 VOUT+.t82 GNDA 0.306738f
C1980 VOUT+.t128 GNDA 0.301601f
C1981 VOUT+.n170 GNDA 0.202214f
C1982 VOUT+.n171 GNDA 0.245051f
C1983 VOUT+.t149 GNDA 0.306738f
C1984 VOUT+.t118 GNDA 0.301601f
C1985 VOUT+.n172 GNDA 0.202214f
C1986 VOUT+.t93 GNDA 0.301601f
C1987 VOUT+.t39 GNDA 0.306738f
C1988 VOUT+.t95 GNDA 0.301601f
C1989 VOUT+.n173 GNDA 0.202214f
C1990 VOUT+.n174 GNDA 0.245051f
C1991 VOUT+.t116 GNDA 0.306738f
C1992 VOUT+.t74 GNDA 0.301601f
C1993 VOUT+.n175 GNDA 0.202214f
C1994 VOUT+.t50 GNDA 0.301601f
C1995 VOUT+.t143 GNDA 0.306738f
C1996 VOUT+.t54 GNDA 0.301601f
C1997 VOUT+.n176 GNDA 0.202214f
C1998 VOUT+.n177 GNDA 0.245051f
C1999 VOUT+.t32 GNDA 0.306738f
C2000 VOUT+.t87 GNDA 0.301601f
C2001 VOUT+.n178 GNDA 0.202214f
C2002 VOUT+.t86 GNDA 0.301601f
C2003 VOUT+.n179 GNDA 0.245051f
C2004 VOUT+.t115 GNDA 0.301601f
C2005 VOUT+.n180 GNDA 0.129123f
C2006 VOUT+.t145 GNDA 0.301601f
C2007 VOUT+.n181 GNDA 0.336474f
C2008 VOUT+.n182 GNDA 0.277096f
C2009 VOUT+.n183 GNDA 0.05655f
C2010 VOUT+.n184 GNDA 0.05655f
C2011 VOUT+.n186 GNDA 0.546652f
C2012 VOUT+.n187 GNDA 0.056967f
C2013 VOUT+.n188 GNDA 1.12158f
C2014 VOUT+.n189 GNDA 0.038454f
C2015 VOUT+.n191 GNDA 0.036192f
C2016 VOUT+.n192 GNDA 1.11215f
C2017 VOUT+.n194 GNDA 0.038454f
C2018 VOUT+.n195 GNDA 0.0754f
C2019 VOUT+.n196 GNDA 0.085956f
C2020 two_stage_opamp_dummy_magic_25_0.VD3.n0 GNDA 0.150417f
C2021 two_stage_opamp_dummy_magic_25_0.VD3.n1 GNDA 0.150417f
C2022 two_stage_opamp_dummy_magic_25_0.VD3.n2 GNDA 0.099935f
C2023 two_stage_opamp_dummy_magic_25_0.VD3.n3 GNDA 0.822594f
C2024 two_stage_opamp_dummy_magic_25_0.VD3.n4 GNDA 0.075209f
C2025 two_stage_opamp_dummy_magic_25_0.VD3.n5 GNDA 0.201695f
C2026 two_stage_opamp_dummy_magic_25_0.VD3.n6 GNDA 0.150417f
C2027 two_stage_opamp_dummy_magic_25_0.VD3.n7 GNDA 0.150417f
C2028 two_stage_opamp_dummy_magic_25_0.VD3.n8 GNDA 0.099935f
C2029 two_stage_opamp_dummy_magic_25_0.VD3.n9 GNDA 0.150417f
C2030 two_stage_opamp_dummy_magic_25_0.VD3.n10 GNDA 0.075209f
C2031 two_stage_opamp_dummy_magic_25_0.VD3.n11 GNDA 0.150417f
C2032 two_stage_opamp_dummy_magic_25_0.VD3.n12 GNDA 0.075209f
C2033 two_stage_opamp_dummy_magic_25_0.VD3.n13 GNDA 0.150417f
C2034 two_stage_opamp_dummy_magic_25_0.VD3.n14 GNDA 0.099935f
C2035 two_stage_opamp_dummy_magic_25_0.VD3.n15 GNDA 0.150417f
C2036 two_stage_opamp_dummy_magic_25_0.VD3.n16 GNDA 0.075209f
C2037 two_stage_opamp_dummy_magic_25_0.VD3.n17 GNDA 0.39821f
C2038 two_stage_opamp_dummy_magic_25_0.VD3.n18 GNDA 0.075209f
C2039 two_stage_opamp_dummy_magic_25_0.VD3.n19 GNDA 0.099935f
C2040 two_stage_opamp_dummy_magic_25_0.VD3.n20 GNDA 0.204473f
C2041 two_stage_opamp_dummy_magic_25_0.VD3.n21 GNDA 0.469399f
C2042 two_stage_opamp_dummy_magic_25_0.VD3.n22 GNDA 0.32328f
C2043 two_stage_opamp_dummy_magic_25_0.VD3.n23 GNDA 0.253736f
C2044 two_stage_opamp_dummy_magic_25_0.VD3.t22 GNDA 0.05484f
C2045 two_stage_opamp_dummy_magic_25_0.VD3.n24 GNDA 0.101472f
C2046 two_stage_opamp_dummy_magic_25_0.VD3.n25 GNDA 0.101472f
C2047 two_stage_opamp_dummy_magic_25_0.VD3.t26 GNDA 0.05484f
C2048 two_stage_opamp_dummy_magic_25_0.VD3.t29 GNDA 0.05484f
C2049 two_stage_opamp_dummy_magic_25_0.VD3.n26 GNDA 0.11218f
C2050 two_stage_opamp_dummy_magic_25_0.VD3.n27 GNDA 0.309358f
C2051 two_stage_opamp_dummy_magic_25_0.VD3.t32 GNDA 0.05484f
C2052 two_stage_opamp_dummy_magic_25_0.VD3.t24 GNDA 0.05484f
C2053 two_stage_opamp_dummy_magic_25_0.VD3.n28 GNDA 0.11218f
C2054 two_stage_opamp_dummy_magic_25_0.VD3.n29 GNDA 0.332049f
C2055 two_stage_opamp_dummy_magic_25_0.VD3.t27 GNDA 0.05484f
C2056 two_stage_opamp_dummy_magic_25_0.VD3.t30 GNDA 0.05484f
C2057 two_stage_opamp_dummy_magic_25_0.VD3.n30 GNDA 0.11218f
C2058 two_stage_opamp_dummy_magic_25_0.VD3.n31 GNDA 0.309358f
C2059 two_stage_opamp_dummy_magic_25_0.VD3.t13 GNDA 0.096159f
C2060 two_stage_opamp_dummy_magic_25_0.VD3.n32 GNDA 0.219169f
C2061 two_stage_opamp_dummy_magic_25_0.VD3.t21 GNDA 0.05484f
C2062 two_stage_opamp_dummy_magic_25_0.VD3.t37 GNDA 0.05484f
C2063 two_stage_opamp_dummy_magic_25_0.VD3.n33 GNDA 0.116347f
C2064 two_stage_opamp_dummy_magic_25_0.VD3.n34 GNDA 0.441622f
C2065 two_stage_opamp_dummy_magic_25_0.VD3.t35 GNDA 0.05484f
C2066 two_stage_opamp_dummy_magic_25_0.VD3.t5 GNDA 0.05484f
C2067 two_stage_opamp_dummy_magic_25_0.VD3.n35 GNDA 0.116347f
C2068 two_stage_opamp_dummy_magic_25_0.VD3.t3 GNDA 0.05484f
C2069 two_stage_opamp_dummy_magic_25_0.VD3.t9 GNDA 0.05484f
C2070 two_stage_opamp_dummy_magic_25_0.VD3.n36 GNDA 0.116347f
C2071 two_stage_opamp_dummy_magic_25_0.VD3.t19 GNDA 0.05484f
C2072 two_stage_opamp_dummy_magic_25_0.VD3.t1 GNDA 0.05484f
C2073 two_stage_opamp_dummy_magic_25_0.VD3.n37 GNDA 0.116347f
C2074 two_stage_opamp_dummy_magic_25_0.VD3.t7 GNDA 0.05484f
C2075 two_stage_opamp_dummy_magic_25_0.VD3.t17 GNDA 0.05484f
C2076 two_stage_opamp_dummy_magic_25_0.VD3.n38 GNDA 0.116347f
C2077 two_stage_opamp_dummy_magic_25_0.VD3.n39 GNDA 0.490884f
C2078 two_stage_opamp_dummy_magic_25_0.VD3.t10 GNDA 0.096159f
C2079 two_stage_opamp_dummy_magic_25_0.VD3.t12 GNDA 0.195072f
C2080 two_stage_opamp_dummy_magic_25_0.VD3.t15 GNDA 0.195072f
C2081 two_stage_opamp_dummy_magic_25_0.VD3.n40 GNDA 0.565887f
C2082 two_stage_opamp_dummy_magic_25_0.VD3.t14 GNDA 0.467448f
C2083 two_stage_opamp_dummy_magic_25_0.VD3.t20 GNDA 0.366642f
C2084 two_stage_opamp_dummy_magic_25_0.VD3.t36 GNDA 0.366642f
C2085 two_stage_opamp_dummy_magic_25_0.VD3.t34 GNDA 0.366642f
C2086 two_stage_opamp_dummy_magic_25_0.VD3.t4 GNDA 0.366642f
C2087 two_stage_opamp_dummy_magic_25_0.VD3.t2 GNDA 0.366642f
C2088 two_stage_opamp_dummy_magic_25_0.VD3.t8 GNDA 0.366642f
C2089 two_stage_opamp_dummy_magic_25_0.VD3.t18 GNDA 0.366642f
C2090 two_stage_opamp_dummy_magic_25_0.VD3.t0 GNDA 0.366642f
C2091 two_stage_opamp_dummy_magic_25_0.VD3.t6 GNDA 0.366642f
C2092 two_stage_opamp_dummy_magic_25_0.VD3.t16 GNDA 0.366642f
C2093 two_stage_opamp_dummy_magic_25_0.VD3.t11 GNDA 0.467448f
C2094 two_stage_opamp_dummy_magic_25_0.VD3.n41 GNDA 0.565887f
C2095 two_stage_opamp_dummy_magic_25_0.VD3.n42 GNDA 0.231296f
C2096 two_stage_opamp_dummy_magic_25_0.VD3.n43 GNDA 0.271333f
C2097 two_stage_opamp_dummy_magic_25_0.VD3.n44 GNDA 0.441622f
C2098 two_stage_opamp_dummy_magic_25_0.VD3.n45 GNDA 0.441622f
C2099 two_stage_opamp_dummy_magic_25_0.VD3.n46 GNDA 0.441622f
C2100 two_stage_opamp_dummy_magic_25_0.VD3.n47 GNDA 0.154506f
C2101 two_stage_opamp_dummy_magic_25_0.VD3.n48 GNDA 0.747385f
C2102 two_stage_opamp_dummy_magic_25_0.VD3.t28 GNDA 0.05484f
C2103 two_stage_opamp_dummy_magic_25_0.VD3.t33 GNDA 0.05484f
C2104 two_stage_opamp_dummy_magic_25_0.VD3.n49 GNDA 0.11218f
C2105 two_stage_opamp_dummy_magic_25_0.VD3.n50 GNDA 0.317096f
C2106 two_stage_opamp_dummy_magic_25_0.VD3.n51 GNDA 0.154506f
C2107 two_stage_opamp_dummy_magic_25_0.VD3.n52 GNDA 0.172095f
C2108 two_stage_opamp_dummy_magic_25_0.VD3.n53 GNDA 0.154506f
C2109 two_stage_opamp_dummy_magic_25_0.VD3.t23 GNDA 0.05484f
C2110 two_stage_opamp_dummy_magic_25_0.VD3.t25 GNDA 0.05484f
C2111 two_stage_opamp_dummy_magic_25_0.VD3.n54 GNDA 0.11218f
C2112 two_stage_opamp_dummy_magic_25_0.VD3.n55 GNDA 0.309358f
C2113 two_stage_opamp_dummy_magic_25_0.VD3.n56 GNDA 0.059483f
C2114 two_stage_opamp_dummy_magic_25_0.VD3.n57 GNDA 0.059483f
C2115 two_stage_opamp_dummy_magic_25_0.VD3.n58 GNDA 0.309358f
C2116 two_stage_opamp_dummy_magic_25_0.VD3.n59 GNDA 0.11218f
C2117 two_stage_opamp_dummy_magic_25_0.VD3.t31 GNDA 0.05484f
C2118 VDDA.n15 GNDA 0.745551f
C2119 VDDA.n16 GNDA 0.676197f
C2120 VDDA.n17 GNDA 2.42737f
C2121 VDDA.n44 GNDA 0.018205f
C2122 VDDA.n48 GNDA 0.017555f
C2123 VDDA.n52 GNDA 0.016255f
C2124 VDDA.n56 GNDA 0.018205f
C2125 VDDA.n60 GNDA 0.017555f
C2126 VDDA.n64 GNDA 0.016255f
C2127 VDDA.n68 GNDA 0.018205f
C2128 VDDA.n72 GNDA 0.017555f
C2129 VDDA.n76 GNDA 0.016255f
C2130 VDDA.n80 GNDA 0.018205f
C2131 VDDA.n84 GNDA 0.017555f
C2132 VDDA.n91 GNDA 0.050713f
C2133 VDDA.n92 GNDA 0.018205f
C2134 VDDA.n98 GNDA 0.016255f
C2135 VDDA.n99 GNDA 0.016255f
C2136 VDDA.n100 GNDA 0.017555f
C2137 VDDA.n106 GNDA 0.018205f
C2138 VDDA.n107 GNDA 0.017555f
C2139 VDDA.n108 GNDA 0.016255f
C2140 VDDA.n114 GNDA 0.017555f
C2141 VDDA.n115 GNDA 0.018205f
C2142 VDDA.n116 GNDA 0.018205f
C2143 VDDA.n122 GNDA 0.016255f
C2144 VDDA.n123 GNDA 0.016255f
C2145 VDDA.n124 GNDA 0.017555f
C2146 VDDA.n130 GNDA 0.018205f
C2147 VDDA.n131 GNDA 0.017555f
C2148 VDDA.n132 GNDA 0.016255f
C2149 VDDA.n138 GNDA 0.017555f
C2150 VDDA.n139 GNDA 0.018205f
C2151 VDDA.n140 GNDA 0.018205f
C2152 VDDA.n146 GNDA 0.016255f
C2153 VDDA.n147 GNDA 0.016255f
C2154 VDDA.n148 GNDA 0.017555f
C2155 VDDA.n154 GNDA 0.018205f
C2156 VDDA.n155 GNDA 0.017555f
C2157 VDDA.n156 GNDA 0.016255f
C2158 VDDA.n162 GNDA 0.017555f
C2159 VDDA.n163 GNDA 0.018205f
C2160 VDDA.n164 GNDA 0.018205f
C2161 VDDA.n170 GNDA 0.016255f
C2162 VDDA.n171 GNDA 0.016255f
C2163 VDDA.n172 GNDA 0.017555f
C2164 VDDA.n178 GNDA 0.018205f
C2165 VDDA.n179 GNDA 0.017555f
C2166 VDDA.n181 GNDA 0.010403f
C2167 VDDA.n182 GNDA 0.010403f
C2168 VDDA.n184 GNDA 0.010403f
C2169 VDDA.n187 GNDA 0.010403f
C2170 VDDA.n190 GNDA 0.040312f
C2171 VDDA.n191 GNDA 0.010403f
C2172 VDDA.n192 GNDA 0.017555f
C2173 VDDA.n195 GNDA 4.6987f
C2174 VDDA.n222 GNDA 0.018205f
C2175 VDDA.n226 GNDA 0.017555f
C2176 VDDA.n230 GNDA 0.016255f
C2177 VDDA.n234 GNDA 0.018205f
C2178 VDDA.n238 GNDA 0.017555f
C2179 VDDA.n242 GNDA 0.016255f
C2180 VDDA.n246 GNDA 0.018205f
C2181 VDDA.n250 GNDA 0.017555f
C2182 VDDA.n254 GNDA 0.016255f
C2183 VDDA.n258 GNDA 0.018205f
C2184 VDDA.n262 GNDA 0.017555f
C2185 VDDA.n269 GNDA 0.050713f
C2186 VDDA.n270 GNDA 0.018205f
C2187 VDDA.n276 GNDA 0.016255f
C2188 VDDA.n277 GNDA 0.016255f
C2189 VDDA.n278 GNDA 0.017555f
C2190 VDDA.n284 GNDA 0.018205f
C2191 VDDA.n285 GNDA 0.017555f
C2192 VDDA.n286 GNDA 0.016255f
C2193 VDDA.n292 GNDA 0.017555f
C2194 VDDA.n293 GNDA 0.018205f
C2195 VDDA.n294 GNDA 0.018205f
C2196 VDDA.n300 GNDA 0.016255f
C2197 VDDA.n301 GNDA 0.016255f
C2198 VDDA.n302 GNDA 0.017555f
C2199 VDDA.n308 GNDA 0.018205f
C2200 VDDA.n309 GNDA 0.017555f
C2201 VDDA.n310 GNDA 0.016255f
C2202 VDDA.n316 GNDA 0.017555f
C2203 VDDA.n317 GNDA 0.018205f
C2204 VDDA.n318 GNDA 0.018205f
C2205 VDDA.n324 GNDA 0.016255f
C2206 VDDA.n325 GNDA 0.016255f
C2207 VDDA.n326 GNDA 0.017555f
C2208 VDDA.n332 GNDA 0.018205f
C2209 VDDA.n333 GNDA 0.017555f
C2210 VDDA.n334 GNDA 0.016255f
C2211 VDDA.n340 GNDA 0.017555f
C2212 VDDA.n341 GNDA 0.018205f
C2213 VDDA.n342 GNDA 0.018205f
C2214 VDDA.n348 GNDA 0.016255f
C2215 VDDA.n349 GNDA 0.016255f
C2216 VDDA.n350 GNDA 0.017555f
C2217 VDDA.n356 GNDA 0.018205f
C2218 VDDA.n357 GNDA 0.017555f
C2219 VDDA.n359 GNDA 0.010403f
C2220 VDDA.n361 GNDA 0.010403f
C2221 VDDA.n364 GNDA 0.098597f
C2222 VDDA.t259 GNDA 0.013301f
C2223 VDDA.n365 GNDA 0.029046f
C2224 VDDA.n366 GNDA 0.010403f
C2225 VDDA.n370 GNDA 0.06957f
C2226 VDDA.n371 GNDA 0.028379f
C2227 VDDA.t280 GNDA 0.014081f
C2228 VDDA.n372 GNDA 0.042396f
C2229 VDDA.t278 GNDA 0.037744f
C2230 VDDA.t25 GNDA 0.028608f
C2231 VDDA.t263 GNDA 0.037744f
C2232 VDDA.t264 GNDA 0.014081f
C2233 VDDA.n373 GNDA 0.042396f
C2234 VDDA.n374 GNDA 0.027863f
C2235 VDDA.n375 GNDA 0.056694f
C2236 VDDA.n376 GNDA 0.090162f
C2237 VDDA.t296 GNDA 0.013433f
C2238 VDDA.n377 GNDA 0.017272f
C2239 VDDA.t270 GNDA 0.034568f
C2240 VDDA.t268 GNDA 0.013433f
C2241 VDDA.n378 GNDA 0.035167f
C2242 VDDA.n379 GNDA 0.086305f
C2243 VDDA.t269 GNDA 0.064659f
C2244 VDDA.t208 GNDA 0.050715f
C2245 VDDA.t297 GNDA 0.064659f
C2246 VDDA.t298 GNDA 0.026983f
C2247 VDDA.n380 GNDA 0.086305f
C2248 VDDA.n381 GNDA 0.034652f
C2249 VDDA.n382 GNDA 0.060372f
C2250 VDDA.n383 GNDA 0.056434f
C2251 VDDA.n384 GNDA 0.343653f
C2252 VDDA.n385 GNDA 0.010403f
C2253 VDDA.n387 GNDA 0.010403f
C2254 VDDA.n388 GNDA 0.010403f
C2255 VDDA.t411 GNDA 0.013004f
C2256 VDDA.t82 GNDA 0.013004f
C2257 VDDA.n389 GNDA 0.033462f
C2258 VDDA.n390 GNDA 0.114131f
C2259 VDDA.t76 GNDA 0.013004f
C2260 VDDA.t168 GNDA 0.013004f
C2261 VDDA.n391 GNDA 0.033462f
C2262 VDDA.n392 GNDA 0.114131f
C2263 VDDA.t36 GNDA 0.013004f
C2264 VDDA.t382 GNDA 0.013004f
C2265 VDDA.n393 GNDA 0.033462f
C2266 VDDA.n394 GNDA 0.114131f
C2267 VDDA.t116 GNDA 0.013004f
C2268 VDDA.t152 GNDA 0.013004f
C2269 VDDA.n395 GNDA 0.033462f
C2270 VDDA.n396 GNDA 0.114131f
C2271 VDDA.t387 GNDA 0.013004f
C2272 VDDA.t74 GNDA 0.013004f
C2273 VDDA.n397 GNDA 0.033462f
C2274 VDDA.n398 GNDA 0.134441f
C2275 VDDA.t338 GNDA 0.015777f
C2276 VDDA.n399 GNDA 0.042161f
C2277 VDDA.t340 GNDA 0.045764f
C2278 VDDA.n400 GNDA 0.153083f
C2279 VDDA.t339 GNDA 0.099148f
C2280 VDDA.t73 GNDA 0.076289f
C2281 VDDA.t386 GNDA 0.076289f
C2282 VDDA.t151 GNDA 0.076289f
C2283 VDDA.t115 GNDA 0.076289f
C2284 VDDA.t381 GNDA 0.076289f
C2285 VDDA.t35 GNDA 0.076289f
C2286 VDDA.t167 GNDA 0.076289f
C2287 VDDA.t75 GNDA 0.076289f
C2288 VDDA.t81 GNDA 0.076289f
C2289 VDDA.t410 GNDA 0.076289f
C2290 VDDA.t324 GNDA 0.099148f
C2291 VDDA.t325 GNDA 0.045764f
C2292 VDDA.n401 GNDA 0.153083f
C2293 VDDA.t323 GNDA 0.015777f
C2294 VDDA.n402 GNDA 0.040896f
C2295 VDDA.n403 GNDA 0.049534f
C2296 VDDA.n405 GNDA 0.010305f
C2297 VDDA.n406 GNDA 0.010403f
C2298 VDDA.n407 GNDA 0.010403f
C2299 VDDA.n408 GNDA 0.010305f
C2300 VDDA.n409 GNDA 0.010403f
C2301 VDDA.n410 GNDA 0.010403f
C2302 VDDA.n411 GNDA 0.010403f
C2303 VDDA.n413 GNDA 0.018392f
C2304 VDDA.n414 GNDA 0.018107f
C2305 VDDA.n415 GNDA 0.142303f
C2306 VDDA.n416 GNDA 0.018107f
C2307 VDDA.n417 GNDA 0.075845f
C2308 VDDA.n418 GNDA 0.018107f
C2309 VDDA.n419 GNDA 0.075845f
C2310 VDDA.n420 GNDA 0.018107f
C2311 VDDA.n421 GNDA 0.075845f
C2312 VDDA.n422 GNDA 0.018107f
C2313 VDDA.n423 GNDA 0.101852f
C2314 VDDA.n424 GNDA 0.045513f
C2315 VDDA.n426 GNDA 0.139141f
C2316 VDDA.n428 GNDA 0.139141f
C2317 VDDA.n430 GNDA 0.056318f
C2318 VDDA.t358 GNDA 0.015464f
C2319 VDDA.n431 GNDA 0.047508f
C2320 VDDA.t357 GNDA 0.038526f
C2321 VDDA.t384 GNDA 0.028608f
C2322 VDDA.t94 GNDA 0.028608f
C2323 VDDA.t14 GNDA 0.028608f
C2324 VDDA.t380 GNDA 0.028608f
C2325 VDDA.t21 GNDA 0.028608f
C2326 VDDA.t83 GNDA 0.028608f
C2327 VDDA.t383 GNDA 0.028608f
C2328 VDDA.t413 GNDA 0.028608f
C2329 VDDA.t412 GNDA 0.028608f
C2330 VDDA.t6 GNDA 0.028608f
C2331 VDDA.t330 GNDA 0.038526f
C2332 VDDA.t331 GNDA 0.015464f
C2333 VDDA.n432 GNDA 0.047508f
C2334 VDDA.n433 GNDA 0.034052f
C2335 VDDA.n434 GNDA 0.197651f
C2336 VDDA.n435 GNDA 0.038361f
C2337 VDDA.n437 GNDA 0.146943f
C2338 VDDA.n438 GNDA 0.018864f
C2339 VDDA.n439 GNDA 0.064144f
C2340 VDDA.n440 GNDA 0.016255f
C2341 VDDA.t288 GNDA 0.038497f
C2342 VDDA.n446 GNDA 0.011823f
C2343 VDDA.n448 GNDA 0.010403f
C2344 VDDA.n450 GNDA 0.169699f
C2345 VDDA.n451 GNDA 0.098597f
C2346 VDDA.t347 GNDA 0.013301f
C2347 VDDA.n452 GNDA 0.029046f
C2348 VDDA.n453 GNDA 0.010403f
C2349 VDDA.n456 GNDA 0.085825f
C2350 VDDA.n457 GNDA 0.010403f
C2351 VDDA.n458 GNDA 0.017555f
C2352 VDDA.n461 GNDA 2.42737f
C2353 VDDA.n488 GNDA 0.018205f
C2354 VDDA.n492 GNDA 0.017555f
C2355 VDDA.n496 GNDA 0.016255f
C2356 VDDA.n500 GNDA 0.018205f
C2357 VDDA.n504 GNDA 0.017555f
C2358 VDDA.n508 GNDA 0.016255f
C2359 VDDA.n512 GNDA 0.018205f
C2360 VDDA.n516 GNDA 0.017555f
C2361 VDDA.n520 GNDA 0.016255f
C2362 VDDA.n524 GNDA 0.018205f
C2363 VDDA.n528 GNDA 0.017555f
C2364 VDDA.n535 GNDA 0.050713f
C2365 VDDA.n536 GNDA 0.018205f
C2366 VDDA.n542 GNDA 0.016255f
C2367 VDDA.n543 GNDA 0.016255f
C2368 VDDA.n544 GNDA 0.017555f
C2369 VDDA.n550 GNDA 0.018205f
C2370 VDDA.n551 GNDA 0.017555f
C2371 VDDA.n552 GNDA 0.016255f
C2372 VDDA.n558 GNDA 0.017555f
C2373 VDDA.n559 GNDA 0.018205f
C2374 VDDA.n560 GNDA 0.018205f
C2375 VDDA.n566 GNDA 0.016255f
C2376 VDDA.n567 GNDA 0.016255f
C2377 VDDA.n568 GNDA 0.017555f
C2378 VDDA.n574 GNDA 0.018205f
C2379 VDDA.n575 GNDA 0.017555f
C2380 VDDA.n576 GNDA 0.016255f
C2381 VDDA.n582 GNDA 0.017555f
C2382 VDDA.n583 GNDA 0.018205f
C2383 VDDA.n584 GNDA 0.018205f
C2384 VDDA.n590 GNDA 0.016255f
C2385 VDDA.n591 GNDA 0.016255f
C2386 VDDA.n592 GNDA 0.017555f
C2387 VDDA.n598 GNDA 0.018205f
C2388 VDDA.n599 GNDA 0.017555f
C2389 VDDA.n600 GNDA 0.016255f
C2390 VDDA.n606 GNDA 0.017555f
C2391 VDDA.n607 GNDA 0.018205f
C2392 VDDA.n608 GNDA 0.018205f
C2393 VDDA.n614 GNDA 0.016255f
C2394 VDDA.n615 GNDA 0.016255f
C2395 VDDA.n616 GNDA 0.017555f
C2396 VDDA.n622 GNDA 0.018205f
C2397 VDDA.n623 GNDA 0.017555f
C2398 VDDA.n625 GNDA 0.010403f
C2399 VDDA.n627 GNDA 0.010403f
C2400 VDDA.n630 GNDA 0.010403f
C2401 VDDA.n633 GNDA 0.040312f
C2402 VDDA.n634 GNDA 0.010403f
C2403 VDDA.n635 GNDA 0.017555f
C2404 VDDA.n664 GNDA 0.018205f
C2405 VDDA.n666 GNDA 0.017555f
C2406 VDDA.n668 GNDA 0.016255f
C2407 VDDA.n670 GNDA 0.018205f
C2408 VDDA.n672 GNDA 0.017555f
C2409 VDDA.n674 GNDA 0.016255f
C2410 VDDA.n676 GNDA 0.018205f
C2411 VDDA.n678 GNDA 0.017555f
C2412 VDDA.n680 GNDA 0.016255f
C2413 VDDA.n682 GNDA 0.018205f
C2414 VDDA.n684 GNDA 0.017555f
C2415 VDDA.n689 GNDA 0.050713f
C2416 VDDA.n690 GNDA 0.018205f
C2417 VDDA.n698 GNDA 0.016255f
C2418 VDDA.n699 GNDA 0.016255f
C2419 VDDA.n700 GNDA 0.017555f
C2420 VDDA.n708 GNDA 0.018205f
C2421 VDDA.n709 GNDA 0.017555f
C2422 VDDA.n710 GNDA 0.016255f
C2423 VDDA.n718 GNDA 0.017555f
C2424 VDDA.n719 GNDA 0.018205f
C2425 VDDA.n720 GNDA 0.018205f
C2426 VDDA.n728 GNDA 0.016255f
C2427 VDDA.n729 GNDA 0.016255f
C2428 VDDA.n730 GNDA 0.017555f
C2429 VDDA.n738 GNDA 0.018205f
C2430 VDDA.n739 GNDA 0.017555f
C2431 VDDA.n740 GNDA 0.016255f
C2432 VDDA.n748 GNDA 0.017555f
C2433 VDDA.n749 GNDA 0.018205f
C2434 VDDA.n750 GNDA 0.018205f
C2435 VDDA.n758 GNDA 0.016255f
C2436 VDDA.n759 GNDA 0.016255f
C2437 VDDA.n760 GNDA 0.017555f
C2438 VDDA.n768 GNDA 0.018205f
C2439 VDDA.n769 GNDA 0.017555f
C2440 VDDA.n770 GNDA 0.016255f
C2441 VDDA.n778 GNDA 0.017555f
C2442 VDDA.n779 GNDA 0.018205f
C2443 VDDA.n780 GNDA 0.018205f
C2444 VDDA.n788 GNDA 0.016255f
C2445 VDDA.n789 GNDA 0.016255f
C2446 VDDA.n790 GNDA 0.017555f
C2447 VDDA.n798 GNDA 0.018205f
C2448 VDDA.n799 GNDA 0.017555f
C2449 VDDA.n800 GNDA 0.010305f
C2450 VDDA.n801 GNDA 0.010403f
C2451 VDDA.n803 GNDA 0.010403f
C2452 VDDA.n804 GNDA 0.010403f
C2453 VDDA.n806 GNDA 0.27503f
C2454 VDDA.n807 GNDA 0.278281f
C2455 VDDA.n810 GNDA 1.62981f
C2456 VDDA.n836 GNDA 0.016255f
C2457 VDDA.n840 GNDA 0.018205f
C2458 VDDA.n844 GNDA 0.017555f
C2459 VDDA.n848 GNDA 0.016255f
C2460 VDDA.n852 GNDA 0.018205f
C2461 VDDA.n856 GNDA 0.017555f
C2462 VDDA.n860 GNDA 0.016255f
C2463 VDDA.n864 GNDA 0.018205f
C2464 VDDA.n868 GNDA 0.017555f
C2465 VDDA.n872 GNDA 0.016255f
C2466 VDDA.n876 GNDA 0.050713f
C2467 VDDA.n884 GNDA 0.018205f
C2468 VDDA.n885 GNDA 0.017555f
C2469 VDDA.n886 GNDA 0.016255f
C2470 VDDA.n892 GNDA 0.017555f
C2471 VDDA.n893 GNDA 0.018205f
C2472 VDDA.n894 GNDA 0.018205f
C2473 VDDA.n900 GNDA 0.016255f
C2474 VDDA.n901 GNDA 0.016255f
C2475 VDDA.n902 GNDA 0.017555f
C2476 VDDA.n908 GNDA 0.018205f
C2477 VDDA.n909 GNDA 0.017555f
C2478 VDDA.n910 GNDA 0.016255f
C2479 VDDA.n916 GNDA 0.017555f
C2480 VDDA.n917 GNDA 0.018205f
C2481 VDDA.n918 GNDA 0.018205f
C2482 VDDA.n924 GNDA 0.016255f
C2483 VDDA.n925 GNDA 0.016255f
C2484 VDDA.n926 GNDA 0.017555f
C2485 VDDA.n932 GNDA 0.018205f
C2486 VDDA.n933 GNDA 0.017555f
C2487 VDDA.n934 GNDA 0.016255f
C2488 VDDA.n940 GNDA 0.017555f
C2489 VDDA.n941 GNDA 0.018205f
C2490 VDDA.n942 GNDA 0.018205f
C2491 VDDA.n948 GNDA 0.016255f
C2492 VDDA.n949 GNDA 0.016255f
C2493 VDDA.n950 GNDA 0.017555f
C2494 VDDA.n956 GNDA 0.018205f
C2495 VDDA.n957 GNDA 0.017555f
C2496 VDDA.n958 GNDA 0.016255f
C2497 VDDA.n964 GNDA 0.017555f
C2498 VDDA.n965 GNDA 0.018205f
C2499 VDDA.n966 GNDA 0.018205f
C2500 VDDA.n970 GNDA 2.42737f
C2501 VDDA.n973 GNDA 0.278281f
C2502 VDDA.n974 GNDA 0.27503f
C2503 VDDA.n976 GNDA 0.040312f
C2504 VDDA.n977 GNDA 0.010403f
C2505 VDDA.n978 GNDA 0.040312f
C2506 VDDA.n979 GNDA 0.010403f
C2507 VDDA.n980 GNDA 0.017555f
C2508 VDDA.n984 GNDA 0.016255f
C2509 VDDA.n988 GNDA 0.018205f
C2510 VDDA.n992 GNDA 0.017555f
C2511 VDDA.n996 GNDA 0.016255f
C2512 VDDA.n1000 GNDA 0.018205f
C2513 VDDA.n1004 GNDA 0.017555f
C2514 VDDA.n1008 GNDA 0.016255f
C2515 VDDA.n1012 GNDA 0.018205f
C2516 VDDA.n1016 GNDA 0.017555f
C2517 VDDA.n1020 GNDA 0.016255f
C2518 VDDA.n1024 GNDA 0.050713f
C2519 VDDA.n1035 GNDA 0.018205f
C2520 VDDA.n1036 GNDA 0.017555f
C2521 VDDA.n1037 GNDA 0.016255f
C2522 VDDA.n1045 GNDA 0.017555f
C2523 VDDA.n1046 GNDA 0.018205f
C2524 VDDA.n1047 GNDA 0.018205f
C2525 VDDA.n1055 GNDA 0.016255f
C2526 VDDA.n1056 GNDA 0.016255f
C2527 VDDA.n1057 GNDA 0.017555f
C2528 VDDA.n1065 GNDA 0.018205f
C2529 VDDA.n1066 GNDA 0.017555f
C2530 VDDA.n1067 GNDA 0.016255f
C2531 VDDA.n1075 GNDA 0.017555f
C2532 VDDA.n1076 GNDA 0.018205f
C2533 VDDA.n1077 GNDA 0.018205f
C2534 VDDA.n1085 GNDA 0.016255f
C2535 VDDA.n1086 GNDA 0.016255f
C2536 VDDA.n1087 GNDA 0.017555f
C2537 VDDA.n1095 GNDA 0.018205f
C2538 VDDA.n1096 GNDA 0.017555f
C2539 VDDA.n1097 GNDA 0.016255f
C2540 VDDA.n1105 GNDA 0.017555f
C2541 VDDA.n1106 GNDA 0.018205f
C2542 VDDA.n1107 GNDA 0.018205f
C2543 VDDA.n1115 GNDA 0.016255f
C2544 VDDA.n1116 GNDA 0.016255f
C2545 VDDA.n1117 GNDA 0.017555f
C2546 VDDA.n1125 GNDA 0.018205f
C2547 VDDA.n1126 GNDA 0.017555f
C2548 VDDA.n1127 GNDA 0.016255f
C2549 VDDA.n1135 GNDA 0.017555f
C2550 VDDA.n1136 GNDA 0.018205f
C2551 VDDA.n1137 GNDA 0.018205f
C2552 VDDA.n1144 GNDA 0.278281f
C2553 VDDA.n1145 GNDA 0.27503f
C2554 VDDA.n1147 GNDA 0.040312f
C2555 VDDA.n1148 GNDA 0.010403f
C2556 VDDA.n1149 GNDA 0.040312f
C2557 VDDA.n1150 GNDA 0.010403f
C2558 VDDA.n1151 GNDA 0.040312f
C2559 VDDA.n1152 GNDA 0.010403f
C2560 VDDA.n1154 GNDA 0.27503f
C2561 VDDA.n1155 GNDA 0.278281f
C2562 VDDA.n1158 GNDA 3.64106f
C2563 VDDA.n1184 GNDA 0.016255f
C2564 VDDA.n1188 GNDA 0.018205f
C2565 VDDA.n1192 GNDA 0.017555f
C2566 VDDA.n1196 GNDA 0.016255f
C2567 VDDA.n1200 GNDA 0.018205f
C2568 VDDA.n1204 GNDA 0.017555f
C2569 VDDA.n1208 GNDA 0.016255f
C2570 VDDA.n1212 GNDA 0.018205f
C2571 VDDA.n1216 GNDA 0.017555f
C2572 VDDA.n1220 GNDA 0.016255f
C2573 VDDA.n1224 GNDA 0.050713f
C2574 VDDA.n1232 GNDA 0.018205f
C2575 VDDA.n1233 GNDA 0.017555f
C2576 VDDA.n1234 GNDA 0.016255f
C2577 VDDA.n1240 GNDA 0.017555f
C2578 VDDA.n1241 GNDA 0.018205f
C2579 VDDA.n1242 GNDA 0.018205f
C2580 VDDA.n1248 GNDA 0.016255f
C2581 VDDA.n1249 GNDA 0.016255f
C2582 VDDA.n1250 GNDA 0.017555f
C2583 VDDA.n1256 GNDA 0.018205f
C2584 VDDA.n1257 GNDA 0.017555f
C2585 VDDA.n1258 GNDA 0.016255f
C2586 VDDA.n1264 GNDA 0.017555f
C2587 VDDA.n1265 GNDA 0.018205f
C2588 VDDA.n1266 GNDA 0.018205f
C2589 VDDA.n1272 GNDA 0.016255f
C2590 VDDA.n1273 GNDA 0.016255f
C2591 VDDA.n1274 GNDA 0.017555f
C2592 VDDA.n1280 GNDA 0.018205f
C2593 VDDA.n1281 GNDA 0.017555f
C2594 VDDA.n1282 GNDA 0.016255f
C2595 VDDA.n1288 GNDA 0.017555f
C2596 VDDA.n1289 GNDA 0.018205f
C2597 VDDA.n1290 GNDA 0.018205f
C2598 VDDA.n1296 GNDA 0.016255f
C2599 VDDA.n1297 GNDA 0.016255f
C2600 VDDA.n1298 GNDA 0.017555f
C2601 VDDA.n1304 GNDA 0.018205f
C2602 VDDA.n1305 GNDA 0.017555f
C2603 VDDA.n1306 GNDA 0.016255f
C2604 VDDA.n1312 GNDA 0.017555f
C2605 VDDA.n1313 GNDA 0.018205f
C2606 VDDA.n1314 GNDA 0.018205f
C2607 VDDA.n1366 GNDA 0.589505f
C2608 VDDA.n1391 GNDA 0.052646f
C2609 VDDA.n1402 GNDA 0.054944f
C2610 VDDA.n1403 GNDA 0.015577f
C2611 VDDA.n1404 GNDA 0.017447f
C2612 VDDA.n1405 GNDA 0.017447f
C2613 VDDA.n1407 GNDA 0.015577f
C2614 VDDA.n1434 GNDA 0.018205f
C2615 VDDA.n1436 GNDA 0.017555f
C2616 VDDA.n1438 GNDA 0.016255f
C2617 VDDA.n1440 GNDA 0.018205f
C2618 VDDA.n1442 GNDA 0.017555f
C2619 VDDA.n1444 GNDA 0.016255f
C2620 VDDA.n1446 GNDA 0.018205f
C2621 VDDA.n1448 GNDA 0.017555f
C2622 VDDA.n1450 GNDA 0.016255f
C2623 VDDA.n1452 GNDA 0.018205f
C2624 VDDA.n1454 GNDA 0.017555f
C2625 VDDA.t420 GNDA 0.121152f
C2626 VDDA.t128 GNDA 0.121591f
C2627 VDDA.t102 GNDA 0.115089f
C2628 VDDA.t103 GNDA 0.121152f
C2629 VDDA.t406 GNDA 0.121591f
C2630 VDDA.t125 GNDA 0.115089f
C2631 VDDA.t391 GNDA 0.121152f
C2632 VDDA.t146 GNDA 0.121591f
C2633 VDDA.t372 GNDA 0.115089f
C2634 VDDA.t388 GNDA 0.121152f
C2635 VDDA.t90 GNDA 0.121591f
C2636 VDDA.t148 GNDA 0.115089f
C2637 VDDA.t101 GNDA 0.121152f
C2638 VDDA.t59 GNDA 0.121591f
C2639 VDDA.t63 GNDA 0.115089f
C2640 VDDA.n1456 GNDA 0.081208f
C2641 VDDA.t91 GNDA 0.06467f
C2642 VDDA.n1457 GNDA 0.088113f
C2643 VDDA.t62 GNDA 0.06467f
C2644 VDDA.n1458 GNDA 0.088113f
C2645 VDDA.t147 GNDA 0.06467f
C2646 VDDA.n1459 GNDA 0.088113f
C2647 VDDA.t145 GNDA 0.06467f
C2648 VDDA.n1460 GNDA 0.088113f
C2649 VDDA.t124 GNDA 0.326117f
C2650 VDDA.n1461 GNDA 1.38805f
C2651 VDDA.n1465 GNDA 0.017555f
C2652 VDDA.n1466 GNDA 0.018205f
C2653 VDDA.n1467 GNDA 0.018205f
C2654 VDDA.n1475 GNDA 0.016255f
C2655 VDDA.n1476 GNDA 0.016255f
C2656 VDDA.n1477 GNDA 0.017555f
C2657 VDDA.n1485 GNDA 0.018205f
C2658 VDDA.n1486 GNDA 0.017555f
C2659 VDDA.n1487 GNDA 0.016255f
C2660 VDDA.n1495 GNDA 0.017555f
C2661 VDDA.n1496 GNDA 0.018205f
C2662 VDDA.n1497 GNDA 0.018205f
C2663 VDDA.n1505 GNDA 0.016255f
C2664 VDDA.n1506 GNDA 0.016255f
C2665 VDDA.n1507 GNDA 0.017555f
C2666 VDDA.n1515 GNDA 0.018205f
C2667 VDDA.n1516 GNDA 0.017555f
C2668 VDDA.n1517 GNDA 0.016255f
C2669 VDDA.n1525 GNDA 0.017555f
C2670 VDDA.n1526 GNDA 0.018205f
C2671 VDDA.n1527 GNDA 0.018205f
C2672 VDDA.n1535 GNDA 0.016255f
C2673 VDDA.n1536 GNDA 0.016255f
C2674 VDDA.n1537 GNDA 0.017555f
C2675 VDDA.n1545 GNDA 0.018205f
C2676 VDDA.n1546 GNDA 0.017555f
C2677 VDDA.n1547 GNDA 0.016255f
C2678 VDDA.n1555 GNDA 0.017555f
C2679 VDDA.n1556 GNDA 0.018205f
C2680 VDDA.n1557 GNDA 0.018205f
C2681 VDDA.n1565 GNDA 0.016255f
C2682 VDDA.n1566 GNDA 0.016255f
C2683 VDDA.n1567 GNDA 0.017555f
C2684 VDDA.n1575 GNDA 0.050713f
C2685 VDDA.n1578 GNDA 5.21885f
C2686 VDDA.n1579 GNDA 3.15559f
C2687 VDDA.n1580 GNDA 0.017447f
C2688 VDDA.n1582 GNDA 0.015577f
C2689 VDDA.n1583 GNDA 0.017447f
C2690 VDDA.n1584 GNDA 0.016824f
C2691 VDDA.n1585 GNDA 0.016824f
C2692 VDDA.n1586 GNDA 0.015577f
C2693 VDDA.n1589 GNDA 0.017447f
C2694 VDDA.n1590 GNDA 0.015577f
C2695 VDDA.n1591 GNDA 0.015577f
C2696 VDDA.n1592 GNDA 0.017447f
C2697 VDDA.n1595 GNDA 0.016824f
C2698 VDDA.n1596 GNDA 0.017447f
C2699 VDDA.n1597 GNDA 0.017447f
C2700 VDDA.n1598 GNDA 0.016824f
C2701 VDDA.n1601 GNDA 0.015577f
C2702 VDDA.n1602 GNDA 0.016824f
C2703 VDDA.n1603 GNDA 0.016824f
C2704 VDDA.n1604 GNDA 0.015577f
C2705 VDDA.n1607 GNDA 0.017447f
C2706 VDDA.n1608 GNDA 0.015577f
C2707 VDDA.n1609 GNDA 0.015577f
C2708 VDDA.n1610 GNDA 0.017447f
C2709 VDDA.n1613 GNDA 0.016824f
C2710 VDDA.n1614 GNDA 0.017447f
C2711 VDDA.n1615 GNDA 0.017447f
C2712 VDDA.n1616 GNDA 0.016824f
C2713 VDDA.n1619 GNDA 0.015577f
C2714 VDDA.n1620 GNDA 0.016824f
C2715 VDDA.n1621 GNDA 0.016824f
C2716 VDDA.n1622 GNDA 0.015577f
C2717 VDDA.n1625 GNDA 0.017447f
C2718 VDDA.n1626 GNDA 0.015577f
C2719 VDDA.n1627 GNDA 0.015577f
C2720 VDDA.n1628 GNDA 0.017447f
C2721 VDDA.n1631 GNDA 0.016824f
C2722 VDDA.n1632 GNDA 0.017447f
C2723 VDDA.n1633 GNDA 0.017447f
C2724 VDDA.n1634 GNDA 0.016824f
C2725 VDDA.n1637 GNDA 0.015577f
C2726 VDDA.n1638 GNDA 0.016824f
C2727 VDDA.n1639 GNDA 0.016824f
C2728 VDDA.n1640 GNDA 0.015577f
C2729 VDDA.n1643 GNDA 0.017447f
C2730 VDDA.n1644 GNDA 0.015908f
C2731 VDDA.n1645 GNDA 0.017447f
C2732 VDDA.n1648 GNDA 0.016824f
C2733 VDDA.n1649 GNDA 0.016824f
C2734 VDDA.n1650 GNDA 0.017743f
C2735 VDDA.n1651 GNDA 0.047352f
C2736 VDDA.n1652 GNDA 0.017447f
C2737 VDDA.n1653 GNDA 0.017447f
C2738 VDDA.n1654 GNDA 0.017447f
C2739 VDDA.n1656 GNDA 0.016824f
C2740 VDDA.n1658 GNDA 0.015577f
C2741 VDDA.n1659 GNDA 0.015577f
C2742 VDDA.n1660 GNDA 0.015577f
C2743 VDDA.n1661 GNDA 0.015577f
C2744 VDDA.n1662 GNDA 0.016824f
C2745 VDDA.n1663 GNDA 0.016824f
C2746 VDDA.n1664 GNDA 0.016824f
C2747 VDDA.n1666 GNDA 0.017447f
C2748 VDDA.n1668 GNDA 0.017447f
C2749 VDDA.n1669 GNDA 0.017447f
C2750 VDDA.n1670 GNDA 0.017447f
C2751 VDDA.n1671 GNDA 0.016824f
C2752 VDDA.n1672 GNDA 0.015577f
C2753 VDDA.n1673 GNDA 0.015577f
C2754 VDDA.n1674 GNDA 0.015577f
C2755 VDDA.n1676 GNDA 0.015577f
C2756 VDDA.n1678 GNDA 0.016824f
C2757 VDDA.n1679 GNDA 0.016824f
C2758 VDDA.n1680 GNDA 0.016824f
C2759 VDDA.n1681 GNDA 0.017447f
C2760 VDDA.n1682 GNDA 0.017447f
C2761 VDDA.n1683 GNDA 0.017447f
C2762 VDDA.n1684 GNDA 0.017447f
C2763 VDDA.n1686 GNDA 0.016824f
C2764 VDDA.n1688 GNDA 0.015577f
C2765 VDDA.n1689 GNDA 0.015577f
C2766 VDDA.n1690 GNDA 0.015577f
C2767 VDDA.n1691 GNDA 0.015577f
C2768 VDDA.n1692 GNDA 0.016824f
C2769 VDDA.n1693 GNDA 0.016824f
C2770 VDDA.n1694 GNDA 0.016824f
C2771 VDDA.n1696 GNDA 0.017447f
C2772 VDDA.n1698 GNDA 0.017447f
C2773 VDDA.n1699 GNDA 0.017447f
C2774 VDDA.n1700 GNDA 0.017447f
C2775 VDDA.n1701 GNDA 0.016824f
C2776 VDDA.n1702 GNDA 0.015577f
C2777 VDDA.n1703 GNDA 0.015577f
C2778 VDDA.n1704 GNDA 0.015577f
C2779 VDDA.n1706 GNDA 0.015577f
C2780 VDDA.n1708 GNDA 0.016824f
C2781 VDDA.n1709 GNDA 0.016824f
C2782 VDDA.n1710 GNDA 0.016824f
C2783 VDDA.n1711 GNDA 0.017447f
C2784 VDDA.n1712 GNDA 0.017447f
C2785 VDDA.n1713 GNDA 0.017447f
C2786 VDDA.n1714 GNDA 0.017447f
C2787 VDDA.n1716 GNDA 0.016824f
C2788 VDDA.n1718 GNDA 0.015577f
C2789 VDDA.n1719 GNDA 0.015577f
C2790 VDDA.n1720 GNDA 0.015577f
C2791 VDDA.n1721 GNDA 0.015577f
C2792 VDDA.n1722 GNDA 0.016824f
C2793 VDDA.n1723 GNDA 0.016824f
C2794 VDDA.n1724 GNDA 0.016824f
C2795 VDDA.n1726 GNDA 0.017447f
C2796 VDDA.n1728 GNDA 0.017447f
C2797 VDDA.n1729 GNDA 0.017447f
C2798 VDDA.n1730 GNDA 0.017447f
C2799 VDDA.n1731 GNDA 0.016824f
C2800 VDDA.n1732 GNDA 0.015577f
C2801 VDDA.n1733 GNDA 0.015577f
C2802 VDDA.n1734 GNDA 0.015577f
C2803 VDDA.n1736 GNDA 0.015577f
C2804 VDDA.n1738 GNDA 0.016824f
C2805 VDDA.n1739 GNDA 0.016824f
C2806 VDDA.n1740 GNDA 0.016824f
C2807 VDDA.n1741 GNDA 0.017447f
C2808 VDDA.n1742 GNDA 0.017447f
C2809 VDDA.n1743 GNDA 0.017447f
C2810 VDDA.n1744 GNDA 0.017447f
C2811 VDDA.n1746 GNDA 0.016824f
C2812 VDDA.n1748 GNDA 0.015577f
C2813 VDDA.n1749 GNDA 0.015577f
C2814 VDDA.n1750 GNDA 0.015577f
C2815 VDDA.n1751 GNDA 0.015577f
C2816 VDDA.n1752 GNDA 0.016824f
C2817 VDDA.n1753 GNDA 0.016824f
C2818 VDDA.n1754 GNDA 0.016824f
C2819 VDDA.n1756 GNDA 0.017447f
C2820 VDDA.n1758 GNDA 0.017447f
C2821 VDDA.n1760 GNDA 0.016824f
C2822 VDDA.n1761 GNDA 0.016824f
C2823 VDDA.n1762 GNDA 0.016824f
C2824 VDDA.n1763 GNDA 0.011839f
C2825 VDDA.n1764 GNDA 0.058863f
C2826 VDDA.n1765 GNDA 0.028615f
C2827 VDDA.n1766 GNDA 0.012288f
C2828 VDDA.t258 GNDA 0.011428f
C2829 VDDA.n1775 GNDA 0.038361f
C2830 VDDA.t256 GNDA 0.031859f
C2831 VDDA.t31 GNDA 0.028608f
C2832 VDDA.t300 GNDA 0.031859f
C2833 VDDA.t301 GNDA 0.011428f
C2834 VDDA.n1783 GNDA 0.038361f
C2835 VDDA.n1787 GNDA 0.012197f
C2836 VDDA.n1788 GNDA 0.030485f
C2837 VDDA.n1789 GNDA 0.034036f
C2838 VDDA.n1903 GNDA 0.022051f
C2839 VDDA.n1906 GNDA 11.7728f
C2840 VDDA.n1909 GNDA 0.018205f
C2841 VDDA.n1911 GNDA 0.017555f
C2842 VDDA.n1913 GNDA 0.016255f
C2843 VDDA.n1915 GNDA 0.018205f
C2844 VDDA.n1917 GNDA 0.017555f
C2845 VDDA.n1919 GNDA 0.016255f
C2846 VDDA.n1921 GNDA 0.018205f
C2847 VDDA.n1923 GNDA 0.017555f
C2848 VDDA.n1925 GNDA 0.016255f
C2849 VDDA.n1927 GNDA 0.018205f
C2850 VDDA.n1929 GNDA 0.017555f
C2851 VDDA.n1932 GNDA 0.010305f
C2852 VDDA.n1934 GNDA 0.010305f
C2853 VDDA.n1936 GNDA 0.010305f
C2854 VDDA.n1938 GNDA 0.010403f
C2855 VDDA.t422 GNDA 0.256028f
C2856 VDDA.t424 GNDA 0.256028f
C2857 VDDA.t421 GNDA 0.243239f
C2858 VDDA.n1939 GNDA 0.47078f
C2859 VDDA.n1940 GNDA 0.248571f
C2860 VDDA.t423 GNDA 0.240274f
C2861 VDDA.n1941 GNDA 0.312969f
C2862 VDDA.n1942 GNDA 0.161948f
C2863 VDDA.n1943 GNDA 0.010305f
C2864 VDDA.n1944 GNDA 0.010403f
C2865 VDDA.n1945 GNDA 0.010403f
C2866 VDDA.n1947 GNDA 0.105331f
C2867 VDDA.n1948 GNDA 0.105331f
C2868 VDDA.n1950 GNDA 0.053169f
C2869 VDDA.n1953 GNDA 0.053169f
C2870 VDDA.n1955 GNDA 0.053169f
C2871 VDDA.n1957 GNDA 0.053169f
C2872 VDDA.n1959 GNDA 0.053169f
C2873 VDDA.n1961 GNDA 0.053169f
C2874 VDDA.n1963 GNDA 0.053169f
C2875 VDDA.n1965 GNDA 0.053169f
C2876 VDDA.n1967 GNDA 0.053169f
C2877 VDDA.n1969 GNDA 0.053169f
C2878 VDDA.n1973 GNDA 0.053169f
C2879 VDDA.n1975 GNDA 0.053169f
C2880 VDDA.n1977 GNDA 0.053169f
C2881 VDDA.n1979 GNDA 0.053169f
C2882 VDDA.n1981 GNDA 0.053169f
C2883 VDDA.n1983 GNDA 0.053169f
C2884 VDDA.n1985 GNDA 0.053169f
C2885 VDDA.n1987 GNDA 0.085609f
C2886 VDDA.n1990 GNDA 0.014509f
C2887 VDDA.n1991 GNDA 0.026716f
C2888 VDDA.t327 GNDA 0.022492f
C2889 VDDA.t9 GNDA 0.018205f
C2890 VDDA.t172 GNDA 0.018205f
C2891 VDDA.t57 GNDA 0.018205f
C2892 VDDA.t131 GNDA 0.018205f
C2893 VDDA.t365 GNDA 0.018205f
C2894 VDDA.t139 GNDA 0.018205f
C2895 VDDA.t163 GNDA 0.018205f
C2896 VDDA.t11 GNDA 0.018205f
C2897 VDDA.t122 GNDA 0.018205f
C2898 VDDA.t170 GNDA 0.018205f
C2899 VDDA.t141 GNDA 0.018205f
C2900 VDDA.t37 GNDA 0.018205f
C2901 VDDA.t186 GNDA 0.018205f
C2902 VDDA.t143 GNDA 0.018205f
C2903 VDDA.t133 GNDA 0.018205f
C2904 VDDA.t55 GNDA 0.018205f
C2905 VDDA.t15 GNDA 0.018205f
C2906 VDDA.t161 GNDA 0.018205f
C2907 VDDA.t243 GNDA 0.027242f
C2908 VDDA.n1992 GNDA 0.021966f
C2909 VDDA.n1993 GNDA 0.01445f
C2910 VDDA.n1995 GNDA 0.069215f
C2911 VDDA.n1996 GNDA 0.069215f
C2912 VDDA.n1998 GNDA 0.03954f
C2913 VDDA.t333 GNDA 0.02777f
C2914 VDDA.t51 GNDA 0.018205f
C2915 VDDA.t361 GNDA 0.018205f
C2916 VDDA.t359 GNDA 0.018205f
C2917 VDDA.t0 GNDA 0.018205f
C2918 VDDA.t157 GNDA 0.018205f
C2919 VDDA.t368 GNDA 0.018205f
C2920 VDDA.t77 GNDA 0.018205f
C2921 VDDA.t69 GNDA 0.018205f
C2922 VDDA.t79 GNDA 0.018205f
C2923 VDDA.t64 GNDA 0.018205f
C2924 VDDA.t194 GNDA 0.018205f
C2925 VDDA.t190 GNDA 0.018205f
C2926 VDDA.t184 GNDA 0.018205f
C2927 VDDA.t188 GNDA 0.018205f
C2928 VDDA.t4 GNDA 0.018205f
C2929 VDDA.t192 GNDA 0.018205f
C2930 VDDA.t7 GNDA 0.018205f
C2931 VDDA.t198 GNDA 0.018205f
C2932 VDDA.t291 GNDA 0.027242f
C2933 VDDA.n1999 GNDA 0.021966f
C2934 VDDA.n2000 GNDA 0.01445f
C2935 VDDA.n2002 GNDA 0.126432f
C2936 VDDA.n2003 GNDA 0.10403f
C2937 VDDA.n2005 GNDA 0.010403f
C2938 VDDA.n2006 GNDA 0.010403f
C2939 VDDA.n2008 GNDA 0.087776f
C2940 VDDA.n2009 GNDA 0.087776f
C2941 VDDA.t293 GNDA 0.031004f
C2942 VDDA.n2010 GNDA 0.011885f
C2943 VDDA.n2011 GNDA 0.025298f
C2944 VDDA.n2012 GNDA 0.025298f
C2945 VDDA.n2013 GNDA 0.025298f
C2946 VDDA.n2014 GNDA 0.025298f
C2947 VDDA.n2015 GNDA 0.025298f
C2948 VDDA.n2016 GNDA 0.025298f
C2949 VDDA.n2017 GNDA 0.025298f
C2950 VDDA.n2018 GNDA 0.025298f
C2951 VDDA.n2044 GNDA 0.060793f
C2952 VDDA.t294 GNDA 0.064477f
C2953 VDDA.t414 GNDA 0.066319f
C2954 VDDA.t416 GNDA 0.066319f
C2955 VDDA.t17 GNDA 0.066319f
C2956 VDDA.t404 GNDA 0.066319f
C2957 VDDA.t126 GNDA 0.066319f
C2958 VDDA.t135 GNDA 0.066319f
C2959 VDDA.t137 GNDA 0.066319f
C2960 VDDA.t92 GNDA 0.066319f
C2961 VDDA.t389 GNDA 0.066319f
C2962 VDDA.t392 GNDA 0.066319f
C2963 VDDA.t19 GNDA 0.066319f
C2964 VDDA.t60 GNDA 0.066319f
C2965 VDDA.t88 GNDA 0.066319f
C2966 VDDA.t104 GNDA 0.066319f
C2967 VDDA.t418 GNDA 0.066319f
C2968 VDDA.t373 GNDA 0.066319f
C2969 VDDA.t266 GNDA 0.064477f
C2970 VDDA.n2061 GNDA 0.060793f
C2971 VDDA.t265 GNDA 0.031004f
C2972 VDDA.n2064 GNDA 0.012522f
C2973 VDDA.n2065 GNDA 0.123905f
C2974 VDDA.n2066 GNDA 0.086968f
C2975 VDDA.n2067 GNDA 0.086968f
C2976 VDDA.n2068 GNDA 0.086968f
C2977 VDDA.n2069 GNDA 0.086968f
C2978 VDDA.n2070 GNDA 0.086968f
C2979 VDDA.n2071 GNDA 0.086968f
C2980 VDDA.n2072 GNDA 0.086968f
C2981 VDDA.n2073 GNDA 0.073335f
C2982 VDDA.n2074 GNDA 0.083621f
C2983 VDDA.n2076 GNDA 0.039775f
C2984 VDDA.t272 GNDA 0.026878f
C2985 VDDA.t84 GNDA 0.016688f
C2986 VDDA.t396 GNDA 0.016688f
C2987 VDDA.t336 GNDA 0.026299f
C2988 VDDA.n2077 GNDA 0.037977f
C2989 VDDA.n2079 GNDA 0.143438f
C2990 VDDA.n2080 GNDA 0.105981f
C2991 VDDA.n2082 GNDA 0.010403f
C2992 VDDA.n2083 GNDA 0.010403f
C2993 VDDA.n2085 GNDA 0.041612f
C2994 VDDA.n2086 GNDA 0.041612f
C2995 VDDA.n2089 GNDA 0.037768f
C2996 VDDA.t246 GNDA 0.026297f
C2997 VDDA.t182 GNDA 0.016688f
C2998 VDDA.t112 GNDA 0.016688f
C2999 VDDA.t285 GNDA 0.026297f
C3000 VDDA.n2090 GNDA 0.037768f
C3001 VDDA.n2095 GNDA 0.02256f
C3002 VDDA.t303 GNDA 0.023775f
C3003 VDDA.t33 GNDA 0.016688f
C3004 VDDA.t174 GNDA 0.016688f
C3005 VDDA.t45 GNDA 0.016688f
C3006 VDDA.t39 GNDA 0.016688f
C3007 VDDA.t275 GNDA 0.023775f
C3008 VDDA.n2096 GNDA 0.02256f
C3009 VDDA.n2104 GNDA 0.037768f
C3010 VDDA.t342 GNDA 0.026297f
C3011 VDDA.t159 GNDA 0.016688f
C3012 VDDA.t176 GNDA 0.016688f
C3013 VDDA.t155 GNDA 0.016688f
C3014 VDDA.t377 GNDA 0.016688f
C3015 VDDA.t394 GNDA 0.016688f
C3016 VDDA.t370 GNDA 0.016688f
C3017 VDDA.t43 GNDA 0.016688f
C3018 VDDA.t110 GNDA 0.016688f
C3019 VDDA.t252 GNDA 0.026297f
C3020 VDDA.n2105 GNDA 0.037768f
C3021 VDDA.n2110 GNDA 0.022564f
C3022 VDDA.t312 GNDA 0.023775f
C3023 VDDA.t108 GNDA 0.016688f
C3024 VDDA.t407 GNDA 0.016688f
C3025 VDDA.t2 GNDA 0.016688f
C3026 VDDA.t178 GNDA 0.016688f
C3027 VDDA.t354 GNDA 0.023775f
C3028 VDDA.n2111 GNDA 0.022564f
C3029 VDDA.n2113 GNDA 0.076379f
C3030 VDDA.n2114 GNDA 0.048204f
C3031 VDDA.n2115 GNDA 0.059681f
C3032 VDDA.n2116 GNDA 0.053829f
C3033 VDDA.n2117 GNDA 0.042364f
C3034 VDDA.n2118 GNDA 0.048215f
C3035 VDDA.n2119 GNDA 0.048215f
C3036 VDDA.n2120 GNDA 0.048215f
C3037 VDDA.n2121 GNDA 0.042364f
C3038 VDDA.n2122 GNDA 0.053829f
C3039 VDDA.n2123 GNDA 0.059681f
C3040 VDDA.n2124 GNDA 0.048202f
C3041 VDDA.n2125 GNDA 0.048202f
C3042 VDDA.n2126 GNDA 0.059681f
C3043 VDDA.n2127 GNDA 0.060982f
C3044 VDDA.n2128 GNDA 0.050816f
C3045 VDDA.n2129 GNDA 0.116248f
C3046 VDDA.n2130 GNDA 0.096878f
C3047 VDDA.n2132 GNDA 0.010403f
C3048 VDDA.n2133 GNDA 0.010403f
C3049 VDDA.n2135 GNDA 0.039662f
C3050 VDDA.n2136 GNDA 0.042912f
C3051 VDDA.n2140 GNDA 0.017555f
C3052 VDDA.n2141 GNDA 0.018205f
C3053 VDDA.n2142 GNDA 0.018205f
C3054 VDDA.n2150 GNDA 0.016255f
C3055 VDDA.n2151 GNDA 0.016255f
C3056 VDDA.n2152 GNDA 0.017555f
C3057 VDDA.n2160 GNDA 0.018205f
C3058 VDDA.n2161 GNDA 0.017555f
C3059 VDDA.n2162 GNDA 0.016255f
C3060 VDDA.n2170 GNDA 0.017555f
C3061 VDDA.n2171 GNDA 0.018205f
C3062 VDDA.n2172 GNDA 0.018205f
C3063 VDDA.n2180 GNDA 0.016255f
C3064 VDDA.n2181 GNDA 0.016255f
C3065 VDDA.n2182 GNDA 0.017555f
C3066 VDDA.n2190 GNDA 0.018205f
C3067 VDDA.n2191 GNDA 0.017555f
C3068 VDDA.n2192 GNDA 0.016255f
C3069 VDDA.n2200 GNDA 0.017555f
C3070 VDDA.n2201 GNDA 0.018205f
C3071 VDDA.n2202 GNDA 0.018205f
C3072 VDDA.n2210 GNDA 0.016255f
C3073 VDDA.n2211 GNDA 0.016255f
C3074 VDDA.n2212 GNDA 0.017555f
C3075 VDDA.n2220 GNDA 0.018205f
C3076 VDDA.n2221 GNDA 0.017555f
C3077 VDDA.n2222 GNDA 0.016255f
C3078 VDDA.n2230 GNDA 0.017555f
C3079 VDDA.n2231 GNDA 0.018205f
C3080 VDDA.n2232 GNDA 0.018205f
C3081 VDDA.n2240 GNDA 0.016255f
C3082 VDDA.n2241 GNDA 0.016255f
C3083 VDDA.n2242 GNDA 0.017555f
C3084 VDDA.n2250 GNDA 0.050713f
C3085 VDDA.n2253 GNDA 13.6106f
C3086 VDDA.n2254 GNDA 4.64669f
C3087 VDDA.n2257 GNDA 0.278281f
C3088 VDDA.n2258 GNDA 0.27503f
C3089 VDDA.n2260 GNDA 0.085825f
C3090 VDDA.n2261 GNDA 0.010403f
C3091 VDDA.n2262 GNDA 0.066319f
C3092 VDDA.n2263 GNDA 0.112901f
C3093 VDDA.t281 GNDA 0.013301f
C3094 VDDA.t349 GNDA 0.026983f
C3095 VDDA.n2264 GNDA 0.078275f
C3096 VDDA.t348 GNDA 0.064659f
C3097 VDDA.t224 GNDA 0.050715f
C3098 VDDA.t230 GNDA 0.050715f
C3099 VDDA.t218 GNDA 0.050715f
C3100 VDDA.t214 GNDA 0.050715f
C3101 VDDA.t210 GNDA 0.050715f
C3102 VDDA.t204 GNDA 0.050715f
C3103 VDDA.t238 GNDA 0.050715f
C3104 VDDA.t226 GNDA 0.050715f
C3105 VDDA.t216 GNDA 0.050715f
C3106 VDDA.t212 GNDA 0.050715f
C3107 VDDA.t282 GNDA 0.064659f
C3108 VDDA.t283 GNDA 0.026983f
C3109 VDDA.n2265 GNDA 0.078275f
C3110 VDDA.n2266 GNDA 0.029046f
C3111 VDDA.n2267 GNDA 0.027711f
C3112 VDDA.n2268 GNDA 0.018957f
C3113 VDDA.n2269 GNDA 0.055722f
C3114 VDDA.n2270 GNDA 0.018957f
C3115 VDDA.n2271 GNDA 0.051155f
C3116 VDDA.n2272 GNDA 0.015979f
C3117 VDDA.n2273 GNDA 0.065635f
C3118 VDDA.n2275 GNDA 0.018957f
C3119 VDDA.n2276 GNDA 0.051155f
C3120 VDDA.n2277 GNDA 0.018957f
C3121 VDDA.n2278 GNDA 0.055722f
C3122 VDDA.n2279 GNDA 0.027711f
C3123 VDDA.n2280 GNDA 0.081042f
C3124 VDDA.n2281 GNDA 0.010403f
C3125 VDDA.n2282 GNDA 0.010403f
C3126 VDDA.n2283 GNDA 0.010305f
C3127 VDDA.n2285 GNDA 0.03446f
C3128 VDDA.n2286 GNDA 0.120285f
C3129 VDDA.n2287 GNDA 0.010403f
C3130 VDDA.t87 GNDA 0.013004f
C3131 VDDA.t401 GNDA 0.013004f
C3132 VDDA.n2288 GNDA 0.033462f
C3133 VDDA.n2289 GNDA 0.114131f
C3134 VDDA.t307 GNDA 0.045764f
C3135 VDDA.t100 GNDA 0.013004f
C3136 VDDA.t376 GNDA 0.013004f
C3137 VDDA.n2290 GNDA 0.033462f
C3138 VDDA.n2291 GNDA 0.114131f
C3139 VDDA.t28 GNDA 0.013004f
C3140 VDDA.t72 GNDA 0.013004f
C3141 VDDA.n2292 GNDA 0.033462f
C3142 VDDA.n2293 GNDA 0.114131f
C3143 VDDA.t49 GNDA 0.013004f
C3144 VDDA.t98 GNDA 0.013004f
C3145 VDDA.n2294 GNDA 0.033462f
C3146 VDDA.n2295 GNDA 0.114131f
C3147 VDDA.t154 GNDA 0.013004f
C3148 VDDA.t150 GNDA 0.013004f
C3149 VDDA.n2296 GNDA 0.033462f
C3150 VDDA.n2297 GNDA 0.134441f
C3151 VDDA.t305 GNDA 0.015777f
C3152 VDDA.n2298 GNDA 0.042161f
C3153 VDDA.n2299 GNDA 0.153083f
C3154 VDDA.t306 GNDA 0.099148f
C3155 VDDA.t153 GNDA 0.076289f
C3156 VDDA.t149 GNDA 0.075806f
C3157 VDDA.t48 GNDA 0.075254f
C3158 VDDA.t97 GNDA 0.076289f
C3159 VDDA.t27 GNDA 0.076289f
C3160 VDDA.t71 GNDA 0.076289f
C3161 VDDA.t99 GNDA 0.076289f
C3162 VDDA.t375 GNDA 0.076289f
C3163 VDDA.t86 GNDA 0.076289f
C3164 VDDA.t400 GNDA 0.076289f
C3165 VDDA.t318 GNDA 0.099148f
C3166 VDDA.t319 GNDA 0.045764f
C3167 VDDA.n2300 GNDA 0.153083f
C3168 VDDA.t317 GNDA 0.015777f
C3169 VDDA.n2301 GNDA 0.040896f
C3170 VDDA.n2302 GNDA 0.049534f
C3171 VDDA.n2304 GNDA 0.010403f
C3172 VDDA.n2305 GNDA 0.010403f
C3173 VDDA.n2307 GNDA 0.010403f
C3174 VDDA.n2308 GNDA 0.010403f
C3175 VDDA.n2309 GNDA 0.018342f
C3176 VDDA.n2310 GNDA 0.018059f
C3177 VDDA.n2311 GNDA 0.14175f
C3178 VDDA.n2312 GNDA 0.018059f
C3179 VDDA.n2313 GNDA 0.075568f
C3180 VDDA.n2314 GNDA 0.018059f
C3181 VDDA.n2315 GNDA 0.075568f
C3182 VDDA.n2316 GNDA 0.018059f
C3183 VDDA.n2317 GNDA 0.075568f
C3184 VDDA.n2318 GNDA 0.018059f
C3185 VDDA.n2319 GNDA 0.101576f
C3186 VDDA.n2320 GNDA 0.045513f
C3187 VDDA.n2321 GNDA 0.010305f
C3188 VDDA.n2322 GNDA 0.010403f
C3189 VDDA.n2324 GNDA 0.13849f
C3190 VDDA.n2325 GNDA 0.056318f
C3191 VDDA.t316 GNDA 0.015464f
C3192 VDDA.n2326 GNDA 0.047508f
C3193 VDDA.t315 GNDA 0.038526f
C3194 VDDA.t165 GNDA 0.028608f
C3195 VDDA.t130 GNDA 0.028608f
C3196 VDDA.t23 GNDA 0.028608f
C3197 VDDA.t54 GNDA 0.028608f
C3198 VDDA.t106 GNDA 0.028608f
C3199 VDDA.t166 GNDA 0.028608f
C3200 VDDA.t53 GNDA 0.028608f
C3201 VDDA.t402 GNDA 0.028608f
C3202 VDDA.t403 GNDA 0.028608f
C3203 VDDA.t399 GNDA 0.028608f
C3204 VDDA.t321 GNDA 0.038526f
C3205 VDDA.t322 GNDA 0.015464f
C3206 VDDA.n2327 GNDA 0.047508f
C3207 VDDA.n2328 GNDA 0.034052f
C3208 VDDA.n2329 GNDA 0.197651f
C3209 VDDA.n2330 GNDA 0.038361f
C3210 VDDA.n2332 GNDA 0.13849f
C3211 VDDA.n2333 GNDA 0.010305f
C3212 VDDA.n2335 GNDA 0.146943f
C3213 VDDA.n2336 GNDA 0.146943f
C3214 VDDA.n2338 GNDA 0.038361f
C3215 VDDA.n2340 GNDA 0.120285f
C3216 VDDA.n2342 GNDA 0.121585f
C3217 VDDA.t364 GNDA 0.034568f
C3218 VDDA.t41 GNDA 0.034568f
C3219 VDDA.t66 GNDA 0.034568f
C3220 VDDA.t68 GNDA 0.034568f
C3221 VDDA.t249 GNDA 0.038497f
C3222 VDDA.n2352 GNDA 0.046353f
C3223 VDDA.n2355 GNDA 0.016255f
C3224 VDDA.n2357 GNDA 0.01204f
C3225 VDDA.n2358 GNDA 0.146807f
C3226 VDDA.n2359 GNDA 0.018864f
C3227 VDDA.n2360 GNDA 0.064144f
C3228 VDDA.n2361 GNDA 0.040826f
C3229 VDDA.n2362 GNDA 0.040826f
C3230 VDDA.n2363 GNDA 0.011823f
C3231 VDDA.n2366 GNDA 0.01192f
C3232 VDDA.n2369 GNDA 0.01192f
C3233 VDDA.n2370 GNDA 0.01192f
C3234 VDDA.n2372 GNDA 0.016255f
C3235 VDDA.n2373 GNDA 0.011699f
C3236 VDDA.n2375 GNDA 0.016255f
C3237 VDDA.n2378 GNDA 0.042425f
C3238 VDDA.t345 GNDA 0.038497f
C3239 VDDA.t363 GNDA 0.034568f
C3240 VDDA.t397 GNDA 0.034568f
C3241 VDDA.t180 GNDA 0.034568f
C3242 VDDA.t24 GNDA 0.034568f
C3243 VDDA.t351 GNDA 0.038497f
C3244 VDDA.n2386 GNDA 0.046353f
C3245 VDDA.n2389 GNDA 0.01204f
C3246 VDDA.n2390 GNDA 0.146807f
C3247 VDDA.n2391 GNDA 0.121585f
C3248 VDDA.n2392 GNDA 0.146943f
C3249 VDDA.n2393 GNDA 0.038361f
C3250 VDDA.n2395 GNDA 0.120285f
C3251 VDDA.n2396 GNDA 0.120285f
C3252 VDDA.n2398 GNDA 0.169699f
C3253 VDDA.n2399 GNDA 0.010403f
C3254 VDDA.n2400 GNDA 0.03446f
C3255 VDDA.n2401 GNDA 0.081042f
C3256 VDDA.t308 GNDA 0.013301f
C3257 VDDA.t261 GNDA 0.026983f
C3258 VDDA.n2402 GNDA 0.078275f
C3259 VDDA.t260 GNDA 0.064659f
C3260 VDDA.t240 GNDA 0.050715f
C3261 VDDA.t228 GNDA 0.050715f
C3262 VDDA.t234 GNDA 0.050715f
C3263 VDDA.t222 GNDA 0.050715f
C3264 VDDA.t206 GNDA 0.050715f
C3265 VDDA.t202 GNDA 0.050715f
C3266 VDDA.t236 GNDA 0.050715f
C3267 VDDA.t200 GNDA 0.050715f
C3268 VDDA.t232 GNDA 0.050715f
C3269 VDDA.t220 GNDA 0.050715f
C3270 VDDA.t309 GNDA 0.064659f
C3271 VDDA.t310 GNDA 0.026983f
C3272 VDDA.n2403 GNDA 0.078275f
C3273 VDDA.n2404 GNDA 0.029046f
C3274 VDDA.n2405 GNDA 0.027711f
C3275 VDDA.n2406 GNDA 0.018957f
C3276 VDDA.n2407 GNDA 0.055722f
C3277 VDDA.n2408 GNDA 0.018957f
C3278 VDDA.n2409 GNDA 0.051155f
C3279 VDDA.n2410 GNDA 0.015979f
C3280 VDDA.n2411 GNDA 0.065635f
C3281 VDDA.n2413 GNDA 0.018957f
C3282 VDDA.n2414 GNDA 0.051155f
C3283 VDDA.n2415 GNDA 0.018957f
C3284 VDDA.n2416 GNDA 0.055722f
C3285 VDDA.n2417 GNDA 0.027711f
C3286 VDDA.n2418 GNDA 0.112901f
C3287 VDDA.n2419 GNDA 0.010403f
C3288 VDDA.n2420 GNDA 0.017555f
C3289 VDDA.n2424 GNDA 0.016255f
C3290 VDDA.n2428 GNDA 0.018205f
C3291 VDDA.n2432 GNDA 0.017555f
C3292 VDDA.n2436 GNDA 0.016255f
C3293 VDDA.n2440 GNDA 0.018205f
C3294 VDDA.n2444 GNDA 0.017555f
C3295 VDDA.n2448 GNDA 0.016255f
C3296 VDDA.n2452 GNDA 0.018205f
C3297 VDDA.n2456 GNDA 0.017555f
C3298 VDDA.n2460 GNDA 0.016255f
C3299 VDDA.n2464 GNDA 0.050713f
C3300 VDDA.n2475 GNDA 0.018205f
C3301 VDDA.n2476 GNDA 0.017555f
C3302 VDDA.n2477 GNDA 0.016255f
C3303 VDDA.n2485 GNDA 0.017555f
C3304 VDDA.n2486 GNDA 0.018205f
C3305 VDDA.n2487 GNDA 0.018205f
C3306 VDDA.n2495 GNDA 0.016255f
C3307 VDDA.n2496 GNDA 0.016255f
C3308 VDDA.n2497 GNDA 0.017555f
C3309 VDDA.n2505 GNDA 0.018205f
C3310 VDDA.n2506 GNDA 0.017555f
C3311 VDDA.n2507 GNDA 0.016255f
C3312 VDDA.n2515 GNDA 0.017555f
C3313 VDDA.n2516 GNDA 0.018205f
C3314 VDDA.n2517 GNDA 0.018205f
C3315 VDDA.n2525 GNDA 0.016255f
C3316 VDDA.n2526 GNDA 0.016255f
C3317 VDDA.n2527 GNDA 0.017555f
C3318 VDDA.n2535 GNDA 0.018205f
C3319 VDDA.n2536 GNDA 0.017555f
C3320 VDDA.n2537 GNDA 0.016255f
C3321 VDDA.n2545 GNDA 0.017555f
C3322 VDDA.n2546 GNDA 0.018205f
C3323 VDDA.n2547 GNDA 0.018205f
C3324 VDDA.n2555 GNDA 0.016255f
C3325 VDDA.n2556 GNDA 0.016255f
C3326 VDDA.n2557 GNDA 0.017555f
C3327 VDDA.n2565 GNDA 0.018205f
C3328 VDDA.n2566 GNDA 0.017555f
C3329 VDDA.n2567 GNDA 0.016255f
C3330 VDDA.n2575 GNDA 0.017555f
C3331 VDDA.n2576 GNDA 0.018205f
C3332 VDDA.n2577 GNDA 0.018205f
C3333 VDDA.n2584 GNDA 0.278281f
C3334 VDDA.n2585 GNDA 0.27503f
C3335 VDDA.n2587 GNDA 0.066319f
C3336 VDDA.n2588 GNDA 0.010403f
C3337 VDDA.n2589 GNDA 0.085825f
C3338 VDDA.n2590 GNDA 0.010403f
C3339 VDDA.n2591 GNDA 0.085825f
C3340 VDDA.n2592 GNDA 0.010403f
C3341 VDDA.n2594 GNDA 0.27503f
C3342 VDDA.n2595 GNDA 0.278281f
C3343 VDDA.n2598 GNDA 3.64106f
C3344 VDDA.n2624 GNDA 0.016255f
C3345 VDDA.n2628 GNDA 0.018205f
C3346 VDDA.n2632 GNDA 0.017555f
C3347 VDDA.n2636 GNDA 0.016255f
C3348 VDDA.n2640 GNDA 0.018205f
C3349 VDDA.n2644 GNDA 0.017555f
C3350 VDDA.n2648 GNDA 0.016255f
C3351 VDDA.n2652 GNDA 0.018205f
C3352 VDDA.n2656 GNDA 0.017555f
C3353 VDDA.n2660 GNDA 0.016255f
C3354 VDDA.n2664 GNDA 0.050713f
C3355 VDDA.n2672 GNDA 0.018205f
C3356 VDDA.n2673 GNDA 0.017555f
C3357 VDDA.n2674 GNDA 0.016255f
C3358 VDDA.n2680 GNDA 0.017555f
C3359 VDDA.n2681 GNDA 0.018205f
C3360 VDDA.n2682 GNDA 0.018205f
C3361 VDDA.n2688 GNDA 0.016255f
C3362 VDDA.n2689 GNDA 0.016255f
C3363 VDDA.n2690 GNDA 0.017555f
C3364 VDDA.n2696 GNDA 0.018205f
C3365 VDDA.n2697 GNDA 0.017555f
C3366 VDDA.n2698 GNDA 0.016255f
C3367 VDDA.n2704 GNDA 0.017555f
C3368 VDDA.n2705 GNDA 0.018205f
C3369 VDDA.n2706 GNDA 0.018205f
C3370 VDDA.n2712 GNDA 0.016255f
C3371 VDDA.n2713 GNDA 0.016255f
C3372 VDDA.n2714 GNDA 0.017555f
C3373 VDDA.n2720 GNDA 0.018205f
C3374 VDDA.n2721 GNDA 0.017555f
C3375 VDDA.n2722 GNDA 0.016255f
C3376 VDDA.n2728 GNDA 0.017555f
C3377 VDDA.n2729 GNDA 0.018205f
C3378 VDDA.n2730 GNDA 0.018205f
C3379 VDDA.n2736 GNDA 0.016255f
C3380 VDDA.n2737 GNDA 0.016255f
C3381 VDDA.n2738 GNDA 0.017555f
C3382 VDDA.n2744 GNDA 0.018205f
C3383 VDDA.n2745 GNDA 0.017555f
C3384 VDDA.n2746 GNDA 0.016255f
C3385 VDDA.n2752 GNDA 0.017555f
C3386 VDDA.n2753 GNDA 0.018205f
C3387 VDDA.n2754 GNDA 0.018205f
C3388 VDDA.n2758 GNDA 2.42737f
C3389 VDDA.n2761 GNDA 0.278281f
C3390 VDDA.n2762 GNDA 0.27503f
C3391 VDDA.n2764 GNDA 0.040312f
C3392 VDDA.n2765 GNDA 0.010403f
C3393 VDDA.n2766 GNDA 0.040312f
C3394 VDDA.n2767 GNDA 0.010403f
C3395 VDDA.n2768 GNDA 0.017555f
C3396 VDDA.n2772 GNDA 0.016255f
C3397 VDDA.n2776 GNDA 0.018205f
C3398 VDDA.n2780 GNDA 0.017555f
C3399 VDDA.n2784 GNDA 0.016255f
C3400 VDDA.n2788 GNDA 0.018205f
C3401 VDDA.n2792 GNDA 0.017555f
C3402 VDDA.n2796 GNDA 0.016255f
C3403 VDDA.n2800 GNDA 0.018205f
C3404 VDDA.n2804 GNDA 0.017555f
C3405 VDDA.n2808 GNDA 0.016255f
C3406 VDDA.n2812 GNDA 0.050713f
C3407 VDDA.n2823 GNDA 0.018205f
C3408 VDDA.n2824 GNDA 0.017555f
C3409 VDDA.n2825 GNDA 0.016255f
C3410 VDDA.n2833 GNDA 0.017555f
C3411 VDDA.n2834 GNDA 0.018205f
C3412 VDDA.n2835 GNDA 0.018205f
C3413 VDDA.n2843 GNDA 0.016255f
C3414 VDDA.n2844 GNDA 0.016255f
C3415 VDDA.n2845 GNDA 0.017555f
C3416 VDDA.n2853 GNDA 0.018205f
C3417 VDDA.n2854 GNDA 0.017555f
C3418 VDDA.n2855 GNDA 0.016255f
C3419 VDDA.n2863 GNDA 0.017555f
C3420 VDDA.n2864 GNDA 0.018205f
C3421 VDDA.n2865 GNDA 0.018205f
C3422 VDDA.n2873 GNDA 0.016255f
C3423 VDDA.n2874 GNDA 0.016255f
C3424 VDDA.n2875 GNDA 0.017555f
C3425 VDDA.n2883 GNDA 0.018205f
C3426 VDDA.n2884 GNDA 0.017555f
C3427 VDDA.n2885 GNDA 0.016255f
C3428 VDDA.n2893 GNDA 0.017555f
C3429 VDDA.n2894 GNDA 0.018205f
C3430 VDDA.n2895 GNDA 0.018205f
C3431 VDDA.n2903 GNDA 0.016255f
C3432 VDDA.n2904 GNDA 0.016255f
C3433 VDDA.n2905 GNDA 0.017555f
C3434 VDDA.n2913 GNDA 0.018205f
C3435 VDDA.n2914 GNDA 0.017555f
C3436 VDDA.n2915 GNDA 0.016255f
C3437 VDDA.n2923 GNDA 0.017555f
C3438 VDDA.n2924 GNDA 0.018205f
C3439 VDDA.n2925 GNDA 0.018205f
C3440 VDDA.n2932 GNDA 0.278281f
C3441 VDDA.n2933 GNDA 0.27503f
C3442 VDDA.n2935 GNDA 0.040312f
C3443 VDDA.n2936 GNDA 0.010403f
C3444 VDDA.n2937 GNDA 0.040312f
C3445 VDDA.n2938 GNDA 0.040312f
C3446 VDDA.n2939 GNDA 0.010403f
C3447 VDDA.n2940 GNDA 0.010403f
C3448 VDDA.n2942 GNDA 0.27503f
C3449 VDDA.n2943 GNDA 0.278281f
C3450 VDDA.n2946 GNDA 6.90068f
C3451 VDDA.n2947 GNDA 0.658859f
C3452 VDDA.n2948 GNDA 0.728212f
C3453 VDDA.n2949 GNDA 0.658859f
C3454 VDDA.n2950 GNDA 0.728212f
C3455 VDDA.n2951 GNDA 0.658859f
C3456 VDDA.n2952 GNDA 0.728212f
C3457 VDDA.n2953 GNDA 0.658859f
C3458 VDDA.n2954 GNDA 0.728212f
C3459 VDDA.n2955 GNDA 0.658859f
C3460 VDDA.n2956 GNDA 0.728212f
C3461 VDDA.n2957 GNDA 0.658859f
C3462 VDDA.n2958 GNDA 0.728212f
C3463 VDDA.n2959 GNDA 0.658859f
C3464 VDDA.n2960 GNDA 0.728212f
C3465 VDDA.n2961 GNDA 0.658859f
C3466 VDDA.n2962 GNDA 0.658859f
C3467 VDDA.n2964 GNDA 0.658859f
C3468 VDDA.n2967 GNDA 0.728212f
C3469 VDDA.n2970 GNDA 0.658859f
C3470 VDDA.n2973 GNDA 0.728212f
C3471 VDDA.n2976 GNDA 0.658859f
C3472 VDDA.n2979 GNDA 0.728212f
C3473 VDDA.n2982 GNDA 0.658859f
C3474 VDDA.n2985 GNDA 0.728212f
C3475 VDDA.n2988 GNDA 0.658859f
C3476 VDDA.n2991 GNDA 0.728212f
C3477 VDDA.n2994 GNDA 0.658859f
C3478 VDDA.n2997 GNDA 0.728212f
C3479 VDDA.n3000 GNDA 0.658859f
C3480 VDDA.n3003 GNDA 0.728212f
C3481 VDDA.n3006 GNDA 0.658859f
C3482 VDDA.n3009 GNDA 0.693535f
C3483 VDDA.n3010 GNDA 0.676197f
C3484 VDDA.n3011 GNDA 0.745551f
C3485 VDDA.n3012 GNDA 0.658859f
C3486 VDDA.n3013 GNDA 0.693535f
C3487 VDDA.n3014 GNDA 0.676197f
C3488 VDDA.n3015 GNDA 0.745551f
C3489 VDDA.n3016 GNDA 0.658859f
C3490 VDDA.n3017 GNDA 0.693535f
C3491 VDDA.n3018 GNDA 0.676197f
C3492 VDDA.n3019 GNDA 0.745551f
C3493 VDDA.n3020 GNDA 0.658859f
C3494 VDDA.n3021 GNDA 0.693535f
C3495 VDDA.n3022 GNDA 0.676197f
C3496 VDDA.n3023 GNDA 0.658859f
C3497 VDDA.n3026 GNDA 0.693535f
C3498 VDDA.n3028 GNDA 0.676197f
C3499 VDDA.n3030 GNDA 0.745551f
C3500 VDDA.n3032 GNDA 0.658859f
C3501 VDDA.n3034 GNDA 0.693535f
C3502 VDDA.n3036 GNDA 0.676197f
C3503 VDDA.n3038 GNDA 0.745551f
C3504 VDDA.n3040 GNDA 0.658859f
C3505 VDDA.n3042 GNDA 0.693535f
C3506 VDDA.n3044 GNDA 0.676197f
C3507 VDDA.n3046 GNDA 0.745551f
C3508 VDDA.n3048 GNDA 0.658859f
C3509 VDDA.n3050 GNDA 0.693535f
C3510 VDDA.n3051 GNDA 0.728212f
C3511 VDDA.n3052 GNDA 6.01642f
C3512 VDDA.n3053 GNDA 2.27133f
C3513 two_stage_opamp_dummy_magic_25_0.VD4.n0 GNDA 0.548627f
C3514 two_stage_opamp_dummy_magic_25_0.VD4.n1 GNDA 1.36659f
C3515 two_stage_opamp_dummy_magic_25_0.VD4.n2 GNDA 2.16604f
C3516 two_stage_opamp_dummy_magic_25_0.VD4.n3 GNDA 0.936914f
C3517 two_stage_opamp_dummy_magic_25_0.VD4.n4 GNDA 0.84648f
C3518 two_stage_opamp_dummy_magic_25_0.VD4.n5 GNDA 1.2192f
C3519 two_stage_opamp_dummy_magic_25_0.VD4.n6 GNDA 0.223288f
C3520 two_stage_opamp_dummy_magic_25_0.VD4.n7 GNDA 0.219626f
C3521 two_stage_opamp_dummy_magic_25_0.VD4.n8 GNDA 0.223288f
C3522 two_stage_opamp_dummy_magic_25_0.VD4.t12 GNDA 0.05484f
C3523 two_stage_opamp_dummy_magic_25_0.VD4.t36 GNDA 0.05484f
C3524 two_stage_opamp_dummy_magic_25_0.VD4.t16 GNDA 0.05484f
C3525 two_stage_opamp_dummy_magic_25_0.VD4.n9 GNDA 0.116347f
C3526 two_stage_opamp_dummy_magic_25_0.VD4.t4 GNDA 0.05484f
C3527 two_stage_opamp_dummy_magic_25_0.VD4.t6 GNDA 0.05484f
C3528 two_stage_opamp_dummy_magic_25_0.VD4.n10 GNDA 0.116347f
C3529 two_stage_opamp_dummy_magic_25_0.VD4.t14 GNDA 0.05484f
C3530 two_stage_opamp_dummy_magic_25_0.VD4.t8 GNDA 0.05484f
C3531 two_stage_opamp_dummy_magic_25_0.VD4.n11 GNDA 0.116347f
C3532 two_stage_opamp_dummy_magic_25_0.VD4.t37 GNDA 0.05484f
C3533 two_stage_opamp_dummy_magic_25_0.VD4.t21 GNDA 0.05484f
C3534 two_stage_opamp_dummy_magic_25_0.VD4.n12 GNDA 0.11218f
C3535 two_stage_opamp_dummy_magic_25_0.VD4.n13 GNDA 0.320708f
C3536 two_stage_opamp_dummy_magic_25_0.VD4.n14 GNDA 0.228605f
C3537 two_stage_opamp_dummy_magic_25_0.VD4.t28 GNDA 0.05484f
C3538 two_stage_opamp_dummy_magic_25_0.VD4.t20 GNDA 0.05484f
C3539 two_stage_opamp_dummy_magic_25_0.VD4.n15 GNDA 0.11218f
C3540 two_stage_opamp_dummy_magic_25_0.VD4.n16 GNDA 0.320077f
C3541 two_stage_opamp_dummy_magic_25_0.VD4.t23 GNDA 0.05484f
C3542 two_stage_opamp_dummy_magic_25_0.VD4.t22 GNDA 0.05484f
C3543 two_stage_opamp_dummy_magic_25_0.VD4.n17 GNDA 0.11218f
C3544 two_stage_opamp_dummy_magic_25_0.VD4.n18 GNDA 0.315749f
C3545 two_stage_opamp_dummy_magic_25_0.VD4.n19 GNDA 0.228531f
C3546 two_stage_opamp_dummy_magic_25_0.VD4.t26 GNDA 0.05484f
C3547 two_stage_opamp_dummy_magic_25_0.VD4.t24 GNDA 0.05484f
C3548 two_stage_opamp_dummy_magic_25_0.VD4.n20 GNDA 0.11218f
C3549 two_stage_opamp_dummy_magic_25_0.VD4.n21 GNDA 0.309358f
C3550 two_stage_opamp_dummy_magic_25_0.VD4.n22 GNDA 0.101472f
C3551 two_stage_opamp_dummy_magic_25_0.VD4.n23 GNDA 0.059483f
C3552 two_stage_opamp_dummy_magic_25_0.VD4.n24 GNDA 0.059483f
C3553 two_stage_opamp_dummy_magic_25_0.VD4.t27 GNDA 0.05484f
C3554 two_stage_opamp_dummy_magic_25_0.VD4.t19 GNDA 0.05484f
C3555 two_stage_opamp_dummy_magic_25_0.VD4.n25 GNDA 0.11218f
C3556 two_stage_opamp_dummy_magic_25_0.VD4.n26 GNDA 0.309358f
C3557 two_stage_opamp_dummy_magic_25_0.VD4.n27 GNDA 0.101472f
C3558 two_stage_opamp_dummy_magic_25_0.VD4.t25 GNDA 0.05484f
C3559 two_stage_opamp_dummy_magic_25_0.VD4.t0 GNDA 0.05484f
C3560 two_stage_opamp_dummy_magic_25_0.VD4.n28 GNDA 0.11218f
C3561 two_stage_opamp_dummy_magic_25_0.VD4.n29 GNDA 0.326446f
C3562 two_stage_opamp_dummy_magic_25_0.VD4.n30 GNDA 0.271333f
C3563 two_stage_opamp_dummy_magic_25_0.VD4.t32 GNDA 0.096159f
C3564 two_stage_opamp_dummy_magic_25_0.VD4.t34 GNDA 0.195072f
C3565 two_stage_opamp_dummy_magic_25_0.VD4.t18 GNDA 0.05484f
C3566 two_stage_opamp_dummy_magic_25_0.VD4.t10 GNDA 0.05484f
C3567 two_stage_opamp_dummy_magic_25_0.VD4.n31 GNDA 0.116347f
C3568 two_stage_opamp_dummy_magic_25_0.VD4.t29 GNDA 0.096159f
C3569 two_stage_opamp_dummy_magic_25_0.VD4.n32 GNDA 0.30186f
C3570 two_stage_opamp_dummy_magic_25_0.VD4.t31 GNDA 0.195072f
C3571 two_stage_opamp_dummy_magic_25_0.VD4.n33 GNDA 0.565887f
C3572 two_stage_opamp_dummy_magic_25_0.VD4.t30 GNDA 0.467448f
C3573 two_stage_opamp_dummy_magic_25_0.VD4.t17 GNDA 0.366642f
C3574 two_stage_opamp_dummy_magic_25_0.VD4.t9 GNDA 0.366642f
C3575 two_stage_opamp_dummy_magic_25_0.VD4.t1 GNDA 0.366642f
C3576 two_stage_opamp_dummy_magic_25_0.VD4.t11 GNDA 0.366642f
C3577 two_stage_opamp_dummy_magic_25_0.VD4.t35 GNDA 0.366642f
C3578 two_stage_opamp_dummy_magic_25_0.VD4.t15 GNDA 0.366642f
C3579 two_stage_opamp_dummy_magic_25_0.VD4.t3 GNDA 0.366642f
C3580 two_stage_opamp_dummy_magic_25_0.VD4.t5 GNDA 0.366642f
C3581 two_stage_opamp_dummy_magic_25_0.VD4.t13 GNDA 0.366642f
C3582 two_stage_opamp_dummy_magic_25_0.VD4.t7 GNDA 0.366642f
C3583 two_stage_opamp_dummy_magic_25_0.VD4.t33 GNDA 0.467448f
C3584 two_stage_opamp_dummy_magic_25_0.VD4.n34 GNDA 0.565887f
C3585 two_stage_opamp_dummy_magic_25_0.VD4.n35 GNDA 0.219169f
C3586 two_stage_opamp_dummy_magic_25_0.VD4.n36 GNDA 0.116347f
C3587 two_stage_opamp_dummy_magic_25_0.VD4.t2 GNDA 0.05484f
C3588 two_stage_opamp_dummy_magic_25_0.Vb3.t7 GNDA 0.019017f
C3589 two_stage_opamp_dummy_magic_25_0.Vb3.t4 GNDA 0.019017f
C3590 two_stage_opamp_dummy_magic_25_0.Vb3.n0 GNDA 0.061257f
C3591 two_stage_opamp_dummy_magic_25_0.Vb3.t3 GNDA 0.019017f
C3592 two_stage_opamp_dummy_magic_25_0.Vb3.t2 GNDA 0.019017f
C3593 two_stage_opamp_dummy_magic_25_0.Vb3.n1 GNDA 0.061257f
C3594 two_stage_opamp_dummy_magic_25_0.Vb3.n2 GNDA 0.337708f
C3595 two_stage_opamp_dummy_magic_25_0.Vb3.t5 GNDA 0.019017f
C3596 two_stage_opamp_dummy_magic_25_0.Vb3.t1 GNDA 0.019017f
C3597 two_stage_opamp_dummy_magic_25_0.Vb3.n3 GNDA 0.057441f
C3598 two_stage_opamp_dummy_magic_25_0.Vb3.n4 GNDA 1.05286f
C3599 two_stage_opamp_dummy_magic_25_0.Vb3.t0 GNDA 0.066561f
C3600 two_stage_opamp_dummy_magic_25_0.Vb3.t6 GNDA 0.066561f
C3601 two_stage_opamp_dummy_magic_25_0.Vb3.n5 GNDA 0.183572f
C3602 two_stage_opamp_dummy_magic_25_0.Vb3.t23 GNDA 0.094136f
C3603 two_stage_opamp_dummy_magic_25_0.Vb3.t21 GNDA 0.094136f
C3604 two_stage_opamp_dummy_magic_25_0.Vb3.t19 GNDA 0.094136f
C3605 two_stage_opamp_dummy_magic_25_0.Vb3.t13 GNDA 0.094136f
C3606 two_stage_opamp_dummy_magic_25_0.Vb3.t16 GNDA 0.108633f
C3607 two_stage_opamp_dummy_magic_25_0.Vb3.n6 GNDA 0.088198f
C3608 two_stage_opamp_dummy_magic_25_0.Vb3.n7 GNDA 0.0542f
C3609 two_stage_opamp_dummy_magic_25_0.Vb3.n8 GNDA 0.0542f
C3610 two_stage_opamp_dummy_magic_25_0.Vb3.n9 GNDA 0.047522f
C3611 two_stage_opamp_dummy_magic_25_0.Vb3.t26 GNDA 0.094136f
C3612 two_stage_opamp_dummy_magic_25_0.Vb3.t9 GNDA 0.094136f
C3613 two_stage_opamp_dummy_magic_25_0.Vb3.t15 GNDA 0.094136f
C3614 two_stage_opamp_dummy_magic_25_0.Vb3.t20 GNDA 0.094136f
C3615 two_stage_opamp_dummy_magic_25_0.Vb3.t22 GNDA 0.108633f
C3616 two_stage_opamp_dummy_magic_25_0.Vb3.n10 GNDA 0.088198f
C3617 two_stage_opamp_dummy_magic_25_0.Vb3.n11 GNDA 0.0542f
C3618 two_stage_opamp_dummy_magic_25_0.Vb3.n12 GNDA 0.0542f
C3619 two_stage_opamp_dummy_magic_25_0.Vb3.n13 GNDA 0.047522f
C3620 two_stage_opamp_dummy_magic_25_0.Vb3.n14 GNDA 0.051559f
C3621 two_stage_opamp_dummy_magic_25_0.Vb3.t25 GNDA 0.094136f
C3622 two_stage_opamp_dummy_magic_25_0.Vb3.t17 GNDA 0.094136f
C3623 two_stage_opamp_dummy_magic_25_0.Vb3.t11 GNDA 0.094136f
C3624 two_stage_opamp_dummy_magic_25_0.Vb3.t14 GNDA 0.094136f
C3625 two_stage_opamp_dummy_magic_25_0.Vb3.t8 GNDA 0.108633f
C3626 two_stage_opamp_dummy_magic_25_0.Vb3.n15 GNDA 0.088198f
C3627 two_stage_opamp_dummy_magic_25_0.Vb3.n16 GNDA 0.0542f
C3628 two_stage_opamp_dummy_magic_25_0.Vb3.n17 GNDA 0.0542f
C3629 two_stage_opamp_dummy_magic_25_0.Vb3.n18 GNDA 0.047522f
C3630 two_stage_opamp_dummy_magic_25_0.Vb3.t27 GNDA 0.094136f
C3631 two_stage_opamp_dummy_magic_25_0.Vb3.t10 GNDA 0.094136f
C3632 two_stage_opamp_dummy_magic_25_0.Vb3.t28 GNDA 0.094136f
C3633 two_stage_opamp_dummy_magic_25_0.Vb3.t12 GNDA 0.094136f
C3634 two_stage_opamp_dummy_magic_25_0.Vb3.t18 GNDA 0.108633f
C3635 two_stage_opamp_dummy_magic_25_0.Vb3.n19 GNDA 0.088198f
C3636 two_stage_opamp_dummy_magic_25_0.Vb3.n20 GNDA 0.0542f
C3637 two_stage_opamp_dummy_magic_25_0.Vb3.n21 GNDA 0.0542f
C3638 two_stage_opamp_dummy_magic_25_0.Vb3.n22 GNDA 0.047522f
C3639 two_stage_opamp_dummy_magic_25_0.Vb3.n23 GNDA 0.052638f
C3640 two_stage_opamp_dummy_magic_25_0.Vb3.n24 GNDA 1.88628f
C3641 two_stage_opamp_dummy_magic_25_0.Vb3.t24 GNDA 0.122973f
C3642 two_stage_opamp_dummy_magic_25_0.Vb3.n25 GNDA 0.467586f
C3643 two_stage_opamp_dummy_magic_25_0.Vb3.n26 GNDA 1.88739f
C3644 bgr_11_0.VB3_CUR_BIAS GNDA 2.91306f
C3645 two_stage_opamp_dummy_magic_25_0.cap_res_X.t56 GNDA 0.412258f
C3646 two_stage_opamp_dummy_magic_25_0.cap_res_X.t92 GNDA 0.413752f
C3647 two_stage_opamp_dummy_magic_25_0.cap_res_X.t24 GNDA 0.412258f
C3648 two_stage_opamp_dummy_magic_25_0.cap_res_X.t61 GNDA 0.413752f
C3649 two_stage_opamp_dummy_magic_25_0.cap_res_X.t114 GNDA 0.412258f
C3650 two_stage_opamp_dummy_magic_25_0.cap_res_X.t78 GNDA 0.413752f
C3651 two_stage_opamp_dummy_magic_25_0.cap_res_X.t53 GNDA 0.412258f
C3652 two_stage_opamp_dummy_magic_25_0.cap_res_X.t87 GNDA 0.413752f
C3653 two_stage_opamp_dummy_magic_25_0.cap_res_X.t70 GNDA 0.412258f
C3654 two_stage_opamp_dummy_magic_25_0.cap_res_X.t36 GNDA 0.413752f
C3655 two_stage_opamp_dummy_magic_25_0.cap_res_X.t89 GNDA 0.412258f
C3656 two_stage_opamp_dummy_magic_25_0.cap_res_X.t129 GNDA 0.413752f
C3657 two_stage_opamp_dummy_magic_25_0.cap_res_X.t108 GNDA 0.412258f
C3658 two_stage_opamp_dummy_magic_25_0.cap_res_X.t74 GNDA 0.413752f
C3659 two_stage_opamp_dummy_magic_25_0.cap_res_X.t58 GNDA 0.412258f
C3660 two_stage_opamp_dummy_magic_25_0.cap_res_X.t91 GNDA 0.413752f
C3661 two_stage_opamp_dummy_magic_25_0.cap_res_X.t76 GNDA 0.412258f
C3662 two_stage_opamp_dummy_magic_25_0.cap_res_X.t43 GNDA 0.413752f
C3663 two_stage_opamp_dummy_magic_25_0.cap_res_X.t95 GNDA 0.412258f
C3664 two_stage_opamp_dummy_magic_25_0.cap_res_X.t132 GNDA 0.413752f
C3665 two_stage_opamp_dummy_magic_25_0.cap_res_X.t113 GNDA 0.412258f
C3666 two_stage_opamp_dummy_magic_25_0.cap_res_X.t80 GNDA 0.413752f
C3667 two_stage_opamp_dummy_magic_25_0.cap_res_X.t137 GNDA 0.412258f
C3668 two_stage_opamp_dummy_magic_25_0.cap_res_X.t33 GNDA 0.413752f
C3669 two_stage_opamp_dummy_magic_25_0.cap_res_X.t14 GNDA 0.412258f
C3670 two_stage_opamp_dummy_magic_25_0.cap_res_X.t119 GNDA 0.413752f
C3671 two_stage_opamp_dummy_magic_25_0.cap_res_X.t101 GNDA 0.412258f
C3672 two_stage_opamp_dummy_magic_25_0.cap_res_X.t0 GNDA 0.413752f
C3673 two_stage_opamp_dummy_magic_25_0.cap_res_X.t120 GNDA 0.412258f
C3674 two_stage_opamp_dummy_magic_25_0.cap_res_X.t84 GNDA 0.413752f
C3675 two_stage_opamp_dummy_magic_25_0.cap_res_X.t5 GNDA 0.412258f
C3676 two_stage_opamp_dummy_magic_25_0.cap_res_X.t41 GNDA 0.413752f
C3677 two_stage_opamp_dummy_magic_25_0.cap_res_X.t22 GNDA 0.412258f
C3678 two_stage_opamp_dummy_magic_25_0.cap_res_X.t125 GNDA 0.413752f
C3679 two_stage_opamp_dummy_magic_25_0.cap_res_X.t45 GNDA 0.412258f
C3680 two_stage_opamp_dummy_magic_25_0.cap_res_X.t79 GNDA 0.413752f
C3681 two_stage_opamp_dummy_magic_25_0.cap_res_X.t59 GNDA 0.412258f
C3682 two_stage_opamp_dummy_magic_25_0.cap_res_X.t27 GNDA 0.413752f
C3683 two_stage_opamp_dummy_magic_25_0.cap_res_X.t82 GNDA 0.412258f
C3684 two_stage_opamp_dummy_magic_25_0.cap_res_X.t116 GNDA 0.413752f
C3685 two_stage_opamp_dummy_magic_25_0.cap_res_X.t97 GNDA 0.412258f
C3686 two_stage_opamp_dummy_magic_25_0.cap_res_X.t63 GNDA 0.413752f
C3687 two_stage_opamp_dummy_magic_25_0.cap_res_X.t48 GNDA 0.412258f
C3688 two_stage_opamp_dummy_magic_25_0.cap_res_X.t83 GNDA 0.413752f
C3689 two_stage_opamp_dummy_magic_25_0.cap_res_X.t64 GNDA 0.412258f
C3690 two_stage_opamp_dummy_magic_25_0.cap_res_X.t32 GNDA 0.413752f
C3691 two_stage_opamp_dummy_magic_25_0.cap_res_X.t86 GNDA 0.412258f
C3692 two_stage_opamp_dummy_magic_25_0.cap_res_X.t122 GNDA 0.413752f
C3693 two_stage_opamp_dummy_magic_25_0.cap_res_X.t103 GNDA 0.412258f
C3694 two_stage_opamp_dummy_magic_25_0.cap_res_X.t69 GNDA 0.413752f
C3695 two_stage_opamp_dummy_magic_25_0.cap_res_X.t127 GNDA 0.412258f
C3696 two_stage_opamp_dummy_magic_25_0.cap_res_X.t23 GNDA 0.413752f
C3697 two_stage_opamp_dummy_magic_25_0.cap_res_X.t6 GNDA 0.412258f
C3698 two_stage_opamp_dummy_magic_25_0.cap_res_X.t107 GNDA 0.413752f
C3699 two_stage_opamp_dummy_magic_25_0.cap_res_X.t90 GNDA 0.412258f
C3700 two_stage_opamp_dummy_magic_25_0.cap_res_X.t128 GNDA 0.413752f
C3701 two_stage_opamp_dummy_magic_25_0.cap_res_X.t109 GNDA 0.412258f
C3702 two_stage_opamp_dummy_magic_25_0.cap_res_X.t75 GNDA 0.413752f
C3703 two_stage_opamp_dummy_magic_25_0.cap_res_X.t94 GNDA 0.412258f
C3704 two_stage_opamp_dummy_magic_25_0.cap_res_X.t46 GNDA 0.413752f
C3705 two_stage_opamp_dummy_magic_25_0.cap_res_X.t126 GNDA 0.412258f
C3706 two_stage_opamp_dummy_magic_25_0.cap_res_X.t42 GNDA 0.413752f
C3707 two_stage_opamp_dummy_magic_25_0.cap_res_X.t3 GNDA 0.412258f
C3708 two_stage_opamp_dummy_magic_25_0.cap_res_X.t40 GNDA 0.413752f
C3709 two_stage_opamp_dummy_magic_25_0.cap_res_X.t20 GNDA 0.412258f
C3710 two_stage_opamp_dummy_magic_25_0.cap_res_X.t123 GNDA 0.413752f
C3711 two_stage_opamp_dummy_magic_25_0.cap_res_X.t39 GNDA 0.412258f
C3712 two_stage_opamp_dummy_magic_25_0.cap_res_X.t71 GNDA 0.413752f
C3713 two_stage_opamp_dummy_magic_25_0.cap_res_X.t54 GNDA 0.412258f
C3714 two_stage_opamp_dummy_magic_25_0.cap_res_X.t19 GNDA 0.413752f
C3715 two_stage_opamp_dummy_magic_25_0.cap_res_X.t98 GNDA 0.412258f
C3716 two_stage_opamp_dummy_magic_25_0.cap_res_X.t136 GNDA 0.413752f
C3717 two_stage_opamp_dummy_magic_25_0.cap_res_X.t10 GNDA 0.412258f
C3718 two_stage_opamp_dummy_magic_25_0.cap_res_X.t52 GNDA 0.432471f
C3719 two_stage_opamp_dummy_magic_25_0.cap_res_X.t37 GNDA 0.412258f
C3720 two_stage_opamp_dummy_magic_25_0.cap_res_X.t77 GNDA 0.221432f
C3721 two_stage_opamp_dummy_magic_25_0.cap_res_X.n0 GNDA 0.236987f
C3722 two_stage_opamp_dummy_magic_25_0.cap_res_X.t17 GNDA 0.412258f
C3723 two_stage_opamp_dummy_magic_25_0.cap_res_X.t55 GNDA 0.221432f
C3724 two_stage_opamp_dummy_magic_25_0.cap_res_X.n1 GNDA 0.235076f
C3725 two_stage_opamp_dummy_magic_25_0.cap_res_X.t118 GNDA 0.412258f
C3726 two_stage_opamp_dummy_magic_25_0.cap_res_X.t21 GNDA 0.221432f
C3727 two_stage_opamp_dummy_magic_25_0.cap_res_X.n2 GNDA 0.235076f
C3728 two_stage_opamp_dummy_magic_25_0.cap_res_X.t2 GNDA 0.412258f
C3729 two_stage_opamp_dummy_magic_25_0.cap_res_X.t44 GNDA 0.221432f
C3730 two_stage_opamp_dummy_magic_25_0.cap_res_X.n3 GNDA 0.235076f
C3731 two_stage_opamp_dummy_magic_25_0.cap_res_X.t100 GNDA 0.412258f
C3732 two_stage_opamp_dummy_magic_25_0.cap_res_X.t4 GNDA 0.221432f
C3733 two_stage_opamp_dummy_magic_25_0.cap_res_X.n4 GNDA 0.235076f
C3734 two_stage_opamp_dummy_magic_25_0.cap_res_X.t65 GNDA 0.412258f
C3735 two_stage_opamp_dummy_magic_25_0.cap_res_X.t105 GNDA 0.221432f
C3736 two_stage_opamp_dummy_magic_25_0.cap_res_X.n5 GNDA 0.235076f
C3737 two_stage_opamp_dummy_magic_25_0.cap_res_X.t29 GNDA 0.412258f
C3738 two_stage_opamp_dummy_magic_25_0.cap_res_X.t67 GNDA 0.221432f
C3739 two_stage_opamp_dummy_magic_25_0.cap_res_X.n6 GNDA 0.235076f
C3740 two_stage_opamp_dummy_magic_25_0.cap_res_X.t49 GNDA 0.412258f
C3741 two_stage_opamp_dummy_magic_25_0.cap_res_X.t88 GNDA 0.221432f
C3742 two_stage_opamp_dummy_magic_25_0.cap_res_X.n7 GNDA 0.235076f
C3743 two_stage_opamp_dummy_magic_25_0.cap_res_X.t8 GNDA 0.412258f
C3744 two_stage_opamp_dummy_magic_25_0.cap_res_X.t51 GNDA 0.221432f
C3745 two_stage_opamp_dummy_magic_25_0.cap_res_X.n8 GNDA 0.235076f
C3746 two_stage_opamp_dummy_magic_25_0.cap_res_X.t111 GNDA 0.412258f
C3747 two_stage_opamp_dummy_magic_25_0.cap_res_X.t12 GNDA 0.221432f
C3748 two_stage_opamp_dummy_magic_25_0.cap_res_X.n9 GNDA 0.235076f
C3749 two_stage_opamp_dummy_magic_25_0.cap_res_X.t60 GNDA 0.412258f
C3750 two_stage_opamp_dummy_magic_25_0.cap_res_X.t93 GNDA 0.413752f
C3751 two_stage_opamp_dummy_magic_25_0.cap_res_X.t134 GNDA 0.199307f
C3752 two_stage_opamp_dummy_magic_25_0.cap_res_X.n10 GNDA 0.257077f
C3753 two_stage_opamp_dummy_magic_25_0.cap_res_X.t38 GNDA 0.220062f
C3754 two_stage_opamp_dummy_magic_25_0.cap_res_X.n11 GNDA 0.279201f
C3755 two_stage_opamp_dummy_magic_25_0.cap_res_X.t106 GNDA 0.220062f
C3756 two_stage_opamp_dummy_magic_25_0.cap_res_X.n12 GNDA 0.299832f
C3757 two_stage_opamp_dummy_magic_25_0.cap_res_X.t72 GNDA 0.220062f
C3758 two_stage_opamp_dummy_magic_25_0.cap_res_X.n13 GNDA 0.299832f
C3759 two_stage_opamp_dummy_magic_25_0.cap_res_X.t135 GNDA 0.220062f
C3760 two_stage_opamp_dummy_magic_25_0.cap_res_X.n14 GNDA 0.299832f
C3761 two_stage_opamp_dummy_magic_25_0.cap_res_X.t26 GNDA 0.220062f
C3762 two_stage_opamp_dummy_magic_25_0.cap_res_X.n15 GNDA 0.299832f
C3763 two_stage_opamp_dummy_magic_25_0.cap_res_X.t57 GNDA 0.220062f
C3764 two_stage_opamp_dummy_magic_25_0.cap_res_X.n16 GNDA 0.299832f
C3765 two_stage_opamp_dummy_magic_25_0.cap_res_X.t18 GNDA 0.220062f
C3766 two_stage_opamp_dummy_magic_25_0.cap_res_X.n17 GNDA 0.299832f
C3767 two_stage_opamp_dummy_magic_25_0.cap_res_X.t117 GNDA 0.220062f
C3768 two_stage_opamp_dummy_magic_25_0.cap_res_X.n18 GNDA 0.299832f
C3769 two_stage_opamp_dummy_magic_25_0.cap_res_X.t13 GNDA 0.220062f
C3770 two_stage_opamp_dummy_magic_25_0.cap_res_X.n19 GNDA 0.299832f
C3771 two_stage_opamp_dummy_magic_25_0.cap_res_X.t112 GNDA 0.220062f
C3772 two_stage_opamp_dummy_magic_25_0.cap_res_X.n20 GNDA 0.299832f
C3773 two_stage_opamp_dummy_magic_25_0.cap_res_X.t73 GNDA 0.220062f
C3774 two_stage_opamp_dummy_magic_25_0.cap_res_X.n21 GNDA 0.299832f
C3775 two_stage_opamp_dummy_magic_25_0.cap_res_X.t35 GNDA 0.220062f
C3776 two_stage_opamp_dummy_magic_25_0.cap_res_X.n22 GNDA 0.299832f
C3777 two_stage_opamp_dummy_magic_25_0.cap_res_X.t68 GNDA 0.220062f
C3778 two_stage_opamp_dummy_magic_25_0.cap_res_X.n23 GNDA 0.299832f
C3779 two_stage_opamp_dummy_magic_25_0.cap_res_X.t30 GNDA 0.220062f
C3780 two_stage_opamp_dummy_magic_25_0.cap_res_X.n24 GNDA 0.299832f
C3781 two_stage_opamp_dummy_magic_25_0.cap_res_X.t130 GNDA 0.220062f
C3782 two_stage_opamp_dummy_magic_25_0.cap_res_X.n25 GNDA 0.299832f
C3783 two_stage_opamp_dummy_magic_25_0.cap_res_X.t25 GNDA 0.220062f
C3784 two_stage_opamp_dummy_magic_25_0.cap_res_X.n26 GNDA 0.299832f
C3785 two_stage_opamp_dummy_magic_25_0.cap_res_X.t124 GNDA 0.220062f
C3786 two_stage_opamp_dummy_magic_25_0.cap_res_X.n27 GNDA 0.299832f
C3787 two_stage_opamp_dummy_magic_25_0.cap_res_X.t96 GNDA 0.220062f
C3788 two_stage_opamp_dummy_magic_25_0.cap_res_X.n28 GNDA 0.299832f
C3789 two_stage_opamp_dummy_magic_25_0.cap_res_X.t133 GNDA 0.220062f
C3790 two_stage_opamp_dummy_magic_25_0.cap_res_X.n29 GNDA 0.276337f
C3791 two_stage_opamp_dummy_magic_25_0.cap_res_X.t110 GNDA 0.413752f
C3792 two_stage_opamp_dummy_magic_25_0.cap_res_X.t7 GNDA 0.413752f
C3793 two_stage_opamp_dummy_magic_25_0.cap_res_X.t102 GNDA 0.412258f
C3794 two_stage_opamp_dummy_magic_25_0.cap_res_X.t11 GNDA 0.434383f
C3795 two_stage_opamp_dummy_magic_25_0.cap_res_X.t47 GNDA 0.221432f
C3796 two_stage_opamp_dummy_magic_25_0.cap_res_X.n30 GNDA 0.255706f
C3797 two_stage_opamp_dummy_magic_25_0.cap_res_X.t9 GNDA 0.412258f
C3798 two_stage_opamp_dummy_magic_25_0.cap_res_X.t34 GNDA 0.434383f
C3799 two_stage_opamp_dummy_magic_25_0.cap_res_X.t16 GNDA 0.413752f
C3800 two_stage_opamp_dummy_magic_25_0.cap_res_X.t81 GNDA 0.412258f
C3801 two_stage_opamp_dummy_magic_25_0.cap_res_X.t115 GNDA 0.221432f
C3802 two_stage_opamp_dummy_magic_25_0.cap_res_X.n31 GNDA 0.255706f
C3803 two_stage_opamp_dummy_magic_25_0.cap_res_X.t121 GNDA 0.412258f
C3804 two_stage_opamp_dummy_magic_25_0.cap_res_X.t104 GNDA 0.434383f
C3805 two_stage_opamp_dummy_magic_25_0.cap_res_X.t1 GNDA 0.221432f
C3806 two_stage_opamp_dummy_magic_25_0.cap_res_X.n32 GNDA 0.235076f
C3807 two_stage_opamp_dummy_magic_25_0.cap_res_X.t85 GNDA 0.412258f
C3808 two_stage_opamp_dummy_magic_25_0.cap_res_X.t66 GNDA 0.434383f
C3809 two_stage_opamp_dummy_magic_25_0.cap_res_X.t99 GNDA 0.221432f
C3810 two_stage_opamp_dummy_magic_25_0.cap_res_X.n33 GNDA 0.235076f
C3811 two_stage_opamp_dummy_magic_25_0.cap_res_X.t50 GNDA 0.412258f
C3812 two_stage_opamp_dummy_magic_25_0.cap_res_X.t31 GNDA 0.434383f
C3813 two_stage_opamp_dummy_magic_25_0.cap_res_X.t62 GNDA 0.221432f
C3814 two_stage_opamp_dummy_magic_25_0.cap_res_X.n34 GNDA 0.235076f
C3815 two_stage_opamp_dummy_magic_25_0.cap_res_X.n35 GNDA 0.235076f
C3816 two_stage_opamp_dummy_magic_25_0.cap_res_X.t28 GNDA 0.221432f
C3817 two_stage_opamp_dummy_magic_25_0.cap_res_X.t131 GNDA 0.434383f
C3818 two_stage_opamp_dummy_magic_25_0.cap_res_X.t15 GNDA 0.590705f
C3819 two_stage_opamp_dummy_magic_25_0.cap_res_X.t138 GNDA 0.355569f
C3820 VOUT-.n1 GNDA 0.075396f
C3821 VOUT-.n4 GNDA 0.056547f
C3822 VOUT-.n5 GNDA 0.094246f
C3823 VOUT-.n6 GNDA 0.056547f
C3824 VOUT-.n7 GNDA 0.056547f
C3825 VOUT-.n9 GNDA 0.038452f
C3826 VOUT-.n11 GNDA 0.038452f
C3827 VOUT-.n13 GNDA 0.075396f
C3828 VOUT-.n14 GNDA 0.038452f
C3829 VOUT-.n16 GNDA 0.038452f
C3830 VOUT-.n18 GNDA 0.049762f
C3831 VOUT-.n19 GNDA 0.071794f
C3832 VOUT-.n20 GNDA 0.069867f
C3833 VOUT-.n21 GNDA 0.049762f
C3834 VOUT-.n22 GNDA 0.049762f
C3835 VOUT-.n23 GNDA 0.069867f
C3836 VOUT-.n24 GNDA 0.069867f
C3837 VOUT-.n25 GNDA 0.049762f
C3838 VOUT-.n26 GNDA 0.079664f
C3839 VOUT-.t0 GNDA 0.045238f
C3840 VOUT-.t11 GNDA 0.045238f
C3841 VOUT-.n27 GNDA 0.092692f
C3842 VOUT-.n28 GNDA 0.239266f
C3843 VOUT-.t10 GNDA 0.045238f
C3844 VOUT-.t2 GNDA 0.045238f
C3845 VOUT-.n29 GNDA 0.092692f
C3846 VOUT-.n30 GNDA 0.236855f
C3847 VOUT-.n31 GNDA 0.057525f
C3848 VOUT-.t6 GNDA 0.045238f
C3849 VOUT-.t1 GNDA 0.045238f
C3850 VOUT-.n32 GNDA 0.092692f
C3851 VOUT-.n33 GNDA 0.236855f
C3852 VOUT-.n34 GNDA 0.032607f
C3853 VOUT-.t4 GNDA 0.045238f
C3854 VOUT-.t7 GNDA 0.045238f
C3855 VOUT-.n35 GNDA 0.092692f
C3856 VOUT-.n36 GNDA 0.236855f
C3857 VOUT-.n37 GNDA 0.032607f
C3858 VOUT-.t17 GNDA 0.045238f
C3859 VOUT-.t12 GNDA 0.045238f
C3860 VOUT-.n38 GNDA 0.092692f
C3861 VOUT-.n39 GNDA 0.239266f
C3862 VOUT-.n40 GNDA 0.057525f
C3863 VOUT-.t16 GNDA 0.045238f
C3864 VOUT-.t5 GNDA 0.045238f
C3865 VOUT-.n41 GNDA 0.092692f
C3866 VOUT-.n42 GNDA 0.236855f
C3867 VOUT-.n43 GNDA 0.038033f
C3868 VOUT-.n44 GNDA 0.022619f
C3869 VOUT-.n45 GNDA 0.022619f
C3870 VOUT-.n46 GNDA 0.038033f
C3871 VOUT-.n47 GNDA 0.069867f
C3872 VOUT-.n48 GNDA 0.0978f
C3873 VOUT-.n49 GNDA 0.121863f
C3874 VOUT-.n50 GNDA 0.170559f
C3875 VOUT-.n51 GNDA 0.049762f
C3876 VOUT-.n52 GNDA 0.081428f
C3877 VOUT-.n53 GNDA 0.049762f
C3878 VOUT-.n54 GNDA 0.081428f
C3879 VOUT-.n55 GNDA 0.049762f
C3880 VOUT-.n56 GNDA 0.049762f
C3881 VOUT-.n57 GNDA 0.049762f
C3882 VOUT-.n58 GNDA 0.081428f
C3883 VOUT-.n59 GNDA 0.049762f
C3884 VOUT-.n60 GNDA 0.074642f
C3885 VOUT-.n61 GNDA 0.239761f
C3886 VOUT-.n62 GNDA 0.232975f
C3887 VOUT-.n64 GNDA 0.075396f
C3888 VOUT-.n65 GNDA 0.03619f
C3889 VOUT-.n66 GNDA 0.537199f
C3890 VOUT-.n69 GNDA 0.056547f
C3891 VOUT-.n70 GNDA 0.056547f
C3892 VOUT-.t96 GNDA 0.306722f
C3893 VOUT-.t63 GNDA 0.301586f
C3894 VOUT-.n71 GNDA 0.202203f
C3895 VOUT-.t22 GNDA 0.301586f
C3896 VOUT-.n72 GNDA 0.131944f
C3897 VOUT-.t58 GNDA 0.306722f
C3898 VOUT-.t20 GNDA 0.301586f
C3899 VOUT-.n73 GNDA 0.202203f
C3900 VOUT-.t118 GNDA 0.301586f
C3901 VOUT-.t45 GNDA 0.306079f
C3902 VOUT-.t148 GNDA 0.306079f
C3903 VOUT-.t107 GNDA 0.306079f
C3904 VOUT-.t127 GNDA 0.306079f
C3905 VOUT-.t91 GNDA 0.306079f
C3906 VOUT-.t56 GNDA 0.306079f
C3907 VOUT-.t154 GNDA 0.306079f
C3908 VOUT-.t38 GNDA 0.306079f
C3909 VOUT-.t139 GNDA 0.306079f
C3910 VOUT-.t119 GNDA 0.306079f
C3911 VOUT-.t146 GNDA 0.306079f
C3912 VOUT-.t104 GNDA 0.301586f
C3913 VOUT-.n74 GNDA 0.202846f
C3914 VOUT-.t79 GNDA 0.301586f
C3915 VOUT-.n75 GNDA 0.259394f
C3916 VOUT-.t101 GNDA 0.301586f
C3917 VOUT-.n76 GNDA 0.259394f
C3918 VOUT-.t135 GNDA 0.301586f
C3919 VOUT-.n77 GNDA 0.259394f
C3920 VOUT-.t112 GNDA 0.301586f
C3921 VOUT-.n78 GNDA 0.259394f
C3922 VOUT-.t152 GNDA 0.301586f
C3923 VOUT-.n79 GNDA 0.259394f
C3924 VOUT-.t51 GNDA 0.301586f
C3925 VOUT-.n80 GNDA 0.259394f
C3926 VOUT-.t89 GNDA 0.301586f
C3927 VOUT-.n81 GNDA 0.259394f
C3928 VOUT-.t68 GNDA 0.301586f
C3929 VOUT-.n82 GNDA 0.259394f
C3930 VOUT-.t105 GNDA 0.301586f
C3931 VOUT-.n83 GNDA 0.259394f
C3932 VOUT-.t144 GNDA 0.301586f
C3933 VOUT-.n84 GNDA 0.259394f
C3934 VOUT-.n85 GNDA 0.245038f
C3935 VOUT-.t117 GNDA 0.306722f
C3936 VOUT-.t85 GNDA 0.301586f
C3937 VOUT-.n86 GNDA 0.202203f
C3938 VOUT-.t50 GNDA 0.301586f
C3939 VOUT-.t102 GNDA 0.306722f
C3940 VOUT-.t137 GNDA 0.301586f
C3941 VOUT-.n87 GNDA 0.202203f
C3942 VOUT-.n88 GNDA 0.245038f
C3943 VOUT-.t153 GNDA 0.306722f
C3944 VOUT-.t116 GNDA 0.301586f
C3945 VOUT-.n89 GNDA 0.202203f
C3946 VOUT-.t84 GNDA 0.301586f
C3947 VOUT-.t136 GNDA 0.306722f
C3948 VOUT-.t33 GNDA 0.301586f
C3949 VOUT-.n90 GNDA 0.202203f
C3950 VOUT-.n91 GNDA 0.245038f
C3951 VOUT-.t62 GNDA 0.306722f
C3952 VOUT-.t110 GNDA 0.301586f
C3953 VOUT-.n92 GNDA 0.202203f
C3954 VOUT-.t21 GNDA 0.301586f
C3955 VOUT-.t30 GNDA 0.306722f
C3956 VOUT-.t114 GNDA 0.301586f
C3957 VOUT-.n93 GNDA 0.202203f
C3958 VOUT-.n94 GNDA 0.245038f
C3959 VOUT-.t66 GNDA 0.306722f
C3960 VOUT-.t28 GNDA 0.301586f
C3961 VOUT-.n95 GNDA 0.202203f
C3962 VOUT-.t130 GNDA 0.301586f
C3963 VOUT-.t47 GNDA 0.306722f
C3964 VOUT-.t81 GNDA 0.301586f
C3965 VOUT-.n96 GNDA 0.202203f
C3966 VOUT-.n97 GNDA 0.245038f
C3967 VOUT-.t29 GNDA 0.306722f
C3968 VOUT-.t133 GNDA 0.301586f
C3969 VOUT-.n98 GNDA 0.202203f
C3970 VOUT-.t99 GNDA 0.301586f
C3971 VOUT-.t150 GNDA 0.306722f
C3972 VOUT-.t49 GNDA 0.301586f
C3973 VOUT-.n99 GNDA 0.202203f
C3974 VOUT-.n100 GNDA 0.245038f
C3975 VOUT-.t70 GNDA 0.306722f
C3976 VOUT-.t34 GNDA 0.301586f
C3977 VOUT-.n101 GNDA 0.202203f
C3978 VOUT-.t138 GNDA 0.301586f
C3979 VOUT-.t53 GNDA 0.306722f
C3980 VOUT-.t87 GNDA 0.301586f
C3981 VOUT-.n102 GNDA 0.202203f
C3982 VOUT-.n103 GNDA 0.245038f
C3983 VOUT-.t100 GNDA 0.306722f
C3984 VOUT-.t64 GNDA 0.301586f
C3985 VOUT-.n104 GNDA 0.202203f
C3986 VOUT-.t23 GNDA 0.301586f
C3987 VOUT-.t54 GNDA 0.306722f
C3988 VOUT-.t145 GNDA 0.301586f
C3989 VOUT-.n105 GNDA 0.197491f
C3990 VOUT-.t141 GNDA 0.306722f
C3991 VOUT-.t25 GNDA 0.301586f
C3992 VOUT-.n106 GNDA 0.197491f
C3993 VOUT-.t106 GNDA 0.306722f
C3994 VOUT-.t125 GNDA 0.301586f
C3995 VOUT-.n107 GNDA 0.197491f
C3996 VOUT-.t71 GNDA 0.306722f
C3997 VOUT-.t90 GNDA 0.301586f
C3998 VOUT-.n108 GNDA 0.197491f
C3999 VOUT-.t35 GNDA 0.306722f
C4000 VOUT-.t52 GNDA 0.301586f
C4001 VOUT-.n109 GNDA 0.199376f
C4002 VOUT-.t75 GNDA 0.306332f
C4003 VOUT-.t147 GNDA 0.306722f
C4004 VOUT-.t122 GNDA 0.301586f
C4005 VOUT-.n110 GNDA 0.202203f
C4006 VOUT-.t140 GNDA 0.301586f
C4007 VOUT-.n111 GNDA 0.131944f
C4008 VOUT-.t41 GNDA 0.301586f
C4009 VOUT-.n112 GNDA 0.262911f
C4010 VOUT-.t155 GNDA 0.301586f
C4011 VOUT-.n113 GNDA 0.195088f
C4012 VOUT-.t57 GNDA 0.301586f
C4013 VOUT-.n114 GNDA 0.193203f
C4014 VOUT-.t94 GNDA 0.301586f
C4015 VOUT-.n115 GNDA 0.193203f
C4016 VOUT-.t128 GNDA 0.301586f
C4017 VOUT-.n116 GNDA 0.193203f
C4018 VOUT-.t109 GNDA 0.301586f
C4019 VOUT-.n117 GNDA 0.193203f
C4020 VOUT-.t149 GNDA 0.301586f
C4021 VOUT-.n118 GNDA 0.131944f
C4022 VOUT-.t46 GNDA 0.301586f
C4023 VOUT-.n119 GNDA 0.131944f
C4024 VOUT-.n120 GNDA 0.188491f
C4025 VOUT-.t132 GNDA 0.306722f
C4026 VOUT-.t95 GNDA 0.301586f
C4027 VOUT-.n121 GNDA 0.202203f
C4028 VOUT-.t60 GNDA 0.301586f
C4029 VOUT-.t42 GNDA 0.306722f
C4030 VOUT-.t78 GNDA 0.301586f
C4031 VOUT-.n122 GNDA 0.202203f
C4032 VOUT-.n123 GNDA 0.245038f
C4033 VOUT-.t103 GNDA 0.306722f
C4034 VOUT-.t69 GNDA 0.301586f
C4035 VOUT-.n124 GNDA 0.202203f
C4036 VOUT-.t32 GNDA 0.301586f
C4037 VOUT-.t86 GNDA 0.306722f
C4038 VOUT-.t120 GNDA 0.301586f
C4039 VOUT-.n125 GNDA 0.202203f
C4040 VOUT-.n126 GNDA 0.245038f
C4041 VOUT-.t67 GNDA 0.306722f
C4042 VOUT-.t27 GNDA 0.301586f
C4043 VOUT-.n127 GNDA 0.202203f
C4044 VOUT-.t131 GNDA 0.301586f
C4045 VOUT-.t48 GNDA 0.306722f
C4046 VOUT-.t82 GNDA 0.301586f
C4047 VOUT-.n128 GNDA 0.202203f
C4048 VOUT-.n129 GNDA 0.245038f
C4049 VOUT-.t98 GNDA 0.306722f
C4050 VOUT-.t65 GNDA 0.301586f
C4051 VOUT-.n130 GNDA 0.202203f
C4052 VOUT-.t26 GNDA 0.301586f
C4053 VOUT-.t80 GNDA 0.306722f
C4054 VOUT-.t113 GNDA 0.301586f
C4055 VOUT-.n131 GNDA 0.202203f
C4056 VOUT-.n132 GNDA 0.245038f
C4057 VOUT-.t61 GNDA 0.306722f
C4058 VOUT-.t24 GNDA 0.301586f
C4059 VOUT-.n133 GNDA 0.202203f
C4060 VOUT-.t126 GNDA 0.301586f
C4061 VOUT-.t43 GNDA 0.306722f
C4062 VOUT-.t76 GNDA 0.301586f
C4063 VOUT-.n134 GNDA 0.202203f
C4064 VOUT-.n135 GNDA 0.245038f
C4065 VOUT-.t19 GNDA 0.306722f
C4066 VOUT-.t123 GNDA 0.301586f
C4067 VOUT-.n136 GNDA 0.202203f
C4068 VOUT-.t88 GNDA 0.301586f
C4069 VOUT-.t142 GNDA 0.306722f
C4070 VOUT-.t37 GNDA 0.301586f
C4071 VOUT-.n137 GNDA 0.202203f
C4072 VOUT-.n138 GNDA 0.245038f
C4073 VOUT-.t55 GNDA 0.306722f
C4074 VOUT-.t156 GNDA 0.301586f
C4075 VOUT-.n139 GNDA 0.202203f
C4076 VOUT-.t121 GNDA 0.301586f
C4077 VOUT-.t36 GNDA 0.306722f
C4078 VOUT-.t72 GNDA 0.301586f
C4079 VOUT-.n140 GNDA 0.202203f
C4080 VOUT-.n141 GNDA 0.245038f
C4081 VOUT-.t151 GNDA 0.306722f
C4082 VOUT-.t115 GNDA 0.301586f
C4083 VOUT-.n142 GNDA 0.202203f
C4084 VOUT-.t83 GNDA 0.301586f
C4085 VOUT-.t134 GNDA 0.306722f
C4086 VOUT-.t31 GNDA 0.301586f
C4087 VOUT-.n143 GNDA 0.202203f
C4088 VOUT-.n144 GNDA 0.245038f
C4089 VOUT-.t111 GNDA 0.306722f
C4090 VOUT-.t77 GNDA 0.301586f
C4091 VOUT-.n145 GNDA 0.202203f
C4092 VOUT-.t44 GNDA 0.301586f
C4093 VOUT-.t97 GNDA 0.306722f
C4094 VOUT-.t129 GNDA 0.301586f
C4095 VOUT-.n146 GNDA 0.202203f
C4096 VOUT-.n147 GNDA 0.245038f
C4097 VOUT-.t74 GNDA 0.306722f
C4098 VOUT-.t40 GNDA 0.301586f
C4099 VOUT-.n148 GNDA 0.202203f
C4100 VOUT-.t143 GNDA 0.301586f
C4101 VOUT-.t59 GNDA 0.306722f
C4102 VOUT-.t93 GNDA 0.301586f
C4103 VOUT-.n149 GNDA 0.202203f
C4104 VOUT-.n150 GNDA 0.245038f
C4105 VOUT-.t108 GNDA 0.306722f
C4106 VOUT-.t73 GNDA 0.301586f
C4107 VOUT-.n151 GNDA 0.202203f
C4108 VOUT-.t39 GNDA 0.301586f
C4109 VOUT-.n152 GNDA 0.245038f
C4110 VOUT-.t124 GNDA 0.301586f
C4111 VOUT-.n153 GNDA 0.128631f
C4112 VOUT-.t92 GNDA 0.301586f
C4113 VOUT-.n154 GNDA 0.340712f
C4114 VOUT-.n155 GNDA 0.277082f
C4115 VOUT-.n156 GNDA 0.056547f
C4116 VOUT-.n157 GNDA 0.056547f
C4117 VOUT-.n158 GNDA 0.056547f
C4118 VOUT-.n159 GNDA 0.165862f
C4119 VOUT-.n160 GNDA 0.05991f
C4120 VOUT-.n161 GNDA 0.056964f
C4121 VOUT-.n163 GNDA 0.546624f
C4122 VOUT-.n164 GNDA 0.056547f
C4123 VOUT-.n165 GNDA 1.12152f
C4124 VOUT-.n169 GNDA 0.038452f
C4125 VOUT-.n170 GNDA 0.038452f
C4126 VOUT-.n171 GNDA 0.03619f
C4127 VOUT-.n172 GNDA 0.075396f
C4128 VOUT-.n173 GNDA 0.038452f
C4129 VOUT-.n174 GNDA 0.038452f
C4130 VOUT-.n176 GNDA 1.1121f
C4131 VOUT-.n177 GNDA 0.101785f
C4132 VOUT-.t9 GNDA 0.086084f
C4133 VOUT-.n178 GNDA 0.251692f
C4134 VOUT-.n179 GNDA 0.03619f
C4135 VOUT-.t8 GNDA 0.052778f
C4136 VOUT-.t15 GNDA 0.052778f
C4137 VOUT-.n180 GNDA 0.113399f
C4138 VOUT-.n181 GNDA 0.272721f
C4139 VOUT-.n182 GNDA 0.03619f
C4140 VOUT-.n183 GNDA 0.233708f
C4141 VOUT-.t3 GNDA 0.052778f
C4142 VOUT-.t18 GNDA 0.052778f
C4143 VOUT-.n184 GNDA 0.113399f
C4144 VOUT-.n185 GNDA 0.282248f
C4145 VOUT-.n186 GNDA 0.161331f
C4146 VOUT-.t13 GNDA 0.052778f
C4147 VOUT-.t14 GNDA 0.052778f
C4148 VOUT-.n187 GNDA 0.113399f
C4149 VOUT-.n188 GNDA 0.268133f
C4150 VOUT-.n189 GNDA 0.123053f
C4151 VOUT-.n190 GNDA 0.03619f
C4152 VOUT-.n191 GNDA 0.186745f
C4153 VOUT-.n192 GNDA 0.03619f
C4154 VOUT-.n193 GNDA 0.03619f
C4155 VOUT-.n194 GNDA 0.03619f
C4156 VOUT-.n195 GNDA 0.03619f
C4157 VOUT-.n196 GNDA 0.07747f
C4158 VOUT-.n197 GNDA 0.097261f
.ends

