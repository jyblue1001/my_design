magic
tech sky130A
timestamp 1722808426
<< nwell >>
rect -90 205 170 395
<< nmos >>
rect 30 50 45 150
rect 85 50 100 150
<< pmos >>
rect 30 225 45 375
rect 85 225 100 375
<< ndiff >>
rect -20 130 30 150
rect -20 110 -5 130
rect 15 110 30 130
rect -20 90 30 110
rect -20 70 -5 90
rect 15 70 30 90
rect -20 50 30 70
rect 45 50 85 150
rect 100 130 150 150
rect 100 110 115 130
rect 135 110 150 130
rect 100 90 150 110
rect 100 70 115 90
rect 135 70 150 90
rect 100 50 150 70
<< pdiff >>
rect -20 345 30 375
rect -20 325 -5 345
rect 15 325 30 345
rect -20 305 30 325
rect -20 285 -5 305
rect 15 285 30 305
rect -20 265 30 285
rect -20 245 -5 265
rect 15 245 30 265
rect -20 225 30 245
rect 45 345 85 375
rect 45 325 55 345
rect 75 325 85 345
rect 45 305 85 325
rect 45 285 55 305
rect 75 285 85 305
rect 45 265 85 285
rect 45 245 55 265
rect 75 245 85 265
rect 45 225 85 245
rect 100 345 150 375
rect 100 325 115 345
rect 135 325 150 345
rect 100 305 150 325
rect 100 285 115 305
rect 135 285 150 305
rect 100 265 150 285
rect 100 245 115 265
rect 135 245 150 265
rect 100 225 150 245
<< ndiffc >>
rect -5 110 15 130
rect -5 70 15 90
rect 115 110 135 130
rect 115 70 135 90
<< pdiffc >>
rect -5 325 15 345
rect -5 285 15 305
rect -5 245 15 265
rect 55 325 75 345
rect 55 285 75 305
rect 55 245 75 265
rect 115 325 135 345
rect 115 285 135 305
rect 115 245 135 265
<< psubdiff >>
rect -60 130 -20 150
rect -60 110 -50 130
rect -30 110 -20 130
rect -60 90 -20 110
rect -60 70 -50 90
rect -30 70 -20 90
rect -60 50 -20 70
<< nsubdiff >>
rect -70 345 -20 375
rect -70 325 -50 345
rect -30 325 -20 345
rect -70 305 -20 325
rect -70 285 -50 305
rect -30 285 -20 305
rect -70 265 -20 285
rect -70 245 -50 265
rect -30 245 -20 265
rect -70 225 -20 245
<< psubdiffcont >>
rect -50 110 -30 130
rect -50 70 -30 90
<< nsubdiffcont >>
rect -50 325 -30 345
rect -50 285 -30 305
rect -50 245 -30 265
<< poly >>
rect 30 375 45 390
rect 85 375 100 390
rect 30 200 45 225
rect -10 190 45 200
rect -10 170 0 190
rect 20 170 45 190
rect -10 160 45 170
rect 30 150 45 160
rect 85 200 100 225
rect 85 190 140 200
rect 85 170 110 190
rect 130 170 140 190
rect 85 160 140 170
rect 85 150 100 160
rect 30 35 45 50
rect 85 35 100 50
<< polycont >>
rect 0 170 20 190
rect 110 170 130 190
<< locali >>
rect -60 385 -50 405
rect -30 385 -5 405
rect 15 385 55 405
rect 75 385 115 405
rect 135 385 160 405
rect -50 365 -30 385
rect 110 365 140 385
rect -60 345 20 365
rect -60 325 -50 345
rect -30 325 -5 345
rect 15 325 20 345
rect -60 305 20 325
rect -60 285 -50 305
rect -30 285 -5 305
rect 15 285 20 305
rect -60 265 20 285
rect -60 245 -50 265
rect -30 245 -5 265
rect 15 245 20 265
rect -60 230 20 245
rect 50 345 80 365
rect 50 325 55 345
rect 75 325 80 345
rect 50 305 80 325
rect 50 285 55 305
rect 75 285 80 305
rect 50 265 80 285
rect 50 245 55 265
rect 75 245 80 265
rect -10 190 30 200
rect -10 170 0 190
rect 20 170 30 190
rect -10 160 30 170
rect 50 140 80 245
rect 110 345 145 365
rect 110 325 115 345
rect 135 325 145 345
rect 110 305 145 325
rect 110 285 115 305
rect 135 285 145 305
rect 110 265 145 285
rect 110 245 115 265
rect 135 245 145 265
rect 110 235 145 245
rect 100 190 140 200
rect 100 170 110 190
rect 130 170 140 190
rect 100 160 140 170
rect -60 130 20 140
rect -60 110 -50 130
rect -30 110 -5 130
rect 15 110 20 130
rect -60 90 20 110
rect -60 70 -50 90
rect -30 70 -5 90
rect 15 70 20 90
rect -60 55 20 70
rect 50 130 140 140
rect 50 110 115 130
rect 135 110 140 130
rect 50 90 140 110
rect 50 70 115 90
rect 135 70 140 90
rect 50 60 140 70
rect -50 30 -30 55
rect -55 10 -50 30
rect -30 10 -5 30
rect 15 10 55 30
rect 75 10 115 30
rect 135 10 140 30
<< viali >>
rect -50 385 -30 405
rect -5 385 15 405
rect 55 385 75 405
rect 115 385 135 405
rect -50 10 -30 30
rect -5 10 15 30
rect 55 10 75 30
rect 115 10 135 30
<< metal1 >>
rect -70 405 165 425
rect -70 385 -50 405
rect -30 385 -5 405
rect 15 385 55 405
rect 75 385 115 405
rect 135 385 165 405
rect -70 365 165 385
rect -60 30 150 50
rect -60 10 -50 30
rect -30 10 -5 30
rect 15 10 55 30
rect 75 10 115 30
rect 135 10 150 30
rect -60 -10 150 10
<< end >>
