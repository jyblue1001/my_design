magic
tech sky130A
timestamp 1756070869
<< metal1 >>
rect 2070 19310 2190 19325
rect 2070 19280 2115 19310
rect 2145 19280 2190 19310
rect 2070 19245 2190 19280
rect 2070 19215 2115 19245
rect 2145 19215 2190 19245
rect 2070 19175 2190 19215
rect 2070 19145 2115 19175
rect 2145 19145 2190 19175
rect 2070 19105 2190 19145
rect 2070 19075 2115 19105
rect 2145 19075 2190 19105
rect 2070 19035 2190 19075
rect 2070 19005 2115 19035
rect 2145 19005 2190 19035
rect 2070 18970 2190 19005
rect 2070 18940 2115 18970
rect 2145 18940 2190 18970
rect 2070 18910 2190 18940
rect 2070 18880 2115 18910
rect 2145 18880 2190 18910
rect 2070 18845 2190 18880
rect 2070 18815 2115 18845
rect 2145 18815 2190 18845
rect 2070 18775 2190 18815
rect 2070 18745 2115 18775
rect 2145 18745 2190 18775
rect 2070 18705 2190 18745
rect 2070 18675 2115 18705
rect 2145 18675 2190 18705
rect 2070 18635 2190 18675
rect 2070 18605 2115 18635
rect 2145 18605 2190 18635
rect 2070 18570 2190 18605
rect 2070 18540 2115 18570
rect 2145 18540 2190 18570
rect 2070 18510 2190 18540
rect 2070 18480 2115 18510
rect 2145 18480 2190 18510
rect 2070 18445 2190 18480
rect 2070 18415 2115 18445
rect 2145 18415 2190 18445
rect 2070 18375 2190 18415
rect 2070 18345 2115 18375
rect 2145 18345 2190 18375
rect 2070 18305 2190 18345
rect 2070 18275 2115 18305
rect 2145 18275 2190 18305
rect 2070 18235 2190 18275
rect 2070 18205 2115 18235
rect 2145 18205 2190 18235
rect 2070 18170 2190 18205
rect 2070 18140 2115 18170
rect 2145 18140 2190 18170
rect 2070 18110 2190 18140
rect 2070 18080 2115 18110
rect 2145 18080 2190 18110
rect 2070 18045 2190 18080
rect 2070 18015 2115 18045
rect 2145 18015 2190 18045
rect 2070 17975 2190 18015
rect 2070 17945 2115 17975
rect 2145 17945 2190 17975
rect 2070 17905 2190 17945
rect 2070 17875 2115 17905
rect 2145 17875 2190 17905
rect 2070 17835 2190 17875
rect 2070 17805 2115 17835
rect 2145 17805 2190 17835
rect 2070 17770 2190 17805
rect 2070 17740 2115 17770
rect 2145 17740 2190 17770
rect 2070 15690 2190 17740
rect 6690 19310 6750 19325
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2070 15660 2075 15690
rect 2105 15660 2115 15690
rect 2145 15660 2155 15690
rect 2185 15660 2190 15690
rect 2070 15650 2190 15660
rect 2070 15620 2075 15650
rect 2105 15620 2115 15650
rect 2145 15620 2155 15650
rect 2185 15620 2190 15650
rect 2070 15610 2190 15620
rect 2070 15580 2075 15610
rect 2105 15580 2115 15610
rect 2145 15580 2155 15610
rect 2185 15580 2190 15610
rect 2070 12710 2190 15580
rect 2070 12680 2075 12710
rect 2105 12680 2115 12710
rect 2145 12680 2155 12710
rect 2185 12680 2190 12710
rect 2070 12670 2190 12680
rect 2070 12640 2075 12670
rect 2105 12640 2115 12670
rect 2145 12640 2155 12670
rect 2185 12640 2190 12670
rect 2070 12550 2190 12640
rect 2070 12520 2075 12550
rect 2105 12520 2115 12550
rect 2145 12520 2155 12550
rect 2185 12520 2190 12550
rect 2070 12510 2190 12520
rect 2070 12480 2075 12510
rect 2105 12480 2115 12510
rect 2145 12480 2155 12510
rect 2185 12480 2190 12510
rect 2070 12470 2190 12480
rect 2070 12440 2075 12470
rect 2105 12440 2115 12470
rect 2145 12440 2155 12470
rect 2185 12440 2190 12470
rect 2070 12435 2190 12440
rect 2205 15925 2325 15930
rect 2205 15895 2210 15925
rect 2240 15895 2250 15925
rect 2280 15895 2290 15925
rect 2320 15895 2325 15925
rect 1280 9635 1400 9650
rect 1280 9605 1325 9635
rect 1355 9605 1400 9635
rect 1280 9570 1400 9605
rect 1280 9540 1325 9570
rect 1355 9540 1400 9570
rect 1280 9500 1400 9540
rect 1280 9470 1325 9500
rect 1355 9470 1400 9500
rect 1280 9430 1400 9470
rect 1280 9400 1325 9430
rect 1355 9400 1400 9430
rect 1280 9360 1400 9400
rect 1280 9330 1325 9360
rect 1355 9330 1400 9360
rect 1280 9295 1400 9330
rect 1280 9265 1325 9295
rect 1355 9265 1400 9295
rect 1280 9235 1400 9265
rect 1280 9205 1325 9235
rect 1355 9205 1400 9235
rect 1280 9170 1400 9205
rect 1280 9140 1325 9170
rect 1355 9140 1400 9170
rect 1280 9100 1400 9140
rect 1280 9070 1325 9100
rect 1355 9070 1400 9100
rect 1280 9030 1400 9070
rect 1280 9000 1325 9030
rect 1355 9000 1400 9030
rect 1280 8960 1400 9000
rect 1280 8930 1325 8960
rect 1355 8930 1400 8960
rect 1280 8895 1400 8930
rect 1280 8865 1325 8895
rect 1355 8865 1400 8895
rect 1280 8835 1400 8865
rect 1280 8805 1325 8835
rect 1355 8805 1400 8835
rect 1280 8770 1400 8805
rect 1280 8740 1325 8770
rect 1355 8740 1400 8770
rect 1280 8700 1400 8740
rect 1280 8670 1325 8700
rect 1355 8670 1400 8700
rect 1280 8630 1400 8670
rect 1280 8600 1325 8630
rect 1355 8600 1400 8630
rect 1280 8560 1400 8600
rect 1280 8530 1325 8560
rect 1355 8530 1400 8560
rect 1280 8495 1400 8530
rect 1280 8465 1325 8495
rect 1355 8465 1400 8495
rect 1280 8435 1400 8465
rect 1280 8405 1325 8435
rect 1355 8405 1400 8435
rect 1280 8370 1400 8405
rect 1280 8340 1325 8370
rect 1355 8340 1400 8370
rect 1280 8300 1400 8340
rect 1280 8270 1325 8300
rect 1355 8270 1400 8300
rect 1280 8230 1400 8270
rect 1280 8200 1325 8230
rect 1355 8200 1400 8230
rect 1280 8160 1400 8200
rect 1280 8130 1325 8160
rect 1355 8130 1400 8160
rect 1280 6195 1400 8130
rect 2205 9635 2325 15895
rect 6660 15595 6780 17725
rect 6660 15565 6665 15595
rect 6695 15565 6705 15595
rect 6735 15565 6745 15595
rect 6775 15565 6780 15595
rect 6660 15555 6780 15565
rect 6660 15525 6665 15555
rect 6695 15525 6705 15555
rect 6735 15525 6745 15555
rect 6775 15525 6780 15555
rect 6660 15515 6780 15525
rect 6660 15485 6665 15515
rect 6695 15485 6705 15515
rect 6735 15485 6745 15515
rect 6775 15485 6780 15515
rect 2205 9605 2250 9635
rect 2280 9605 2325 9635
rect 2205 9570 2325 9605
rect 2205 9540 2250 9570
rect 2280 9540 2325 9570
rect 2205 9500 2325 9540
rect 2205 9470 2250 9500
rect 2280 9470 2325 9500
rect 2205 9430 2325 9470
rect 2205 9400 2250 9430
rect 2280 9400 2325 9430
rect 2205 9360 2325 9400
rect 2205 9330 2250 9360
rect 2280 9330 2325 9360
rect 2205 9295 2325 9330
rect 2205 9265 2250 9295
rect 2280 9265 2325 9295
rect 2205 9235 2325 9265
rect 2205 9205 2250 9235
rect 2280 9205 2325 9235
rect 2205 9170 2325 9205
rect 2205 9140 2250 9170
rect 2280 9140 2325 9170
rect 2205 9100 2325 9140
rect 2205 9070 2250 9100
rect 2280 9070 2325 9100
rect 2205 9030 2325 9070
rect 2205 9000 2250 9030
rect 2280 9000 2325 9030
rect 2205 8960 2325 9000
rect 2205 8930 2250 8960
rect 2280 8930 2325 8960
rect 2205 8895 2325 8930
rect 2205 8865 2250 8895
rect 2280 8865 2325 8895
rect 2205 8835 2325 8865
rect 2205 8805 2250 8835
rect 2280 8805 2325 8835
rect 2205 8770 2325 8805
rect 2205 8740 2250 8770
rect 2280 8740 2325 8770
rect 2205 8700 2325 8740
rect 2205 8670 2250 8700
rect 2280 8670 2325 8700
rect 2205 8630 2325 8670
rect 2205 8600 2250 8630
rect 2280 8600 2325 8630
rect 2205 8560 2325 8600
rect 2205 8530 2250 8560
rect 2280 8530 2325 8560
rect 2205 8495 2325 8530
rect 2205 8465 2250 8495
rect 2280 8465 2325 8495
rect 2205 8435 2325 8465
rect 2205 8405 2250 8435
rect 2280 8405 2325 8435
rect 2205 8370 2325 8405
rect 2205 8340 2250 8370
rect 2280 8340 2325 8370
rect 2205 8300 2325 8340
rect 2205 8270 2250 8300
rect 2280 8270 2325 8300
rect 2205 8230 2325 8270
rect 2205 8200 2250 8230
rect 2280 8200 2325 8230
rect 2205 8160 2325 8200
rect 2205 8130 2250 8160
rect 2280 8130 2325 8160
rect 2205 8105 2325 8130
rect 1980 8085 2100 8090
rect 1980 8055 1985 8085
rect 2015 8055 2025 8085
rect 2055 8055 2065 8085
rect 2095 8055 2100 8085
rect 1630 8030 1750 8035
rect 1630 8000 1635 8030
rect 1665 8000 1675 8030
rect 1705 8000 1715 8030
rect 1745 8000 1750 8030
rect 1630 6195 1750 8000
rect 1980 6195 2100 8055
rect 2475 8085 2515 13175
rect 2475 8055 2480 8085
rect 2510 8055 2515 8085
rect 2475 8050 2515 8055
rect 2725 6310 2745 9735
rect 2855 6420 2875 9735
rect 3175 7980 3215 10325
rect 3235 7980 3275 10325
rect 3165 7955 3280 7980
rect 3165 7925 3180 7955
rect 3210 7925 3240 7955
rect 3270 7925 3280 7955
rect 3165 7885 3280 7925
rect 3165 7855 3180 7885
rect 3210 7855 3240 7885
rect 3270 7855 3280 7885
rect 3165 7815 3280 7855
rect 3165 7785 3180 7815
rect 3210 7785 3240 7815
rect 3270 7785 3280 7815
rect 3165 7745 3280 7785
rect 3165 7715 3180 7745
rect 3210 7715 3240 7745
rect 3270 7715 3280 7745
rect 3165 7680 3280 7715
rect 3165 7650 3180 7680
rect 3210 7650 3240 7680
rect 3270 7650 3280 7680
rect 3165 7620 3280 7650
rect 3165 7590 3180 7620
rect 3210 7590 3240 7620
rect 3270 7590 3280 7620
rect 3165 7555 3280 7590
rect 3165 7525 3180 7555
rect 3210 7525 3240 7555
rect 3270 7525 3280 7555
rect 3165 7485 3280 7525
rect 3165 7455 3180 7485
rect 3210 7455 3240 7485
rect 3270 7455 3280 7485
rect 3165 7415 3280 7455
rect 3165 7385 3180 7415
rect 3210 7385 3240 7415
rect 3270 7385 3280 7415
rect 3165 7345 3280 7385
rect 3165 7315 3180 7345
rect 3210 7315 3240 7345
rect 3270 7315 3280 7345
rect 3165 7280 3280 7315
rect 3165 7250 3180 7280
rect 3210 7250 3240 7280
rect 3270 7250 3280 7280
rect 3165 7220 3280 7250
rect 3165 7190 3180 7220
rect 3210 7190 3240 7220
rect 3270 7190 3280 7220
rect 3165 7155 3280 7190
rect 3165 7125 3180 7155
rect 3210 7125 3240 7155
rect 3270 7125 3280 7155
rect 3165 7085 3280 7125
rect 3165 7055 3180 7085
rect 3210 7055 3240 7085
rect 3270 7055 3280 7085
rect 3165 7015 3280 7055
rect 3165 6985 3180 7015
rect 3210 6985 3240 7015
rect 3270 6985 3280 7015
rect 3165 6945 3280 6985
rect 3165 6915 3180 6945
rect 3210 6915 3240 6945
rect 3270 6915 3280 6945
rect 3165 6880 3280 6915
rect 3165 6850 3180 6880
rect 3210 6850 3240 6880
rect 3270 6850 3280 6880
rect 3165 6820 3280 6850
rect 3165 6790 3180 6820
rect 3210 6790 3240 6820
rect 3270 6790 3280 6820
rect 3165 6755 3280 6790
rect 3165 6725 3180 6755
rect 3210 6725 3240 6755
rect 3270 6725 3280 6755
rect 3165 6685 3280 6725
rect 3165 6655 3180 6685
rect 3210 6655 3240 6685
rect 3270 6655 3280 6685
rect 3165 6615 3280 6655
rect 3165 6585 3180 6615
rect 3210 6585 3240 6615
rect 3270 6585 3280 6615
rect 3165 6545 3280 6585
rect 3165 6515 3180 6545
rect 3210 6515 3240 6545
rect 3270 6515 3280 6545
rect 3165 6480 3280 6515
rect 3165 6450 3180 6480
rect 3210 6450 3240 6480
rect 3270 6450 3280 6480
rect 3165 6435 3280 6450
rect 2845 6415 2885 6420
rect 2845 6385 2850 6415
rect 2880 6385 2885 6415
rect 2845 6380 2885 6385
rect 2715 6305 2755 6310
rect 2715 6275 2720 6305
rect 2750 6275 2755 6305
rect 2715 6270 2755 6275
rect 3075 6305 3115 6310
rect 3295 6305 3325 9740
rect 3345 7980 3385 10325
rect 3630 8030 3670 9735
rect 3630 8000 3635 8030
rect 3665 8000 3670 8030
rect 3630 7995 3670 8000
rect 3850 8030 3890 9735
rect 3850 8000 3855 8030
rect 3885 8000 3890 8030
rect 3850 7995 3890 8000
rect 3340 7955 3390 7980
rect 3340 7925 3350 7955
rect 3380 7925 3390 7955
rect 3340 7885 3390 7925
rect 3340 7855 3350 7885
rect 3380 7855 3390 7885
rect 3340 7815 3390 7855
rect 3340 7785 3350 7815
rect 3380 7785 3390 7815
rect 3340 7745 3390 7785
rect 3340 7715 3350 7745
rect 3380 7715 3390 7745
rect 3340 7680 3390 7715
rect 3340 7650 3350 7680
rect 3380 7650 3390 7680
rect 3340 7620 3390 7650
rect 3340 7590 3350 7620
rect 3380 7590 3390 7620
rect 3340 7555 3390 7590
rect 3340 7525 3350 7555
rect 3380 7525 3390 7555
rect 3340 7485 3390 7525
rect 3340 7455 3350 7485
rect 3380 7455 3390 7485
rect 3340 7415 3390 7455
rect 3340 7385 3350 7415
rect 3380 7385 3390 7415
rect 3340 7345 3390 7385
rect 3340 7315 3350 7345
rect 3380 7315 3390 7345
rect 3340 7280 3390 7315
rect 3340 7250 3350 7280
rect 3380 7250 3390 7280
rect 3340 7220 3390 7250
rect 3340 7190 3350 7220
rect 3380 7190 3390 7220
rect 3340 7155 3390 7190
rect 3340 7125 3350 7155
rect 3380 7125 3390 7155
rect 3340 7085 3390 7125
rect 3340 7055 3350 7085
rect 3380 7055 3390 7085
rect 3340 7015 3390 7055
rect 3340 6985 3350 7015
rect 3380 6985 3390 7015
rect 3340 6945 3390 6985
rect 3340 6915 3350 6945
rect 3380 6915 3390 6945
rect 3340 6880 3390 6915
rect 3340 6850 3350 6880
rect 3380 6850 3390 6880
rect 3340 6820 3390 6850
rect 3340 6790 3350 6820
rect 3380 6790 3390 6820
rect 3340 6755 3390 6790
rect 3340 6725 3350 6755
rect 3380 6725 3390 6755
rect 3340 6685 3390 6725
rect 3340 6655 3350 6685
rect 3380 6655 3390 6685
rect 3340 6615 3390 6655
rect 3340 6585 3350 6615
rect 3380 6585 3390 6615
rect 3340 6545 3390 6585
rect 3340 6515 3350 6545
rect 3380 6515 3390 6545
rect 3340 6480 3390 6515
rect 3340 6450 3350 6480
rect 3380 6450 3390 6480
rect 3340 6435 3390 6450
rect 3380 6415 3420 6420
rect 3380 6385 3385 6415
rect 3415 6385 3420 6415
rect 3380 6380 3420 6385
rect 3075 6275 3080 6305
rect 3110 6275 3115 6305
rect 3075 6270 3115 6275
rect 3290 6300 3330 6305
rect 3290 6270 3295 6300
rect 3325 6270 3330 6300
rect 930 6190 1050 6195
rect 930 6160 935 6190
rect 965 6160 975 6190
rect 1005 6160 1015 6190
rect 1045 6160 1050 6190
rect 930 6150 1050 6160
rect 930 6120 935 6150
rect 965 6120 975 6150
rect 1005 6120 1015 6150
rect 1045 6120 1050 6150
rect 930 6110 1050 6120
rect 930 6080 935 6110
rect 965 6080 975 6110
rect 1005 6080 1015 6110
rect 1045 6080 1050 6110
rect 930 1145 1050 6080
rect 3085 5080 3105 6270
rect 3290 6265 3330 6270
rect 3075 5075 3115 5080
rect 3075 5045 3080 5075
rect 3110 5045 3115 5075
rect 3075 5040 3115 5045
rect 3390 3795 3410 6380
rect 3435 6245 3475 6250
rect 3435 6215 3440 6245
rect 3470 6215 3475 6245
rect 3380 3790 3420 3795
rect 3380 3760 3385 3790
rect 3415 3760 3420 3790
rect 3380 3755 3420 3760
rect 3435 3110 3475 6215
rect 4310 6190 4340 9740
rect 4310 6150 4340 6160
rect 4310 6110 4340 6120
rect 4310 6075 4340 6080
rect 4420 6190 4450 9740
rect 4470 6300 4510 6305
rect 4470 6270 4475 6300
rect 4505 6270 4510 6300
rect 4470 6245 4510 6270
rect 4470 6215 4475 6245
rect 4505 6215 4510 6245
rect 4470 6210 4510 6215
rect 4420 6150 4450 6160
rect 4420 6110 4450 6120
rect 4420 6075 4450 6080
rect 4530 6190 4560 9740
rect 4530 6150 4560 6160
rect 4530 6110 4560 6120
rect 4530 6075 4560 6080
rect 4640 6190 4670 9740
rect 5310 8015 5350 9735
rect 5310 7985 5315 8015
rect 5345 7985 5350 8015
rect 5310 7980 5350 7985
rect 6155 6420 6175 9740
rect 5470 6415 5510 6420
rect 5470 6385 5475 6415
rect 5505 6385 5510 6415
rect 5470 6380 5510 6385
rect 6145 6415 6185 6420
rect 6145 6385 6150 6415
rect 6180 6385 6185 6415
rect 6145 6380 6185 6385
rect 4640 6150 4670 6160
rect 4640 6110 4670 6120
rect 4640 6075 4670 6080
rect 5480 3855 5500 6380
rect 5545 6245 5585 6250
rect 5545 6215 5550 6245
rect 5580 6215 5585 6245
rect 5475 3850 5505 3855
rect 5475 3815 5505 3820
rect 3435 3080 3440 3110
rect 3470 3080 3475 3110
rect 3435 3075 3475 3080
rect 4470 3110 4510 3115
rect 4470 3080 4475 3110
rect 4505 3080 4510 3110
rect 4470 2890 4510 3080
rect 5545 3110 5585 6215
rect 5870 5420 5910 5425
rect 5870 5390 5875 5420
rect 5905 5390 5910 5420
rect 5620 5020 5660 5025
rect 5620 4990 5625 5020
rect 5655 4990 5660 5020
rect 5620 4425 5660 4990
rect 5870 5020 5910 5390
rect 6220 5420 6260 13120
rect 6465 8070 6505 13175
rect 6660 12925 6780 15485
rect 6660 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6745 12925
rect 6775 12895 6780 12925
rect 6660 12885 6780 12895
rect 6660 12855 6665 12885
rect 6695 12855 6705 12885
rect 6735 12855 6745 12885
rect 6775 12855 6780 12885
rect 6660 12845 6780 12855
rect 6660 12815 6665 12845
rect 6695 12815 6705 12845
rect 6735 12815 6745 12845
rect 6775 12815 6780 12845
rect 6660 12810 6780 12815
rect 6660 12150 6780 12155
rect 6660 12120 6665 12150
rect 6695 12120 6705 12150
rect 6735 12120 6745 12150
rect 6775 12120 6780 12150
rect 6660 12110 6780 12120
rect 6660 12080 6665 12110
rect 6695 12080 6705 12110
rect 6735 12080 6745 12110
rect 6775 12080 6780 12110
rect 6660 12070 6780 12080
rect 6660 12040 6665 12070
rect 6695 12040 6705 12070
rect 6735 12040 6745 12070
rect 6775 12040 6780 12070
rect 6660 11165 6780 12040
rect 6660 11135 6665 11165
rect 6695 11135 6705 11165
rect 6735 11135 6745 11165
rect 6775 11135 6780 11165
rect 6660 11125 6780 11135
rect 6660 11095 6665 11125
rect 6695 11095 6705 11125
rect 6735 11095 6745 11125
rect 6775 11095 6780 11125
rect 6660 11085 6780 11095
rect 6660 11055 6665 11085
rect 6695 11055 6705 11085
rect 6735 11055 6745 11085
rect 6775 11055 6780 11085
rect 6660 10440 6780 11055
rect 6660 10410 6665 10440
rect 6695 10410 6705 10440
rect 6735 10410 6745 10440
rect 6775 10410 6780 10440
rect 6660 10400 6780 10410
rect 6660 10370 6665 10400
rect 6695 10370 6705 10400
rect 6735 10370 6745 10400
rect 6775 10370 6780 10400
rect 6660 10360 6780 10370
rect 6660 10330 6665 10360
rect 6695 10330 6705 10360
rect 6735 10330 6745 10360
rect 6775 10330 6780 10360
rect 6660 10080 6780 10330
rect 6660 10050 6665 10080
rect 6695 10050 6705 10080
rect 6735 10050 6745 10080
rect 6775 10050 6780 10080
rect 6660 10040 6780 10050
rect 6660 10010 6665 10040
rect 6695 10010 6705 10040
rect 6735 10010 6745 10040
rect 6775 10010 6780 10040
rect 6660 10000 6780 10010
rect 6660 9970 6665 10000
rect 6695 9970 6705 10000
rect 6735 9970 6745 10000
rect 6775 9970 6780 10000
rect 6660 9570 6780 9970
rect 6660 9540 6705 9570
rect 6735 9540 6780 9570
rect 6660 9500 6780 9540
rect 6660 9470 6705 9500
rect 6735 9470 6780 9500
rect 6660 9430 6780 9470
rect 6660 9400 6705 9430
rect 6735 9400 6780 9430
rect 6660 9360 6780 9400
rect 6660 9330 6705 9360
rect 6735 9330 6780 9360
rect 6660 9295 6780 9330
rect 6660 9265 6705 9295
rect 6735 9265 6780 9295
rect 6660 9235 6780 9265
rect 6660 9205 6705 9235
rect 6735 9205 6780 9235
rect 6660 9170 6780 9205
rect 6660 9140 6705 9170
rect 6735 9140 6780 9170
rect 6660 9100 6780 9140
rect 6660 9070 6705 9100
rect 6735 9070 6780 9100
rect 6660 9030 6780 9070
rect 6660 9000 6705 9030
rect 6735 9000 6780 9030
rect 6660 8960 6780 9000
rect 6660 8930 6705 8960
rect 6735 8930 6780 8960
rect 6660 8895 6780 8930
rect 6660 8865 6705 8895
rect 6735 8865 6780 8895
rect 6660 8835 6780 8865
rect 6660 8805 6705 8835
rect 6735 8805 6780 8835
rect 6660 8770 6780 8805
rect 6660 8740 6705 8770
rect 6735 8740 6780 8770
rect 6660 8700 6780 8740
rect 6660 8670 6705 8700
rect 6735 8670 6780 8700
rect 6660 8630 6780 8670
rect 6660 8600 6705 8630
rect 6735 8600 6780 8630
rect 6660 8560 6780 8600
rect 6660 8530 6705 8560
rect 6735 8530 6780 8560
rect 6660 8495 6780 8530
rect 6660 8465 6705 8495
rect 6735 8465 6780 8495
rect 6660 8435 6780 8465
rect 6660 8405 6705 8435
rect 6735 8405 6780 8435
rect 6660 8370 6780 8405
rect 6660 8340 6705 8370
rect 6735 8340 6780 8370
rect 6660 8300 6780 8340
rect 6660 8270 6705 8300
rect 6735 8270 6780 8300
rect 6660 8230 6780 8270
rect 6660 8200 6705 8230
rect 6735 8200 6780 8230
rect 6660 8160 6780 8200
rect 6660 8130 6705 8160
rect 6735 8130 6780 8160
rect 6660 8105 6780 8130
rect 7580 9635 7700 9650
rect 7580 9605 7625 9635
rect 7655 9605 7700 9635
rect 7580 9570 7700 9605
rect 7580 9540 7625 9570
rect 7655 9540 7700 9570
rect 7580 9500 7700 9540
rect 7580 9470 7625 9500
rect 7655 9470 7700 9500
rect 7580 9430 7700 9470
rect 7580 9400 7625 9430
rect 7655 9400 7700 9430
rect 7580 9360 7700 9400
rect 7580 9330 7625 9360
rect 7655 9330 7700 9360
rect 7580 9295 7700 9330
rect 7580 9265 7625 9295
rect 7655 9265 7700 9295
rect 7580 9235 7700 9265
rect 7580 9205 7625 9235
rect 7655 9205 7700 9235
rect 7580 9170 7700 9205
rect 7580 9140 7625 9170
rect 7655 9140 7700 9170
rect 7580 9100 7700 9140
rect 7580 9070 7625 9100
rect 7655 9070 7700 9100
rect 7580 9030 7700 9070
rect 7580 9000 7625 9030
rect 7655 9000 7700 9030
rect 7580 8960 7700 9000
rect 7580 8930 7625 8960
rect 7655 8930 7700 8960
rect 7580 8895 7700 8930
rect 7580 8865 7625 8895
rect 7655 8865 7700 8895
rect 7580 8835 7700 8865
rect 7580 8805 7625 8835
rect 7655 8805 7700 8835
rect 7580 8770 7700 8805
rect 7580 8740 7625 8770
rect 7655 8740 7700 8770
rect 7580 8700 7700 8740
rect 7580 8670 7625 8700
rect 7655 8670 7700 8700
rect 7580 8630 7700 8670
rect 7580 8600 7625 8630
rect 7655 8600 7700 8630
rect 7580 8560 7700 8600
rect 7580 8530 7625 8560
rect 7655 8530 7700 8560
rect 7580 8495 7700 8530
rect 7580 8465 7625 8495
rect 7655 8465 7700 8495
rect 7580 8435 7700 8465
rect 7580 8405 7625 8435
rect 7655 8405 7700 8435
rect 7580 8370 7700 8405
rect 7580 8340 7625 8370
rect 7655 8340 7700 8370
rect 7580 8300 7700 8340
rect 7580 8270 7625 8300
rect 7655 8270 7700 8300
rect 7580 8230 7700 8270
rect 7580 8200 7625 8230
rect 7655 8200 7700 8230
rect 7580 8160 7700 8200
rect 7580 8130 7625 8160
rect 7655 8130 7700 8160
rect 6465 8040 6470 8070
rect 6500 8040 6505 8070
rect 6465 8035 6505 8040
rect 6880 8070 7000 8075
rect 6880 8040 6885 8070
rect 6915 8040 6925 8070
rect 6955 8040 6965 8070
rect 6995 8040 7000 8070
rect 6880 6195 7000 8040
rect 7230 8015 7350 8020
rect 7230 7985 7235 8015
rect 7265 7985 7275 8015
rect 7305 7985 7315 8015
rect 7345 7985 7350 8015
rect 7230 6195 7350 7985
rect 7580 6195 7700 8130
rect 6220 5390 6225 5420
rect 6255 5390 6260 5420
rect 6220 5385 6260 5390
rect 7930 6190 8050 6195
rect 7930 6160 7935 6190
rect 7965 6160 7975 6190
rect 8005 6160 8015 6190
rect 8045 6160 8050 6190
rect 7930 6150 8050 6160
rect 7930 6120 7935 6150
rect 7965 6120 7975 6150
rect 8005 6120 8015 6150
rect 8045 6120 8050 6150
rect 7930 6110 8050 6120
rect 7930 6080 7935 6110
rect 7965 6080 7975 6110
rect 8005 6080 8015 6110
rect 8045 6080 8050 6110
rect 5870 4990 5875 5020
rect 5905 4990 5910 5020
rect 5870 4985 5910 4990
rect 5620 4395 5625 4425
rect 5655 4395 5660 4425
rect 5620 4390 5660 4395
rect 5545 3080 5550 3110
rect 5580 3080 5585 3110
rect 5545 3075 5585 3080
rect 4470 2860 4475 2890
rect 4505 2860 4510 2890
rect 4470 2855 4510 2860
rect 930 1115 935 1145
rect 965 1115 975 1145
rect 1005 1115 1015 1145
rect 1045 1115 1050 1145
rect 930 1105 1050 1115
rect 930 1075 935 1105
rect 965 1075 975 1105
rect 1005 1075 1015 1105
rect 1045 1075 1050 1105
rect 930 1065 1050 1075
rect 930 1035 935 1065
rect 965 1035 975 1065
rect 1005 1035 1015 1065
rect 1045 1035 1050 1065
rect 930 1030 1050 1035
rect 4415 1145 4455 1150
rect 4415 1115 4420 1145
rect 4450 1115 4455 1145
rect 4415 1105 4455 1115
rect 4415 1075 4420 1105
rect 4450 1075 4455 1105
rect 4415 1065 4455 1075
rect 4415 1035 4420 1065
rect 4450 1035 4455 1065
rect 4415 1030 4455 1035
rect 4525 1145 4565 1150
rect 4525 1115 4530 1145
rect 4560 1115 4565 1145
rect 4525 1105 4565 1115
rect 4525 1075 4530 1105
rect 4560 1075 4565 1105
rect 4525 1065 4565 1075
rect 4525 1035 4530 1065
rect 4560 1035 4565 1065
rect 4525 1030 4565 1035
rect 7930 1145 8050 6080
rect 7930 1115 7935 1145
rect 7965 1115 7975 1145
rect 8005 1115 8015 1145
rect 8045 1115 8050 1145
rect 7930 1105 8050 1115
rect 7930 1075 7935 1105
rect 7965 1075 7975 1105
rect 8005 1075 8015 1105
rect 8045 1075 8050 1105
rect 7930 1065 8050 1075
rect 7930 1035 7935 1065
rect 7965 1035 7975 1065
rect 8005 1035 8015 1065
rect 8045 1035 8050 1065
rect 7930 1030 8050 1035
rect -120 -1320 0 -1225
rect -120 -1350 -75 -1320
rect -45 -1350 0 -1320
rect -120 -1385 0 -1350
rect -120 -1415 -75 -1385
rect -45 -1415 0 -1385
rect -120 -1455 0 -1415
rect -120 -1485 -75 -1455
rect -45 -1485 0 -1455
rect -120 -1525 0 -1485
rect -120 -1555 -75 -1525
rect -45 -1555 0 -1525
rect -120 -1595 0 -1555
rect -120 -1625 -75 -1595
rect -45 -1625 0 -1595
rect -120 -1660 0 -1625
rect -120 -1690 -75 -1660
rect -45 -1690 0 -1660
rect -120 -1720 0 -1690
rect -120 -1750 -75 -1720
rect -45 -1750 0 -1720
rect -120 -1785 0 -1750
rect -120 -1815 -75 -1785
rect -45 -1815 0 -1785
rect -120 -1855 0 -1815
rect -120 -1885 -75 -1855
rect -45 -1885 0 -1855
rect -120 -1925 0 -1885
rect -120 -1955 -75 -1925
rect -45 -1955 0 -1925
rect -120 -1995 0 -1955
rect -120 -2025 -75 -1995
rect -45 -2025 0 -1995
rect -120 -2060 0 -2025
rect -120 -2090 -75 -2060
rect -45 -2090 0 -2060
rect -120 -2120 0 -2090
rect -120 -2150 -75 -2120
rect -45 -2150 0 -2120
rect -120 -2185 0 -2150
rect -120 -2215 -75 -2185
rect -45 -2215 0 -2185
rect -120 -2255 0 -2215
rect -120 -2285 -75 -2255
rect -45 -2285 0 -2255
rect -120 -2325 0 -2285
rect -120 -2355 -75 -2325
rect -45 -2355 0 -2325
rect -120 -2395 0 -2355
rect -120 -2425 -75 -2395
rect -45 -2425 0 -2395
rect -120 -2460 0 -2425
rect -120 -2490 -75 -2460
rect -45 -2490 0 -2460
rect -120 -2520 0 -2490
rect -120 -2550 -75 -2520
rect -45 -2550 0 -2520
rect -120 -2585 0 -2550
rect -120 -2615 -75 -2585
rect -45 -2615 0 -2585
rect -120 -2655 0 -2615
rect -120 -2685 -75 -2655
rect -45 -2685 0 -2655
rect -120 -2725 0 -2685
rect -120 -2755 -75 -2725
rect -45 -2755 0 -2725
rect -120 -2795 0 -2755
rect -120 -2825 -75 -2795
rect -45 -2825 0 -2795
rect -120 -2860 0 -2825
rect -120 -2890 -75 -2860
rect -45 -2890 0 -2860
rect -120 -2905 0 -2890
rect 230 -1320 350 -1225
rect 230 -1350 275 -1320
rect 305 -1350 350 -1320
rect 230 -1385 350 -1350
rect 230 -1415 275 -1385
rect 305 -1415 350 -1385
rect 230 -1455 350 -1415
rect 230 -1485 275 -1455
rect 305 -1485 350 -1455
rect 230 -1525 350 -1485
rect 230 -1555 275 -1525
rect 305 -1555 350 -1525
rect 230 -1595 350 -1555
rect 230 -1625 275 -1595
rect 305 -1625 350 -1595
rect 230 -1660 350 -1625
rect 230 -1690 275 -1660
rect 305 -1690 350 -1660
rect 230 -1720 350 -1690
rect 230 -1750 275 -1720
rect 305 -1750 350 -1720
rect 230 -1785 350 -1750
rect 230 -1815 275 -1785
rect 305 -1815 350 -1785
rect 230 -1855 350 -1815
rect 230 -1885 275 -1855
rect 305 -1885 350 -1855
rect 230 -1925 350 -1885
rect 230 -1955 275 -1925
rect 305 -1955 350 -1925
rect 230 -1995 350 -1955
rect 230 -2025 275 -1995
rect 305 -2025 350 -1995
rect 230 -2060 350 -2025
rect 230 -2090 275 -2060
rect 305 -2090 350 -2060
rect 230 -2120 350 -2090
rect 230 -2150 275 -2120
rect 305 -2150 350 -2120
rect 230 -2185 350 -2150
rect 230 -2215 275 -2185
rect 305 -2215 350 -2185
rect 230 -2255 350 -2215
rect 230 -2285 275 -2255
rect 305 -2285 350 -2255
rect 230 -2325 350 -2285
rect 230 -2355 275 -2325
rect 305 -2355 350 -2325
rect 230 -2395 350 -2355
rect 230 -2425 275 -2395
rect 305 -2425 350 -2395
rect 230 -2460 350 -2425
rect 230 -2490 275 -2460
rect 305 -2490 350 -2460
rect 230 -2520 350 -2490
rect 230 -2550 275 -2520
rect 305 -2550 350 -2520
rect 230 -2585 350 -2550
rect 230 -2615 275 -2585
rect 305 -2615 350 -2585
rect 230 -2655 350 -2615
rect 230 -2685 275 -2655
rect 305 -2685 350 -2655
rect 230 -2725 350 -2685
rect 230 -2755 275 -2725
rect 305 -2755 350 -2725
rect 230 -2795 350 -2755
rect 230 -2825 275 -2795
rect 305 -2825 350 -2795
rect 230 -2860 350 -2825
rect 230 -2890 275 -2860
rect 305 -2890 350 -2860
rect 230 -2905 350 -2890
rect 580 -1320 700 -1225
rect 580 -1350 625 -1320
rect 655 -1350 700 -1320
rect 580 -1385 700 -1350
rect 580 -1415 625 -1385
rect 655 -1415 700 -1385
rect 580 -1455 700 -1415
rect 580 -1485 625 -1455
rect 655 -1485 700 -1455
rect 580 -1525 700 -1485
rect 580 -1555 625 -1525
rect 655 -1555 700 -1525
rect 580 -1595 700 -1555
rect 580 -1625 625 -1595
rect 655 -1625 700 -1595
rect 580 -1660 700 -1625
rect 580 -1690 625 -1660
rect 655 -1690 700 -1660
rect 580 -1720 700 -1690
rect 580 -1750 625 -1720
rect 655 -1750 700 -1720
rect 580 -1785 700 -1750
rect 580 -1815 625 -1785
rect 655 -1815 700 -1785
rect 580 -1855 700 -1815
rect 580 -1885 625 -1855
rect 655 -1885 700 -1855
rect 580 -1925 700 -1885
rect 580 -1955 625 -1925
rect 655 -1955 700 -1925
rect 580 -1995 700 -1955
rect 580 -2025 625 -1995
rect 655 -2025 700 -1995
rect 580 -2060 700 -2025
rect 580 -2090 625 -2060
rect 655 -2090 700 -2060
rect 580 -2120 700 -2090
rect 580 -2150 625 -2120
rect 655 -2150 700 -2120
rect 580 -2185 700 -2150
rect 580 -2215 625 -2185
rect 655 -2215 700 -2185
rect 580 -2255 700 -2215
rect 580 -2285 625 -2255
rect 655 -2285 700 -2255
rect 580 -2325 700 -2285
rect 580 -2355 625 -2325
rect 655 -2355 700 -2325
rect 580 -2395 700 -2355
rect 580 -2425 625 -2395
rect 655 -2425 700 -2395
rect 580 -2460 700 -2425
rect 580 -2490 625 -2460
rect 655 -2490 700 -2460
rect 580 -2520 700 -2490
rect 580 -2550 625 -2520
rect 655 -2550 700 -2520
rect 580 -2585 700 -2550
rect 580 -2615 625 -2585
rect 655 -2615 700 -2585
rect 580 -2655 700 -2615
rect 580 -2685 625 -2655
rect 655 -2685 700 -2655
rect 580 -2725 700 -2685
rect 580 -2755 625 -2725
rect 655 -2755 700 -2725
rect 580 -2795 700 -2755
rect 580 -2825 625 -2795
rect 655 -2825 700 -2795
rect 580 -2860 700 -2825
rect 580 -2890 625 -2860
rect 655 -2890 700 -2860
rect 580 -2905 700 -2890
rect 930 -1320 1050 -1225
rect 930 -1350 975 -1320
rect 1005 -1350 1050 -1320
rect 930 -1385 1050 -1350
rect 930 -1415 975 -1385
rect 1005 -1415 1050 -1385
rect 930 -1455 1050 -1415
rect 930 -1485 975 -1455
rect 1005 -1485 1050 -1455
rect 930 -1525 1050 -1485
rect 930 -1555 975 -1525
rect 1005 -1555 1050 -1525
rect 930 -1595 1050 -1555
rect 930 -1625 975 -1595
rect 1005 -1625 1050 -1595
rect 930 -1660 1050 -1625
rect 930 -1690 975 -1660
rect 1005 -1690 1050 -1660
rect 930 -1720 1050 -1690
rect 930 -1750 975 -1720
rect 1005 -1750 1050 -1720
rect 930 -1785 1050 -1750
rect 930 -1815 975 -1785
rect 1005 -1815 1050 -1785
rect 930 -1855 1050 -1815
rect 930 -1885 975 -1855
rect 1005 -1885 1050 -1855
rect 930 -1925 1050 -1885
rect 930 -1955 975 -1925
rect 1005 -1955 1050 -1925
rect 930 -1995 1050 -1955
rect 930 -2025 975 -1995
rect 1005 -2025 1050 -1995
rect 930 -2060 1050 -2025
rect 930 -2090 975 -2060
rect 1005 -2090 1050 -2060
rect 930 -2120 1050 -2090
rect 930 -2150 975 -2120
rect 1005 -2150 1050 -2120
rect 930 -2185 1050 -2150
rect 930 -2215 975 -2185
rect 1005 -2215 1050 -2185
rect 930 -2255 1050 -2215
rect 930 -2285 975 -2255
rect 1005 -2285 1050 -2255
rect 930 -2325 1050 -2285
rect 930 -2355 975 -2325
rect 1005 -2355 1050 -2325
rect 930 -2395 1050 -2355
rect 930 -2425 975 -2395
rect 1005 -2425 1050 -2395
rect 930 -2460 1050 -2425
rect 930 -2490 975 -2460
rect 1005 -2490 1050 -2460
rect 930 -2520 1050 -2490
rect 930 -2550 975 -2520
rect 1005 -2550 1050 -2520
rect 930 -2585 1050 -2550
rect 930 -2615 975 -2585
rect 1005 -2615 1050 -2585
rect 930 -2655 1050 -2615
rect 930 -2685 975 -2655
rect 1005 -2685 1050 -2655
rect 930 -2725 1050 -2685
rect 930 -2755 975 -2725
rect 1005 -2755 1050 -2725
rect 930 -2795 1050 -2755
rect 930 -2825 975 -2795
rect 1005 -2825 1050 -2795
rect 930 -2860 1050 -2825
rect 930 -2890 975 -2860
rect 1005 -2890 1050 -2860
rect 930 -2905 1050 -2890
rect 1280 -1320 1400 -1225
rect 1280 -1350 1325 -1320
rect 1355 -1350 1400 -1320
rect 1280 -1385 1400 -1350
rect 1280 -1415 1325 -1385
rect 1355 -1415 1400 -1385
rect 1280 -1455 1400 -1415
rect 1280 -1485 1325 -1455
rect 1355 -1485 1400 -1455
rect 1280 -1525 1400 -1485
rect 1280 -1555 1325 -1525
rect 1355 -1555 1400 -1525
rect 1280 -1595 1400 -1555
rect 1280 -1625 1325 -1595
rect 1355 -1625 1400 -1595
rect 1280 -1660 1400 -1625
rect 1280 -1690 1325 -1660
rect 1355 -1690 1400 -1660
rect 1280 -1720 1400 -1690
rect 1280 -1750 1325 -1720
rect 1355 -1750 1400 -1720
rect 1280 -1785 1400 -1750
rect 1280 -1815 1325 -1785
rect 1355 -1815 1400 -1785
rect 1280 -1855 1400 -1815
rect 1280 -1885 1325 -1855
rect 1355 -1885 1400 -1855
rect 1280 -1925 1400 -1885
rect 1280 -1955 1325 -1925
rect 1355 -1955 1400 -1925
rect 1280 -1995 1400 -1955
rect 1280 -2025 1325 -1995
rect 1355 -2025 1400 -1995
rect 1280 -2060 1400 -2025
rect 1280 -2090 1325 -2060
rect 1355 -2090 1400 -2060
rect 1280 -2120 1400 -2090
rect 1280 -2150 1325 -2120
rect 1355 -2150 1400 -2120
rect 1280 -2185 1400 -2150
rect 1280 -2215 1325 -2185
rect 1355 -2215 1400 -2185
rect 1280 -2255 1400 -2215
rect 1280 -2285 1325 -2255
rect 1355 -2285 1400 -2255
rect 1280 -2325 1400 -2285
rect 1280 -2355 1325 -2325
rect 1355 -2355 1400 -2325
rect 1280 -2395 1400 -2355
rect 1280 -2425 1325 -2395
rect 1355 -2425 1400 -2395
rect 1280 -2460 1400 -2425
rect 1280 -2490 1325 -2460
rect 1355 -2490 1400 -2460
rect 1280 -2520 1400 -2490
rect 1280 -2550 1325 -2520
rect 1355 -2550 1400 -2520
rect 1280 -2585 1400 -2550
rect 1280 -2615 1325 -2585
rect 1355 -2615 1400 -2585
rect 1280 -2655 1400 -2615
rect 1280 -2685 1325 -2655
rect 1355 -2685 1400 -2655
rect 1280 -2725 1400 -2685
rect 1280 -2755 1325 -2725
rect 1355 -2755 1400 -2725
rect 1280 -2795 1400 -2755
rect 1280 -2825 1325 -2795
rect 1355 -2825 1400 -2795
rect 1280 -2860 1400 -2825
rect 1280 -2890 1325 -2860
rect 1355 -2890 1400 -2860
rect 1280 -2905 1400 -2890
rect 1630 -1320 1750 -1225
rect 1630 -1350 1675 -1320
rect 1705 -1350 1750 -1320
rect 1630 -1385 1750 -1350
rect 1630 -1415 1675 -1385
rect 1705 -1415 1750 -1385
rect 1630 -1455 1750 -1415
rect 1630 -1485 1675 -1455
rect 1705 -1485 1750 -1455
rect 1630 -1525 1750 -1485
rect 1630 -1555 1675 -1525
rect 1705 -1555 1750 -1525
rect 1630 -1595 1750 -1555
rect 1630 -1625 1675 -1595
rect 1705 -1625 1750 -1595
rect 1630 -1660 1750 -1625
rect 1630 -1690 1675 -1660
rect 1705 -1690 1750 -1660
rect 1630 -1720 1750 -1690
rect 1630 -1750 1675 -1720
rect 1705 -1750 1750 -1720
rect 1630 -1785 1750 -1750
rect 1630 -1815 1675 -1785
rect 1705 -1815 1750 -1785
rect 1630 -1855 1750 -1815
rect 1630 -1885 1675 -1855
rect 1705 -1885 1750 -1855
rect 1630 -1925 1750 -1885
rect 1630 -1955 1675 -1925
rect 1705 -1955 1750 -1925
rect 1630 -1995 1750 -1955
rect 1630 -2025 1675 -1995
rect 1705 -2025 1750 -1995
rect 1630 -2060 1750 -2025
rect 1630 -2090 1675 -2060
rect 1705 -2090 1750 -2060
rect 1630 -2120 1750 -2090
rect 1630 -2150 1675 -2120
rect 1705 -2150 1750 -2120
rect 1630 -2185 1750 -2150
rect 1630 -2215 1675 -2185
rect 1705 -2215 1750 -2185
rect 1630 -2255 1750 -2215
rect 1630 -2285 1675 -2255
rect 1705 -2285 1750 -2255
rect 1630 -2325 1750 -2285
rect 1630 -2355 1675 -2325
rect 1705 -2355 1750 -2325
rect 1630 -2395 1750 -2355
rect 1630 -2425 1675 -2395
rect 1705 -2425 1750 -2395
rect 1630 -2460 1750 -2425
rect 1630 -2490 1675 -2460
rect 1705 -2490 1750 -2460
rect 1630 -2520 1750 -2490
rect 1630 -2550 1675 -2520
rect 1705 -2550 1750 -2520
rect 1630 -2585 1750 -2550
rect 1630 -2615 1675 -2585
rect 1705 -2615 1750 -2585
rect 1630 -2655 1750 -2615
rect 1630 -2685 1675 -2655
rect 1705 -2685 1750 -2655
rect 1630 -2725 1750 -2685
rect 1630 -2755 1675 -2725
rect 1705 -2755 1750 -2725
rect 1630 -2795 1750 -2755
rect 1630 -2825 1675 -2795
rect 1705 -2825 1750 -2795
rect 1630 -2860 1750 -2825
rect 1630 -2890 1675 -2860
rect 1705 -2890 1750 -2860
rect 1630 -2905 1750 -2890
rect 1980 -1320 2100 -1225
rect 1980 -1350 2025 -1320
rect 2055 -1350 2100 -1320
rect 1980 -1385 2100 -1350
rect 1980 -1415 2025 -1385
rect 2055 -1415 2100 -1385
rect 1980 -1455 2100 -1415
rect 1980 -1485 2025 -1455
rect 2055 -1485 2100 -1455
rect 1980 -1525 2100 -1485
rect 1980 -1555 2025 -1525
rect 2055 -1555 2100 -1525
rect 1980 -1595 2100 -1555
rect 1980 -1625 2025 -1595
rect 2055 -1625 2100 -1595
rect 1980 -1660 2100 -1625
rect 1980 -1690 2025 -1660
rect 2055 -1690 2100 -1660
rect 1980 -1720 2100 -1690
rect 1980 -1750 2025 -1720
rect 2055 -1750 2100 -1720
rect 1980 -1785 2100 -1750
rect 1980 -1815 2025 -1785
rect 2055 -1815 2100 -1785
rect 1980 -1855 2100 -1815
rect 1980 -1885 2025 -1855
rect 2055 -1885 2100 -1855
rect 1980 -1925 2100 -1885
rect 1980 -1955 2025 -1925
rect 2055 -1955 2100 -1925
rect 1980 -1995 2100 -1955
rect 1980 -2025 2025 -1995
rect 2055 -2025 2100 -1995
rect 1980 -2060 2100 -2025
rect 1980 -2090 2025 -2060
rect 2055 -2090 2100 -2060
rect 1980 -2120 2100 -2090
rect 1980 -2150 2025 -2120
rect 2055 -2150 2100 -2120
rect 1980 -2185 2100 -2150
rect 1980 -2215 2025 -2185
rect 2055 -2215 2100 -2185
rect 1980 -2255 2100 -2215
rect 1980 -2285 2025 -2255
rect 2055 -2285 2100 -2255
rect 1980 -2325 2100 -2285
rect 1980 -2355 2025 -2325
rect 2055 -2355 2100 -2325
rect 1980 -2395 2100 -2355
rect 1980 -2425 2025 -2395
rect 2055 -2425 2100 -2395
rect 1980 -2460 2100 -2425
rect 1980 -2490 2025 -2460
rect 2055 -2490 2100 -2460
rect 1980 -2520 2100 -2490
rect 1980 -2550 2025 -2520
rect 2055 -2550 2100 -2520
rect 1980 -2585 2100 -2550
rect 1980 -2615 2025 -2585
rect 2055 -2615 2100 -2585
rect 1980 -2655 2100 -2615
rect 1980 -2685 2025 -2655
rect 2055 -2685 2100 -2655
rect 1980 -2725 2100 -2685
rect 1980 -2755 2025 -2725
rect 2055 -2755 2100 -2725
rect 1980 -2795 2100 -2755
rect 1980 -2825 2025 -2795
rect 2055 -2825 2100 -2795
rect 1980 -2860 2100 -2825
rect 1980 -2890 2025 -2860
rect 2055 -2890 2100 -2860
rect 1980 -2905 2100 -2890
rect 2330 -1320 2450 -1225
rect 2330 -1350 2375 -1320
rect 2405 -1350 2450 -1320
rect 2330 -1385 2450 -1350
rect 2330 -1415 2375 -1385
rect 2405 -1415 2450 -1385
rect 2330 -1455 2450 -1415
rect 2330 -1485 2375 -1455
rect 2405 -1485 2450 -1455
rect 2330 -1525 2450 -1485
rect 2330 -1555 2375 -1525
rect 2405 -1555 2450 -1525
rect 2330 -1595 2450 -1555
rect 2330 -1625 2375 -1595
rect 2405 -1625 2450 -1595
rect 2330 -1660 2450 -1625
rect 2330 -1690 2375 -1660
rect 2405 -1690 2450 -1660
rect 2330 -1720 2450 -1690
rect 2330 -1750 2375 -1720
rect 2405 -1750 2450 -1720
rect 2330 -1785 2450 -1750
rect 2330 -1815 2375 -1785
rect 2405 -1815 2450 -1785
rect 2330 -1855 2450 -1815
rect 2330 -1885 2375 -1855
rect 2405 -1885 2450 -1855
rect 2330 -1925 2450 -1885
rect 2330 -1955 2375 -1925
rect 2405 -1955 2450 -1925
rect 2330 -1995 2450 -1955
rect 2330 -2025 2375 -1995
rect 2405 -2025 2450 -1995
rect 2330 -2060 2450 -2025
rect 2330 -2090 2375 -2060
rect 2405 -2090 2450 -2060
rect 2330 -2120 2450 -2090
rect 2330 -2150 2375 -2120
rect 2405 -2150 2450 -2120
rect 2330 -2185 2450 -2150
rect 2330 -2215 2375 -2185
rect 2405 -2215 2450 -2185
rect 2330 -2255 2450 -2215
rect 2330 -2285 2375 -2255
rect 2405 -2285 2450 -2255
rect 2330 -2325 2450 -2285
rect 2330 -2355 2375 -2325
rect 2405 -2355 2450 -2325
rect 2330 -2395 2450 -2355
rect 2330 -2425 2375 -2395
rect 2405 -2425 2450 -2395
rect 2330 -2460 2450 -2425
rect 2330 -2490 2375 -2460
rect 2405 -2490 2450 -2460
rect 2330 -2520 2450 -2490
rect 2330 -2550 2375 -2520
rect 2405 -2550 2450 -2520
rect 2330 -2585 2450 -2550
rect 2330 -2615 2375 -2585
rect 2405 -2615 2450 -2585
rect 2330 -2655 2450 -2615
rect 2330 -2685 2375 -2655
rect 2405 -2685 2450 -2655
rect 2330 -2725 2450 -2685
rect 2330 -2755 2375 -2725
rect 2405 -2755 2450 -2725
rect 2330 -2795 2450 -2755
rect 2330 -2825 2375 -2795
rect 2405 -2825 2450 -2795
rect 2330 -2860 2450 -2825
rect 2330 -2890 2375 -2860
rect 2405 -2890 2450 -2860
rect 2330 -2905 2450 -2890
rect 2680 -1320 2800 -1225
rect 2680 -1350 2725 -1320
rect 2755 -1350 2800 -1320
rect 2680 -1385 2800 -1350
rect 2680 -1415 2725 -1385
rect 2755 -1415 2800 -1385
rect 2680 -1455 2800 -1415
rect 2680 -1485 2725 -1455
rect 2755 -1485 2800 -1455
rect 2680 -1525 2800 -1485
rect 2680 -1555 2725 -1525
rect 2755 -1555 2800 -1525
rect 2680 -1595 2800 -1555
rect 2680 -1625 2725 -1595
rect 2755 -1625 2800 -1595
rect 2680 -1660 2800 -1625
rect 2680 -1690 2725 -1660
rect 2755 -1690 2800 -1660
rect 2680 -1720 2800 -1690
rect 2680 -1750 2725 -1720
rect 2755 -1750 2800 -1720
rect 2680 -1785 2800 -1750
rect 2680 -1815 2725 -1785
rect 2755 -1815 2800 -1785
rect 2680 -1855 2800 -1815
rect 2680 -1885 2725 -1855
rect 2755 -1885 2800 -1855
rect 2680 -1925 2800 -1885
rect 2680 -1955 2725 -1925
rect 2755 -1955 2800 -1925
rect 2680 -1995 2800 -1955
rect 2680 -2025 2725 -1995
rect 2755 -2025 2800 -1995
rect 2680 -2060 2800 -2025
rect 2680 -2090 2725 -2060
rect 2755 -2090 2800 -2060
rect 2680 -2120 2800 -2090
rect 2680 -2150 2725 -2120
rect 2755 -2150 2800 -2120
rect 2680 -2185 2800 -2150
rect 2680 -2215 2725 -2185
rect 2755 -2215 2800 -2185
rect 2680 -2255 2800 -2215
rect 2680 -2285 2725 -2255
rect 2755 -2285 2800 -2255
rect 2680 -2325 2800 -2285
rect 2680 -2355 2725 -2325
rect 2755 -2355 2800 -2325
rect 2680 -2395 2800 -2355
rect 2680 -2425 2725 -2395
rect 2755 -2425 2800 -2395
rect 2680 -2460 2800 -2425
rect 2680 -2490 2725 -2460
rect 2755 -2490 2800 -2460
rect 2680 -2520 2800 -2490
rect 2680 -2550 2725 -2520
rect 2755 -2550 2800 -2520
rect 2680 -2585 2800 -2550
rect 2680 -2615 2725 -2585
rect 2755 -2615 2800 -2585
rect 2680 -2655 2800 -2615
rect 2680 -2685 2725 -2655
rect 2755 -2685 2800 -2655
rect 2680 -2725 2800 -2685
rect 2680 -2755 2725 -2725
rect 2755 -2755 2800 -2725
rect 2680 -2795 2800 -2755
rect 2680 -2825 2725 -2795
rect 2755 -2825 2800 -2795
rect 2680 -2860 2800 -2825
rect 2680 -2890 2725 -2860
rect 2755 -2890 2800 -2860
rect 2680 -2905 2800 -2890
rect 3030 -1320 3150 -1225
rect 3030 -1350 3075 -1320
rect 3105 -1350 3150 -1320
rect 3030 -1385 3150 -1350
rect 3030 -1415 3075 -1385
rect 3105 -1415 3150 -1385
rect 3030 -1455 3150 -1415
rect 3030 -1485 3075 -1455
rect 3105 -1485 3150 -1455
rect 3030 -1525 3150 -1485
rect 3030 -1555 3075 -1525
rect 3105 -1555 3150 -1525
rect 3030 -1595 3150 -1555
rect 3030 -1625 3075 -1595
rect 3105 -1625 3150 -1595
rect 3030 -1660 3150 -1625
rect 3030 -1690 3075 -1660
rect 3105 -1690 3150 -1660
rect 3030 -1720 3150 -1690
rect 3030 -1750 3075 -1720
rect 3105 -1750 3150 -1720
rect 3030 -1785 3150 -1750
rect 3030 -1815 3075 -1785
rect 3105 -1815 3150 -1785
rect 3030 -1855 3150 -1815
rect 3030 -1885 3075 -1855
rect 3105 -1885 3150 -1855
rect 3030 -1925 3150 -1885
rect 3030 -1955 3075 -1925
rect 3105 -1955 3150 -1925
rect 3030 -1995 3150 -1955
rect 3030 -2025 3075 -1995
rect 3105 -2025 3150 -1995
rect 3030 -2060 3150 -2025
rect 3030 -2090 3075 -2060
rect 3105 -2090 3150 -2060
rect 3030 -2120 3150 -2090
rect 3030 -2150 3075 -2120
rect 3105 -2150 3150 -2120
rect 3030 -2185 3150 -2150
rect 3030 -2215 3075 -2185
rect 3105 -2215 3150 -2185
rect 3030 -2255 3150 -2215
rect 3030 -2285 3075 -2255
rect 3105 -2285 3150 -2255
rect 3030 -2325 3150 -2285
rect 3030 -2355 3075 -2325
rect 3105 -2355 3150 -2325
rect 3030 -2395 3150 -2355
rect 3030 -2425 3075 -2395
rect 3105 -2425 3150 -2395
rect 3030 -2460 3150 -2425
rect 3030 -2490 3075 -2460
rect 3105 -2490 3150 -2460
rect 3030 -2520 3150 -2490
rect 3030 -2550 3075 -2520
rect 3105 -2550 3150 -2520
rect 3030 -2585 3150 -2550
rect 3030 -2615 3075 -2585
rect 3105 -2615 3150 -2585
rect 3030 -2655 3150 -2615
rect 3030 -2685 3075 -2655
rect 3105 -2685 3150 -2655
rect 3030 -2725 3150 -2685
rect 3030 -2755 3075 -2725
rect 3105 -2755 3150 -2725
rect 3030 -2795 3150 -2755
rect 3030 -2825 3075 -2795
rect 3105 -2825 3150 -2795
rect 3030 -2860 3150 -2825
rect 3030 -2890 3075 -2860
rect 3105 -2890 3150 -2860
rect 3030 -2905 3150 -2890
rect 3380 -3020 3500 -1250
rect 3380 -3050 3425 -3020
rect 3455 -3050 3500 -3020
rect 3380 -3085 3500 -3050
rect 3380 -3115 3425 -3085
rect 3455 -3115 3500 -3085
rect 3380 -3155 3500 -3115
rect 3380 -3185 3425 -3155
rect 3455 -3185 3500 -3155
rect 3380 -3225 3500 -3185
rect 3380 -3255 3425 -3225
rect 3455 -3255 3500 -3225
rect 3380 -3295 3500 -3255
rect 3380 -3325 3425 -3295
rect 3455 -3325 3500 -3295
rect 3380 -3360 3500 -3325
rect 3380 -3390 3425 -3360
rect 3455 -3390 3500 -3360
rect 3380 -3420 3500 -3390
rect 3380 -3450 3425 -3420
rect 3455 -3450 3500 -3420
rect 3380 -3485 3500 -3450
rect 3380 -3515 3425 -3485
rect 3455 -3515 3500 -3485
rect 3380 -3555 3500 -3515
rect 3380 -3585 3425 -3555
rect 3455 -3585 3500 -3555
rect 3380 -3625 3500 -3585
rect 3380 -3655 3425 -3625
rect 3455 -3655 3500 -3625
rect 3380 -3695 3500 -3655
rect 3380 -3725 3425 -3695
rect 3455 -3725 3500 -3695
rect 3380 -3760 3500 -3725
rect 3380 -3790 3425 -3760
rect 3455 -3790 3500 -3760
rect 3380 -3820 3500 -3790
rect 3380 -3850 3425 -3820
rect 3455 -3850 3500 -3820
rect 3380 -3885 3500 -3850
rect 3380 -3915 3425 -3885
rect 3455 -3915 3500 -3885
rect 3380 -3955 3500 -3915
rect 3380 -3985 3425 -3955
rect 3455 -3985 3500 -3955
rect 3380 -4025 3500 -3985
rect 3380 -4055 3425 -4025
rect 3455 -4055 3500 -4025
rect 3380 -4095 3500 -4055
rect 3380 -4125 3425 -4095
rect 3455 -4125 3500 -4095
rect 3380 -4160 3500 -4125
rect 3380 -4190 3425 -4160
rect 3455 -4190 3500 -4160
rect 3380 -4220 3500 -4190
rect 3380 -4250 3425 -4220
rect 3455 -4250 3500 -4220
rect 3380 -4285 3500 -4250
rect 3380 -4315 3425 -4285
rect 3455 -4315 3500 -4285
rect 3380 -4355 3500 -4315
rect 3380 -4385 3425 -4355
rect 3455 -4385 3500 -4355
rect 3380 -4425 3500 -4385
rect 3380 -4455 3425 -4425
rect 3455 -4455 3500 -4425
rect 3380 -4495 3500 -4455
rect 3380 -4525 3425 -4495
rect 3455 -4525 3500 -4495
rect 3380 -4560 3500 -4525
rect 3380 -4590 3425 -4560
rect 3455 -4590 3500 -4560
rect 3380 -4605 3500 -4590
rect 3730 -3020 3850 -1250
rect 3730 -3050 3775 -3020
rect 3805 -3050 3850 -3020
rect 3730 -3085 3850 -3050
rect 3730 -3115 3775 -3085
rect 3805 -3115 3850 -3085
rect 3730 -3155 3850 -3115
rect 3730 -3185 3775 -3155
rect 3805 -3185 3850 -3155
rect 3730 -3225 3850 -3185
rect 3730 -3255 3775 -3225
rect 3805 -3255 3850 -3225
rect 3730 -3295 3850 -3255
rect 3730 -3325 3775 -3295
rect 3805 -3325 3850 -3295
rect 3730 -3360 3850 -3325
rect 3730 -3390 3775 -3360
rect 3805 -3390 3850 -3360
rect 3730 -3420 3850 -3390
rect 3730 -3450 3775 -3420
rect 3805 -3450 3850 -3420
rect 3730 -3485 3850 -3450
rect 3730 -3515 3775 -3485
rect 3805 -3515 3850 -3485
rect 3730 -3555 3850 -3515
rect 3730 -3585 3775 -3555
rect 3805 -3585 3850 -3555
rect 3730 -3625 3850 -3585
rect 3730 -3655 3775 -3625
rect 3805 -3655 3850 -3625
rect 3730 -3695 3850 -3655
rect 3730 -3725 3775 -3695
rect 3805 -3725 3850 -3695
rect 3730 -3760 3850 -3725
rect 3730 -3790 3775 -3760
rect 3805 -3790 3850 -3760
rect 3730 -3820 3850 -3790
rect 3730 -3850 3775 -3820
rect 3805 -3850 3850 -3820
rect 3730 -3885 3850 -3850
rect 3730 -3915 3775 -3885
rect 3805 -3915 3850 -3885
rect 3730 -3955 3850 -3915
rect 3730 -3985 3775 -3955
rect 3805 -3985 3850 -3955
rect 3730 -4025 3850 -3985
rect 3730 -4055 3775 -4025
rect 3805 -4055 3850 -4025
rect 3730 -4095 3850 -4055
rect 3730 -4125 3775 -4095
rect 3805 -4125 3850 -4095
rect 3730 -4160 3850 -4125
rect 3730 -4190 3775 -4160
rect 3805 -4190 3850 -4160
rect 3730 -4220 3850 -4190
rect 3730 -4250 3775 -4220
rect 3805 -4250 3850 -4220
rect 3730 -4285 3850 -4250
rect 3730 -4315 3775 -4285
rect 3805 -4315 3850 -4285
rect 3730 -4355 3850 -4315
rect 3730 -4385 3775 -4355
rect 3805 -4385 3850 -4355
rect 3730 -4425 3850 -4385
rect 3730 -4455 3775 -4425
rect 3805 -4455 3850 -4425
rect 3730 -4495 3850 -4455
rect 3730 -4525 3775 -4495
rect 3805 -4525 3850 -4495
rect 3730 -4560 3850 -4525
rect 3730 -4590 3775 -4560
rect 3805 -4590 3850 -4560
rect 3730 -4605 3850 -4590
rect 4080 -3020 4200 -1250
rect 4080 -3050 4125 -3020
rect 4155 -3050 4200 -3020
rect 4080 -3085 4200 -3050
rect 4080 -3115 4125 -3085
rect 4155 -3115 4200 -3085
rect 4080 -3155 4200 -3115
rect 4080 -3185 4125 -3155
rect 4155 -3185 4200 -3155
rect 4080 -3225 4200 -3185
rect 4080 -3255 4125 -3225
rect 4155 -3255 4200 -3225
rect 4080 -3295 4200 -3255
rect 4080 -3325 4125 -3295
rect 4155 -3325 4200 -3295
rect 4080 -3360 4200 -3325
rect 4080 -3390 4125 -3360
rect 4155 -3390 4200 -3360
rect 4080 -3420 4200 -3390
rect 4080 -3450 4125 -3420
rect 4155 -3450 4200 -3420
rect 4080 -3485 4200 -3450
rect 4080 -3515 4125 -3485
rect 4155 -3515 4200 -3485
rect 4080 -3555 4200 -3515
rect 4080 -3585 4125 -3555
rect 4155 -3585 4200 -3555
rect 4080 -3625 4200 -3585
rect 4080 -3655 4125 -3625
rect 4155 -3655 4200 -3625
rect 4080 -3695 4200 -3655
rect 4080 -3725 4125 -3695
rect 4155 -3725 4200 -3695
rect 4080 -3760 4200 -3725
rect 4080 -3790 4125 -3760
rect 4155 -3790 4200 -3760
rect 4080 -3820 4200 -3790
rect 4080 -3850 4125 -3820
rect 4155 -3850 4200 -3820
rect 4080 -3885 4200 -3850
rect 4080 -3915 4125 -3885
rect 4155 -3915 4200 -3885
rect 4080 -3955 4200 -3915
rect 4080 -3985 4125 -3955
rect 4155 -3985 4200 -3955
rect 4080 -4025 4200 -3985
rect 4080 -4055 4125 -4025
rect 4155 -4055 4200 -4025
rect 4080 -4095 4200 -4055
rect 4080 -4125 4125 -4095
rect 4155 -4125 4200 -4095
rect 4080 -4160 4200 -4125
rect 4080 -4190 4125 -4160
rect 4155 -4190 4200 -4160
rect 4080 -4220 4200 -4190
rect 4080 -4250 4125 -4220
rect 4155 -4250 4200 -4220
rect 4080 -4285 4200 -4250
rect 4080 -4315 4125 -4285
rect 4155 -4315 4200 -4285
rect 4080 -4355 4200 -4315
rect 4080 -4385 4125 -4355
rect 4155 -4385 4200 -4355
rect 4080 -4425 4200 -4385
rect 4080 -4455 4125 -4425
rect 4155 -4455 4200 -4425
rect 4080 -4495 4200 -4455
rect 4080 -4525 4125 -4495
rect 4155 -4525 4200 -4495
rect 4080 -4560 4200 -4525
rect 4080 -4590 4125 -4560
rect 4155 -4590 4200 -4560
rect 4080 -4605 4200 -4590
rect 4430 -3020 4550 -1250
rect 4430 -3050 4475 -3020
rect 4505 -3050 4550 -3020
rect 4430 -3085 4550 -3050
rect 4430 -3115 4475 -3085
rect 4505 -3115 4550 -3085
rect 4430 -3155 4550 -3115
rect 4430 -3185 4475 -3155
rect 4505 -3185 4550 -3155
rect 4430 -3225 4550 -3185
rect 4430 -3255 4475 -3225
rect 4505 -3255 4550 -3225
rect 4430 -3295 4550 -3255
rect 4430 -3325 4475 -3295
rect 4505 -3325 4550 -3295
rect 4430 -3360 4550 -3325
rect 4430 -3390 4475 -3360
rect 4505 -3390 4550 -3360
rect 4430 -3420 4550 -3390
rect 4430 -3450 4475 -3420
rect 4505 -3450 4550 -3420
rect 4430 -3485 4550 -3450
rect 4430 -3515 4475 -3485
rect 4505 -3515 4550 -3485
rect 4430 -3555 4550 -3515
rect 4430 -3585 4475 -3555
rect 4505 -3585 4550 -3555
rect 4430 -3625 4550 -3585
rect 4430 -3655 4475 -3625
rect 4505 -3655 4550 -3625
rect 4430 -3695 4550 -3655
rect 4430 -3725 4475 -3695
rect 4505 -3725 4550 -3695
rect 4430 -3760 4550 -3725
rect 4430 -3790 4475 -3760
rect 4505 -3790 4550 -3760
rect 4430 -3820 4550 -3790
rect 4430 -3850 4475 -3820
rect 4505 -3850 4550 -3820
rect 4430 -3885 4550 -3850
rect 4430 -3915 4475 -3885
rect 4505 -3915 4550 -3885
rect 4430 -3955 4550 -3915
rect 4430 -3985 4475 -3955
rect 4505 -3985 4550 -3955
rect 4430 -4025 4550 -3985
rect 4430 -4055 4475 -4025
rect 4505 -4055 4550 -4025
rect 4430 -4095 4550 -4055
rect 4430 -4125 4475 -4095
rect 4505 -4125 4550 -4095
rect 4430 -4160 4550 -4125
rect 4430 -4190 4475 -4160
rect 4505 -4190 4550 -4160
rect 4430 -4220 4550 -4190
rect 4430 -4250 4475 -4220
rect 4505 -4250 4550 -4220
rect 4430 -4285 4550 -4250
rect 4430 -4315 4475 -4285
rect 4505 -4315 4550 -4285
rect 4430 -4355 4550 -4315
rect 4430 -4385 4475 -4355
rect 4505 -4385 4550 -4355
rect 4430 -4425 4550 -4385
rect 4430 -4455 4475 -4425
rect 4505 -4455 4550 -4425
rect 4430 -4495 4550 -4455
rect 4430 -4525 4475 -4495
rect 4505 -4525 4550 -4495
rect 4430 -4560 4550 -4525
rect 4430 -4590 4475 -4560
rect 4505 -4590 4550 -4560
rect 4430 -4605 4550 -4590
rect 4780 -3020 4900 -1250
rect 4780 -3050 4825 -3020
rect 4855 -3050 4900 -3020
rect 4780 -3085 4900 -3050
rect 4780 -3115 4825 -3085
rect 4855 -3115 4900 -3085
rect 4780 -3155 4900 -3115
rect 4780 -3185 4825 -3155
rect 4855 -3185 4900 -3155
rect 4780 -3225 4900 -3185
rect 4780 -3255 4825 -3225
rect 4855 -3255 4900 -3225
rect 4780 -3295 4900 -3255
rect 4780 -3325 4825 -3295
rect 4855 -3325 4900 -3295
rect 4780 -3360 4900 -3325
rect 4780 -3390 4825 -3360
rect 4855 -3390 4900 -3360
rect 4780 -3420 4900 -3390
rect 4780 -3450 4825 -3420
rect 4855 -3450 4900 -3420
rect 4780 -3485 4900 -3450
rect 4780 -3515 4825 -3485
rect 4855 -3515 4900 -3485
rect 4780 -3555 4900 -3515
rect 4780 -3585 4825 -3555
rect 4855 -3585 4900 -3555
rect 4780 -3625 4900 -3585
rect 4780 -3655 4825 -3625
rect 4855 -3655 4900 -3625
rect 4780 -3695 4900 -3655
rect 4780 -3725 4825 -3695
rect 4855 -3725 4900 -3695
rect 4780 -3760 4900 -3725
rect 4780 -3790 4825 -3760
rect 4855 -3790 4900 -3760
rect 4780 -3820 4900 -3790
rect 4780 -3850 4825 -3820
rect 4855 -3850 4900 -3820
rect 4780 -3885 4900 -3850
rect 4780 -3915 4825 -3885
rect 4855 -3915 4900 -3885
rect 4780 -3955 4900 -3915
rect 4780 -3985 4825 -3955
rect 4855 -3985 4900 -3955
rect 4780 -4025 4900 -3985
rect 4780 -4055 4825 -4025
rect 4855 -4055 4900 -4025
rect 4780 -4095 4900 -4055
rect 4780 -4125 4825 -4095
rect 4855 -4125 4900 -4095
rect 4780 -4160 4900 -4125
rect 4780 -4190 4825 -4160
rect 4855 -4190 4900 -4160
rect 4780 -4220 4900 -4190
rect 4780 -4250 4825 -4220
rect 4855 -4250 4900 -4220
rect 4780 -4285 4900 -4250
rect 4780 -4315 4825 -4285
rect 4855 -4315 4900 -4285
rect 4780 -4355 4900 -4315
rect 4780 -4385 4825 -4355
rect 4855 -4385 4900 -4355
rect 4780 -4425 4900 -4385
rect 4780 -4455 4825 -4425
rect 4855 -4455 4900 -4425
rect 4780 -4495 4900 -4455
rect 4780 -4525 4825 -4495
rect 4855 -4525 4900 -4495
rect 4780 -4560 4900 -4525
rect 4780 -4590 4825 -4560
rect 4855 -4590 4900 -4560
rect 4780 -4605 4900 -4590
rect 5130 -3020 5250 -1250
rect 5130 -3050 5175 -3020
rect 5205 -3050 5250 -3020
rect 5130 -3085 5250 -3050
rect 5130 -3115 5175 -3085
rect 5205 -3115 5250 -3085
rect 5130 -3155 5250 -3115
rect 5130 -3185 5175 -3155
rect 5205 -3185 5250 -3155
rect 5130 -3225 5250 -3185
rect 5130 -3255 5175 -3225
rect 5205 -3255 5250 -3225
rect 5130 -3295 5250 -3255
rect 5130 -3325 5175 -3295
rect 5205 -3325 5250 -3295
rect 5130 -3360 5250 -3325
rect 5130 -3390 5175 -3360
rect 5205 -3390 5250 -3360
rect 5130 -3420 5250 -3390
rect 5130 -3450 5175 -3420
rect 5205 -3450 5250 -3420
rect 5130 -3485 5250 -3450
rect 5130 -3515 5175 -3485
rect 5205 -3515 5250 -3485
rect 5130 -3555 5250 -3515
rect 5130 -3585 5175 -3555
rect 5205 -3585 5250 -3555
rect 5130 -3625 5250 -3585
rect 5130 -3655 5175 -3625
rect 5205 -3655 5250 -3625
rect 5130 -3695 5250 -3655
rect 5130 -3725 5175 -3695
rect 5205 -3725 5250 -3695
rect 5130 -3760 5250 -3725
rect 5130 -3790 5175 -3760
rect 5205 -3790 5250 -3760
rect 5130 -3820 5250 -3790
rect 5130 -3850 5175 -3820
rect 5205 -3850 5250 -3820
rect 5130 -3885 5250 -3850
rect 5130 -3915 5175 -3885
rect 5205 -3915 5250 -3885
rect 5130 -3955 5250 -3915
rect 5130 -3985 5175 -3955
rect 5205 -3985 5250 -3955
rect 5130 -4025 5250 -3985
rect 5130 -4055 5175 -4025
rect 5205 -4055 5250 -4025
rect 5130 -4095 5250 -4055
rect 5130 -4125 5175 -4095
rect 5205 -4125 5250 -4095
rect 5130 -4160 5250 -4125
rect 5130 -4190 5175 -4160
rect 5205 -4190 5250 -4160
rect 5130 -4220 5250 -4190
rect 5130 -4250 5175 -4220
rect 5205 -4250 5250 -4220
rect 5130 -4285 5250 -4250
rect 5130 -4315 5175 -4285
rect 5205 -4315 5250 -4285
rect 5130 -4355 5250 -4315
rect 5130 -4385 5175 -4355
rect 5205 -4385 5250 -4355
rect 5130 -4425 5250 -4385
rect 5130 -4455 5175 -4425
rect 5205 -4455 5250 -4425
rect 5130 -4495 5250 -4455
rect 5130 -4525 5175 -4495
rect 5205 -4525 5250 -4495
rect 5130 -4560 5250 -4525
rect 5130 -4590 5175 -4560
rect 5205 -4590 5250 -4560
rect 5130 -4605 5250 -4590
rect 5480 -3020 5600 -1250
rect 5830 -1320 5950 -1225
rect 5830 -1350 5875 -1320
rect 5905 -1350 5950 -1320
rect 5830 -1385 5950 -1350
rect 5830 -1415 5875 -1385
rect 5905 -1415 5950 -1385
rect 5830 -1455 5950 -1415
rect 5830 -1485 5875 -1455
rect 5905 -1485 5950 -1455
rect 5830 -1525 5950 -1485
rect 5830 -1555 5875 -1525
rect 5905 -1555 5950 -1525
rect 5830 -1595 5950 -1555
rect 5830 -1625 5875 -1595
rect 5905 -1625 5950 -1595
rect 5830 -1660 5950 -1625
rect 5830 -1690 5875 -1660
rect 5905 -1690 5950 -1660
rect 5830 -1720 5950 -1690
rect 5830 -1750 5875 -1720
rect 5905 -1750 5950 -1720
rect 5830 -1785 5950 -1750
rect 5830 -1815 5875 -1785
rect 5905 -1815 5950 -1785
rect 5830 -1855 5950 -1815
rect 5830 -1885 5875 -1855
rect 5905 -1885 5950 -1855
rect 5830 -1925 5950 -1885
rect 5830 -1955 5875 -1925
rect 5905 -1955 5950 -1925
rect 5830 -1995 5950 -1955
rect 5830 -2025 5875 -1995
rect 5905 -2025 5950 -1995
rect 5830 -2060 5950 -2025
rect 5830 -2090 5875 -2060
rect 5905 -2090 5950 -2060
rect 5830 -2120 5950 -2090
rect 5830 -2150 5875 -2120
rect 5905 -2150 5950 -2120
rect 5830 -2185 5950 -2150
rect 5830 -2215 5875 -2185
rect 5905 -2215 5950 -2185
rect 5830 -2255 5950 -2215
rect 5830 -2285 5875 -2255
rect 5905 -2285 5950 -2255
rect 5830 -2325 5950 -2285
rect 5830 -2355 5875 -2325
rect 5905 -2355 5950 -2325
rect 5830 -2395 5950 -2355
rect 5830 -2425 5875 -2395
rect 5905 -2425 5950 -2395
rect 5830 -2460 5950 -2425
rect 5830 -2490 5875 -2460
rect 5905 -2490 5950 -2460
rect 5830 -2520 5950 -2490
rect 5830 -2550 5875 -2520
rect 5905 -2550 5950 -2520
rect 5830 -2585 5950 -2550
rect 5830 -2615 5875 -2585
rect 5905 -2615 5950 -2585
rect 5830 -2655 5950 -2615
rect 5830 -2685 5875 -2655
rect 5905 -2685 5950 -2655
rect 5830 -2725 5950 -2685
rect 5830 -2755 5875 -2725
rect 5905 -2755 5950 -2725
rect 5830 -2795 5950 -2755
rect 5830 -2825 5875 -2795
rect 5905 -2825 5950 -2795
rect 5830 -2860 5950 -2825
rect 5830 -2890 5875 -2860
rect 5905 -2890 5950 -2860
rect 5830 -2905 5950 -2890
rect 6180 -1320 6300 -1225
rect 6180 -1350 6225 -1320
rect 6255 -1350 6300 -1320
rect 6180 -1385 6300 -1350
rect 6180 -1415 6225 -1385
rect 6255 -1415 6300 -1385
rect 6180 -1455 6300 -1415
rect 6180 -1485 6225 -1455
rect 6255 -1485 6300 -1455
rect 6180 -1525 6300 -1485
rect 6180 -1555 6225 -1525
rect 6255 -1555 6300 -1525
rect 6180 -1595 6300 -1555
rect 6180 -1625 6225 -1595
rect 6255 -1625 6300 -1595
rect 6180 -1660 6300 -1625
rect 6180 -1690 6225 -1660
rect 6255 -1690 6300 -1660
rect 6180 -1720 6300 -1690
rect 6180 -1750 6225 -1720
rect 6255 -1750 6300 -1720
rect 6180 -1785 6300 -1750
rect 6180 -1815 6225 -1785
rect 6255 -1815 6300 -1785
rect 6180 -1855 6300 -1815
rect 6180 -1885 6225 -1855
rect 6255 -1885 6300 -1855
rect 6180 -1925 6300 -1885
rect 6180 -1955 6225 -1925
rect 6255 -1955 6300 -1925
rect 6180 -1995 6300 -1955
rect 6180 -2025 6225 -1995
rect 6255 -2025 6300 -1995
rect 6180 -2060 6300 -2025
rect 6180 -2090 6225 -2060
rect 6255 -2090 6300 -2060
rect 6180 -2120 6300 -2090
rect 6180 -2150 6225 -2120
rect 6255 -2150 6300 -2120
rect 6180 -2185 6300 -2150
rect 6180 -2215 6225 -2185
rect 6255 -2215 6300 -2185
rect 6180 -2255 6300 -2215
rect 6180 -2285 6225 -2255
rect 6255 -2285 6300 -2255
rect 6180 -2325 6300 -2285
rect 6180 -2355 6225 -2325
rect 6255 -2355 6300 -2325
rect 6180 -2395 6300 -2355
rect 6180 -2425 6225 -2395
rect 6255 -2425 6300 -2395
rect 6180 -2460 6300 -2425
rect 6180 -2490 6225 -2460
rect 6255 -2490 6300 -2460
rect 6180 -2520 6300 -2490
rect 6180 -2550 6225 -2520
rect 6255 -2550 6300 -2520
rect 6180 -2585 6300 -2550
rect 6180 -2615 6225 -2585
rect 6255 -2615 6300 -2585
rect 6180 -2655 6300 -2615
rect 6180 -2685 6225 -2655
rect 6255 -2685 6300 -2655
rect 6180 -2725 6300 -2685
rect 6180 -2755 6225 -2725
rect 6255 -2755 6300 -2725
rect 6180 -2795 6300 -2755
rect 6180 -2825 6225 -2795
rect 6255 -2825 6300 -2795
rect 6180 -2860 6300 -2825
rect 6180 -2890 6225 -2860
rect 6255 -2890 6300 -2860
rect 6180 -2905 6300 -2890
rect 6530 -1320 6650 -1225
rect 6530 -1350 6575 -1320
rect 6605 -1350 6650 -1320
rect 6530 -1385 6650 -1350
rect 6530 -1415 6575 -1385
rect 6605 -1415 6650 -1385
rect 6530 -1455 6650 -1415
rect 6530 -1485 6575 -1455
rect 6605 -1485 6650 -1455
rect 6530 -1525 6650 -1485
rect 6530 -1555 6575 -1525
rect 6605 -1555 6650 -1525
rect 6530 -1595 6650 -1555
rect 6530 -1625 6575 -1595
rect 6605 -1625 6650 -1595
rect 6530 -1660 6650 -1625
rect 6530 -1690 6575 -1660
rect 6605 -1690 6650 -1660
rect 6530 -1720 6650 -1690
rect 6530 -1750 6575 -1720
rect 6605 -1750 6650 -1720
rect 6530 -1785 6650 -1750
rect 6530 -1815 6575 -1785
rect 6605 -1815 6650 -1785
rect 6530 -1855 6650 -1815
rect 6530 -1885 6575 -1855
rect 6605 -1885 6650 -1855
rect 6530 -1925 6650 -1885
rect 6530 -1955 6575 -1925
rect 6605 -1955 6650 -1925
rect 6530 -1995 6650 -1955
rect 6530 -2025 6575 -1995
rect 6605 -2025 6650 -1995
rect 6530 -2060 6650 -2025
rect 6530 -2090 6575 -2060
rect 6605 -2090 6650 -2060
rect 6530 -2120 6650 -2090
rect 6530 -2150 6575 -2120
rect 6605 -2150 6650 -2120
rect 6530 -2185 6650 -2150
rect 6530 -2215 6575 -2185
rect 6605 -2215 6650 -2185
rect 6530 -2255 6650 -2215
rect 6530 -2285 6575 -2255
rect 6605 -2285 6650 -2255
rect 6530 -2325 6650 -2285
rect 6530 -2355 6575 -2325
rect 6605 -2355 6650 -2325
rect 6530 -2395 6650 -2355
rect 6530 -2425 6575 -2395
rect 6605 -2425 6650 -2395
rect 6530 -2460 6650 -2425
rect 6530 -2490 6575 -2460
rect 6605 -2490 6650 -2460
rect 6530 -2520 6650 -2490
rect 6530 -2550 6575 -2520
rect 6605 -2550 6650 -2520
rect 6530 -2585 6650 -2550
rect 6530 -2615 6575 -2585
rect 6605 -2615 6650 -2585
rect 6530 -2655 6650 -2615
rect 6530 -2685 6575 -2655
rect 6605 -2685 6650 -2655
rect 6530 -2725 6650 -2685
rect 6530 -2755 6575 -2725
rect 6605 -2755 6650 -2725
rect 6530 -2795 6650 -2755
rect 6530 -2825 6575 -2795
rect 6605 -2825 6650 -2795
rect 6530 -2860 6650 -2825
rect 6530 -2890 6575 -2860
rect 6605 -2890 6650 -2860
rect 6530 -2905 6650 -2890
rect 6880 -1320 7000 -1225
rect 6880 -1350 6925 -1320
rect 6955 -1350 7000 -1320
rect 6880 -1385 7000 -1350
rect 6880 -1415 6925 -1385
rect 6955 -1415 7000 -1385
rect 6880 -1455 7000 -1415
rect 6880 -1485 6925 -1455
rect 6955 -1485 7000 -1455
rect 6880 -1525 7000 -1485
rect 6880 -1555 6925 -1525
rect 6955 -1555 7000 -1525
rect 6880 -1595 7000 -1555
rect 6880 -1625 6925 -1595
rect 6955 -1625 7000 -1595
rect 6880 -1660 7000 -1625
rect 6880 -1690 6925 -1660
rect 6955 -1690 7000 -1660
rect 6880 -1720 7000 -1690
rect 6880 -1750 6925 -1720
rect 6955 -1750 7000 -1720
rect 6880 -1785 7000 -1750
rect 6880 -1815 6925 -1785
rect 6955 -1815 7000 -1785
rect 6880 -1855 7000 -1815
rect 6880 -1885 6925 -1855
rect 6955 -1885 7000 -1855
rect 6880 -1925 7000 -1885
rect 6880 -1955 6925 -1925
rect 6955 -1955 7000 -1925
rect 6880 -1995 7000 -1955
rect 6880 -2025 6925 -1995
rect 6955 -2025 7000 -1995
rect 6880 -2060 7000 -2025
rect 6880 -2090 6925 -2060
rect 6955 -2090 7000 -2060
rect 6880 -2120 7000 -2090
rect 6880 -2150 6925 -2120
rect 6955 -2150 7000 -2120
rect 6880 -2185 7000 -2150
rect 6880 -2215 6925 -2185
rect 6955 -2215 7000 -2185
rect 6880 -2255 7000 -2215
rect 6880 -2285 6925 -2255
rect 6955 -2285 7000 -2255
rect 6880 -2325 7000 -2285
rect 6880 -2355 6925 -2325
rect 6955 -2355 7000 -2325
rect 6880 -2395 7000 -2355
rect 6880 -2425 6925 -2395
rect 6955 -2425 7000 -2395
rect 6880 -2460 7000 -2425
rect 6880 -2490 6925 -2460
rect 6955 -2490 7000 -2460
rect 6880 -2520 7000 -2490
rect 6880 -2550 6925 -2520
rect 6955 -2550 7000 -2520
rect 6880 -2585 7000 -2550
rect 6880 -2615 6925 -2585
rect 6955 -2615 7000 -2585
rect 6880 -2655 7000 -2615
rect 6880 -2685 6925 -2655
rect 6955 -2685 7000 -2655
rect 6880 -2725 7000 -2685
rect 6880 -2755 6925 -2725
rect 6955 -2755 7000 -2725
rect 6880 -2795 7000 -2755
rect 6880 -2825 6925 -2795
rect 6955 -2825 7000 -2795
rect 6880 -2860 7000 -2825
rect 6880 -2890 6925 -2860
rect 6955 -2890 7000 -2860
rect 6880 -2905 7000 -2890
rect 7230 -1320 7350 -1225
rect 7230 -1350 7275 -1320
rect 7305 -1350 7350 -1320
rect 7230 -1385 7350 -1350
rect 7230 -1415 7275 -1385
rect 7305 -1415 7350 -1385
rect 7230 -1455 7350 -1415
rect 7230 -1485 7275 -1455
rect 7305 -1485 7350 -1455
rect 7230 -1525 7350 -1485
rect 7230 -1555 7275 -1525
rect 7305 -1555 7350 -1525
rect 7230 -1595 7350 -1555
rect 7230 -1625 7275 -1595
rect 7305 -1625 7350 -1595
rect 7230 -1660 7350 -1625
rect 7230 -1690 7275 -1660
rect 7305 -1690 7350 -1660
rect 7230 -1720 7350 -1690
rect 7230 -1750 7275 -1720
rect 7305 -1750 7350 -1720
rect 7230 -1785 7350 -1750
rect 7230 -1815 7275 -1785
rect 7305 -1815 7350 -1785
rect 7230 -1855 7350 -1815
rect 7230 -1885 7275 -1855
rect 7305 -1885 7350 -1855
rect 7230 -1925 7350 -1885
rect 7230 -1955 7275 -1925
rect 7305 -1955 7350 -1925
rect 7230 -1995 7350 -1955
rect 7230 -2025 7275 -1995
rect 7305 -2025 7350 -1995
rect 7230 -2060 7350 -2025
rect 7230 -2090 7275 -2060
rect 7305 -2090 7350 -2060
rect 7230 -2120 7350 -2090
rect 7230 -2150 7275 -2120
rect 7305 -2150 7350 -2120
rect 7230 -2185 7350 -2150
rect 7230 -2215 7275 -2185
rect 7305 -2215 7350 -2185
rect 7230 -2255 7350 -2215
rect 7230 -2285 7275 -2255
rect 7305 -2285 7350 -2255
rect 7230 -2325 7350 -2285
rect 7230 -2355 7275 -2325
rect 7305 -2355 7350 -2325
rect 7230 -2395 7350 -2355
rect 7230 -2425 7275 -2395
rect 7305 -2425 7350 -2395
rect 7230 -2460 7350 -2425
rect 7230 -2490 7275 -2460
rect 7305 -2490 7350 -2460
rect 7230 -2520 7350 -2490
rect 7230 -2550 7275 -2520
rect 7305 -2550 7350 -2520
rect 7230 -2585 7350 -2550
rect 7230 -2615 7275 -2585
rect 7305 -2615 7350 -2585
rect 7230 -2655 7350 -2615
rect 7230 -2685 7275 -2655
rect 7305 -2685 7350 -2655
rect 7230 -2725 7350 -2685
rect 7230 -2755 7275 -2725
rect 7305 -2755 7350 -2725
rect 7230 -2795 7350 -2755
rect 7230 -2825 7275 -2795
rect 7305 -2825 7350 -2795
rect 7230 -2860 7350 -2825
rect 7230 -2890 7275 -2860
rect 7305 -2890 7350 -2860
rect 7230 -2905 7350 -2890
rect 7580 -1320 7700 -1225
rect 7580 -1350 7625 -1320
rect 7655 -1350 7700 -1320
rect 7580 -1385 7700 -1350
rect 7580 -1415 7625 -1385
rect 7655 -1415 7700 -1385
rect 7580 -1455 7700 -1415
rect 7580 -1485 7625 -1455
rect 7655 -1485 7700 -1455
rect 7580 -1525 7700 -1485
rect 7580 -1555 7625 -1525
rect 7655 -1555 7700 -1525
rect 7580 -1595 7700 -1555
rect 7580 -1625 7625 -1595
rect 7655 -1625 7700 -1595
rect 7580 -1660 7700 -1625
rect 7580 -1690 7625 -1660
rect 7655 -1690 7700 -1660
rect 7580 -1720 7700 -1690
rect 7580 -1750 7625 -1720
rect 7655 -1750 7700 -1720
rect 7580 -1785 7700 -1750
rect 7580 -1815 7625 -1785
rect 7655 -1815 7700 -1785
rect 7580 -1855 7700 -1815
rect 7580 -1885 7625 -1855
rect 7655 -1885 7700 -1855
rect 7580 -1925 7700 -1885
rect 7580 -1955 7625 -1925
rect 7655 -1955 7700 -1925
rect 7580 -1995 7700 -1955
rect 7580 -2025 7625 -1995
rect 7655 -2025 7700 -1995
rect 7580 -2060 7700 -2025
rect 7580 -2090 7625 -2060
rect 7655 -2090 7700 -2060
rect 7580 -2120 7700 -2090
rect 7580 -2150 7625 -2120
rect 7655 -2150 7700 -2120
rect 7580 -2185 7700 -2150
rect 7580 -2215 7625 -2185
rect 7655 -2215 7700 -2185
rect 7580 -2255 7700 -2215
rect 7580 -2285 7625 -2255
rect 7655 -2285 7700 -2255
rect 7580 -2325 7700 -2285
rect 7580 -2355 7625 -2325
rect 7655 -2355 7700 -2325
rect 7580 -2395 7700 -2355
rect 7580 -2425 7625 -2395
rect 7655 -2425 7700 -2395
rect 7580 -2460 7700 -2425
rect 7580 -2490 7625 -2460
rect 7655 -2490 7700 -2460
rect 7580 -2520 7700 -2490
rect 7580 -2550 7625 -2520
rect 7655 -2550 7700 -2520
rect 7580 -2585 7700 -2550
rect 7580 -2615 7625 -2585
rect 7655 -2615 7700 -2585
rect 7580 -2655 7700 -2615
rect 7580 -2685 7625 -2655
rect 7655 -2685 7700 -2655
rect 7580 -2725 7700 -2685
rect 7580 -2755 7625 -2725
rect 7655 -2755 7700 -2725
rect 7580 -2795 7700 -2755
rect 7580 -2825 7625 -2795
rect 7655 -2825 7700 -2795
rect 7580 -2860 7700 -2825
rect 7580 -2890 7625 -2860
rect 7655 -2890 7700 -2860
rect 7580 -2905 7700 -2890
rect 7930 -1320 8050 -1225
rect 7930 -1350 7975 -1320
rect 8005 -1350 8050 -1320
rect 7930 -1385 8050 -1350
rect 7930 -1415 7975 -1385
rect 8005 -1415 8050 -1385
rect 7930 -1455 8050 -1415
rect 7930 -1485 7975 -1455
rect 8005 -1485 8050 -1455
rect 7930 -1525 8050 -1485
rect 7930 -1555 7975 -1525
rect 8005 -1555 8050 -1525
rect 7930 -1595 8050 -1555
rect 7930 -1625 7975 -1595
rect 8005 -1625 8050 -1595
rect 7930 -1660 8050 -1625
rect 7930 -1690 7975 -1660
rect 8005 -1690 8050 -1660
rect 7930 -1720 8050 -1690
rect 7930 -1750 7975 -1720
rect 8005 -1750 8050 -1720
rect 7930 -1785 8050 -1750
rect 7930 -1815 7975 -1785
rect 8005 -1815 8050 -1785
rect 7930 -1855 8050 -1815
rect 7930 -1885 7975 -1855
rect 8005 -1885 8050 -1855
rect 7930 -1925 8050 -1885
rect 7930 -1955 7975 -1925
rect 8005 -1955 8050 -1925
rect 7930 -1995 8050 -1955
rect 7930 -2025 7975 -1995
rect 8005 -2025 8050 -1995
rect 7930 -2060 8050 -2025
rect 7930 -2090 7975 -2060
rect 8005 -2090 8050 -2060
rect 7930 -2120 8050 -2090
rect 7930 -2150 7975 -2120
rect 8005 -2150 8050 -2120
rect 7930 -2185 8050 -2150
rect 7930 -2215 7975 -2185
rect 8005 -2215 8050 -2185
rect 7930 -2255 8050 -2215
rect 7930 -2285 7975 -2255
rect 8005 -2285 8050 -2255
rect 7930 -2325 8050 -2285
rect 7930 -2355 7975 -2325
rect 8005 -2355 8050 -2325
rect 7930 -2395 8050 -2355
rect 7930 -2425 7975 -2395
rect 8005 -2425 8050 -2395
rect 7930 -2460 8050 -2425
rect 7930 -2490 7975 -2460
rect 8005 -2490 8050 -2460
rect 7930 -2520 8050 -2490
rect 7930 -2550 7975 -2520
rect 8005 -2550 8050 -2520
rect 7930 -2585 8050 -2550
rect 7930 -2615 7975 -2585
rect 8005 -2615 8050 -2585
rect 7930 -2655 8050 -2615
rect 7930 -2685 7975 -2655
rect 8005 -2685 8050 -2655
rect 7930 -2725 8050 -2685
rect 7930 -2755 7975 -2725
rect 8005 -2755 8050 -2725
rect 7930 -2795 8050 -2755
rect 7930 -2825 7975 -2795
rect 8005 -2825 8050 -2795
rect 7930 -2860 8050 -2825
rect 7930 -2890 7975 -2860
rect 8005 -2890 8050 -2860
rect 7930 -2905 8050 -2890
rect 8280 -1320 8400 -1225
rect 8280 -1350 8325 -1320
rect 8355 -1350 8400 -1320
rect 8280 -1385 8400 -1350
rect 8280 -1415 8325 -1385
rect 8355 -1415 8400 -1385
rect 8280 -1455 8400 -1415
rect 8280 -1485 8325 -1455
rect 8355 -1485 8400 -1455
rect 8280 -1525 8400 -1485
rect 8280 -1555 8325 -1525
rect 8355 -1555 8400 -1525
rect 8280 -1595 8400 -1555
rect 8280 -1625 8325 -1595
rect 8355 -1625 8400 -1595
rect 8280 -1660 8400 -1625
rect 8280 -1690 8325 -1660
rect 8355 -1690 8400 -1660
rect 8280 -1720 8400 -1690
rect 8280 -1750 8325 -1720
rect 8355 -1750 8400 -1720
rect 8280 -1785 8400 -1750
rect 8280 -1815 8325 -1785
rect 8355 -1815 8400 -1785
rect 8280 -1855 8400 -1815
rect 8280 -1885 8325 -1855
rect 8355 -1885 8400 -1855
rect 8280 -1925 8400 -1885
rect 8280 -1955 8325 -1925
rect 8355 -1955 8400 -1925
rect 8280 -1995 8400 -1955
rect 8280 -2025 8325 -1995
rect 8355 -2025 8400 -1995
rect 8280 -2060 8400 -2025
rect 8280 -2090 8325 -2060
rect 8355 -2090 8400 -2060
rect 8280 -2120 8400 -2090
rect 8280 -2150 8325 -2120
rect 8355 -2150 8400 -2120
rect 8280 -2185 8400 -2150
rect 8280 -2215 8325 -2185
rect 8355 -2215 8400 -2185
rect 8280 -2255 8400 -2215
rect 8280 -2285 8325 -2255
rect 8355 -2285 8400 -2255
rect 8280 -2325 8400 -2285
rect 8280 -2355 8325 -2325
rect 8355 -2355 8400 -2325
rect 8280 -2395 8400 -2355
rect 8280 -2425 8325 -2395
rect 8355 -2425 8400 -2395
rect 8280 -2460 8400 -2425
rect 8280 -2490 8325 -2460
rect 8355 -2490 8400 -2460
rect 8280 -2520 8400 -2490
rect 8280 -2550 8325 -2520
rect 8355 -2550 8400 -2520
rect 8280 -2585 8400 -2550
rect 8280 -2615 8325 -2585
rect 8355 -2615 8400 -2585
rect 8280 -2655 8400 -2615
rect 8280 -2685 8325 -2655
rect 8355 -2685 8400 -2655
rect 8280 -2725 8400 -2685
rect 8280 -2755 8325 -2725
rect 8355 -2755 8400 -2725
rect 8280 -2795 8400 -2755
rect 8280 -2825 8325 -2795
rect 8355 -2825 8400 -2795
rect 8280 -2860 8400 -2825
rect 8280 -2890 8325 -2860
rect 8355 -2890 8400 -2860
rect 8280 -2905 8400 -2890
rect 8630 -1320 8750 -1225
rect 8630 -1350 8675 -1320
rect 8705 -1350 8750 -1320
rect 8630 -1385 8750 -1350
rect 8630 -1415 8675 -1385
rect 8705 -1415 8750 -1385
rect 8630 -1455 8750 -1415
rect 8630 -1485 8675 -1455
rect 8705 -1485 8750 -1455
rect 8630 -1525 8750 -1485
rect 8630 -1555 8675 -1525
rect 8705 -1555 8750 -1525
rect 8630 -1595 8750 -1555
rect 8630 -1625 8675 -1595
rect 8705 -1625 8750 -1595
rect 8630 -1660 8750 -1625
rect 8630 -1690 8675 -1660
rect 8705 -1690 8750 -1660
rect 8630 -1720 8750 -1690
rect 8630 -1750 8675 -1720
rect 8705 -1750 8750 -1720
rect 8630 -1785 8750 -1750
rect 8630 -1815 8675 -1785
rect 8705 -1815 8750 -1785
rect 8630 -1855 8750 -1815
rect 8630 -1885 8675 -1855
rect 8705 -1885 8750 -1855
rect 8630 -1925 8750 -1885
rect 8630 -1955 8675 -1925
rect 8705 -1955 8750 -1925
rect 8630 -1995 8750 -1955
rect 8630 -2025 8675 -1995
rect 8705 -2025 8750 -1995
rect 8630 -2060 8750 -2025
rect 8630 -2090 8675 -2060
rect 8705 -2090 8750 -2060
rect 8630 -2120 8750 -2090
rect 8630 -2150 8675 -2120
rect 8705 -2150 8750 -2120
rect 8630 -2185 8750 -2150
rect 8630 -2215 8675 -2185
rect 8705 -2215 8750 -2185
rect 8630 -2255 8750 -2215
rect 8630 -2285 8675 -2255
rect 8705 -2285 8750 -2255
rect 8630 -2325 8750 -2285
rect 8630 -2355 8675 -2325
rect 8705 -2355 8750 -2325
rect 8630 -2395 8750 -2355
rect 8630 -2425 8675 -2395
rect 8705 -2425 8750 -2395
rect 8630 -2460 8750 -2425
rect 8630 -2490 8675 -2460
rect 8705 -2490 8750 -2460
rect 8630 -2520 8750 -2490
rect 8630 -2550 8675 -2520
rect 8705 -2550 8750 -2520
rect 8630 -2585 8750 -2550
rect 8630 -2615 8675 -2585
rect 8705 -2615 8750 -2585
rect 8630 -2655 8750 -2615
rect 8630 -2685 8675 -2655
rect 8705 -2685 8750 -2655
rect 8630 -2725 8750 -2685
rect 8630 -2755 8675 -2725
rect 8705 -2755 8750 -2725
rect 8630 -2795 8750 -2755
rect 8630 -2825 8675 -2795
rect 8705 -2825 8750 -2795
rect 8630 -2860 8750 -2825
rect 8630 -2890 8675 -2860
rect 8705 -2890 8750 -2860
rect 8630 -2905 8750 -2890
rect 8980 -1320 9100 -1225
rect 8980 -1350 9025 -1320
rect 9055 -1350 9100 -1320
rect 8980 -1385 9100 -1350
rect 8980 -1415 9025 -1385
rect 9055 -1415 9100 -1385
rect 8980 -1455 9100 -1415
rect 8980 -1485 9025 -1455
rect 9055 -1485 9100 -1455
rect 8980 -1525 9100 -1485
rect 8980 -1555 9025 -1525
rect 9055 -1555 9100 -1525
rect 8980 -1595 9100 -1555
rect 8980 -1625 9025 -1595
rect 9055 -1625 9100 -1595
rect 8980 -1660 9100 -1625
rect 8980 -1690 9025 -1660
rect 9055 -1690 9100 -1660
rect 8980 -1720 9100 -1690
rect 8980 -1750 9025 -1720
rect 9055 -1750 9100 -1720
rect 8980 -1785 9100 -1750
rect 8980 -1815 9025 -1785
rect 9055 -1815 9100 -1785
rect 8980 -1855 9100 -1815
rect 8980 -1885 9025 -1855
rect 9055 -1885 9100 -1855
rect 8980 -1925 9100 -1885
rect 8980 -1955 9025 -1925
rect 9055 -1955 9100 -1925
rect 8980 -1995 9100 -1955
rect 8980 -2025 9025 -1995
rect 9055 -2025 9100 -1995
rect 8980 -2060 9100 -2025
rect 8980 -2090 9025 -2060
rect 9055 -2090 9100 -2060
rect 8980 -2120 9100 -2090
rect 8980 -2150 9025 -2120
rect 9055 -2150 9100 -2120
rect 8980 -2185 9100 -2150
rect 8980 -2215 9025 -2185
rect 9055 -2215 9100 -2185
rect 8980 -2255 9100 -2215
rect 8980 -2285 9025 -2255
rect 9055 -2285 9100 -2255
rect 8980 -2325 9100 -2285
rect 8980 -2355 9025 -2325
rect 9055 -2355 9100 -2325
rect 8980 -2395 9100 -2355
rect 8980 -2425 9025 -2395
rect 9055 -2425 9100 -2395
rect 8980 -2460 9100 -2425
rect 8980 -2490 9025 -2460
rect 9055 -2490 9100 -2460
rect 8980 -2520 9100 -2490
rect 8980 -2550 9025 -2520
rect 9055 -2550 9100 -2520
rect 8980 -2585 9100 -2550
rect 8980 -2615 9025 -2585
rect 9055 -2615 9100 -2585
rect 8980 -2655 9100 -2615
rect 8980 -2685 9025 -2655
rect 9055 -2685 9100 -2655
rect 8980 -2725 9100 -2685
rect 8980 -2755 9025 -2725
rect 9055 -2755 9100 -2725
rect 8980 -2795 9100 -2755
rect 8980 -2825 9025 -2795
rect 9055 -2825 9100 -2795
rect 8980 -2860 9100 -2825
rect 8980 -2890 9025 -2860
rect 9055 -2890 9100 -2860
rect 8980 -2905 9100 -2890
rect 5480 -3050 5525 -3020
rect 5555 -3050 5600 -3020
rect 5480 -3085 5600 -3050
rect 5480 -3115 5525 -3085
rect 5555 -3115 5600 -3085
rect 5480 -3155 5600 -3115
rect 5480 -3185 5525 -3155
rect 5555 -3185 5600 -3155
rect 5480 -3225 5600 -3185
rect 5480 -3255 5525 -3225
rect 5555 -3255 5600 -3225
rect 5480 -3295 5600 -3255
rect 5480 -3325 5525 -3295
rect 5555 -3325 5600 -3295
rect 5480 -3360 5600 -3325
rect 5480 -3390 5525 -3360
rect 5555 -3390 5600 -3360
rect 5480 -3420 5600 -3390
rect 5480 -3450 5525 -3420
rect 5555 -3450 5600 -3420
rect 5480 -3485 5600 -3450
rect 5480 -3515 5525 -3485
rect 5555 -3515 5600 -3485
rect 5480 -3555 5600 -3515
rect 5480 -3585 5525 -3555
rect 5555 -3585 5600 -3555
rect 5480 -3625 5600 -3585
rect 5480 -3655 5525 -3625
rect 5555 -3655 5600 -3625
rect 5480 -3695 5600 -3655
rect 5480 -3725 5525 -3695
rect 5555 -3725 5600 -3695
rect 5480 -3760 5600 -3725
rect 5480 -3790 5525 -3760
rect 5555 -3790 5600 -3760
rect 5480 -3820 5600 -3790
rect 5480 -3850 5525 -3820
rect 5555 -3850 5600 -3820
rect 5480 -3885 5600 -3850
rect 5480 -3915 5525 -3885
rect 5555 -3915 5600 -3885
rect 5480 -3955 5600 -3915
rect 5480 -3985 5525 -3955
rect 5555 -3985 5600 -3955
rect 5480 -4025 5600 -3985
rect 5480 -4055 5525 -4025
rect 5555 -4055 5600 -4025
rect 5480 -4095 5600 -4055
rect 5480 -4125 5525 -4095
rect 5555 -4125 5600 -4095
rect 5480 -4160 5600 -4125
rect 5480 -4190 5525 -4160
rect 5555 -4190 5600 -4160
rect 5480 -4220 5600 -4190
rect 5480 -4250 5525 -4220
rect 5555 -4250 5600 -4220
rect 5480 -4285 5600 -4250
rect 5480 -4315 5525 -4285
rect 5555 -4315 5600 -4285
rect 5480 -4355 5600 -4315
rect 5480 -4385 5525 -4355
rect 5555 -4385 5600 -4355
rect 5480 -4425 5600 -4385
rect 5480 -4455 5525 -4425
rect 5555 -4455 5600 -4425
rect 5480 -4495 5600 -4455
rect 5480 -4525 5525 -4495
rect 5555 -4525 5600 -4495
rect 5480 -4560 5600 -4525
rect 5480 -4590 5525 -4560
rect 5555 -4590 5600 -4560
rect 5480 -4605 5600 -4590
<< via1 >>
rect 2115 19280 2145 19310
rect 2115 19215 2145 19245
rect 2115 19145 2145 19175
rect 2115 19075 2145 19105
rect 2115 19005 2145 19035
rect 2115 18940 2145 18970
rect 2115 18880 2145 18910
rect 2115 18815 2145 18845
rect 2115 18745 2145 18775
rect 2115 18675 2145 18705
rect 2115 18605 2145 18635
rect 2115 18540 2145 18570
rect 2115 18480 2145 18510
rect 2115 18415 2145 18445
rect 2115 18345 2145 18375
rect 2115 18275 2145 18305
rect 2115 18205 2145 18235
rect 2115 18140 2145 18170
rect 2115 18080 2145 18110
rect 2115 18015 2145 18045
rect 2115 17945 2145 17975
rect 2115 17875 2145 17905
rect 2115 17805 2145 17835
rect 2115 17740 2145 17770
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 2075 15660 2105 15690
rect 2115 15660 2145 15690
rect 2155 15660 2185 15690
rect 2075 15620 2105 15650
rect 2115 15620 2145 15650
rect 2155 15620 2185 15650
rect 2075 15580 2105 15610
rect 2115 15580 2145 15610
rect 2155 15580 2185 15610
rect 2075 12680 2105 12710
rect 2115 12680 2145 12710
rect 2155 12680 2185 12710
rect 2075 12640 2105 12670
rect 2115 12640 2145 12670
rect 2155 12640 2185 12670
rect 2075 12520 2105 12550
rect 2115 12520 2145 12550
rect 2155 12520 2185 12550
rect 2075 12480 2105 12510
rect 2115 12480 2145 12510
rect 2155 12480 2185 12510
rect 2075 12440 2105 12470
rect 2115 12440 2145 12470
rect 2155 12440 2185 12470
rect 2210 15895 2240 15925
rect 2250 15895 2280 15925
rect 2290 15895 2320 15925
rect 1325 9605 1355 9635
rect 1325 9540 1355 9570
rect 1325 9470 1355 9500
rect 1325 9400 1355 9430
rect 1325 9330 1355 9360
rect 1325 9265 1355 9295
rect 1325 9205 1355 9235
rect 1325 9140 1355 9170
rect 1325 9070 1355 9100
rect 1325 9000 1355 9030
rect 1325 8930 1355 8960
rect 1325 8865 1355 8895
rect 1325 8805 1355 8835
rect 1325 8740 1355 8770
rect 1325 8670 1355 8700
rect 1325 8600 1355 8630
rect 1325 8530 1355 8560
rect 1325 8465 1355 8495
rect 1325 8405 1355 8435
rect 1325 8340 1355 8370
rect 1325 8270 1355 8300
rect 1325 8200 1355 8230
rect 1325 8130 1355 8160
rect 6665 15565 6695 15595
rect 6705 15565 6735 15595
rect 6745 15565 6775 15595
rect 6665 15525 6695 15555
rect 6705 15525 6735 15555
rect 6745 15525 6775 15555
rect 6665 15485 6695 15515
rect 6705 15485 6735 15515
rect 6745 15485 6775 15515
rect 2250 9605 2280 9635
rect 2250 9540 2280 9570
rect 2250 9470 2280 9500
rect 2250 9400 2280 9430
rect 2250 9330 2280 9360
rect 2250 9265 2280 9295
rect 2250 9205 2280 9235
rect 2250 9140 2280 9170
rect 2250 9070 2280 9100
rect 2250 9000 2280 9030
rect 2250 8930 2280 8960
rect 2250 8865 2280 8895
rect 2250 8805 2280 8835
rect 2250 8740 2280 8770
rect 2250 8670 2280 8700
rect 2250 8600 2280 8630
rect 2250 8530 2280 8560
rect 2250 8465 2280 8495
rect 2250 8405 2280 8435
rect 2250 8340 2280 8370
rect 2250 8270 2280 8300
rect 2250 8200 2280 8230
rect 2250 8130 2280 8160
rect 1985 8055 2015 8085
rect 2025 8055 2055 8085
rect 2065 8055 2095 8085
rect 1635 8000 1665 8030
rect 1675 8000 1705 8030
rect 1715 8000 1745 8030
rect 2480 8055 2510 8085
rect 3180 7925 3210 7955
rect 3240 7925 3270 7955
rect 3180 7855 3210 7885
rect 3240 7855 3270 7885
rect 3180 7785 3210 7815
rect 3240 7785 3270 7815
rect 3180 7715 3210 7745
rect 3240 7715 3270 7745
rect 3180 7650 3210 7680
rect 3240 7650 3270 7680
rect 3180 7590 3210 7620
rect 3240 7590 3270 7620
rect 3180 7525 3210 7555
rect 3240 7525 3270 7555
rect 3180 7455 3210 7485
rect 3240 7455 3270 7485
rect 3180 7385 3210 7415
rect 3240 7385 3270 7415
rect 3180 7315 3210 7345
rect 3240 7315 3270 7345
rect 3180 7250 3210 7280
rect 3240 7250 3270 7280
rect 3180 7190 3210 7220
rect 3240 7190 3270 7220
rect 3180 7125 3210 7155
rect 3240 7125 3270 7155
rect 3180 7055 3210 7085
rect 3240 7055 3270 7085
rect 3180 6985 3210 7015
rect 3240 6985 3270 7015
rect 3180 6915 3210 6945
rect 3240 6915 3270 6945
rect 3180 6850 3210 6880
rect 3240 6850 3270 6880
rect 3180 6790 3210 6820
rect 3240 6790 3270 6820
rect 3180 6725 3210 6755
rect 3240 6725 3270 6755
rect 3180 6655 3210 6685
rect 3240 6655 3270 6685
rect 3180 6585 3210 6615
rect 3240 6585 3270 6615
rect 3180 6515 3210 6545
rect 3240 6515 3270 6545
rect 3180 6450 3210 6480
rect 3240 6450 3270 6480
rect 2850 6385 2880 6415
rect 2720 6275 2750 6305
rect 3635 8000 3665 8030
rect 3855 8000 3885 8030
rect 3350 7925 3380 7955
rect 3350 7855 3380 7885
rect 3350 7785 3380 7815
rect 3350 7715 3380 7745
rect 3350 7650 3380 7680
rect 3350 7590 3380 7620
rect 3350 7525 3380 7555
rect 3350 7455 3380 7485
rect 3350 7385 3380 7415
rect 3350 7315 3380 7345
rect 3350 7250 3380 7280
rect 3350 7190 3380 7220
rect 3350 7125 3380 7155
rect 3350 7055 3380 7085
rect 3350 6985 3380 7015
rect 3350 6915 3380 6945
rect 3350 6850 3380 6880
rect 3350 6790 3380 6820
rect 3350 6725 3380 6755
rect 3350 6655 3380 6685
rect 3350 6585 3380 6615
rect 3350 6515 3380 6545
rect 3350 6450 3380 6480
rect 3385 6385 3415 6415
rect 3080 6275 3110 6305
rect 3295 6270 3325 6300
rect 935 6160 965 6190
rect 975 6160 1005 6190
rect 1015 6160 1045 6190
rect 935 6120 965 6150
rect 975 6120 1005 6150
rect 1015 6120 1045 6150
rect 935 6080 965 6110
rect 975 6080 1005 6110
rect 1015 6080 1045 6110
rect 3080 5045 3110 5075
rect 3440 6215 3470 6245
rect 3385 3760 3415 3790
rect 4310 6160 4340 6190
rect 4310 6120 4340 6150
rect 4310 6080 4340 6110
rect 4475 6270 4505 6300
rect 4475 6215 4505 6245
rect 4420 6160 4450 6190
rect 4420 6120 4450 6150
rect 4420 6080 4450 6110
rect 4530 6160 4560 6190
rect 4530 6120 4560 6150
rect 4530 6080 4560 6110
rect 5315 7985 5345 8015
rect 5475 6385 5505 6415
rect 6150 6385 6180 6415
rect 4640 6160 4670 6190
rect 4640 6120 4670 6150
rect 4640 6080 4670 6110
rect 5550 6215 5580 6245
rect 5475 3820 5505 3850
rect 3440 3080 3470 3110
rect 4475 3080 4505 3110
rect 5875 5390 5905 5420
rect 5625 4990 5655 5020
rect 6665 12895 6695 12925
rect 6705 12895 6735 12925
rect 6745 12895 6775 12925
rect 6665 12855 6695 12885
rect 6705 12855 6735 12885
rect 6745 12855 6775 12885
rect 6665 12815 6695 12845
rect 6705 12815 6735 12845
rect 6745 12815 6775 12845
rect 6665 12120 6695 12150
rect 6705 12120 6735 12150
rect 6745 12120 6775 12150
rect 6665 12080 6695 12110
rect 6705 12080 6735 12110
rect 6745 12080 6775 12110
rect 6665 12040 6695 12070
rect 6705 12040 6735 12070
rect 6745 12040 6775 12070
rect 6665 11135 6695 11165
rect 6705 11135 6735 11165
rect 6745 11135 6775 11165
rect 6665 11095 6695 11125
rect 6705 11095 6735 11125
rect 6745 11095 6775 11125
rect 6665 11055 6695 11085
rect 6705 11055 6735 11085
rect 6745 11055 6775 11085
rect 6665 10410 6695 10440
rect 6705 10410 6735 10440
rect 6745 10410 6775 10440
rect 6665 10370 6695 10400
rect 6705 10370 6735 10400
rect 6745 10370 6775 10400
rect 6665 10330 6695 10360
rect 6705 10330 6735 10360
rect 6745 10330 6775 10360
rect 6665 10050 6695 10080
rect 6705 10050 6735 10080
rect 6745 10050 6775 10080
rect 6665 10010 6695 10040
rect 6705 10010 6735 10040
rect 6745 10010 6775 10040
rect 6665 9970 6695 10000
rect 6705 9970 6735 10000
rect 6745 9970 6775 10000
rect 6705 9540 6735 9570
rect 6705 9470 6735 9500
rect 6705 9400 6735 9430
rect 6705 9330 6735 9360
rect 6705 9265 6735 9295
rect 6705 9205 6735 9235
rect 6705 9140 6735 9170
rect 6705 9070 6735 9100
rect 6705 9000 6735 9030
rect 6705 8930 6735 8960
rect 6705 8865 6735 8895
rect 6705 8805 6735 8835
rect 6705 8740 6735 8770
rect 6705 8670 6735 8700
rect 6705 8600 6735 8630
rect 6705 8530 6735 8560
rect 6705 8465 6735 8495
rect 6705 8405 6735 8435
rect 6705 8340 6735 8370
rect 6705 8270 6735 8300
rect 6705 8200 6735 8230
rect 6705 8130 6735 8160
rect 7625 9605 7655 9635
rect 7625 9540 7655 9570
rect 7625 9470 7655 9500
rect 7625 9400 7655 9430
rect 7625 9330 7655 9360
rect 7625 9265 7655 9295
rect 7625 9205 7655 9235
rect 7625 9140 7655 9170
rect 7625 9070 7655 9100
rect 7625 9000 7655 9030
rect 7625 8930 7655 8960
rect 7625 8865 7655 8895
rect 7625 8805 7655 8835
rect 7625 8740 7655 8770
rect 7625 8670 7655 8700
rect 7625 8600 7655 8630
rect 7625 8530 7655 8560
rect 7625 8465 7655 8495
rect 7625 8405 7655 8435
rect 7625 8340 7655 8370
rect 7625 8270 7655 8300
rect 7625 8200 7655 8230
rect 7625 8130 7655 8160
rect 6470 8040 6500 8070
rect 6885 8040 6915 8070
rect 6925 8040 6955 8070
rect 6965 8040 6995 8070
rect 7235 7985 7265 8015
rect 7275 7985 7305 8015
rect 7315 7985 7345 8015
rect 6225 5390 6255 5420
rect 7935 6160 7965 6190
rect 7975 6160 8005 6190
rect 8015 6160 8045 6190
rect 7935 6120 7965 6150
rect 7975 6120 8005 6150
rect 8015 6120 8045 6150
rect 7935 6080 7965 6110
rect 7975 6080 8005 6110
rect 8015 6080 8045 6110
rect 5875 4990 5905 5020
rect 5625 4395 5655 4425
rect 5550 3080 5580 3110
rect 4475 2860 4505 2890
rect 935 1115 965 1145
rect 975 1115 1005 1145
rect 1015 1115 1045 1145
rect 935 1075 965 1105
rect 975 1075 1005 1105
rect 1015 1075 1045 1105
rect 935 1035 965 1065
rect 975 1035 1005 1065
rect 1015 1035 1045 1065
rect 4420 1115 4450 1145
rect 4420 1075 4450 1105
rect 4420 1035 4450 1065
rect 4530 1115 4560 1145
rect 4530 1075 4560 1105
rect 4530 1035 4560 1065
rect 7935 1115 7965 1145
rect 7975 1115 8005 1145
rect 8015 1115 8045 1145
rect 7935 1075 7965 1105
rect 7975 1075 8005 1105
rect 8015 1075 8045 1105
rect 7935 1035 7965 1065
rect 7975 1035 8005 1065
rect 8015 1035 8045 1065
rect -75 -1350 -45 -1320
rect -75 -1415 -45 -1385
rect -75 -1485 -45 -1455
rect -75 -1555 -45 -1525
rect -75 -1625 -45 -1595
rect -75 -1690 -45 -1660
rect -75 -1750 -45 -1720
rect -75 -1815 -45 -1785
rect -75 -1885 -45 -1855
rect -75 -1955 -45 -1925
rect -75 -2025 -45 -1995
rect -75 -2090 -45 -2060
rect -75 -2150 -45 -2120
rect -75 -2215 -45 -2185
rect -75 -2285 -45 -2255
rect -75 -2355 -45 -2325
rect -75 -2425 -45 -2395
rect -75 -2490 -45 -2460
rect -75 -2550 -45 -2520
rect -75 -2615 -45 -2585
rect -75 -2685 -45 -2655
rect -75 -2755 -45 -2725
rect -75 -2825 -45 -2795
rect -75 -2890 -45 -2860
rect 275 -1350 305 -1320
rect 275 -1415 305 -1385
rect 275 -1485 305 -1455
rect 275 -1555 305 -1525
rect 275 -1625 305 -1595
rect 275 -1690 305 -1660
rect 275 -1750 305 -1720
rect 275 -1815 305 -1785
rect 275 -1885 305 -1855
rect 275 -1955 305 -1925
rect 275 -2025 305 -1995
rect 275 -2090 305 -2060
rect 275 -2150 305 -2120
rect 275 -2215 305 -2185
rect 275 -2285 305 -2255
rect 275 -2355 305 -2325
rect 275 -2425 305 -2395
rect 275 -2490 305 -2460
rect 275 -2550 305 -2520
rect 275 -2615 305 -2585
rect 275 -2685 305 -2655
rect 275 -2755 305 -2725
rect 275 -2825 305 -2795
rect 275 -2890 305 -2860
rect 625 -1350 655 -1320
rect 625 -1415 655 -1385
rect 625 -1485 655 -1455
rect 625 -1555 655 -1525
rect 625 -1625 655 -1595
rect 625 -1690 655 -1660
rect 625 -1750 655 -1720
rect 625 -1815 655 -1785
rect 625 -1885 655 -1855
rect 625 -1955 655 -1925
rect 625 -2025 655 -1995
rect 625 -2090 655 -2060
rect 625 -2150 655 -2120
rect 625 -2215 655 -2185
rect 625 -2285 655 -2255
rect 625 -2355 655 -2325
rect 625 -2425 655 -2395
rect 625 -2490 655 -2460
rect 625 -2550 655 -2520
rect 625 -2615 655 -2585
rect 625 -2685 655 -2655
rect 625 -2755 655 -2725
rect 625 -2825 655 -2795
rect 625 -2890 655 -2860
rect 975 -1350 1005 -1320
rect 975 -1415 1005 -1385
rect 975 -1485 1005 -1455
rect 975 -1555 1005 -1525
rect 975 -1625 1005 -1595
rect 975 -1690 1005 -1660
rect 975 -1750 1005 -1720
rect 975 -1815 1005 -1785
rect 975 -1885 1005 -1855
rect 975 -1955 1005 -1925
rect 975 -2025 1005 -1995
rect 975 -2090 1005 -2060
rect 975 -2150 1005 -2120
rect 975 -2215 1005 -2185
rect 975 -2285 1005 -2255
rect 975 -2355 1005 -2325
rect 975 -2425 1005 -2395
rect 975 -2490 1005 -2460
rect 975 -2550 1005 -2520
rect 975 -2615 1005 -2585
rect 975 -2685 1005 -2655
rect 975 -2755 1005 -2725
rect 975 -2825 1005 -2795
rect 975 -2890 1005 -2860
rect 1325 -1350 1355 -1320
rect 1325 -1415 1355 -1385
rect 1325 -1485 1355 -1455
rect 1325 -1555 1355 -1525
rect 1325 -1625 1355 -1595
rect 1325 -1690 1355 -1660
rect 1325 -1750 1355 -1720
rect 1325 -1815 1355 -1785
rect 1325 -1885 1355 -1855
rect 1325 -1955 1355 -1925
rect 1325 -2025 1355 -1995
rect 1325 -2090 1355 -2060
rect 1325 -2150 1355 -2120
rect 1325 -2215 1355 -2185
rect 1325 -2285 1355 -2255
rect 1325 -2355 1355 -2325
rect 1325 -2425 1355 -2395
rect 1325 -2490 1355 -2460
rect 1325 -2550 1355 -2520
rect 1325 -2615 1355 -2585
rect 1325 -2685 1355 -2655
rect 1325 -2755 1355 -2725
rect 1325 -2825 1355 -2795
rect 1325 -2890 1355 -2860
rect 1675 -1350 1705 -1320
rect 1675 -1415 1705 -1385
rect 1675 -1485 1705 -1455
rect 1675 -1555 1705 -1525
rect 1675 -1625 1705 -1595
rect 1675 -1690 1705 -1660
rect 1675 -1750 1705 -1720
rect 1675 -1815 1705 -1785
rect 1675 -1885 1705 -1855
rect 1675 -1955 1705 -1925
rect 1675 -2025 1705 -1995
rect 1675 -2090 1705 -2060
rect 1675 -2150 1705 -2120
rect 1675 -2215 1705 -2185
rect 1675 -2285 1705 -2255
rect 1675 -2355 1705 -2325
rect 1675 -2425 1705 -2395
rect 1675 -2490 1705 -2460
rect 1675 -2550 1705 -2520
rect 1675 -2615 1705 -2585
rect 1675 -2685 1705 -2655
rect 1675 -2755 1705 -2725
rect 1675 -2825 1705 -2795
rect 1675 -2890 1705 -2860
rect 2025 -1350 2055 -1320
rect 2025 -1415 2055 -1385
rect 2025 -1485 2055 -1455
rect 2025 -1555 2055 -1525
rect 2025 -1625 2055 -1595
rect 2025 -1690 2055 -1660
rect 2025 -1750 2055 -1720
rect 2025 -1815 2055 -1785
rect 2025 -1885 2055 -1855
rect 2025 -1955 2055 -1925
rect 2025 -2025 2055 -1995
rect 2025 -2090 2055 -2060
rect 2025 -2150 2055 -2120
rect 2025 -2215 2055 -2185
rect 2025 -2285 2055 -2255
rect 2025 -2355 2055 -2325
rect 2025 -2425 2055 -2395
rect 2025 -2490 2055 -2460
rect 2025 -2550 2055 -2520
rect 2025 -2615 2055 -2585
rect 2025 -2685 2055 -2655
rect 2025 -2755 2055 -2725
rect 2025 -2825 2055 -2795
rect 2025 -2890 2055 -2860
rect 2375 -1350 2405 -1320
rect 2375 -1415 2405 -1385
rect 2375 -1485 2405 -1455
rect 2375 -1555 2405 -1525
rect 2375 -1625 2405 -1595
rect 2375 -1690 2405 -1660
rect 2375 -1750 2405 -1720
rect 2375 -1815 2405 -1785
rect 2375 -1885 2405 -1855
rect 2375 -1955 2405 -1925
rect 2375 -2025 2405 -1995
rect 2375 -2090 2405 -2060
rect 2375 -2150 2405 -2120
rect 2375 -2215 2405 -2185
rect 2375 -2285 2405 -2255
rect 2375 -2355 2405 -2325
rect 2375 -2425 2405 -2395
rect 2375 -2490 2405 -2460
rect 2375 -2550 2405 -2520
rect 2375 -2615 2405 -2585
rect 2375 -2685 2405 -2655
rect 2375 -2755 2405 -2725
rect 2375 -2825 2405 -2795
rect 2375 -2890 2405 -2860
rect 2725 -1350 2755 -1320
rect 2725 -1415 2755 -1385
rect 2725 -1485 2755 -1455
rect 2725 -1555 2755 -1525
rect 2725 -1625 2755 -1595
rect 2725 -1690 2755 -1660
rect 2725 -1750 2755 -1720
rect 2725 -1815 2755 -1785
rect 2725 -1885 2755 -1855
rect 2725 -1955 2755 -1925
rect 2725 -2025 2755 -1995
rect 2725 -2090 2755 -2060
rect 2725 -2150 2755 -2120
rect 2725 -2215 2755 -2185
rect 2725 -2285 2755 -2255
rect 2725 -2355 2755 -2325
rect 2725 -2425 2755 -2395
rect 2725 -2490 2755 -2460
rect 2725 -2550 2755 -2520
rect 2725 -2615 2755 -2585
rect 2725 -2685 2755 -2655
rect 2725 -2755 2755 -2725
rect 2725 -2825 2755 -2795
rect 2725 -2890 2755 -2860
rect 3075 -1350 3105 -1320
rect 3075 -1415 3105 -1385
rect 3075 -1485 3105 -1455
rect 3075 -1555 3105 -1525
rect 3075 -1625 3105 -1595
rect 3075 -1690 3105 -1660
rect 3075 -1750 3105 -1720
rect 3075 -1815 3105 -1785
rect 3075 -1885 3105 -1855
rect 3075 -1955 3105 -1925
rect 3075 -2025 3105 -1995
rect 3075 -2090 3105 -2060
rect 3075 -2150 3105 -2120
rect 3075 -2215 3105 -2185
rect 3075 -2285 3105 -2255
rect 3075 -2355 3105 -2325
rect 3075 -2425 3105 -2395
rect 3075 -2490 3105 -2460
rect 3075 -2550 3105 -2520
rect 3075 -2615 3105 -2585
rect 3075 -2685 3105 -2655
rect 3075 -2755 3105 -2725
rect 3075 -2825 3105 -2795
rect 3075 -2890 3105 -2860
rect 3425 -3050 3455 -3020
rect 3425 -3115 3455 -3085
rect 3425 -3185 3455 -3155
rect 3425 -3255 3455 -3225
rect 3425 -3325 3455 -3295
rect 3425 -3390 3455 -3360
rect 3425 -3450 3455 -3420
rect 3425 -3515 3455 -3485
rect 3425 -3585 3455 -3555
rect 3425 -3655 3455 -3625
rect 3425 -3725 3455 -3695
rect 3425 -3790 3455 -3760
rect 3425 -3850 3455 -3820
rect 3425 -3915 3455 -3885
rect 3425 -3985 3455 -3955
rect 3425 -4055 3455 -4025
rect 3425 -4125 3455 -4095
rect 3425 -4190 3455 -4160
rect 3425 -4250 3455 -4220
rect 3425 -4315 3455 -4285
rect 3425 -4385 3455 -4355
rect 3425 -4455 3455 -4425
rect 3425 -4525 3455 -4495
rect 3425 -4590 3455 -4560
rect 3775 -3050 3805 -3020
rect 3775 -3115 3805 -3085
rect 3775 -3185 3805 -3155
rect 3775 -3255 3805 -3225
rect 3775 -3325 3805 -3295
rect 3775 -3390 3805 -3360
rect 3775 -3450 3805 -3420
rect 3775 -3515 3805 -3485
rect 3775 -3585 3805 -3555
rect 3775 -3655 3805 -3625
rect 3775 -3725 3805 -3695
rect 3775 -3790 3805 -3760
rect 3775 -3850 3805 -3820
rect 3775 -3915 3805 -3885
rect 3775 -3985 3805 -3955
rect 3775 -4055 3805 -4025
rect 3775 -4125 3805 -4095
rect 3775 -4190 3805 -4160
rect 3775 -4250 3805 -4220
rect 3775 -4315 3805 -4285
rect 3775 -4385 3805 -4355
rect 3775 -4455 3805 -4425
rect 3775 -4525 3805 -4495
rect 3775 -4590 3805 -4560
rect 4125 -3050 4155 -3020
rect 4125 -3115 4155 -3085
rect 4125 -3185 4155 -3155
rect 4125 -3255 4155 -3225
rect 4125 -3325 4155 -3295
rect 4125 -3390 4155 -3360
rect 4125 -3450 4155 -3420
rect 4125 -3515 4155 -3485
rect 4125 -3585 4155 -3555
rect 4125 -3655 4155 -3625
rect 4125 -3725 4155 -3695
rect 4125 -3790 4155 -3760
rect 4125 -3850 4155 -3820
rect 4125 -3915 4155 -3885
rect 4125 -3985 4155 -3955
rect 4125 -4055 4155 -4025
rect 4125 -4125 4155 -4095
rect 4125 -4190 4155 -4160
rect 4125 -4250 4155 -4220
rect 4125 -4315 4155 -4285
rect 4125 -4385 4155 -4355
rect 4125 -4455 4155 -4425
rect 4125 -4525 4155 -4495
rect 4125 -4590 4155 -4560
rect 4475 -3050 4505 -3020
rect 4475 -3115 4505 -3085
rect 4475 -3185 4505 -3155
rect 4475 -3255 4505 -3225
rect 4475 -3325 4505 -3295
rect 4475 -3390 4505 -3360
rect 4475 -3450 4505 -3420
rect 4475 -3515 4505 -3485
rect 4475 -3585 4505 -3555
rect 4475 -3655 4505 -3625
rect 4475 -3725 4505 -3695
rect 4475 -3790 4505 -3760
rect 4475 -3850 4505 -3820
rect 4475 -3915 4505 -3885
rect 4475 -3985 4505 -3955
rect 4475 -4055 4505 -4025
rect 4475 -4125 4505 -4095
rect 4475 -4190 4505 -4160
rect 4475 -4250 4505 -4220
rect 4475 -4315 4505 -4285
rect 4475 -4385 4505 -4355
rect 4475 -4455 4505 -4425
rect 4475 -4525 4505 -4495
rect 4475 -4590 4505 -4560
rect 4825 -3050 4855 -3020
rect 4825 -3115 4855 -3085
rect 4825 -3185 4855 -3155
rect 4825 -3255 4855 -3225
rect 4825 -3325 4855 -3295
rect 4825 -3390 4855 -3360
rect 4825 -3450 4855 -3420
rect 4825 -3515 4855 -3485
rect 4825 -3585 4855 -3555
rect 4825 -3655 4855 -3625
rect 4825 -3725 4855 -3695
rect 4825 -3790 4855 -3760
rect 4825 -3850 4855 -3820
rect 4825 -3915 4855 -3885
rect 4825 -3985 4855 -3955
rect 4825 -4055 4855 -4025
rect 4825 -4125 4855 -4095
rect 4825 -4190 4855 -4160
rect 4825 -4250 4855 -4220
rect 4825 -4315 4855 -4285
rect 4825 -4385 4855 -4355
rect 4825 -4455 4855 -4425
rect 4825 -4525 4855 -4495
rect 4825 -4590 4855 -4560
rect 5175 -3050 5205 -3020
rect 5175 -3115 5205 -3085
rect 5175 -3185 5205 -3155
rect 5175 -3255 5205 -3225
rect 5175 -3325 5205 -3295
rect 5175 -3390 5205 -3360
rect 5175 -3450 5205 -3420
rect 5175 -3515 5205 -3485
rect 5175 -3585 5205 -3555
rect 5175 -3655 5205 -3625
rect 5175 -3725 5205 -3695
rect 5175 -3790 5205 -3760
rect 5175 -3850 5205 -3820
rect 5175 -3915 5205 -3885
rect 5175 -3985 5205 -3955
rect 5175 -4055 5205 -4025
rect 5175 -4125 5205 -4095
rect 5175 -4190 5205 -4160
rect 5175 -4250 5205 -4220
rect 5175 -4315 5205 -4285
rect 5175 -4385 5205 -4355
rect 5175 -4455 5205 -4425
rect 5175 -4525 5205 -4495
rect 5175 -4590 5205 -4560
rect 5875 -1350 5905 -1320
rect 5875 -1415 5905 -1385
rect 5875 -1485 5905 -1455
rect 5875 -1555 5905 -1525
rect 5875 -1625 5905 -1595
rect 5875 -1690 5905 -1660
rect 5875 -1750 5905 -1720
rect 5875 -1815 5905 -1785
rect 5875 -1885 5905 -1855
rect 5875 -1955 5905 -1925
rect 5875 -2025 5905 -1995
rect 5875 -2090 5905 -2060
rect 5875 -2150 5905 -2120
rect 5875 -2215 5905 -2185
rect 5875 -2285 5905 -2255
rect 5875 -2355 5905 -2325
rect 5875 -2425 5905 -2395
rect 5875 -2490 5905 -2460
rect 5875 -2550 5905 -2520
rect 5875 -2615 5905 -2585
rect 5875 -2685 5905 -2655
rect 5875 -2755 5905 -2725
rect 5875 -2825 5905 -2795
rect 5875 -2890 5905 -2860
rect 6225 -1350 6255 -1320
rect 6225 -1415 6255 -1385
rect 6225 -1485 6255 -1455
rect 6225 -1555 6255 -1525
rect 6225 -1625 6255 -1595
rect 6225 -1690 6255 -1660
rect 6225 -1750 6255 -1720
rect 6225 -1815 6255 -1785
rect 6225 -1885 6255 -1855
rect 6225 -1955 6255 -1925
rect 6225 -2025 6255 -1995
rect 6225 -2090 6255 -2060
rect 6225 -2150 6255 -2120
rect 6225 -2215 6255 -2185
rect 6225 -2285 6255 -2255
rect 6225 -2355 6255 -2325
rect 6225 -2425 6255 -2395
rect 6225 -2490 6255 -2460
rect 6225 -2550 6255 -2520
rect 6225 -2615 6255 -2585
rect 6225 -2685 6255 -2655
rect 6225 -2755 6255 -2725
rect 6225 -2825 6255 -2795
rect 6225 -2890 6255 -2860
rect 6575 -1350 6605 -1320
rect 6575 -1415 6605 -1385
rect 6575 -1485 6605 -1455
rect 6575 -1555 6605 -1525
rect 6575 -1625 6605 -1595
rect 6575 -1690 6605 -1660
rect 6575 -1750 6605 -1720
rect 6575 -1815 6605 -1785
rect 6575 -1885 6605 -1855
rect 6575 -1955 6605 -1925
rect 6575 -2025 6605 -1995
rect 6575 -2090 6605 -2060
rect 6575 -2150 6605 -2120
rect 6575 -2215 6605 -2185
rect 6575 -2285 6605 -2255
rect 6575 -2355 6605 -2325
rect 6575 -2425 6605 -2395
rect 6575 -2490 6605 -2460
rect 6575 -2550 6605 -2520
rect 6575 -2615 6605 -2585
rect 6575 -2685 6605 -2655
rect 6575 -2755 6605 -2725
rect 6575 -2825 6605 -2795
rect 6575 -2890 6605 -2860
rect 6925 -1350 6955 -1320
rect 6925 -1415 6955 -1385
rect 6925 -1485 6955 -1455
rect 6925 -1555 6955 -1525
rect 6925 -1625 6955 -1595
rect 6925 -1690 6955 -1660
rect 6925 -1750 6955 -1720
rect 6925 -1815 6955 -1785
rect 6925 -1885 6955 -1855
rect 6925 -1955 6955 -1925
rect 6925 -2025 6955 -1995
rect 6925 -2090 6955 -2060
rect 6925 -2150 6955 -2120
rect 6925 -2215 6955 -2185
rect 6925 -2285 6955 -2255
rect 6925 -2355 6955 -2325
rect 6925 -2425 6955 -2395
rect 6925 -2490 6955 -2460
rect 6925 -2550 6955 -2520
rect 6925 -2615 6955 -2585
rect 6925 -2685 6955 -2655
rect 6925 -2755 6955 -2725
rect 6925 -2825 6955 -2795
rect 6925 -2890 6955 -2860
rect 7275 -1350 7305 -1320
rect 7275 -1415 7305 -1385
rect 7275 -1485 7305 -1455
rect 7275 -1555 7305 -1525
rect 7275 -1625 7305 -1595
rect 7275 -1690 7305 -1660
rect 7275 -1750 7305 -1720
rect 7275 -1815 7305 -1785
rect 7275 -1885 7305 -1855
rect 7275 -1955 7305 -1925
rect 7275 -2025 7305 -1995
rect 7275 -2090 7305 -2060
rect 7275 -2150 7305 -2120
rect 7275 -2215 7305 -2185
rect 7275 -2285 7305 -2255
rect 7275 -2355 7305 -2325
rect 7275 -2425 7305 -2395
rect 7275 -2490 7305 -2460
rect 7275 -2550 7305 -2520
rect 7275 -2615 7305 -2585
rect 7275 -2685 7305 -2655
rect 7275 -2755 7305 -2725
rect 7275 -2825 7305 -2795
rect 7275 -2890 7305 -2860
rect 7625 -1350 7655 -1320
rect 7625 -1415 7655 -1385
rect 7625 -1485 7655 -1455
rect 7625 -1555 7655 -1525
rect 7625 -1625 7655 -1595
rect 7625 -1690 7655 -1660
rect 7625 -1750 7655 -1720
rect 7625 -1815 7655 -1785
rect 7625 -1885 7655 -1855
rect 7625 -1955 7655 -1925
rect 7625 -2025 7655 -1995
rect 7625 -2090 7655 -2060
rect 7625 -2150 7655 -2120
rect 7625 -2215 7655 -2185
rect 7625 -2285 7655 -2255
rect 7625 -2355 7655 -2325
rect 7625 -2425 7655 -2395
rect 7625 -2490 7655 -2460
rect 7625 -2550 7655 -2520
rect 7625 -2615 7655 -2585
rect 7625 -2685 7655 -2655
rect 7625 -2755 7655 -2725
rect 7625 -2825 7655 -2795
rect 7625 -2890 7655 -2860
rect 7975 -1350 8005 -1320
rect 7975 -1415 8005 -1385
rect 7975 -1485 8005 -1455
rect 7975 -1555 8005 -1525
rect 7975 -1625 8005 -1595
rect 7975 -1690 8005 -1660
rect 7975 -1750 8005 -1720
rect 7975 -1815 8005 -1785
rect 7975 -1885 8005 -1855
rect 7975 -1955 8005 -1925
rect 7975 -2025 8005 -1995
rect 7975 -2090 8005 -2060
rect 7975 -2150 8005 -2120
rect 7975 -2215 8005 -2185
rect 7975 -2285 8005 -2255
rect 7975 -2355 8005 -2325
rect 7975 -2425 8005 -2395
rect 7975 -2490 8005 -2460
rect 7975 -2550 8005 -2520
rect 7975 -2615 8005 -2585
rect 7975 -2685 8005 -2655
rect 7975 -2755 8005 -2725
rect 7975 -2825 8005 -2795
rect 7975 -2890 8005 -2860
rect 8325 -1350 8355 -1320
rect 8325 -1415 8355 -1385
rect 8325 -1485 8355 -1455
rect 8325 -1555 8355 -1525
rect 8325 -1625 8355 -1595
rect 8325 -1690 8355 -1660
rect 8325 -1750 8355 -1720
rect 8325 -1815 8355 -1785
rect 8325 -1885 8355 -1855
rect 8325 -1955 8355 -1925
rect 8325 -2025 8355 -1995
rect 8325 -2090 8355 -2060
rect 8325 -2150 8355 -2120
rect 8325 -2215 8355 -2185
rect 8325 -2285 8355 -2255
rect 8325 -2355 8355 -2325
rect 8325 -2425 8355 -2395
rect 8325 -2490 8355 -2460
rect 8325 -2550 8355 -2520
rect 8325 -2615 8355 -2585
rect 8325 -2685 8355 -2655
rect 8325 -2755 8355 -2725
rect 8325 -2825 8355 -2795
rect 8325 -2890 8355 -2860
rect 8675 -1350 8705 -1320
rect 8675 -1415 8705 -1385
rect 8675 -1485 8705 -1455
rect 8675 -1555 8705 -1525
rect 8675 -1625 8705 -1595
rect 8675 -1690 8705 -1660
rect 8675 -1750 8705 -1720
rect 8675 -1815 8705 -1785
rect 8675 -1885 8705 -1855
rect 8675 -1955 8705 -1925
rect 8675 -2025 8705 -1995
rect 8675 -2090 8705 -2060
rect 8675 -2150 8705 -2120
rect 8675 -2215 8705 -2185
rect 8675 -2285 8705 -2255
rect 8675 -2355 8705 -2325
rect 8675 -2425 8705 -2395
rect 8675 -2490 8705 -2460
rect 8675 -2550 8705 -2520
rect 8675 -2615 8705 -2585
rect 8675 -2685 8705 -2655
rect 8675 -2755 8705 -2725
rect 8675 -2825 8705 -2795
rect 8675 -2890 8705 -2860
rect 9025 -1350 9055 -1320
rect 9025 -1415 9055 -1385
rect 9025 -1485 9055 -1455
rect 9025 -1555 9055 -1525
rect 9025 -1625 9055 -1595
rect 9025 -1690 9055 -1660
rect 9025 -1750 9055 -1720
rect 9025 -1815 9055 -1785
rect 9025 -1885 9055 -1855
rect 9025 -1955 9055 -1925
rect 9025 -2025 9055 -1995
rect 9025 -2090 9055 -2060
rect 9025 -2150 9055 -2120
rect 9025 -2215 9055 -2185
rect 9025 -2285 9055 -2255
rect 9025 -2355 9055 -2325
rect 9025 -2425 9055 -2395
rect 9025 -2490 9055 -2460
rect 9025 -2550 9055 -2520
rect 9025 -2615 9055 -2585
rect 9025 -2685 9055 -2655
rect 9025 -2755 9055 -2725
rect 9025 -2825 9055 -2795
rect 9025 -2890 9055 -2860
rect 5525 -3050 5555 -3020
rect 5525 -3115 5555 -3085
rect 5525 -3185 5555 -3155
rect 5525 -3255 5555 -3225
rect 5525 -3325 5555 -3295
rect 5525 -3390 5555 -3360
rect 5525 -3450 5555 -3420
rect 5525 -3515 5555 -3485
rect 5525 -3585 5555 -3555
rect 5525 -3655 5555 -3625
rect 5525 -3725 5555 -3695
rect 5525 -3790 5555 -3760
rect 5525 -3850 5555 -3820
rect 5525 -3915 5555 -3885
rect 5525 -3985 5555 -3955
rect 5525 -4055 5555 -4025
rect 5525 -4125 5555 -4095
rect 5525 -4190 5555 -4160
rect 5525 -4250 5555 -4220
rect 5525 -4315 5555 -4285
rect 5525 -4385 5555 -4355
rect 5525 -4455 5555 -4425
rect 5525 -4525 5555 -4495
rect 5525 -4590 5555 -4560
<< metal2 >>
rect 2100 19310 2160 19325
rect 2100 19280 2115 19310
rect 2145 19280 2160 19310
rect 2100 19245 2160 19280
rect 2100 19215 2115 19245
rect 2145 19215 2160 19245
rect 2100 19175 2160 19215
rect 2100 19145 2115 19175
rect 2145 19145 2160 19175
rect 2100 19105 2160 19145
rect 2100 19075 2115 19105
rect 2145 19075 2160 19105
rect 2100 19035 2160 19075
rect 2100 19005 2115 19035
rect 2145 19005 2160 19035
rect 2100 18970 2160 19005
rect 2100 18940 2115 18970
rect 2145 18940 2160 18970
rect 2100 18910 2160 18940
rect 2100 18880 2115 18910
rect 2145 18880 2160 18910
rect 2100 18845 2160 18880
rect 2100 18815 2115 18845
rect 2145 18815 2160 18845
rect 2100 18775 2160 18815
rect 2100 18745 2115 18775
rect 2145 18745 2160 18775
rect 2100 18705 2160 18745
rect 2100 18675 2115 18705
rect 2145 18675 2160 18705
rect 2100 18635 2160 18675
rect 2100 18605 2115 18635
rect 2145 18605 2160 18635
rect 2100 18570 2160 18605
rect 2100 18540 2115 18570
rect 2145 18540 2160 18570
rect 2100 18510 2160 18540
rect 2100 18480 2115 18510
rect 2145 18480 2160 18510
rect 2100 18445 2160 18480
rect 2100 18415 2115 18445
rect 2145 18415 2160 18445
rect 2100 18375 2160 18415
rect 2100 18345 2115 18375
rect 2145 18345 2160 18375
rect 2100 18305 2160 18345
rect 2100 18275 2115 18305
rect 2145 18275 2160 18305
rect 2100 18235 2160 18275
rect 2100 18205 2115 18235
rect 2145 18205 2160 18235
rect 2100 18170 2160 18205
rect 2100 18140 2115 18170
rect 2145 18140 2160 18170
rect 2100 18110 2160 18140
rect 2100 18080 2115 18110
rect 2145 18080 2160 18110
rect 2100 18045 2160 18080
rect 2100 18015 2115 18045
rect 2145 18015 2160 18045
rect 2100 17975 2160 18015
rect 2100 17945 2115 17975
rect 2145 17945 2160 17975
rect 2100 17905 2160 17945
rect 2100 17875 2115 17905
rect 2145 17875 2160 17905
rect 2100 17835 2160 17875
rect 2100 17805 2115 17835
rect 2145 17805 2160 17835
rect 2100 17770 2160 17805
rect 2100 17740 2115 17770
rect 2145 17740 2160 17770
rect 2100 17725 2160 17740
rect 6690 19310 6750 19325
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2205 15925 2325 15930
rect 2205 15895 2210 15925
rect 2240 15895 2250 15925
rect 2280 15895 2290 15925
rect 2320 15920 2325 15925
rect 2320 15900 2385 15920
rect 2320 15895 2325 15900
rect 2205 15890 2325 15895
rect 2070 15690 2970 15695
rect 2070 15660 2075 15690
rect 2105 15660 2115 15690
rect 2145 15660 2155 15690
rect 2185 15660 2970 15690
rect 2070 15650 2970 15660
rect 2070 15620 2075 15650
rect 2105 15620 2115 15650
rect 2145 15620 2155 15650
rect 2185 15620 2970 15650
rect 2070 15610 2970 15620
rect 2070 15580 2075 15610
rect 2105 15580 2115 15610
rect 2145 15580 2155 15610
rect 2185 15580 2970 15610
rect 2070 15575 2970 15580
rect 6650 15595 6780 15600
rect 6650 15565 6665 15595
rect 6695 15565 6705 15595
rect 6735 15565 6745 15595
rect 6775 15565 6780 15595
rect 6650 15555 6780 15565
rect 6650 15525 6665 15555
rect 6695 15525 6705 15555
rect 6735 15525 6745 15555
rect 6775 15525 6780 15555
rect 6650 15515 6780 15525
rect 6650 15485 6665 15515
rect 6695 15485 6705 15515
rect 6735 15485 6745 15515
rect 6775 15485 6780 15515
rect 6650 15480 6780 15485
rect 5690 12925 6780 12930
rect 5690 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6745 12925
rect 6775 12895 6780 12925
rect 5690 12885 6780 12895
rect 5690 12855 6665 12885
rect 6695 12855 6705 12885
rect 6735 12855 6745 12885
rect 6775 12855 6780 12885
rect 5690 12845 6780 12855
rect 5690 12815 6665 12845
rect 6695 12815 6705 12845
rect 6735 12815 6745 12845
rect 6775 12815 6780 12845
rect 5690 12810 6780 12815
rect 2070 12710 3355 12715
rect 2070 12680 2075 12710
rect 2105 12680 2115 12710
rect 2145 12680 2155 12710
rect 2185 12680 3355 12710
rect 2070 12670 3355 12680
rect 2070 12640 2075 12670
rect 2105 12640 2115 12670
rect 2145 12640 2155 12670
rect 2185 12640 3355 12670
rect 2070 12635 3355 12640
rect 2070 12550 3800 12555
rect 2070 12520 2075 12550
rect 2105 12520 2115 12550
rect 2145 12520 2155 12550
rect 2185 12520 3800 12550
rect 2070 12510 3800 12520
rect 2070 12480 2075 12510
rect 2105 12480 2115 12510
rect 2145 12480 2155 12510
rect 2185 12480 3800 12510
rect 2070 12470 3800 12480
rect 2070 12440 2075 12470
rect 2105 12440 2115 12470
rect 2145 12440 2155 12470
rect 2185 12440 3800 12470
rect 2070 12435 3800 12440
rect 5670 12150 6780 12155
rect 5670 12120 6665 12150
rect 6695 12120 6705 12150
rect 6735 12120 6745 12150
rect 6775 12120 6780 12150
rect 5670 12110 6780 12120
rect 5670 12080 6665 12110
rect 6695 12080 6705 12110
rect 6735 12080 6745 12110
rect 6775 12080 6780 12110
rect 5670 12070 6780 12080
rect 5670 12040 6665 12070
rect 6695 12040 6705 12070
rect 6735 12040 6745 12070
rect 6775 12040 6780 12070
rect 5670 12035 6780 12040
rect 5870 11165 6780 11170
rect 5870 11135 6665 11165
rect 6695 11135 6705 11165
rect 6735 11135 6745 11165
rect 6775 11135 6780 11165
rect 5870 11125 6780 11135
rect 5870 11095 6665 11125
rect 6695 11095 6705 11125
rect 6735 11095 6745 11125
rect 6775 11095 6780 11125
rect 5870 11085 6780 11095
rect 5870 11055 6665 11085
rect 6695 11055 6705 11085
rect 6735 11055 6745 11085
rect 6775 11055 6780 11085
rect 5870 11050 6780 11055
rect 5855 10440 6780 10445
rect 5855 10410 6665 10440
rect 6695 10410 6705 10440
rect 6735 10410 6745 10440
rect 6775 10410 6780 10440
rect 5855 10400 6780 10410
rect 5855 10370 6665 10400
rect 6695 10370 6705 10400
rect 6735 10370 6745 10400
rect 6775 10370 6780 10400
rect 5855 10360 6780 10370
rect 5855 10330 6665 10360
rect 6695 10330 6705 10360
rect 6735 10330 6745 10360
rect 6775 10330 6780 10360
rect 5855 10325 6780 10330
rect 5925 10080 6780 10085
rect 5925 10050 6665 10080
rect 6695 10050 6705 10080
rect 6735 10050 6745 10080
rect 6775 10050 6780 10080
rect 5925 10040 6780 10050
rect 5925 10010 6665 10040
rect 6695 10010 6705 10040
rect 6735 10010 6745 10040
rect 6775 10010 6780 10040
rect 5925 10000 6780 10010
rect 5925 9970 6665 10000
rect 6695 9970 6705 10000
rect 6735 9970 6745 10000
rect 6775 9970 6780 10000
rect 5925 9965 6780 9970
rect 1310 9635 1370 9650
rect 1310 9605 1325 9635
rect 1355 9605 1370 9635
rect 1310 9570 1370 9605
rect 1310 9540 1325 9570
rect 1355 9540 1370 9570
rect 1310 9500 1370 9540
rect 1310 9470 1325 9500
rect 1355 9470 1370 9500
rect 1310 9430 1370 9470
rect 1310 9400 1325 9430
rect 1355 9400 1370 9430
rect 1310 9360 1370 9400
rect 1310 9330 1325 9360
rect 1355 9330 1370 9360
rect 1310 9295 1370 9330
rect 1310 9265 1325 9295
rect 1355 9265 1370 9295
rect 1310 9235 1370 9265
rect 1310 9205 1325 9235
rect 1355 9205 1370 9235
rect 1310 9170 1370 9205
rect 1310 9140 1325 9170
rect 1355 9140 1370 9170
rect 1310 9100 1370 9140
rect 1310 9070 1325 9100
rect 1355 9070 1370 9100
rect 1310 9030 1370 9070
rect 1310 9000 1325 9030
rect 1355 9000 1370 9030
rect 1310 8960 1370 9000
rect 1310 8930 1325 8960
rect 1355 8930 1370 8960
rect 1310 8895 1370 8930
rect 1310 8865 1325 8895
rect 1355 8865 1370 8895
rect 1310 8835 1370 8865
rect 1310 8805 1325 8835
rect 1355 8805 1370 8835
rect 1310 8770 1370 8805
rect 1310 8740 1325 8770
rect 1355 8740 1370 8770
rect 1310 8700 1370 8740
rect 1310 8670 1325 8700
rect 1355 8670 1370 8700
rect 1310 8630 1370 8670
rect 1310 8600 1325 8630
rect 1355 8600 1370 8630
rect 1310 8560 1370 8600
rect 1310 8530 1325 8560
rect 1355 8530 1370 8560
rect 1310 8495 1370 8530
rect 1310 8465 1325 8495
rect 1355 8465 1370 8495
rect 1310 8435 1370 8465
rect 1310 8405 1325 8435
rect 1355 8405 1370 8435
rect 1310 8370 1370 8405
rect 1310 8340 1325 8370
rect 1355 8340 1370 8370
rect 1310 8300 1370 8340
rect 1310 8270 1325 8300
rect 1355 8270 1370 8300
rect 1310 8230 1370 8270
rect 1310 8200 1325 8230
rect 1355 8200 1370 8230
rect 1310 8160 1370 8200
rect 1310 8130 1325 8160
rect 1355 8130 1370 8160
rect 1310 8105 1370 8130
rect 2235 9635 2295 9650
rect 2235 9605 2250 9635
rect 2280 9605 2295 9635
rect 2235 9570 2295 9605
rect 2235 9540 2250 9570
rect 2280 9540 2295 9570
rect 2235 9500 2295 9540
rect 2235 9470 2250 9500
rect 2280 9470 2295 9500
rect 2235 9430 2295 9470
rect 2235 9400 2250 9430
rect 2280 9400 2295 9430
rect 2235 9360 2295 9400
rect 2235 9330 2250 9360
rect 2280 9330 2295 9360
rect 2235 9295 2295 9330
rect 2235 9265 2250 9295
rect 2280 9265 2295 9295
rect 2235 9235 2295 9265
rect 2235 9205 2250 9235
rect 2280 9205 2295 9235
rect 2235 9170 2295 9205
rect 2235 9140 2250 9170
rect 2280 9140 2295 9170
rect 2235 9100 2295 9140
rect 2235 9070 2250 9100
rect 2280 9070 2295 9100
rect 2235 9030 2295 9070
rect 2235 9000 2250 9030
rect 2280 9000 2295 9030
rect 2235 8960 2295 9000
rect 2235 8930 2250 8960
rect 2280 8930 2295 8960
rect 2235 8895 2295 8930
rect 2235 8865 2250 8895
rect 2280 8865 2295 8895
rect 2235 8835 2295 8865
rect 2235 8805 2250 8835
rect 2280 8805 2295 8835
rect 2235 8770 2295 8805
rect 2235 8740 2250 8770
rect 2280 8740 2295 8770
rect 2235 8700 2295 8740
rect 2235 8670 2250 8700
rect 2280 8670 2295 8700
rect 2235 8630 2295 8670
rect 2235 8600 2250 8630
rect 2280 8600 2295 8630
rect 2235 8560 2295 8600
rect 2235 8530 2250 8560
rect 2280 8530 2295 8560
rect 2235 8495 2295 8530
rect 2235 8465 2250 8495
rect 2280 8465 2295 8495
rect 2235 8435 2295 8465
rect 2235 8405 2250 8435
rect 2280 8405 2295 8435
rect 2235 8370 2295 8405
rect 2235 8340 2250 8370
rect 2280 8340 2295 8370
rect 2235 8300 2295 8340
rect 2235 8270 2250 8300
rect 2280 8270 2295 8300
rect 2235 8230 2295 8270
rect 2235 8200 2250 8230
rect 2280 8200 2295 8230
rect 2235 8160 2295 8200
rect 2235 8130 2250 8160
rect 2280 8130 2295 8160
rect 2235 8105 2295 8130
rect 6690 9635 6750 9650
rect 6690 9605 6705 9635
rect 6735 9605 6750 9635
rect 6690 9570 6750 9605
rect 6690 9540 6705 9570
rect 6735 9540 6750 9570
rect 6690 9500 6750 9540
rect 6690 9470 6705 9500
rect 6735 9470 6750 9500
rect 6690 9430 6750 9470
rect 6690 9400 6705 9430
rect 6735 9400 6750 9430
rect 6690 9360 6750 9400
rect 6690 9330 6705 9360
rect 6735 9330 6750 9360
rect 6690 9295 6750 9330
rect 6690 9265 6705 9295
rect 6735 9265 6750 9295
rect 6690 9235 6750 9265
rect 6690 9205 6705 9235
rect 6735 9205 6750 9235
rect 6690 9170 6750 9205
rect 6690 9140 6705 9170
rect 6735 9140 6750 9170
rect 6690 9100 6750 9140
rect 6690 9070 6705 9100
rect 6735 9070 6750 9100
rect 6690 9030 6750 9070
rect 6690 9000 6705 9030
rect 6735 9000 6750 9030
rect 6690 8960 6750 9000
rect 6690 8930 6705 8960
rect 6735 8930 6750 8960
rect 6690 8895 6750 8930
rect 6690 8865 6705 8895
rect 6735 8865 6750 8895
rect 6690 8835 6750 8865
rect 6690 8805 6705 8835
rect 6735 8805 6750 8835
rect 6690 8770 6750 8805
rect 6690 8740 6705 8770
rect 6735 8740 6750 8770
rect 6690 8700 6750 8740
rect 6690 8670 6705 8700
rect 6735 8670 6750 8700
rect 6690 8630 6750 8670
rect 6690 8600 6705 8630
rect 6735 8600 6750 8630
rect 6690 8560 6750 8600
rect 6690 8530 6705 8560
rect 6735 8530 6750 8560
rect 6690 8495 6750 8530
rect 6690 8465 6705 8495
rect 6735 8465 6750 8495
rect 6690 8435 6750 8465
rect 6690 8405 6705 8435
rect 6735 8405 6750 8435
rect 6690 8370 6750 8405
rect 6690 8340 6705 8370
rect 6735 8340 6750 8370
rect 6690 8300 6750 8340
rect 6690 8270 6705 8300
rect 6735 8270 6750 8300
rect 6690 8230 6750 8270
rect 6690 8200 6705 8230
rect 6735 8200 6750 8230
rect 6690 8160 6750 8200
rect 6690 8130 6705 8160
rect 6735 8130 6750 8160
rect 6690 8105 6750 8130
rect 7610 9635 7670 9650
rect 7610 9605 7625 9635
rect 7655 9605 7670 9635
rect 7610 9570 7670 9605
rect 7610 9540 7625 9570
rect 7655 9540 7670 9570
rect 7610 9500 7670 9540
rect 7610 9470 7625 9500
rect 7655 9470 7670 9500
rect 7610 9430 7670 9470
rect 7610 9400 7625 9430
rect 7655 9400 7670 9430
rect 7610 9360 7670 9400
rect 7610 9330 7625 9360
rect 7655 9330 7670 9360
rect 7610 9295 7670 9330
rect 7610 9265 7625 9295
rect 7655 9265 7670 9295
rect 7610 9235 7670 9265
rect 7610 9205 7625 9235
rect 7655 9205 7670 9235
rect 7610 9170 7670 9205
rect 7610 9140 7625 9170
rect 7655 9140 7670 9170
rect 7610 9100 7670 9140
rect 7610 9070 7625 9100
rect 7655 9070 7670 9100
rect 7610 9030 7670 9070
rect 7610 9000 7625 9030
rect 7655 9000 7670 9030
rect 7610 8960 7670 9000
rect 7610 8930 7625 8960
rect 7655 8930 7670 8960
rect 7610 8895 7670 8930
rect 7610 8865 7625 8895
rect 7655 8865 7670 8895
rect 7610 8835 7670 8865
rect 7610 8805 7625 8835
rect 7655 8805 7670 8835
rect 7610 8770 7670 8805
rect 7610 8740 7625 8770
rect 7655 8740 7670 8770
rect 7610 8700 7670 8740
rect 7610 8670 7625 8700
rect 7655 8670 7670 8700
rect 7610 8630 7670 8670
rect 7610 8600 7625 8630
rect 7655 8600 7670 8630
rect 7610 8560 7670 8600
rect 7610 8530 7625 8560
rect 7655 8530 7670 8560
rect 7610 8495 7670 8530
rect 7610 8465 7625 8495
rect 7655 8465 7670 8495
rect 7610 8435 7670 8465
rect 7610 8405 7625 8435
rect 7655 8405 7670 8435
rect 7610 8370 7670 8405
rect 7610 8340 7625 8370
rect 7655 8340 7670 8370
rect 7610 8300 7670 8340
rect 7610 8270 7625 8300
rect 7655 8270 7670 8300
rect 7610 8230 7670 8270
rect 7610 8200 7625 8230
rect 7655 8200 7670 8230
rect 7610 8160 7670 8200
rect 7610 8130 7625 8160
rect 7655 8130 7670 8160
rect 7610 8105 7670 8130
rect 1980 8085 2515 8090
rect 1980 8055 1985 8085
rect 2015 8055 2025 8085
rect 2055 8055 2065 8085
rect 2095 8055 2480 8085
rect 2510 8055 2515 8085
rect 1980 8050 2515 8055
rect 6465 8070 7000 8075
rect 6465 8040 6470 8070
rect 6500 8040 6885 8070
rect 6915 8040 6925 8070
rect 6955 8040 6965 8070
rect 6995 8040 7000 8070
rect 6465 8035 7000 8040
rect 1630 8030 3890 8035
rect 1630 8000 1635 8030
rect 1665 8000 1675 8030
rect 1705 8000 1715 8030
rect 1745 8000 3635 8030
rect 3665 8000 3855 8030
rect 3885 8000 3890 8030
rect 1630 7995 3890 8000
rect 5310 8015 7350 8020
rect 5310 7985 5315 8015
rect 5345 7985 7235 8015
rect 7265 7985 7275 8015
rect 7305 7985 7315 8015
rect 7345 7985 7350 8015
rect 5310 7980 7350 7985
rect 3165 7955 3280 7980
rect 3165 7925 3180 7955
rect 3210 7925 3240 7955
rect 3270 7925 3280 7955
rect 3165 7885 3280 7925
rect 3165 7855 3180 7885
rect 3210 7855 3240 7885
rect 3270 7855 3280 7885
rect 3165 7815 3280 7855
rect 3165 7785 3180 7815
rect 3210 7785 3240 7815
rect 3270 7785 3280 7815
rect 3165 7745 3280 7785
rect 3165 7715 3180 7745
rect 3210 7715 3240 7745
rect 3270 7715 3280 7745
rect 3165 7680 3280 7715
rect 3165 7650 3180 7680
rect 3210 7650 3240 7680
rect 3270 7650 3280 7680
rect 3165 7620 3280 7650
rect 3165 7590 3180 7620
rect 3210 7590 3240 7620
rect 3270 7590 3280 7620
rect 3165 7555 3280 7590
rect 3165 7525 3180 7555
rect 3210 7525 3240 7555
rect 3270 7525 3280 7555
rect 3165 7485 3280 7525
rect 3165 7455 3180 7485
rect 3210 7455 3240 7485
rect 3270 7455 3280 7485
rect 3165 7415 3280 7455
rect 3165 7385 3180 7415
rect 3210 7385 3240 7415
rect 3270 7385 3280 7415
rect 3165 7345 3280 7385
rect 3165 7315 3180 7345
rect 3210 7315 3240 7345
rect 3270 7315 3280 7345
rect 3165 7280 3280 7315
rect 3165 7250 3180 7280
rect 3210 7250 3240 7280
rect 3270 7250 3280 7280
rect 3165 7220 3280 7250
rect 3165 7190 3180 7220
rect 3210 7190 3240 7220
rect 3270 7190 3280 7220
rect 3165 7155 3280 7190
rect 3165 7125 3180 7155
rect 3210 7125 3240 7155
rect 3270 7125 3280 7155
rect 3165 7085 3280 7125
rect 3165 7055 3180 7085
rect 3210 7055 3240 7085
rect 3270 7055 3280 7085
rect 3165 7015 3280 7055
rect 3165 6985 3180 7015
rect 3210 6985 3240 7015
rect 3270 6985 3280 7015
rect 3165 6945 3280 6985
rect 3165 6915 3180 6945
rect 3210 6915 3240 6945
rect 3270 6915 3280 6945
rect 3165 6880 3280 6915
rect 3165 6850 3180 6880
rect 3210 6850 3240 6880
rect 3270 6850 3280 6880
rect 3165 6820 3280 6850
rect 3165 6790 3180 6820
rect 3210 6790 3240 6820
rect 3270 6790 3280 6820
rect 3165 6755 3280 6790
rect 3165 6725 3180 6755
rect 3210 6725 3240 6755
rect 3270 6725 3280 6755
rect 3165 6685 3280 6725
rect 3165 6655 3180 6685
rect 3210 6655 3240 6685
rect 3270 6655 3280 6685
rect 3165 6615 3280 6655
rect 3165 6585 3180 6615
rect 3210 6585 3240 6615
rect 3270 6585 3280 6615
rect 3165 6545 3280 6585
rect 3165 6515 3180 6545
rect 3210 6515 3240 6545
rect 3270 6515 3280 6545
rect 3165 6480 3280 6515
rect 3165 6450 3180 6480
rect 3210 6450 3240 6480
rect 3270 6450 3280 6480
rect 3165 6435 3280 6450
rect 3340 7955 3390 7980
rect 3340 7925 3350 7955
rect 3380 7925 3390 7955
rect 3340 7885 3390 7925
rect 3340 7855 3350 7885
rect 3380 7855 3390 7885
rect 3340 7815 3390 7855
rect 3340 7785 3350 7815
rect 3380 7785 3390 7815
rect 3340 7745 3390 7785
rect 3340 7715 3350 7745
rect 3380 7715 3390 7745
rect 3340 7680 3390 7715
rect 3340 7650 3350 7680
rect 3380 7650 3390 7680
rect 3340 7620 3390 7650
rect 3340 7590 3350 7620
rect 3380 7590 3390 7620
rect 3340 7555 3390 7590
rect 3340 7525 3350 7555
rect 3380 7525 3390 7555
rect 3340 7485 3390 7525
rect 3340 7455 3350 7485
rect 3380 7455 3390 7485
rect 3340 7415 3390 7455
rect 3340 7385 3350 7415
rect 3380 7385 3390 7415
rect 3340 7345 3390 7385
rect 3340 7315 3350 7345
rect 3380 7315 3390 7345
rect 3340 7280 3390 7315
rect 3340 7250 3350 7280
rect 3380 7250 3390 7280
rect 3340 7220 3390 7250
rect 3340 7190 3350 7220
rect 3380 7190 3390 7220
rect 3340 7155 3390 7190
rect 3340 7125 3350 7155
rect 3380 7125 3390 7155
rect 3340 7085 3390 7125
rect 3340 7055 3350 7085
rect 3380 7055 3390 7085
rect 3340 7015 3390 7055
rect 3340 6985 3350 7015
rect 3380 6985 3390 7015
rect 3340 6945 3390 6985
rect 3340 6915 3350 6945
rect 3380 6915 3390 6945
rect 3340 6880 3390 6915
rect 3340 6850 3350 6880
rect 3380 6850 3390 6880
rect 3340 6820 3390 6850
rect 3340 6790 3350 6820
rect 3380 6790 3390 6820
rect 3340 6755 3390 6790
rect 3340 6725 3350 6755
rect 3380 6725 3390 6755
rect 3340 6685 3390 6725
rect 3340 6655 3350 6685
rect 3380 6655 3390 6685
rect 3340 6615 3390 6655
rect 3340 6585 3350 6615
rect 3380 6585 3390 6615
rect 3340 6545 3390 6585
rect 3340 6515 3350 6545
rect 3380 6515 3390 6545
rect 3340 6480 3390 6515
rect 3340 6450 3350 6480
rect 3380 6450 3390 6480
rect 3340 6435 3390 6450
rect 2845 6415 2885 6420
rect 2845 6385 2850 6415
rect 2880 6410 2885 6415
rect 3380 6415 3420 6420
rect 3380 6410 3385 6415
rect 2880 6390 3385 6410
rect 2880 6385 2885 6390
rect 2845 6380 2885 6385
rect 3380 6385 3385 6390
rect 3415 6385 3420 6415
rect 3380 6380 3420 6385
rect 5470 6415 5510 6420
rect 5470 6385 5475 6415
rect 5505 6410 5510 6415
rect 6145 6415 6185 6420
rect 6145 6410 6150 6415
rect 5505 6390 6150 6410
rect 5505 6385 5510 6390
rect 5470 6380 5510 6385
rect 6145 6385 6150 6390
rect 6180 6385 6185 6415
rect 6145 6380 6185 6385
rect 2715 6305 2755 6310
rect 2715 6275 2720 6305
rect 2750 6300 2755 6305
rect 3075 6305 3115 6310
rect 3075 6300 3080 6305
rect 2750 6280 3080 6300
rect 2750 6275 2755 6280
rect 2715 6270 2755 6275
rect 3075 6275 3080 6280
rect 3110 6275 3115 6305
rect 3075 6270 3115 6275
rect 3290 6300 4510 6305
rect 3290 6270 3295 6300
rect 3325 6270 4475 6300
rect 4505 6270 4510 6300
rect 3290 6265 4510 6270
rect 3435 6245 5585 6250
rect 3435 6215 3440 6245
rect 3470 6215 4475 6245
rect 4505 6215 5550 6245
rect 5580 6215 5585 6245
rect 3435 6210 5585 6215
rect 930 6190 8050 6195
rect 930 6160 935 6190
rect 965 6160 975 6190
rect 1005 6160 1015 6190
rect 1045 6160 4310 6190
rect 4340 6160 4420 6190
rect 4450 6160 4530 6190
rect 4560 6160 4640 6190
rect 4670 6160 7935 6190
rect 7965 6160 7975 6190
rect 8005 6160 8015 6190
rect 8045 6160 8050 6190
rect 930 6150 8050 6160
rect 930 6120 935 6150
rect 965 6120 975 6150
rect 1005 6120 1015 6150
rect 1045 6120 4310 6150
rect 4340 6120 4420 6150
rect 4450 6120 4530 6150
rect 4560 6120 4640 6150
rect 4670 6120 7935 6150
rect 7965 6120 7975 6150
rect 8005 6120 8015 6150
rect 8045 6120 8050 6150
rect 930 6110 8050 6120
rect 930 6080 935 6110
rect 965 6080 975 6110
rect 1005 6080 1015 6110
rect 1045 6080 4310 6110
rect 4340 6080 4420 6110
rect 4450 6080 4530 6110
rect 4560 6080 4640 6110
rect 4670 6080 7935 6110
rect 7965 6080 7975 6110
rect 8005 6080 8015 6110
rect 8045 6080 8050 6110
rect 930 6075 8050 6080
rect 5870 5420 6260 5425
rect 5870 5390 5875 5420
rect 5905 5390 6225 5420
rect 6255 5390 6260 5420
rect 5870 5385 6260 5390
rect 3075 5075 3115 5080
rect 3075 5045 3080 5075
rect 3110 5045 3115 5075
rect 3075 5040 3115 5045
rect 5620 5020 5910 5025
rect 5620 4990 5625 5020
rect 5655 4990 5875 5020
rect 5905 4990 5910 5020
rect 5620 4985 5910 4990
rect 5620 4425 5660 4430
rect 5620 4395 5625 4425
rect 5655 4395 5660 4425
rect 5620 4390 5660 4395
rect 5475 3850 5505 3855
rect 4720 3825 5475 3845
rect 5475 3815 5505 3820
rect 3380 3790 3420 3795
rect 3380 3760 3385 3790
rect 3415 3785 3420 3790
rect 3415 3765 3955 3785
rect 3415 3760 3420 3765
rect 3380 3755 3420 3760
rect 3435 3110 5585 3115
rect 3435 3080 3440 3110
rect 3470 3080 4475 3110
rect 4505 3080 5550 3110
rect 5580 3080 5585 3110
rect 3435 3075 5585 3080
rect 4470 2890 4510 2895
rect 4470 2860 4475 2890
rect 4505 2860 4510 2890
rect 4470 2855 4510 2860
rect 2045 2295 2085 2305
rect 2120 2295 2160 2305
rect 2045 2275 2160 2295
rect 2045 2265 2085 2275
rect 2120 2265 2160 2275
rect 2000 2240 2040 2250
rect 2075 2240 2115 2250
rect 2000 2220 2115 2240
rect 2000 2210 2040 2220
rect 2075 2210 2115 2220
rect 3605 1580 3625 1600
rect 5355 1580 5375 1600
rect 930 1145 8050 1150
rect 930 1115 935 1145
rect 965 1115 975 1145
rect 1005 1115 1015 1145
rect 1045 1115 4420 1145
rect 4450 1115 4530 1145
rect 4560 1115 7935 1145
rect 7965 1115 7975 1145
rect 8005 1115 8015 1145
rect 8045 1115 8050 1145
rect 930 1105 8050 1115
rect 930 1075 935 1105
rect 965 1075 975 1105
rect 1005 1075 1015 1105
rect 1045 1075 4420 1105
rect 4450 1075 4530 1105
rect 4560 1075 7935 1105
rect 7965 1075 7975 1105
rect 8005 1075 8015 1105
rect 8045 1075 8050 1105
rect 930 1065 8050 1075
rect 930 1035 935 1065
rect 965 1035 975 1065
rect 1005 1035 1015 1065
rect 1045 1035 4420 1065
rect 4450 1035 4530 1065
rect 4560 1035 7935 1065
rect 7965 1035 7975 1065
rect 8005 1035 8015 1065
rect 8045 1035 8050 1065
rect 930 1030 8050 1035
rect 2175 840 2195 860
rect 6785 840 6805 860
rect -90 -1320 -30 -1305
rect -90 -1350 -75 -1320
rect -45 -1350 -30 -1320
rect -90 -1385 -30 -1350
rect -90 -1415 -75 -1385
rect -45 -1415 -30 -1385
rect -90 -1455 -30 -1415
rect -90 -1485 -75 -1455
rect -45 -1485 -30 -1455
rect -90 -1525 -30 -1485
rect -90 -1555 -75 -1525
rect -45 -1555 -30 -1525
rect -90 -1595 -30 -1555
rect -90 -1625 -75 -1595
rect -45 -1625 -30 -1595
rect -90 -1660 -30 -1625
rect -90 -1690 -75 -1660
rect -45 -1690 -30 -1660
rect -90 -1720 -30 -1690
rect -90 -1750 -75 -1720
rect -45 -1750 -30 -1720
rect -90 -1785 -30 -1750
rect -90 -1815 -75 -1785
rect -45 -1815 -30 -1785
rect -90 -1855 -30 -1815
rect -90 -1885 -75 -1855
rect -45 -1885 -30 -1855
rect -90 -1925 -30 -1885
rect -90 -1955 -75 -1925
rect -45 -1955 -30 -1925
rect -90 -1995 -30 -1955
rect -90 -2025 -75 -1995
rect -45 -2025 -30 -1995
rect -90 -2060 -30 -2025
rect -90 -2090 -75 -2060
rect -45 -2090 -30 -2060
rect -90 -2120 -30 -2090
rect -90 -2150 -75 -2120
rect -45 -2150 -30 -2120
rect -90 -2185 -30 -2150
rect -90 -2215 -75 -2185
rect -45 -2215 -30 -2185
rect -90 -2255 -30 -2215
rect -90 -2285 -75 -2255
rect -45 -2285 -30 -2255
rect -90 -2325 -30 -2285
rect -90 -2355 -75 -2325
rect -45 -2355 -30 -2325
rect -90 -2395 -30 -2355
rect -90 -2425 -75 -2395
rect -45 -2425 -30 -2395
rect -90 -2460 -30 -2425
rect -90 -2490 -75 -2460
rect -45 -2490 -30 -2460
rect -90 -2520 -30 -2490
rect -90 -2550 -75 -2520
rect -45 -2550 -30 -2520
rect -90 -2585 -30 -2550
rect -90 -2615 -75 -2585
rect -45 -2615 -30 -2585
rect -90 -2655 -30 -2615
rect -90 -2685 -75 -2655
rect -45 -2685 -30 -2655
rect -90 -2725 -30 -2685
rect -90 -2755 -75 -2725
rect -45 -2755 -30 -2725
rect -90 -2795 -30 -2755
rect -90 -2825 -75 -2795
rect -45 -2825 -30 -2795
rect -90 -2860 -30 -2825
rect -90 -2890 -75 -2860
rect -45 -2890 -30 -2860
rect -90 -2905 -30 -2890
rect 260 -1320 320 -1305
rect 260 -1350 275 -1320
rect 305 -1350 320 -1320
rect 260 -1385 320 -1350
rect 260 -1415 275 -1385
rect 305 -1415 320 -1385
rect 260 -1455 320 -1415
rect 260 -1485 275 -1455
rect 305 -1485 320 -1455
rect 260 -1525 320 -1485
rect 260 -1555 275 -1525
rect 305 -1555 320 -1525
rect 260 -1595 320 -1555
rect 260 -1625 275 -1595
rect 305 -1625 320 -1595
rect 260 -1660 320 -1625
rect 260 -1690 275 -1660
rect 305 -1690 320 -1660
rect 260 -1720 320 -1690
rect 260 -1750 275 -1720
rect 305 -1750 320 -1720
rect 260 -1785 320 -1750
rect 260 -1815 275 -1785
rect 305 -1815 320 -1785
rect 260 -1855 320 -1815
rect 260 -1885 275 -1855
rect 305 -1885 320 -1855
rect 260 -1925 320 -1885
rect 260 -1955 275 -1925
rect 305 -1955 320 -1925
rect 260 -1995 320 -1955
rect 260 -2025 275 -1995
rect 305 -2025 320 -1995
rect 260 -2060 320 -2025
rect 260 -2090 275 -2060
rect 305 -2090 320 -2060
rect 260 -2120 320 -2090
rect 260 -2150 275 -2120
rect 305 -2150 320 -2120
rect 260 -2185 320 -2150
rect 260 -2215 275 -2185
rect 305 -2215 320 -2185
rect 260 -2255 320 -2215
rect 260 -2285 275 -2255
rect 305 -2285 320 -2255
rect 260 -2325 320 -2285
rect 260 -2355 275 -2325
rect 305 -2355 320 -2325
rect 260 -2395 320 -2355
rect 260 -2425 275 -2395
rect 305 -2425 320 -2395
rect 260 -2460 320 -2425
rect 260 -2490 275 -2460
rect 305 -2490 320 -2460
rect 260 -2520 320 -2490
rect 260 -2550 275 -2520
rect 305 -2550 320 -2520
rect 260 -2585 320 -2550
rect 260 -2615 275 -2585
rect 305 -2615 320 -2585
rect 260 -2655 320 -2615
rect 260 -2685 275 -2655
rect 305 -2685 320 -2655
rect 260 -2725 320 -2685
rect 260 -2755 275 -2725
rect 305 -2755 320 -2725
rect 260 -2795 320 -2755
rect 260 -2825 275 -2795
rect 305 -2825 320 -2795
rect 260 -2860 320 -2825
rect 260 -2890 275 -2860
rect 305 -2890 320 -2860
rect 260 -2905 320 -2890
rect 610 -1320 670 -1305
rect 610 -1350 625 -1320
rect 655 -1350 670 -1320
rect 610 -1385 670 -1350
rect 610 -1415 625 -1385
rect 655 -1415 670 -1385
rect 610 -1455 670 -1415
rect 610 -1485 625 -1455
rect 655 -1485 670 -1455
rect 610 -1525 670 -1485
rect 610 -1555 625 -1525
rect 655 -1555 670 -1525
rect 610 -1595 670 -1555
rect 610 -1625 625 -1595
rect 655 -1625 670 -1595
rect 610 -1660 670 -1625
rect 610 -1690 625 -1660
rect 655 -1690 670 -1660
rect 610 -1720 670 -1690
rect 610 -1750 625 -1720
rect 655 -1750 670 -1720
rect 610 -1785 670 -1750
rect 610 -1815 625 -1785
rect 655 -1815 670 -1785
rect 610 -1855 670 -1815
rect 610 -1885 625 -1855
rect 655 -1885 670 -1855
rect 610 -1925 670 -1885
rect 610 -1955 625 -1925
rect 655 -1955 670 -1925
rect 610 -1995 670 -1955
rect 610 -2025 625 -1995
rect 655 -2025 670 -1995
rect 610 -2060 670 -2025
rect 610 -2090 625 -2060
rect 655 -2090 670 -2060
rect 610 -2120 670 -2090
rect 610 -2150 625 -2120
rect 655 -2150 670 -2120
rect 610 -2185 670 -2150
rect 610 -2215 625 -2185
rect 655 -2215 670 -2185
rect 610 -2255 670 -2215
rect 610 -2285 625 -2255
rect 655 -2285 670 -2255
rect 610 -2325 670 -2285
rect 610 -2355 625 -2325
rect 655 -2355 670 -2325
rect 610 -2395 670 -2355
rect 610 -2425 625 -2395
rect 655 -2425 670 -2395
rect 610 -2460 670 -2425
rect 610 -2490 625 -2460
rect 655 -2490 670 -2460
rect 610 -2520 670 -2490
rect 610 -2550 625 -2520
rect 655 -2550 670 -2520
rect 610 -2585 670 -2550
rect 610 -2615 625 -2585
rect 655 -2615 670 -2585
rect 610 -2655 670 -2615
rect 610 -2685 625 -2655
rect 655 -2685 670 -2655
rect 610 -2725 670 -2685
rect 610 -2755 625 -2725
rect 655 -2755 670 -2725
rect 610 -2795 670 -2755
rect 610 -2825 625 -2795
rect 655 -2825 670 -2795
rect 610 -2860 670 -2825
rect 610 -2890 625 -2860
rect 655 -2890 670 -2860
rect 610 -2905 670 -2890
rect 960 -1320 1020 -1305
rect 960 -1350 975 -1320
rect 1005 -1350 1020 -1320
rect 960 -1385 1020 -1350
rect 960 -1415 975 -1385
rect 1005 -1415 1020 -1385
rect 960 -1455 1020 -1415
rect 960 -1485 975 -1455
rect 1005 -1485 1020 -1455
rect 960 -1525 1020 -1485
rect 960 -1555 975 -1525
rect 1005 -1555 1020 -1525
rect 960 -1595 1020 -1555
rect 960 -1625 975 -1595
rect 1005 -1625 1020 -1595
rect 960 -1660 1020 -1625
rect 960 -1690 975 -1660
rect 1005 -1690 1020 -1660
rect 960 -1720 1020 -1690
rect 960 -1750 975 -1720
rect 1005 -1750 1020 -1720
rect 960 -1785 1020 -1750
rect 960 -1815 975 -1785
rect 1005 -1815 1020 -1785
rect 960 -1855 1020 -1815
rect 960 -1885 975 -1855
rect 1005 -1885 1020 -1855
rect 960 -1925 1020 -1885
rect 960 -1955 975 -1925
rect 1005 -1955 1020 -1925
rect 960 -1995 1020 -1955
rect 960 -2025 975 -1995
rect 1005 -2025 1020 -1995
rect 960 -2060 1020 -2025
rect 960 -2090 975 -2060
rect 1005 -2090 1020 -2060
rect 960 -2120 1020 -2090
rect 960 -2150 975 -2120
rect 1005 -2150 1020 -2120
rect 960 -2185 1020 -2150
rect 960 -2215 975 -2185
rect 1005 -2215 1020 -2185
rect 960 -2255 1020 -2215
rect 960 -2285 975 -2255
rect 1005 -2285 1020 -2255
rect 960 -2325 1020 -2285
rect 960 -2355 975 -2325
rect 1005 -2355 1020 -2325
rect 960 -2395 1020 -2355
rect 960 -2425 975 -2395
rect 1005 -2425 1020 -2395
rect 960 -2460 1020 -2425
rect 960 -2490 975 -2460
rect 1005 -2490 1020 -2460
rect 960 -2520 1020 -2490
rect 960 -2550 975 -2520
rect 1005 -2550 1020 -2520
rect 960 -2585 1020 -2550
rect 960 -2615 975 -2585
rect 1005 -2615 1020 -2585
rect 960 -2655 1020 -2615
rect 960 -2685 975 -2655
rect 1005 -2685 1020 -2655
rect 960 -2725 1020 -2685
rect 960 -2755 975 -2725
rect 1005 -2755 1020 -2725
rect 960 -2795 1020 -2755
rect 960 -2825 975 -2795
rect 1005 -2825 1020 -2795
rect 960 -2860 1020 -2825
rect 960 -2890 975 -2860
rect 1005 -2890 1020 -2860
rect 960 -2905 1020 -2890
rect 1310 -1320 1370 -1305
rect 1310 -1350 1325 -1320
rect 1355 -1350 1370 -1320
rect 1310 -1385 1370 -1350
rect 1310 -1415 1325 -1385
rect 1355 -1415 1370 -1385
rect 1310 -1455 1370 -1415
rect 1310 -1485 1325 -1455
rect 1355 -1485 1370 -1455
rect 1310 -1525 1370 -1485
rect 1310 -1555 1325 -1525
rect 1355 -1555 1370 -1525
rect 1310 -1595 1370 -1555
rect 1310 -1625 1325 -1595
rect 1355 -1625 1370 -1595
rect 1310 -1660 1370 -1625
rect 1310 -1690 1325 -1660
rect 1355 -1690 1370 -1660
rect 1310 -1720 1370 -1690
rect 1310 -1750 1325 -1720
rect 1355 -1750 1370 -1720
rect 1310 -1785 1370 -1750
rect 1310 -1815 1325 -1785
rect 1355 -1815 1370 -1785
rect 1310 -1855 1370 -1815
rect 1310 -1885 1325 -1855
rect 1355 -1885 1370 -1855
rect 1310 -1925 1370 -1885
rect 1310 -1955 1325 -1925
rect 1355 -1955 1370 -1925
rect 1310 -1995 1370 -1955
rect 1310 -2025 1325 -1995
rect 1355 -2025 1370 -1995
rect 1310 -2060 1370 -2025
rect 1310 -2090 1325 -2060
rect 1355 -2090 1370 -2060
rect 1310 -2120 1370 -2090
rect 1310 -2150 1325 -2120
rect 1355 -2150 1370 -2120
rect 1310 -2185 1370 -2150
rect 1310 -2215 1325 -2185
rect 1355 -2215 1370 -2185
rect 1310 -2255 1370 -2215
rect 1310 -2285 1325 -2255
rect 1355 -2285 1370 -2255
rect 1310 -2325 1370 -2285
rect 1310 -2355 1325 -2325
rect 1355 -2355 1370 -2325
rect 1310 -2395 1370 -2355
rect 1310 -2425 1325 -2395
rect 1355 -2425 1370 -2395
rect 1310 -2460 1370 -2425
rect 1310 -2490 1325 -2460
rect 1355 -2490 1370 -2460
rect 1310 -2520 1370 -2490
rect 1310 -2550 1325 -2520
rect 1355 -2550 1370 -2520
rect 1310 -2585 1370 -2550
rect 1310 -2615 1325 -2585
rect 1355 -2615 1370 -2585
rect 1310 -2655 1370 -2615
rect 1310 -2685 1325 -2655
rect 1355 -2685 1370 -2655
rect 1310 -2725 1370 -2685
rect 1310 -2755 1325 -2725
rect 1355 -2755 1370 -2725
rect 1310 -2795 1370 -2755
rect 1310 -2825 1325 -2795
rect 1355 -2825 1370 -2795
rect 1310 -2860 1370 -2825
rect 1310 -2890 1325 -2860
rect 1355 -2890 1370 -2860
rect 1310 -2905 1370 -2890
rect 1660 -1320 1720 -1305
rect 1660 -1350 1675 -1320
rect 1705 -1350 1720 -1320
rect 1660 -1385 1720 -1350
rect 1660 -1415 1675 -1385
rect 1705 -1415 1720 -1385
rect 1660 -1455 1720 -1415
rect 1660 -1485 1675 -1455
rect 1705 -1485 1720 -1455
rect 1660 -1525 1720 -1485
rect 1660 -1555 1675 -1525
rect 1705 -1555 1720 -1525
rect 1660 -1595 1720 -1555
rect 1660 -1625 1675 -1595
rect 1705 -1625 1720 -1595
rect 1660 -1660 1720 -1625
rect 1660 -1690 1675 -1660
rect 1705 -1690 1720 -1660
rect 1660 -1720 1720 -1690
rect 1660 -1750 1675 -1720
rect 1705 -1750 1720 -1720
rect 1660 -1785 1720 -1750
rect 1660 -1815 1675 -1785
rect 1705 -1815 1720 -1785
rect 1660 -1855 1720 -1815
rect 1660 -1885 1675 -1855
rect 1705 -1885 1720 -1855
rect 1660 -1925 1720 -1885
rect 1660 -1955 1675 -1925
rect 1705 -1955 1720 -1925
rect 1660 -1995 1720 -1955
rect 1660 -2025 1675 -1995
rect 1705 -2025 1720 -1995
rect 1660 -2060 1720 -2025
rect 1660 -2090 1675 -2060
rect 1705 -2090 1720 -2060
rect 1660 -2120 1720 -2090
rect 1660 -2150 1675 -2120
rect 1705 -2150 1720 -2120
rect 1660 -2185 1720 -2150
rect 1660 -2215 1675 -2185
rect 1705 -2215 1720 -2185
rect 1660 -2255 1720 -2215
rect 1660 -2285 1675 -2255
rect 1705 -2285 1720 -2255
rect 1660 -2325 1720 -2285
rect 1660 -2355 1675 -2325
rect 1705 -2355 1720 -2325
rect 1660 -2395 1720 -2355
rect 1660 -2425 1675 -2395
rect 1705 -2425 1720 -2395
rect 1660 -2460 1720 -2425
rect 1660 -2490 1675 -2460
rect 1705 -2490 1720 -2460
rect 1660 -2520 1720 -2490
rect 1660 -2550 1675 -2520
rect 1705 -2550 1720 -2520
rect 1660 -2585 1720 -2550
rect 1660 -2615 1675 -2585
rect 1705 -2615 1720 -2585
rect 1660 -2655 1720 -2615
rect 1660 -2685 1675 -2655
rect 1705 -2685 1720 -2655
rect 1660 -2725 1720 -2685
rect 1660 -2755 1675 -2725
rect 1705 -2755 1720 -2725
rect 1660 -2795 1720 -2755
rect 1660 -2825 1675 -2795
rect 1705 -2825 1720 -2795
rect 1660 -2860 1720 -2825
rect 1660 -2890 1675 -2860
rect 1705 -2890 1720 -2860
rect 1660 -2905 1720 -2890
rect 2010 -1320 2070 -1305
rect 2010 -1350 2025 -1320
rect 2055 -1350 2070 -1320
rect 2010 -1385 2070 -1350
rect 2010 -1415 2025 -1385
rect 2055 -1415 2070 -1385
rect 2010 -1455 2070 -1415
rect 2010 -1485 2025 -1455
rect 2055 -1485 2070 -1455
rect 2010 -1525 2070 -1485
rect 2010 -1555 2025 -1525
rect 2055 -1555 2070 -1525
rect 2010 -1595 2070 -1555
rect 2010 -1625 2025 -1595
rect 2055 -1625 2070 -1595
rect 2010 -1660 2070 -1625
rect 2010 -1690 2025 -1660
rect 2055 -1690 2070 -1660
rect 2010 -1720 2070 -1690
rect 2010 -1750 2025 -1720
rect 2055 -1750 2070 -1720
rect 2010 -1785 2070 -1750
rect 2010 -1815 2025 -1785
rect 2055 -1815 2070 -1785
rect 2010 -1855 2070 -1815
rect 2010 -1885 2025 -1855
rect 2055 -1885 2070 -1855
rect 2010 -1925 2070 -1885
rect 2010 -1955 2025 -1925
rect 2055 -1955 2070 -1925
rect 2010 -1995 2070 -1955
rect 2010 -2025 2025 -1995
rect 2055 -2025 2070 -1995
rect 2010 -2060 2070 -2025
rect 2010 -2090 2025 -2060
rect 2055 -2090 2070 -2060
rect 2010 -2120 2070 -2090
rect 2010 -2150 2025 -2120
rect 2055 -2150 2070 -2120
rect 2010 -2185 2070 -2150
rect 2010 -2215 2025 -2185
rect 2055 -2215 2070 -2185
rect 2010 -2255 2070 -2215
rect 2010 -2285 2025 -2255
rect 2055 -2285 2070 -2255
rect 2010 -2325 2070 -2285
rect 2010 -2355 2025 -2325
rect 2055 -2355 2070 -2325
rect 2010 -2395 2070 -2355
rect 2010 -2425 2025 -2395
rect 2055 -2425 2070 -2395
rect 2010 -2460 2070 -2425
rect 2010 -2490 2025 -2460
rect 2055 -2490 2070 -2460
rect 2010 -2520 2070 -2490
rect 2010 -2550 2025 -2520
rect 2055 -2550 2070 -2520
rect 2010 -2585 2070 -2550
rect 2010 -2615 2025 -2585
rect 2055 -2615 2070 -2585
rect 2010 -2655 2070 -2615
rect 2010 -2685 2025 -2655
rect 2055 -2685 2070 -2655
rect 2010 -2725 2070 -2685
rect 2010 -2755 2025 -2725
rect 2055 -2755 2070 -2725
rect 2010 -2795 2070 -2755
rect 2010 -2825 2025 -2795
rect 2055 -2825 2070 -2795
rect 2010 -2860 2070 -2825
rect 2010 -2890 2025 -2860
rect 2055 -2890 2070 -2860
rect 2010 -2905 2070 -2890
rect 2360 -1320 2420 -1305
rect 2360 -1350 2375 -1320
rect 2405 -1350 2420 -1320
rect 2360 -1385 2420 -1350
rect 2360 -1415 2375 -1385
rect 2405 -1415 2420 -1385
rect 2360 -1455 2420 -1415
rect 2360 -1485 2375 -1455
rect 2405 -1485 2420 -1455
rect 2360 -1525 2420 -1485
rect 2360 -1555 2375 -1525
rect 2405 -1555 2420 -1525
rect 2360 -1595 2420 -1555
rect 2360 -1625 2375 -1595
rect 2405 -1625 2420 -1595
rect 2360 -1660 2420 -1625
rect 2360 -1690 2375 -1660
rect 2405 -1690 2420 -1660
rect 2360 -1720 2420 -1690
rect 2360 -1750 2375 -1720
rect 2405 -1750 2420 -1720
rect 2360 -1785 2420 -1750
rect 2360 -1815 2375 -1785
rect 2405 -1815 2420 -1785
rect 2360 -1855 2420 -1815
rect 2360 -1885 2375 -1855
rect 2405 -1885 2420 -1855
rect 2360 -1925 2420 -1885
rect 2360 -1955 2375 -1925
rect 2405 -1955 2420 -1925
rect 2360 -1995 2420 -1955
rect 2360 -2025 2375 -1995
rect 2405 -2025 2420 -1995
rect 2360 -2060 2420 -2025
rect 2360 -2090 2375 -2060
rect 2405 -2090 2420 -2060
rect 2360 -2120 2420 -2090
rect 2360 -2150 2375 -2120
rect 2405 -2150 2420 -2120
rect 2360 -2185 2420 -2150
rect 2360 -2215 2375 -2185
rect 2405 -2215 2420 -2185
rect 2360 -2255 2420 -2215
rect 2360 -2285 2375 -2255
rect 2405 -2285 2420 -2255
rect 2360 -2325 2420 -2285
rect 2360 -2355 2375 -2325
rect 2405 -2355 2420 -2325
rect 2360 -2395 2420 -2355
rect 2360 -2425 2375 -2395
rect 2405 -2425 2420 -2395
rect 2360 -2460 2420 -2425
rect 2360 -2490 2375 -2460
rect 2405 -2490 2420 -2460
rect 2360 -2520 2420 -2490
rect 2360 -2550 2375 -2520
rect 2405 -2550 2420 -2520
rect 2360 -2585 2420 -2550
rect 2360 -2615 2375 -2585
rect 2405 -2615 2420 -2585
rect 2360 -2655 2420 -2615
rect 2360 -2685 2375 -2655
rect 2405 -2685 2420 -2655
rect 2360 -2725 2420 -2685
rect 2360 -2755 2375 -2725
rect 2405 -2755 2420 -2725
rect 2360 -2795 2420 -2755
rect 2360 -2825 2375 -2795
rect 2405 -2825 2420 -2795
rect 2360 -2860 2420 -2825
rect 2360 -2890 2375 -2860
rect 2405 -2890 2420 -2860
rect 2360 -2905 2420 -2890
rect 2710 -1320 2770 -1305
rect 2710 -1350 2725 -1320
rect 2755 -1350 2770 -1320
rect 2710 -1385 2770 -1350
rect 2710 -1415 2725 -1385
rect 2755 -1415 2770 -1385
rect 2710 -1455 2770 -1415
rect 2710 -1485 2725 -1455
rect 2755 -1485 2770 -1455
rect 2710 -1525 2770 -1485
rect 2710 -1555 2725 -1525
rect 2755 -1555 2770 -1525
rect 2710 -1595 2770 -1555
rect 2710 -1625 2725 -1595
rect 2755 -1625 2770 -1595
rect 2710 -1660 2770 -1625
rect 2710 -1690 2725 -1660
rect 2755 -1690 2770 -1660
rect 2710 -1720 2770 -1690
rect 2710 -1750 2725 -1720
rect 2755 -1750 2770 -1720
rect 2710 -1785 2770 -1750
rect 2710 -1815 2725 -1785
rect 2755 -1815 2770 -1785
rect 2710 -1855 2770 -1815
rect 2710 -1885 2725 -1855
rect 2755 -1885 2770 -1855
rect 2710 -1925 2770 -1885
rect 2710 -1955 2725 -1925
rect 2755 -1955 2770 -1925
rect 2710 -1995 2770 -1955
rect 2710 -2025 2725 -1995
rect 2755 -2025 2770 -1995
rect 2710 -2060 2770 -2025
rect 2710 -2090 2725 -2060
rect 2755 -2090 2770 -2060
rect 2710 -2120 2770 -2090
rect 2710 -2150 2725 -2120
rect 2755 -2150 2770 -2120
rect 2710 -2185 2770 -2150
rect 2710 -2215 2725 -2185
rect 2755 -2215 2770 -2185
rect 2710 -2255 2770 -2215
rect 2710 -2285 2725 -2255
rect 2755 -2285 2770 -2255
rect 2710 -2325 2770 -2285
rect 2710 -2355 2725 -2325
rect 2755 -2355 2770 -2325
rect 2710 -2395 2770 -2355
rect 2710 -2425 2725 -2395
rect 2755 -2425 2770 -2395
rect 2710 -2460 2770 -2425
rect 2710 -2490 2725 -2460
rect 2755 -2490 2770 -2460
rect 2710 -2520 2770 -2490
rect 2710 -2550 2725 -2520
rect 2755 -2550 2770 -2520
rect 2710 -2585 2770 -2550
rect 2710 -2615 2725 -2585
rect 2755 -2615 2770 -2585
rect 2710 -2655 2770 -2615
rect 2710 -2685 2725 -2655
rect 2755 -2685 2770 -2655
rect 2710 -2725 2770 -2685
rect 2710 -2755 2725 -2725
rect 2755 -2755 2770 -2725
rect 2710 -2795 2770 -2755
rect 2710 -2825 2725 -2795
rect 2755 -2825 2770 -2795
rect 2710 -2860 2770 -2825
rect 2710 -2890 2725 -2860
rect 2755 -2890 2770 -2860
rect 2710 -2905 2770 -2890
rect 3060 -1320 3120 -1305
rect 3060 -1350 3075 -1320
rect 3105 -1350 3120 -1320
rect 3060 -1385 3120 -1350
rect 3060 -1415 3075 -1385
rect 3105 -1415 3120 -1385
rect 3060 -1455 3120 -1415
rect 3060 -1485 3075 -1455
rect 3105 -1485 3120 -1455
rect 3060 -1525 3120 -1485
rect 3060 -1555 3075 -1525
rect 3105 -1555 3120 -1525
rect 3060 -1595 3120 -1555
rect 3060 -1625 3075 -1595
rect 3105 -1625 3120 -1595
rect 3060 -1660 3120 -1625
rect 3060 -1690 3075 -1660
rect 3105 -1690 3120 -1660
rect 3060 -1720 3120 -1690
rect 3060 -1750 3075 -1720
rect 3105 -1750 3120 -1720
rect 3060 -1785 3120 -1750
rect 3060 -1815 3075 -1785
rect 3105 -1815 3120 -1785
rect 3060 -1855 3120 -1815
rect 3060 -1885 3075 -1855
rect 3105 -1885 3120 -1855
rect 3060 -1925 3120 -1885
rect 3060 -1955 3075 -1925
rect 3105 -1955 3120 -1925
rect 3060 -1995 3120 -1955
rect 3060 -2025 3075 -1995
rect 3105 -2025 3120 -1995
rect 3060 -2060 3120 -2025
rect 3060 -2090 3075 -2060
rect 3105 -2090 3120 -2060
rect 3060 -2120 3120 -2090
rect 3060 -2150 3075 -2120
rect 3105 -2150 3120 -2120
rect 3060 -2185 3120 -2150
rect 3060 -2215 3075 -2185
rect 3105 -2215 3120 -2185
rect 3060 -2255 3120 -2215
rect 3060 -2285 3075 -2255
rect 3105 -2285 3120 -2255
rect 3060 -2325 3120 -2285
rect 3060 -2355 3075 -2325
rect 3105 -2355 3120 -2325
rect 3060 -2395 3120 -2355
rect 3060 -2425 3075 -2395
rect 3105 -2425 3120 -2395
rect 3060 -2460 3120 -2425
rect 3060 -2490 3075 -2460
rect 3105 -2490 3120 -2460
rect 3060 -2520 3120 -2490
rect 3060 -2550 3075 -2520
rect 3105 -2550 3120 -2520
rect 3060 -2585 3120 -2550
rect 3060 -2615 3075 -2585
rect 3105 -2615 3120 -2585
rect 3060 -2655 3120 -2615
rect 3060 -2685 3075 -2655
rect 3105 -2685 3120 -2655
rect 3060 -2725 3120 -2685
rect 3060 -2755 3075 -2725
rect 3105 -2755 3120 -2725
rect 3060 -2795 3120 -2755
rect 3060 -2825 3075 -2795
rect 3105 -2825 3120 -2795
rect 3060 -2860 3120 -2825
rect 3060 -2890 3075 -2860
rect 3105 -2890 3120 -2860
rect 3060 -2905 3120 -2890
rect 5860 -1320 5920 -1305
rect 5860 -1350 5875 -1320
rect 5905 -1350 5920 -1320
rect 5860 -1385 5920 -1350
rect 5860 -1415 5875 -1385
rect 5905 -1415 5920 -1385
rect 5860 -1455 5920 -1415
rect 5860 -1485 5875 -1455
rect 5905 -1485 5920 -1455
rect 5860 -1525 5920 -1485
rect 5860 -1555 5875 -1525
rect 5905 -1555 5920 -1525
rect 5860 -1595 5920 -1555
rect 5860 -1625 5875 -1595
rect 5905 -1625 5920 -1595
rect 5860 -1660 5920 -1625
rect 5860 -1690 5875 -1660
rect 5905 -1690 5920 -1660
rect 5860 -1720 5920 -1690
rect 5860 -1750 5875 -1720
rect 5905 -1750 5920 -1720
rect 5860 -1785 5920 -1750
rect 5860 -1815 5875 -1785
rect 5905 -1815 5920 -1785
rect 5860 -1855 5920 -1815
rect 5860 -1885 5875 -1855
rect 5905 -1885 5920 -1855
rect 5860 -1925 5920 -1885
rect 5860 -1955 5875 -1925
rect 5905 -1955 5920 -1925
rect 5860 -1995 5920 -1955
rect 5860 -2025 5875 -1995
rect 5905 -2025 5920 -1995
rect 5860 -2060 5920 -2025
rect 5860 -2090 5875 -2060
rect 5905 -2090 5920 -2060
rect 5860 -2120 5920 -2090
rect 5860 -2150 5875 -2120
rect 5905 -2150 5920 -2120
rect 5860 -2185 5920 -2150
rect 5860 -2215 5875 -2185
rect 5905 -2215 5920 -2185
rect 5860 -2255 5920 -2215
rect 5860 -2285 5875 -2255
rect 5905 -2285 5920 -2255
rect 5860 -2325 5920 -2285
rect 5860 -2355 5875 -2325
rect 5905 -2355 5920 -2325
rect 5860 -2395 5920 -2355
rect 5860 -2425 5875 -2395
rect 5905 -2425 5920 -2395
rect 5860 -2460 5920 -2425
rect 5860 -2490 5875 -2460
rect 5905 -2490 5920 -2460
rect 5860 -2520 5920 -2490
rect 5860 -2550 5875 -2520
rect 5905 -2550 5920 -2520
rect 5860 -2585 5920 -2550
rect 5860 -2615 5875 -2585
rect 5905 -2615 5920 -2585
rect 5860 -2655 5920 -2615
rect 5860 -2685 5875 -2655
rect 5905 -2685 5920 -2655
rect 5860 -2725 5920 -2685
rect 5860 -2755 5875 -2725
rect 5905 -2755 5920 -2725
rect 5860 -2795 5920 -2755
rect 5860 -2825 5875 -2795
rect 5905 -2825 5920 -2795
rect 5860 -2860 5920 -2825
rect 5860 -2890 5875 -2860
rect 5905 -2890 5920 -2860
rect 5860 -2905 5920 -2890
rect 6210 -1320 6270 -1305
rect 6210 -1350 6225 -1320
rect 6255 -1350 6270 -1320
rect 6210 -1385 6270 -1350
rect 6210 -1415 6225 -1385
rect 6255 -1415 6270 -1385
rect 6210 -1455 6270 -1415
rect 6210 -1485 6225 -1455
rect 6255 -1485 6270 -1455
rect 6210 -1525 6270 -1485
rect 6210 -1555 6225 -1525
rect 6255 -1555 6270 -1525
rect 6210 -1595 6270 -1555
rect 6210 -1625 6225 -1595
rect 6255 -1625 6270 -1595
rect 6210 -1660 6270 -1625
rect 6210 -1690 6225 -1660
rect 6255 -1690 6270 -1660
rect 6210 -1720 6270 -1690
rect 6210 -1750 6225 -1720
rect 6255 -1750 6270 -1720
rect 6210 -1785 6270 -1750
rect 6210 -1815 6225 -1785
rect 6255 -1815 6270 -1785
rect 6210 -1855 6270 -1815
rect 6210 -1885 6225 -1855
rect 6255 -1885 6270 -1855
rect 6210 -1925 6270 -1885
rect 6210 -1955 6225 -1925
rect 6255 -1955 6270 -1925
rect 6210 -1995 6270 -1955
rect 6210 -2025 6225 -1995
rect 6255 -2025 6270 -1995
rect 6210 -2060 6270 -2025
rect 6210 -2090 6225 -2060
rect 6255 -2090 6270 -2060
rect 6210 -2120 6270 -2090
rect 6210 -2150 6225 -2120
rect 6255 -2150 6270 -2120
rect 6210 -2185 6270 -2150
rect 6210 -2215 6225 -2185
rect 6255 -2215 6270 -2185
rect 6210 -2255 6270 -2215
rect 6210 -2285 6225 -2255
rect 6255 -2285 6270 -2255
rect 6210 -2325 6270 -2285
rect 6210 -2355 6225 -2325
rect 6255 -2355 6270 -2325
rect 6210 -2395 6270 -2355
rect 6210 -2425 6225 -2395
rect 6255 -2425 6270 -2395
rect 6210 -2460 6270 -2425
rect 6210 -2490 6225 -2460
rect 6255 -2490 6270 -2460
rect 6210 -2520 6270 -2490
rect 6210 -2550 6225 -2520
rect 6255 -2550 6270 -2520
rect 6210 -2585 6270 -2550
rect 6210 -2615 6225 -2585
rect 6255 -2615 6270 -2585
rect 6210 -2655 6270 -2615
rect 6210 -2685 6225 -2655
rect 6255 -2685 6270 -2655
rect 6210 -2725 6270 -2685
rect 6210 -2755 6225 -2725
rect 6255 -2755 6270 -2725
rect 6210 -2795 6270 -2755
rect 6210 -2825 6225 -2795
rect 6255 -2825 6270 -2795
rect 6210 -2860 6270 -2825
rect 6210 -2890 6225 -2860
rect 6255 -2890 6270 -2860
rect 6210 -2905 6270 -2890
rect 6560 -1320 6620 -1305
rect 6560 -1350 6575 -1320
rect 6605 -1350 6620 -1320
rect 6560 -1385 6620 -1350
rect 6560 -1415 6575 -1385
rect 6605 -1415 6620 -1385
rect 6560 -1455 6620 -1415
rect 6560 -1485 6575 -1455
rect 6605 -1485 6620 -1455
rect 6560 -1525 6620 -1485
rect 6560 -1555 6575 -1525
rect 6605 -1555 6620 -1525
rect 6560 -1595 6620 -1555
rect 6560 -1625 6575 -1595
rect 6605 -1625 6620 -1595
rect 6560 -1660 6620 -1625
rect 6560 -1690 6575 -1660
rect 6605 -1690 6620 -1660
rect 6560 -1720 6620 -1690
rect 6560 -1750 6575 -1720
rect 6605 -1750 6620 -1720
rect 6560 -1785 6620 -1750
rect 6560 -1815 6575 -1785
rect 6605 -1815 6620 -1785
rect 6560 -1855 6620 -1815
rect 6560 -1885 6575 -1855
rect 6605 -1885 6620 -1855
rect 6560 -1925 6620 -1885
rect 6560 -1955 6575 -1925
rect 6605 -1955 6620 -1925
rect 6560 -1995 6620 -1955
rect 6560 -2025 6575 -1995
rect 6605 -2025 6620 -1995
rect 6560 -2060 6620 -2025
rect 6560 -2090 6575 -2060
rect 6605 -2090 6620 -2060
rect 6560 -2120 6620 -2090
rect 6560 -2150 6575 -2120
rect 6605 -2150 6620 -2120
rect 6560 -2185 6620 -2150
rect 6560 -2215 6575 -2185
rect 6605 -2215 6620 -2185
rect 6560 -2255 6620 -2215
rect 6560 -2285 6575 -2255
rect 6605 -2285 6620 -2255
rect 6560 -2325 6620 -2285
rect 6560 -2355 6575 -2325
rect 6605 -2355 6620 -2325
rect 6560 -2395 6620 -2355
rect 6560 -2425 6575 -2395
rect 6605 -2425 6620 -2395
rect 6560 -2460 6620 -2425
rect 6560 -2490 6575 -2460
rect 6605 -2490 6620 -2460
rect 6560 -2520 6620 -2490
rect 6560 -2550 6575 -2520
rect 6605 -2550 6620 -2520
rect 6560 -2585 6620 -2550
rect 6560 -2615 6575 -2585
rect 6605 -2615 6620 -2585
rect 6560 -2655 6620 -2615
rect 6560 -2685 6575 -2655
rect 6605 -2685 6620 -2655
rect 6560 -2725 6620 -2685
rect 6560 -2755 6575 -2725
rect 6605 -2755 6620 -2725
rect 6560 -2795 6620 -2755
rect 6560 -2825 6575 -2795
rect 6605 -2825 6620 -2795
rect 6560 -2860 6620 -2825
rect 6560 -2890 6575 -2860
rect 6605 -2890 6620 -2860
rect 6560 -2905 6620 -2890
rect 6910 -1320 6970 -1305
rect 6910 -1350 6925 -1320
rect 6955 -1350 6970 -1320
rect 6910 -1385 6970 -1350
rect 6910 -1415 6925 -1385
rect 6955 -1415 6970 -1385
rect 6910 -1455 6970 -1415
rect 6910 -1485 6925 -1455
rect 6955 -1485 6970 -1455
rect 6910 -1525 6970 -1485
rect 6910 -1555 6925 -1525
rect 6955 -1555 6970 -1525
rect 6910 -1595 6970 -1555
rect 6910 -1625 6925 -1595
rect 6955 -1625 6970 -1595
rect 6910 -1660 6970 -1625
rect 6910 -1690 6925 -1660
rect 6955 -1690 6970 -1660
rect 6910 -1720 6970 -1690
rect 6910 -1750 6925 -1720
rect 6955 -1750 6970 -1720
rect 6910 -1785 6970 -1750
rect 6910 -1815 6925 -1785
rect 6955 -1815 6970 -1785
rect 6910 -1855 6970 -1815
rect 6910 -1885 6925 -1855
rect 6955 -1885 6970 -1855
rect 6910 -1925 6970 -1885
rect 6910 -1955 6925 -1925
rect 6955 -1955 6970 -1925
rect 6910 -1995 6970 -1955
rect 6910 -2025 6925 -1995
rect 6955 -2025 6970 -1995
rect 6910 -2060 6970 -2025
rect 6910 -2090 6925 -2060
rect 6955 -2090 6970 -2060
rect 6910 -2120 6970 -2090
rect 6910 -2150 6925 -2120
rect 6955 -2150 6970 -2120
rect 6910 -2185 6970 -2150
rect 6910 -2215 6925 -2185
rect 6955 -2215 6970 -2185
rect 6910 -2255 6970 -2215
rect 6910 -2285 6925 -2255
rect 6955 -2285 6970 -2255
rect 6910 -2325 6970 -2285
rect 6910 -2355 6925 -2325
rect 6955 -2355 6970 -2325
rect 6910 -2395 6970 -2355
rect 6910 -2425 6925 -2395
rect 6955 -2425 6970 -2395
rect 6910 -2460 6970 -2425
rect 6910 -2490 6925 -2460
rect 6955 -2490 6970 -2460
rect 6910 -2520 6970 -2490
rect 6910 -2550 6925 -2520
rect 6955 -2550 6970 -2520
rect 6910 -2585 6970 -2550
rect 6910 -2615 6925 -2585
rect 6955 -2615 6970 -2585
rect 6910 -2655 6970 -2615
rect 6910 -2685 6925 -2655
rect 6955 -2685 6970 -2655
rect 6910 -2725 6970 -2685
rect 6910 -2755 6925 -2725
rect 6955 -2755 6970 -2725
rect 6910 -2795 6970 -2755
rect 6910 -2825 6925 -2795
rect 6955 -2825 6970 -2795
rect 6910 -2860 6970 -2825
rect 6910 -2890 6925 -2860
rect 6955 -2890 6970 -2860
rect 6910 -2905 6970 -2890
rect 7260 -1320 7320 -1305
rect 7260 -1350 7275 -1320
rect 7305 -1350 7320 -1320
rect 7260 -1385 7320 -1350
rect 7260 -1415 7275 -1385
rect 7305 -1415 7320 -1385
rect 7260 -1455 7320 -1415
rect 7260 -1485 7275 -1455
rect 7305 -1485 7320 -1455
rect 7260 -1525 7320 -1485
rect 7260 -1555 7275 -1525
rect 7305 -1555 7320 -1525
rect 7260 -1595 7320 -1555
rect 7260 -1625 7275 -1595
rect 7305 -1625 7320 -1595
rect 7260 -1660 7320 -1625
rect 7260 -1690 7275 -1660
rect 7305 -1690 7320 -1660
rect 7260 -1720 7320 -1690
rect 7260 -1750 7275 -1720
rect 7305 -1750 7320 -1720
rect 7260 -1785 7320 -1750
rect 7260 -1815 7275 -1785
rect 7305 -1815 7320 -1785
rect 7260 -1855 7320 -1815
rect 7260 -1885 7275 -1855
rect 7305 -1885 7320 -1855
rect 7260 -1925 7320 -1885
rect 7260 -1955 7275 -1925
rect 7305 -1955 7320 -1925
rect 7260 -1995 7320 -1955
rect 7260 -2025 7275 -1995
rect 7305 -2025 7320 -1995
rect 7260 -2060 7320 -2025
rect 7260 -2090 7275 -2060
rect 7305 -2090 7320 -2060
rect 7260 -2120 7320 -2090
rect 7260 -2150 7275 -2120
rect 7305 -2150 7320 -2120
rect 7260 -2185 7320 -2150
rect 7260 -2215 7275 -2185
rect 7305 -2215 7320 -2185
rect 7260 -2255 7320 -2215
rect 7260 -2285 7275 -2255
rect 7305 -2285 7320 -2255
rect 7260 -2325 7320 -2285
rect 7260 -2355 7275 -2325
rect 7305 -2355 7320 -2325
rect 7260 -2395 7320 -2355
rect 7260 -2425 7275 -2395
rect 7305 -2425 7320 -2395
rect 7260 -2460 7320 -2425
rect 7260 -2490 7275 -2460
rect 7305 -2490 7320 -2460
rect 7260 -2520 7320 -2490
rect 7260 -2550 7275 -2520
rect 7305 -2550 7320 -2520
rect 7260 -2585 7320 -2550
rect 7260 -2615 7275 -2585
rect 7305 -2615 7320 -2585
rect 7260 -2655 7320 -2615
rect 7260 -2685 7275 -2655
rect 7305 -2685 7320 -2655
rect 7260 -2725 7320 -2685
rect 7260 -2755 7275 -2725
rect 7305 -2755 7320 -2725
rect 7260 -2795 7320 -2755
rect 7260 -2825 7275 -2795
rect 7305 -2825 7320 -2795
rect 7260 -2860 7320 -2825
rect 7260 -2890 7275 -2860
rect 7305 -2890 7320 -2860
rect 7260 -2905 7320 -2890
rect 7610 -1320 7670 -1305
rect 7610 -1350 7625 -1320
rect 7655 -1350 7670 -1320
rect 7610 -1385 7670 -1350
rect 7610 -1415 7625 -1385
rect 7655 -1415 7670 -1385
rect 7610 -1455 7670 -1415
rect 7610 -1485 7625 -1455
rect 7655 -1485 7670 -1455
rect 7610 -1525 7670 -1485
rect 7610 -1555 7625 -1525
rect 7655 -1555 7670 -1525
rect 7610 -1595 7670 -1555
rect 7610 -1625 7625 -1595
rect 7655 -1625 7670 -1595
rect 7610 -1660 7670 -1625
rect 7610 -1690 7625 -1660
rect 7655 -1690 7670 -1660
rect 7610 -1720 7670 -1690
rect 7610 -1750 7625 -1720
rect 7655 -1750 7670 -1720
rect 7610 -1785 7670 -1750
rect 7610 -1815 7625 -1785
rect 7655 -1815 7670 -1785
rect 7610 -1855 7670 -1815
rect 7610 -1885 7625 -1855
rect 7655 -1885 7670 -1855
rect 7610 -1925 7670 -1885
rect 7610 -1955 7625 -1925
rect 7655 -1955 7670 -1925
rect 7610 -1995 7670 -1955
rect 7610 -2025 7625 -1995
rect 7655 -2025 7670 -1995
rect 7610 -2060 7670 -2025
rect 7610 -2090 7625 -2060
rect 7655 -2090 7670 -2060
rect 7610 -2120 7670 -2090
rect 7610 -2150 7625 -2120
rect 7655 -2150 7670 -2120
rect 7610 -2185 7670 -2150
rect 7610 -2215 7625 -2185
rect 7655 -2215 7670 -2185
rect 7610 -2255 7670 -2215
rect 7610 -2285 7625 -2255
rect 7655 -2285 7670 -2255
rect 7610 -2325 7670 -2285
rect 7610 -2355 7625 -2325
rect 7655 -2355 7670 -2325
rect 7610 -2395 7670 -2355
rect 7610 -2425 7625 -2395
rect 7655 -2425 7670 -2395
rect 7610 -2460 7670 -2425
rect 7610 -2490 7625 -2460
rect 7655 -2490 7670 -2460
rect 7610 -2520 7670 -2490
rect 7610 -2550 7625 -2520
rect 7655 -2550 7670 -2520
rect 7610 -2585 7670 -2550
rect 7610 -2615 7625 -2585
rect 7655 -2615 7670 -2585
rect 7610 -2655 7670 -2615
rect 7610 -2685 7625 -2655
rect 7655 -2685 7670 -2655
rect 7610 -2725 7670 -2685
rect 7610 -2755 7625 -2725
rect 7655 -2755 7670 -2725
rect 7610 -2795 7670 -2755
rect 7610 -2825 7625 -2795
rect 7655 -2825 7670 -2795
rect 7610 -2860 7670 -2825
rect 7610 -2890 7625 -2860
rect 7655 -2890 7670 -2860
rect 7610 -2905 7670 -2890
rect 7960 -1320 8020 -1305
rect 7960 -1350 7975 -1320
rect 8005 -1350 8020 -1320
rect 7960 -1385 8020 -1350
rect 7960 -1415 7975 -1385
rect 8005 -1415 8020 -1385
rect 7960 -1455 8020 -1415
rect 7960 -1485 7975 -1455
rect 8005 -1485 8020 -1455
rect 7960 -1525 8020 -1485
rect 7960 -1555 7975 -1525
rect 8005 -1555 8020 -1525
rect 7960 -1595 8020 -1555
rect 7960 -1625 7975 -1595
rect 8005 -1625 8020 -1595
rect 7960 -1660 8020 -1625
rect 7960 -1690 7975 -1660
rect 8005 -1690 8020 -1660
rect 7960 -1720 8020 -1690
rect 7960 -1750 7975 -1720
rect 8005 -1750 8020 -1720
rect 7960 -1785 8020 -1750
rect 7960 -1815 7975 -1785
rect 8005 -1815 8020 -1785
rect 7960 -1855 8020 -1815
rect 7960 -1885 7975 -1855
rect 8005 -1885 8020 -1855
rect 7960 -1925 8020 -1885
rect 7960 -1955 7975 -1925
rect 8005 -1955 8020 -1925
rect 7960 -1995 8020 -1955
rect 7960 -2025 7975 -1995
rect 8005 -2025 8020 -1995
rect 7960 -2060 8020 -2025
rect 7960 -2090 7975 -2060
rect 8005 -2090 8020 -2060
rect 7960 -2120 8020 -2090
rect 7960 -2150 7975 -2120
rect 8005 -2150 8020 -2120
rect 7960 -2185 8020 -2150
rect 7960 -2215 7975 -2185
rect 8005 -2215 8020 -2185
rect 7960 -2255 8020 -2215
rect 7960 -2285 7975 -2255
rect 8005 -2285 8020 -2255
rect 7960 -2325 8020 -2285
rect 7960 -2355 7975 -2325
rect 8005 -2355 8020 -2325
rect 7960 -2395 8020 -2355
rect 7960 -2425 7975 -2395
rect 8005 -2425 8020 -2395
rect 7960 -2460 8020 -2425
rect 7960 -2490 7975 -2460
rect 8005 -2490 8020 -2460
rect 7960 -2520 8020 -2490
rect 7960 -2550 7975 -2520
rect 8005 -2550 8020 -2520
rect 7960 -2585 8020 -2550
rect 7960 -2615 7975 -2585
rect 8005 -2615 8020 -2585
rect 7960 -2655 8020 -2615
rect 7960 -2685 7975 -2655
rect 8005 -2685 8020 -2655
rect 7960 -2725 8020 -2685
rect 7960 -2755 7975 -2725
rect 8005 -2755 8020 -2725
rect 7960 -2795 8020 -2755
rect 7960 -2825 7975 -2795
rect 8005 -2825 8020 -2795
rect 7960 -2860 8020 -2825
rect 7960 -2890 7975 -2860
rect 8005 -2890 8020 -2860
rect 7960 -2905 8020 -2890
rect 8310 -1320 8370 -1305
rect 8310 -1350 8325 -1320
rect 8355 -1350 8370 -1320
rect 8310 -1385 8370 -1350
rect 8310 -1415 8325 -1385
rect 8355 -1415 8370 -1385
rect 8310 -1455 8370 -1415
rect 8310 -1485 8325 -1455
rect 8355 -1485 8370 -1455
rect 8310 -1525 8370 -1485
rect 8310 -1555 8325 -1525
rect 8355 -1555 8370 -1525
rect 8310 -1595 8370 -1555
rect 8310 -1625 8325 -1595
rect 8355 -1625 8370 -1595
rect 8310 -1660 8370 -1625
rect 8310 -1690 8325 -1660
rect 8355 -1690 8370 -1660
rect 8310 -1720 8370 -1690
rect 8310 -1750 8325 -1720
rect 8355 -1750 8370 -1720
rect 8310 -1785 8370 -1750
rect 8310 -1815 8325 -1785
rect 8355 -1815 8370 -1785
rect 8310 -1855 8370 -1815
rect 8310 -1885 8325 -1855
rect 8355 -1885 8370 -1855
rect 8310 -1925 8370 -1885
rect 8310 -1955 8325 -1925
rect 8355 -1955 8370 -1925
rect 8310 -1995 8370 -1955
rect 8310 -2025 8325 -1995
rect 8355 -2025 8370 -1995
rect 8310 -2060 8370 -2025
rect 8310 -2090 8325 -2060
rect 8355 -2090 8370 -2060
rect 8310 -2120 8370 -2090
rect 8310 -2150 8325 -2120
rect 8355 -2150 8370 -2120
rect 8310 -2185 8370 -2150
rect 8310 -2215 8325 -2185
rect 8355 -2215 8370 -2185
rect 8310 -2255 8370 -2215
rect 8310 -2285 8325 -2255
rect 8355 -2285 8370 -2255
rect 8310 -2325 8370 -2285
rect 8310 -2355 8325 -2325
rect 8355 -2355 8370 -2325
rect 8310 -2395 8370 -2355
rect 8310 -2425 8325 -2395
rect 8355 -2425 8370 -2395
rect 8310 -2460 8370 -2425
rect 8310 -2490 8325 -2460
rect 8355 -2490 8370 -2460
rect 8310 -2520 8370 -2490
rect 8310 -2550 8325 -2520
rect 8355 -2550 8370 -2520
rect 8310 -2585 8370 -2550
rect 8310 -2615 8325 -2585
rect 8355 -2615 8370 -2585
rect 8310 -2655 8370 -2615
rect 8310 -2685 8325 -2655
rect 8355 -2685 8370 -2655
rect 8310 -2725 8370 -2685
rect 8310 -2755 8325 -2725
rect 8355 -2755 8370 -2725
rect 8310 -2795 8370 -2755
rect 8310 -2825 8325 -2795
rect 8355 -2825 8370 -2795
rect 8310 -2860 8370 -2825
rect 8310 -2890 8325 -2860
rect 8355 -2890 8370 -2860
rect 8310 -2905 8370 -2890
rect 8660 -1320 8720 -1305
rect 8660 -1350 8675 -1320
rect 8705 -1350 8720 -1320
rect 8660 -1385 8720 -1350
rect 8660 -1415 8675 -1385
rect 8705 -1415 8720 -1385
rect 8660 -1455 8720 -1415
rect 8660 -1485 8675 -1455
rect 8705 -1485 8720 -1455
rect 8660 -1525 8720 -1485
rect 8660 -1555 8675 -1525
rect 8705 -1555 8720 -1525
rect 8660 -1595 8720 -1555
rect 8660 -1625 8675 -1595
rect 8705 -1625 8720 -1595
rect 8660 -1660 8720 -1625
rect 8660 -1690 8675 -1660
rect 8705 -1690 8720 -1660
rect 8660 -1720 8720 -1690
rect 8660 -1750 8675 -1720
rect 8705 -1750 8720 -1720
rect 8660 -1785 8720 -1750
rect 8660 -1815 8675 -1785
rect 8705 -1815 8720 -1785
rect 8660 -1855 8720 -1815
rect 8660 -1885 8675 -1855
rect 8705 -1885 8720 -1855
rect 8660 -1925 8720 -1885
rect 8660 -1955 8675 -1925
rect 8705 -1955 8720 -1925
rect 8660 -1995 8720 -1955
rect 8660 -2025 8675 -1995
rect 8705 -2025 8720 -1995
rect 8660 -2060 8720 -2025
rect 8660 -2090 8675 -2060
rect 8705 -2090 8720 -2060
rect 8660 -2120 8720 -2090
rect 8660 -2150 8675 -2120
rect 8705 -2150 8720 -2120
rect 8660 -2185 8720 -2150
rect 8660 -2215 8675 -2185
rect 8705 -2215 8720 -2185
rect 8660 -2255 8720 -2215
rect 8660 -2285 8675 -2255
rect 8705 -2285 8720 -2255
rect 8660 -2325 8720 -2285
rect 8660 -2355 8675 -2325
rect 8705 -2355 8720 -2325
rect 8660 -2395 8720 -2355
rect 8660 -2425 8675 -2395
rect 8705 -2425 8720 -2395
rect 8660 -2460 8720 -2425
rect 8660 -2490 8675 -2460
rect 8705 -2490 8720 -2460
rect 8660 -2520 8720 -2490
rect 8660 -2550 8675 -2520
rect 8705 -2550 8720 -2520
rect 8660 -2585 8720 -2550
rect 8660 -2615 8675 -2585
rect 8705 -2615 8720 -2585
rect 8660 -2655 8720 -2615
rect 8660 -2685 8675 -2655
rect 8705 -2685 8720 -2655
rect 8660 -2725 8720 -2685
rect 8660 -2755 8675 -2725
rect 8705 -2755 8720 -2725
rect 8660 -2795 8720 -2755
rect 8660 -2825 8675 -2795
rect 8705 -2825 8720 -2795
rect 8660 -2860 8720 -2825
rect 8660 -2890 8675 -2860
rect 8705 -2890 8720 -2860
rect 8660 -2905 8720 -2890
rect 9010 -1320 9070 -1305
rect 9010 -1350 9025 -1320
rect 9055 -1350 9070 -1320
rect 9010 -1385 9070 -1350
rect 9010 -1415 9025 -1385
rect 9055 -1415 9070 -1385
rect 9010 -1455 9070 -1415
rect 9010 -1485 9025 -1455
rect 9055 -1485 9070 -1455
rect 9010 -1525 9070 -1485
rect 9010 -1555 9025 -1525
rect 9055 -1555 9070 -1525
rect 9010 -1595 9070 -1555
rect 9010 -1625 9025 -1595
rect 9055 -1625 9070 -1595
rect 9010 -1660 9070 -1625
rect 9010 -1690 9025 -1660
rect 9055 -1690 9070 -1660
rect 9010 -1720 9070 -1690
rect 9010 -1750 9025 -1720
rect 9055 -1750 9070 -1720
rect 9010 -1785 9070 -1750
rect 9010 -1815 9025 -1785
rect 9055 -1815 9070 -1785
rect 9010 -1855 9070 -1815
rect 9010 -1885 9025 -1855
rect 9055 -1885 9070 -1855
rect 9010 -1925 9070 -1885
rect 9010 -1955 9025 -1925
rect 9055 -1955 9070 -1925
rect 9010 -1995 9070 -1955
rect 9010 -2025 9025 -1995
rect 9055 -2025 9070 -1995
rect 9010 -2060 9070 -2025
rect 9010 -2090 9025 -2060
rect 9055 -2090 9070 -2060
rect 9010 -2120 9070 -2090
rect 9010 -2150 9025 -2120
rect 9055 -2150 9070 -2120
rect 9010 -2185 9070 -2150
rect 9010 -2215 9025 -2185
rect 9055 -2215 9070 -2185
rect 9010 -2255 9070 -2215
rect 9010 -2285 9025 -2255
rect 9055 -2285 9070 -2255
rect 9010 -2325 9070 -2285
rect 9010 -2355 9025 -2325
rect 9055 -2355 9070 -2325
rect 9010 -2395 9070 -2355
rect 9010 -2425 9025 -2395
rect 9055 -2425 9070 -2395
rect 9010 -2460 9070 -2425
rect 9010 -2490 9025 -2460
rect 9055 -2490 9070 -2460
rect 9010 -2520 9070 -2490
rect 9010 -2550 9025 -2520
rect 9055 -2550 9070 -2520
rect 9010 -2585 9070 -2550
rect 9010 -2615 9025 -2585
rect 9055 -2615 9070 -2585
rect 9010 -2655 9070 -2615
rect 9010 -2685 9025 -2655
rect 9055 -2685 9070 -2655
rect 9010 -2725 9070 -2685
rect 9010 -2755 9025 -2725
rect 9055 -2755 9070 -2725
rect 9010 -2795 9070 -2755
rect 9010 -2825 9025 -2795
rect 9055 -2825 9070 -2795
rect 9010 -2860 9070 -2825
rect 9010 -2890 9025 -2860
rect 9055 -2890 9070 -2860
rect 9010 -2905 9070 -2890
rect 3410 -3020 3470 -3005
rect 3410 -3050 3425 -3020
rect 3455 -3050 3470 -3020
rect 3410 -3085 3470 -3050
rect 3410 -3115 3425 -3085
rect 3455 -3115 3470 -3085
rect 3410 -3155 3470 -3115
rect 3410 -3185 3425 -3155
rect 3455 -3185 3470 -3155
rect 3410 -3225 3470 -3185
rect 3410 -3255 3425 -3225
rect 3455 -3255 3470 -3225
rect 3410 -3295 3470 -3255
rect 3410 -3325 3425 -3295
rect 3455 -3325 3470 -3295
rect 3410 -3360 3470 -3325
rect 3410 -3390 3425 -3360
rect 3455 -3390 3470 -3360
rect 3410 -3420 3470 -3390
rect 3410 -3450 3425 -3420
rect 3455 -3450 3470 -3420
rect 3410 -3485 3470 -3450
rect 3410 -3515 3425 -3485
rect 3455 -3515 3470 -3485
rect 3410 -3555 3470 -3515
rect 3410 -3585 3425 -3555
rect 3455 -3585 3470 -3555
rect 3410 -3625 3470 -3585
rect 3410 -3655 3425 -3625
rect 3455 -3655 3470 -3625
rect 3410 -3695 3470 -3655
rect 3410 -3725 3425 -3695
rect 3455 -3725 3470 -3695
rect 3410 -3760 3470 -3725
rect 3410 -3790 3425 -3760
rect 3455 -3790 3470 -3760
rect 3410 -3820 3470 -3790
rect 3410 -3850 3425 -3820
rect 3455 -3850 3470 -3820
rect 3410 -3885 3470 -3850
rect 3410 -3915 3425 -3885
rect 3455 -3915 3470 -3885
rect 3410 -3955 3470 -3915
rect 3410 -3985 3425 -3955
rect 3455 -3985 3470 -3955
rect 3410 -4025 3470 -3985
rect 3410 -4055 3425 -4025
rect 3455 -4055 3470 -4025
rect 3410 -4095 3470 -4055
rect 3410 -4125 3425 -4095
rect 3455 -4125 3470 -4095
rect 3410 -4160 3470 -4125
rect 3410 -4190 3425 -4160
rect 3455 -4190 3470 -4160
rect 3410 -4220 3470 -4190
rect 3410 -4250 3425 -4220
rect 3455 -4250 3470 -4220
rect 3410 -4285 3470 -4250
rect 3410 -4315 3425 -4285
rect 3455 -4315 3470 -4285
rect 3410 -4355 3470 -4315
rect 3410 -4385 3425 -4355
rect 3455 -4385 3470 -4355
rect 3410 -4425 3470 -4385
rect 3410 -4455 3425 -4425
rect 3455 -4455 3470 -4425
rect 3410 -4495 3470 -4455
rect 3410 -4525 3425 -4495
rect 3455 -4525 3470 -4495
rect 3410 -4560 3470 -4525
rect 3410 -4590 3425 -4560
rect 3455 -4590 3470 -4560
rect 3410 -4605 3470 -4590
rect 3760 -3020 3820 -3005
rect 3760 -3050 3775 -3020
rect 3805 -3050 3820 -3020
rect 3760 -3085 3820 -3050
rect 3760 -3115 3775 -3085
rect 3805 -3115 3820 -3085
rect 3760 -3155 3820 -3115
rect 3760 -3185 3775 -3155
rect 3805 -3185 3820 -3155
rect 3760 -3225 3820 -3185
rect 3760 -3255 3775 -3225
rect 3805 -3255 3820 -3225
rect 3760 -3295 3820 -3255
rect 3760 -3325 3775 -3295
rect 3805 -3325 3820 -3295
rect 3760 -3360 3820 -3325
rect 3760 -3390 3775 -3360
rect 3805 -3390 3820 -3360
rect 3760 -3420 3820 -3390
rect 3760 -3450 3775 -3420
rect 3805 -3450 3820 -3420
rect 3760 -3485 3820 -3450
rect 3760 -3515 3775 -3485
rect 3805 -3515 3820 -3485
rect 3760 -3555 3820 -3515
rect 3760 -3585 3775 -3555
rect 3805 -3585 3820 -3555
rect 3760 -3625 3820 -3585
rect 3760 -3655 3775 -3625
rect 3805 -3655 3820 -3625
rect 3760 -3695 3820 -3655
rect 3760 -3725 3775 -3695
rect 3805 -3725 3820 -3695
rect 3760 -3760 3820 -3725
rect 3760 -3790 3775 -3760
rect 3805 -3790 3820 -3760
rect 3760 -3820 3820 -3790
rect 3760 -3850 3775 -3820
rect 3805 -3850 3820 -3820
rect 3760 -3885 3820 -3850
rect 3760 -3915 3775 -3885
rect 3805 -3915 3820 -3885
rect 3760 -3955 3820 -3915
rect 3760 -3985 3775 -3955
rect 3805 -3985 3820 -3955
rect 3760 -4025 3820 -3985
rect 3760 -4055 3775 -4025
rect 3805 -4055 3820 -4025
rect 3760 -4095 3820 -4055
rect 3760 -4125 3775 -4095
rect 3805 -4125 3820 -4095
rect 3760 -4160 3820 -4125
rect 3760 -4190 3775 -4160
rect 3805 -4190 3820 -4160
rect 3760 -4220 3820 -4190
rect 3760 -4250 3775 -4220
rect 3805 -4250 3820 -4220
rect 3760 -4285 3820 -4250
rect 3760 -4315 3775 -4285
rect 3805 -4315 3820 -4285
rect 3760 -4355 3820 -4315
rect 3760 -4385 3775 -4355
rect 3805 -4385 3820 -4355
rect 3760 -4425 3820 -4385
rect 3760 -4455 3775 -4425
rect 3805 -4455 3820 -4425
rect 3760 -4495 3820 -4455
rect 3760 -4525 3775 -4495
rect 3805 -4525 3820 -4495
rect 3760 -4560 3820 -4525
rect 3760 -4590 3775 -4560
rect 3805 -4590 3820 -4560
rect 3760 -4605 3820 -4590
rect 4110 -3020 4170 -3005
rect 4110 -3050 4125 -3020
rect 4155 -3050 4170 -3020
rect 4110 -3085 4170 -3050
rect 4110 -3115 4125 -3085
rect 4155 -3115 4170 -3085
rect 4110 -3155 4170 -3115
rect 4110 -3185 4125 -3155
rect 4155 -3185 4170 -3155
rect 4110 -3225 4170 -3185
rect 4110 -3255 4125 -3225
rect 4155 -3255 4170 -3225
rect 4110 -3295 4170 -3255
rect 4110 -3325 4125 -3295
rect 4155 -3325 4170 -3295
rect 4110 -3360 4170 -3325
rect 4110 -3390 4125 -3360
rect 4155 -3390 4170 -3360
rect 4110 -3420 4170 -3390
rect 4110 -3450 4125 -3420
rect 4155 -3450 4170 -3420
rect 4110 -3485 4170 -3450
rect 4110 -3515 4125 -3485
rect 4155 -3515 4170 -3485
rect 4110 -3555 4170 -3515
rect 4110 -3585 4125 -3555
rect 4155 -3585 4170 -3555
rect 4110 -3625 4170 -3585
rect 4110 -3655 4125 -3625
rect 4155 -3655 4170 -3625
rect 4110 -3695 4170 -3655
rect 4110 -3725 4125 -3695
rect 4155 -3725 4170 -3695
rect 4110 -3760 4170 -3725
rect 4110 -3790 4125 -3760
rect 4155 -3790 4170 -3760
rect 4110 -3820 4170 -3790
rect 4110 -3850 4125 -3820
rect 4155 -3850 4170 -3820
rect 4110 -3885 4170 -3850
rect 4110 -3915 4125 -3885
rect 4155 -3915 4170 -3885
rect 4110 -3955 4170 -3915
rect 4110 -3985 4125 -3955
rect 4155 -3985 4170 -3955
rect 4110 -4025 4170 -3985
rect 4110 -4055 4125 -4025
rect 4155 -4055 4170 -4025
rect 4110 -4095 4170 -4055
rect 4110 -4125 4125 -4095
rect 4155 -4125 4170 -4095
rect 4110 -4160 4170 -4125
rect 4110 -4190 4125 -4160
rect 4155 -4190 4170 -4160
rect 4110 -4220 4170 -4190
rect 4110 -4250 4125 -4220
rect 4155 -4250 4170 -4220
rect 4110 -4285 4170 -4250
rect 4110 -4315 4125 -4285
rect 4155 -4315 4170 -4285
rect 4110 -4355 4170 -4315
rect 4110 -4385 4125 -4355
rect 4155 -4385 4170 -4355
rect 4110 -4425 4170 -4385
rect 4110 -4455 4125 -4425
rect 4155 -4455 4170 -4425
rect 4110 -4495 4170 -4455
rect 4110 -4525 4125 -4495
rect 4155 -4525 4170 -4495
rect 4110 -4560 4170 -4525
rect 4110 -4590 4125 -4560
rect 4155 -4590 4170 -4560
rect 4110 -4605 4170 -4590
rect 4460 -3020 4520 -3005
rect 4460 -3050 4475 -3020
rect 4505 -3050 4520 -3020
rect 4460 -3085 4520 -3050
rect 4460 -3115 4475 -3085
rect 4505 -3115 4520 -3085
rect 4460 -3155 4520 -3115
rect 4460 -3185 4475 -3155
rect 4505 -3185 4520 -3155
rect 4460 -3225 4520 -3185
rect 4460 -3255 4475 -3225
rect 4505 -3255 4520 -3225
rect 4460 -3295 4520 -3255
rect 4460 -3325 4475 -3295
rect 4505 -3325 4520 -3295
rect 4460 -3360 4520 -3325
rect 4460 -3390 4475 -3360
rect 4505 -3390 4520 -3360
rect 4460 -3420 4520 -3390
rect 4460 -3450 4475 -3420
rect 4505 -3450 4520 -3420
rect 4460 -3485 4520 -3450
rect 4460 -3515 4475 -3485
rect 4505 -3515 4520 -3485
rect 4460 -3555 4520 -3515
rect 4460 -3585 4475 -3555
rect 4505 -3585 4520 -3555
rect 4460 -3625 4520 -3585
rect 4460 -3655 4475 -3625
rect 4505 -3655 4520 -3625
rect 4460 -3695 4520 -3655
rect 4460 -3725 4475 -3695
rect 4505 -3725 4520 -3695
rect 4460 -3760 4520 -3725
rect 4460 -3790 4475 -3760
rect 4505 -3790 4520 -3760
rect 4460 -3820 4520 -3790
rect 4460 -3850 4475 -3820
rect 4505 -3850 4520 -3820
rect 4460 -3885 4520 -3850
rect 4460 -3915 4475 -3885
rect 4505 -3915 4520 -3885
rect 4460 -3955 4520 -3915
rect 4460 -3985 4475 -3955
rect 4505 -3985 4520 -3955
rect 4460 -4025 4520 -3985
rect 4460 -4055 4475 -4025
rect 4505 -4055 4520 -4025
rect 4460 -4095 4520 -4055
rect 4460 -4125 4475 -4095
rect 4505 -4125 4520 -4095
rect 4460 -4160 4520 -4125
rect 4460 -4190 4475 -4160
rect 4505 -4190 4520 -4160
rect 4460 -4220 4520 -4190
rect 4460 -4250 4475 -4220
rect 4505 -4250 4520 -4220
rect 4460 -4285 4520 -4250
rect 4460 -4315 4475 -4285
rect 4505 -4315 4520 -4285
rect 4460 -4355 4520 -4315
rect 4460 -4385 4475 -4355
rect 4505 -4385 4520 -4355
rect 4460 -4425 4520 -4385
rect 4460 -4455 4475 -4425
rect 4505 -4455 4520 -4425
rect 4460 -4495 4520 -4455
rect 4460 -4525 4475 -4495
rect 4505 -4525 4520 -4495
rect 4460 -4560 4520 -4525
rect 4460 -4590 4475 -4560
rect 4505 -4590 4520 -4560
rect 4460 -4605 4520 -4590
rect 4810 -3020 4870 -3005
rect 4810 -3050 4825 -3020
rect 4855 -3050 4870 -3020
rect 4810 -3085 4870 -3050
rect 4810 -3115 4825 -3085
rect 4855 -3115 4870 -3085
rect 4810 -3155 4870 -3115
rect 4810 -3185 4825 -3155
rect 4855 -3185 4870 -3155
rect 4810 -3225 4870 -3185
rect 4810 -3255 4825 -3225
rect 4855 -3255 4870 -3225
rect 4810 -3295 4870 -3255
rect 4810 -3325 4825 -3295
rect 4855 -3325 4870 -3295
rect 4810 -3360 4870 -3325
rect 4810 -3390 4825 -3360
rect 4855 -3390 4870 -3360
rect 4810 -3420 4870 -3390
rect 4810 -3450 4825 -3420
rect 4855 -3450 4870 -3420
rect 4810 -3485 4870 -3450
rect 4810 -3515 4825 -3485
rect 4855 -3515 4870 -3485
rect 4810 -3555 4870 -3515
rect 4810 -3585 4825 -3555
rect 4855 -3585 4870 -3555
rect 4810 -3625 4870 -3585
rect 4810 -3655 4825 -3625
rect 4855 -3655 4870 -3625
rect 4810 -3695 4870 -3655
rect 4810 -3725 4825 -3695
rect 4855 -3725 4870 -3695
rect 4810 -3760 4870 -3725
rect 4810 -3790 4825 -3760
rect 4855 -3790 4870 -3760
rect 4810 -3820 4870 -3790
rect 4810 -3850 4825 -3820
rect 4855 -3850 4870 -3820
rect 4810 -3885 4870 -3850
rect 4810 -3915 4825 -3885
rect 4855 -3915 4870 -3885
rect 4810 -3955 4870 -3915
rect 4810 -3985 4825 -3955
rect 4855 -3985 4870 -3955
rect 4810 -4025 4870 -3985
rect 4810 -4055 4825 -4025
rect 4855 -4055 4870 -4025
rect 4810 -4095 4870 -4055
rect 4810 -4125 4825 -4095
rect 4855 -4125 4870 -4095
rect 4810 -4160 4870 -4125
rect 4810 -4190 4825 -4160
rect 4855 -4190 4870 -4160
rect 4810 -4220 4870 -4190
rect 4810 -4250 4825 -4220
rect 4855 -4250 4870 -4220
rect 4810 -4285 4870 -4250
rect 4810 -4315 4825 -4285
rect 4855 -4315 4870 -4285
rect 4810 -4355 4870 -4315
rect 4810 -4385 4825 -4355
rect 4855 -4385 4870 -4355
rect 4810 -4425 4870 -4385
rect 4810 -4455 4825 -4425
rect 4855 -4455 4870 -4425
rect 4810 -4495 4870 -4455
rect 4810 -4525 4825 -4495
rect 4855 -4525 4870 -4495
rect 4810 -4560 4870 -4525
rect 4810 -4590 4825 -4560
rect 4855 -4590 4870 -4560
rect 4810 -4605 4870 -4590
rect 5160 -3020 5220 -3005
rect 5160 -3050 5175 -3020
rect 5205 -3050 5220 -3020
rect 5160 -3085 5220 -3050
rect 5160 -3115 5175 -3085
rect 5205 -3115 5220 -3085
rect 5160 -3155 5220 -3115
rect 5160 -3185 5175 -3155
rect 5205 -3185 5220 -3155
rect 5160 -3225 5220 -3185
rect 5160 -3255 5175 -3225
rect 5205 -3255 5220 -3225
rect 5160 -3295 5220 -3255
rect 5160 -3325 5175 -3295
rect 5205 -3325 5220 -3295
rect 5160 -3360 5220 -3325
rect 5160 -3390 5175 -3360
rect 5205 -3390 5220 -3360
rect 5160 -3420 5220 -3390
rect 5160 -3450 5175 -3420
rect 5205 -3450 5220 -3420
rect 5160 -3485 5220 -3450
rect 5160 -3515 5175 -3485
rect 5205 -3515 5220 -3485
rect 5160 -3555 5220 -3515
rect 5160 -3585 5175 -3555
rect 5205 -3585 5220 -3555
rect 5160 -3625 5220 -3585
rect 5160 -3655 5175 -3625
rect 5205 -3655 5220 -3625
rect 5160 -3695 5220 -3655
rect 5160 -3725 5175 -3695
rect 5205 -3725 5220 -3695
rect 5160 -3760 5220 -3725
rect 5160 -3790 5175 -3760
rect 5205 -3790 5220 -3760
rect 5160 -3820 5220 -3790
rect 5160 -3850 5175 -3820
rect 5205 -3850 5220 -3820
rect 5160 -3885 5220 -3850
rect 5160 -3915 5175 -3885
rect 5205 -3915 5220 -3885
rect 5160 -3955 5220 -3915
rect 5160 -3985 5175 -3955
rect 5205 -3985 5220 -3955
rect 5160 -4025 5220 -3985
rect 5160 -4055 5175 -4025
rect 5205 -4055 5220 -4025
rect 5160 -4095 5220 -4055
rect 5160 -4125 5175 -4095
rect 5205 -4125 5220 -4095
rect 5160 -4160 5220 -4125
rect 5160 -4190 5175 -4160
rect 5205 -4190 5220 -4160
rect 5160 -4220 5220 -4190
rect 5160 -4250 5175 -4220
rect 5205 -4250 5220 -4220
rect 5160 -4285 5220 -4250
rect 5160 -4315 5175 -4285
rect 5205 -4315 5220 -4285
rect 5160 -4355 5220 -4315
rect 5160 -4385 5175 -4355
rect 5205 -4385 5220 -4355
rect 5160 -4425 5220 -4385
rect 5160 -4455 5175 -4425
rect 5205 -4455 5220 -4425
rect 5160 -4495 5220 -4455
rect 5160 -4525 5175 -4495
rect 5205 -4525 5220 -4495
rect 5160 -4560 5220 -4525
rect 5160 -4590 5175 -4560
rect 5205 -4590 5220 -4560
rect 5160 -4605 5220 -4590
rect 5510 -3020 5570 -3005
rect 5510 -3050 5525 -3020
rect 5555 -3050 5570 -3020
rect 5510 -3085 5570 -3050
rect 5510 -3115 5525 -3085
rect 5555 -3115 5570 -3085
rect 5510 -3155 5570 -3115
rect 5510 -3185 5525 -3155
rect 5555 -3185 5570 -3155
rect 5510 -3225 5570 -3185
rect 5510 -3255 5525 -3225
rect 5555 -3255 5570 -3225
rect 5510 -3295 5570 -3255
rect 5510 -3325 5525 -3295
rect 5555 -3325 5570 -3295
rect 5510 -3360 5570 -3325
rect 5510 -3390 5525 -3360
rect 5555 -3390 5570 -3360
rect 5510 -3420 5570 -3390
rect 5510 -3450 5525 -3420
rect 5555 -3450 5570 -3420
rect 5510 -3485 5570 -3450
rect 5510 -3515 5525 -3485
rect 5555 -3515 5570 -3485
rect 5510 -3555 5570 -3515
rect 5510 -3585 5525 -3555
rect 5555 -3585 5570 -3555
rect 5510 -3625 5570 -3585
rect 5510 -3655 5525 -3625
rect 5555 -3655 5570 -3625
rect 5510 -3695 5570 -3655
rect 5510 -3725 5525 -3695
rect 5555 -3725 5570 -3695
rect 5510 -3760 5570 -3725
rect 5510 -3790 5525 -3760
rect 5555 -3790 5570 -3760
rect 5510 -3820 5570 -3790
rect 5510 -3850 5525 -3820
rect 5555 -3850 5570 -3820
rect 5510 -3885 5570 -3850
rect 5510 -3915 5525 -3885
rect 5555 -3915 5570 -3885
rect 5510 -3955 5570 -3915
rect 5510 -3985 5525 -3955
rect 5555 -3985 5570 -3955
rect 5510 -4025 5570 -3985
rect 5510 -4055 5525 -4025
rect 5555 -4055 5570 -4025
rect 5510 -4095 5570 -4055
rect 5510 -4125 5525 -4095
rect 5555 -4125 5570 -4095
rect 5510 -4160 5570 -4125
rect 5510 -4190 5525 -4160
rect 5555 -4190 5570 -4160
rect 5510 -4220 5570 -4190
rect 5510 -4250 5525 -4220
rect 5555 -4250 5570 -4220
rect 5510 -4285 5570 -4250
rect 5510 -4315 5525 -4285
rect 5555 -4315 5570 -4285
rect 5510 -4355 5570 -4315
rect 5510 -4385 5525 -4355
rect 5555 -4385 5570 -4355
rect 5510 -4425 5570 -4385
rect 5510 -4455 5525 -4425
rect 5555 -4455 5570 -4425
rect 5510 -4495 5570 -4455
rect 5510 -4525 5525 -4495
rect 5555 -4525 5570 -4495
rect 5510 -4560 5570 -4525
rect 5510 -4590 5525 -4560
rect 5555 -4590 5570 -4560
rect 5510 -4605 5570 -4590
<< via2 >>
rect 2115 19280 2145 19310
rect 2115 19215 2145 19245
rect 2115 19145 2145 19175
rect 2115 19075 2145 19105
rect 2115 19005 2145 19035
rect 2115 18940 2145 18970
rect 2115 18880 2145 18910
rect 2115 18815 2145 18845
rect 2115 18745 2145 18775
rect 2115 18675 2145 18705
rect 2115 18605 2145 18635
rect 2115 18540 2145 18570
rect 2115 18480 2145 18510
rect 2115 18415 2145 18445
rect 2115 18345 2145 18375
rect 2115 18275 2145 18305
rect 2115 18205 2145 18235
rect 2115 18140 2145 18170
rect 2115 18080 2145 18110
rect 2115 18015 2145 18045
rect 2115 17945 2145 17975
rect 2115 17875 2145 17905
rect 2115 17805 2145 17835
rect 2115 17740 2145 17770
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 1325 9605 1355 9635
rect 1325 9540 1355 9570
rect 1325 9470 1355 9500
rect 1325 9400 1355 9430
rect 1325 9330 1355 9360
rect 1325 9265 1355 9295
rect 1325 9205 1355 9235
rect 1325 9140 1355 9170
rect 1325 9070 1355 9100
rect 1325 9000 1355 9030
rect 1325 8930 1355 8960
rect 1325 8865 1355 8895
rect 1325 8805 1355 8835
rect 1325 8740 1355 8770
rect 1325 8670 1355 8700
rect 1325 8600 1355 8630
rect 1325 8530 1355 8560
rect 1325 8465 1355 8495
rect 1325 8405 1355 8435
rect 1325 8340 1355 8370
rect 1325 8270 1355 8300
rect 1325 8200 1355 8230
rect 1325 8130 1355 8160
rect 2250 9605 2280 9635
rect 2250 9540 2280 9570
rect 2250 9470 2280 9500
rect 2250 9400 2280 9430
rect 2250 9330 2280 9360
rect 2250 9265 2280 9295
rect 2250 9205 2280 9235
rect 2250 9140 2280 9170
rect 2250 9070 2280 9100
rect 2250 9000 2280 9030
rect 2250 8930 2280 8960
rect 2250 8865 2280 8895
rect 2250 8805 2280 8835
rect 2250 8740 2280 8770
rect 2250 8670 2280 8700
rect 2250 8600 2280 8630
rect 2250 8530 2280 8560
rect 2250 8465 2280 8495
rect 2250 8405 2280 8435
rect 2250 8340 2280 8370
rect 2250 8270 2280 8300
rect 2250 8200 2280 8230
rect 2250 8130 2280 8160
rect 6705 9605 6735 9635
rect 6705 9540 6735 9570
rect 6705 9470 6735 9500
rect 6705 9400 6735 9430
rect 6705 9330 6735 9360
rect 6705 9265 6735 9295
rect 6705 9205 6735 9235
rect 6705 9140 6735 9170
rect 6705 9070 6735 9100
rect 6705 9000 6735 9030
rect 6705 8930 6735 8960
rect 6705 8865 6735 8895
rect 6705 8805 6735 8835
rect 6705 8740 6735 8770
rect 6705 8670 6735 8700
rect 6705 8600 6735 8630
rect 6705 8530 6735 8560
rect 6705 8465 6735 8495
rect 6705 8405 6735 8435
rect 6705 8340 6735 8370
rect 6705 8270 6735 8300
rect 6705 8200 6735 8230
rect 6705 8130 6735 8160
rect 7625 9605 7655 9635
rect 7625 9540 7655 9570
rect 7625 9470 7655 9500
rect 7625 9400 7655 9430
rect 7625 9330 7655 9360
rect 7625 9265 7655 9295
rect 7625 9205 7655 9235
rect 7625 9140 7655 9170
rect 7625 9070 7655 9100
rect 7625 9000 7655 9030
rect 7625 8930 7655 8960
rect 7625 8865 7655 8895
rect 7625 8805 7655 8835
rect 7625 8740 7655 8770
rect 7625 8670 7655 8700
rect 7625 8600 7655 8630
rect 7625 8530 7655 8560
rect 7625 8465 7655 8495
rect 7625 8405 7655 8435
rect 7625 8340 7655 8370
rect 7625 8270 7655 8300
rect 7625 8200 7655 8230
rect 7625 8130 7655 8160
rect 3180 7925 3210 7955
rect 3240 7925 3270 7955
rect 3180 7855 3210 7885
rect 3240 7855 3270 7885
rect 3180 7785 3210 7815
rect 3240 7785 3270 7815
rect 3180 7715 3210 7745
rect 3240 7715 3270 7745
rect 3180 7650 3210 7680
rect 3240 7650 3270 7680
rect 3180 7590 3210 7620
rect 3240 7590 3270 7620
rect 3180 7525 3210 7555
rect 3240 7525 3270 7555
rect 3180 7455 3210 7485
rect 3240 7455 3270 7485
rect 3180 7385 3210 7415
rect 3240 7385 3270 7415
rect 3180 7315 3210 7345
rect 3240 7315 3270 7345
rect 3180 7250 3210 7280
rect 3240 7250 3270 7280
rect 3180 7190 3210 7220
rect 3240 7190 3270 7220
rect 3180 7125 3210 7155
rect 3240 7125 3270 7155
rect 3180 7055 3210 7085
rect 3240 7055 3270 7085
rect 3180 6985 3210 7015
rect 3240 6985 3270 7015
rect 3180 6915 3210 6945
rect 3240 6915 3270 6945
rect 3180 6850 3210 6880
rect 3240 6850 3270 6880
rect 3180 6790 3210 6820
rect 3240 6790 3270 6820
rect 3180 6725 3210 6755
rect 3240 6725 3270 6755
rect 3180 6655 3210 6685
rect 3240 6655 3270 6685
rect 3180 6585 3210 6615
rect 3240 6585 3270 6615
rect 3180 6515 3210 6545
rect 3240 6515 3270 6545
rect 3180 6450 3210 6480
rect 3240 6450 3270 6480
rect 3350 7925 3380 7955
rect 3350 7855 3380 7885
rect 3350 7785 3380 7815
rect 3350 7715 3380 7745
rect 3350 7650 3380 7680
rect 3350 7590 3380 7620
rect 3350 7525 3380 7555
rect 3350 7455 3380 7485
rect 3350 7385 3380 7415
rect 3350 7315 3380 7345
rect 3350 7250 3380 7280
rect 3350 7190 3380 7220
rect 3350 7125 3380 7155
rect 3350 7055 3380 7085
rect 3350 6985 3380 7015
rect 3350 6915 3380 6945
rect 3350 6850 3380 6880
rect 3350 6790 3380 6820
rect 3350 6725 3380 6755
rect 3350 6655 3380 6685
rect 3350 6585 3380 6615
rect 3350 6515 3380 6545
rect 3350 6450 3380 6480
rect -75 -1350 -45 -1320
rect -75 -1415 -45 -1385
rect -75 -1485 -45 -1455
rect -75 -1555 -45 -1525
rect -75 -1625 -45 -1595
rect -75 -1690 -45 -1660
rect -75 -1750 -45 -1720
rect -75 -1815 -45 -1785
rect -75 -1885 -45 -1855
rect -75 -1955 -45 -1925
rect -75 -2025 -45 -1995
rect -75 -2090 -45 -2060
rect -75 -2150 -45 -2120
rect -75 -2215 -45 -2185
rect -75 -2285 -45 -2255
rect -75 -2355 -45 -2325
rect -75 -2425 -45 -2395
rect -75 -2490 -45 -2460
rect -75 -2550 -45 -2520
rect -75 -2615 -45 -2585
rect -75 -2685 -45 -2655
rect -75 -2755 -45 -2725
rect -75 -2825 -45 -2795
rect -75 -2890 -45 -2860
rect 275 -1350 305 -1320
rect 275 -1415 305 -1385
rect 275 -1485 305 -1455
rect 275 -1555 305 -1525
rect 275 -1625 305 -1595
rect 275 -1690 305 -1660
rect 275 -1750 305 -1720
rect 275 -1815 305 -1785
rect 275 -1885 305 -1855
rect 275 -1955 305 -1925
rect 275 -2025 305 -1995
rect 275 -2090 305 -2060
rect 275 -2150 305 -2120
rect 275 -2215 305 -2185
rect 275 -2285 305 -2255
rect 275 -2355 305 -2325
rect 275 -2425 305 -2395
rect 275 -2490 305 -2460
rect 275 -2550 305 -2520
rect 275 -2615 305 -2585
rect 275 -2685 305 -2655
rect 275 -2755 305 -2725
rect 275 -2825 305 -2795
rect 275 -2890 305 -2860
rect 625 -1350 655 -1320
rect 625 -1415 655 -1385
rect 625 -1485 655 -1455
rect 625 -1555 655 -1525
rect 625 -1625 655 -1595
rect 625 -1690 655 -1660
rect 625 -1750 655 -1720
rect 625 -1815 655 -1785
rect 625 -1885 655 -1855
rect 625 -1955 655 -1925
rect 625 -2025 655 -1995
rect 625 -2090 655 -2060
rect 625 -2150 655 -2120
rect 625 -2215 655 -2185
rect 625 -2285 655 -2255
rect 625 -2355 655 -2325
rect 625 -2425 655 -2395
rect 625 -2490 655 -2460
rect 625 -2550 655 -2520
rect 625 -2615 655 -2585
rect 625 -2685 655 -2655
rect 625 -2755 655 -2725
rect 625 -2825 655 -2795
rect 625 -2890 655 -2860
rect 975 -1350 1005 -1320
rect 975 -1415 1005 -1385
rect 975 -1485 1005 -1455
rect 975 -1555 1005 -1525
rect 975 -1625 1005 -1595
rect 975 -1690 1005 -1660
rect 975 -1750 1005 -1720
rect 975 -1815 1005 -1785
rect 975 -1885 1005 -1855
rect 975 -1955 1005 -1925
rect 975 -2025 1005 -1995
rect 975 -2090 1005 -2060
rect 975 -2150 1005 -2120
rect 975 -2215 1005 -2185
rect 975 -2285 1005 -2255
rect 975 -2355 1005 -2325
rect 975 -2425 1005 -2395
rect 975 -2490 1005 -2460
rect 975 -2550 1005 -2520
rect 975 -2615 1005 -2585
rect 975 -2685 1005 -2655
rect 975 -2755 1005 -2725
rect 975 -2825 1005 -2795
rect 975 -2890 1005 -2860
rect 1325 -1350 1355 -1320
rect 1325 -1415 1355 -1385
rect 1325 -1485 1355 -1455
rect 1325 -1555 1355 -1525
rect 1325 -1625 1355 -1595
rect 1325 -1690 1355 -1660
rect 1325 -1750 1355 -1720
rect 1325 -1815 1355 -1785
rect 1325 -1885 1355 -1855
rect 1325 -1955 1355 -1925
rect 1325 -2025 1355 -1995
rect 1325 -2090 1355 -2060
rect 1325 -2150 1355 -2120
rect 1325 -2215 1355 -2185
rect 1325 -2285 1355 -2255
rect 1325 -2355 1355 -2325
rect 1325 -2425 1355 -2395
rect 1325 -2490 1355 -2460
rect 1325 -2550 1355 -2520
rect 1325 -2615 1355 -2585
rect 1325 -2685 1355 -2655
rect 1325 -2755 1355 -2725
rect 1325 -2825 1355 -2795
rect 1325 -2890 1355 -2860
rect 1675 -1350 1705 -1320
rect 1675 -1415 1705 -1385
rect 1675 -1485 1705 -1455
rect 1675 -1555 1705 -1525
rect 1675 -1625 1705 -1595
rect 1675 -1690 1705 -1660
rect 1675 -1750 1705 -1720
rect 1675 -1815 1705 -1785
rect 1675 -1885 1705 -1855
rect 1675 -1955 1705 -1925
rect 1675 -2025 1705 -1995
rect 1675 -2090 1705 -2060
rect 1675 -2150 1705 -2120
rect 1675 -2215 1705 -2185
rect 1675 -2285 1705 -2255
rect 1675 -2355 1705 -2325
rect 1675 -2425 1705 -2395
rect 1675 -2490 1705 -2460
rect 1675 -2550 1705 -2520
rect 1675 -2615 1705 -2585
rect 1675 -2685 1705 -2655
rect 1675 -2755 1705 -2725
rect 1675 -2825 1705 -2795
rect 1675 -2890 1705 -2860
rect 2025 -1350 2055 -1320
rect 2025 -1415 2055 -1385
rect 2025 -1485 2055 -1455
rect 2025 -1555 2055 -1525
rect 2025 -1625 2055 -1595
rect 2025 -1690 2055 -1660
rect 2025 -1750 2055 -1720
rect 2025 -1815 2055 -1785
rect 2025 -1885 2055 -1855
rect 2025 -1955 2055 -1925
rect 2025 -2025 2055 -1995
rect 2025 -2090 2055 -2060
rect 2025 -2150 2055 -2120
rect 2025 -2215 2055 -2185
rect 2025 -2285 2055 -2255
rect 2025 -2355 2055 -2325
rect 2025 -2425 2055 -2395
rect 2025 -2490 2055 -2460
rect 2025 -2550 2055 -2520
rect 2025 -2615 2055 -2585
rect 2025 -2685 2055 -2655
rect 2025 -2755 2055 -2725
rect 2025 -2825 2055 -2795
rect 2025 -2890 2055 -2860
rect 2375 -1350 2405 -1320
rect 2375 -1415 2405 -1385
rect 2375 -1485 2405 -1455
rect 2375 -1555 2405 -1525
rect 2375 -1625 2405 -1595
rect 2375 -1690 2405 -1660
rect 2375 -1750 2405 -1720
rect 2375 -1815 2405 -1785
rect 2375 -1885 2405 -1855
rect 2375 -1955 2405 -1925
rect 2375 -2025 2405 -1995
rect 2375 -2090 2405 -2060
rect 2375 -2150 2405 -2120
rect 2375 -2215 2405 -2185
rect 2375 -2285 2405 -2255
rect 2375 -2355 2405 -2325
rect 2375 -2425 2405 -2395
rect 2375 -2490 2405 -2460
rect 2375 -2550 2405 -2520
rect 2375 -2615 2405 -2585
rect 2375 -2685 2405 -2655
rect 2375 -2755 2405 -2725
rect 2375 -2825 2405 -2795
rect 2375 -2890 2405 -2860
rect 2725 -1350 2755 -1320
rect 2725 -1415 2755 -1385
rect 2725 -1485 2755 -1455
rect 2725 -1555 2755 -1525
rect 2725 -1625 2755 -1595
rect 2725 -1690 2755 -1660
rect 2725 -1750 2755 -1720
rect 2725 -1815 2755 -1785
rect 2725 -1885 2755 -1855
rect 2725 -1955 2755 -1925
rect 2725 -2025 2755 -1995
rect 2725 -2090 2755 -2060
rect 2725 -2150 2755 -2120
rect 2725 -2215 2755 -2185
rect 2725 -2285 2755 -2255
rect 2725 -2355 2755 -2325
rect 2725 -2425 2755 -2395
rect 2725 -2490 2755 -2460
rect 2725 -2550 2755 -2520
rect 2725 -2615 2755 -2585
rect 2725 -2685 2755 -2655
rect 2725 -2755 2755 -2725
rect 2725 -2825 2755 -2795
rect 2725 -2890 2755 -2860
rect 3075 -1350 3105 -1320
rect 3075 -1415 3105 -1385
rect 3075 -1485 3105 -1455
rect 3075 -1555 3105 -1525
rect 3075 -1625 3105 -1595
rect 3075 -1690 3105 -1660
rect 3075 -1750 3105 -1720
rect 3075 -1815 3105 -1785
rect 3075 -1885 3105 -1855
rect 3075 -1955 3105 -1925
rect 3075 -2025 3105 -1995
rect 3075 -2090 3105 -2060
rect 3075 -2150 3105 -2120
rect 3075 -2215 3105 -2185
rect 3075 -2285 3105 -2255
rect 3075 -2355 3105 -2325
rect 3075 -2425 3105 -2395
rect 3075 -2490 3105 -2460
rect 3075 -2550 3105 -2520
rect 3075 -2615 3105 -2585
rect 3075 -2685 3105 -2655
rect 3075 -2755 3105 -2725
rect 3075 -2825 3105 -2795
rect 3075 -2890 3105 -2860
rect 5875 -1350 5905 -1320
rect 5875 -1415 5905 -1385
rect 5875 -1485 5905 -1455
rect 5875 -1555 5905 -1525
rect 5875 -1625 5905 -1595
rect 5875 -1690 5905 -1660
rect 5875 -1750 5905 -1720
rect 5875 -1815 5905 -1785
rect 5875 -1885 5905 -1855
rect 5875 -1955 5905 -1925
rect 5875 -2025 5905 -1995
rect 5875 -2090 5905 -2060
rect 5875 -2150 5905 -2120
rect 5875 -2215 5905 -2185
rect 5875 -2285 5905 -2255
rect 5875 -2355 5905 -2325
rect 5875 -2425 5905 -2395
rect 5875 -2490 5905 -2460
rect 5875 -2550 5905 -2520
rect 5875 -2615 5905 -2585
rect 5875 -2685 5905 -2655
rect 5875 -2755 5905 -2725
rect 5875 -2825 5905 -2795
rect 5875 -2890 5905 -2860
rect 6225 -1350 6255 -1320
rect 6225 -1415 6255 -1385
rect 6225 -1485 6255 -1455
rect 6225 -1555 6255 -1525
rect 6225 -1625 6255 -1595
rect 6225 -1690 6255 -1660
rect 6225 -1750 6255 -1720
rect 6225 -1815 6255 -1785
rect 6225 -1885 6255 -1855
rect 6225 -1955 6255 -1925
rect 6225 -2025 6255 -1995
rect 6225 -2090 6255 -2060
rect 6225 -2150 6255 -2120
rect 6225 -2215 6255 -2185
rect 6225 -2285 6255 -2255
rect 6225 -2355 6255 -2325
rect 6225 -2425 6255 -2395
rect 6225 -2490 6255 -2460
rect 6225 -2550 6255 -2520
rect 6225 -2615 6255 -2585
rect 6225 -2685 6255 -2655
rect 6225 -2755 6255 -2725
rect 6225 -2825 6255 -2795
rect 6225 -2890 6255 -2860
rect 6575 -1350 6605 -1320
rect 6575 -1415 6605 -1385
rect 6575 -1485 6605 -1455
rect 6575 -1555 6605 -1525
rect 6575 -1625 6605 -1595
rect 6575 -1690 6605 -1660
rect 6575 -1750 6605 -1720
rect 6575 -1815 6605 -1785
rect 6575 -1885 6605 -1855
rect 6575 -1955 6605 -1925
rect 6575 -2025 6605 -1995
rect 6575 -2090 6605 -2060
rect 6575 -2150 6605 -2120
rect 6575 -2215 6605 -2185
rect 6575 -2285 6605 -2255
rect 6575 -2355 6605 -2325
rect 6575 -2425 6605 -2395
rect 6575 -2490 6605 -2460
rect 6575 -2550 6605 -2520
rect 6575 -2615 6605 -2585
rect 6575 -2685 6605 -2655
rect 6575 -2755 6605 -2725
rect 6575 -2825 6605 -2795
rect 6575 -2890 6605 -2860
rect 6925 -1350 6955 -1320
rect 6925 -1415 6955 -1385
rect 6925 -1485 6955 -1455
rect 6925 -1555 6955 -1525
rect 6925 -1625 6955 -1595
rect 6925 -1690 6955 -1660
rect 6925 -1750 6955 -1720
rect 6925 -1815 6955 -1785
rect 6925 -1885 6955 -1855
rect 6925 -1955 6955 -1925
rect 6925 -2025 6955 -1995
rect 6925 -2090 6955 -2060
rect 6925 -2150 6955 -2120
rect 6925 -2215 6955 -2185
rect 6925 -2285 6955 -2255
rect 6925 -2355 6955 -2325
rect 6925 -2425 6955 -2395
rect 6925 -2490 6955 -2460
rect 6925 -2550 6955 -2520
rect 6925 -2615 6955 -2585
rect 6925 -2685 6955 -2655
rect 6925 -2755 6955 -2725
rect 6925 -2825 6955 -2795
rect 6925 -2890 6955 -2860
rect 7275 -1350 7305 -1320
rect 7275 -1415 7305 -1385
rect 7275 -1485 7305 -1455
rect 7275 -1555 7305 -1525
rect 7275 -1625 7305 -1595
rect 7275 -1690 7305 -1660
rect 7275 -1750 7305 -1720
rect 7275 -1815 7305 -1785
rect 7275 -1885 7305 -1855
rect 7275 -1955 7305 -1925
rect 7275 -2025 7305 -1995
rect 7275 -2090 7305 -2060
rect 7275 -2150 7305 -2120
rect 7275 -2215 7305 -2185
rect 7275 -2285 7305 -2255
rect 7275 -2355 7305 -2325
rect 7275 -2425 7305 -2395
rect 7275 -2490 7305 -2460
rect 7275 -2550 7305 -2520
rect 7275 -2615 7305 -2585
rect 7275 -2685 7305 -2655
rect 7275 -2755 7305 -2725
rect 7275 -2825 7305 -2795
rect 7275 -2890 7305 -2860
rect 7625 -1350 7655 -1320
rect 7625 -1415 7655 -1385
rect 7625 -1485 7655 -1455
rect 7625 -1555 7655 -1525
rect 7625 -1625 7655 -1595
rect 7625 -1690 7655 -1660
rect 7625 -1750 7655 -1720
rect 7625 -1815 7655 -1785
rect 7625 -1885 7655 -1855
rect 7625 -1955 7655 -1925
rect 7625 -2025 7655 -1995
rect 7625 -2090 7655 -2060
rect 7625 -2150 7655 -2120
rect 7625 -2215 7655 -2185
rect 7625 -2285 7655 -2255
rect 7625 -2355 7655 -2325
rect 7625 -2425 7655 -2395
rect 7625 -2490 7655 -2460
rect 7625 -2550 7655 -2520
rect 7625 -2615 7655 -2585
rect 7625 -2685 7655 -2655
rect 7625 -2755 7655 -2725
rect 7625 -2825 7655 -2795
rect 7625 -2890 7655 -2860
rect 7975 -1350 8005 -1320
rect 7975 -1415 8005 -1385
rect 7975 -1485 8005 -1455
rect 7975 -1555 8005 -1525
rect 7975 -1625 8005 -1595
rect 7975 -1690 8005 -1660
rect 7975 -1750 8005 -1720
rect 7975 -1815 8005 -1785
rect 7975 -1885 8005 -1855
rect 7975 -1955 8005 -1925
rect 7975 -2025 8005 -1995
rect 7975 -2090 8005 -2060
rect 7975 -2150 8005 -2120
rect 7975 -2215 8005 -2185
rect 7975 -2285 8005 -2255
rect 7975 -2355 8005 -2325
rect 7975 -2425 8005 -2395
rect 7975 -2490 8005 -2460
rect 7975 -2550 8005 -2520
rect 7975 -2615 8005 -2585
rect 7975 -2685 8005 -2655
rect 7975 -2755 8005 -2725
rect 7975 -2825 8005 -2795
rect 7975 -2890 8005 -2860
rect 8325 -1350 8355 -1320
rect 8325 -1415 8355 -1385
rect 8325 -1485 8355 -1455
rect 8325 -1555 8355 -1525
rect 8325 -1625 8355 -1595
rect 8325 -1690 8355 -1660
rect 8325 -1750 8355 -1720
rect 8325 -1815 8355 -1785
rect 8325 -1885 8355 -1855
rect 8325 -1955 8355 -1925
rect 8325 -2025 8355 -1995
rect 8325 -2090 8355 -2060
rect 8325 -2150 8355 -2120
rect 8325 -2215 8355 -2185
rect 8325 -2285 8355 -2255
rect 8325 -2355 8355 -2325
rect 8325 -2425 8355 -2395
rect 8325 -2490 8355 -2460
rect 8325 -2550 8355 -2520
rect 8325 -2615 8355 -2585
rect 8325 -2685 8355 -2655
rect 8325 -2755 8355 -2725
rect 8325 -2825 8355 -2795
rect 8325 -2890 8355 -2860
rect 8675 -1350 8705 -1320
rect 8675 -1415 8705 -1385
rect 8675 -1485 8705 -1455
rect 8675 -1555 8705 -1525
rect 8675 -1625 8705 -1595
rect 8675 -1690 8705 -1660
rect 8675 -1750 8705 -1720
rect 8675 -1815 8705 -1785
rect 8675 -1885 8705 -1855
rect 8675 -1955 8705 -1925
rect 8675 -2025 8705 -1995
rect 8675 -2090 8705 -2060
rect 8675 -2150 8705 -2120
rect 8675 -2215 8705 -2185
rect 8675 -2285 8705 -2255
rect 8675 -2355 8705 -2325
rect 8675 -2425 8705 -2395
rect 8675 -2490 8705 -2460
rect 8675 -2550 8705 -2520
rect 8675 -2615 8705 -2585
rect 8675 -2685 8705 -2655
rect 8675 -2755 8705 -2725
rect 8675 -2825 8705 -2795
rect 8675 -2890 8705 -2860
rect 9025 -1350 9055 -1320
rect 9025 -1415 9055 -1385
rect 9025 -1485 9055 -1455
rect 9025 -1555 9055 -1525
rect 9025 -1625 9055 -1595
rect 9025 -1690 9055 -1660
rect 9025 -1750 9055 -1720
rect 9025 -1815 9055 -1785
rect 9025 -1885 9055 -1855
rect 9025 -1955 9055 -1925
rect 9025 -2025 9055 -1995
rect 9025 -2090 9055 -2060
rect 9025 -2150 9055 -2120
rect 9025 -2215 9055 -2185
rect 9025 -2285 9055 -2255
rect 9025 -2355 9055 -2325
rect 9025 -2425 9055 -2395
rect 9025 -2490 9055 -2460
rect 9025 -2550 9055 -2520
rect 9025 -2615 9055 -2585
rect 9025 -2685 9055 -2655
rect 9025 -2755 9055 -2725
rect 9025 -2825 9055 -2795
rect 9025 -2890 9055 -2860
rect 3425 -3050 3455 -3020
rect 3425 -3115 3455 -3085
rect 3425 -3185 3455 -3155
rect 3425 -3255 3455 -3225
rect 3425 -3325 3455 -3295
rect 3425 -3390 3455 -3360
rect 3425 -3450 3455 -3420
rect 3425 -3515 3455 -3485
rect 3425 -3585 3455 -3555
rect 3425 -3655 3455 -3625
rect 3425 -3725 3455 -3695
rect 3425 -3790 3455 -3760
rect 3425 -3850 3455 -3820
rect 3425 -3915 3455 -3885
rect 3425 -3985 3455 -3955
rect 3425 -4055 3455 -4025
rect 3425 -4125 3455 -4095
rect 3425 -4190 3455 -4160
rect 3425 -4250 3455 -4220
rect 3425 -4315 3455 -4285
rect 3425 -4385 3455 -4355
rect 3425 -4455 3455 -4425
rect 3425 -4525 3455 -4495
rect 3425 -4590 3455 -4560
rect 3775 -3050 3805 -3020
rect 3775 -3115 3805 -3085
rect 3775 -3185 3805 -3155
rect 3775 -3255 3805 -3225
rect 3775 -3325 3805 -3295
rect 3775 -3390 3805 -3360
rect 3775 -3450 3805 -3420
rect 3775 -3515 3805 -3485
rect 3775 -3585 3805 -3555
rect 3775 -3655 3805 -3625
rect 3775 -3725 3805 -3695
rect 3775 -3790 3805 -3760
rect 3775 -3850 3805 -3820
rect 3775 -3915 3805 -3885
rect 3775 -3985 3805 -3955
rect 3775 -4055 3805 -4025
rect 3775 -4125 3805 -4095
rect 3775 -4190 3805 -4160
rect 3775 -4250 3805 -4220
rect 3775 -4315 3805 -4285
rect 3775 -4385 3805 -4355
rect 3775 -4455 3805 -4425
rect 3775 -4525 3805 -4495
rect 3775 -4590 3805 -4560
rect 4125 -3050 4155 -3020
rect 4125 -3115 4155 -3085
rect 4125 -3185 4155 -3155
rect 4125 -3255 4155 -3225
rect 4125 -3325 4155 -3295
rect 4125 -3390 4155 -3360
rect 4125 -3450 4155 -3420
rect 4125 -3515 4155 -3485
rect 4125 -3585 4155 -3555
rect 4125 -3655 4155 -3625
rect 4125 -3725 4155 -3695
rect 4125 -3790 4155 -3760
rect 4125 -3850 4155 -3820
rect 4125 -3915 4155 -3885
rect 4125 -3985 4155 -3955
rect 4125 -4055 4155 -4025
rect 4125 -4125 4155 -4095
rect 4125 -4190 4155 -4160
rect 4125 -4250 4155 -4220
rect 4125 -4315 4155 -4285
rect 4125 -4385 4155 -4355
rect 4125 -4455 4155 -4425
rect 4125 -4525 4155 -4495
rect 4125 -4590 4155 -4560
rect 4475 -3050 4505 -3020
rect 4475 -3115 4505 -3085
rect 4475 -3185 4505 -3155
rect 4475 -3255 4505 -3225
rect 4475 -3325 4505 -3295
rect 4475 -3390 4505 -3360
rect 4475 -3450 4505 -3420
rect 4475 -3515 4505 -3485
rect 4475 -3585 4505 -3555
rect 4475 -3655 4505 -3625
rect 4475 -3725 4505 -3695
rect 4475 -3790 4505 -3760
rect 4475 -3850 4505 -3820
rect 4475 -3915 4505 -3885
rect 4475 -3985 4505 -3955
rect 4475 -4055 4505 -4025
rect 4475 -4125 4505 -4095
rect 4475 -4190 4505 -4160
rect 4475 -4250 4505 -4220
rect 4475 -4315 4505 -4285
rect 4475 -4385 4505 -4355
rect 4475 -4455 4505 -4425
rect 4475 -4525 4505 -4495
rect 4475 -4590 4505 -4560
rect 4825 -3050 4855 -3020
rect 4825 -3115 4855 -3085
rect 4825 -3185 4855 -3155
rect 4825 -3255 4855 -3225
rect 4825 -3325 4855 -3295
rect 4825 -3390 4855 -3360
rect 4825 -3450 4855 -3420
rect 4825 -3515 4855 -3485
rect 4825 -3585 4855 -3555
rect 4825 -3655 4855 -3625
rect 4825 -3725 4855 -3695
rect 4825 -3790 4855 -3760
rect 4825 -3850 4855 -3820
rect 4825 -3915 4855 -3885
rect 4825 -3985 4855 -3955
rect 4825 -4055 4855 -4025
rect 4825 -4125 4855 -4095
rect 4825 -4190 4855 -4160
rect 4825 -4250 4855 -4220
rect 4825 -4315 4855 -4285
rect 4825 -4385 4855 -4355
rect 4825 -4455 4855 -4425
rect 4825 -4525 4855 -4495
rect 4825 -4590 4855 -4560
rect 5175 -3050 5205 -3020
rect 5175 -3115 5205 -3085
rect 5175 -3185 5205 -3155
rect 5175 -3255 5205 -3225
rect 5175 -3325 5205 -3295
rect 5175 -3390 5205 -3360
rect 5175 -3450 5205 -3420
rect 5175 -3515 5205 -3485
rect 5175 -3585 5205 -3555
rect 5175 -3655 5205 -3625
rect 5175 -3725 5205 -3695
rect 5175 -3790 5205 -3760
rect 5175 -3850 5205 -3820
rect 5175 -3915 5205 -3885
rect 5175 -3985 5205 -3955
rect 5175 -4055 5205 -4025
rect 5175 -4125 5205 -4095
rect 5175 -4190 5205 -4160
rect 5175 -4250 5205 -4220
rect 5175 -4315 5205 -4285
rect 5175 -4385 5205 -4355
rect 5175 -4455 5205 -4425
rect 5175 -4525 5205 -4495
rect 5175 -4590 5205 -4560
rect 5525 -3050 5555 -3020
rect 5525 -3115 5555 -3085
rect 5525 -3185 5555 -3155
rect 5525 -3255 5555 -3225
rect 5525 -3325 5555 -3295
rect 5525 -3390 5555 -3360
rect 5525 -3450 5555 -3420
rect 5525 -3515 5555 -3485
rect 5525 -3585 5555 -3555
rect 5525 -3655 5555 -3625
rect 5525 -3725 5555 -3695
rect 5525 -3790 5555 -3760
rect 5525 -3850 5555 -3820
rect 5525 -3915 5555 -3885
rect 5525 -3985 5555 -3955
rect 5525 -4055 5555 -4025
rect 5525 -4125 5555 -4095
rect 5525 -4190 5555 -4160
rect 5525 -4250 5555 -4220
rect 5525 -4315 5555 -4285
rect 5525 -4385 5555 -4355
rect 5525 -4455 5555 -4425
rect 5525 -4525 5555 -4495
rect 5525 -4590 5555 -4560
<< metal3 >>
rect 2100 19315 2160 19325
rect 2100 19275 2110 19315
rect 2150 19275 2160 19315
rect 2100 19250 2160 19275
rect 2100 19210 2110 19250
rect 2150 19210 2160 19250
rect 2100 19180 2160 19210
rect 2100 19140 2110 19180
rect 2150 19140 2160 19180
rect 2100 19110 2160 19140
rect 2100 19070 2110 19110
rect 2150 19070 2160 19110
rect 2100 19040 2160 19070
rect 2100 19000 2110 19040
rect 2150 19000 2160 19040
rect 2100 18975 2160 19000
rect 2100 18935 2110 18975
rect 2150 18935 2160 18975
rect 2100 18915 2160 18935
rect 2100 18875 2110 18915
rect 2150 18875 2160 18915
rect 2100 18850 2160 18875
rect 2100 18810 2110 18850
rect 2150 18810 2160 18850
rect 2100 18780 2160 18810
rect 2100 18740 2110 18780
rect 2150 18740 2160 18780
rect 2100 18710 2160 18740
rect 2100 18670 2110 18710
rect 2150 18670 2160 18710
rect 2100 18640 2160 18670
rect 2100 18600 2110 18640
rect 2150 18600 2160 18640
rect 2100 18575 2160 18600
rect 2100 18535 2110 18575
rect 2150 18535 2160 18575
rect 2100 18515 2160 18535
rect 2100 18475 2110 18515
rect 2150 18475 2160 18515
rect 2100 18450 2160 18475
rect 2100 18410 2110 18450
rect 2150 18410 2160 18450
rect 2100 18380 2160 18410
rect 2100 18340 2110 18380
rect 2150 18340 2160 18380
rect 2100 18310 2160 18340
rect 2100 18270 2110 18310
rect 2150 18270 2160 18310
rect 2100 18240 2160 18270
rect 2100 18200 2110 18240
rect 2150 18200 2160 18240
rect 2100 18175 2160 18200
rect 2100 18135 2110 18175
rect 2150 18135 2160 18175
rect 2100 18115 2160 18135
rect 2100 18075 2110 18115
rect 2150 18075 2160 18115
rect 2100 18050 2160 18075
rect 2100 18010 2110 18050
rect 2150 18010 2160 18050
rect 2100 17980 2160 18010
rect 2100 17940 2110 17980
rect 2150 17940 2160 17980
rect 2100 17910 2160 17940
rect 2100 17870 2110 17910
rect 2150 17870 2160 17910
rect 2100 17840 2160 17870
rect 2100 17800 2110 17840
rect 2150 17800 2160 17840
rect 2100 17775 2160 17800
rect 2100 17735 2110 17775
rect 2150 17735 2160 17775
rect 2100 17725 2160 17735
rect 6690 19315 6750 19325
rect 6690 19275 6700 19315
rect 6740 19275 6750 19315
rect 6690 19250 6750 19275
rect 6690 19210 6700 19250
rect 6740 19210 6750 19250
rect 6690 19180 6750 19210
rect 6690 19140 6700 19180
rect 6740 19140 6750 19180
rect 6690 19110 6750 19140
rect 6690 19070 6700 19110
rect 6740 19070 6750 19110
rect 6690 19040 6750 19070
rect 6690 19000 6700 19040
rect 6740 19000 6750 19040
rect 6690 18975 6750 19000
rect 6690 18935 6700 18975
rect 6740 18935 6750 18975
rect 6690 18915 6750 18935
rect 6690 18875 6700 18915
rect 6740 18875 6750 18915
rect 6690 18850 6750 18875
rect 6690 18810 6700 18850
rect 6740 18810 6750 18850
rect 6690 18780 6750 18810
rect 6690 18740 6700 18780
rect 6740 18740 6750 18780
rect 6690 18710 6750 18740
rect 6690 18670 6700 18710
rect 6740 18670 6750 18710
rect 6690 18640 6750 18670
rect 6690 18600 6700 18640
rect 6740 18600 6750 18640
rect 6690 18575 6750 18600
rect 6690 18535 6700 18575
rect 6740 18535 6750 18575
rect 6690 18515 6750 18535
rect 6690 18475 6700 18515
rect 6740 18475 6750 18515
rect 6690 18450 6750 18475
rect 6690 18410 6700 18450
rect 6740 18410 6750 18450
rect 6690 18380 6750 18410
rect 6690 18340 6700 18380
rect 6740 18340 6750 18380
rect 6690 18310 6750 18340
rect 6690 18270 6700 18310
rect 6740 18270 6750 18310
rect 6690 18240 6750 18270
rect 6690 18200 6700 18240
rect 6740 18200 6750 18240
rect 6690 18175 6750 18200
rect 6690 18135 6700 18175
rect 6740 18135 6750 18175
rect 6690 18115 6750 18135
rect 6690 18075 6700 18115
rect 6740 18075 6750 18115
rect 6690 18050 6750 18075
rect 6690 18010 6700 18050
rect 6740 18010 6750 18050
rect 6690 17980 6750 18010
rect 6690 17940 6700 17980
rect 6740 17940 6750 17980
rect 6690 17910 6750 17940
rect 6690 17870 6700 17910
rect 6740 17870 6750 17910
rect 6690 17840 6750 17870
rect 6690 17800 6700 17840
rect 6740 17800 6750 17840
rect 6690 17775 6750 17800
rect 6690 17735 6700 17775
rect 6740 17735 6750 17775
rect 6690 17725 6750 17735
rect 31290 19305 32890 19325
rect 31290 19270 31305 19305
rect 31340 19270 31350 19305
rect 31385 19270 31395 19305
rect 31430 19270 31440 19305
rect 31475 19270 31485 19305
rect 31520 19270 31530 19305
rect 31565 19270 31575 19305
rect 31610 19270 31620 19305
rect 31655 19270 31665 19305
rect 31700 19270 31710 19305
rect 31745 19270 31755 19305
rect 31790 19270 31800 19305
rect 31835 19270 31845 19305
rect 31880 19270 31890 19305
rect 31925 19270 31935 19305
rect 31970 19270 31980 19305
rect 32015 19270 32025 19305
rect 32060 19270 32070 19305
rect 32105 19270 32115 19305
rect 32150 19270 32160 19305
rect 32195 19270 32205 19305
rect 32240 19270 32250 19305
rect 32285 19270 32295 19305
rect 32330 19270 32340 19305
rect 32375 19270 32385 19305
rect 32420 19270 32430 19305
rect 32465 19270 32475 19305
rect 32510 19270 32520 19305
rect 32555 19270 32565 19305
rect 32600 19270 32610 19305
rect 32645 19270 32655 19305
rect 32690 19270 32700 19305
rect 32735 19270 32745 19305
rect 32780 19270 32790 19305
rect 32825 19270 32835 19305
rect 32870 19270 32890 19305
rect 31290 19260 32890 19270
rect 31290 19225 31305 19260
rect 31340 19225 31350 19260
rect 31385 19225 31395 19260
rect 31430 19225 31440 19260
rect 31475 19225 31485 19260
rect 31520 19225 31530 19260
rect 31565 19225 31575 19260
rect 31610 19225 31620 19260
rect 31655 19225 31665 19260
rect 31700 19225 31710 19260
rect 31745 19225 31755 19260
rect 31790 19225 31800 19260
rect 31835 19225 31845 19260
rect 31880 19225 31890 19260
rect 31925 19225 31935 19260
rect 31970 19225 31980 19260
rect 32015 19225 32025 19260
rect 32060 19225 32070 19260
rect 32105 19225 32115 19260
rect 32150 19225 32160 19260
rect 32195 19225 32205 19260
rect 32240 19225 32250 19260
rect 32285 19225 32295 19260
rect 32330 19225 32340 19260
rect 32375 19225 32385 19260
rect 32420 19225 32430 19260
rect 32465 19225 32475 19260
rect 32510 19225 32520 19260
rect 32555 19225 32565 19260
rect 32600 19225 32610 19260
rect 32645 19225 32655 19260
rect 32690 19225 32700 19260
rect 32735 19225 32745 19260
rect 32780 19225 32790 19260
rect 32825 19225 32835 19260
rect 32870 19225 32890 19260
rect 31290 19215 32890 19225
rect 31290 19180 31305 19215
rect 31340 19180 31350 19215
rect 31385 19180 31395 19215
rect 31430 19180 31440 19215
rect 31475 19180 31485 19215
rect 31520 19180 31530 19215
rect 31565 19180 31575 19215
rect 31610 19180 31620 19215
rect 31655 19180 31665 19215
rect 31700 19180 31710 19215
rect 31745 19180 31755 19215
rect 31790 19180 31800 19215
rect 31835 19180 31845 19215
rect 31880 19180 31890 19215
rect 31925 19180 31935 19215
rect 31970 19180 31980 19215
rect 32015 19180 32025 19215
rect 32060 19180 32070 19215
rect 32105 19180 32115 19215
rect 32150 19180 32160 19215
rect 32195 19180 32205 19215
rect 32240 19180 32250 19215
rect 32285 19180 32295 19215
rect 32330 19180 32340 19215
rect 32375 19180 32385 19215
rect 32420 19180 32430 19215
rect 32465 19180 32475 19215
rect 32510 19180 32520 19215
rect 32555 19180 32565 19215
rect 32600 19180 32610 19215
rect 32645 19180 32655 19215
rect 32690 19180 32700 19215
rect 32735 19180 32745 19215
rect 32780 19180 32790 19215
rect 32825 19180 32835 19215
rect 32870 19180 32890 19215
rect 31290 19170 32890 19180
rect 31290 19135 31305 19170
rect 31340 19135 31350 19170
rect 31385 19135 31395 19170
rect 31430 19135 31440 19170
rect 31475 19135 31485 19170
rect 31520 19135 31530 19170
rect 31565 19135 31575 19170
rect 31610 19135 31620 19170
rect 31655 19135 31665 19170
rect 31700 19135 31710 19170
rect 31745 19135 31755 19170
rect 31790 19135 31800 19170
rect 31835 19135 31845 19170
rect 31880 19135 31890 19170
rect 31925 19135 31935 19170
rect 31970 19135 31980 19170
rect 32015 19135 32025 19170
rect 32060 19135 32070 19170
rect 32105 19135 32115 19170
rect 32150 19135 32160 19170
rect 32195 19135 32205 19170
rect 32240 19135 32250 19170
rect 32285 19135 32295 19170
rect 32330 19135 32340 19170
rect 32375 19135 32385 19170
rect 32420 19135 32430 19170
rect 32465 19135 32475 19170
rect 32510 19135 32520 19170
rect 32555 19135 32565 19170
rect 32600 19135 32610 19170
rect 32645 19135 32655 19170
rect 32690 19135 32700 19170
rect 32735 19135 32745 19170
rect 32780 19135 32790 19170
rect 32825 19135 32835 19170
rect 32870 19135 32890 19170
rect 31290 19125 32890 19135
rect 31290 19090 31305 19125
rect 31340 19090 31350 19125
rect 31385 19090 31395 19125
rect 31430 19090 31440 19125
rect 31475 19090 31485 19125
rect 31520 19090 31530 19125
rect 31565 19090 31575 19125
rect 31610 19090 31620 19125
rect 31655 19090 31665 19125
rect 31700 19090 31710 19125
rect 31745 19090 31755 19125
rect 31790 19090 31800 19125
rect 31835 19090 31845 19125
rect 31880 19090 31890 19125
rect 31925 19090 31935 19125
rect 31970 19090 31980 19125
rect 32015 19090 32025 19125
rect 32060 19090 32070 19125
rect 32105 19090 32115 19125
rect 32150 19090 32160 19125
rect 32195 19090 32205 19125
rect 32240 19090 32250 19125
rect 32285 19090 32295 19125
rect 32330 19090 32340 19125
rect 32375 19090 32385 19125
rect 32420 19090 32430 19125
rect 32465 19090 32475 19125
rect 32510 19090 32520 19125
rect 32555 19090 32565 19125
rect 32600 19090 32610 19125
rect 32645 19090 32655 19125
rect 32690 19090 32700 19125
rect 32735 19090 32745 19125
rect 32780 19090 32790 19125
rect 32825 19090 32835 19125
rect 32870 19090 32890 19125
rect 31290 19080 32890 19090
rect 31290 19045 31305 19080
rect 31340 19045 31350 19080
rect 31385 19045 31395 19080
rect 31430 19045 31440 19080
rect 31475 19045 31485 19080
rect 31520 19045 31530 19080
rect 31565 19045 31575 19080
rect 31610 19045 31620 19080
rect 31655 19045 31665 19080
rect 31700 19045 31710 19080
rect 31745 19045 31755 19080
rect 31790 19045 31800 19080
rect 31835 19045 31845 19080
rect 31880 19045 31890 19080
rect 31925 19045 31935 19080
rect 31970 19045 31980 19080
rect 32015 19045 32025 19080
rect 32060 19045 32070 19080
rect 32105 19045 32115 19080
rect 32150 19045 32160 19080
rect 32195 19045 32205 19080
rect 32240 19045 32250 19080
rect 32285 19045 32295 19080
rect 32330 19045 32340 19080
rect 32375 19045 32385 19080
rect 32420 19045 32430 19080
rect 32465 19045 32475 19080
rect 32510 19045 32520 19080
rect 32555 19045 32565 19080
rect 32600 19045 32610 19080
rect 32645 19045 32655 19080
rect 32690 19045 32700 19080
rect 32735 19045 32745 19080
rect 32780 19045 32790 19080
rect 32825 19045 32835 19080
rect 32870 19045 32890 19080
rect 31290 19035 32890 19045
rect 31290 19000 31305 19035
rect 31340 19000 31350 19035
rect 31385 19000 31395 19035
rect 31430 19000 31440 19035
rect 31475 19000 31485 19035
rect 31520 19000 31530 19035
rect 31565 19000 31575 19035
rect 31610 19000 31620 19035
rect 31655 19000 31665 19035
rect 31700 19000 31710 19035
rect 31745 19000 31755 19035
rect 31790 19000 31800 19035
rect 31835 19000 31845 19035
rect 31880 19000 31890 19035
rect 31925 19000 31935 19035
rect 31970 19000 31980 19035
rect 32015 19000 32025 19035
rect 32060 19000 32070 19035
rect 32105 19000 32115 19035
rect 32150 19000 32160 19035
rect 32195 19000 32205 19035
rect 32240 19000 32250 19035
rect 32285 19000 32295 19035
rect 32330 19000 32340 19035
rect 32375 19000 32385 19035
rect 32420 19000 32430 19035
rect 32465 19000 32475 19035
rect 32510 19000 32520 19035
rect 32555 19000 32565 19035
rect 32600 19000 32610 19035
rect 32645 19000 32655 19035
rect 32690 19000 32700 19035
rect 32735 19000 32745 19035
rect 32780 19000 32790 19035
rect 32825 19000 32835 19035
rect 32870 19000 32890 19035
rect 31290 18990 32890 19000
rect 31290 18955 31305 18990
rect 31340 18955 31350 18990
rect 31385 18955 31395 18990
rect 31430 18955 31440 18990
rect 31475 18955 31485 18990
rect 31520 18955 31530 18990
rect 31565 18955 31575 18990
rect 31610 18955 31620 18990
rect 31655 18955 31665 18990
rect 31700 18955 31710 18990
rect 31745 18955 31755 18990
rect 31790 18955 31800 18990
rect 31835 18955 31845 18990
rect 31880 18955 31890 18990
rect 31925 18955 31935 18990
rect 31970 18955 31980 18990
rect 32015 18955 32025 18990
rect 32060 18955 32070 18990
rect 32105 18955 32115 18990
rect 32150 18955 32160 18990
rect 32195 18955 32205 18990
rect 32240 18955 32250 18990
rect 32285 18955 32295 18990
rect 32330 18955 32340 18990
rect 32375 18955 32385 18990
rect 32420 18955 32430 18990
rect 32465 18955 32475 18990
rect 32510 18955 32520 18990
rect 32555 18955 32565 18990
rect 32600 18955 32610 18990
rect 32645 18955 32655 18990
rect 32690 18955 32700 18990
rect 32735 18955 32745 18990
rect 32780 18955 32790 18990
rect 32825 18955 32835 18990
rect 32870 18955 32890 18990
rect 31290 18945 32890 18955
rect 31290 18910 31305 18945
rect 31340 18910 31350 18945
rect 31385 18910 31395 18945
rect 31430 18910 31440 18945
rect 31475 18910 31485 18945
rect 31520 18910 31530 18945
rect 31565 18910 31575 18945
rect 31610 18910 31620 18945
rect 31655 18910 31665 18945
rect 31700 18910 31710 18945
rect 31745 18910 31755 18945
rect 31790 18910 31800 18945
rect 31835 18910 31845 18945
rect 31880 18910 31890 18945
rect 31925 18910 31935 18945
rect 31970 18910 31980 18945
rect 32015 18910 32025 18945
rect 32060 18910 32070 18945
rect 32105 18910 32115 18945
rect 32150 18910 32160 18945
rect 32195 18910 32205 18945
rect 32240 18910 32250 18945
rect 32285 18910 32295 18945
rect 32330 18910 32340 18945
rect 32375 18910 32385 18945
rect 32420 18910 32430 18945
rect 32465 18910 32475 18945
rect 32510 18910 32520 18945
rect 32555 18910 32565 18945
rect 32600 18910 32610 18945
rect 32645 18910 32655 18945
rect 32690 18910 32700 18945
rect 32735 18910 32745 18945
rect 32780 18910 32790 18945
rect 32825 18910 32835 18945
rect 32870 18910 32890 18945
rect 31290 18900 32890 18910
rect 31290 18865 31305 18900
rect 31340 18865 31350 18900
rect 31385 18865 31395 18900
rect 31430 18865 31440 18900
rect 31475 18865 31485 18900
rect 31520 18865 31530 18900
rect 31565 18865 31575 18900
rect 31610 18865 31620 18900
rect 31655 18865 31665 18900
rect 31700 18865 31710 18900
rect 31745 18865 31755 18900
rect 31790 18865 31800 18900
rect 31835 18865 31845 18900
rect 31880 18865 31890 18900
rect 31925 18865 31935 18900
rect 31970 18865 31980 18900
rect 32015 18865 32025 18900
rect 32060 18865 32070 18900
rect 32105 18865 32115 18900
rect 32150 18865 32160 18900
rect 32195 18865 32205 18900
rect 32240 18865 32250 18900
rect 32285 18865 32295 18900
rect 32330 18865 32340 18900
rect 32375 18865 32385 18900
rect 32420 18865 32430 18900
rect 32465 18865 32475 18900
rect 32510 18865 32520 18900
rect 32555 18865 32565 18900
rect 32600 18865 32610 18900
rect 32645 18865 32655 18900
rect 32690 18865 32700 18900
rect 32735 18865 32745 18900
rect 32780 18865 32790 18900
rect 32825 18865 32835 18900
rect 32870 18865 32890 18900
rect 31290 18855 32890 18865
rect 31290 18820 31305 18855
rect 31340 18820 31350 18855
rect 31385 18820 31395 18855
rect 31430 18820 31440 18855
rect 31475 18820 31485 18855
rect 31520 18820 31530 18855
rect 31565 18820 31575 18855
rect 31610 18820 31620 18855
rect 31655 18820 31665 18855
rect 31700 18820 31710 18855
rect 31745 18820 31755 18855
rect 31790 18820 31800 18855
rect 31835 18820 31845 18855
rect 31880 18820 31890 18855
rect 31925 18820 31935 18855
rect 31970 18820 31980 18855
rect 32015 18820 32025 18855
rect 32060 18820 32070 18855
rect 32105 18820 32115 18855
rect 32150 18820 32160 18855
rect 32195 18820 32205 18855
rect 32240 18820 32250 18855
rect 32285 18820 32295 18855
rect 32330 18820 32340 18855
rect 32375 18820 32385 18855
rect 32420 18820 32430 18855
rect 32465 18820 32475 18855
rect 32510 18820 32520 18855
rect 32555 18820 32565 18855
rect 32600 18820 32610 18855
rect 32645 18820 32655 18855
rect 32690 18820 32700 18855
rect 32735 18820 32745 18855
rect 32780 18820 32790 18855
rect 32825 18820 32835 18855
rect 32870 18820 32890 18855
rect 31290 18810 32890 18820
rect 31290 18775 31305 18810
rect 31340 18775 31350 18810
rect 31385 18775 31395 18810
rect 31430 18775 31440 18810
rect 31475 18775 31485 18810
rect 31520 18775 31530 18810
rect 31565 18775 31575 18810
rect 31610 18775 31620 18810
rect 31655 18775 31665 18810
rect 31700 18775 31710 18810
rect 31745 18775 31755 18810
rect 31790 18775 31800 18810
rect 31835 18775 31845 18810
rect 31880 18775 31890 18810
rect 31925 18775 31935 18810
rect 31970 18775 31980 18810
rect 32015 18775 32025 18810
rect 32060 18775 32070 18810
rect 32105 18775 32115 18810
rect 32150 18775 32160 18810
rect 32195 18775 32205 18810
rect 32240 18775 32250 18810
rect 32285 18775 32295 18810
rect 32330 18775 32340 18810
rect 32375 18775 32385 18810
rect 32420 18775 32430 18810
rect 32465 18775 32475 18810
rect 32510 18775 32520 18810
rect 32555 18775 32565 18810
rect 32600 18775 32610 18810
rect 32645 18775 32655 18810
rect 32690 18775 32700 18810
rect 32735 18775 32745 18810
rect 32780 18775 32790 18810
rect 32825 18775 32835 18810
rect 32870 18775 32890 18810
rect 31290 18765 32890 18775
rect 31290 18730 31305 18765
rect 31340 18730 31350 18765
rect 31385 18730 31395 18765
rect 31430 18730 31440 18765
rect 31475 18730 31485 18765
rect 31520 18730 31530 18765
rect 31565 18730 31575 18765
rect 31610 18730 31620 18765
rect 31655 18730 31665 18765
rect 31700 18730 31710 18765
rect 31745 18730 31755 18765
rect 31790 18730 31800 18765
rect 31835 18730 31845 18765
rect 31880 18730 31890 18765
rect 31925 18730 31935 18765
rect 31970 18730 31980 18765
rect 32015 18730 32025 18765
rect 32060 18730 32070 18765
rect 32105 18730 32115 18765
rect 32150 18730 32160 18765
rect 32195 18730 32205 18765
rect 32240 18730 32250 18765
rect 32285 18730 32295 18765
rect 32330 18730 32340 18765
rect 32375 18730 32385 18765
rect 32420 18730 32430 18765
rect 32465 18730 32475 18765
rect 32510 18730 32520 18765
rect 32555 18730 32565 18765
rect 32600 18730 32610 18765
rect 32645 18730 32655 18765
rect 32690 18730 32700 18765
rect 32735 18730 32745 18765
rect 32780 18730 32790 18765
rect 32825 18730 32835 18765
rect 32870 18730 32890 18765
rect 31290 18720 32890 18730
rect 31290 18685 31305 18720
rect 31340 18685 31350 18720
rect 31385 18685 31395 18720
rect 31430 18685 31440 18720
rect 31475 18685 31485 18720
rect 31520 18685 31530 18720
rect 31565 18685 31575 18720
rect 31610 18685 31620 18720
rect 31655 18685 31665 18720
rect 31700 18685 31710 18720
rect 31745 18685 31755 18720
rect 31790 18685 31800 18720
rect 31835 18685 31845 18720
rect 31880 18685 31890 18720
rect 31925 18685 31935 18720
rect 31970 18685 31980 18720
rect 32015 18685 32025 18720
rect 32060 18685 32070 18720
rect 32105 18685 32115 18720
rect 32150 18685 32160 18720
rect 32195 18685 32205 18720
rect 32240 18685 32250 18720
rect 32285 18685 32295 18720
rect 32330 18685 32340 18720
rect 32375 18685 32385 18720
rect 32420 18685 32430 18720
rect 32465 18685 32475 18720
rect 32510 18685 32520 18720
rect 32555 18685 32565 18720
rect 32600 18685 32610 18720
rect 32645 18685 32655 18720
rect 32690 18685 32700 18720
rect 32735 18685 32745 18720
rect 32780 18685 32790 18720
rect 32825 18685 32835 18720
rect 32870 18685 32890 18720
rect 31290 18675 32890 18685
rect 31290 18640 31305 18675
rect 31340 18640 31350 18675
rect 31385 18640 31395 18675
rect 31430 18640 31440 18675
rect 31475 18640 31485 18675
rect 31520 18640 31530 18675
rect 31565 18640 31575 18675
rect 31610 18640 31620 18675
rect 31655 18640 31665 18675
rect 31700 18640 31710 18675
rect 31745 18640 31755 18675
rect 31790 18640 31800 18675
rect 31835 18640 31845 18675
rect 31880 18640 31890 18675
rect 31925 18640 31935 18675
rect 31970 18640 31980 18675
rect 32015 18640 32025 18675
rect 32060 18640 32070 18675
rect 32105 18640 32115 18675
rect 32150 18640 32160 18675
rect 32195 18640 32205 18675
rect 32240 18640 32250 18675
rect 32285 18640 32295 18675
rect 32330 18640 32340 18675
rect 32375 18640 32385 18675
rect 32420 18640 32430 18675
rect 32465 18640 32475 18675
rect 32510 18640 32520 18675
rect 32555 18640 32565 18675
rect 32600 18640 32610 18675
rect 32645 18640 32655 18675
rect 32690 18640 32700 18675
rect 32735 18640 32745 18675
rect 32780 18640 32790 18675
rect 32825 18640 32835 18675
rect 32870 18640 32890 18675
rect 31290 18630 32890 18640
rect 31290 18595 31305 18630
rect 31340 18595 31350 18630
rect 31385 18595 31395 18630
rect 31430 18595 31440 18630
rect 31475 18595 31485 18630
rect 31520 18595 31530 18630
rect 31565 18595 31575 18630
rect 31610 18595 31620 18630
rect 31655 18595 31665 18630
rect 31700 18595 31710 18630
rect 31745 18595 31755 18630
rect 31790 18595 31800 18630
rect 31835 18595 31845 18630
rect 31880 18595 31890 18630
rect 31925 18595 31935 18630
rect 31970 18595 31980 18630
rect 32015 18595 32025 18630
rect 32060 18595 32070 18630
rect 32105 18595 32115 18630
rect 32150 18595 32160 18630
rect 32195 18595 32205 18630
rect 32240 18595 32250 18630
rect 32285 18595 32295 18630
rect 32330 18595 32340 18630
rect 32375 18595 32385 18630
rect 32420 18595 32430 18630
rect 32465 18595 32475 18630
rect 32510 18595 32520 18630
rect 32555 18595 32565 18630
rect 32600 18595 32610 18630
rect 32645 18595 32655 18630
rect 32690 18595 32700 18630
rect 32735 18595 32745 18630
rect 32780 18595 32790 18630
rect 32825 18595 32835 18630
rect 32870 18595 32890 18630
rect 31290 18585 32890 18595
rect 31290 18550 31305 18585
rect 31340 18550 31350 18585
rect 31385 18550 31395 18585
rect 31430 18550 31440 18585
rect 31475 18550 31485 18585
rect 31520 18550 31530 18585
rect 31565 18550 31575 18585
rect 31610 18550 31620 18585
rect 31655 18550 31665 18585
rect 31700 18550 31710 18585
rect 31745 18550 31755 18585
rect 31790 18550 31800 18585
rect 31835 18550 31845 18585
rect 31880 18550 31890 18585
rect 31925 18550 31935 18585
rect 31970 18550 31980 18585
rect 32015 18550 32025 18585
rect 32060 18550 32070 18585
rect 32105 18550 32115 18585
rect 32150 18550 32160 18585
rect 32195 18550 32205 18585
rect 32240 18550 32250 18585
rect 32285 18550 32295 18585
rect 32330 18550 32340 18585
rect 32375 18550 32385 18585
rect 32420 18550 32430 18585
rect 32465 18550 32475 18585
rect 32510 18550 32520 18585
rect 32555 18550 32565 18585
rect 32600 18550 32610 18585
rect 32645 18550 32655 18585
rect 32690 18550 32700 18585
rect 32735 18550 32745 18585
rect 32780 18550 32790 18585
rect 32825 18550 32835 18585
rect 32870 18550 32890 18585
rect 31290 18540 32890 18550
rect 31290 18505 31305 18540
rect 31340 18505 31350 18540
rect 31385 18505 31395 18540
rect 31430 18505 31440 18540
rect 31475 18505 31485 18540
rect 31520 18505 31530 18540
rect 31565 18505 31575 18540
rect 31610 18505 31620 18540
rect 31655 18505 31665 18540
rect 31700 18505 31710 18540
rect 31745 18505 31755 18540
rect 31790 18505 31800 18540
rect 31835 18505 31845 18540
rect 31880 18505 31890 18540
rect 31925 18505 31935 18540
rect 31970 18505 31980 18540
rect 32015 18505 32025 18540
rect 32060 18505 32070 18540
rect 32105 18505 32115 18540
rect 32150 18505 32160 18540
rect 32195 18505 32205 18540
rect 32240 18505 32250 18540
rect 32285 18505 32295 18540
rect 32330 18505 32340 18540
rect 32375 18505 32385 18540
rect 32420 18505 32430 18540
rect 32465 18505 32475 18540
rect 32510 18505 32520 18540
rect 32555 18505 32565 18540
rect 32600 18505 32610 18540
rect 32645 18505 32655 18540
rect 32690 18505 32700 18540
rect 32735 18505 32745 18540
rect 32780 18505 32790 18540
rect 32825 18505 32835 18540
rect 32870 18505 32890 18540
rect 31290 18495 32890 18505
rect 31290 18460 31305 18495
rect 31340 18460 31350 18495
rect 31385 18460 31395 18495
rect 31430 18460 31440 18495
rect 31475 18460 31485 18495
rect 31520 18460 31530 18495
rect 31565 18460 31575 18495
rect 31610 18460 31620 18495
rect 31655 18460 31665 18495
rect 31700 18460 31710 18495
rect 31745 18460 31755 18495
rect 31790 18460 31800 18495
rect 31835 18460 31845 18495
rect 31880 18460 31890 18495
rect 31925 18460 31935 18495
rect 31970 18460 31980 18495
rect 32015 18460 32025 18495
rect 32060 18460 32070 18495
rect 32105 18460 32115 18495
rect 32150 18460 32160 18495
rect 32195 18460 32205 18495
rect 32240 18460 32250 18495
rect 32285 18460 32295 18495
rect 32330 18460 32340 18495
rect 32375 18460 32385 18495
rect 32420 18460 32430 18495
rect 32465 18460 32475 18495
rect 32510 18460 32520 18495
rect 32555 18460 32565 18495
rect 32600 18460 32610 18495
rect 32645 18460 32655 18495
rect 32690 18460 32700 18495
rect 32735 18460 32745 18495
rect 32780 18460 32790 18495
rect 32825 18460 32835 18495
rect 32870 18460 32890 18495
rect 31290 18450 32890 18460
rect 31290 18415 31305 18450
rect 31340 18415 31350 18450
rect 31385 18415 31395 18450
rect 31430 18415 31440 18450
rect 31475 18415 31485 18450
rect 31520 18415 31530 18450
rect 31565 18415 31575 18450
rect 31610 18415 31620 18450
rect 31655 18415 31665 18450
rect 31700 18415 31710 18450
rect 31745 18415 31755 18450
rect 31790 18415 31800 18450
rect 31835 18415 31845 18450
rect 31880 18415 31890 18450
rect 31925 18415 31935 18450
rect 31970 18415 31980 18450
rect 32015 18415 32025 18450
rect 32060 18415 32070 18450
rect 32105 18415 32115 18450
rect 32150 18415 32160 18450
rect 32195 18415 32205 18450
rect 32240 18415 32250 18450
rect 32285 18415 32295 18450
rect 32330 18415 32340 18450
rect 32375 18415 32385 18450
rect 32420 18415 32430 18450
rect 32465 18415 32475 18450
rect 32510 18415 32520 18450
rect 32555 18415 32565 18450
rect 32600 18415 32610 18450
rect 32645 18415 32655 18450
rect 32690 18415 32700 18450
rect 32735 18415 32745 18450
rect 32780 18415 32790 18450
rect 32825 18415 32835 18450
rect 32870 18415 32890 18450
rect 31290 18405 32890 18415
rect 31290 18370 31305 18405
rect 31340 18370 31350 18405
rect 31385 18370 31395 18405
rect 31430 18370 31440 18405
rect 31475 18370 31485 18405
rect 31520 18370 31530 18405
rect 31565 18370 31575 18405
rect 31610 18370 31620 18405
rect 31655 18370 31665 18405
rect 31700 18370 31710 18405
rect 31745 18370 31755 18405
rect 31790 18370 31800 18405
rect 31835 18370 31845 18405
rect 31880 18370 31890 18405
rect 31925 18370 31935 18405
rect 31970 18370 31980 18405
rect 32015 18370 32025 18405
rect 32060 18370 32070 18405
rect 32105 18370 32115 18405
rect 32150 18370 32160 18405
rect 32195 18370 32205 18405
rect 32240 18370 32250 18405
rect 32285 18370 32295 18405
rect 32330 18370 32340 18405
rect 32375 18370 32385 18405
rect 32420 18370 32430 18405
rect 32465 18370 32475 18405
rect 32510 18370 32520 18405
rect 32555 18370 32565 18405
rect 32600 18370 32610 18405
rect 32645 18370 32655 18405
rect 32690 18370 32700 18405
rect 32735 18370 32745 18405
rect 32780 18370 32790 18405
rect 32825 18370 32835 18405
rect 32870 18370 32890 18405
rect 31290 18360 32890 18370
rect 31290 18325 31305 18360
rect 31340 18325 31350 18360
rect 31385 18325 31395 18360
rect 31430 18325 31440 18360
rect 31475 18325 31485 18360
rect 31520 18325 31530 18360
rect 31565 18325 31575 18360
rect 31610 18325 31620 18360
rect 31655 18325 31665 18360
rect 31700 18325 31710 18360
rect 31745 18325 31755 18360
rect 31790 18325 31800 18360
rect 31835 18325 31845 18360
rect 31880 18325 31890 18360
rect 31925 18325 31935 18360
rect 31970 18325 31980 18360
rect 32015 18325 32025 18360
rect 32060 18325 32070 18360
rect 32105 18325 32115 18360
rect 32150 18325 32160 18360
rect 32195 18325 32205 18360
rect 32240 18325 32250 18360
rect 32285 18325 32295 18360
rect 32330 18325 32340 18360
rect 32375 18325 32385 18360
rect 32420 18325 32430 18360
rect 32465 18325 32475 18360
rect 32510 18325 32520 18360
rect 32555 18325 32565 18360
rect 32600 18325 32610 18360
rect 32645 18325 32655 18360
rect 32690 18325 32700 18360
rect 32735 18325 32745 18360
rect 32780 18325 32790 18360
rect 32825 18325 32835 18360
rect 32870 18325 32890 18360
rect 31290 18315 32890 18325
rect 31290 18280 31305 18315
rect 31340 18280 31350 18315
rect 31385 18280 31395 18315
rect 31430 18280 31440 18315
rect 31475 18280 31485 18315
rect 31520 18280 31530 18315
rect 31565 18280 31575 18315
rect 31610 18280 31620 18315
rect 31655 18280 31665 18315
rect 31700 18280 31710 18315
rect 31745 18280 31755 18315
rect 31790 18280 31800 18315
rect 31835 18280 31845 18315
rect 31880 18280 31890 18315
rect 31925 18280 31935 18315
rect 31970 18280 31980 18315
rect 32015 18280 32025 18315
rect 32060 18280 32070 18315
rect 32105 18280 32115 18315
rect 32150 18280 32160 18315
rect 32195 18280 32205 18315
rect 32240 18280 32250 18315
rect 32285 18280 32295 18315
rect 32330 18280 32340 18315
rect 32375 18280 32385 18315
rect 32420 18280 32430 18315
rect 32465 18280 32475 18315
rect 32510 18280 32520 18315
rect 32555 18280 32565 18315
rect 32600 18280 32610 18315
rect 32645 18280 32655 18315
rect 32690 18280 32700 18315
rect 32735 18280 32745 18315
rect 32780 18280 32790 18315
rect 32825 18280 32835 18315
rect 32870 18280 32890 18315
rect 31290 18270 32890 18280
rect 31290 18235 31305 18270
rect 31340 18235 31350 18270
rect 31385 18235 31395 18270
rect 31430 18235 31440 18270
rect 31475 18235 31485 18270
rect 31520 18235 31530 18270
rect 31565 18235 31575 18270
rect 31610 18235 31620 18270
rect 31655 18235 31665 18270
rect 31700 18235 31710 18270
rect 31745 18235 31755 18270
rect 31790 18235 31800 18270
rect 31835 18235 31845 18270
rect 31880 18235 31890 18270
rect 31925 18235 31935 18270
rect 31970 18235 31980 18270
rect 32015 18235 32025 18270
rect 32060 18235 32070 18270
rect 32105 18235 32115 18270
rect 32150 18235 32160 18270
rect 32195 18235 32205 18270
rect 32240 18235 32250 18270
rect 32285 18235 32295 18270
rect 32330 18235 32340 18270
rect 32375 18235 32385 18270
rect 32420 18235 32430 18270
rect 32465 18235 32475 18270
rect 32510 18235 32520 18270
rect 32555 18235 32565 18270
rect 32600 18235 32610 18270
rect 32645 18235 32655 18270
rect 32690 18235 32700 18270
rect 32735 18235 32745 18270
rect 32780 18235 32790 18270
rect 32825 18235 32835 18270
rect 32870 18235 32890 18270
rect 31290 18225 32890 18235
rect 31290 18190 31305 18225
rect 31340 18190 31350 18225
rect 31385 18190 31395 18225
rect 31430 18190 31440 18225
rect 31475 18190 31485 18225
rect 31520 18190 31530 18225
rect 31565 18190 31575 18225
rect 31610 18190 31620 18225
rect 31655 18190 31665 18225
rect 31700 18190 31710 18225
rect 31745 18190 31755 18225
rect 31790 18190 31800 18225
rect 31835 18190 31845 18225
rect 31880 18190 31890 18225
rect 31925 18190 31935 18225
rect 31970 18190 31980 18225
rect 32015 18190 32025 18225
rect 32060 18190 32070 18225
rect 32105 18190 32115 18225
rect 32150 18190 32160 18225
rect 32195 18190 32205 18225
rect 32240 18190 32250 18225
rect 32285 18190 32295 18225
rect 32330 18190 32340 18225
rect 32375 18190 32385 18225
rect 32420 18190 32430 18225
rect 32465 18190 32475 18225
rect 32510 18190 32520 18225
rect 32555 18190 32565 18225
rect 32600 18190 32610 18225
rect 32645 18190 32655 18225
rect 32690 18190 32700 18225
rect 32735 18190 32745 18225
rect 32780 18190 32790 18225
rect 32825 18190 32835 18225
rect 32870 18190 32890 18225
rect 31290 18180 32890 18190
rect 31290 18145 31305 18180
rect 31340 18145 31350 18180
rect 31385 18145 31395 18180
rect 31430 18145 31440 18180
rect 31475 18145 31485 18180
rect 31520 18145 31530 18180
rect 31565 18145 31575 18180
rect 31610 18145 31620 18180
rect 31655 18145 31665 18180
rect 31700 18145 31710 18180
rect 31745 18145 31755 18180
rect 31790 18145 31800 18180
rect 31835 18145 31845 18180
rect 31880 18145 31890 18180
rect 31925 18145 31935 18180
rect 31970 18145 31980 18180
rect 32015 18145 32025 18180
rect 32060 18145 32070 18180
rect 32105 18145 32115 18180
rect 32150 18145 32160 18180
rect 32195 18145 32205 18180
rect 32240 18145 32250 18180
rect 32285 18145 32295 18180
rect 32330 18145 32340 18180
rect 32375 18145 32385 18180
rect 32420 18145 32430 18180
rect 32465 18145 32475 18180
rect 32510 18145 32520 18180
rect 32555 18145 32565 18180
rect 32600 18145 32610 18180
rect 32645 18145 32655 18180
rect 32690 18145 32700 18180
rect 32735 18145 32745 18180
rect 32780 18145 32790 18180
rect 32825 18145 32835 18180
rect 32870 18145 32890 18180
rect 31290 18135 32890 18145
rect 31290 18100 31305 18135
rect 31340 18100 31350 18135
rect 31385 18100 31395 18135
rect 31430 18100 31440 18135
rect 31475 18100 31485 18135
rect 31520 18100 31530 18135
rect 31565 18100 31575 18135
rect 31610 18100 31620 18135
rect 31655 18100 31665 18135
rect 31700 18100 31710 18135
rect 31745 18100 31755 18135
rect 31790 18100 31800 18135
rect 31835 18100 31845 18135
rect 31880 18100 31890 18135
rect 31925 18100 31935 18135
rect 31970 18100 31980 18135
rect 32015 18100 32025 18135
rect 32060 18100 32070 18135
rect 32105 18100 32115 18135
rect 32150 18100 32160 18135
rect 32195 18100 32205 18135
rect 32240 18100 32250 18135
rect 32285 18100 32295 18135
rect 32330 18100 32340 18135
rect 32375 18100 32385 18135
rect 32420 18100 32430 18135
rect 32465 18100 32475 18135
rect 32510 18100 32520 18135
rect 32555 18100 32565 18135
rect 32600 18100 32610 18135
rect 32645 18100 32655 18135
rect 32690 18100 32700 18135
rect 32735 18100 32745 18135
rect 32780 18100 32790 18135
rect 32825 18100 32835 18135
rect 32870 18100 32890 18135
rect 31290 18090 32890 18100
rect 31290 18055 31305 18090
rect 31340 18055 31350 18090
rect 31385 18055 31395 18090
rect 31430 18055 31440 18090
rect 31475 18055 31485 18090
rect 31520 18055 31530 18090
rect 31565 18055 31575 18090
rect 31610 18055 31620 18090
rect 31655 18055 31665 18090
rect 31700 18055 31710 18090
rect 31745 18055 31755 18090
rect 31790 18055 31800 18090
rect 31835 18055 31845 18090
rect 31880 18055 31890 18090
rect 31925 18055 31935 18090
rect 31970 18055 31980 18090
rect 32015 18055 32025 18090
rect 32060 18055 32070 18090
rect 32105 18055 32115 18090
rect 32150 18055 32160 18090
rect 32195 18055 32205 18090
rect 32240 18055 32250 18090
rect 32285 18055 32295 18090
rect 32330 18055 32340 18090
rect 32375 18055 32385 18090
rect 32420 18055 32430 18090
rect 32465 18055 32475 18090
rect 32510 18055 32520 18090
rect 32555 18055 32565 18090
rect 32600 18055 32610 18090
rect 32645 18055 32655 18090
rect 32690 18055 32700 18090
rect 32735 18055 32745 18090
rect 32780 18055 32790 18090
rect 32825 18055 32835 18090
rect 32870 18055 32890 18090
rect 31290 18045 32890 18055
rect 31290 18010 31305 18045
rect 31340 18010 31350 18045
rect 31385 18010 31395 18045
rect 31430 18010 31440 18045
rect 31475 18010 31485 18045
rect 31520 18010 31530 18045
rect 31565 18010 31575 18045
rect 31610 18010 31620 18045
rect 31655 18010 31665 18045
rect 31700 18010 31710 18045
rect 31745 18010 31755 18045
rect 31790 18010 31800 18045
rect 31835 18010 31845 18045
rect 31880 18010 31890 18045
rect 31925 18010 31935 18045
rect 31970 18010 31980 18045
rect 32015 18010 32025 18045
rect 32060 18010 32070 18045
rect 32105 18010 32115 18045
rect 32150 18010 32160 18045
rect 32195 18010 32205 18045
rect 32240 18010 32250 18045
rect 32285 18010 32295 18045
rect 32330 18010 32340 18045
rect 32375 18010 32385 18045
rect 32420 18010 32430 18045
rect 32465 18010 32475 18045
rect 32510 18010 32520 18045
rect 32555 18010 32565 18045
rect 32600 18010 32610 18045
rect 32645 18010 32655 18045
rect 32690 18010 32700 18045
rect 32735 18010 32745 18045
rect 32780 18010 32790 18045
rect 32825 18010 32835 18045
rect 32870 18010 32890 18045
rect 31290 18000 32890 18010
rect 31290 17965 31305 18000
rect 31340 17965 31350 18000
rect 31385 17965 31395 18000
rect 31430 17965 31440 18000
rect 31475 17965 31485 18000
rect 31520 17965 31530 18000
rect 31565 17965 31575 18000
rect 31610 17965 31620 18000
rect 31655 17965 31665 18000
rect 31700 17965 31710 18000
rect 31745 17965 31755 18000
rect 31790 17965 31800 18000
rect 31835 17965 31845 18000
rect 31880 17965 31890 18000
rect 31925 17965 31935 18000
rect 31970 17965 31980 18000
rect 32015 17965 32025 18000
rect 32060 17965 32070 18000
rect 32105 17965 32115 18000
rect 32150 17965 32160 18000
rect 32195 17965 32205 18000
rect 32240 17965 32250 18000
rect 32285 17965 32295 18000
rect 32330 17965 32340 18000
rect 32375 17965 32385 18000
rect 32420 17965 32430 18000
rect 32465 17965 32475 18000
rect 32510 17965 32520 18000
rect 32555 17965 32565 18000
rect 32600 17965 32610 18000
rect 32645 17965 32655 18000
rect 32690 17965 32700 18000
rect 32735 17965 32745 18000
rect 32780 17965 32790 18000
rect 32825 17965 32835 18000
rect 32870 17965 32890 18000
rect 31290 17955 32890 17965
rect 31290 17920 31305 17955
rect 31340 17920 31350 17955
rect 31385 17920 31395 17955
rect 31430 17920 31440 17955
rect 31475 17920 31485 17955
rect 31520 17920 31530 17955
rect 31565 17920 31575 17955
rect 31610 17920 31620 17955
rect 31655 17920 31665 17955
rect 31700 17920 31710 17955
rect 31745 17920 31755 17955
rect 31790 17920 31800 17955
rect 31835 17920 31845 17955
rect 31880 17920 31890 17955
rect 31925 17920 31935 17955
rect 31970 17920 31980 17955
rect 32015 17920 32025 17955
rect 32060 17920 32070 17955
rect 32105 17920 32115 17955
rect 32150 17920 32160 17955
rect 32195 17920 32205 17955
rect 32240 17920 32250 17955
rect 32285 17920 32295 17955
rect 32330 17920 32340 17955
rect 32375 17920 32385 17955
rect 32420 17920 32430 17955
rect 32465 17920 32475 17955
rect 32510 17920 32520 17955
rect 32555 17920 32565 17955
rect 32600 17920 32610 17955
rect 32645 17920 32655 17955
rect 32690 17920 32700 17955
rect 32735 17920 32745 17955
rect 32780 17920 32790 17955
rect 32825 17920 32835 17955
rect 32870 17920 32890 17955
rect 31290 17910 32890 17920
rect 31290 17875 31305 17910
rect 31340 17875 31350 17910
rect 31385 17875 31395 17910
rect 31430 17875 31440 17910
rect 31475 17875 31485 17910
rect 31520 17875 31530 17910
rect 31565 17875 31575 17910
rect 31610 17875 31620 17910
rect 31655 17875 31665 17910
rect 31700 17875 31710 17910
rect 31745 17875 31755 17910
rect 31790 17875 31800 17910
rect 31835 17875 31845 17910
rect 31880 17875 31890 17910
rect 31925 17875 31935 17910
rect 31970 17875 31980 17910
rect 32015 17875 32025 17910
rect 32060 17875 32070 17910
rect 32105 17875 32115 17910
rect 32150 17875 32160 17910
rect 32195 17875 32205 17910
rect 32240 17875 32250 17910
rect 32285 17875 32295 17910
rect 32330 17875 32340 17910
rect 32375 17875 32385 17910
rect 32420 17875 32430 17910
rect 32465 17875 32475 17910
rect 32510 17875 32520 17910
rect 32555 17875 32565 17910
rect 32600 17875 32610 17910
rect 32645 17875 32655 17910
rect 32690 17875 32700 17910
rect 32735 17875 32745 17910
rect 32780 17875 32790 17910
rect 32825 17875 32835 17910
rect 32870 17875 32890 17910
rect 31290 17865 32890 17875
rect 31290 17830 31305 17865
rect 31340 17830 31350 17865
rect 31385 17830 31395 17865
rect 31430 17830 31440 17865
rect 31475 17830 31485 17865
rect 31520 17830 31530 17865
rect 31565 17830 31575 17865
rect 31610 17830 31620 17865
rect 31655 17830 31665 17865
rect 31700 17830 31710 17865
rect 31745 17830 31755 17865
rect 31790 17830 31800 17865
rect 31835 17830 31845 17865
rect 31880 17830 31890 17865
rect 31925 17830 31935 17865
rect 31970 17830 31980 17865
rect 32015 17830 32025 17865
rect 32060 17830 32070 17865
rect 32105 17830 32115 17865
rect 32150 17830 32160 17865
rect 32195 17830 32205 17865
rect 32240 17830 32250 17865
rect 32285 17830 32295 17865
rect 32330 17830 32340 17865
rect 32375 17830 32385 17865
rect 32420 17830 32430 17865
rect 32465 17830 32475 17865
rect 32510 17830 32520 17865
rect 32555 17830 32565 17865
rect 32600 17830 32610 17865
rect 32645 17830 32655 17865
rect 32690 17830 32700 17865
rect 32735 17830 32745 17865
rect 32780 17830 32790 17865
rect 32825 17830 32835 17865
rect 32870 17830 32890 17865
rect 31290 17820 32890 17830
rect 31290 17785 31305 17820
rect 31340 17785 31350 17820
rect 31385 17785 31395 17820
rect 31430 17785 31440 17820
rect 31475 17785 31485 17820
rect 31520 17785 31530 17820
rect 31565 17785 31575 17820
rect 31610 17785 31620 17820
rect 31655 17785 31665 17820
rect 31700 17785 31710 17820
rect 31745 17785 31755 17820
rect 31790 17785 31800 17820
rect 31835 17785 31845 17820
rect 31880 17785 31890 17820
rect 31925 17785 31935 17820
rect 31970 17785 31980 17820
rect 32015 17785 32025 17820
rect 32060 17785 32070 17820
rect 32105 17785 32115 17820
rect 32150 17785 32160 17820
rect 32195 17785 32205 17820
rect 32240 17785 32250 17820
rect 32285 17785 32295 17820
rect 32330 17785 32340 17820
rect 32375 17785 32385 17820
rect 32420 17785 32430 17820
rect 32465 17785 32475 17820
rect 32510 17785 32520 17820
rect 32555 17785 32565 17820
rect 32600 17785 32610 17820
rect 32645 17785 32655 17820
rect 32690 17785 32700 17820
rect 32735 17785 32745 17820
rect 32780 17785 32790 17820
rect 32825 17785 32835 17820
rect 32870 17785 32890 17820
rect 31290 17775 32890 17785
rect 31290 17740 31305 17775
rect 31340 17740 31350 17775
rect 31385 17740 31395 17775
rect 31430 17740 31440 17775
rect 31475 17740 31485 17775
rect 31520 17740 31530 17775
rect 31565 17740 31575 17775
rect 31610 17740 31620 17775
rect 31655 17740 31665 17775
rect 31700 17740 31710 17775
rect 31745 17740 31755 17775
rect 31790 17740 31800 17775
rect 31835 17740 31845 17775
rect 31880 17740 31890 17775
rect 31925 17740 31935 17775
rect 31970 17740 31980 17775
rect 32015 17740 32025 17775
rect 32060 17740 32070 17775
rect 32105 17740 32115 17775
rect 32150 17740 32160 17775
rect 32195 17740 32205 17775
rect 32240 17740 32250 17775
rect 32285 17740 32295 17775
rect 32330 17740 32340 17775
rect 32375 17740 32385 17775
rect 32420 17740 32430 17775
rect 32465 17740 32475 17775
rect 32510 17740 32520 17775
rect 32555 17740 32565 17775
rect 32600 17740 32610 17775
rect 32645 17740 32655 17775
rect 32690 17740 32700 17775
rect 32735 17740 32745 17775
rect 32780 17740 32790 17775
rect 32825 17740 32835 17775
rect 32870 17740 32890 17775
rect -38770 9630 -37170 10155
rect -38770 9595 -38755 9630
rect -38720 9595 -38710 9630
rect -38675 9595 -38665 9630
rect -38630 9595 -38620 9630
rect -38585 9595 -38575 9630
rect -38540 9595 -38530 9630
rect -38495 9595 -38485 9630
rect -38450 9595 -38440 9630
rect -38405 9595 -38395 9630
rect -38360 9595 -38350 9630
rect -38315 9595 -38305 9630
rect -38270 9595 -38260 9630
rect -38225 9595 -38215 9630
rect -38180 9595 -38170 9630
rect -38135 9595 -38125 9630
rect -38090 9595 -38080 9630
rect -38045 9595 -38035 9630
rect -38000 9595 -37990 9630
rect -37955 9595 -37945 9630
rect -37910 9595 -37900 9630
rect -37865 9595 -37855 9630
rect -37820 9595 -37810 9630
rect -37775 9595 -37765 9630
rect -37730 9595 -37720 9630
rect -37685 9595 -37675 9630
rect -37640 9595 -37630 9630
rect -37595 9595 -37585 9630
rect -37550 9595 -37540 9630
rect -37505 9595 -37495 9630
rect -37460 9595 -37450 9630
rect -37415 9595 -37405 9630
rect -37370 9595 -37360 9630
rect -37325 9595 -37315 9630
rect -37280 9595 -37270 9630
rect -37235 9595 -37225 9630
rect -37190 9595 -37170 9630
rect -38770 9585 -37170 9595
rect -38770 9550 -38755 9585
rect -38720 9550 -38710 9585
rect -38675 9550 -38665 9585
rect -38630 9550 -38620 9585
rect -38585 9550 -38575 9585
rect -38540 9550 -38530 9585
rect -38495 9550 -38485 9585
rect -38450 9550 -38440 9585
rect -38405 9550 -38395 9585
rect -38360 9550 -38350 9585
rect -38315 9550 -38305 9585
rect -38270 9550 -38260 9585
rect -38225 9550 -38215 9585
rect -38180 9550 -38170 9585
rect -38135 9550 -38125 9585
rect -38090 9550 -38080 9585
rect -38045 9550 -38035 9585
rect -38000 9550 -37990 9585
rect -37955 9550 -37945 9585
rect -37910 9550 -37900 9585
rect -37865 9550 -37855 9585
rect -37820 9550 -37810 9585
rect -37775 9550 -37765 9585
rect -37730 9550 -37720 9585
rect -37685 9550 -37675 9585
rect -37640 9550 -37630 9585
rect -37595 9550 -37585 9585
rect -37550 9550 -37540 9585
rect -37505 9550 -37495 9585
rect -37460 9550 -37450 9585
rect -37415 9550 -37405 9585
rect -37370 9550 -37360 9585
rect -37325 9550 -37315 9585
rect -37280 9550 -37270 9585
rect -37235 9550 -37225 9585
rect -37190 9550 -37170 9585
rect -38770 9540 -37170 9550
rect -38770 9505 -38755 9540
rect -38720 9505 -38710 9540
rect -38675 9505 -38665 9540
rect -38630 9505 -38620 9540
rect -38585 9505 -38575 9540
rect -38540 9505 -38530 9540
rect -38495 9505 -38485 9540
rect -38450 9505 -38440 9540
rect -38405 9505 -38395 9540
rect -38360 9505 -38350 9540
rect -38315 9505 -38305 9540
rect -38270 9505 -38260 9540
rect -38225 9505 -38215 9540
rect -38180 9505 -38170 9540
rect -38135 9505 -38125 9540
rect -38090 9505 -38080 9540
rect -38045 9505 -38035 9540
rect -38000 9505 -37990 9540
rect -37955 9505 -37945 9540
rect -37910 9505 -37900 9540
rect -37865 9505 -37855 9540
rect -37820 9505 -37810 9540
rect -37775 9505 -37765 9540
rect -37730 9505 -37720 9540
rect -37685 9505 -37675 9540
rect -37640 9505 -37630 9540
rect -37595 9505 -37585 9540
rect -37550 9505 -37540 9540
rect -37505 9505 -37495 9540
rect -37460 9505 -37450 9540
rect -37415 9505 -37405 9540
rect -37370 9505 -37360 9540
rect -37325 9505 -37315 9540
rect -37280 9505 -37270 9540
rect -37235 9505 -37225 9540
rect -37190 9505 -37170 9540
rect -38770 9495 -37170 9505
rect -38770 9460 -38755 9495
rect -38720 9460 -38710 9495
rect -38675 9460 -38665 9495
rect -38630 9460 -38620 9495
rect -38585 9460 -38575 9495
rect -38540 9460 -38530 9495
rect -38495 9460 -38485 9495
rect -38450 9460 -38440 9495
rect -38405 9460 -38395 9495
rect -38360 9460 -38350 9495
rect -38315 9460 -38305 9495
rect -38270 9460 -38260 9495
rect -38225 9460 -38215 9495
rect -38180 9460 -38170 9495
rect -38135 9460 -38125 9495
rect -38090 9460 -38080 9495
rect -38045 9460 -38035 9495
rect -38000 9460 -37990 9495
rect -37955 9460 -37945 9495
rect -37910 9460 -37900 9495
rect -37865 9460 -37855 9495
rect -37820 9460 -37810 9495
rect -37775 9460 -37765 9495
rect -37730 9460 -37720 9495
rect -37685 9460 -37675 9495
rect -37640 9460 -37630 9495
rect -37595 9460 -37585 9495
rect -37550 9460 -37540 9495
rect -37505 9460 -37495 9495
rect -37460 9460 -37450 9495
rect -37415 9460 -37405 9495
rect -37370 9460 -37360 9495
rect -37325 9460 -37315 9495
rect -37280 9460 -37270 9495
rect -37235 9460 -37225 9495
rect -37190 9460 -37170 9495
rect -38770 9450 -37170 9460
rect -38770 9415 -38755 9450
rect -38720 9415 -38710 9450
rect -38675 9415 -38665 9450
rect -38630 9415 -38620 9450
rect -38585 9415 -38575 9450
rect -38540 9415 -38530 9450
rect -38495 9415 -38485 9450
rect -38450 9415 -38440 9450
rect -38405 9415 -38395 9450
rect -38360 9415 -38350 9450
rect -38315 9415 -38305 9450
rect -38270 9415 -38260 9450
rect -38225 9415 -38215 9450
rect -38180 9415 -38170 9450
rect -38135 9415 -38125 9450
rect -38090 9415 -38080 9450
rect -38045 9415 -38035 9450
rect -38000 9415 -37990 9450
rect -37955 9415 -37945 9450
rect -37910 9415 -37900 9450
rect -37865 9415 -37855 9450
rect -37820 9415 -37810 9450
rect -37775 9415 -37765 9450
rect -37730 9415 -37720 9450
rect -37685 9415 -37675 9450
rect -37640 9415 -37630 9450
rect -37595 9415 -37585 9450
rect -37550 9415 -37540 9450
rect -37505 9415 -37495 9450
rect -37460 9415 -37450 9450
rect -37415 9415 -37405 9450
rect -37370 9415 -37360 9450
rect -37325 9415 -37315 9450
rect -37280 9415 -37270 9450
rect -37235 9415 -37225 9450
rect -37190 9415 -37170 9450
rect -38770 9405 -37170 9415
rect -38770 9370 -38755 9405
rect -38720 9370 -38710 9405
rect -38675 9370 -38665 9405
rect -38630 9370 -38620 9405
rect -38585 9370 -38575 9405
rect -38540 9370 -38530 9405
rect -38495 9370 -38485 9405
rect -38450 9370 -38440 9405
rect -38405 9370 -38395 9405
rect -38360 9370 -38350 9405
rect -38315 9370 -38305 9405
rect -38270 9370 -38260 9405
rect -38225 9370 -38215 9405
rect -38180 9370 -38170 9405
rect -38135 9370 -38125 9405
rect -38090 9370 -38080 9405
rect -38045 9370 -38035 9405
rect -38000 9370 -37990 9405
rect -37955 9370 -37945 9405
rect -37910 9370 -37900 9405
rect -37865 9370 -37855 9405
rect -37820 9370 -37810 9405
rect -37775 9370 -37765 9405
rect -37730 9370 -37720 9405
rect -37685 9370 -37675 9405
rect -37640 9370 -37630 9405
rect -37595 9370 -37585 9405
rect -37550 9370 -37540 9405
rect -37505 9370 -37495 9405
rect -37460 9370 -37450 9405
rect -37415 9370 -37405 9405
rect -37370 9370 -37360 9405
rect -37325 9370 -37315 9405
rect -37280 9370 -37270 9405
rect -37235 9370 -37225 9405
rect -37190 9370 -37170 9405
rect -38770 9360 -37170 9370
rect -38770 9325 -38755 9360
rect -38720 9325 -38710 9360
rect -38675 9325 -38665 9360
rect -38630 9325 -38620 9360
rect -38585 9325 -38575 9360
rect -38540 9325 -38530 9360
rect -38495 9325 -38485 9360
rect -38450 9325 -38440 9360
rect -38405 9325 -38395 9360
rect -38360 9325 -38350 9360
rect -38315 9325 -38305 9360
rect -38270 9325 -38260 9360
rect -38225 9325 -38215 9360
rect -38180 9325 -38170 9360
rect -38135 9325 -38125 9360
rect -38090 9325 -38080 9360
rect -38045 9325 -38035 9360
rect -38000 9325 -37990 9360
rect -37955 9325 -37945 9360
rect -37910 9325 -37900 9360
rect -37865 9325 -37855 9360
rect -37820 9325 -37810 9360
rect -37775 9325 -37765 9360
rect -37730 9325 -37720 9360
rect -37685 9325 -37675 9360
rect -37640 9325 -37630 9360
rect -37595 9325 -37585 9360
rect -37550 9325 -37540 9360
rect -37505 9325 -37495 9360
rect -37460 9325 -37450 9360
rect -37415 9325 -37405 9360
rect -37370 9325 -37360 9360
rect -37325 9325 -37315 9360
rect -37280 9325 -37270 9360
rect -37235 9325 -37225 9360
rect -37190 9325 -37170 9360
rect -38770 9315 -37170 9325
rect -38770 9280 -38755 9315
rect -38720 9280 -38710 9315
rect -38675 9280 -38665 9315
rect -38630 9280 -38620 9315
rect -38585 9280 -38575 9315
rect -38540 9280 -38530 9315
rect -38495 9280 -38485 9315
rect -38450 9280 -38440 9315
rect -38405 9280 -38395 9315
rect -38360 9280 -38350 9315
rect -38315 9280 -38305 9315
rect -38270 9280 -38260 9315
rect -38225 9280 -38215 9315
rect -38180 9280 -38170 9315
rect -38135 9280 -38125 9315
rect -38090 9280 -38080 9315
rect -38045 9280 -38035 9315
rect -38000 9280 -37990 9315
rect -37955 9280 -37945 9315
rect -37910 9280 -37900 9315
rect -37865 9280 -37855 9315
rect -37820 9280 -37810 9315
rect -37775 9280 -37765 9315
rect -37730 9280 -37720 9315
rect -37685 9280 -37675 9315
rect -37640 9280 -37630 9315
rect -37595 9280 -37585 9315
rect -37550 9280 -37540 9315
rect -37505 9280 -37495 9315
rect -37460 9280 -37450 9315
rect -37415 9280 -37405 9315
rect -37370 9280 -37360 9315
rect -37325 9280 -37315 9315
rect -37280 9280 -37270 9315
rect -37235 9280 -37225 9315
rect -37190 9280 -37170 9315
rect -38770 9270 -37170 9280
rect -38770 9235 -38755 9270
rect -38720 9235 -38710 9270
rect -38675 9235 -38665 9270
rect -38630 9235 -38620 9270
rect -38585 9235 -38575 9270
rect -38540 9235 -38530 9270
rect -38495 9235 -38485 9270
rect -38450 9235 -38440 9270
rect -38405 9235 -38395 9270
rect -38360 9235 -38350 9270
rect -38315 9235 -38305 9270
rect -38270 9235 -38260 9270
rect -38225 9235 -38215 9270
rect -38180 9235 -38170 9270
rect -38135 9235 -38125 9270
rect -38090 9235 -38080 9270
rect -38045 9235 -38035 9270
rect -38000 9235 -37990 9270
rect -37955 9235 -37945 9270
rect -37910 9235 -37900 9270
rect -37865 9235 -37855 9270
rect -37820 9235 -37810 9270
rect -37775 9235 -37765 9270
rect -37730 9235 -37720 9270
rect -37685 9235 -37675 9270
rect -37640 9235 -37630 9270
rect -37595 9235 -37585 9270
rect -37550 9235 -37540 9270
rect -37505 9235 -37495 9270
rect -37460 9235 -37450 9270
rect -37415 9235 -37405 9270
rect -37370 9235 -37360 9270
rect -37325 9235 -37315 9270
rect -37280 9235 -37270 9270
rect -37235 9235 -37225 9270
rect -37190 9235 -37170 9270
rect -38770 9225 -37170 9235
rect -38770 9190 -38755 9225
rect -38720 9190 -38710 9225
rect -38675 9190 -38665 9225
rect -38630 9190 -38620 9225
rect -38585 9190 -38575 9225
rect -38540 9190 -38530 9225
rect -38495 9190 -38485 9225
rect -38450 9190 -38440 9225
rect -38405 9190 -38395 9225
rect -38360 9190 -38350 9225
rect -38315 9190 -38305 9225
rect -38270 9190 -38260 9225
rect -38225 9190 -38215 9225
rect -38180 9190 -38170 9225
rect -38135 9190 -38125 9225
rect -38090 9190 -38080 9225
rect -38045 9190 -38035 9225
rect -38000 9190 -37990 9225
rect -37955 9190 -37945 9225
rect -37910 9190 -37900 9225
rect -37865 9190 -37855 9225
rect -37820 9190 -37810 9225
rect -37775 9190 -37765 9225
rect -37730 9190 -37720 9225
rect -37685 9190 -37675 9225
rect -37640 9190 -37630 9225
rect -37595 9190 -37585 9225
rect -37550 9190 -37540 9225
rect -37505 9190 -37495 9225
rect -37460 9190 -37450 9225
rect -37415 9190 -37405 9225
rect -37370 9190 -37360 9225
rect -37325 9190 -37315 9225
rect -37280 9190 -37270 9225
rect -37235 9190 -37225 9225
rect -37190 9190 -37170 9225
rect -38770 9180 -37170 9190
rect -38770 9145 -38755 9180
rect -38720 9145 -38710 9180
rect -38675 9145 -38665 9180
rect -38630 9145 -38620 9180
rect -38585 9145 -38575 9180
rect -38540 9145 -38530 9180
rect -38495 9145 -38485 9180
rect -38450 9145 -38440 9180
rect -38405 9145 -38395 9180
rect -38360 9145 -38350 9180
rect -38315 9145 -38305 9180
rect -38270 9145 -38260 9180
rect -38225 9145 -38215 9180
rect -38180 9145 -38170 9180
rect -38135 9145 -38125 9180
rect -38090 9145 -38080 9180
rect -38045 9145 -38035 9180
rect -38000 9145 -37990 9180
rect -37955 9145 -37945 9180
rect -37910 9145 -37900 9180
rect -37865 9145 -37855 9180
rect -37820 9145 -37810 9180
rect -37775 9145 -37765 9180
rect -37730 9145 -37720 9180
rect -37685 9145 -37675 9180
rect -37640 9145 -37630 9180
rect -37595 9145 -37585 9180
rect -37550 9145 -37540 9180
rect -37505 9145 -37495 9180
rect -37460 9145 -37450 9180
rect -37415 9145 -37405 9180
rect -37370 9145 -37360 9180
rect -37325 9145 -37315 9180
rect -37280 9145 -37270 9180
rect -37235 9145 -37225 9180
rect -37190 9145 -37170 9180
rect -38770 9135 -37170 9145
rect -38770 9100 -38755 9135
rect -38720 9100 -38710 9135
rect -38675 9100 -38665 9135
rect -38630 9100 -38620 9135
rect -38585 9100 -38575 9135
rect -38540 9100 -38530 9135
rect -38495 9100 -38485 9135
rect -38450 9100 -38440 9135
rect -38405 9100 -38395 9135
rect -38360 9100 -38350 9135
rect -38315 9100 -38305 9135
rect -38270 9100 -38260 9135
rect -38225 9100 -38215 9135
rect -38180 9100 -38170 9135
rect -38135 9100 -38125 9135
rect -38090 9100 -38080 9135
rect -38045 9100 -38035 9135
rect -38000 9100 -37990 9135
rect -37955 9100 -37945 9135
rect -37910 9100 -37900 9135
rect -37865 9100 -37855 9135
rect -37820 9100 -37810 9135
rect -37775 9100 -37765 9135
rect -37730 9100 -37720 9135
rect -37685 9100 -37675 9135
rect -37640 9100 -37630 9135
rect -37595 9100 -37585 9135
rect -37550 9100 -37540 9135
rect -37505 9100 -37495 9135
rect -37460 9100 -37450 9135
rect -37415 9100 -37405 9135
rect -37370 9100 -37360 9135
rect -37325 9100 -37315 9135
rect -37280 9100 -37270 9135
rect -37235 9100 -37225 9135
rect -37190 9100 -37170 9135
rect -38770 9090 -37170 9100
rect -38770 9055 -38755 9090
rect -38720 9055 -38710 9090
rect -38675 9055 -38665 9090
rect -38630 9055 -38620 9090
rect -38585 9055 -38575 9090
rect -38540 9055 -38530 9090
rect -38495 9055 -38485 9090
rect -38450 9055 -38440 9090
rect -38405 9055 -38395 9090
rect -38360 9055 -38350 9090
rect -38315 9055 -38305 9090
rect -38270 9055 -38260 9090
rect -38225 9055 -38215 9090
rect -38180 9055 -38170 9090
rect -38135 9055 -38125 9090
rect -38090 9055 -38080 9090
rect -38045 9055 -38035 9090
rect -38000 9055 -37990 9090
rect -37955 9055 -37945 9090
rect -37910 9055 -37900 9090
rect -37865 9055 -37855 9090
rect -37820 9055 -37810 9090
rect -37775 9055 -37765 9090
rect -37730 9055 -37720 9090
rect -37685 9055 -37675 9090
rect -37640 9055 -37630 9090
rect -37595 9055 -37585 9090
rect -37550 9055 -37540 9090
rect -37505 9055 -37495 9090
rect -37460 9055 -37450 9090
rect -37415 9055 -37405 9090
rect -37370 9055 -37360 9090
rect -37325 9055 -37315 9090
rect -37280 9055 -37270 9090
rect -37235 9055 -37225 9090
rect -37190 9055 -37170 9090
rect -38770 9045 -37170 9055
rect -38770 9010 -38755 9045
rect -38720 9010 -38710 9045
rect -38675 9010 -38665 9045
rect -38630 9010 -38620 9045
rect -38585 9010 -38575 9045
rect -38540 9010 -38530 9045
rect -38495 9010 -38485 9045
rect -38450 9010 -38440 9045
rect -38405 9010 -38395 9045
rect -38360 9010 -38350 9045
rect -38315 9010 -38305 9045
rect -38270 9010 -38260 9045
rect -38225 9010 -38215 9045
rect -38180 9010 -38170 9045
rect -38135 9010 -38125 9045
rect -38090 9010 -38080 9045
rect -38045 9010 -38035 9045
rect -38000 9010 -37990 9045
rect -37955 9010 -37945 9045
rect -37910 9010 -37900 9045
rect -37865 9010 -37855 9045
rect -37820 9010 -37810 9045
rect -37775 9010 -37765 9045
rect -37730 9010 -37720 9045
rect -37685 9010 -37675 9045
rect -37640 9010 -37630 9045
rect -37595 9010 -37585 9045
rect -37550 9010 -37540 9045
rect -37505 9010 -37495 9045
rect -37460 9010 -37450 9045
rect -37415 9010 -37405 9045
rect -37370 9010 -37360 9045
rect -37325 9010 -37315 9045
rect -37280 9010 -37270 9045
rect -37235 9010 -37225 9045
rect -37190 9010 -37170 9045
rect -38770 9000 -37170 9010
rect -38770 8965 -38755 9000
rect -38720 8965 -38710 9000
rect -38675 8965 -38665 9000
rect -38630 8965 -38620 9000
rect -38585 8965 -38575 9000
rect -38540 8965 -38530 9000
rect -38495 8965 -38485 9000
rect -38450 8965 -38440 9000
rect -38405 8965 -38395 9000
rect -38360 8965 -38350 9000
rect -38315 8965 -38305 9000
rect -38270 8965 -38260 9000
rect -38225 8965 -38215 9000
rect -38180 8965 -38170 9000
rect -38135 8965 -38125 9000
rect -38090 8965 -38080 9000
rect -38045 8965 -38035 9000
rect -38000 8965 -37990 9000
rect -37955 8965 -37945 9000
rect -37910 8965 -37900 9000
rect -37865 8965 -37855 9000
rect -37820 8965 -37810 9000
rect -37775 8965 -37765 9000
rect -37730 8965 -37720 9000
rect -37685 8965 -37675 9000
rect -37640 8965 -37630 9000
rect -37595 8965 -37585 9000
rect -37550 8965 -37540 9000
rect -37505 8965 -37495 9000
rect -37460 8965 -37450 9000
rect -37415 8965 -37405 9000
rect -37370 8965 -37360 9000
rect -37325 8965 -37315 9000
rect -37280 8965 -37270 9000
rect -37235 8965 -37225 9000
rect -37190 8965 -37170 9000
rect -38770 8955 -37170 8965
rect -38770 8920 -38755 8955
rect -38720 8920 -38710 8955
rect -38675 8920 -38665 8955
rect -38630 8920 -38620 8955
rect -38585 8920 -38575 8955
rect -38540 8920 -38530 8955
rect -38495 8920 -38485 8955
rect -38450 8920 -38440 8955
rect -38405 8920 -38395 8955
rect -38360 8920 -38350 8955
rect -38315 8920 -38305 8955
rect -38270 8920 -38260 8955
rect -38225 8920 -38215 8955
rect -38180 8920 -38170 8955
rect -38135 8920 -38125 8955
rect -38090 8920 -38080 8955
rect -38045 8920 -38035 8955
rect -38000 8920 -37990 8955
rect -37955 8920 -37945 8955
rect -37910 8920 -37900 8955
rect -37865 8920 -37855 8955
rect -37820 8920 -37810 8955
rect -37775 8920 -37765 8955
rect -37730 8920 -37720 8955
rect -37685 8920 -37675 8955
rect -37640 8920 -37630 8955
rect -37595 8920 -37585 8955
rect -37550 8920 -37540 8955
rect -37505 8920 -37495 8955
rect -37460 8920 -37450 8955
rect -37415 8920 -37405 8955
rect -37370 8920 -37360 8955
rect -37325 8920 -37315 8955
rect -37280 8920 -37270 8955
rect -37235 8920 -37225 8955
rect -37190 8920 -37170 8955
rect -38770 8910 -37170 8920
rect -38770 8875 -38755 8910
rect -38720 8875 -38710 8910
rect -38675 8875 -38665 8910
rect -38630 8875 -38620 8910
rect -38585 8875 -38575 8910
rect -38540 8875 -38530 8910
rect -38495 8875 -38485 8910
rect -38450 8875 -38440 8910
rect -38405 8875 -38395 8910
rect -38360 8875 -38350 8910
rect -38315 8875 -38305 8910
rect -38270 8875 -38260 8910
rect -38225 8875 -38215 8910
rect -38180 8875 -38170 8910
rect -38135 8875 -38125 8910
rect -38090 8875 -38080 8910
rect -38045 8875 -38035 8910
rect -38000 8875 -37990 8910
rect -37955 8875 -37945 8910
rect -37910 8875 -37900 8910
rect -37865 8875 -37855 8910
rect -37820 8875 -37810 8910
rect -37775 8875 -37765 8910
rect -37730 8875 -37720 8910
rect -37685 8875 -37675 8910
rect -37640 8875 -37630 8910
rect -37595 8875 -37585 8910
rect -37550 8875 -37540 8910
rect -37505 8875 -37495 8910
rect -37460 8875 -37450 8910
rect -37415 8875 -37405 8910
rect -37370 8875 -37360 8910
rect -37325 8875 -37315 8910
rect -37280 8875 -37270 8910
rect -37235 8875 -37225 8910
rect -37190 8875 -37170 8910
rect -38770 8865 -37170 8875
rect -38770 8830 -38755 8865
rect -38720 8830 -38710 8865
rect -38675 8830 -38665 8865
rect -38630 8830 -38620 8865
rect -38585 8830 -38575 8865
rect -38540 8830 -38530 8865
rect -38495 8830 -38485 8865
rect -38450 8830 -38440 8865
rect -38405 8830 -38395 8865
rect -38360 8830 -38350 8865
rect -38315 8830 -38305 8865
rect -38270 8830 -38260 8865
rect -38225 8830 -38215 8865
rect -38180 8830 -38170 8865
rect -38135 8830 -38125 8865
rect -38090 8830 -38080 8865
rect -38045 8830 -38035 8865
rect -38000 8830 -37990 8865
rect -37955 8830 -37945 8865
rect -37910 8830 -37900 8865
rect -37865 8830 -37855 8865
rect -37820 8830 -37810 8865
rect -37775 8830 -37765 8865
rect -37730 8830 -37720 8865
rect -37685 8830 -37675 8865
rect -37640 8830 -37630 8865
rect -37595 8830 -37585 8865
rect -37550 8830 -37540 8865
rect -37505 8830 -37495 8865
rect -37460 8830 -37450 8865
rect -37415 8830 -37405 8865
rect -37370 8830 -37360 8865
rect -37325 8830 -37315 8865
rect -37280 8830 -37270 8865
rect -37235 8830 -37225 8865
rect -37190 8830 -37170 8865
rect -38770 8820 -37170 8830
rect -38770 8785 -38755 8820
rect -38720 8785 -38710 8820
rect -38675 8785 -38665 8820
rect -38630 8785 -38620 8820
rect -38585 8785 -38575 8820
rect -38540 8785 -38530 8820
rect -38495 8785 -38485 8820
rect -38450 8785 -38440 8820
rect -38405 8785 -38395 8820
rect -38360 8785 -38350 8820
rect -38315 8785 -38305 8820
rect -38270 8785 -38260 8820
rect -38225 8785 -38215 8820
rect -38180 8785 -38170 8820
rect -38135 8785 -38125 8820
rect -38090 8785 -38080 8820
rect -38045 8785 -38035 8820
rect -38000 8785 -37990 8820
rect -37955 8785 -37945 8820
rect -37910 8785 -37900 8820
rect -37865 8785 -37855 8820
rect -37820 8785 -37810 8820
rect -37775 8785 -37765 8820
rect -37730 8785 -37720 8820
rect -37685 8785 -37675 8820
rect -37640 8785 -37630 8820
rect -37595 8785 -37585 8820
rect -37550 8785 -37540 8820
rect -37505 8785 -37495 8820
rect -37460 8785 -37450 8820
rect -37415 8785 -37405 8820
rect -37370 8785 -37360 8820
rect -37325 8785 -37315 8820
rect -37280 8785 -37270 8820
rect -37235 8785 -37225 8820
rect -37190 8785 -37170 8820
rect -38770 8775 -37170 8785
rect -38770 8740 -38755 8775
rect -38720 8740 -38710 8775
rect -38675 8740 -38665 8775
rect -38630 8740 -38620 8775
rect -38585 8740 -38575 8775
rect -38540 8740 -38530 8775
rect -38495 8740 -38485 8775
rect -38450 8740 -38440 8775
rect -38405 8740 -38395 8775
rect -38360 8740 -38350 8775
rect -38315 8740 -38305 8775
rect -38270 8740 -38260 8775
rect -38225 8740 -38215 8775
rect -38180 8740 -38170 8775
rect -38135 8740 -38125 8775
rect -38090 8740 -38080 8775
rect -38045 8740 -38035 8775
rect -38000 8740 -37990 8775
rect -37955 8740 -37945 8775
rect -37910 8740 -37900 8775
rect -37865 8740 -37855 8775
rect -37820 8740 -37810 8775
rect -37775 8740 -37765 8775
rect -37730 8740 -37720 8775
rect -37685 8740 -37675 8775
rect -37640 8740 -37630 8775
rect -37595 8740 -37585 8775
rect -37550 8740 -37540 8775
rect -37505 8740 -37495 8775
rect -37460 8740 -37450 8775
rect -37415 8740 -37405 8775
rect -37370 8740 -37360 8775
rect -37325 8740 -37315 8775
rect -37280 8740 -37270 8775
rect -37235 8740 -37225 8775
rect -37190 8740 -37170 8775
rect -38770 8730 -37170 8740
rect -38770 8695 -38755 8730
rect -38720 8695 -38710 8730
rect -38675 8695 -38665 8730
rect -38630 8695 -38620 8730
rect -38585 8695 -38575 8730
rect -38540 8695 -38530 8730
rect -38495 8695 -38485 8730
rect -38450 8695 -38440 8730
rect -38405 8695 -38395 8730
rect -38360 8695 -38350 8730
rect -38315 8695 -38305 8730
rect -38270 8695 -38260 8730
rect -38225 8695 -38215 8730
rect -38180 8695 -38170 8730
rect -38135 8695 -38125 8730
rect -38090 8695 -38080 8730
rect -38045 8695 -38035 8730
rect -38000 8695 -37990 8730
rect -37955 8695 -37945 8730
rect -37910 8695 -37900 8730
rect -37865 8695 -37855 8730
rect -37820 8695 -37810 8730
rect -37775 8695 -37765 8730
rect -37730 8695 -37720 8730
rect -37685 8695 -37675 8730
rect -37640 8695 -37630 8730
rect -37595 8695 -37585 8730
rect -37550 8695 -37540 8730
rect -37505 8695 -37495 8730
rect -37460 8695 -37450 8730
rect -37415 8695 -37405 8730
rect -37370 8695 -37360 8730
rect -37325 8695 -37315 8730
rect -37280 8695 -37270 8730
rect -37235 8695 -37225 8730
rect -37190 8695 -37170 8730
rect -38770 8685 -37170 8695
rect -38770 8650 -38755 8685
rect -38720 8650 -38710 8685
rect -38675 8650 -38665 8685
rect -38630 8650 -38620 8685
rect -38585 8650 -38575 8685
rect -38540 8650 -38530 8685
rect -38495 8650 -38485 8685
rect -38450 8650 -38440 8685
rect -38405 8650 -38395 8685
rect -38360 8650 -38350 8685
rect -38315 8650 -38305 8685
rect -38270 8650 -38260 8685
rect -38225 8650 -38215 8685
rect -38180 8650 -38170 8685
rect -38135 8650 -38125 8685
rect -38090 8650 -38080 8685
rect -38045 8650 -38035 8685
rect -38000 8650 -37990 8685
rect -37955 8650 -37945 8685
rect -37910 8650 -37900 8685
rect -37865 8650 -37855 8685
rect -37820 8650 -37810 8685
rect -37775 8650 -37765 8685
rect -37730 8650 -37720 8685
rect -37685 8650 -37675 8685
rect -37640 8650 -37630 8685
rect -37595 8650 -37585 8685
rect -37550 8650 -37540 8685
rect -37505 8650 -37495 8685
rect -37460 8650 -37450 8685
rect -37415 8650 -37405 8685
rect -37370 8650 -37360 8685
rect -37325 8650 -37315 8685
rect -37280 8650 -37270 8685
rect -37235 8650 -37225 8685
rect -37190 8650 -37170 8685
rect -38770 8640 -37170 8650
rect -38770 8605 -38755 8640
rect -38720 8605 -38710 8640
rect -38675 8605 -38665 8640
rect -38630 8605 -38620 8640
rect -38585 8605 -38575 8640
rect -38540 8605 -38530 8640
rect -38495 8605 -38485 8640
rect -38450 8605 -38440 8640
rect -38405 8605 -38395 8640
rect -38360 8605 -38350 8640
rect -38315 8605 -38305 8640
rect -38270 8605 -38260 8640
rect -38225 8605 -38215 8640
rect -38180 8605 -38170 8640
rect -38135 8605 -38125 8640
rect -38090 8605 -38080 8640
rect -38045 8605 -38035 8640
rect -38000 8605 -37990 8640
rect -37955 8605 -37945 8640
rect -37910 8605 -37900 8640
rect -37865 8605 -37855 8640
rect -37820 8605 -37810 8640
rect -37775 8605 -37765 8640
rect -37730 8605 -37720 8640
rect -37685 8605 -37675 8640
rect -37640 8605 -37630 8640
rect -37595 8605 -37585 8640
rect -37550 8605 -37540 8640
rect -37505 8605 -37495 8640
rect -37460 8605 -37450 8640
rect -37415 8605 -37405 8640
rect -37370 8605 -37360 8640
rect -37325 8605 -37315 8640
rect -37280 8605 -37270 8640
rect -37235 8605 -37225 8640
rect -37190 8605 -37170 8640
rect -38770 8595 -37170 8605
rect -38770 8560 -38755 8595
rect -38720 8560 -38710 8595
rect -38675 8560 -38665 8595
rect -38630 8560 -38620 8595
rect -38585 8560 -38575 8595
rect -38540 8560 -38530 8595
rect -38495 8560 -38485 8595
rect -38450 8560 -38440 8595
rect -38405 8560 -38395 8595
rect -38360 8560 -38350 8595
rect -38315 8560 -38305 8595
rect -38270 8560 -38260 8595
rect -38225 8560 -38215 8595
rect -38180 8560 -38170 8595
rect -38135 8560 -38125 8595
rect -38090 8560 -38080 8595
rect -38045 8560 -38035 8595
rect -38000 8560 -37990 8595
rect -37955 8560 -37945 8595
rect -37910 8560 -37900 8595
rect -37865 8560 -37855 8595
rect -37820 8560 -37810 8595
rect -37775 8560 -37765 8595
rect -37730 8560 -37720 8595
rect -37685 8560 -37675 8595
rect -37640 8560 -37630 8595
rect -37595 8560 -37585 8595
rect -37550 8560 -37540 8595
rect -37505 8560 -37495 8595
rect -37460 8560 -37450 8595
rect -37415 8560 -37405 8595
rect -37370 8560 -37360 8595
rect -37325 8560 -37315 8595
rect -37280 8560 -37270 8595
rect -37235 8560 -37225 8595
rect -37190 8560 -37170 8595
rect -38770 8550 -37170 8560
rect -38770 8515 -38755 8550
rect -38720 8515 -38710 8550
rect -38675 8515 -38665 8550
rect -38630 8515 -38620 8550
rect -38585 8515 -38575 8550
rect -38540 8515 -38530 8550
rect -38495 8515 -38485 8550
rect -38450 8515 -38440 8550
rect -38405 8515 -38395 8550
rect -38360 8515 -38350 8550
rect -38315 8515 -38305 8550
rect -38270 8515 -38260 8550
rect -38225 8515 -38215 8550
rect -38180 8515 -38170 8550
rect -38135 8515 -38125 8550
rect -38090 8515 -38080 8550
rect -38045 8515 -38035 8550
rect -38000 8515 -37990 8550
rect -37955 8515 -37945 8550
rect -37910 8515 -37900 8550
rect -37865 8515 -37855 8550
rect -37820 8515 -37810 8550
rect -37775 8515 -37765 8550
rect -37730 8515 -37720 8550
rect -37685 8515 -37675 8550
rect -37640 8515 -37630 8550
rect -37595 8515 -37585 8550
rect -37550 8515 -37540 8550
rect -37505 8515 -37495 8550
rect -37460 8515 -37450 8550
rect -37415 8515 -37405 8550
rect -37370 8515 -37360 8550
rect -37325 8515 -37315 8550
rect -37280 8515 -37270 8550
rect -37235 8515 -37225 8550
rect -37190 8515 -37170 8550
rect -38770 8505 -37170 8515
rect -38770 8470 -38755 8505
rect -38720 8470 -38710 8505
rect -38675 8470 -38665 8505
rect -38630 8470 -38620 8505
rect -38585 8470 -38575 8505
rect -38540 8470 -38530 8505
rect -38495 8470 -38485 8505
rect -38450 8470 -38440 8505
rect -38405 8470 -38395 8505
rect -38360 8470 -38350 8505
rect -38315 8470 -38305 8505
rect -38270 8470 -38260 8505
rect -38225 8470 -38215 8505
rect -38180 8470 -38170 8505
rect -38135 8470 -38125 8505
rect -38090 8470 -38080 8505
rect -38045 8470 -38035 8505
rect -38000 8470 -37990 8505
rect -37955 8470 -37945 8505
rect -37910 8470 -37900 8505
rect -37865 8470 -37855 8505
rect -37820 8470 -37810 8505
rect -37775 8470 -37765 8505
rect -37730 8470 -37720 8505
rect -37685 8470 -37675 8505
rect -37640 8470 -37630 8505
rect -37595 8470 -37585 8505
rect -37550 8470 -37540 8505
rect -37505 8470 -37495 8505
rect -37460 8470 -37450 8505
rect -37415 8470 -37405 8505
rect -37370 8470 -37360 8505
rect -37325 8470 -37315 8505
rect -37280 8470 -37270 8505
rect -37235 8470 -37225 8505
rect -37190 8470 -37170 8505
rect -38770 8460 -37170 8470
rect -38770 8425 -38755 8460
rect -38720 8425 -38710 8460
rect -38675 8425 -38665 8460
rect -38630 8425 -38620 8460
rect -38585 8425 -38575 8460
rect -38540 8425 -38530 8460
rect -38495 8425 -38485 8460
rect -38450 8425 -38440 8460
rect -38405 8425 -38395 8460
rect -38360 8425 -38350 8460
rect -38315 8425 -38305 8460
rect -38270 8425 -38260 8460
rect -38225 8425 -38215 8460
rect -38180 8425 -38170 8460
rect -38135 8425 -38125 8460
rect -38090 8425 -38080 8460
rect -38045 8425 -38035 8460
rect -38000 8425 -37990 8460
rect -37955 8425 -37945 8460
rect -37910 8425 -37900 8460
rect -37865 8425 -37855 8460
rect -37820 8425 -37810 8460
rect -37775 8425 -37765 8460
rect -37730 8425 -37720 8460
rect -37685 8425 -37675 8460
rect -37640 8425 -37630 8460
rect -37595 8425 -37585 8460
rect -37550 8425 -37540 8460
rect -37505 8425 -37495 8460
rect -37460 8425 -37450 8460
rect -37415 8425 -37405 8460
rect -37370 8425 -37360 8460
rect -37325 8425 -37315 8460
rect -37280 8425 -37270 8460
rect -37235 8425 -37225 8460
rect -37190 8425 -37170 8460
rect -38770 8415 -37170 8425
rect -38770 8380 -38755 8415
rect -38720 8380 -38710 8415
rect -38675 8380 -38665 8415
rect -38630 8380 -38620 8415
rect -38585 8380 -38575 8415
rect -38540 8380 -38530 8415
rect -38495 8380 -38485 8415
rect -38450 8380 -38440 8415
rect -38405 8380 -38395 8415
rect -38360 8380 -38350 8415
rect -38315 8380 -38305 8415
rect -38270 8380 -38260 8415
rect -38225 8380 -38215 8415
rect -38180 8380 -38170 8415
rect -38135 8380 -38125 8415
rect -38090 8380 -38080 8415
rect -38045 8380 -38035 8415
rect -38000 8380 -37990 8415
rect -37955 8380 -37945 8415
rect -37910 8380 -37900 8415
rect -37865 8380 -37855 8415
rect -37820 8380 -37810 8415
rect -37775 8380 -37765 8415
rect -37730 8380 -37720 8415
rect -37685 8380 -37675 8415
rect -37640 8380 -37630 8415
rect -37595 8380 -37585 8415
rect -37550 8380 -37540 8415
rect -37505 8380 -37495 8415
rect -37460 8380 -37450 8415
rect -37415 8380 -37405 8415
rect -37370 8380 -37360 8415
rect -37325 8380 -37315 8415
rect -37280 8380 -37270 8415
rect -37235 8380 -37225 8415
rect -37190 8380 -37170 8415
rect -38770 8370 -37170 8380
rect -38770 8335 -38755 8370
rect -38720 8335 -38710 8370
rect -38675 8335 -38665 8370
rect -38630 8335 -38620 8370
rect -38585 8335 -38575 8370
rect -38540 8335 -38530 8370
rect -38495 8335 -38485 8370
rect -38450 8335 -38440 8370
rect -38405 8335 -38395 8370
rect -38360 8335 -38350 8370
rect -38315 8335 -38305 8370
rect -38270 8335 -38260 8370
rect -38225 8335 -38215 8370
rect -38180 8335 -38170 8370
rect -38135 8335 -38125 8370
rect -38090 8335 -38080 8370
rect -38045 8335 -38035 8370
rect -38000 8335 -37990 8370
rect -37955 8335 -37945 8370
rect -37910 8335 -37900 8370
rect -37865 8335 -37855 8370
rect -37820 8335 -37810 8370
rect -37775 8335 -37765 8370
rect -37730 8335 -37720 8370
rect -37685 8335 -37675 8370
rect -37640 8335 -37630 8370
rect -37595 8335 -37585 8370
rect -37550 8335 -37540 8370
rect -37505 8335 -37495 8370
rect -37460 8335 -37450 8370
rect -37415 8335 -37405 8370
rect -37370 8335 -37360 8370
rect -37325 8335 -37315 8370
rect -37280 8335 -37270 8370
rect -37235 8335 -37225 8370
rect -37190 8335 -37170 8370
rect -38770 8325 -37170 8335
rect -38770 8290 -38755 8325
rect -38720 8290 -38710 8325
rect -38675 8290 -38665 8325
rect -38630 8290 -38620 8325
rect -38585 8290 -38575 8325
rect -38540 8290 -38530 8325
rect -38495 8290 -38485 8325
rect -38450 8290 -38440 8325
rect -38405 8290 -38395 8325
rect -38360 8290 -38350 8325
rect -38315 8290 -38305 8325
rect -38270 8290 -38260 8325
rect -38225 8290 -38215 8325
rect -38180 8290 -38170 8325
rect -38135 8290 -38125 8325
rect -38090 8290 -38080 8325
rect -38045 8290 -38035 8325
rect -38000 8290 -37990 8325
rect -37955 8290 -37945 8325
rect -37910 8290 -37900 8325
rect -37865 8290 -37855 8325
rect -37820 8290 -37810 8325
rect -37775 8290 -37765 8325
rect -37730 8290 -37720 8325
rect -37685 8290 -37675 8325
rect -37640 8290 -37630 8325
rect -37595 8290 -37585 8325
rect -37550 8290 -37540 8325
rect -37505 8290 -37495 8325
rect -37460 8290 -37450 8325
rect -37415 8290 -37405 8325
rect -37370 8290 -37360 8325
rect -37325 8290 -37315 8325
rect -37280 8290 -37270 8325
rect -37235 8290 -37225 8325
rect -37190 8290 -37170 8325
rect -38770 8280 -37170 8290
rect -38770 8245 -38755 8280
rect -38720 8245 -38710 8280
rect -38675 8245 -38665 8280
rect -38630 8245 -38620 8280
rect -38585 8245 -38575 8280
rect -38540 8245 -38530 8280
rect -38495 8245 -38485 8280
rect -38450 8245 -38440 8280
rect -38405 8245 -38395 8280
rect -38360 8245 -38350 8280
rect -38315 8245 -38305 8280
rect -38270 8245 -38260 8280
rect -38225 8245 -38215 8280
rect -38180 8245 -38170 8280
rect -38135 8245 -38125 8280
rect -38090 8245 -38080 8280
rect -38045 8245 -38035 8280
rect -38000 8245 -37990 8280
rect -37955 8245 -37945 8280
rect -37910 8245 -37900 8280
rect -37865 8245 -37855 8280
rect -37820 8245 -37810 8280
rect -37775 8245 -37765 8280
rect -37730 8245 -37720 8280
rect -37685 8245 -37675 8280
rect -37640 8245 -37630 8280
rect -37595 8245 -37585 8280
rect -37550 8245 -37540 8280
rect -37505 8245 -37495 8280
rect -37460 8245 -37450 8280
rect -37415 8245 -37405 8280
rect -37370 8245 -37360 8280
rect -37325 8245 -37315 8280
rect -37280 8245 -37270 8280
rect -37235 8245 -37225 8280
rect -37190 8245 -37170 8280
rect -38770 8235 -37170 8245
rect -38770 8200 -38755 8235
rect -38720 8200 -38710 8235
rect -38675 8200 -38665 8235
rect -38630 8200 -38620 8235
rect -38585 8200 -38575 8235
rect -38540 8200 -38530 8235
rect -38495 8200 -38485 8235
rect -38450 8200 -38440 8235
rect -38405 8200 -38395 8235
rect -38360 8200 -38350 8235
rect -38315 8200 -38305 8235
rect -38270 8200 -38260 8235
rect -38225 8200 -38215 8235
rect -38180 8200 -38170 8235
rect -38135 8200 -38125 8235
rect -38090 8200 -38080 8235
rect -38045 8200 -38035 8235
rect -38000 8200 -37990 8235
rect -37955 8200 -37945 8235
rect -37910 8200 -37900 8235
rect -37865 8200 -37855 8235
rect -37820 8200 -37810 8235
rect -37775 8200 -37765 8235
rect -37730 8200 -37720 8235
rect -37685 8200 -37675 8235
rect -37640 8200 -37630 8235
rect -37595 8200 -37585 8235
rect -37550 8200 -37540 8235
rect -37505 8200 -37495 8235
rect -37460 8200 -37450 8235
rect -37415 8200 -37405 8235
rect -37370 8200 -37360 8235
rect -37325 8200 -37315 8235
rect -37280 8200 -37270 8235
rect -37235 8200 -37225 8235
rect -37190 8200 -37170 8235
rect -38770 8190 -37170 8200
rect -38770 8155 -38755 8190
rect -38720 8155 -38710 8190
rect -38675 8155 -38665 8190
rect -38630 8155 -38620 8190
rect -38585 8155 -38575 8190
rect -38540 8155 -38530 8190
rect -38495 8155 -38485 8190
rect -38450 8155 -38440 8190
rect -38405 8155 -38395 8190
rect -38360 8155 -38350 8190
rect -38315 8155 -38305 8190
rect -38270 8155 -38260 8190
rect -38225 8155 -38215 8190
rect -38180 8155 -38170 8190
rect -38135 8155 -38125 8190
rect -38090 8155 -38080 8190
rect -38045 8155 -38035 8190
rect -38000 8155 -37990 8190
rect -37955 8155 -37945 8190
rect -37910 8155 -37900 8190
rect -37865 8155 -37855 8190
rect -37820 8155 -37810 8190
rect -37775 8155 -37765 8190
rect -37730 8155 -37720 8190
rect -37685 8155 -37675 8190
rect -37640 8155 -37630 8190
rect -37595 8155 -37585 8190
rect -37550 8155 -37540 8190
rect -37505 8155 -37495 8190
rect -37460 8155 -37450 8190
rect -37415 8155 -37405 8190
rect -37370 8155 -37360 8190
rect -37325 8155 -37315 8190
rect -37280 8155 -37270 8190
rect -37235 8155 -37225 8190
rect -37190 8155 -37170 8190
rect -38770 8145 -37170 8155
rect -38770 8110 -38755 8145
rect -38720 8110 -38710 8145
rect -38675 8110 -38665 8145
rect -38630 8110 -38620 8145
rect -38585 8110 -38575 8145
rect -38540 8110 -38530 8145
rect -38495 8110 -38485 8145
rect -38450 8110 -38440 8145
rect -38405 8110 -38395 8145
rect -38360 8110 -38350 8145
rect -38315 8110 -38305 8145
rect -38270 8110 -38260 8145
rect -38225 8110 -38215 8145
rect -38180 8110 -38170 8145
rect -38135 8110 -38125 8145
rect -38090 8110 -38080 8145
rect -38045 8110 -38035 8145
rect -38000 8110 -37990 8145
rect -37955 8110 -37945 8145
rect -37910 8110 -37900 8145
rect -37865 8110 -37855 8145
rect -37820 8110 -37810 8145
rect -37775 8110 -37765 8145
rect -37730 8110 -37720 8145
rect -37685 8110 -37675 8145
rect -37640 8110 -37630 8145
rect -37595 8110 -37585 8145
rect -37550 8110 -37540 8145
rect -37505 8110 -37495 8145
rect -37460 8110 -37450 8145
rect -37415 8110 -37405 8145
rect -37370 8110 -37360 8145
rect -37325 8110 -37315 8145
rect -37280 8110 -37270 8145
rect -37235 8110 -37225 8145
rect -37190 8110 -37170 8145
rect -38770 8105 -37170 8110
rect 1310 9640 1370 9650
rect 1310 9600 1320 9640
rect 1360 9600 1370 9640
rect 1310 9575 1370 9600
rect 1310 9535 1320 9575
rect 1360 9535 1370 9575
rect 1310 9505 1370 9535
rect 1310 9465 1320 9505
rect 1360 9465 1370 9505
rect 1310 9435 1370 9465
rect 1310 9395 1320 9435
rect 1360 9395 1370 9435
rect 1310 9365 1370 9395
rect 1310 9325 1320 9365
rect 1360 9325 1370 9365
rect 1310 9300 1370 9325
rect 1310 9260 1320 9300
rect 1360 9260 1370 9300
rect 1310 9240 1370 9260
rect 1310 9200 1320 9240
rect 1360 9200 1370 9240
rect 1310 9175 1370 9200
rect 1310 9135 1320 9175
rect 1360 9135 1370 9175
rect 1310 9105 1370 9135
rect 1310 9065 1320 9105
rect 1360 9065 1370 9105
rect 1310 9035 1370 9065
rect 1310 8995 1320 9035
rect 1360 8995 1370 9035
rect 1310 8965 1370 8995
rect 1310 8925 1320 8965
rect 1360 8925 1370 8965
rect 1310 8900 1370 8925
rect 1310 8860 1320 8900
rect 1360 8860 1370 8900
rect 1310 8840 1370 8860
rect 1310 8800 1320 8840
rect 1360 8800 1370 8840
rect 1310 8775 1370 8800
rect 1310 8735 1320 8775
rect 1360 8735 1370 8775
rect 1310 8705 1370 8735
rect 1310 8665 1320 8705
rect 1360 8665 1370 8705
rect 1310 8635 1370 8665
rect 1310 8595 1320 8635
rect 1360 8595 1370 8635
rect 1310 8565 1370 8595
rect 1310 8525 1320 8565
rect 1360 8525 1370 8565
rect 1310 8500 1370 8525
rect 1310 8460 1320 8500
rect 1360 8460 1370 8500
rect 1310 8440 1370 8460
rect 1310 8400 1320 8440
rect 1360 8400 1370 8440
rect 1310 8375 1370 8400
rect 1310 8335 1320 8375
rect 1360 8335 1370 8375
rect 1310 8305 1370 8335
rect 1310 8265 1320 8305
rect 1360 8265 1370 8305
rect 1310 8235 1370 8265
rect 1310 8195 1320 8235
rect 1360 8195 1370 8235
rect 1310 8165 1370 8195
rect 1310 8125 1320 8165
rect 1360 8125 1370 8165
rect 1310 8105 1370 8125
rect 2235 9640 2295 9650
rect 2235 9600 2245 9640
rect 2285 9600 2295 9640
rect 2235 9575 2295 9600
rect 2235 9535 2245 9575
rect 2285 9535 2295 9575
rect 2235 9505 2295 9535
rect 2235 9465 2245 9505
rect 2285 9465 2295 9505
rect 2235 9435 2295 9465
rect 2235 9395 2245 9435
rect 2285 9395 2295 9435
rect 2235 9365 2295 9395
rect 2235 9325 2245 9365
rect 2285 9325 2295 9365
rect 2235 9300 2295 9325
rect 2235 9260 2245 9300
rect 2285 9260 2295 9300
rect 2235 9240 2295 9260
rect 2235 9200 2245 9240
rect 2285 9200 2295 9240
rect 2235 9175 2295 9200
rect 2235 9135 2245 9175
rect 2285 9135 2295 9175
rect 2235 9105 2295 9135
rect 2235 9065 2245 9105
rect 2285 9065 2295 9105
rect 2235 9035 2295 9065
rect 2235 8995 2245 9035
rect 2285 8995 2295 9035
rect 2235 8965 2295 8995
rect 2235 8925 2245 8965
rect 2285 8925 2295 8965
rect 2235 8900 2295 8925
rect 2235 8860 2245 8900
rect 2285 8860 2295 8900
rect 2235 8840 2295 8860
rect 2235 8800 2245 8840
rect 2285 8800 2295 8840
rect 2235 8775 2295 8800
rect 2235 8735 2245 8775
rect 2285 8735 2295 8775
rect 2235 8705 2295 8735
rect 2235 8665 2245 8705
rect 2285 8665 2295 8705
rect 2235 8635 2295 8665
rect 2235 8595 2245 8635
rect 2285 8595 2295 8635
rect 2235 8565 2295 8595
rect 2235 8525 2245 8565
rect 2285 8525 2295 8565
rect 2235 8500 2295 8525
rect 2235 8460 2245 8500
rect 2285 8460 2295 8500
rect 2235 8440 2295 8460
rect 2235 8400 2245 8440
rect 2285 8400 2295 8440
rect 2235 8375 2295 8400
rect 2235 8335 2245 8375
rect 2285 8335 2295 8375
rect 2235 8305 2295 8335
rect 2235 8265 2245 8305
rect 2285 8265 2295 8305
rect 2235 8235 2295 8265
rect 2235 8195 2245 8235
rect 2285 8195 2295 8235
rect 2235 8165 2295 8195
rect 2235 8125 2245 8165
rect 2285 8125 2295 8165
rect 2235 8105 2295 8125
rect 6690 9640 6750 9650
rect 6690 9600 6700 9640
rect 6740 9600 6750 9640
rect 6690 9575 6750 9600
rect 6690 9535 6700 9575
rect 6740 9535 6750 9575
rect 6690 9505 6750 9535
rect 6690 9465 6700 9505
rect 6740 9465 6750 9505
rect 6690 9435 6750 9465
rect 6690 9395 6700 9435
rect 6740 9395 6750 9435
rect 6690 9365 6750 9395
rect 6690 9325 6700 9365
rect 6740 9325 6750 9365
rect 6690 9300 6750 9325
rect 6690 9260 6700 9300
rect 6740 9260 6750 9300
rect 6690 9240 6750 9260
rect 6690 9200 6700 9240
rect 6740 9200 6750 9240
rect 6690 9175 6750 9200
rect 6690 9135 6700 9175
rect 6740 9135 6750 9175
rect 6690 9105 6750 9135
rect 6690 9065 6700 9105
rect 6740 9065 6750 9105
rect 6690 9035 6750 9065
rect 6690 8995 6700 9035
rect 6740 8995 6750 9035
rect 6690 8965 6750 8995
rect 6690 8925 6700 8965
rect 6740 8925 6750 8965
rect 6690 8900 6750 8925
rect 6690 8860 6700 8900
rect 6740 8860 6750 8900
rect 6690 8840 6750 8860
rect 6690 8800 6700 8840
rect 6740 8800 6750 8840
rect 6690 8775 6750 8800
rect 6690 8735 6700 8775
rect 6740 8735 6750 8775
rect 6690 8705 6750 8735
rect 6690 8665 6700 8705
rect 6740 8665 6750 8705
rect 6690 8635 6750 8665
rect 6690 8595 6700 8635
rect 6740 8595 6750 8635
rect 6690 8565 6750 8595
rect 6690 8525 6700 8565
rect 6740 8525 6750 8565
rect 6690 8500 6750 8525
rect 6690 8460 6700 8500
rect 6740 8460 6750 8500
rect 6690 8440 6750 8460
rect 6690 8400 6700 8440
rect 6740 8400 6750 8440
rect 6690 8375 6750 8400
rect 6690 8335 6700 8375
rect 6740 8335 6750 8375
rect 6690 8305 6750 8335
rect 6690 8265 6700 8305
rect 6740 8265 6750 8305
rect 6690 8235 6750 8265
rect 6690 8195 6700 8235
rect 6740 8195 6750 8235
rect 6690 8165 6750 8195
rect 6690 8125 6700 8165
rect 6740 8125 6750 8165
rect 6690 8105 6750 8125
rect 7610 9640 7670 9650
rect 7610 9600 7620 9640
rect 7660 9600 7670 9640
rect 7610 9575 7670 9600
rect 7610 9535 7620 9575
rect 7660 9535 7670 9575
rect 7610 9505 7670 9535
rect 7610 9465 7620 9505
rect 7660 9465 7670 9505
rect 7610 9435 7670 9465
rect 7610 9395 7620 9435
rect 7660 9395 7670 9435
rect 7610 9365 7670 9395
rect 7610 9325 7620 9365
rect 7660 9325 7670 9365
rect 7610 9300 7670 9325
rect 7610 9260 7620 9300
rect 7660 9260 7670 9300
rect 7610 9240 7670 9260
rect 7610 9200 7620 9240
rect 7660 9200 7670 9240
rect 7610 9175 7670 9200
rect 7610 9135 7620 9175
rect 7660 9135 7670 9175
rect 7610 9105 7670 9135
rect 7610 9065 7620 9105
rect 7660 9065 7670 9105
rect 7610 9035 7670 9065
rect 7610 8995 7620 9035
rect 7660 8995 7670 9035
rect 7610 8965 7670 8995
rect 7610 8925 7620 8965
rect 7660 8925 7670 8965
rect 7610 8900 7670 8925
rect 7610 8860 7620 8900
rect 7660 8860 7670 8900
rect 7610 8840 7670 8860
rect 7610 8800 7620 8840
rect 7660 8800 7670 8840
rect 7610 8775 7670 8800
rect 7610 8735 7620 8775
rect 7660 8735 7670 8775
rect 7610 8705 7670 8735
rect 7610 8665 7620 8705
rect 7660 8665 7670 8705
rect 7610 8635 7670 8665
rect 7610 8595 7620 8635
rect 7660 8595 7670 8635
rect 7610 8565 7670 8595
rect 7610 8525 7620 8565
rect 7660 8525 7670 8565
rect 7610 8500 7670 8525
rect 7610 8460 7620 8500
rect 7660 8460 7670 8500
rect 7610 8440 7670 8460
rect 7610 8400 7620 8440
rect 7660 8400 7670 8440
rect 7610 8375 7670 8400
rect 7610 8335 7620 8375
rect 7660 8335 7670 8375
rect 7610 8305 7670 8335
rect 7610 8265 7620 8305
rect 7660 8265 7670 8305
rect 7610 8235 7670 8265
rect 7610 8195 7620 8235
rect 7660 8195 7670 8235
rect 7610 8165 7670 8195
rect 7610 8125 7620 8165
rect 7660 8125 7670 8165
rect 7610 8105 7670 8125
rect 31290 8030 32890 17740
rect 31290 7995 31305 8030
rect 31340 7995 31350 8030
rect 31385 7995 31395 8030
rect 31430 7995 31440 8030
rect 31475 7995 31485 8030
rect 31520 7995 31530 8030
rect 31565 7995 31575 8030
rect 31610 7995 31620 8030
rect 31655 7995 31665 8030
rect 31700 7995 31710 8030
rect 31745 7995 31755 8030
rect 31790 7995 31800 8030
rect 31835 7995 31845 8030
rect 31880 7995 31890 8030
rect 31925 7995 31935 8030
rect 31970 7995 31980 8030
rect 32015 7995 32025 8030
rect 32060 7995 32070 8030
rect 32105 7995 32115 8030
rect 32150 7995 32160 8030
rect 32195 7995 32205 8030
rect 32240 7995 32250 8030
rect 32285 7995 32295 8030
rect 32330 7995 32340 8030
rect 32375 7995 32385 8030
rect 32420 7995 32430 8030
rect 32465 7995 32475 8030
rect 32510 7995 32520 8030
rect 32555 7995 32565 8030
rect 32600 7995 32610 8030
rect 32645 7995 32655 8030
rect 32690 7995 32700 8030
rect 32735 7995 32745 8030
rect 32780 7995 32790 8030
rect 32825 7995 32835 8030
rect 32870 7995 32890 8030
rect 31290 7985 32890 7995
rect -38770 7970 -37170 7980
rect -38770 7935 -38755 7970
rect -38720 7935 -38710 7970
rect -38675 7935 -38665 7970
rect -38630 7935 -38620 7970
rect -38585 7935 -38575 7970
rect -38540 7935 -38530 7970
rect -38495 7935 -38485 7970
rect -38450 7935 -38440 7970
rect -38405 7935 -38395 7970
rect -38360 7935 -38350 7970
rect -38315 7935 -38305 7970
rect -38270 7935 -38260 7970
rect -38225 7935 -38215 7970
rect -38180 7935 -38170 7970
rect -38135 7935 -38125 7970
rect -38090 7935 -38080 7970
rect -38045 7935 -38035 7970
rect -38000 7935 -37990 7970
rect -37955 7935 -37945 7970
rect -37910 7935 -37900 7970
rect -37865 7935 -37855 7970
rect -37820 7935 -37810 7970
rect -37775 7935 -37765 7970
rect -37730 7935 -37720 7970
rect -37685 7935 -37675 7970
rect -37640 7935 -37630 7970
rect -37595 7935 -37585 7970
rect -37550 7935 -37540 7970
rect -37505 7935 -37495 7970
rect -37460 7935 -37450 7970
rect -37415 7935 -37405 7970
rect -37370 7935 -37360 7970
rect -37325 7935 -37315 7970
rect -37280 7935 -37270 7970
rect -37235 7935 -37225 7970
rect -37190 7935 -37170 7970
rect -38770 7925 -37170 7935
rect -38770 7890 -38755 7925
rect -38720 7890 -38710 7925
rect -38675 7890 -38665 7925
rect -38630 7890 -38620 7925
rect -38585 7890 -38575 7925
rect -38540 7890 -38530 7925
rect -38495 7890 -38485 7925
rect -38450 7890 -38440 7925
rect -38405 7890 -38395 7925
rect -38360 7890 -38350 7925
rect -38315 7890 -38305 7925
rect -38270 7890 -38260 7925
rect -38225 7890 -38215 7925
rect -38180 7890 -38170 7925
rect -38135 7890 -38125 7925
rect -38090 7890 -38080 7925
rect -38045 7890 -38035 7925
rect -38000 7890 -37990 7925
rect -37955 7890 -37945 7925
rect -37910 7890 -37900 7925
rect -37865 7890 -37855 7925
rect -37820 7890 -37810 7925
rect -37775 7890 -37765 7925
rect -37730 7890 -37720 7925
rect -37685 7890 -37675 7925
rect -37640 7890 -37630 7925
rect -37595 7890 -37585 7925
rect -37550 7890 -37540 7925
rect -37505 7890 -37495 7925
rect -37460 7890 -37450 7925
rect -37415 7890 -37405 7925
rect -37370 7890 -37360 7925
rect -37325 7890 -37315 7925
rect -37280 7890 -37270 7925
rect -37235 7890 -37225 7925
rect -37190 7890 -37170 7925
rect -38770 7880 -37170 7890
rect -38770 7845 -38755 7880
rect -38720 7845 -38710 7880
rect -38675 7845 -38665 7880
rect -38630 7845 -38620 7880
rect -38585 7845 -38575 7880
rect -38540 7845 -38530 7880
rect -38495 7845 -38485 7880
rect -38450 7845 -38440 7880
rect -38405 7845 -38395 7880
rect -38360 7845 -38350 7880
rect -38315 7845 -38305 7880
rect -38270 7845 -38260 7880
rect -38225 7845 -38215 7880
rect -38180 7845 -38170 7880
rect -38135 7845 -38125 7880
rect -38090 7845 -38080 7880
rect -38045 7845 -38035 7880
rect -38000 7845 -37990 7880
rect -37955 7845 -37945 7880
rect -37910 7845 -37900 7880
rect -37865 7845 -37855 7880
rect -37820 7845 -37810 7880
rect -37775 7845 -37765 7880
rect -37730 7845 -37720 7880
rect -37685 7845 -37675 7880
rect -37640 7845 -37630 7880
rect -37595 7845 -37585 7880
rect -37550 7845 -37540 7880
rect -37505 7845 -37495 7880
rect -37460 7845 -37450 7880
rect -37415 7845 -37405 7880
rect -37370 7845 -37360 7880
rect -37325 7845 -37315 7880
rect -37280 7845 -37270 7880
rect -37235 7845 -37225 7880
rect -37190 7845 -37170 7880
rect -38770 7835 -37170 7845
rect -38770 7800 -38755 7835
rect -38720 7800 -38710 7835
rect -38675 7800 -38665 7835
rect -38630 7800 -38620 7835
rect -38585 7800 -38575 7835
rect -38540 7800 -38530 7835
rect -38495 7800 -38485 7835
rect -38450 7800 -38440 7835
rect -38405 7800 -38395 7835
rect -38360 7800 -38350 7835
rect -38315 7800 -38305 7835
rect -38270 7800 -38260 7835
rect -38225 7800 -38215 7835
rect -38180 7800 -38170 7835
rect -38135 7800 -38125 7835
rect -38090 7800 -38080 7835
rect -38045 7800 -38035 7835
rect -38000 7800 -37990 7835
rect -37955 7800 -37945 7835
rect -37910 7800 -37900 7835
rect -37865 7800 -37855 7835
rect -37820 7800 -37810 7835
rect -37775 7800 -37765 7835
rect -37730 7800 -37720 7835
rect -37685 7800 -37675 7835
rect -37640 7800 -37630 7835
rect -37595 7800 -37585 7835
rect -37550 7800 -37540 7835
rect -37505 7800 -37495 7835
rect -37460 7800 -37450 7835
rect -37415 7800 -37405 7835
rect -37370 7800 -37360 7835
rect -37325 7800 -37315 7835
rect -37280 7800 -37270 7835
rect -37235 7800 -37225 7835
rect -37190 7800 -37170 7835
rect -38770 7790 -37170 7800
rect -38770 7755 -38755 7790
rect -38720 7755 -38710 7790
rect -38675 7755 -38665 7790
rect -38630 7755 -38620 7790
rect -38585 7755 -38575 7790
rect -38540 7755 -38530 7790
rect -38495 7755 -38485 7790
rect -38450 7755 -38440 7790
rect -38405 7755 -38395 7790
rect -38360 7755 -38350 7790
rect -38315 7755 -38305 7790
rect -38270 7755 -38260 7790
rect -38225 7755 -38215 7790
rect -38180 7755 -38170 7790
rect -38135 7755 -38125 7790
rect -38090 7755 -38080 7790
rect -38045 7755 -38035 7790
rect -38000 7755 -37990 7790
rect -37955 7755 -37945 7790
rect -37910 7755 -37900 7790
rect -37865 7755 -37855 7790
rect -37820 7755 -37810 7790
rect -37775 7755 -37765 7790
rect -37730 7755 -37720 7790
rect -37685 7755 -37675 7790
rect -37640 7755 -37630 7790
rect -37595 7755 -37585 7790
rect -37550 7755 -37540 7790
rect -37505 7755 -37495 7790
rect -37460 7755 -37450 7790
rect -37415 7755 -37405 7790
rect -37370 7755 -37360 7790
rect -37325 7755 -37315 7790
rect -37280 7755 -37270 7790
rect -37235 7755 -37225 7790
rect -37190 7755 -37170 7790
rect -38770 7745 -37170 7755
rect -38770 7710 -38755 7745
rect -38720 7710 -38710 7745
rect -38675 7710 -38665 7745
rect -38630 7710 -38620 7745
rect -38585 7710 -38575 7745
rect -38540 7710 -38530 7745
rect -38495 7710 -38485 7745
rect -38450 7710 -38440 7745
rect -38405 7710 -38395 7745
rect -38360 7710 -38350 7745
rect -38315 7710 -38305 7745
rect -38270 7710 -38260 7745
rect -38225 7710 -38215 7745
rect -38180 7710 -38170 7745
rect -38135 7710 -38125 7745
rect -38090 7710 -38080 7745
rect -38045 7710 -38035 7745
rect -38000 7710 -37990 7745
rect -37955 7710 -37945 7745
rect -37910 7710 -37900 7745
rect -37865 7710 -37855 7745
rect -37820 7710 -37810 7745
rect -37775 7710 -37765 7745
rect -37730 7710 -37720 7745
rect -37685 7710 -37675 7745
rect -37640 7710 -37630 7745
rect -37595 7710 -37585 7745
rect -37550 7710 -37540 7745
rect -37505 7710 -37495 7745
rect -37460 7710 -37450 7745
rect -37415 7710 -37405 7745
rect -37370 7710 -37360 7745
rect -37325 7710 -37315 7745
rect -37280 7710 -37270 7745
rect -37235 7710 -37225 7745
rect -37190 7710 -37170 7745
rect -38770 7700 -37170 7710
rect -38770 7665 -38755 7700
rect -38720 7665 -38710 7700
rect -38675 7665 -38665 7700
rect -38630 7665 -38620 7700
rect -38585 7665 -38575 7700
rect -38540 7665 -38530 7700
rect -38495 7665 -38485 7700
rect -38450 7665 -38440 7700
rect -38405 7665 -38395 7700
rect -38360 7665 -38350 7700
rect -38315 7665 -38305 7700
rect -38270 7665 -38260 7700
rect -38225 7665 -38215 7700
rect -38180 7665 -38170 7700
rect -38135 7665 -38125 7700
rect -38090 7665 -38080 7700
rect -38045 7665 -38035 7700
rect -38000 7665 -37990 7700
rect -37955 7665 -37945 7700
rect -37910 7665 -37900 7700
rect -37865 7665 -37855 7700
rect -37820 7665 -37810 7700
rect -37775 7665 -37765 7700
rect -37730 7665 -37720 7700
rect -37685 7665 -37675 7700
rect -37640 7665 -37630 7700
rect -37595 7665 -37585 7700
rect -37550 7665 -37540 7700
rect -37505 7665 -37495 7700
rect -37460 7665 -37450 7700
rect -37415 7665 -37405 7700
rect -37370 7665 -37360 7700
rect -37325 7665 -37315 7700
rect -37280 7665 -37270 7700
rect -37235 7665 -37225 7700
rect -37190 7665 -37170 7700
rect -38770 7655 -37170 7665
rect -38770 7620 -38755 7655
rect -38720 7620 -38710 7655
rect -38675 7620 -38665 7655
rect -38630 7620 -38620 7655
rect -38585 7620 -38575 7655
rect -38540 7620 -38530 7655
rect -38495 7620 -38485 7655
rect -38450 7620 -38440 7655
rect -38405 7620 -38395 7655
rect -38360 7620 -38350 7655
rect -38315 7620 -38305 7655
rect -38270 7620 -38260 7655
rect -38225 7620 -38215 7655
rect -38180 7620 -38170 7655
rect -38135 7620 -38125 7655
rect -38090 7620 -38080 7655
rect -38045 7620 -38035 7655
rect -38000 7620 -37990 7655
rect -37955 7620 -37945 7655
rect -37910 7620 -37900 7655
rect -37865 7620 -37855 7655
rect -37820 7620 -37810 7655
rect -37775 7620 -37765 7655
rect -37730 7620 -37720 7655
rect -37685 7620 -37675 7655
rect -37640 7620 -37630 7655
rect -37595 7620 -37585 7655
rect -37550 7620 -37540 7655
rect -37505 7620 -37495 7655
rect -37460 7620 -37450 7655
rect -37415 7620 -37405 7655
rect -37370 7620 -37360 7655
rect -37325 7620 -37315 7655
rect -37280 7620 -37270 7655
rect -37235 7620 -37225 7655
rect -37190 7620 -37170 7655
rect -38770 7610 -37170 7620
rect -38770 7575 -38755 7610
rect -38720 7575 -38710 7610
rect -38675 7575 -38665 7610
rect -38630 7575 -38620 7610
rect -38585 7575 -38575 7610
rect -38540 7575 -38530 7610
rect -38495 7575 -38485 7610
rect -38450 7575 -38440 7610
rect -38405 7575 -38395 7610
rect -38360 7575 -38350 7610
rect -38315 7575 -38305 7610
rect -38270 7575 -38260 7610
rect -38225 7575 -38215 7610
rect -38180 7575 -38170 7610
rect -38135 7575 -38125 7610
rect -38090 7575 -38080 7610
rect -38045 7575 -38035 7610
rect -38000 7575 -37990 7610
rect -37955 7575 -37945 7610
rect -37910 7575 -37900 7610
rect -37865 7575 -37855 7610
rect -37820 7575 -37810 7610
rect -37775 7575 -37765 7610
rect -37730 7575 -37720 7610
rect -37685 7575 -37675 7610
rect -37640 7575 -37630 7610
rect -37595 7575 -37585 7610
rect -37550 7575 -37540 7610
rect -37505 7575 -37495 7610
rect -37460 7575 -37450 7610
rect -37415 7575 -37405 7610
rect -37370 7575 -37360 7610
rect -37325 7575 -37315 7610
rect -37280 7575 -37270 7610
rect -37235 7575 -37225 7610
rect -37190 7575 -37170 7610
rect -38770 7565 -37170 7575
rect -38770 7530 -38755 7565
rect -38720 7530 -38710 7565
rect -38675 7530 -38665 7565
rect -38630 7530 -38620 7565
rect -38585 7530 -38575 7565
rect -38540 7530 -38530 7565
rect -38495 7530 -38485 7565
rect -38450 7530 -38440 7565
rect -38405 7530 -38395 7565
rect -38360 7530 -38350 7565
rect -38315 7530 -38305 7565
rect -38270 7530 -38260 7565
rect -38225 7530 -38215 7565
rect -38180 7530 -38170 7565
rect -38135 7530 -38125 7565
rect -38090 7530 -38080 7565
rect -38045 7530 -38035 7565
rect -38000 7530 -37990 7565
rect -37955 7530 -37945 7565
rect -37910 7530 -37900 7565
rect -37865 7530 -37855 7565
rect -37820 7530 -37810 7565
rect -37775 7530 -37765 7565
rect -37730 7530 -37720 7565
rect -37685 7530 -37675 7565
rect -37640 7530 -37630 7565
rect -37595 7530 -37585 7565
rect -37550 7530 -37540 7565
rect -37505 7530 -37495 7565
rect -37460 7530 -37450 7565
rect -37415 7530 -37405 7565
rect -37370 7530 -37360 7565
rect -37325 7530 -37315 7565
rect -37280 7530 -37270 7565
rect -37235 7530 -37225 7565
rect -37190 7530 -37170 7565
rect -38770 7520 -37170 7530
rect -38770 7485 -38755 7520
rect -38720 7485 -38710 7520
rect -38675 7485 -38665 7520
rect -38630 7485 -38620 7520
rect -38585 7485 -38575 7520
rect -38540 7485 -38530 7520
rect -38495 7485 -38485 7520
rect -38450 7485 -38440 7520
rect -38405 7485 -38395 7520
rect -38360 7485 -38350 7520
rect -38315 7485 -38305 7520
rect -38270 7485 -38260 7520
rect -38225 7485 -38215 7520
rect -38180 7485 -38170 7520
rect -38135 7485 -38125 7520
rect -38090 7485 -38080 7520
rect -38045 7485 -38035 7520
rect -38000 7485 -37990 7520
rect -37955 7485 -37945 7520
rect -37910 7485 -37900 7520
rect -37865 7485 -37855 7520
rect -37820 7485 -37810 7520
rect -37775 7485 -37765 7520
rect -37730 7485 -37720 7520
rect -37685 7485 -37675 7520
rect -37640 7485 -37630 7520
rect -37595 7485 -37585 7520
rect -37550 7485 -37540 7520
rect -37505 7485 -37495 7520
rect -37460 7485 -37450 7520
rect -37415 7485 -37405 7520
rect -37370 7485 -37360 7520
rect -37325 7485 -37315 7520
rect -37280 7485 -37270 7520
rect -37235 7485 -37225 7520
rect -37190 7485 -37170 7520
rect -38770 7475 -37170 7485
rect -38770 7440 -38755 7475
rect -38720 7440 -38710 7475
rect -38675 7440 -38665 7475
rect -38630 7440 -38620 7475
rect -38585 7440 -38575 7475
rect -38540 7440 -38530 7475
rect -38495 7440 -38485 7475
rect -38450 7440 -38440 7475
rect -38405 7440 -38395 7475
rect -38360 7440 -38350 7475
rect -38315 7440 -38305 7475
rect -38270 7440 -38260 7475
rect -38225 7440 -38215 7475
rect -38180 7440 -38170 7475
rect -38135 7440 -38125 7475
rect -38090 7440 -38080 7475
rect -38045 7440 -38035 7475
rect -38000 7440 -37990 7475
rect -37955 7440 -37945 7475
rect -37910 7440 -37900 7475
rect -37865 7440 -37855 7475
rect -37820 7440 -37810 7475
rect -37775 7440 -37765 7475
rect -37730 7440 -37720 7475
rect -37685 7440 -37675 7475
rect -37640 7440 -37630 7475
rect -37595 7440 -37585 7475
rect -37550 7440 -37540 7475
rect -37505 7440 -37495 7475
rect -37460 7440 -37450 7475
rect -37415 7440 -37405 7475
rect -37370 7440 -37360 7475
rect -37325 7440 -37315 7475
rect -37280 7440 -37270 7475
rect -37235 7440 -37225 7475
rect -37190 7440 -37170 7475
rect -38770 7430 -37170 7440
rect -38770 7395 -38755 7430
rect -38720 7395 -38710 7430
rect -38675 7395 -38665 7430
rect -38630 7395 -38620 7430
rect -38585 7395 -38575 7430
rect -38540 7395 -38530 7430
rect -38495 7395 -38485 7430
rect -38450 7395 -38440 7430
rect -38405 7395 -38395 7430
rect -38360 7395 -38350 7430
rect -38315 7395 -38305 7430
rect -38270 7395 -38260 7430
rect -38225 7395 -38215 7430
rect -38180 7395 -38170 7430
rect -38135 7395 -38125 7430
rect -38090 7395 -38080 7430
rect -38045 7395 -38035 7430
rect -38000 7395 -37990 7430
rect -37955 7395 -37945 7430
rect -37910 7395 -37900 7430
rect -37865 7395 -37855 7430
rect -37820 7395 -37810 7430
rect -37775 7395 -37765 7430
rect -37730 7395 -37720 7430
rect -37685 7395 -37675 7430
rect -37640 7395 -37630 7430
rect -37595 7395 -37585 7430
rect -37550 7395 -37540 7430
rect -37505 7395 -37495 7430
rect -37460 7395 -37450 7430
rect -37415 7395 -37405 7430
rect -37370 7395 -37360 7430
rect -37325 7395 -37315 7430
rect -37280 7395 -37270 7430
rect -37235 7395 -37225 7430
rect -37190 7395 -37170 7430
rect -38770 7385 -37170 7395
rect -38770 7350 -38755 7385
rect -38720 7350 -38710 7385
rect -38675 7350 -38665 7385
rect -38630 7350 -38620 7385
rect -38585 7350 -38575 7385
rect -38540 7350 -38530 7385
rect -38495 7350 -38485 7385
rect -38450 7350 -38440 7385
rect -38405 7350 -38395 7385
rect -38360 7350 -38350 7385
rect -38315 7350 -38305 7385
rect -38270 7350 -38260 7385
rect -38225 7350 -38215 7385
rect -38180 7350 -38170 7385
rect -38135 7350 -38125 7385
rect -38090 7350 -38080 7385
rect -38045 7350 -38035 7385
rect -38000 7350 -37990 7385
rect -37955 7350 -37945 7385
rect -37910 7350 -37900 7385
rect -37865 7350 -37855 7385
rect -37820 7350 -37810 7385
rect -37775 7350 -37765 7385
rect -37730 7350 -37720 7385
rect -37685 7350 -37675 7385
rect -37640 7350 -37630 7385
rect -37595 7350 -37585 7385
rect -37550 7350 -37540 7385
rect -37505 7350 -37495 7385
rect -37460 7350 -37450 7385
rect -37415 7350 -37405 7385
rect -37370 7350 -37360 7385
rect -37325 7350 -37315 7385
rect -37280 7350 -37270 7385
rect -37235 7350 -37225 7385
rect -37190 7350 -37170 7385
rect -38770 7340 -37170 7350
rect -38770 7305 -38755 7340
rect -38720 7305 -38710 7340
rect -38675 7305 -38665 7340
rect -38630 7305 -38620 7340
rect -38585 7305 -38575 7340
rect -38540 7305 -38530 7340
rect -38495 7305 -38485 7340
rect -38450 7305 -38440 7340
rect -38405 7305 -38395 7340
rect -38360 7305 -38350 7340
rect -38315 7305 -38305 7340
rect -38270 7305 -38260 7340
rect -38225 7305 -38215 7340
rect -38180 7305 -38170 7340
rect -38135 7305 -38125 7340
rect -38090 7305 -38080 7340
rect -38045 7305 -38035 7340
rect -38000 7305 -37990 7340
rect -37955 7305 -37945 7340
rect -37910 7305 -37900 7340
rect -37865 7305 -37855 7340
rect -37820 7305 -37810 7340
rect -37775 7305 -37765 7340
rect -37730 7305 -37720 7340
rect -37685 7305 -37675 7340
rect -37640 7305 -37630 7340
rect -37595 7305 -37585 7340
rect -37550 7305 -37540 7340
rect -37505 7305 -37495 7340
rect -37460 7305 -37450 7340
rect -37415 7305 -37405 7340
rect -37370 7305 -37360 7340
rect -37325 7305 -37315 7340
rect -37280 7305 -37270 7340
rect -37235 7305 -37225 7340
rect -37190 7305 -37170 7340
rect -38770 7295 -37170 7305
rect -38770 7260 -38755 7295
rect -38720 7260 -38710 7295
rect -38675 7260 -38665 7295
rect -38630 7260 -38620 7295
rect -38585 7260 -38575 7295
rect -38540 7260 -38530 7295
rect -38495 7260 -38485 7295
rect -38450 7260 -38440 7295
rect -38405 7260 -38395 7295
rect -38360 7260 -38350 7295
rect -38315 7260 -38305 7295
rect -38270 7260 -38260 7295
rect -38225 7260 -38215 7295
rect -38180 7260 -38170 7295
rect -38135 7260 -38125 7295
rect -38090 7260 -38080 7295
rect -38045 7260 -38035 7295
rect -38000 7260 -37990 7295
rect -37955 7260 -37945 7295
rect -37910 7260 -37900 7295
rect -37865 7260 -37855 7295
rect -37820 7260 -37810 7295
rect -37775 7260 -37765 7295
rect -37730 7260 -37720 7295
rect -37685 7260 -37675 7295
rect -37640 7260 -37630 7295
rect -37595 7260 -37585 7295
rect -37550 7260 -37540 7295
rect -37505 7260 -37495 7295
rect -37460 7260 -37450 7295
rect -37415 7260 -37405 7295
rect -37370 7260 -37360 7295
rect -37325 7260 -37315 7295
rect -37280 7260 -37270 7295
rect -37235 7260 -37225 7295
rect -37190 7260 -37170 7295
rect -38770 7250 -37170 7260
rect -38770 7215 -38755 7250
rect -38720 7215 -38710 7250
rect -38675 7215 -38665 7250
rect -38630 7215 -38620 7250
rect -38585 7215 -38575 7250
rect -38540 7215 -38530 7250
rect -38495 7215 -38485 7250
rect -38450 7215 -38440 7250
rect -38405 7215 -38395 7250
rect -38360 7215 -38350 7250
rect -38315 7215 -38305 7250
rect -38270 7215 -38260 7250
rect -38225 7215 -38215 7250
rect -38180 7215 -38170 7250
rect -38135 7215 -38125 7250
rect -38090 7215 -38080 7250
rect -38045 7215 -38035 7250
rect -38000 7215 -37990 7250
rect -37955 7215 -37945 7250
rect -37910 7215 -37900 7250
rect -37865 7215 -37855 7250
rect -37820 7215 -37810 7250
rect -37775 7215 -37765 7250
rect -37730 7215 -37720 7250
rect -37685 7215 -37675 7250
rect -37640 7215 -37630 7250
rect -37595 7215 -37585 7250
rect -37550 7215 -37540 7250
rect -37505 7215 -37495 7250
rect -37460 7215 -37450 7250
rect -37415 7215 -37405 7250
rect -37370 7215 -37360 7250
rect -37325 7215 -37315 7250
rect -37280 7215 -37270 7250
rect -37235 7215 -37225 7250
rect -37190 7215 -37170 7250
rect -38770 7205 -37170 7215
rect -38770 7170 -38755 7205
rect -38720 7170 -38710 7205
rect -38675 7170 -38665 7205
rect -38630 7170 -38620 7205
rect -38585 7170 -38575 7205
rect -38540 7170 -38530 7205
rect -38495 7170 -38485 7205
rect -38450 7170 -38440 7205
rect -38405 7170 -38395 7205
rect -38360 7170 -38350 7205
rect -38315 7170 -38305 7205
rect -38270 7170 -38260 7205
rect -38225 7170 -38215 7205
rect -38180 7170 -38170 7205
rect -38135 7170 -38125 7205
rect -38090 7170 -38080 7205
rect -38045 7170 -38035 7205
rect -38000 7170 -37990 7205
rect -37955 7170 -37945 7205
rect -37910 7170 -37900 7205
rect -37865 7170 -37855 7205
rect -37820 7170 -37810 7205
rect -37775 7170 -37765 7205
rect -37730 7170 -37720 7205
rect -37685 7170 -37675 7205
rect -37640 7170 -37630 7205
rect -37595 7170 -37585 7205
rect -37550 7170 -37540 7205
rect -37505 7170 -37495 7205
rect -37460 7170 -37450 7205
rect -37415 7170 -37405 7205
rect -37370 7170 -37360 7205
rect -37325 7170 -37315 7205
rect -37280 7170 -37270 7205
rect -37235 7170 -37225 7205
rect -37190 7170 -37170 7205
rect -38770 7160 -37170 7170
rect -38770 7125 -38755 7160
rect -38720 7125 -38710 7160
rect -38675 7125 -38665 7160
rect -38630 7125 -38620 7160
rect -38585 7125 -38575 7160
rect -38540 7125 -38530 7160
rect -38495 7125 -38485 7160
rect -38450 7125 -38440 7160
rect -38405 7125 -38395 7160
rect -38360 7125 -38350 7160
rect -38315 7125 -38305 7160
rect -38270 7125 -38260 7160
rect -38225 7125 -38215 7160
rect -38180 7125 -38170 7160
rect -38135 7125 -38125 7160
rect -38090 7125 -38080 7160
rect -38045 7125 -38035 7160
rect -38000 7125 -37990 7160
rect -37955 7125 -37945 7160
rect -37910 7125 -37900 7160
rect -37865 7125 -37855 7160
rect -37820 7125 -37810 7160
rect -37775 7125 -37765 7160
rect -37730 7125 -37720 7160
rect -37685 7125 -37675 7160
rect -37640 7125 -37630 7160
rect -37595 7125 -37585 7160
rect -37550 7125 -37540 7160
rect -37505 7125 -37495 7160
rect -37460 7125 -37450 7160
rect -37415 7125 -37405 7160
rect -37370 7125 -37360 7160
rect -37325 7125 -37315 7160
rect -37280 7125 -37270 7160
rect -37235 7125 -37225 7160
rect -37190 7125 -37170 7160
rect -38770 7115 -37170 7125
rect -38770 7080 -38755 7115
rect -38720 7080 -38710 7115
rect -38675 7080 -38665 7115
rect -38630 7080 -38620 7115
rect -38585 7080 -38575 7115
rect -38540 7080 -38530 7115
rect -38495 7080 -38485 7115
rect -38450 7080 -38440 7115
rect -38405 7080 -38395 7115
rect -38360 7080 -38350 7115
rect -38315 7080 -38305 7115
rect -38270 7080 -38260 7115
rect -38225 7080 -38215 7115
rect -38180 7080 -38170 7115
rect -38135 7080 -38125 7115
rect -38090 7080 -38080 7115
rect -38045 7080 -38035 7115
rect -38000 7080 -37990 7115
rect -37955 7080 -37945 7115
rect -37910 7080 -37900 7115
rect -37865 7080 -37855 7115
rect -37820 7080 -37810 7115
rect -37775 7080 -37765 7115
rect -37730 7080 -37720 7115
rect -37685 7080 -37675 7115
rect -37640 7080 -37630 7115
rect -37595 7080 -37585 7115
rect -37550 7080 -37540 7115
rect -37505 7080 -37495 7115
rect -37460 7080 -37450 7115
rect -37415 7080 -37405 7115
rect -37370 7080 -37360 7115
rect -37325 7080 -37315 7115
rect -37280 7080 -37270 7115
rect -37235 7080 -37225 7115
rect -37190 7080 -37170 7115
rect -38770 7070 -37170 7080
rect -38770 7035 -38755 7070
rect -38720 7035 -38710 7070
rect -38675 7035 -38665 7070
rect -38630 7035 -38620 7070
rect -38585 7035 -38575 7070
rect -38540 7035 -38530 7070
rect -38495 7035 -38485 7070
rect -38450 7035 -38440 7070
rect -38405 7035 -38395 7070
rect -38360 7035 -38350 7070
rect -38315 7035 -38305 7070
rect -38270 7035 -38260 7070
rect -38225 7035 -38215 7070
rect -38180 7035 -38170 7070
rect -38135 7035 -38125 7070
rect -38090 7035 -38080 7070
rect -38045 7035 -38035 7070
rect -38000 7035 -37990 7070
rect -37955 7035 -37945 7070
rect -37910 7035 -37900 7070
rect -37865 7035 -37855 7070
rect -37820 7035 -37810 7070
rect -37775 7035 -37765 7070
rect -37730 7035 -37720 7070
rect -37685 7035 -37675 7070
rect -37640 7035 -37630 7070
rect -37595 7035 -37585 7070
rect -37550 7035 -37540 7070
rect -37505 7035 -37495 7070
rect -37460 7035 -37450 7070
rect -37415 7035 -37405 7070
rect -37370 7035 -37360 7070
rect -37325 7035 -37315 7070
rect -37280 7035 -37270 7070
rect -37235 7035 -37225 7070
rect -37190 7035 -37170 7070
rect -38770 7025 -37170 7035
rect -38770 6990 -38755 7025
rect -38720 6990 -38710 7025
rect -38675 6990 -38665 7025
rect -38630 6990 -38620 7025
rect -38585 6990 -38575 7025
rect -38540 6990 -38530 7025
rect -38495 6990 -38485 7025
rect -38450 6990 -38440 7025
rect -38405 6990 -38395 7025
rect -38360 6990 -38350 7025
rect -38315 6990 -38305 7025
rect -38270 6990 -38260 7025
rect -38225 6990 -38215 7025
rect -38180 6990 -38170 7025
rect -38135 6990 -38125 7025
rect -38090 6990 -38080 7025
rect -38045 6990 -38035 7025
rect -38000 6990 -37990 7025
rect -37955 6990 -37945 7025
rect -37910 6990 -37900 7025
rect -37865 6990 -37855 7025
rect -37820 6990 -37810 7025
rect -37775 6990 -37765 7025
rect -37730 6990 -37720 7025
rect -37685 6990 -37675 7025
rect -37640 6990 -37630 7025
rect -37595 6990 -37585 7025
rect -37550 6990 -37540 7025
rect -37505 6990 -37495 7025
rect -37460 6990 -37450 7025
rect -37415 6990 -37405 7025
rect -37370 6990 -37360 7025
rect -37325 6990 -37315 7025
rect -37280 6990 -37270 7025
rect -37235 6990 -37225 7025
rect -37190 6990 -37170 7025
rect -38770 6980 -37170 6990
rect -38770 6945 -38755 6980
rect -38720 6945 -38710 6980
rect -38675 6945 -38665 6980
rect -38630 6945 -38620 6980
rect -38585 6945 -38575 6980
rect -38540 6945 -38530 6980
rect -38495 6945 -38485 6980
rect -38450 6945 -38440 6980
rect -38405 6945 -38395 6980
rect -38360 6945 -38350 6980
rect -38315 6945 -38305 6980
rect -38270 6945 -38260 6980
rect -38225 6945 -38215 6980
rect -38180 6945 -38170 6980
rect -38135 6945 -38125 6980
rect -38090 6945 -38080 6980
rect -38045 6945 -38035 6980
rect -38000 6945 -37990 6980
rect -37955 6945 -37945 6980
rect -37910 6945 -37900 6980
rect -37865 6945 -37855 6980
rect -37820 6945 -37810 6980
rect -37775 6945 -37765 6980
rect -37730 6945 -37720 6980
rect -37685 6945 -37675 6980
rect -37640 6945 -37630 6980
rect -37595 6945 -37585 6980
rect -37550 6945 -37540 6980
rect -37505 6945 -37495 6980
rect -37460 6945 -37450 6980
rect -37415 6945 -37405 6980
rect -37370 6945 -37360 6980
rect -37325 6945 -37315 6980
rect -37280 6945 -37270 6980
rect -37235 6945 -37225 6980
rect -37190 6945 -37170 6980
rect -38770 6935 -37170 6945
rect -38770 6900 -38755 6935
rect -38720 6900 -38710 6935
rect -38675 6900 -38665 6935
rect -38630 6900 -38620 6935
rect -38585 6900 -38575 6935
rect -38540 6900 -38530 6935
rect -38495 6900 -38485 6935
rect -38450 6900 -38440 6935
rect -38405 6900 -38395 6935
rect -38360 6900 -38350 6935
rect -38315 6900 -38305 6935
rect -38270 6900 -38260 6935
rect -38225 6900 -38215 6935
rect -38180 6900 -38170 6935
rect -38135 6900 -38125 6935
rect -38090 6900 -38080 6935
rect -38045 6900 -38035 6935
rect -38000 6900 -37990 6935
rect -37955 6900 -37945 6935
rect -37910 6900 -37900 6935
rect -37865 6900 -37855 6935
rect -37820 6900 -37810 6935
rect -37775 6900 -37765 6935
rect -37730 6900 -37720 6935
rect -37685 6900 -37675 6935
rect -37640 6900 -37630 6935
rect -37595 6900 -37585 6935
rect -37550 6900 -37540 6935
rect -37505 6900 -37495 6935
rect -37460 6900 -37450 6935
rect -37415 6900 -37405 6935
rect -37370 6900 -37360 6935
rect -37325 6900 -37315 6935
rect -37280 6900 -37270 6935
rect -37235 6900 -37225 6935
rect -37190 6900 -37170 6935
rect -38770 6890 -37170 6900
rect -38770 6855 -38755 6890
rect -38720 6855 -38710 6890
rect -38675 6855 -38665 6890
rect -38630 6855 -38620 6890
rect -38585 6855 -38575 6890
rect -38540 6855 -38530 6890
rect -38495 6855 -38485 6890
rect -38450 6855 -38440 6890
rect -38405 6855 -38395 6890
rect -38360 6855 -38350 6890
rect -38315 6855 -38305 6890
rect -38270 6855 -38260 6890
rect -38225 6855 -38215 6890
rect -38180 6855 -38170 6890
rect -38135 6855 -38125 6890
rect -38090 6855 -38080 6890
rect -38045 6855 -38035 6890
rect -38000 6855 -37990 6890
rect -37955 6855 -37945 6890
rect -37910 6855 -37900 6890
rect -37865 6855 -37855 6890
rect -37820 6855 -37810 6890
rect -37775 6855 -37765 6890
rect -37730 6855 -37720 6890
rect -37685 6855 -37675 6890
rect -37640 6855 -37630 6890
rect -37595 6855 -37585 6890
rect -37550 6855 -37540 6890
rect -37505 6855 -37495 6890
rect -37460 6855 -37450 6890
rect -37415 6855 -37405 6890
rect -37370 6855 -37360 6890
rect -37325 6855 -37315 6890
rect -37280 6855 -37270 6890
rect -37235 6855 -37225 6890
rect -37190 6855 -37170 6890
rect -38770 6845 -37170 6855
rect -38770 6810 -38755 6845
rect -38720 6810 -38710 6845
rect -38675 6810 -38665 6845
rect -38630 6810 -38620 6845
rect -38585 6810 -38575 6845
rect -38540 6810 -38530 6845
rect -38495 6810 -38485 6845
rect -38450 6810 -38440 6845
rect -38405 6810 -38395 6845
rect -38360 6810 -38350 6845
rect -38315 6810 -38305 6845
rect -38270 6810 -38260 6845
rect -38225 6810 -38215 6845
rect -38180 6810 -38170 6845
rect -38135 6810 -38125 6845
rect -38090 6810 -38080 6845
rect -38045 6810 -38035 6845
rect -38000 6810 -37990 6845
rect -37955 6810 -37945 6845
rect -37910 6810 -37900 6845
rect -37865 6810 -37855 6845
rect -37820 6810 -37810 6845
rect -37775 6810 -37765 6845
rect -37730 6810 -37720 6845
rect -37685 6810 -37675 6845
rect -37640 6810 -37630 6845
rect -37595 6810 -37585 6845
rect -37550 6810 -37540 6845
rect -37505 6810 -37495 6845
rect -37460 6810 -37450 6845
rect -37415 6810 -37405 6845
rect -37370 6810 -37360 6845
rect -37325 6810 -37315 6845
rect -37280 6810 -37270 6845
rect -37235 6810 -37225 6845
rect -37190 6810 -37170 6845
rect -38770 6800 -37170 6810
rect -38770 6765 -38755 6800
rect -38720 6765 -38710 6800
rect -38675 6765 -38665 6800
rect -38630 6765 -38620 6800
rect -38585 6765 -38575 6800
rect -38540 6765 -38530 6800
rect -38495 6765 -38485 6800
rect -38450 6765 -38440 6800
rect -38405 6765 -38395 6800
rect -38360 6765 -38350 6800
rect -38315 6765 -38305 6800
rect -38270 6765 -38260 6800
rect -38225 6765 -38215 6800
rect -38180 6765 -38170 6800
rect -38135 6765 -38125 6800
rect -38090 6765 -38080 6800
rect -38045 6765 -38035 6800
rect -38000 6765 -37990 6800
rect -37955 6765 -37945 6800
rect -37910 6765 -37900 6800
rect -37865 6765 -37855 6800
rect -37820 6765 -37810 6800
rect -37775 6765 -37765 6800
rect -37730 6765 -37720 6800
rect -37685 6765 -37675 6800
rect -37640 6765 -37630 6800
rect -37595 6765 -37585 6800
rect -37550 6765 -37540 6800
rect -37505 6765 -37495 6800
rect -37460 6765 -37450 6800
rect -37415 6765 -37405 6800
rect -37370 6765 -37360 6800
rect -37325 6765 -37315 6800
rect -37280 6765 -37270 6800
rect -37235 6765 -37225 6800
rect -37190 6765 -37170 6800
rect -38770 6755 -37170 6765
rect -38770 6720 -38755 6755
rect -38720 6720 -38710 6755
rect -38675 6720 -38665 6755
rect -38630 6720 -38620 6755
rect -38585 6720 -38575 6755
rect -38540 6720 -38530 6755
rect -38495 6720 -38485 6755
rect -38450 6720 -38440 6755
rect -38405 6720 -38395 6755
rect -38360 6720 -38350 6755
rect -38315 6720 -38305 6755
rect -38270 6720 -38260 6755
rect -38225 6720 -38215 6755
rect -38180 6720 -38170 6755
rect -38135 6720 -38125 6755
rect -38090 6720 -38080 6755
rect -38045 6720 -38035 6755
rect -38000 6720 -37990 6755
rect -37955 6720 -37945 6755
rect -37910 6720 -37900 6755
rect -37865 6720 -37855 6755
rect -37820 6720 -37810 6755
rect -37775 6720 -37765 6755
rect -37730 6720 -37720 6755
rect -37685 6720 -37675 6755
rect -37640 6720 -37630 6755
rect -37595 6720 -37585 6755
rect -37550 6720 -37540 6755
rect -37505 6720 -37495 6755
rect -37460 6720 -37450 6755
rect -37415 6720 -37405 6755
rect -37370 6720 -37360 6755
rect -37325 6720 -37315 6755
rect -37280 6720 -37270 6755
rect -37235 6720 -37225 6755
rect -37190 6720 -37170 6755
rect -38770 6710 -37170 6720
rect -38770 6675 -38755 6710
rect -38720 6675 -38710 6710
rect -38675 6675 -38665 6710
rect -38630 6675 -38620 6710
rect -38585 6675 -38575 6710
rect -38540 6675 -38530 6710
rect -38495 6675 -38485 6710
rect -38450 6675 -38440 6710
rect -38405 6675 -38395 6710
rect -38360 6675 -38350 6710
rect -38315 6675 -38305 6710
rect -38270 6675 -38260 6710
rect -38225 6675 -38215 6710
rect -38180 6675 -38170 6710
rect -38135 6675 -38125 6710
rect -38090 6675 -38080 6710
rect -38045 6675 -38035 6710
rect -38000 6675 -37990 6710
rect -37955 6675 -37945 6710
rect -37910 6675 -37900 6710
rect -37865 6675 -37855 6710
rect -37820 6675 -37810 6710
rect -37775 6675 -37765 6710
rect -37730 6675 -37720 6710
rect -37685 6675 -37675 6710
rect -37640 6675 -37630 6710
rect -37595 6675 -37585 6710
rect -37550 6675 -37540 6710
rect -37505 6675 -37495 6710
rect -37460 6675 -37450 6710
rect -37415 6675 -37405 6710
rect -37370 6675 -37360 6710
rect -37325 6675 -37315 6710
rect -37280 6675 -37270 6710
rect -37235 6675 -37225 6710
rect -37190 6675 -37170 6710
rect -38770 6665 -37170 6675
rect -38770 6630 -38755 6665
rect -38720 6630 -38710 6665
rect -38675 6630 -38665 6665
rect -38630 6630 -38620 6665
rect -38585 6630 -38575 6665
rect -38540 6630 -38530 6665
rect -38495 6630 -38485 6665
rect -38450 6630 -38440 6665
rect -38405 6630 -38395 6665
rect -38360 6630 -38350 6665
rect -38315 6630 -38305 6665
rect -38270 6630 -38260 6665
rect -38225 6630 -38215 6665
rect -38180 6630 -38170 6665
rect -38135 6630 -38125 6665
rect -38090 6630 -38080 6665
rect -38045 6630 -38035 6665
rect -38000 6630 -37990 6665
rect -37955 6630 -37945 6665
rect -37910 6630 -37900 6665
rect -37865 6630 -37855 6665
rect -37820 6630 -37810 6665
rect -37775 6630 -37765 6665
rect -37730 6630 -37720 6665
rect -37685 6630 -37675 6665
rect -37640 6630 -37630 6665
rect -37595 6630 -37585 6665
rect -37550 6630 -37540 6665
rect -37505 6630 -37495 6665
rect -37460 6630 -37450 6665
rect -37415 6630 -37405 6665
rect -37370 6630 -37360 6665
rect -37325 6630 -37315 6665
rect -37280 6630 -37270 6665
rect -37235 6630 -37225 6665
rect -37190 6630 -37170 6665
rect -38770 6620 -37170 6630
rect -38770 6585 -38755 6620
rect -38720 6585 -38710 6620
rect -38675 6585 -38665 6620
rect -38630 6585 -38620 6620
rect -38585 6585 -38575 6620
rect -38540 6585 -38530 6620
rect -38495 6585 -38485 6620
rect -38450 6585 -38440 6620
rect -38405 6585 -38395 6620
rect -38360 6585 -38350 6620
rect -38315 6585 -38305 6620
rect -38270 6585 -38260 6620
rect -38225 6585 -38215 6620
rect -38180 6585 -38170 6620
rect -38135 6585 -38125 6620
rect -38090 6585 -38080 6620
rect -38045 6585 -38035 6620
rect -38000 6585 -37990 6620
rect -37955 6585 -37945 6620
rect -37910 6585 -37900 6620
rect -37865 6585 -37855 6620
rect -37820 6585 -37810 6620
rect -37775 6585 -37765 6620
rect -37730 6585 -37720 6620
rect -37685 6585 -37675 6620
rect -37640 6585 -37630 6620
rect -37595 6585 -37585 6620
rect -37550 6585 -37540 6620
rect -37505 6585 -37495 6620
rect -37460 6585 -37450 6620
rect -37415 6585 -37405 6620
rect -37370 6585 -37360 6620
rect -37325 6585 -37315 6620
rect -37280 6585 -37270 6620
rect -37235 6585 -37225 6620
rect -37190 6585 -37170 6620
rect -38770 6575 -37170 6585
rect -38770 6540 -38755 6575
rect -38720 6540 -38710 6575
rect -38675 6540 -38665 6575
rect -38630 6540 -38620 6575
rect -38585 6540 -38575 6575
rect -38540 6540 -38530 6575
rect -38495 6540 -38485 6575
rect -38450 6540 -38440 6575
rect -38405 6540 -38395 6575
rect -38360 6540 -38350 6575
rect -38315 6540 -38305 6575
rect -38270 6540 -38260 6575
rect -38225 6540 -38215 6575
rect -38180 6540 -38170 6575
rect -38135 6540 -38125 6575
rect -38090 6540 -38080 6575
rect -38045 6540 -38035 6575
rect -38000 6540 -37990 6575
rect -37955 6540 -37945 6575
rect -37910 6540 -37900 6575
rect -37865 6540 -37855 6575
rect -37820 6540 -37810 6575
rect -37775 6540 -37765 6575
rect -37730 6540 -37720 6575
rect -37685 6540 -37675 6575
rect -37640 6540 -37630 6575
rect -37595 6540 -37585 6575
rect -37550 6540 -37540 6575
rect -37505 6540 -37495 6575
rect -37460 6540 -37450 6575
rect -37415 6540 -37405 6575
rect -37370 6540 -37360 6575
rect -37325 6540 -37315 6575
rect -37280 6540 -37270 6575
rect -37235 6540 -37225 6575
rect -37190 6540 -37170 6575
rect -38770 6530 -37170 6540
rect -38770 6495 -38755 6530
rect -38720 6495 -38710 6530
rect -38675 6495 -38665 6530
rect -38630 6495 -38620 6530
rect -38585 6495 -38575 6530
rect -38540 6495 -38530 6530
rect -38495 6495 -38485 6530
rect -38450 6495 -38440 6530
rect -38405 6495 -38395 6530
rect -38360 6495 -38350 6530
rect -38315 6495 -38305 6530
rect -38270 6495 -38260 6530
rect -38225 6495 -38215 6530
rect -38180 6495 -38170 6530
rect -38135 6495 -38125 6530
rect -38090 6495 -38080 6530
rect -38045 6495 -38035 6530
rect -38000 6495 -37990 6530
rect -37955 6495 -37945 6530
rect -37910 6495 -37900 6530
rect -37865 6495 -37855 6530
rect -37820 6495 -37810 6530
rect -37775 6495 -37765 6530
rect -37730 6495 -37720 6530
rect -37685 6495 -37675 6530
rect -37640 6495 -37630 6530
rect -37595 6495 -37585 6530
rect -37550 6495 -37540 6530
rect -37505 6495 -37495 6530
rect -37460 6495 -37450 6530
rect -37415 6495 -37405 6530
rect -37370 6495 -37360 6530
rect -37325 6495 -37315 6530
rect -37280 6495 -37270 6530
rect -37235 6495 -37225 6530
rect -37190 6495 -37170 6530
rect -38770 6485 -37170 6495
rect -38770 6450 -38755 6485
rect -38720 6450 -38710 6485
rect -38675 6450 -38665 6485
rect -38630 6450 -38620 6485
rect -38585 6450 -38575 6485
rect -38540 6450 -38530 6485
rect -38495 6450 -38485 6485
rect -38450 6450 -38440 6485
rect -38405 6450 -38395 6485
rect -38360 6450 -38350 6485
rect -38315 6450 -38305 6485
rect -38270 6450 -38260 6485
rect -38225 6450 -38215 6485
rect -38180 6450 -38170 6485
rect -38135 6450 -38125 6485
rect -38090 6450 -38080 6485
rect -38045 6450 -38035 6485
rect -38000 6450 -37990 6485
rect -37955 6450 -37945 6485
rect -37910 6450 -37900 6485
rect -37865 6450 -37855 6485
rect -37820 6450 -37810 6485
rect -37775 6450 -37765 6485
rect -37730 6450 -37720 6485
rect -37685 6450 -37675 6485
rect -37640 6450 -37630 6485
rect -37595 6450 -37585 6485
rect -37550 6450 -37540 6485
rect -37505 6450 -37495 6485
rect -37460 6450 -37450 6485
rect -37415 6450 -37405 6485
rect -37370 6450 -37360 6485
rect -37325 6450 -37315 6485
rect -37280 6450 -37270 6485
rect -37235 6450 -37225 6485
rect -37190 6450 -37170 6485
rect -38770 5940 -37170 6450
rect 3165 7960 3280 7980
rect 3165 7920 3175 7960
rect 3215 7920 3235 7960
rect 3275 7920 3280 7960
rect 3165 7890 3280 7920
rect 3165 7850 3175 7890
rect 3215 7850 3235 7890
rect 3275 7850 3280 7890
rect 3165 7820 3280 7850
rect 3165 7780 3175 7820
rect 3215 7780 3235 7820
rect 3275 7780 3280 7820
rect 3165 7750 3280 7780
rect 3165 7710 3175 7750
rect 3215 7710 3235 7750
rect 3275 7710 3280 7750
rect 3165 7685 3280 7710
rect 3165 7645 3175 7685
rect 3215 7645 3235 7685
rect 3275 7645 3280 7685
rect 3165 7625 3280 7645
rect 3165 7585 3175 7625
rect 3215 7585 3235 7625
rect 3275 7585 3280 7625
rect 3165 7560 3280 7585
rect 3165 7520 3175 7560
rect 3215 7520 3235 7560
rect 3275 7520 3280 7560
rect 3165 7490 3280 7520
rect 3165 7450 3175 7490
rect 3215 7450 3235 7490
rect 3275 7450 3280 7490
rect 3165 7420 3280 7450
rect 3165 7380 3175 7420
rect 3215 7380 3235 7420
rect 3275 7380 3280 7420
rect 3165 7350 3280 7380
rect 3165 7310 3175 7350
rect 3215 7310 3235 7350
rect 3275 7310 3280 7350
rect 3165 7285 3280 7310
rect 3165 7245 3175 7285
rect 3215 7245 3235 7285
rect 3275 7245 3280 7285
rect 3165 7225 3280 7245
rect 3165 7185 3175 7225
rect 3215 7185 3235 7225
rect 3275 7185 3280 7225
rect 3165 7160 3280 7185
rect 3165 7120 3175 7160
rect 3215 7120 3235 7160
rect 3275 7120 3280 7160
rect 3165 7090 3280 7120
rect 3165 7050 3175 7090
rect 3215 7050 3235 7090
rect 3275 7050 3280 7090
rect 3165 7020 3280 7050
rect 3165 6980 3175 7020
rect 3215 6980 3235 7020
rect 3275 6980 3280 7020
rect 3165 6950 3280 6980
rect 3165 6910 3175 6950
rect 3215 6910 3235 6950
rect 3275 6910 3280 6950
rect 3165 6885 3280 6910
rect 3165 6845 3175 6885
rect 3215 6845 3235 6885
rect 3275 6845 3280 6885
rect 3165 6825 3280 6845
rect 3165 6785 3175 6825
rect 3215 6785 3235 6825
rect 3275 6785 3280 6825
rect 3165 6760 3280 6785
rect 3165 6720 3175 6760
rect 3215 6720 3235 6760
rect 3275 6720 3280 6760
rect 3165 6690 3280 6720
rect 3165 6650 3175 6690
rect 3215 6650 3235 6690
rect 3275 6650 3280 6690
rect 3165 6620 3280 6650
rect 3165 6580 3175 6620
rect 3215 6580 3235 6620
rect 3275 6580 3280 6620
rect 3165 6550 3280 6580
rect 3165 6510 3175 6550
rect 3215 6510 3235 6550
rect 3275 6510 3280 6550
rect 3165 6485 3280 6510
rect 3165 6445 3175 6485
rect 3215 6445 3235 6485
rect 3275 6445 3280 6485
rect 3165 6435 3280 6445
rect 3340 7960 3390 7980
rect 3340 7920 3345 7960
rect 3385 7920 3390 7960
rect 3340 7890 3390 7920
rect 3340 7850 3345 7890
rect 3385 7850 3390 7890
rect 3340 7820 3390 7850
rect 3340 7780 3345 7820
rect 3385 7780 3390 7820
rect 3340 7750 3390 7780
rect 3340 7710 3345 7750
rect 3385 7710 3390 7750
rect 3340 7685 3390 7710
rect 3340 7645 3345 7685
rect 3385 7645 3390 7685
rect 3340 7625 3390 7645
rect 3340 7585 3345 7625
rect 3385 7585 3390 7625
rect 3340 7560 3390 7585
rect 3340 7520 3345 7560
rect 3385 7520 3390 7560
rect 3340 7490 3390 7520
rect 3340 7450 3345 7490
rect 3385 7450 3390 7490
rect 3340 7420 3390 7450
rect 3340 7380 3345 7420
rect 3385 7380 3390 7420
rect 3340 7350 3390 7380
rect 3340 7310 3345 7350
rect 3385 7310 3390 7350
rect 3340 7285 3390 7310
rect 3340 7245 3345 7285
rect 3385 7245 3390 7285
rect 3340 7225 3390 7245
rect 3340 7185 3345 7225
rect 3385 7185 3390 7225
rect 3340 7160 3390 7185
rect 3340 7120 3345 7160
rect 3385 7120 3390 7160
rect 3340 7090 3390 7120
rect 3340 7050 3345 7090
rect 3385 7050 3390 7090
rect 3340 7020 3390 7050
rect 3340 6980 3345 7020
rect 3385 6980 3390 7020
rect 3340 6950 3390 6980
rect 3340 6910 3345 6950
rect 3385 6910 3390 6950
rect 3340 6885 3390 6910
rect 3340 6845 3345 6885
rect 3385 6845 3390 6885
rect 3340 6825 3390 6845
rect 3340 6785 3345 6825
rect 3385 6785 3390 6825
rect 3340 6760 3390 6785
rect 3340 6720 3345 6760
rect 3385 6720 3390 6760
rect 3340 6690 3390 6720
rect 3340 6650 3345 6690
rect 3385 6650 3390 6690
rect 3340 6620 3390 6650
rect 3340 6580 3345 6620
rect 3385 6580 3390 6620
rect 3340 6550 3390 6580
rect 3340 6510 3345 6550
rect 3385 6510 3390 6550
rect 3340 6485 3390 6510
rect 3340 6445 3345 6485
rect 3385 6445 3390 6485
rect 3340 6435 3390 6445
rect 31290 7950 31305 7985
rect 31340 7950 31350 7985
rect 31385 7950 31395 7985
rect 31430 7950 31440 7985
rect 31475 7950 31485 7985
rect 31520 7950 31530 7985
rect 31565 7950 31575 7985
rect 31610 7950 31620 7985
rect 31655 7950 31665 7985
rect 31700 7950 31710 7985
rect 31745 7950 31755 7985
rect 31790 7950 31800 7985
rect 31835 7950 31845 7985
rect 31880 7950 31890 7985
rect 31925 7950 31935 7985
rect 31970 7950 31980 7985
rect 32015 7950 32025 7985
rect 32060 7950 32070 7985
rect 32105 7950 32115 7985
rect 32150 7950 32160 7985
rect 32195 7950 32205 7985
rect 32240 7950 32250 7985
rect 32285 7950 32295 7985
rect 32330 7950 32340 7985
rect 32375 7950 32385 7985
rect 32420 7950 32430 7985
rect 32465 7950 32475 7985
rect 32510 7950 32520 7985
rect 32555 7950 32565 7985
rect 32600 7950 32610 7985
rect 32645 7950 32655 7985
rect 32690 7950 32700 7985
rect 32735 7950 32745 7985
rect 32780 7950 32790 7985
rect 32825 7950 32835 7985
rect 32870 7950 32890 7985
rect 31290 7940 32890 7950
rect 31290 7905 31305 7940
rect 31340 7905 31350 7940
rect 31385 7905 31395 7940
rect 31430 7905 31440 7940
rect 31475 7905 31485 7940
rect 31520 7905 31530 7940
rect 31565 7905 31575 7940
rect 31610 7905 31620 7940
rect 31655 7905 31665 7940
rect 31700 7905 31710 7940
rect 31745 7905 31755 7940
rect 31790 7905 31800 7940
rect 31835 7905 31845 7940
rect 31880 7905 31890 7940
rect 31925 7905 31935 7940
rect 31970 7905 31980 7940
rect 32015 7905 32025 7940
rect 32060 7905 32070 7940
rect 32105 7905 32115 7940
rect 32150 7905 32160 7940
rect 32195 7905 32205 7940
rect 32240 7905 32250 7940
rect 32285 7905 32295 7940
rect 32330 7905 32340 7940
rect 32375 7905 32385 7940
rect 32420 7905 32430 7940
rect 32465 7905 32475 7940
rect 32510 7905 32520 7940
rect 32555 7905 32565 7940
rect 32600 7905 32610 7940
rect 32645 7905 32655 7940
rect 32690 7905 32700 7940
rect 32735 7905 32745 7940
rect 32780 7905 32790 7940
rect 32825 7905 32835 7940
rect 32870 7905 32890 7940
rect 31290 7895 32890 7905
rect 31290 7860 31305 7895
rect 31340 7860 31350 7895
rect 31385 7860 31395 7895
rect 31430 7860 31440 7895
rect 31475 7860 31485 7895
rect 31520 7860 31530 7895
rect 31565 7860 31575 7895
rect 31610 7860 31620 7895
rect 31655 7860 31665 7895
rect 31700 7860 31710 7895
rect 31745 7860 31755 7895
rect 31790 7860 31800 7895
rect 31835 7860 31845 7895
rect 31880 7860 31890 7895
rect 31925 7860 31935 7895
rect 31970 7860 31980 7895
rect 32015 7860 32025 7895
rect 32060 7860 32070 7895
rect 32105 7860 32115 7895
rect 32150 7860 32160 7895
rect 32195 7860 32205 7895
rect 32240 7860 32250 7895
rect 32285 7860 32295 7895
rect 32330 7860 32340 7895
rect 32375 7860 32385 7895
rect 32420 7860 32430 7895
rect 32465 7860 32475 7895
rect 32510 7860 32520 7895
rect 32555 7860 32565 7895
rect 32600 7860 32610 7895
rect 32645 7860 32655 7895
rect 32690 7860 32700 7895
rect 32735 7860 32745 7895
rect 32780 7860 32790 7895
rect 32825 7860 32835 7895
rect 32870 7860 32890 7895
rect 31290 7850 32890 7860
rect 31290 7815 31305 7850
rect 31340 7815 31350 7850
rect 31385 7815 31395 7850
rect 31430 7815 31440 7850
rect 31475 7815 31485 7850
rect 31520 7815 31530 7850
rect 31565 7815 31575 7850
rect 31610 7815 31620 7850
rect 31655 7815 31665 7850
rect 31700 7815 31710 7850
rect 31745 7815 31755 7850
rect 31790 7815 31800 7850
rect 31835 7815 31845 7850
rect 31880 7815 31890 7850
rect 31925 7815 31935 7850
rect 31970 7815 31980 7850
rect 32015 7815 32025 7850
rect 32060 7815 32070 7850
rect 32105 7815 32115 7850
rect 32150 7815 32160 7850
rect 32195 7815 32205 7850
rect 32240 7815 32250 7850
rect 32285 7815 32295 7850
rect 32330 7815 32340 7850
rect 32375 7815 32385 7850
rect 32420 7815 32430 7850
rect 32465 7815 32475 7850
rect 32510 7815 32520 7850
rect 32555 7815 32565 7850
rect 32600 7815 32610 7850
rect 32645 7815 32655 7850
rect 32690 7815 32700 7850
rect 32735 7815 32745 7850
rect 32780 7815 32790 7850
rect 32825 7815 32835 7850
rect 32870 7815 32890 7850
rect 31290 7805 32890 7815
rect 31290 7770 31305 7805
rect 31340 7770 31350 7805
rect 31385 7770 31395 7805
rect 31430 7770 31440 7805
rect 31475 7770 31485 7805
rect 31520 7770 31530 7805
rect 31565 7770 31575 7805
rect 31610 7770 31620 7805
rect 31655 7770 31665 7805
rect 31700 7770 31710 7805
rect 31745 7770 31755 7805
rect 31790 7770 31800 7805
rect 31835 7770 31845 7805
rect 31880 7770 31890 7805
rect 31925 7770 31935 7805
rect 31970 7770 31980 7805
rect 32015 7770 32025 7805
rect 32060 7770 32070 7805
rect 32105 7770 32115 7805
rect 32150 7770 32160 7805
rect 32195 7770 32205 7805
rect 32240 7770 32250 7805
rect 32285 7770 32295 7805
rect 32330 7770 32340 7805
rect 32375 7770 32385 7805
rect 32420 7770 32430 7805
rect 32465 7770 32475 7805
rect 32510 7770 32520 7805
rect 32555 7770 32565 7805
rect 32600 7770 32610 7805
rect 32645 7770 32655 7805
rect 32690 7770 32700 7805
rect 32735 7770 32745 7805
rect 32780 7770 32790 7805
rect 32825 7770 32835 7805
rect 32870 7770 32890 7805
rect 31290 7760 32890 7770
rect 31290 7725 31305 7760
rect 31340 7725 31350 7760
rect 31385 7725 31395 7760
rect 31430 7725 31440 7760
rect 31475 7725 31485 7760
rect 31520 7725 31530 7760
rect 31565 7725 31575 7760
rect 31610 7725 31620 7760
rect 31655 7725 31665 7760
rect 31700 7725 31710 7760
rect 31745 7725 31755 7760
rect 31790 7725 31800 7760
rect 31835 7725 31845 7760
rect 31880 7725 31890 7760
rect 31925 7725 31935 7760
rect 31970 7725 31980 7760
rect 32015 7725 32025 7760
rect 32060 7725 32070 7760
rect 32105 7725 32115 7760
rect 32150 7725 32160 7760
rect 32195 7725 32205 7760
rect 32240 7725 32250 7760
rect 32285 7725 32295 7760
rect 32330 7725 32340 7760
rect 32375 7725 32385 7760
rect 32420 7725 32430 7760
rect 32465 7725 32475 7760
rect 32510 7725 32520 7760
rect 32555 7725 32565 7760
rect 32600 7725 32610 7760
rect 32645 7725 32655 7760
rect 32690 7725 32700 7760
rect 32735 7725 32745 7760
rect 32780 7725 32790 7760
rect 32825 7725 32835 7760
rect 32870 7725 32890 7760
rect 31290 7715 32890 7725
rect 31290 7680 31305 7715
rect 31340 7680 31350 7715
rect 31385 7680 31395 7715
rect 31430 7680 31440 7715
rect 31475 7680 31485 7715
rect 31520 7680 31530 7715
rect 31565 7680 31575 7715
rect 31610 7680 31620 7715
rect 31655 7680 31665 7715
rect 31700 7680 31710 7715
rect 31745 7680 31755 7715
rect 31790 7680 31800 7715
rect 31835 7680 31845 7715
rect 31880 7680 31890 7715
rect 31925 7680 31935 7715
rect 31970 7680 31980 7715
rect 32015 7680 32025 7715
rect 32060 7680 32070 7715
rect 32105 7680 32115 7715
rect 32150 7680 32160 7715
rect 32195 7680 32205 7715
rect 32240 7680 32250 7715
rect 32285 7680 32295 7715
rect 32330 7680 32340 7715
rect 32375 7680 32385 7715
rect 32420 7680 32430 7715
rect 32465 7680 32475 7715
rect 32510 7680 32520 7715
rect 32555 7680 32565 7715
rect 32600 7680 32610 7715
rect 32645 7680 32655 7715
rect 32690 7680 32700 7715
rect 32735 7680 32745 7715
rect 32780 7680 32790 7715
rect 32825 7680 32835 7715
rect 32870 7680 32890 7715
rect 31290 7670 32890 7680
rect 31290 7635 31305 7670
rect 31340 7635 31350 7670
rect 31385 7635 31395 7670
rect 31430 7635 31440 7670
rect 31475 7635 31485 7670
rect 31520 7635 31530 7670
rect 31565 7635 31575 7670
rect 31610 7635 31620 7670
rect 31655 7635 31665 7670
rect 31700 7635 31710 7670
rect 31745 7635 31755 7670
rect 31790 7635 31800 7670
rect 31835 7635 31845 7670
rect 31880 7635 31890 7670
rect 31925 7635 31935 7670
rect 31970 7635 31980 7670
rect 32015 7635 32025 7670
rect 32060 7635 32070 7670
rect 32105 7635 32115 7670
rect 32150 7635 32160 7670
rect 32195 7635 32205 7670
rect 32240 7635 32250 7670
rect 32285 7635 32295 7670
rect 32330 7635 32340 7670
rect 32375 7635 32385 7670
rect 32420 7635 32430 7670
rect 32465 7635 32475 7670
rect 32510 7635 32520 7670
rect 32555 7635 32565 7670
rect 32600 7635 32610 7670
rect 32645 7635 32655 7670
rect 32690 7635 32700 7670
rect 32735 7635 32745 7670
rect 32780 7635 32790 7670
rect 32825 7635 32835 7670
rect 32870 7635 32890 7670
rect 31290 7625 32890 7635
rect 31290 7590 31305 7625
rect 31340 7590 31350 7625
rect 31385 7590 31395 7625
rect 31430 7590 31440 7625
rect 31475 7590 31485 7625
rect 31520 7590 31530 7625
rect 31565 7590 31575 7625
rect 31610 7590 31620 7625
rect 31655 7590 31665 7625
rect 31700 7590 31710 7625
rect 31745 7590 31755 7625
rect 31790 7590 31800 7625
rect 31835 7590 31845 7625
rect 31880 7590 31890 7625
rect 31925 7590 31935 7625
rect 31970 7590 31980 7625
rect 32015 7590 32025 7625
rect 32060 7590 32070 7625
rect 32105 7590 32115 7625
rect 32150 7590 32160 7625
rect 32195 7590 32205 7625
rect 32240 7590 32250 7625
rect 32285 7590 32295 7625
rect 32330 7590 32340 7625
rect 32375 7590 32385 7625
rect 32420 7590 32430 7625
rect 32465 7590 32475 7625
rect 32510 7590 32520 7625
rect 32555 7590 32565 7625
rect 32600 7590 32610 7625
rect 32645 7590 32655 7625
rect 32690 7590 32700 7625
rect 32735 7590 32745 7625
rect 32780 7590 32790 7625
rect 32825 7590 32835 7625
rect 32870 7590 32890 7625
rect 31290 7580 32890 7590
rect 31290 7545 31305 7580
rect 31340 7545 31350 7580
rect 31385 7545 31395 7580
rect 31430 7545 31440 7580
rect 31475 7545 31485 7580
rect 31520 7545 31530 7580
rect 31565 7545 31575 7580
rect 31610 7545 31620 7580
rect 31655 7545 31665 7580
rect 31700 7545 31710 7580
rect 31745 7545 31755 7580
rect 31790 7545 31800 7580
rect 31835 7545 31845 7580
rect 31880 7545 31890 7580
rect 31925 7545 31935 7580
rect 31970 7545 31980 7580
rect 32015 7545 32025 7580
rect 32060 7545 32070 7580
rect 32105 7545 32115 7580
rect 32150 7545 32160 7580
rect 32195 7545 32205 7580
rect 32240 7545 32250 7580
rect 32285 7545 32295 7580
rect 32330 7545 32340 7580
rect 32375 7545 32385 7580
rect 32420 7545 32430 7580
rect 32465 7545 32475 7580
rect 32510 7545 32520 7580
rect 32555 7545 32565 7580
rect 32600 7545 32610 7580
rect 32645 7545 32655 7580
rect 32690 7545 32700 7580
rect 32735 7545 32745 7580
rect 32780 7545 32790 7580
rect 32825 7545 32835 7580
rect 32870 7545 32890 7580
rect 31290 7535 32890 7545
rect 31290 7500 31305 7535
rect 31340 7500 31350 7535
rect 31385 7500 31395 7535
rect 31430 7500 31440 7535
rect 31475 7500 31485 7535
rect 31520 7500 31530 7535
rect 31565 7500 31575 7535
rect 31610 7500 31620 7535
rect 31655 7500 31665 7535
rect 31700 7500 31710 7535
rect 31745 7500 31755 7535
rect 31790 7500 31800 7535
rect 31835 7500 31845 7535
rect 31880 7500 31890 7535
rect 31925 7500 31935 7535
rect 31970 7500 31980 7535
rect 32015 7500 32025 7535
rect 32060 7500 32070 7535
rect 32105 7500 32115 7535
rect 32150 7500 32160 7535
rect 32195 7500 32205 7535
rect 32240 7500 32250 7535
rect 32285 7500 32295 7535
rect 32330 7500 32340 7535
rect 32375 7500 32385 7535
rect 32420 7500 32430 7535
rect 32465 7500 32475 7535
rect 32510 7500 32520 7535
rect 32555 7500 32565 7535
rect 32600 7500 32610 7535
rect 32645 7500 32655 7535
rect 32690 7500 32700 7535
rect 32735 7500 32745 7535
rect 32780 7500 32790 7535
rect 32825 7500 32835 7535
rect 32870 7500 32890 7535
rect 31290 7490 32890 7500
rect 31290 7455 31305 7490
rect 31340 7455 31350 7490
rect 31385 7455 31395 7490
rect 31430 7455 31440 7490
rect 31475 7455 31485 7490
rect 31520 7455 31530 7490
rect 31565 7455 31575 7490
rect 31610 7455 31620 7490
rect 31655 7455 31665 7490
rect 31700 7455 31710 7490
rect 31745 7455 31755 7490
rect 31790 7455 31800 7490
rect 31835 7455 31845 7490
rect 31880 7455 31890 7490
rect 31925 7455 31935 7490
rect 31970 7455 31980 7490
rect 32015 7455 32025 7490
rect 32060 7455 32070 7490
rect 32105 7455 32115 7490
rect 32150 7455 32160 7490
rect 32195 7455 32205 7490
rect 32240 7455 32250 7490
rect 32285 7455 32295 7490
rect 32330 7455 32340 7490
rect 32375 7455 32385 7490
rect 32420 7455 32430 7490
rect 32465 7455 32475 7490
rect 32510 7455 32520 7490
rect 32555 7455 32565 7490
rect 32600 7455 32610 7490
rect 32645 7455 32655 7490
rect 32690 7455 32700 7490
rect 32735 7455 32745 7490
rect 32780 7455 32790 7490
rect 32825 7455 32835 7490
rect 32870 7455 32890 7490
rect 31290 7445 32890 7455
rect 31290 7410 31305 7445
rect 31340 7410 31350 7445
rect 31385 7410 31395 7445
rect 31430 7410 31440 7445
rect 31475 7410 31485 7445
rect 31520 7410 31530 7445
rect 31565 7410 31575 7445
rect 31610 7410 31620 7445
rect 31655 7410 31665 7445
rect 31700 7410 31710 7445
rect 31745 7410 31755 7445
rect 31790 7410 31800 7445
rect 31835 7410 31845 7445
rect 31880 7410 31890 7445
rect 31925 7410 31935 7445
rect 31970 7410 31980 7445
rect 32015 7410 32025 7445
rect 32060 7410 32070 7445
rect 32105 7410 32115 7445
rect 32150 7410 32160 7445
rect 32195 7410 32205 7445
rect 32240 7410 32250 7445
rect 32285 7410 32295 7445
rect 32330 7410 32340 7445
rect 32375 7410 32385 7445
rect 32420 7410 32430 7445
rect 32465 7410 32475 7445
rect 32510 7410 32520 7445
rect 32555 7410 32565 7445
rect 32600 7410 32610 7445
rect 32645 7410 32655 7445
rect 32690 7410 32700 7445
rect 32735 7410 32745 7445
rect 32780 7410 32790 7445
rect 32825 7410 32835 7445
rect 32870 7410 32890 7445
rect 31290 7400 32890 7410
rect 31290 7365 31305 7400
rect 31340 7365 31350 7400
rect 31385 7365 31395 7400
rect 31430 7365 31440 7400
rect 31475 7365 31485 7400
rect 31520 7365 31530 7400
rect 31565 7365 31575 7400
rect 31610 7365 31620 7400
rect 31655 7365 31665 7400
rect 31700 7365 31710 7400
rect 31745 7365 31755 7400
rect 31790 7365 31800 7400
rect 31835 7365 31845 7400
rect 31880 7365 31890 7400
rect 31925 7365 31935 7400
rect 31970 7365 31980 7400
rect 32015 7365 32025 7400
rect 32060 7365 32070 7400
rect 32105 7365 32115 7400
rect 32150 7365 32160 7400
rect 32195 7365 32205 7400
rect 32240 7365 32250 7400
rect 32285 7365 32295 7400
rect 32330 7365 32340 7400
rect 32375 7365 32385 7400
rect 32420 7365 32430 7400
rect 32465 7365 32475 7400
rect 32510 7365 32520 7400
rect 32555 7365 32565 7400
rect 32600 7365 32610 7400
rect 32645 7365 32655 7400
rect 32690 7365 32700 7400
rect 32735 7365 32745 7400
rect 32780 7365 32790 7400
rect 32825 7365 32835 7400
rect 32870 7365 32890 7400
rect 31290 7355 32890 7365
rect 31290 7320 31305 7355
rect 31340 7320 31350 7355
rect 31385 7320 31395 7355
rect 31430 7320 31440 7355
rect 31475 7320 31485 7355
rect 31520 7320 31530 7355
rect 31565 7320 31575 7355
rect 31610 7320 31620 7355
rect 31655 7320 31665 7355
rect 31700 7320 31710 7355
rect 31745 7320 31755 7355
rect 31790 7320 31800 7355
rect 31835 7320 31845 7355
rect 31880 7320 31890 7355
rect 31925 7320 31935 7355
rect 31970 7320 31980 7355
rect 32015 7320 32025 7355
rect 32060 7320 32070 7355
rect 32105 7320 32115 7355
rect 32150 7320 32160 7355
rect 32195 7320 32205 7355
rect 32240 7320 32250 7355
rect 32285 7320 32295 7355
rect 32330 7320 32340 7355
rect 32375 7320 32385 7355
rect 32420 7320 32430 7355
rect 32465 7320 32475 7355
rect 32510 7320 32520 7355
rect 32555 7320 32565 7355
rect 32600 7320 32610 7355
rect 32645 7320 32655 7355
rect 32690 7320 32700 7355
rect 32735 7320 32745 7355
rect 32780 7320 32790 7355
rect 32825 7320 32835 7355
rect 32870 7320 32890 7355
rect 31290 7310 32890 7320
rect 31290 7275 31305 7310
rect 31340 7275 31350 7310
rect 31385 7275 31395 7310
rect 31430 7275 31440 7310
rect 31475 7275 31485 7310
rect 31520 7275 31530 7310
rect 31565 7275 31575 7310
rect 31610 7275 31620 7310
rect 31655 7275 31665 7310
rect 31700 7275 31710 7310
rect 31745 7275 31755 7310
rect 31790 7275 31800 7310
rect 31835 7275 31845 7310
rect 31880 7275 31890 7310
rect 31925 7275 31935 7310
rect 31970 7275 31980 7310
rect 32015 7275 32025 7310
rect 32060 7275 32070 7310
rect 32105 7275 32115 7310
rect 32150 7275 32160 7310
rect 32195 7275 32205 7310
rect 32240 7275 32250 7310
rect 32285 7275 32295 7310
rect 32330 7275 32340 7310
rect 32375 7275 32385 7310
rect 32420 7275 32430 7310
rect 32465 7275 32475 7310
rect 32510 7275 32520 7310
rect 32555 7275 32565 7310
rect 32600 7275 32610 7310
rect 32645 7275 32655 7310
rect 32690 7275 32700 7310
rect 32735 7275 32745 7310
rect 32780 7275 32790 7310
rect 32825 7275 32835 7310
rect 32870 7275 32890 7310
rect 31290 7265 32890 7275
rect 31290 7230 31305 7265
rect 31340 7230 31350 7265
rect 31385 7230 31395 7265
rect 31430 7230 31440 7265
rect 31475 7230 31485 7265
rect 31520 7230 31530 7265
rect 31565 7230 31575 7265
rect 31610 7230 31620 7265
rect 31655 7230 31665 7265
rect 31700 7230 31710 7265
rect 31745 7230 31755 7265
rect 31790 7230 31800 7265
rect 31835 7230 31845 7265
rect 31880 7230 31890 7265
rect 31925 7230 31935 7265
rect 31970 7230 31980 7265
rect 32015 7230 32025 7265
rect 32060 7230 32070 7265
rect 32105 7230 32115 7265
rect 32150 7230 32160 7265
rect 32195 7230 32205 7265
rect 32240 7230 32250 7265
rect 32285 7230 32295 7265
rect 32330 7230 32340 7265
rect 32375 7230 32385 7265
rect 32420 7230 32430 7265
rect 32465 7230 32475 7265
rect 32510 7230 32520 7265
rect 32555 7230 32565 7265
rect 32600 7230 32610 7265
rect 32645 7230 32655 7265
rect 32690 7230 32700 7265
rect 32735 7230 32745 7265
rect 32780 7230 32790 7265
rect 32825 7230 32835 7265
rect 32870 7230 32890 7265
rect 31290 7220 32890 7230
rect 31290 7185 31305 7220
rect 31340 7185 31350 7220
rect 31385 7185 31395 7220
rect 31430 7185 31440 7220
rect 31475 7185 31485 7220
rect 31520 7185 31530 7220
rect 31565 7185 31575 7220
rect 31610 7185 31620 7220
rect 31655 7185 31665 7220
rect 31700 7185 31710 7220
rect 31745 7185 31755 7220
rect 31790 7185 31800 7220
rect 31835 7185 31845 7220
rect 31880 7185 31890 7220
rect 31925 7185 31935 7220
rect 31970 7185 31980 7220
rect 32015 7185 32025 7220
rect 32060 7185 32070 7220
rect 32105 7185 32115 7220
rect 32150 7185 32160 7220
rect 32195 7185 32205 7220
rect 32240 7185 32250 7220
rect 32285 7185 32295 7220
rect 32330 7185 32340 7220
rect 32375 7185 32385 7220
rect 32420 7185 32430 7220
rect 32465 7185 32475 7220
rect 32510 7185 32520 7220
rect 32555 7185 32565 7220
rect 32600 7185 32610 7220
rect 32645 7185 32655 7220
rect 32690 7185 32700 7220
rect 32735 7185 32745 7220
rect 32780 7185 32790 7220
rect 32825 7185 32835 7220
rect 32870 7185 32890 7220
rect 31290 7175 32890 7185
rect 31290 7140 31305 7175
rect 31340 7140 31350 7175
rect 31385 7140 31395 7175
rect 31430 7140 31440 7175
rect 31475 7140 31485 7175
rect 31520 7140 31530 7175
rect 31565 7140 31575 7175
rect 31610 7140 31620 7175
rect 31655 7140 31665 7175
rect 31700 7140 31710 7175
rect 31745 7140 31755 7175
rect 31790 7140 31800 7175
rect 31835 7140 31845 7175
rect 31880 7140 31890 7175
rect 31925 7140 31935 7175
rect 31970 7140 31980 7175
rect 32015 7140 32025 7175
rect 32060 7140 32070 7175
rect 32105 7140 32115 7175
rect 32150 7140 32160 7175
rect 32195 7140 32205 7175
rect 32240 7140 32250 7175
rect 32285 7140 32295 7175
rect 32330 7140 32340 7175
rect 32375 7140 32385 7175
rect 32420 7140 32430 7175
rect 32465 7140 32475 7175
rect 32510 7140 32520 7175
rect 32555 7140 32565 7175
rect 32600 7140 32610 7175
rect 32645 7140 32655 7175
rect 32690 7140 32700 7175
rect 32735 7140 32745 7175
rect 32780 7140 32790 7175
rect 32825 7140 32835 7175
rect 32870 7140 32890 7175
rect 31290 7130 32890 7140
rect 31290 7095 31305 7130
rect 31340 7095 31350 7130
rect 31385 7095 31395 7130
rect 31430 7095 31440 7130
rect 31475 7095 31485 7130
rect 31520 7095 31530 7130
rect 31565 7095 31575 7130
rect 31610 7095 31620 7130
rect 31655 7095 31665 7130
rect 31700 7095 31710 7130
rect 31745 7095 31755 7130
rect 31790 7095 31800 7130
rect 31835 7095 31845 7130
rect 31880 7095 31890 7130
rect 31925 7095 31935 7130
rect 31970 7095 31980 7130
rect 32015 7095 32025 7130
rect 32060 7095 32070 7130
rect 32105 7095 32115 7130
rect 32150 7095 32160 7130
rect 32195 7095 32205 7130
rect 32240 7095 32250 7130
rect 32285 7095 32295 7130
rect 32330 7095 32340 7130
rect 32375 7095 32385 7130
rect 32420 7095 32430 7130
rect 32465 7095 32475 7130
rect 32510 7095 32520 7130
rect 32555 7095 32565 7130
rect 32600 7095 32610 7130
rect 32645 7095 32655 7130
rect 32690 7095 32700 7130
rect 32735 7095 32745 7130
rect 32780 7095 32790 7130
rect 32825 7095 32835 7130
rect 32870 7095 32890 7130
rect 31290 7085 32890 7095
rect 31290 7050 31305 7085
rect 31340 7050 31350 7085
rect 31385 7050 31395 7085
rect 31430 7050 31440 7085
rect 31475 7050 31485 7085
rect 31520 7050 31530 7085
rect 31565 7050 31575 7085
rect 31610 7050 31620 7085
rect 31655 7050 31665 7085
rect 31700 7050 31710 7085
rect 31745 7050 31755 7085
rect 31790 7050 31800 7085
rect 31835 7050 31845 7085
rect 31880 7050 31890 7085
rect 31925 7050 31935 7085
rect 31970 7050 31980 7085
rect 32015 7050 32025 7085
rect 32060 7050 32070 7085
rect 32105 7050 32115 7085
rect 32150 7050 32160 7085
rect 32195 7050 32205 7085
rect 32240 7050 32250 7085
rect 32285 7050 32295 7085
rect 32330 7050 32340 7085
rect 32375 7050 32385 7085
rect 32420 7050 32430 7085
rect 32465 7050 32475 7085
rect 32510 7050 32520 7085
rect 32555 7050 32565 7085
rect 32600 7050 32610 7085
rect 32645 7050 32655 7085
rect 32690 7050 32700 7085
rect 32735 7050 32745 7085
rect 32780 7050 32790 7085
rect 32825 7050 32835 7085
rect 32870 7050 32890 7085
rect 31290 7040 32890 7050
rect 31290 7005 31305 7040
rect 31340 7005 31350 7040
rect 31385 7005 31395 7040
rect 31430 7005 31440 7040
rect 31475 7005 31485 7040
rect 31520 7005 31530 7040
rect 31565 7005 31575 7040
rect 31610 7005 31620 7040
rect 31655 7005 31665 7040
rect 31700 7005 31710 7040
rect 31745 7005 31755 7040
rect 31790 7005 31800 7040
rect 31835 7005 31845 7040
rect 31880 7005 31890 7040
rect 31925 7005 31935 7040
rect 31970 7005 31980 7040
rect 32015 7005 32025 7040
rect 32060 7005 32070 7040
rect 32105 7005 32115 7040
rect 32150 7005 32160 7040
rect 32195 7005 32205 7040
rect 32240 7005 32250 7040
rect 32285 7005 32295 7040
rect 32330 7005 32340 7040
rect 32375 7005 32385 7040
rect 32420 7005 32430 7040
rect 32465 7005 32475 7040
rect 32510 7005 32520 7040
rect 32555 7005 32565 7040
rect 32600 7005 32610 7040
rect 32645 7005 32655 7040
rect 32690 7005 32700 7040
rect 32735 7005 32745 7040
rect 32780 7005 32790 7040
rect 32825 7005 32835 7040
rect 32870 7005 32890 7040
rect 31290 6995 32890 7005
rect 31290 6960 31305 6995
rect 31340 6960 31350 6995
rect 31385 6960 31395 6995
rect 31430 6960 31440 6995
rect 31475 6960 31485 6995
rect 31520 6960 31530 6995
rect 31565 6960 31575 6995
rect 31610 6960 31620 6995
rect 31655 6960 31665 6995
rect 31700 6960 31710 6995
rect 31745 6960 31755 6995
rect 31790 6960 31800 6995
rect 31835 6960 31845 6995
rect 31880 6960 31890 6995
rect 31925 6960 31935 6995
rect 31970 6960 31980 6995
rect 32015 6960 32025 6995
rect 32060 6960 32070 6995
rect 32105 6960 32115 6995
rect 32150 6960 32160 6995
rect 32195 6960 32205 6995
rect 32240 6960 32250 6995
rect 32285 6960 32295 6995
rect 32330 6960 32340 6995
rect 32375 6960 32385 6995
rect 32420 6960 32430 6995
rect 32465 6960 32475 6995
rect 32510 6960 32520 6995
rect 32555 6960 32565 6995
rect 32600 6960 32610 6995
rect 32645 6960 32655 6995
rect 32690 6960 32700 6995
rect 32735 6960 32745 6995
rect 32780 6960 32790 6995
rect 32825 6960 32835 6995
rect 32870 6960 32890 6995
rect 31290 6950 32890 6960
rect 31290 6915 31305 6950
rect 31340 6915 31350 6950
rect 31385 6915 31395 6950
rect 31430 6915 31440 6950
rect 31475 6915 31485 6950
rect 31520 6915 31530 6950
rect 31565 6915 31575 6950
rect 31610 6915 31620 6950
rect 31655 6915 31665 6950
rect 31700 6915 31710 6950
rect 31745 6915 31755 6950
rect 31790 6915 31800 6950
rect 31835 6915 31845 6950
rect 31880 6915 31890 6950
rect 31925 6915 31935 6950
rect 31970 6915 31980 6950
rect 32015 6915 32025 6950
rect 32060 6915 32070 6950
rect 32105 6915 32115 6950
rect 32150 6915 32160 6950
rect 32195 6915 32205 6950
rect 32240 6915 32250 6950
rect 32285 6915 32295 6950
rect 32330 6915 32340 6950
rect 32375 6915 32385 6950
rect 32420 6915 32430 6950
rect 32465 6915 32475 6950
rect 32510 6915 32520 6950
rect 32555 6915 32565 6950
rect 32600 6915 32610 6950
rect 32645 6915 32655 6950
rect 32690 6915 32700 6950
rect 32735 6915 32745 6950
rect 32780 6915 32790 6950
rect 32825 6915 32835 6950
rect 32870 6915 32890 6950
rect 31290 6905 32890 6915
rect 31290 6870 31305 6905
rect 31340 6870 31350 6905
rect 31385 6870 31395 6905
rect 31430 6870 31440 6905
rect 31475 6870 31485 6905
rect 31520 6870 31530 6905
rect 31565 6870 31575 6905
rect 31610 6870 31620 6905
rect 31655 6870 31665 6905
rect 31700 6870 31710 6905
rect 31745 6870 31755 6905
rect 31790 6870 31800 6905
rect 31835 6870 31845 6905
rect 31880 6870 31890 6905
rect 31925 6870 31935 6905
rect 31970 6870 31980 6905
rect 32015 6870 32025 6905
rect 32060 6870 32070 6905
rect 32105 6870 32115 6905
rect 32150 6870 32160 6905
rect 32195 6870 32205 6905
rect 32240 6870 32250 6905
rect 32285 6870 32295 6905
rect 32330 6870 32340 6905
rect 32375 6870 32385 6905
rect 32420 6870 32430 6905
rect 32465 6870 32475 6905
rect 32510 6870 32520 6905
rect 32555 6870 32565 6905
rect 32600 6870 32610 6905
rect 32645 6870 32655 6905
rect 32690 6870 32700 6905
rect 32735 6870 32745 6905
rect 32780 6870 32790 6905
rect 32825 6870 32835 6905
rect 32870 6870 32890 6905
rect 31290 6860 32890 6870
rect 31290 6825 31305 6860
rect 31340 6825 31350 6860
rect 31385 6825 31395 6860
rect 31430 6825 31440 6860
rect 31475 6825 31485 6860
rect 31520 6825 31530 6860
rect 31565 6825 31575 6860
rect 31610 6825 31620 6860
rect 31655 6825 31665 6860
rect 31700 6825 31710 6860
rect 31745 6825 31755 6860
rect 31790 6825 31800 6860
rect 31835 6825 31845 6860
rect 31880 6825 31890 6860
rect 31925 6825 31935 6860
rect 31970 6825 31980 6860
rect 32015 6825 32025 6860
rect 32060 6825 32070 6860
rect 32105 6825 32115 6860
rect 32150 6825 32160 6860
rect 32195 6825 32205 6860
rect 32240 6825 32250 6860
rect 32285 6825 32295 6860
rect 32330 6825 32340 6860
rect 32375 6825 32385 6860
rect 32420 6825 32430 6860
rect 32465 6825 32475 6860
rect 32510 6825 32520 6860
rect 32555 6825 32565 6860
rect 32600 6825 32610 6860
rect 32645 6825 32655 6860
rect 32690 6825 32700 6860
rect 32735 6825 32745 6860
rect 32780 6825 32790 6860
rect 32825 6825 32835 6860
rect 32870 6825 32890 6860
rect 31290 6815 32890 6825
rect 31290 6780 31305 6815
rect 31340 6780 31350 6815
rect 31385 6780 31395 6815
rect 31430 6780 31440 6815
rect 31475 6780 31485 6815
rect 31520 6780 31530 6815
rect 31565 6780 31575 6815
rect 31610 6780 31620 6815
rect 31655 6780 31665 6815
rect 31700 6780 31710 6815
rect 31745 6780 31755 6815
rect 31790 6780 31800 6815
rect 31835 6780 31845 6815
rect 31880 6780 31890 6815
rect 31925 6780 31935 6815
rect 31970 6780 31980 6815
rect 32015 6780 32025 6815
rect 32060 6780 32070 6815
rect 32105 6780 32115 6815
rect 32150 6780 32160 6815
rect 32195 6780 32205 6815
rect 32240 6780 32250 6815
rect 32285 6780 32295 6815
rect 32330 6780 32340 6815
rect 32375 6780 32385 6815
rect 32420 6780 32430 6815
rect 32465 6780 32475 6815
rect 32510 6780 32520 6815
rect 32555 6780 32565 6815
rect 32600 6780 32610 6815
rect 32645 6780 32655 6815
rect 32690 6780 32700 6815
rect 32735 6780 32745 6815
rect 32780 6780 32790 6815
rect 32825 6780 32835 6815
rect 32870 6780 32890 6815
rect 31290 6770 32890 6780
rect 31290 6735 31305 6770
rect 31340 6735 31350 6770
rect 31385 6735 31395 6770
rect 31430 6735 31440 6770
rect 31475 6735 31485 6770
rect 31520 6735 31530 6770
rect 31565 6735 31575 6770
rect 31610 6735 31620 6770
rect 31655 6735 31665 6770
rect 31700 6735 31710 6770
rect 31745 6735 31755 6770
rect 31790 6735 31800 6770
rect 31835 6735 31845 6770
rect 31880 6735 31890 6770
rect 31925 6735 31935 6770
rect 31970 6735 31980 6770
rect 32015 6735 32025 6770
rect 32060 6735 32070 6770
rect 32105 6735 32115 6770
rect 32150 6735 32160 6770
rect 32195 6735 32205 6770
rect 32240 6735 32250 6770
rect 32285 6735 32295 6770
rect 32330 6735 32340 6770
rect 32375 6735 32385 6770
rect 32420 6735 32430 6770
rect 32465 6735 32475 6770
rect 32510 6735 32520 6770
rect 32555 6735 32565 6770
rect 32600 6735 32610 6770
rect 32645 6735 32655 6770
rect 32690 6735 32700 6770
rect 32735 6735 32745 6770
rect 32780 6735 32790 6770
rect 32825 6735 32835 6770
rect 32870 6735 32890 6770
rect 31290 6725 32890 6735
rect 31290 6690 31305 6725
rect 31340 6690 31350 6725
rect 31385 6690 31395 6725
rect 31430 6690 31440 6725
rect 31475 6690 31485 6725
rect 31520 6690 31530 6725
rect 31565 6690 31575 6725
rect 31610 6690 31620 6725
rect 31655 6690 31665 6725
rect 31700 6690 31710 6725
rect 31745 6690 31755 6725
rect 31790 6690 31800 6725
rect 31835 6690 31845 6725
rect 31880 6690 31890 6725
rect 31925 6690 31935 6725
rect 31970 6690 31980 6725
rect 32015 6690 32025 6725
rect 32060 6690 32070 6725
rect 32105 6690 32115 6725
rect 32150 6690 32160 6725
rect 32195 6690 32205 6725
rect 32240 6690 32250 6725
rect 32285 6690 32295 6725
rect 32330 6690 32340 6725
rect 32375 6690 32385 6725
rect 32420 6690 32430 6725
rect 32465 6690 32475 6725
rect 32510 6690 32520 6725
rect 32555 6690 32565 6725
rect 32600 6690 32610 6725
rect 32645 6690 32655 6725
rect 32690 6690 32700 6725
rect 32735 6690 32745 6725
rect 32780 6690 32790 6725
rect 32825 6690 32835 6725
rect 32870 6690 32890 6725
rect 31290 6680 32890 6690
rect 31290 6645 31305 6680
rect 31340 6645 31350 6680
rect 31385 6645 31395 6680
rect 31430 6645 31440 6680
rect 31475 6645 31485 6680
rect 31520 6645 31530 6680
rect 31565 6645 31575 6680
rect 31610 6645 31620 6680
rect 31655 6645 31665 6680
rect 31700 6645 31710 6680
rect 31745 6645 31755 6680
rect 31790 6645 31800 6680
rect 31835 6645 31845 6680
rect 31880 6645 31890 6680
rect 31925 6645 31935 6680
rect 31970 6645 31980 6680
rect 32015 6645 32025 6680
rect 32060 6645 32070 6680
rect 32105 6645 32115 6680
rect 32150 6645 32160 6680
rect 32195 6645 32205 6680
rect 32240 6645 32250 6680
rect 32285 6645 32295 6680
rect 32330 6645 32340 6680
rect 32375 6645 32385 6680
rect 32420 6645 32430 6680
rect 32465 6645 32475 6680
rect 32510 6645 32520 6680
rect 32555 6645 32565 6680
rect 32600 6645 32610 6680
rect 32645 6645 32655 6680
rect 32690 6645 32700 6680
rect 32735 6645 32745 6680
rect 32780 6645 32790 6680
rect 32825 6645 32835 6680
rect 32870 6645 32890 6680
rect 31290 6635 32890 6645
rect 31290 6600 31305 6635
rect 31340 6600 31350 6635
rect 31385 6600 31395 6635
rect 31430 6600 31440 6635
rect 31475 6600 31485 6635
rect 31520 6600 31530 6635
rect 31565 6600 31575 6635
rect 31610 6600 31620 6635
rect 31655 6600 31665 6635
rect 31700 6600 31710 6635
rect 31745 6600 31755 6635
rect 31790 6600 31800 6635
rect 31835 6600 31845 6635
rect 31880 6600 31890 6635
rect 31925 6600 31935 6635
rect 31970 6600 31980 6635
rect 32015 6600 32025 6635
rect 32060 6600 32070 6635
rect 32105 6600 32115 6635
rect 32150 6600 32160 6635
rect 32195 6600 32205 6635
rect 32240 6600 32250 6635
rect 32285 6600 32295 6635
rect 32330 6600 32340 6635
rect 32375 6600 32385 6635
rect 32420 6600 32430 6635
rect 32465 6600 32475 6635
rect 32510 6600 32520 6635
rect 32555 6600 32565 6635
rect 32600 6600 32610 6635
rect 32645 6600 32655 6635
rect 32690 6600 32700 6635
rect 32735 6600 32745 6635
rect 32780 6600 32790 6635
rect 32825 6600 32835 6635
rect 32870 6600 32890 6635
rect 31290 6590 32890 6600
rect 31290 6555 31305 6590
rect 31340 6555 31350 6590
rect 31385 6555 31395 6590
rect 31430 6555 31440 6590
rect 31475 6555 31485 6590
rect 31520 6555 31530 6590
rect 31565 6555 31575 6590
rect 31610 6555 31620 6590
rect 31655 6555 31665 6590
rect 31700 6555 31710 6590
rect 31745 6555 31755 6590
rect 31790 6555 31800 6590
rect 31835 6555 31845 6590
rect 31880 6555 31890 6590
rect 31925 6555 31935 6590
rect 31970 6555 31980 6590
rect 32015 6555 32025 6590
rect 32060 6555 32070 6590
rect 32105 6555 32115 6590
rect 32150 6555 32160 6590
rect 32195 6555 32205 6590
rect 32240 6555 32250 6590
rect 32285 6555 32295 6590
rect 32330 6555 32340 6590
rect 32375 6555 32385 6590
rect 32420 6555 32430 6590
rect 32465 6555 32475 6590
rect 32510 6555 32520 6590
rect 32555 6555 32565 6590
rect 32600 6555 32610 6590
rect 32645 6555 32655 6590
rect 32690 6555 32700 6590
rect 32735 6555 32745 6590
rect 32780 6555 32790 6590
rect 32825 6555 32835 6590
rect 32870 6555 32890 6590
rect 31290 6545 32890 6555
rect 31290 6510 31305 6545
rect 31340 6510 31350 6545
rect 31385 6510 31395 6545
rect 31430 6510 31440 6545
rect 31475 6510 31485 6545
rect 31520 6510 31530 6545
rect 31565 6510 31575 6545
rect 31610 6510 31620 6545
rect 31655 6510 31665 6545
rect 31700 6510 31710 6545
rect 31745 6510 31755 6545
rect 31790 6510 31800 6545
rect 31835 6510 31845 6545
rect 31880 6510 31890 6545
rect 31925 6510 31935 6545
rect 31970 6510 31980 6545
rect 32015 6510 32025 6545
rect 32060 6510 32070 6545
rect 32105 6510 32115 6545
rect 32150 6510 32160 6545
rect 32195 6510 32205 6545
rect 32240 6510 32250 6545
rect 32285 6510 32295 6545
rect 32330 6510 32340 6545
rect 32375 6510 32385 6545
rect 32420 6510 32430 6545
rect 32465 6510 32475 6545
rect 32510 6510 32520 6545
rect 32555 6510 32565 6545
rect 32600 6510 32610 6545
rect 32645 6510 32655 6545
rect 32690 6510 32700 6545
rect 32735 6510 32745 6545
rect 32780 6510 32790 6545
rect 32825 6510 32835 6545
rect 32870 6510 32890 6545
rect 31290 6500 32890 6510
rect 31290 6465 31305 6500
rect 31340 6465 31350 6500
rect 31385 6465 31395 6500
rect 31430 6465 31440 6500
rect 31475 6465 31485 6500
rect 31520 6465 31530 6500
rect 31565 6465 31575 6500
rect 31610 6465 31620 6500
rect 31655 6465 31665 6500
rect 31700 6465 31710 6500
rect 31745 6465 31755 6500
rect 31790 6465 31800 6500
rect 31835 6465 31845 6500
rect 31880 6465 31890 6500
rect 31925 6465 31935 6500
rect 31970 6465 31980 6500
rect 32015 6465 32025 6500
rect 32060 6465 32070 6500
rect 32105 6465 32115 6500
rect 32150 6465 32160 6500
rect 32195 6465 32205 6500
rect 32240 6465 32250 6500
rect 32285 6465 32295 6500
rect 32330 6465 32340 6500
rect 32375 6465 32385 6500
rect 32420 6465 32430 6500
rect 32465 6465 32475 6500
rect 32510 6465 32520 6500
rect 32555 6465 32565 6500
rect 32600 6465 32610 6500
rect 32645 6465 32655 6500
rect 32690 6465 32700 6500
rect 32735 6465 32745 6500
rect 32780 6465 32790 6500
rect 32825 6465 32835 6500
rect 32870 6465 32890 6500
rect -90 -1315 -30 -1305
rect -90 -1355 -80 -1315
rect -40 -1355 -30 -1315
rect -90 -1380 -30 -1355
rect -90 -1420 -80 -1380
rect -40 -1420 -30 -1380
rect -90 -1450 -30 -1420
rect -90 -1490 -80 -1450
rect -40 -1490 -30 -1450
rect -90 -1520 -30 -1490
rect -90 -1560 -80 -1520
rect -40 -1560 -30 -1520
rect -90 -1590 -30 -1560
rect -90 -1630 -80 -1590
rect -40 -1630 -30 -1590
rect -90 -1655 -30 -1630
rect -90 -1695 -80 -1655
rect -40 -1695 -30 -1655
rect -90 -1715 -30 -1695
rect -90 -1755 -80 -1715
rect -40 -1755 -30 -1715
rect -90 -1780 -30 -1755
rect -90 -1820 -80 -1780
rect -40 -1820 -30 -1780
rect -90 -1850 -30 -1820
rect -90 -1890 -80 -1850
rect -40 -1890 -30 -1850
rect -90 -1920 -30 -1890
rect -90 -1960 -80 -1920
rect -40 -1960 -30 -1920
rect -90 -1990 -30 -1960
rect -90 -2030 -80 -1990
rect -40 -2030 -30 -1990
rect -90 -2055 -30 -2030
rect -90 -2095 -80 -2055
rect -40 -2095 -30 -2055
rect -90 -2115 -30 -2095
rect -90 -2155 -80 -2115
rect -40 -2155 -30 -2115
rect -90 -2180 -30 -2155
rect -90 -2220 -80 -2180
rect -40 -2220 -30 -2180
rect -90 -2250 -30 -2220
rect -90 -2290 -80 -2250
rect -40 -2290 -30 -2250
rect -90 -2320 -30 -2290
rect -90 -2360 -80 -2320
rect -40 -2360 -30 -2320
rect -90 -2390 -30 -2360
rect -90 -2430 -80 -2390
rect -40 -2430 -30 -2390
rect -90 -2455 -30 -2430
rect -90 -2495 -80 -2455
rect -40 -2495 -30 -2455
rect -90 -2515 -30 -2495
rect -90 -2555 -80 -2515
rect -40 -2555 -30 -2515
rect -90 -2580 -30 -2555
rect -90 -2620 -80 -2580
rect -40 -2620 -30 -2580
rect -90 -2650 -30 -2620
rect -90 -2690 -80 -2650
rect -40 -2690 -30 -2650
rect -90 -2720 -30 -2690
rect -90 -2760 -80 -2720
rect -40 -2760 -30 -2720
rect -90 -2790 -30 -2760
rect -90 -2830 -80 -2790
rect -40 -2830 -30 -2790
rect -90 -2855 -30 -2830
rect -90 -2895 -80 -2855
rect -40 -2895 -30 -2855
rect -90 -2905 -30 -2895
rect 260 -1315 320 -1305
rect 260 -1355 270 -1315
rect 310 -1355 320 -1315
rect 260 -1380 320 -1355
rect 260 -1420 270 -1380
rect 310 -1420 320 -1380
rect 260 -1450 320 -1420
rect 260 -1490 270 -1450
rect 310 -1490 320 -1450
rect 260 -1520 320 -1490
rect 260 -1560 270 -1520
rect 310 -1560 320 -1520
rect 260 -1590 320 -1560
rect 260 -1630 270 -1590
rect 310 -1630 320 -1590
rect 260 -1655 320 -1630
rect 260 -1695 270 -1655
rect 310 -1695 320 -1655
rect 260 -1715 320 -1695
rect 260 -1755 270 -1715
rect 310 -1755 320 -1715
rect 260 -1780 320 -1755
rect 260 -1820 270 -1780
rect 310 -1820 320 -1780
rect 260 -1850 320 -1820
rect 260 -1890 270 -1850
rect 310 -1890 320 -1850
rect 260 -1920 320 -1890
rect 260 -1960 270 -1920
rect 310 -1960 320 -1920
rect 260 -1990 320 -1960
rect 260 -2030 270 -1990
rect 310 -2030 320 -1990
rect 260 -2055 320 -2030
rect 260 -2095 270 -2055
rect 310 -2095 320 -2055
rect 260 -2115 320 -2095
rect 260 -2155 270 -2115
rect 310 -2155 320 -2115
rect 260 -2180 320 -2155
rect 260 -2220 270 -2180
rect 310 -2220 320 -2180
rect 260 -2250 320 -2220
rect 260 -2290 270 -2250
rect 310 -2290 320 -2250
rect 260 -2320 320 -2290
rect 260 -2360 270 -2320
rect 310 -2360 320 -2320
rect 260 -2390 320 -2360
rect 260 -2430 270 -2390
rect 310 -2430 320 -2390
rect 260 -2455 320 -2430
rect 260 -2495 270 -2455
rect 310 -2495 320 -2455
rect 260 -2515 320 -2495
rect 260 -2555 270 -2515
rect 310 -2555 320 -2515
rect 260 -2580 320 -2555
rect 260 -2620 270 -2580
rect 310 -2620 320 -2580
rect 260 -2650 320 -2620
rect 260 -2690 270 -2650
rect 310 -2690 320 -2650
rect 260 -2720 320 -2690
rect 260 -2760 270 -2720
rect 310 -2760 320 -2720
rect 260 -2790 320 -2760
rect 260 -2830 270 -2790
rect 310 -2830 320 -2790
rect 260 -2855 320 -2830
rect 260 -2895 270 -2855
rect 310 -2895 320 -2855
rect 260 -2905 320 -2895
rect 610 -1315 670 -1305
rect 610 -1355 620 -1315
rect 660 -1355 670 -1315
rect 610 -1380 670 -1355
rect 610 -1420 620 -1380
rect 660 -1420 670 -1380
rect 610 -1450 670 -1420
rect 610 -1490 620 -1450
rect 660 -1490 670 -1450
rect 610 -1520 670 -1490
rect 610 -1560 620 -1520
rect 660 -1560 670 -1520
rect 610 -1590 670 -1560
rect 610 -1630 620 -1590
rect 660 -1630 670 -1590
rect 610 -1655 670 -1630
rect 610 -1695 620 -1655
rect 660 -1695 670 -1655
rect 610 -1715 670 -1695
rect 610 -1755 620 -1715
rect 660 -1755 670 -1715
rect 610 -1780 670 -1755
rect 610 -1820 620 -1780
rect 660 -1820 670 -1780
rect 610 -1850 670 -1820
rect 610 -1890 620 -1850
rect 660 -1890 670 -1850
rect 610 -1920 670 -1890
rect 610 -1960 620 -1920
rect 660 -1960 670 -1920
rect 610 -1990 670 -1960
rect 610 -2030 620 -1990
rect 660 -2030 670 -1990
rect 610 -2055 670 -2030
rect 610 -2095 620 -2055
rect 660 -2095 670 -2055
rect 610 -2115 670 -2095
rect 610 -2155 620 -2115
rect 660 -2155 670 -2115
rect 610 -2180 670 -2155
rect 610 -2220 620 -2180
rect 660 -2220 670 -2180
rect 610 -2250 670 -2220
rect 610 -2290 620 -2250
rect 660 -2290 670 -2250
rect 610 -2320 670 -2290
rect 610 -2360 620 -2320
rect 660 -2360 670 -2320
rect 610 -2390 670 -2360
rect 610 -2430 620 -2390
rect 660 -2430 670 -2390
rect 610 -2455 670 -2430
rect 610 -2495 620 -2455
rect 660 -2495 670 -2455
rect 610 -2515 670 -2495
rect 610 -2555 620 -2515
rect 660 -2555 670 -2515
rect 610 -2580 670 -2555
rect 610 -2620 620 -2580
rect 660 -2620 670 -2580
rect 610 -2650 670 -2620
rect 610 -2690 620 -2650
rect 660 -2690 670 -2650
rect 610 -2720 670 -2690
rect 610 -2760 620 -2720
rect 660 -2760 670 -2720
rect 610 -2790 670 -2760
rect 610 -2830 620 -2790
rect 660 -2830 670 -2790
rect 610 -2855 670 -2830
rect 610 -2895 620 -2855
rect 660 -2895 670 -2855
rect 610 -2905 670 -2895
rect 960 -1315 1020 -1305
rect 960 -1355 970 -1315
rect 1010 -1355 1020 -1315
rect 960 -1380 1020 -1355
rect 960 -1420 970 -1380
rect 1010 -1420 1020 -1380
rect 960 -1450 1020 -1420
rect 960 -1490 970 -1450
rect 1010 -1490 1020 -1450
rect 960 -1520 1020 -1490
rect 960 -1560 970 -1520
rect 1010 -1560 1020 -1520
rect 960 -1590 1020 -1560
rect 960 -1630 970 -1590
rect 1010 -1630 1020 -1590
rect 960 -1655 1020 -1630
rect 960 -1695 970 -1655
rect 1010 -1695 1020 -1655
rect 960 -1715 1020 -1695
rect 960 -1755 970 -1715
rect 1010 -1755 1020 -1715
rect 960 -1780 1020 -1755
rect 960 -1820 970 -1780
rect 1010 -1820 1020 -1780
rect 960 -1850 1020 -1820
rect 960 -1890 970 -1850
rect 1010 -1890 1020 -1850
rect 960 -1920 1020 -1890
rect 960 -1960 970 -1920
rect 1010 -1960 1020 -1920
rect 960 -1990 1020 -1960
rect 960 -2030 970 -1990
rect 1010 -2030 1020 -1990
rect 960 -2055 1020 -2030
rect 960 -2095 970 -2055
rect 1010 -2095 1020 -2055
rect 960 -2115 1020 -2095
rect 960 -2155 970 -2115
rect 1010 -2155 1020 -2115
rect 960 -2180 1020 -2155
rect 960 -2220 970 -2180
rect 1010 -2220 1020 -2180
rect 960 -2250 1020 -2220
rect 960 -2290 970 -2250
rect 1010 -2290 1020 -2250
rect 960 -2320 1020 -2290
rect 960 -2360 970 -2320
rect 1010 -2360 1020 -2320
rect 960 -2390 1020 -2360
rect 960 -2430 970 -2390
rect 1010 -2430 1020 -2390
rect 960 -2455 1020 -2430
rect 960 -2495 970 -2455
rect 1010 -2495 1020 -2455
rect 960 -2515 1020 -2495
rect 960 -2555 970 -2515
rect 1010 -2555 1020 -2515
rect 960 -2580 1020 -2555
rect 960 -2620 970 -2580
rect 1010 -2620 1020 -2580
rect 960 -2650 1020 -2620
rect 960 -2690 970 -2650
rect 1010 -2690 1020 -2650
rect 960 -2720 1020 -2690
rect 960 -2760 970 -2720
rect 1010 -2760 1020 -2720
rect 960 -2790 1020 -2760
rect 960 -2830 970 -2790
rect 1010 -2830 1020 -2790
rect 960 -2855 1020 -2830
rect 960 -2895 970 -2855
rect 1010 -2895 1020 -2855
rect 960 -2905 1020 -2895
rect 1310 -1315 1370 -1305
rect 1310 -1355 1320 -1315
rect 1360 -1355 1370 -1315
rect 1310 -1380 1370 -1355
rect 1310 -1420 1320 -1380
rect 1360 -1420 1370 -1380
rect 1310 -1450 1370 -1420
rect 1310 -1490 1320 -1450
rect 1360 -1490 1370 -1450
rect 1310 -1520 1370 -1490
rect 1310 -1560 1320 -1520
rect 1360 -1560 1370 -1520
rect 1310 -1590 1370 -1560
rect 1310 -1630 1320 -1590
rect 1360 -1630 1370 -1590
rect 1310 -1655 1370 -1630
rect 1310 -1695 1320 -1655
rect 1360 -1695 1370 -1655
rect 1310 -1715 1370 -1695
rect 1310 -1755 1320 -1715
rect 1360 -1755 1370 -1715
rect 1310 -1780 1370 -1755
rect 1310 -1820 1320 -1780
rect 1360 -1820 1370 -1780
rect 1310 -1850 1370 -1820
rect 1310 -1890 1320 -1850
rect 1360 -1890 1370 -1850
rect 1310 -1920 1370 -1890
rect 1310 -1960 1320 -1920
rect 1360 -1960 1370 -1920
rect 1310 -1990 1370 -1960
rect 1310 -2030 1320 -1990
rect 1360 -2030 1370 -1990
rect 1310 -2055 1370 -2030
rect 1310 -2095 1320 -2055
rect 1360 -2095 1370 -2055
rect 1310 -2115 1370 -2095
rect 1310 -2155 1320 -2115
rect 1360 -2155 1370 -2115
rect 1310 -2180 1370 -2155
rect 1310 -2220 1320 -2180
rect 1360 -2220 1370 -2180
rect 1310 -2250 1370 -2220
rect 1310 -2290 1320 -2250
rect 1360 -2290 1370 -2250
rect 1310 -2320 1370 -2290
rect 1310 -2360 1320 -2320
rect 1360 -2360 1370 -2320
rect 1310 -2390 1370 -2360
rect 1310 -2430 1320 -2390
rect 1360 -2430 1370 -2390
rect 1310 -2455 1370 -2430
rect 1310 -2495 1320 -2455
rect 1360 -2495 1370 -2455
rect 1310 -2515 1370 -2495
rect 1310 -2555 1320 -2515
rect 1360 -2555 1370 -2515
rect 1310 -2580 1370 -2555
rect 1310 -2620 1320 -2580
rect 1360 -2620 1370 -2580
rect 1310 -2650 1370 -2620
rect 1310 -2690 1320 -2650
rect 1360 -2690 1370 -2650
rect 1310 -2720 1370 -2690
rect 1310 -2760 1320 -2720
rect 1360 -2760 1370 -2720
rect 1310 -2790 1370 -2760
rect 1310 -2830 1320 -2790
rect 1360 -2830 1370 -2790
rect 1310 -2855 1370 -2830
rect 1310 -2895 1320 -2855
rect 1360 -2895 1370 -2855
rect 1310 -2905 1370 -2895
rect 1660 -1315 1720 -1305
rect 1660 -1355 1670 -1315
rect 1710 -1355 1720 -1315
rect 1660 -1380 1720 -1355
rect 1660 -1420 1670 -1380
rect 1710 -1420 1720 -1380
rect 1660 -1450 1720 -1420
rect 1660 -1490 1670 -1450
rect 1710 -1490 1720 -1450
rect 1660 -1520 1720 -1490
rect 1660 -1560 1670 -1520
rect 1710 -1560 1720 -1520
rect 1660 -1590 1720 -1560
rect 1660 -1630 1670 -1590
rect 1710 -1630 1720 -1590
rect 1660 -1655 1720 -1630
rect 1660 -1695 1670 -1655
rect 1710 -1695 1720 -1655
rect 1660 -1715 1720 -1695
rect 1660 -1755 1670 -1715
rect 1710 -1755 1720 -1715
rect 1660 -1780 1720 -1755
rect 1660 -1820 1670 -1780
rect 1710 -1820 1720 -1780
rect 1660 -1850 1720 -1820
rect 1660 -1890 1670 -1850
rect 1710 -1890 1720 -1850
rect 1660 -1920 1720 -1890
rect 1660 -1960 1670 -1920
rect 1710 -1960 1720 -1920
rect 1660 -1990 1720 -1960
rect 1660 -2030 1670 -1990
rect 1710 -2030 1720 -1990
rect 1660 -2055 1720 -2030
rect 1660 -2095 1670 -2055
rect 1710 -2095 1720 -2055
rect 1660 -2115 1720 -2095
rect 1660 -2155 1670 -2115
rect 1710 -2155 1720 -2115
rect 1660 -2180 1720 -2155
rect 1660 -2220 1670 -2180
rect 1710 -2220 1720 -2180
rect 1660 -2250 1720 -2220
rect 1660 -2290 1670 -2250
rect 1710 -2290 1720 -2250
rect 1660 -2320 1720 -2290
rect 1660 -2360 1670 -2320
rect 1710 -2360 1720 -2320
rect 1660 -2390 1720 -2360
rect 1660 -2430 1670 -2390
rect 1710 -2430 1720 -2390
rect 1660 -2455 1720 -2430
rect 1660 -2495 1670 -2455
rect 1710 -2495 1720 -2455
rect 1660 -2515 1720 -2495
rect 1660 -2555 1670 -2515
rect 1710 -2555 1720 -2515
rect 1660 -2580 1720 -2555
rect 1660 -2620 1670 -2580
rect 1710 -2620 1720 -2580
rect 1660 -2650 1720 -2620
rect 1660 -2690 1670 -2650
rect 1710 -2690 1720 -2650
rect 1660 -2720 1720 -2690
rect 1660 -2760 1670 -2720
rect 1710 -2760 1720 -2720
rect 1660 -2790 1720 -2760
rect 1660 -2830 1670 -2790
rect 1710 -2830 1720 -2790
rect 1660 -2855 1720 -2830
rect 1660 -2895 1670 -2855
rect 1710 -2895 1720 -2855
rect 1660 -2905 1720 -2895
rect 2010 -1315 2070 -1305
rect 2010 -1355 2020 -1315
rect 2060 -1355 2070 -1315
rect 2010 -1380 2070 -1355
rect 2010 -1420 2020 -1380
rect 2060 -1420 2070 -1380
rect 2010 -1450 2070 -1420
rect 2010 -1490 2020 -1450
rect 2060 -1490 2070 -1450
rect 2010 -1520 2070 -1490
rect 2010 -1560 2020 -1520
rect 2060 -1560 2070 -1520
rect 2010 -1590 2070 -1560
rect 2010 -1630 2020 -1590
rect 2060 -1630 2070 -1590
rect 2010 -1655 2070 -1630
rect 2010 -1695 2020 -1655
rect 2060 -1695 2070 -1655
rect 2010 -1715 2070 -1695
rect 2010 -1755 2020 -1715
rect 2060 -1755 2070 -1715
rect 2010 -1780 2070 -1755
rect 2010 -1820 2020 -1780
rect 2060 -1820 2070 -1780
rect 2010 -1850 2070 -1820
rect 2010 -1890 2020 -1850
rect 2060 -1890 2070 -1850
rect 2010 -1920 2070 -1890
rect 2010 -1960 2020 -1920
rect 2060 -1960 2070 -1920
rect 2010 -1990 2070 -1960
rect 2010 -2030 2020 -1990
rect 2060 -2030 2070 -1990
rect 2010 -2055 2070 -2030
rect 2010 -2095 2020 -2055
rect 2060 -2095 2070 -2055
rect 2010 -2115 2070 -2095
rect 2010 -2155 2020 -2115
rect 2060 -2155 2070 -2115
rect 2010 -2180 2070 -2155
rect 2010 -2220 2020 -2180
rect 2060 -2220 2070 -2180
rect 2010 -2250 2070 -2220
rect 2010 -2290 2020 -2250
rect 2060 -2290 2070 -2250
rect 2010 -2320 2070 -2290
rect 2010 -2360 2020 -2320
rect 2060 -2360 2070 -2320
rect 2010 -2390 2070 -2360
rect 2010 -2430 2020 -2390
rect 2060 -2430 2070 -2390
rect 2010 -2455 2070 -2430
rect 2010 -2495 2020 -2455
rect 2060 -2495 2070 -2455
rect 2010 -2515 2070 -2495
rect 2010 -2555 2020 -2515
rect 2060 -2555 2070 -2515
rect 2010 -2580 2070 -2555
rect 2010 -2620 2020 -2580
rect 2060 -2620 2070 -2580
rect 2010 -2650 2070 -2620
rect 2010 -2690 2020 -2650
rect 2060 -2690 2070 -2650
rect 2010 -2720 2070 -2690
rect 2010 -2760 2020 -2720
rect 2060 -2760 2070 -2720
rect 2010 -2790 2070 -2760
rect 2010 -2830 2020 -2790
rect 2060 -2830 2070 -2790
rect 2010 -2855 2070 -2830
rect 2010 -2895 2020 -2855
rect 2060 -2895 2070 -2855
rect 2010 -2905 2070 -2895
rect 2360 -1315 2420 -1305
rect 2360 -1355 2370 -1315
rect 2410 -1355 2420 -1315
rect 2360 -1380 2420 -1355
rect 2360 -1420 2370 -1380
rect 2410 -1420 2420 -1380
rect 2360 -1450 2420 -1420
rect 2360 -1490 2370 -1450
rect 2410 -1490 2420 -1450
rect 2360 -1520 2420 -1490
rect 2360 -1560 2370 -1520
rect 2410 -1560 2420 -1520
rect 2360 -1590 2420 -1560
rect 2360 -1630 2370 -1590
rect 2410 -1630 2420 -1590
rect 2360 -1655 2420 -1630
rect 2360 -1695 2370 -1655
rect 2410 -1695 2420 -1655
rect 2360 -1715 2420 -1695
rect 2360 -1755 2370 -1715
rect 2410 -1755 2420 -1715
rect 2360 -1780 2420 -1755
rect 2360 -1820 2370 -1780
rect 2410 -1820 2420 -1780
rect 2360 -1850 2420 -1820
rect 2360 -1890 2370 -1850
rect 2410 -1890 2420 -1850
rect 2360 -1920 2420 -1890
rect 2360 -1960 2370 -1920
rect 2410 -1960 2420 -1920
rect 2360 -1990 2420 -1960
rect 2360 -2030 2370 -1990
rect 2410 -2030 2420 -1990
rect 2360 -2055 2420 -2030
rect 2360 -2095 2370 -2055
rect 2410 -2095 2420 -2055
rect 2360 -2115 2420 -2095
rect 2360 -2155 2370 -2115
rect 2410 -2155 2420 -2115
rect 2360 -2180 2420 -2155
rect 2360 -2220 2370 -2180
rect 2410 -2220 2420 -2180
rect 2360 -2250 2420 -2220
rect 2360 -2290 2370 -2250
rect 2410 -2290 2420 -2250
rect 2360 -2320 2420 -2290
rect 2360 -2360 2370 -2320
rect 2410 -2360 2420 -2320
rect 2360 -2390 2420 -2360
rect 2360 -2430 2370 -2390
rect 2410 -2430 2420 -2390
rect 2360 -2455 2420 -2430
rect 2360 -2495 2370 -2455
rect 2410 -2495 2420 -2455
rect 2360 -2515 2420 -2495
rect 2360 -2555 2370 -2515
rect 2410 -2555 2420 -2515
rect 2360 -2580 2420 -2555
rect 2360 -2620 2370 -2580
rect 2410 -2620 2420 -2580
rect 2360 -2650 2420 -2620
rect 2360 -2690 2370 -2650
rect 2410 -2690 2420 -2650
rect 2360 -2720 2420 -2690
rect 2360 -2760 2370 -2720
rect 2410 -2760 2420 -2720
rect 2360 -2790 2420 -2760
rect 2360 -2830 2370 -2790
rect 2410 -2830 2420 -2790
rect 2360 -2855 2420 -2830
rect 2360 -2895 2370 -2855
rect 2410 -2895 2420 -2855
rect 2360 -2905 2420 -2895
rect 2710 -1315 2770 -1305
rect 2710 -1355 2720 -1315
rect 2760 -1355 2770 -1315
rect 2710 -1380 2770 -1355
rect 2710 -1420 2720 -1380
rect 2760 -1420 2770 -1380
rect 2710 -1450 2770 -1420
rect 2710 -1490 2720 -1450
rect 2760 -1490 2770 -1450
rect 2710 -1520 2770 -1490
rect 2710 -1560 2720 -1520
rect 2760 -1560 2770 -1520
rect 2710 -1590 2770 -1560
rect 2710 -1630 2720 -1590
rect 2760 -1630 2770 -1590
rect 2710 -1655 2770 -1630
rect 2710 -1695 2720 -1655
rect 2760 -1695 2770 -1655
rect 2710 -1715 2770 -1695
rect 2710 -1755 2720 -1715
rect 2760 -1755 2770 -1715
rect 2710 -1780 2770 -1755
rect 2710 -1820 2720 -1780
rect 2760 -1820 2770 -1780
rect 2710 -1850 2770 -1820
rect 2710 -1890 2720 -1850
rect 2760 -1890 2770 -1850
rect 2710 -1920 2770 -1890
rect 2710 -1960 2720 -1920
rect 2760 -1960 2770 -1920
rect 2710 -1990 2770 -1960
rect 2710 -2030 2720 -1990
rect 2760 -2030 2770 -1990
rect 2710 -2055 2770 -2030
rect 2710 -2095 2720 -2055
rect 2760 -2095 2770 -2055
rect 2710 -2115 2770 -2095
rect 2710 -2155 2720 -2115
rect 2760 -2155 2770 -2115
rect 2710 -2180 2770 -2155
rect 2710 -2220 2720 -2180
rect 2760 -2220 2770 -2180
rect 2710 -2250 2770 -2220
rect 2710 -2290 2720 -2250
rect 2760 -2290 2770 -2250
rect 2710 -2320 2770 -2290
rect 2710 -2360 2720 -2320
rect 2760 -2360 2770 -2320
rect 2710 -2390 2770 -2360
rect 2710 -2430 2720 -2390
rect 2760 -2430 2770 -2390
rect 2710 -2455 2770 -2430
rect 2710 -2495 2720 -2455
rect 2760 -2495 2770 -2455
rect 2710 -2515 2770 -2495
rect 2710 -2555 2720 -2515
rect 2760 -2555 2770 -2515
rect 2710 -2580 2770 -2555
rect 2710 -2620 2720 -2580
rect 2760 -2620 2770 -2580
rect 2710 -2650 2770 -2620
rect 2710 -2690 2720 -2650
rect 2760 -2690 2770 -2650
rect 2710 -2720 2770 -2690
rect 2710 -2760 2720 -2720
rect 2760 -2760 2770 -2720
rect 2710 -2790 2770 -2760
rect 2710 -2830 2720 -2790
rect 2760 -2830 2770 -2790
rect 2710 -2855 2770 -2830
rect 2710 -2895 2720 -2855
rect 2760 -2895 2770 -2855
rect 2710 -2905 2770 -2895
rect 3060 -1315 3120 -1305
rect 3060 -1355 3070 -1315
rect 3110 -1355 3120 -1315
rect 3060 -1380 3120 -1355
rect 3060 -1420 3070 -1380
rect 3110 -1420 3120 -1380
rect 3060 -1450 3120 -1420
rect 3060 -1490 3070 -1450
rect 3110 -1490 3120 -1450
rect 3060 -1520 3120 -1490
rect 3060 -1560 3070 -1520
rect 3110 -1560 3120 -1520
rect 3060 -1590 3120 -1560
rect 3060 -1630 3070 -1590
rect 3110 -1630 3120 -1590
rect 3060 -1655 3120 -1630
rect 3060 -1695 3070 -1655
rect 3110 -1695 3120 -1655
rect 3060 -1715 3120 -1695
rect 3060 -1755 3070 -1715
rect 3110 -1755 3120 -1715
rect 3060 -1780 3120 -1755
rect 3060 -1820 3070 -1780
rect 3110 -1820 3120 -1780
rect 3060 -1850 3120 -1820
rect 3060 -1890 3070 -1850
rect 3110 -1890 3120 -1850
rect 3060 -1920 3120 -1890
rect 3060 -1960 3070 -1920
rect 3110 -1960 3120 -1920
rect 3060 -1990 3120 -1960
rect 3060 -2030 3070 -1990
rect 3110 -2030 3120 -1990
rect 3060 -2055 3120 -2030
rect 3060 -2095 3070 -2055
rect 3110 -2095 3120 -2055
rect 3060 -2115 3120 -2095
rect 3060 -2155 3070 -2115
rect 3110 -2155 3120 -2115
rect 3060 -2180 3120 -2155
rect 3060 -2220 3070 -2180
rect 3110 -2220 3120 -2180
rect 3060 -2250 3120 -2220
rect 3060 -2290 3070 -2250
rect 3110 -2290 3120 -2250
rect 3060 -2320 3120 -2290
rect 3060 -2360 3070 -2320
rect 3110 -2360 3120 -2320
rect 3060 -2390 3120 -2360
rect 3060 -2430 3070 -2390
rect 3110 -2430 3120 -2390
rect 3060 -2455 3120 -2430
rect 3060 -2495 3070 -2455
rect 3110 -2495 3120 -2455
rect 3060 -2515 3120 -2495
rect 3060 -2555 3070 -2515
rect 3110 -2555 3120 -2515
rect 3060 -2580 3120 -2555
rect 3060 -2620 3070 -2580
rect 3110 -2620 3120 -2580
rect 3060 -2650 3120 -2620
rect 3060 -2690 3070 -2650
rect 3110 -2690 3120 -2650
rect 3060 -2720 3120 -2690
rect 3060 -2760 3070 -2720
rect 3110 -2760 3120 -2720
rect 3060 -2790 3120 -2760
rect 3060 -2830 3070 -2790
rect 3110 -2830 3120 -2790
rect 3060 -2855 3120 -2830
rect 3060 -2895 3070 -2855
rect 3110 -2895 3120 -2855
rect 3060 -2905 3120 -2895
rect 5860 -1315 5920 -1305
rect 5860 -1355 5870 -1315
rect 5910 -1355 5920 -1315
rect 5860 -1380 5920 -1355
rect 5860 -1420 5870 -1380
rect 5910 -1420 5920 -1380
rect 5860 -1450 5920 -1420
rect 5860 -1490 5870 -1450
rect 5910 -1490 5920 -1450
rect 5860 -1520 5920 -1490
rect 5860 -1560 5870 -1520
rect 5910 -1560 5920 -1520
rect 5860 -1590 5920 -1560
rect 5860 -1630 5870 -1590
rect 5910 -1630 5920 -1590
rect 5860 -1655 5920 -1630
rect 5860 -1695 5870 -1655
rect 5910 -1695 5920 -1655
rect 5860 -1715 5920 -1695
rect 5860 -1755 5870 -1715
rect 5910 -1755 5920 -1715
rect 5860 -1780 5920 -1755
rect 5860 -1820 5870 -1780
rect 5910 -1820 5920 -1780
rect 5860 -1850 5920 -1820
rect 5860 -1890 5870 -1850
rect 5910 -1890 5920 -1850
rect 5860 -1920 5920 -1890
rect 5860 -1960 5870 -1920
rect 5910 -1960 5920 -1920
rect 5860 -1990 5920 -1960
rect 5860 -2030 5870 -1990
rect 5910 -2030 5920 -1990
rect 5860 -2055 5920 -2030
rect 5860 -2095 5870 -2055
rect 5910 -2095 5920 -2055
rect 5860 -2115 5920 -2095
rect 5860 -2155 5870 -2115
rect 5910 -2155 5920 -2115
rect 5860 -2180 5920 -2155
rect 5860 -2220 5870 -2180
rect 5910 -2220 5920 -2180
rect 5860 -2250 5920 -2220
rect 5860 -2290 5870 -2250
rect 5910 -2290 5920 -2250
rect 5860 -2320 5920 -2290
rect 5860 -2360 5870 -2320
rect 5910 -2360 5920 -2320
rect 5860 -2390 5920 -2360
rect 5860 -2430 5870 -2390
rect 5910 -2430 5920 -2390
rect 5860 -2455 5920 -2430
rect 5860 -2495 5870 -2455
rect 5910 -2495 5920 -2455
rect 5860 -2515 5920 -2495
rect 5860 -2555 5870 -2515
rect 5910 -2555 5920 -2515
rect 5860 -2580 5920 -2555
rect 5860 -2620 5870 -2580
rect 5910 -2620 5920 -2580
rect 5860 -2650 5920 -2620
rect 5860 -2690 5870 -2650
rect 5910 -2690 5920 -2650
rect 5860 -2720 5920 -2690
rect 5860 -2760 5870 -2720
rect 5910 -2760 5920 -2720
rect 5860 -2790 5920 -2760
rect 5860 -2830 5870 -2790
rect 5910 -2830 5920 -2790
rect 5860 -2855 5920 -2830
rect 5860 -2895 5870 -2855
rect 5910 -2895 5920 -2855
rect 5860 -2905 5920 -2895
rect 6210 -1315 6270 -1305
rect 6210 -1355 6220 -1315
rect 6260 -1355 6270 -1315
rect 6210 -1380 6270 -1355
rect 6210 -1420 6220 -1380
rect 6260 -1420 6270 -1380
rect 6210 -1450 6270 -1420
rect 6210 -1490 6220 -1450
rect 6260 -1490 6270 -1450
rect 6210 -1520 6270 -1490
rect 6210 -1560 6220 -1520
rect 6260 -1560 6270 -1520
rect 6210 -1590 6270 -1560
rect 6210 -1630 6220 -1590
rect 6260 -1630 6270 -1590
rect 6210 -1655 6270 -1630
rect 6210 -1695 6220 -1655
rect 6260 -1695 6270 -1655
rect 6210 -1715 6270 -1695
rect 6210 -1755 6220 -1715
rect 6260 -1755 6270 -1715
rect 6210 -1780 6270 -1755
rect 6210 -1820 6220 -1780
rect 6260 -1820 6270 -1780
rect 6210 -1850 6270 -1820
rect 6210 -1890 6220 -1850
rect 6260 -1890 6270 -1850
rect 6210 -1920 6270 -1890
rect 6210 -1960 6220 -1920
rect 6260 -1960 6270 -1920
rect 6210 -1990 6270 -1960
rect 6210 -2030 6220 -1990
rect 6260 -2030 6270 -1990
rect 6210 -2055 6270 -2030
rect 6210 -2095 6220 -2055
rect 6260 -2095 6270 -2055
rect 6210 -2115 6270 -2095
rect 6210 -2155 6220 -2115
rect 6260 -2155 6270 -2115
rect 6210 -2180 6270 -2155
rect 6210 -2220 6220 -2180
rect 6260 -2220 6270 -2180
rect 6210 -2250 6270 -2220
rect 6210 -2290 6220 -2250
rect 6260 -2290 6270 -2250
rect 6210 -2320 6270 -2290
rect 6210 -2360 6220 -2320
rect 6260 -2360 6270 -2320
rect 6210 -2390 6270 -2360
rect 6210 -2430 6220 -2390
rect 6260 -2430 6270 -2390
rect 6210 -2455 6270 -2430
rect 6210 -2495 6220 -2455
rect 6260 -2495 6270 -2455
rect 6210 -2515 6270 -2495
rect 6210 -2555 6220 -2515
rect 6260 -2555 6270 -2515
rect 6210 -2580 6270 -2555
rect 6210 -2620 6220 -2580
rect 6260 -2620 6270 -2580
rect 6210 -2650 6270 -2620
rect 6210 -2690 6220 -2650
rect 6260 -2690 6270 -2650
rect 6210 -2720 6270 -2690
rect 6210 -2760 6220 -2720
rect 6260 -2760 6270 -2720
rect 6210 -2790 6270 -2760
rect 6210 -2830 6220 -2790
rect 6260 -2830 6270 -2790
rect 6210 -2855 6270 -2830
rect 6210 -2895 6220 -2855
rect 6260 -2895 6270 -2855
rect 6210 -2905 6270 -2895
rect 6560 -1315 6620 -1305
rect 6560 -1355 6570 -1315
rect 6610 -1355 6620 -1315
rect 6560 -1380 6620 -1355
rect 6560 -1420 6570 -1380
rect 6610 -1420 6620 -1380
rect 6560 -1450 6620 -1420
rect 6560 -1490 6570 -1450
rect 6610 -1490 6620 -1450
rect 6560 -1520 6620 -1490
rect 6560 -1560 6570 -1520
rect 6610 -1560 6620 -1520
rect 6560 -1590 6620 -1560
rect 6560 -1630 6570 -1590
rect 6610 -1630 6620 -1590
rect 6560 -1655 6620 -1630
rect 6560 -1695 6570 -1655
rect 6610 -1695 6620 -1655
rect 6560 -1715 6620 -1695
rect 6560 -1755 6570 -1715
rect 6610 -1755 6620 -1715
rect 6560 -1780 6620 -1755
rect 6560 -1820 6570 -1780
rect 6610 -1820 6620 -1780
rect 6560 -1850 6620 -1820
rect 6560 -1890 6570 -1850
rect 6610 -1890 6620 -1850
rect 6560 -1920 6620 -1890
rect 6560 -1960 6570 -1920
rect 6610 -1960 6620 -1920
rect 6560 -1990 6620 -1960
rect 6560 -2030 6570 -1990
rect 6610 -2030 6620 -1990
rect 6560 -2055 6620 -2030
rect 6560 -2095 6570 -2055
rect 6610 -2095 6620 -2055
rect 6560 -2115 6620 -2095
rect 6560 -2155 6570 -2115
rect 6610 -2155 6620 -2115
rect 6560 -2180 6620 -2155
rect 6560 -2220 6570 -2180
rect 6610 -2220 6620 -2180
rect 6560 -2250 6620 -2220
rect 6560 -2290 6570 -2250
rect 6610 -2290 6620 -2250
rect 6560 -2320 6620 -2290
rect 6560 -2360 6570 -2320
rect 6610 -2360 6620 -2320
rect 6560 -2390 6620 -2360
rect 6560 -2430 6570 -2390
rect 6610 -2430 6620 -2390
rect 6560 -2455 6620 -2430
rect 6560 -2495 6570 -2455
rect 6610 -2495 6620 -2455
rect 6560 -2515 6620 -2495
rect 6560 -2555 6570 -2515
rect 6610 -2555 6620 -2515
rect 6560 -2580 6620 -2555
rect 6560 -2620 6570 -2580
rect 6610 -2620 6620 -2580
rect 6560 -2650 6620 -2620
rect 6560 -2690 6570 -2650
rect 6610 -2690 6620 -2650
rect 6560 -2720 6620 -2690
rect 6560 -2760 6570 -2720
rect 6610 -2760 6620 -2720
rect 6560 -2790 6620 -2760
rect 6560 -2830 6570 -2790
rect 6610 -2830 6620 -2790
rect 6560 -2855 6620 -2830
rect 6560 -2895 6570 -2855
rect 6610 -2895 6620 -2855
rect 6560 -2905 6620 -2895
rect 6910 -1315 6970 -1305
rect 6910 -1355 6920 -1315
rect 6960 -1355 6970 -1315
rect 6910 -1380 6970 -1355
rect 6910 -1420 6920 -1380
rect 6960 -1420 6970 -1380
rect 6910 -1450 6970 -1420
rect 6910 -1490 6920 -1450
rect 6960 -1490 6970 -1450
rect 6910 -1520 6970 -1490
rect 6910 -1560 6920 -1520
rect 6960 -1560 6970 -1520
rect 6910 -1590 6970 -1560
rect 6910 -1630 6920 -1590
rect 6960 -1630 6970 -1590
rect 6910 -1655 6970 -1630
rect 6910 -1695 6920 -1655
rect 6960 -1695 6970 -1655
rect 6910 -1715 6970 -1695
rect 6910 -1755 6920 -1715
rect 6960 -1755 6970 -1715
rect 6910 -1780 6970 -1755
rect 6910 -1820 6920 -1780
rect 6960 -1820 6970 -1780
rect 6910 -1850 6970 -1820
rect 6910 -1890 6920 -1850
rect 6960 -1890 6970 -1850
rect 6910 -1920 6970 -1890
rect 6910 -1960 6920 -1920
rect 6960 -1960 6970 -1920
rect 6910 -1990 6970 -1960
rect 6910 -2030 6920 -1990
rect 6960 -2030 6970 -1990
rect 6910 -2055 6970 -2030
rect 6910 -2095 6920 -2055
rect 6960 -2095 6970 -2055
rect 6910 -2115 6970 -2095
rect 6910 -2155 6920 -2115
rect 6960 -2155 6970 -2115
rect 6910 -2180 6970 -2155
rect 6910 -2220 6920 -2180
rect 6960 -2220 6970 -2180
rect 6910 -2250 6970 -2220
rect 6910 -2290 6920 -2250
rect 6960 -2290 6970 -2250
rect 6910 -2320 6970 -2290
rect 6910 -2360 6920 -2320
rect 6960 -2360 6970 -2320
rect 6910 -2390 6970 -2360
rect 6910 -2430 6920 -2390
rect 6960 -2430 6970 -2390
rect 6910 -2455 6970 -2430
rect 6910 -2495 6920 -2455
rect 6960 -2495 6970 -2455
rect 6910 -2515 6970 -2495
rect 6910 -2555 6920 -2515
rect 6960 -2555 6970 -2515
rect 6910 -2580 6970 -2555
rect 6910 -2620 6920 -2580
rect 6960 -2620 6970 -2580
rect 6910 -2650 6970 -2620
rect 6910 -2690 6920 -2650
rect 6960 -2690 6970 -2650
rect 6910 -2720 6970 -2690
rect 6910 -2760 6920 -2720
rect 6960 -2760 6970 -2720
rect 6910 -2790 6970 -2760
rect 6910 -2830 6920 -2790
rect 6960 -2830 6970 -2790
rect 6910 -2855 6970 -2830
rect 6910 -2895 6920 -2855
rect 6960 -2895 6970 -2855
rect 6910 -2905 6970 -2895
rect 7260 -1315 7320 -1305
rect 7260 -1355 7270 -1315
rect 7310 -1355 7320 -1315
rect 7260 -1380 7320 -1355
rect 7260 -1420 7270 -1380
rect 7310 -1420 7320 -1380
rect 7260 -1450 7320 -1420
rect 7260 -1490 7270 -1450
rect 7310 -1490 7320 -1450
rect 7260 -1520 7320 -1490
rect 7260 -1560 7270 -1520
rect 7310 -1560 7320 -1520
rect 7260 -1590 7320 -1560
rect 7260 -1630 7270 -1590
rect 7310 -1630 7320 -1590
rect 7260 -1655 7320 -1630
rect 7260 -1695 7270 -1655
rect 7310 -1695 7320 -1655
rect 7260 -1715 7320 -1695
rect 7260 -1755 7270 -1715
rect 7310 -1755 7320 -1715
rect 7260 -1780 7320 -1755
rect 7260 -1820 7270 -1780
rect 7310 -1820 7320 -1780
rect 7260 -1850 7320 -1820
rect 7260 -1890 7270 -1850
rect 7310 -1890 7320 -1850
rect 7260 -1920 7320 -1890
rect 7260 -1960 7270 -1920
rect 7310 -1960 7320 -1920
rect 7260 -1990 7320 -1960
rect 7260 -2030 7270 -1990
rect 7310 -2030 7320 -1990
rect 7260 -2055 7320 -2030
rect 7260 -2095 7270 -2055
rect 7310 -2095 7320 -2055
rect 7260 -2115 7320 -2095
rect 7260 -2155 7270 -2115
rect 7310 -2155 7320 -2115
rect 7260 -2180 7320 -2155
rect 7260 -2220 7270 -2180
rect 7310 -2220 7320 -2180
rect 7260 -2250 7320 -2220
rect 7260 -2290 7270 -2250
rect 7310 -2290 7320 -2250
rect 7260 -2320 7320 -2290
rect 7260 -2360 7270 -2320
rect 7310 -2360 7320 -2320
rect 7260 -2390 7320 -2360
rect 7260 -2430 7270 -2390
rect 7310 -2430 7320 -2390
rect 7260 -2455 7320 -2430
rect 7260 -2495 7270 -2455
rect 7310 -2495 7320 -2455
rect 7260 -2515 7320 -2495
rect 7260 -2555 7270 -2515
rect 7310 -2555 7320 -2515
rect 7260 -2580 7320 -2555
rect 7260 -2620 7270 -2580
rect 7310 -2620 7320 -2580
rect 7260 -2650 7320 -2620
rect 7260 -2690 7270 -2650
rect 7310 -2690 7320 -2650
rect 7260 -2720 7320 -2690
rect 7260 -2760 7270 -2720
rect 7310 -2760 7320 -2720
rect 7260 -2790 7320 -2760
rect 7260 -2830 7270 -2790
rect 7310 -2830 7320 -2790
rect 7260 -2855 7320 -2830
rect 7260 -2895 7270 -2855
rect 7310 -2895 7320 -2855
rect 7260 -2905 7320 -2895
rect 7610 -1315 7670 -1305
rect 7610 -1355 7620 -1315
rect 7660 -1355 7670 -1315
rect 7610 -1380 7670 -1355
rect 7610 -1420 7620 -1380
rect 7660 -1420 7670 -1380
rect 7610 -1450 7670 -1420
rect 7610 -1490 7620 -1450
rect 7660 -1490 7670 -1450
rect 7610 -1520 7670 -1490
rect 7610 -1560 7620 -1520
rect 7660 -1560 7670 -1520
rect 7610 -1590 7670 -1560
rect 7610 -1630 7620 -1590
rect 7660 -1630 7670 -1590
rect 7610 -1655 7670 -1630
rect 7610 -1695 7620 -1655
rect 7660 -1695 7670 -1655
rect 7610 -1715 7670 -1695
rect 7610 -1755 7620 -1715
rect 7660 -1755 7670 -1715
rect 7610 -1780 7670 -1755
rect 7610 -1820 7620 -1780
rect 7660 -1820 7670 -1780
rect 7610 -1850 7670 -1820
rect 7610 -1890 7620 -1850
rect 7660 -1890 7670 -1850
rect 7610 -1920 7670 -1890
rect 7610 -1960 7620 -1920
rect 7660 -1960 7670 -1920
rect 7610 -1990 7670 -1960
rect 7610 -2030 7620 -1990
rect 7660 -2030 7670 -1990
rect 7610 -2055 7670 -2030
rect 7610 -2095 7620 -2055
rect 7660 -2095 7670 -2055
rect 7610 -2115 7670 -2095
rect 7610 -2155 7620 -2115
rect 7660 -2155 7670 -2115
rect 7610 -2180 7670 -2155
rect 7610 -2220 7620 -2180
rect 7660 -2220 7670 -2180
rect 7610 -2250 7670 -2220
rect 7610 -2290 7620 -2250
rect 7660 -2290 7670 -2250
rect 7610 -2320 7670 -2290
rect 7610 -2360 7620 -2320
rect 7660 -2360 7670 -2320
rect 7610 -2390 7670 -2360
rect 7610 -2430 7620 -2390
rect 7660 -2430 7670 -2390
rect 7610 -2455 7670 -2430
rect 7610 -2495 7620 -2455
rect 7660 -2495 7670 -2455
rect 7610 -2515 7670 -2495
rect 7610 -2555 7620 -2515
rect 7660 -2555 7670 -2515
rect 7610 -2580 7670 -2555
rect 7610 -2620 7620 -2580
rect 7660 -2620 7670 -2580
rect 7610 -2650 7670 -2620
rect 7610 -2690 7620 -2650
rect 7660 -2690 7670 -2650
rect 7610 -2720 7670 -2690
rect 7610 -2760 7620 -2720
rect 7660 -2760 7670 -2720
rect 7610 -2790 7670 -2760
rect 7610 -2830 7620 -2790
rect 7660 -2830 7670 -2790
rect 7610 -2855 7670 -2830
rect 7610 -2895 7620 -2855
rect 7660 -2895 7670 -2855
rect 7610 -2905 7670 -2895
rect 7960 -1315 8020 -1305
rect 7960 -1355 7970 -1315
rect 8010 -1355 8020 -1315
rect 7960 -1380 8020 -1355
rect 7960 -1420 7970 -1380
rect 8010 -1420 8020 -1380
rect 7960 -1450 8020 -1420
rect 7960 -1490 7970 -1450
rect 8010 -1490 8020 -1450
rect 7960 -1520 8020 -1490
rect 7960 -1560 7970 -1520
rect 8010 -1560 8020 -1520
rect 7960 -1590 8020 -1560
rect 7960 -1630 7970 -1590
rect 8010 -1630 8020 -1590
rect 7960 -1655 8020 -1630
rect 7960 -1695 7970 -1655
rect 8010 -1695 8020 -1655
rect 7960 -1715 8020 -1695
rect 7960 -1755 7970 -1715
rect 8010 -1755 8020 -1715
rect 7960 -1780 8020 -1755
rect 7960 -1820 7970 -1780
rect 8010 -1820 8020 -1780
rect 7960 -1850 8020 -1820
rect 7960 -1890 7970 -1850
rect 8010 -1890 8020 -1850
rect 7960 -1920 8020 -1890
rect 7960 -1960 7970 -1920
rect 8010 -1960 8020 -1920
rect 7960 -1990 8020 -1960
rect 7960 -2030 7970 -1990
rect 8010 -2030 8020 -1990
rect 7960 -2055 8020 -2030
rect 7960 -2095 7970 -2055
rect 8010 -2095 8020 -2055
rect 7960 -2115 8020 -2095
rect 7960 -2155 7970 -2115
rect 8010 -2155 8020 -2115
rect 7960 -2180 8020 -2155
rect 7960 -2220 7970 -2180
rect 8010 -2220 8020 -2180
rect 7960 -2250 8020 -2220
rect 7960 -2290 7970 -2250
rect 8010 -2290 8020 -2250
rect 7960 -2320 8020 -2290
rect 7960 -2360 7970 -2320
rect 8010 -2360 8020 -2320
rect 7960 -2390 8020 -2360
rect 7960 -2430 7970 -2390
rect 8010 -2430 8020 -2390
rect 7960 -2455 8020 -2430
rect 7960 -2495 7970 -2455
rect 8010 -2495 8020 -2455
rect 7960 -2515 8020 -2495
rect 7960 -2555 7970 -2515
rect 8010 -2555 8020 -2515
rect 7960 -2580 8020 -2555
rect 7960 -2620 7970 -2580
rect 8010 -2620 8020 -2580
rect 7960 -2650 8020 -2620
rect 7960 -2690 7970 -2650
rect 8010 -2690 8020 -2650
rect 7960 -2720 8020 -2690
rect 7960 -2760 7970 -2720
rect 8010 -2760 8020 -2720
rect 7960 -2790 8020 -2760
rect 7960 -2830 7970 -2790
rect 8010 -2830 8020 -2790
rect 7960 -2855 8020 -2830
rect 7960 -2895 7970 -2855
rect 8010 -2895 8020 -2855
rect 7960 -2905 8020 -2895
rect 8310 -1315 8370 -1305
rect 8310 -1355 8320 -1315
rect 8360 -1355 8370 -1315
rect 8310 -1380 8370 -1355
rect 8310 -1420 8320 -1380
rect 8360 -1420 8370 -1380
rect 8310 -1450 8370 -1420
rect 8310 -1490 8320 -1450
rect 8360 -1490 8370 -1450
rect 8310 -1520 8370 -1490
rect 8310 -1560 8320 -1520
rect 8360 -1560 8370 -1520
rect 8310 -1590 8370 -1560
rect 8310 -1630 8320 -1590
rect 8360 -1630 8370 -1590
rect 8310 -1655 8370 -1630
rect 8310 -1695 8320 -1655
rect 8360 -1695 8370 -1655
rect 8310 -1715 8370 -1695
rect 8310 -1755 8320 -1715
rect 8360 -1755 8370 -1715
rect 8310 -1780 8370 -1755
rect 8310 -1820 8320 -1780
rect 8360 -1820 8370 -1780
rect 8310 -1850 8370 -1820
rect 8310 -1890 8320 -1850
rect 8360 -1890 8370 -1850
rect 8310 -1920 8370 -1890
rect 8310 -1960 8320 -1920
rect 8360 -1960 8370 -1920
rect 8310 -1990 8370 -1960
rect 8310 -2030 8320 -1990
rect 8360 -2030 8370 -1990
rect 8310 -2055 8370 -2030
rect 8310 -2095 8320 -2055
rect 8360 -2095 8370 -2055
rect 8310 -2115 8370 -2095
rect 8310 -2155 8320 -2115
rect 8360 -2155 8370 -2115
rect 8310 -2180 8370 -2155
rect 8310 -2220 8320 -2180
rect 8360 -2220 8370 -2180
rect 8310 -2250 8370 -2220
rect 8310 -2290 8320 -2250
rect 8360 -2290 8370 -2250
rect 8310 -2320 8370 -2290
rect 8310 -2360 8320 -2320
rect 8360 -2360 8370 -2320
rect 8310 -2390 8370 -2360
rect 8310 -2430 8320 -2390
rect 8360 -2430 8370 -2390
rect 8310 -2455 8370 -2430
rect 8310 -2495 8320 -2455
rect 8360 -2495 8370 -2455
rect 8310 -2515 8370 -2495
rect 8310 -2555 8320 -2515
rect 8360 -2555 8370 -2515
rect 8310 -2580 8370 -2555
rect 8310 -2620 8320 -2580
rect 8360 -2620 8370 -2580
rect 8310 -2650 8370 -2620
rect 8310 -2690 8320 -2650
rect 8360 -2690 8370 -2650
rect 8310 -2720 8370 -2690
rect 8310 -2760 8320 -2720
rect 8360 -2760 8370 -2720
rect 8310 -2790 8370 -2760
rect 8310 -2830 8320 -2790
rect 8360 -2830 8370 -2790
rect 8310 -2855 8370 -2830
rect 8310 -2895 8320 -2855
rect 8360 -2895 8370 -2855
rect 8310 -2905 8370 -2895
rect 8660 -1315 8720 -1305
rect 8660 -1355 8670 -1315
rect 8710 -1355 8720 -1315
rect 8660 -1380 8720 -1355
rect 8660 -1420 8670 -1380
rect 8710 -1420 8720 -1380
rect 8660 -1450 8720 -1420
rect 8660 -1490 8670 -1450
rect 8710 -1490 8720 -1450
rect 8660 -1520 8720 -1490
rect 8660 -1560 8670 -1520
rect 8710 -1560 8720 -1520
rect 8660 -1590 8720 -1560
rect 8660 -1630 8670 -1590
rect 8710 -1630 8720 -1590
rect 8660 -1655 8720 -1630
rect 8660 -1695 8670 -1655
rect 8710 -1695 8720 -1655
rect 8660 -1715 8720 -1695
rect 8660 -1755 8670 -1715
rect 8710 -1755 8720 -1715
rect 8660 -1780 8720 -1755
rect 8660 -1820 8670 -1780
rect 8710 -1820 8720 -1780
rect 8660 -1850 8720 -1820
rect 8660 -1890 8670 -1850
rect 8710 -1890 8720 -1850
rect 8660 -1920 8720 -1890
rect 8660 -1960 8670 -1920
rect 8710 -1960 8720 -1920
rect 8660 -1990 8720 -1960
rect 8660 -2030 8670 -1990
rect 8710 -2030 8720 -1990
rect 8660 -2055 8720 -2030
rect 8660 -2095 8670 -2055
rect 8710 -2095 8720 -2055
rect 8660 -2115 8720 -2095
rect 8660 -2155 8670 -2115
rect 8710 -2155 8720 -2115
rect 8660 -2180 8720 -2155
rect 8660 -2220 8670 -2180
rect 8710 -2220 8720 -2180
rect 8660 -2250 8720 -2220
rect 8660 -2290 8670 -2250
rect 8710 -2290 8720 -2250
rect 8660 -2320 8720 -2290
rect 8660 -2360 8670 -2320
rect 8710 -2360 8720 -2320
rect 8660 -2390 8720 -2360
rect 8660 -2430 8670 -2390
rect 8710 -2430 8720 -2390
rect 8660 -2455 8720 -2430
rect 8660 -2495 8670 -2455
rect 8710 -2495 8720 -2455
rect 8660 -2515 8720 -2495
rect 8660 -2555 8670 -2515
rect 8710 -2555 8720 -2515
rect 8660 -2580 8720 -2555
rect 8660 -2620 8670 -2580
rect 8710 -2620 8720 -2580
rect 8660 -2650 8720 -2620
rect 8660 -2690 8670 -2650
rect 8710 -2690 8720 -2650
rect 8660 -2720 8720 -2690
rect 8660 -2760 8670 -2720
rect 8710 -2760 8720 -2720
rect 8660 -2790 8720 -2760
rect 8660 -2830 8670 -2790
rect 8710 -2830 8720 -2790
rect 8660 -2855 8720 -2830
rect 8660 -2895 8670 -2855
rect 8710 -2895 8720 -2855
rect 8660 -2905 8720 -2895
rect 9010 -1315 9070 -1305
rect 9010 -1355 9020 -1315
rect 9060 -1355 9070 -1315
rect 9010 -1380 9070 -1355
rect 9010 -1420 9020 -1380
rect 9060 -1420 9070 -1380
rect 9010 -1450 9070 -1420
rect 9010 -1490 9020 -1450
rect 9060 -1490 9070 -1450
rect 9010 -1520 9070 -1490
rect 9010 -1560 9020 -1520
rect 9060 -1560 9070 -1520
rect 9010 -1590 9070 -1560
rect 9010 -1630 9020 -1590
rect 9060 -1630 9070 -1590
rect 9010 -1655 9070 -1630
rect 9010 -1695 9020 -1655
rect 9060 -1695 9070 -1655
rect 9010 -1715 9070 -1695
rect 9010 -1755 9020 -1715
rect 9060 -1755 9070 -1715
rect 9010 -1780 9070 -1755
rect 9010 -1820 9020 -1780
rect 9060 -1820 9070 -1780
rect 9010 -1850 9070 -1820
rect 9010 -1890 9020 -1850
rect 9060 -1890 9070 -1850
rect 9010 -1920 9070 -1890
rect 9010 -1960 9020 -1920
rect 9060 -1960 9070 -1920
rect 9010 -1990 9070 -1960
rect 9010 -2030 9020 -1990
rect 9060 -2030 9070 -1990
rect 9010 -2055 9070 -2030
rect 9010 -2095 9020 -2055
rect 9060 -2095 9070 -2055
rect 9010 -2115 9070 -2095
rect 9010 -2155 9020 -2115
rect 9060 -2155 9070 -2115
rect 9010 -2180 9070 -2155
rect 9010 -2220 9020 -2180
rect 9060 -2220 9070 -2180
rect 9010 -2250 9070 -2220
rect 9010 -2290 9020 -2250
rect 9060 -2290 9070 -2250
rect 9010 -2320 9070 -2290
rect 9010 -2360 9020 -2320
rect 9060 -2360 9070 -2320
rect 9010 -2390 9070 -2360
rect 9010 -2430 9020 -2390
rect 9060 -2430 9070 -2390
rect 9010 -2455 9070 -2430
rect 9010 -2495 9020 -2455
rect 9060 -2495 9070 -2455
rect 9010 -2515 9070 -2495
rect 9010 -2555 9020 -2515
rect 9060 -2555 9070 -2515
rect 9010 -2580 9070 -2555
rect 9010 -2620 9020 -2580
rect 9060 -2620 9070 -2580
rect 9010 -2650 9070 -2620
rect 9010 -2690 9020 -2650
rect 9060 -2690 9070 -2650
rect 9010 -2720 9070 -2690
rect 9010 -2760 9020 -2720
rect 9060 -2760 9070 -2720
rect 9010 -2790 9070 -2760
rect 9010 -2830 9020 -2790
rect 9060 -2830 9070 -2790
rect 9010 -2855 9070 -2830
rect 9010 -2895 9020 -2855
rect 9060 -2895 9070 -2855
rect 9010 -2905 9070 -2895
rect 31290 -1325 32890 6465
rect 31290 -1360 31305 -1325
rect 31340 -1360 31350 -1325
rect 31385 -1360 31395 -1325
rect 31430 -1360 31440 -1325
rect 31475 -1360 31485 -1325
rect 31520 -1360 31530 -1325
rect 31565 -1360 31575 -1325
rect 31610 -1360 31620 -1325
rect 31655 -1360 31665 -1325
rect 31700 -1360 31710 -1325
rect 31745 -1360 31755 -1325
rect 31790 -1360 31800 -1325
rect 31835 -1360 31845 -1325
rect 31880 -1360 31890 -1325
rect 31925 -1360 31935 -1325
rect 31970 -1360 31980 -1325
rect 32015 -1360 32025 -1325
rect 32060 -1360 32070 -1325
rect 32105 -1360 32115 -1325
rect 32150 -1360 32160 -1325
rect 32195 -1360 32205 -1325
rect 32240 -1360 32250 -1325
rect 32285 -1360 32295 -1325
rect 32330 -1360 32340 -1325
rect 32375 -1360 32385 -1325
rect 32420 -1360 32430 -1325
rect 32465 -1360 32475 -1325
rect 32510 -1360 32520 -1325
rect 32555 -1360 32565 -1325
rect 32600 -1360 32610 -1325
rect 32645 -1360 32655 -1325
rect 32690 -1360 32700 -1325
rect 32735 -1360 32745 -1325
rect 32780 -1360 32790 -1325
rect 32825 -1360 32835 -1325
rect 32870 -1360 32890 -1325
rect 31290 -1370 32890 -1360
rect 31290 -1405 31305 -1370
rect 31340 -1405 31350 -1370
rect 31385 -1405 31395 -1370
rect 31430 -1405 31440 -1370
rect 31475 -1405 31485 -1370
rect 31520 -1405 31530 -1370
rect 31565 -1405 31575 -1370
rect 31610 -1405 31620 -1370
rect 31655 -1405 31665 -1370
rect 31700 -1405 31710 -1370
rect 31745 -1405 31755 -1370
rect 31790 -1405 31800 -1370
rect 31835 -1405 31845 -1370
rect 31880 -1405 31890 -1370
rect 31925 -1405 31935 -1370
rect 31970 -1405 31980 -1370
rect 32015 -1405 32025 -1370
rect 32060 -1405 32070 -1370
rect 32105 -1405 32115 -1370
rect 32150 -1405 32160 -1370
rect 32195 -1405 32205 -1370
rect 32240 -1405 32250 -1370
rect 32285 -1405 32295 -1370
rect 32330 -1405 32340 -1370
rect 32375 -1405 32385 -1370
rect 32420 -1405 32430 -1370
rect 32465 -1405 32475 -1370
rect 32510 -1405 32520 -1370
rect 32555 -1405 32565 -1370
rect 32600 -1405 32610 -1370
rect 32645 -1405 32655 -1370
rect 32690 -1405 32700 -1370
rect 32735 -1405 32745 -1370
rect 32780 -1405 32790 -1370
rect 32825 -1405 32835 -1370
rect 32870 -1405 32890 -1370
rect 31290 -1415 32890 -1405
rect 31290 -1450 31305 -1415
rect 31340 -1450 31350 -1415
rect 31385 -1450 31395 -1415
rect 31430 -1450 31440 -1415
rect 31475 -1450 31485 -1415
rect 31520 -1450 31530 -1415
rect 31565 -1450 31575 -1415
rect 31610 -1450 31620 -1415
rect 31655 -1450 31665 -1415
rect 31700 -1450 31710 -1415
rect 31745 -1450 31755 -1415
rect 31790 -1450 31800 -1415
rect 31835 -1450 31845 -1415
rect 31880 -1450 31890 -1415
rect 31925 -1450 31935 -1415
rect 31970 -1450 31980 -1415
rect 32015 -1450 32025 -1415
rect 32060 -1450 32070 -1415
rect 32105 -1450 32115 -1415
rect 32150 -1450 32160 -1415
rect 32195 -1450 32205 -1415
rect 32240 -1450 32250 -1415
rect 32285 -1450 32295 -1415
rect 32330 -1450 32340 -1415
rect 32375 -1450 32385 -1415
rect 32420 -1450 32430 -1415
rect 32465 -1450 32475 -1415
rect 32510 -1450 32520 -1415
rect 32555 -1450 32565 -1415
rect 32600 -1450 32610 -1415
rect 32645 -1450 32655 -1415
rect 32690 -1450 32700 -1415
rect 32735 -1450 32745 -1415
rect 32780 -1450 32790 -1415
rect 32825 -1450 32835 -1415
rect 32870 -1450 32890 -1415
rect 31290 -1460 32890 -1450
rect 31290 -1495 31305 -1460
rect 31340 -1495 31350 -1460
rect 31385 -1495 31395 -1460
rect 31430 -1495 31440 -1460
rect 31475 -1495 31485 -1460
rect 31520 -1495 31530 -1460
rect 31565 -1495 31575 -1460
rect 31610 -1495 31620 -1460
rect 31655 -1495 31665 -1460
rect 31700 -1495 31710 -1460
rect 31745 -1495 31755 -1460
rect 31790 -1495 31800 -1460
rect 31835 -1495 31845 -1460
rect 31880 -1495 31890 -1460
rect 31925 -1495 31935 -1460
rect 31970 -1495 31980 -1460
rect 32015 -1495 32025 -1460
rect 32060 -1495 32070 -1460
rect 32105 -1495 32115 -1460
rect 32150 -1495 32160 -1460
rect 32195 -1495 32205 -1460
rect 32240 -1495 32250 -1460
rect 32285 -1495 32295 -1460
rect 32330 -1495 32340 -1460
rect 32375 -1495 32385 -1460
rect 32420 -1495 32430 -1460
rect 32465 -1495 32475 -1460
rect 32510 -1495 32520 -1460
rect 32555 -1495 32565 -1460
rect 32600 -1495 32610 -1460
rect 32645 -1495 32655 -1460
rect 32690 -1495 32700 -1460
rect 32735 -1495 32745 -1460
rect 32780 -1495 32790 -1460
rect 32825 -1495 32835 -1460
rect 32870 -1495 32890 -1460
rect 31290 -1505 32890 -1495
rect 31290 -1540 31305 -1505
rect 31340 -1540 31350 -1505
rect 31385 -1540 31395 -1505
rect 31430 -1540 31440 -1505
rect 31475 -1540 31485 -1505
rect 31520 -1540 31530 -1505
rect 31565 -1540 31575 -1505
rect 31610 -1540 31620 -1505
rect 31655 -1540 31665 -1505
rect 31700 -1540 31710 -1505
rect 31745 -1540 31755 -1505
rect 31790 -1540 31800 -1505
rect 31835 -1540 31845 -1505
rect 31880 -1540 31890 -1505
rect 31925 -1540 31935 -1505
rect 31970 -1540 31980 -1505
rect 32015 -1540 32025 -1505
rect 32060 -1540 32070 -1505
rect 32105 -1540 32115 -1505
rect 32150 -1540 32160 -1505
rect 32195 -1540 32205 -1505
rect 32240 -1540 32250 -1505
rect 32285 -1540 32295 -1505
rect 32330 -1540 32340 -1505
rect 32375 -1540 32385 -1505
rect 32420 -1540 32430 -1505
rect 32465 -1540 32475 -1505
rect 32510 -1540 32520 -1505
rect 32555 -1540 32565 -1505
rect 32600 -1540 32610 -1505
rect 32645 -1540 32655 -1505
rect 32690 -1540 32700 -1505
rect 32735 -1540 32745 -1505
rect 32780 -1540 32790 -1505
rect 32825 -1540 32835 -1505
rect 32870 -1540 32890 -1505
rect 31290 -1550 32890 -1540
rect 31290 -1585 31305 -1550
rect 31340 -1585 31350 -1550
rect 31385 -1585 31395 -1550
rect 31430 -1585 31440 -1550
rect 31475 -1585 31485 -1550
rect 31520 -1585 31530 -1550
rect 31565 -1585 31575 -1550
rect 31610 -1585 31620 -1550
rect 31655 -1585 31665 -1550
rect 31700 -1585 31710 -1550
rect 31745 -1585 31755 -1550
rect 31790 -1585 31800 -1550
rect 31835 -1585 31845 -1550
rect 31880 -1585 31890 -1550
rect 31925 -1585 31935 -1550
rect 31970 -1585 31980 -1550
rect 32015 -1585 32025 -1550
rect 32060 -1585 32070 -1550
rect 32105 -1585 32115 -1550
rect 32150 -1585 32160 -1550
rect 32195 -1585 32205 -1550
rect 32240 -1585 32250 -1550
rect 32285 -1585 32295 -1550
rect 32330 -1585 32340 -1550
rect 32375 -1585 32385 -1550
rect 32420 -1585 32430 -1550
rect 32465 -1585 32475 -1550
rect 32510 -1585 32520 -1550
rect 32555 -1585 32565 -1550
rect 32600 -1585 32610 -1550
rect 32645 -1585 32655 -1550
rect 32690 -1585 32700 -1550
rect 32735 -1585 32745 -1550
rect 32780 -1585 32790 -1550
rect 32825 -1585 32835 -1550
rect 32870 -1585 32890 -1550
rect 31290 -1595 32890 -1585
rect 31290 -1630 31305 -1595
rect 31340 -1630 31350 -1595
rect 31385 -1630 31395 -1595
rect 31430 -1630 31440 -1595
rect 31475 -1630 31485 -1595
rect 31520 -1630 31530 -1595
rect 31565 -1630 31575 -1595
rect 31610 -1630 31620 -1595
rect 31655 -1630 31665 -1595
rect 31700 -1630 31710 -1595
rect 31745 -1630 31755 -1595
rect 31790 -1630 31800 -1595
rect 31835 -1630 31845 -1595
rect 31880 -1630 31890 -1595
rect 31925 -1630 31935 -1595
rect 31970 -1630 31980 -1595
rect 32015 -1630 32025 -1595
rect 32060 -1630 32070 -1595
rect 32105 -1630 32115 -1595
rect 32150 -1630 32160 -1595
rect 32195 -1630 32205 -1595
rect 32240 -1630 32250 -1595
rect 32285 -1630 32295 -1595
rect 32330 -1630 32340 -1595
rect 32375 -1630 32385 -1595
rect 32420 -1630 32430 -1595
rect 32465 -1630 32475 -1595
rect 32510 -1630 32520 -1595
rect 32555 -1630 32565 -1595
rect 32600 -1630 32610 -1595
rect 32645 -1630 32655 -1595
rect 32690 -1630 32700 -1595
rect 32735 -1630 32745 -1595
rect 32780 -1630 32790 -1595
rect 32825 -1630 32835 -1595
rect 32870 -1630 32890 -1595
rect 31290 -1640 32890 -1630
rect 31290 -1675 31305 -1640
rect 31340 -1675 31350 -1640
rect 31385 -1675 31395 -1640
rect 31430 -1675 31440 -1640
rect 31475 -1675 31485 -1640
rect 31520 -1675 31530 -1640
rect 31565 -1675 31575 -1640
rect 31610 -1675 31620 -1640
rect 31655 -1675 31665 -1640
rect 31700 -1675 31710 -1640
rect 31745 -1675 31755 -1640
rect 31790 -1675 31800 -1640
rect 31835 -1675 31845 -1640
rect 31880 -1675 31890 -1640
rect 31925 -1675 31935 -1640
rect 31970 -1675 31980 -1640
rect 32015 -1675 32025 -1640
rect 32060 -1675 32070 -1640
rect 32105 -1675 32115 -1640
rect 32150 -1675 32160 -1640
rect 32195 -1675 32205 -1640
rect 32240 -1675 32250 -1640
rect 32285 -1675 32295 -1640
rect 32330 -1675 32340 -1640
rect 32375 -1675 32385 -1640
rect 32420 -1675 32430 -1640
rect 32465 -1675 32475 -1640
rect 32510 -1675 32520 -1640
rect 32555 -1675 32565 -1640
rect 32600 -1675 32610 -1640
rect 32645 -1675 32655 -1640
rect 32690 -1675 32700 -1640
rect 32735 -1675 32745 -1640
rect 32780 -1675 32790 -1640
rect 32825 -1675 32835 -1640
rect 32870 -1675 32890 -1640
rect 31290 -1685 32890 -1675
rect 31290 -1720 31305 -1685
rect 31340 -1720 31350 -1685
rect 31385 -1720 31395 -1685
rect 31430 -1720 31440 -1685
rect 31475 -1720 31485 -1685
rect 31520 -1720 31530 -1685
rect 31565 -1720 31575 -1685
rect 31610 -1720 31620 -1685
rect 31655 -1720 31665 -1685
rect 31700 -1720 31710 -1685
rect 31745 -1720 31755 -1685
rect 31790 -1720 31800 -1685
rect 31835 -1720 31845 -1685
rect 31880 -1720 31890 -1685
rect 31925 -1720 31935 -1685
rect 31970 -1720 31980 -1685
rect 32015 -1720 32025 -1685
rect 32060 -1720 32070 -1685
rect 32105 -1720 32115 -1685
rect 32150 -1720 32160 -1685
rect 32195 -1720 32205 -1685
rect 32240 -1720 32250 -1685
rect 32285 -1720 32295 -1685
rect 32330 -1720 32340 -1685
rect 32375 -1720 32385 -1685
rect 32420 -1720 32430 -1685
rect 32465 -1720 32475 -1685
rect 32510 -1720 32520 -1685
rect 32555 -1720 32565 -1685
rect 32600 -1720 32610 -1685
rect 32645 -1720 32655 -1685
rect 32690 -1720 32700 -1685
rect 32735 -1720 32745 -1685
rect 32780 -1720 32790 -1685
rect 32825 -1720 32835 -1685
rect 32870 -1720 32890 -1685
rect 31290 -1730 32890 -1720
rect 31290 -1765 31305 -1730
rect 31340 -1765 31350 -1730
rect 31385 -1765 31395 -1730
rect 31430 -1765 31440 -1730
rect 31475 -1765 31485 -1730
rect 31520 -1765 31530 -1730
rect 31565 -1765 31575 -1730
rect 31610 -1765 31620 -1730
rect 31655 -1765 31665 -1730
rect 31700 -1765 31710 -1730
rect 31745 -1765 31755 -1730
rect 31790 -1765 31800 -1730
rect 31835 -1765 31845 -1730
rect 31880 -1765 31890 -1730
rect 31925 -1765 31935 -1730
rect 31970 -1765 31980 -1730
rect 32015 -1765 32025 -1730
rect 32060 -1765 32070 -1730
rect 32105 -1765 32115 -1730
rect 32150 -1765 32160 -1730
rect 32195 -1765 32205 -1730
rect 32240 -1765 32250 -1730
rect 32285 -1765 32295 -1730
rect 32330 -1765 32340 -1730
rect 32375 -1765 32385 -1730
rect 32420 -1765 32430 -1730
rect 32465 -1765 32475 -1730
rect 32510 -1765 32520 -1730
rect 32555 -1765 32565 -1730
rect 32600 -1765 32610 -1730
rect 32645 -1765 32655 -1730
rect 32690 -1765 32700 -1730
rect 32735 -1765 32745 -1730
rect 32780 -1765 32790 -1730
rect 32825 -1765 32835 -1730
rect 32870 -1765 32890 -1730
rect 31290 -1775 32890 -1765
rect 31290 -1810 31305 -1775
rect 31340 -1810 31350 -1775
rect 31385 -1810 31395 -1775
rect 31430 -1810 31440 -1775
rect 31475 -1810 31485 -1775
rect 31520 -1810 31530 -1775
rect 31565 -1810 31575 -1775
rect 31610 -1810 31620 -1775
rect 31655 -1810 31665 -1775
rect 31700 -1810 31710 -1775
rect 31745 -1810 31755 -1775
rect 31790 -1810 31800 -1775
rect 31835 -1810 31845 -1775
rect 31880 -1810 31890 -1775
rect 31925 -1810 31935 -1775
rect 31970 -1810 31980 -1775
rect 32015 -1810 32025 -1775
rect 32060 -1810 32070 -1775
rect 32105 -1810 32115 -1775
rect 32150 -1810 32160 -1775
rect 32195 -1810 32205 -1775
rect 32240 -1810 32250 -1775
rect 32285 -1810 32295 -1775
rect 32330 -1810 32340 -1775
rect 32375 -1810 32385 -1775
rect 32420 -1810 32430 -1775
rect 32465 -1810 32475 -1775
rect 32510 -1810 32520 -1775
rect 32555 -1810 32565 -1775
rect 32600 -1810 32610 -1775
rect 32645 -1810 32655 -1775
rect 32690 -1810 32700 -1775
rect 32735 -1810 32745 -1775
rect 32780 -1810 32790 -1775
rect 32825 -1810 32835 -1775
rect 32870 -1810 32890 -1775
rect 31290 -1820 32890 -1810
rect 31290 -1855 31305 -1820
rect 31340 -1855 31350 -1820
rect 31385 -1855 31395 -1820
rect 31430 -1855 31440 -1820
rect 31475 -1855 31485 -1820
rect 31520 -1855 31530 -1820
rect 31565 -1855 31575 -1820
rect 31610 -1855 31620 -1820
rect 31655 -1855 31665 -1820
rect 31700 -1855 31710 -1820
rect 31745 -1855 31755 -1820
rect 31790 -1855 31800 -1820
rect 31835 -1855 31845 -1820
rect 31880 -1855 31890 -1820
rect 31925 -1855 31935 -1820
rect 31970 -1855 31980 -1820
rect 32015 -1855 32025 -1820
rect 32060 -1855 32070 -1820
rect 32105 -1855 32115 -1820
rect 32150 -1855 32160 -1820
rect 32195 -1855 32205 -1820
rect 32240 -1855 32250 -1820
rect 32285 -1855 32295 -1820
rect 32330 -1855 32340 -1820
rect 32375 -1855 32385 -1820
rect 32420 -1855 32430 -1820
rect 32465 -1855 32475 -1820
rect 32510 -1855 32520 -1820
rect 32555 -1855 32565 -1820
rect 32600 -1855 32610 -1820
rect 32645 -1855 32655 -1820
rect 32690 -1855 32700 -1820
rect 32735 -1855 32745 -1820
rect 32780 -1855 32790 -1820
rect 32825 -1855 32835 -1820
rect 32870 -1855 32890 -1820
rect 31290 -1865 32890 -1855
rect 31290 -1900 31305 -1865
rect 31340 -1900 31350 -1865
rect 31385 -1900 31395 -1865
rect 31430 -1900 31440 -1865
rect 31475 -1900 31485 -1865
rect 31520 -1900 31530 -1865
rect 31565 -1900 31575 -1865
rect 31610 -1900 31620 -1865
rect 31655 -1900 31665 -1865
rect 31700 -1900 31710 -1865
rect 31745 -1900 31755 -1865
rect 31790 -1900 31800 -1865
rect 31835 -1900 31845 -1865
rect 31880 -1900 31890 -1865
rect 31925 -1900 31935 -1865
rect 31970 -1900 31980 -1865
rect 32015 -1900 32025 -1865
rect 32060 -1900 32070 -1865
rect 32105 -1900 32115 -1865
rect 32150 -1900 32160 -1865
rect 32195 -1900 32205 -1865
rect 32240 -1900 32250 -1865
rect 32285 -1900 32295 -1865
rect 32330 -1900 32340 -1865
rect 32375 -1900 32385 -1865
rect 32420 -1900 32430 -1865
rect 32465 -1900 32475 -1865
rect 32510 -1900 32520 -1865
rect 32555 -1900 32565 -1865
rect 32600 -1900 32610 -1865
rect 32645 -1900 32655 -1865
rect 32690 -1900 32700 -1865
rect 32735 -1900 32745 -1865
rect 32780 -1900 32790 -1865
rect 32825 -1900 32835 -1865
rect 32870 -1900 32890 -1865
rect 31290 -1910 32890 -1900
rect 31290 -1945 31305 -1910
rect 31340 -1945 31350 -1910
rect 31385 -1945 31395 -1910
rect 31430 -1945 31440 -1910
rect 31475 -1945 31485 -1910
rect 31520 -1945 31530 -1910
rect 31565 -1945 31575 -1910
rect 31610 -1945 31620 -1910
rect 31655 -1945 31665 -1910
rect 31700 -1945 31710 -1910
rect 31745 -1945 31755 -1910
rect 31790 -1945 31800 -1910
rect 31835 -1945 31845 -1910
rect 31880 -1945 31890 -1910
rect 31925 -1945 31935 -1910
rect 31970 -1945 31980 -1910
rect 32015 -1945 32025 -1910
rect 32060 -1945 32070 -1910
rect 32105 -1945 32115 -1910
rect 32150 -1945 32160 -1910
rect 32195 -1945 32205 -1910
rect 32240 -1945 32250 -1910
rect 32285 -1945 32295 -1910
rect 32330 -1945 32340 -1910
rect 32375 -1945 32385 -1910
rect 32420 -1945 32430 -1910
rect 32465 -1945 32475 -1910
rect 32510 -1945 32520 -1910
rect 32555 -1945 32565 -1910
rect 32600 -1945 32610 -1910
rect 32645 -1945 32655 -1910
rect 32690 -1945 32700 -1910
rect 32735 -1945 32745 -1910
rect 32780 -1945 32790 -1910
rect 32825 -1945 32835 -1910
rect 32870 -1945 32890 -1910
rect 31290 -1955 32890 -1945
rect 31290 -1990 31305 -1955
rect 31340 -1990 31350 -1955
rect 31385 -1990 31395 -1955
rect 31430 -1990 31440 -1955
rect 31475 -1990 31485 -1955
rect 31520 -1990 31530 -1955
rect 31565 -1990 31575 -1955
rect 31610 -1990 31620 -1955
rect 31655 -1990 31665 -1955
rect 31700 -1990 31710 -1955
rect 31745 -1990 31755 -1955
rect 31790 -1990 31800 -1955
rect 31835 -1990 31845 -1955
rect 31880 -1990 31890 -1955
rect 31925 -1990 31935 -1955
rect 31970 -1990 31980 -1955
rect 32015 -1990 32025 -1955
rect 32060 -1990 32070 -1955
rect 32105 -1990 32115 -1955
rect 32150 -1990 32160 -1955
rect 32195 -1990 32205 -1955
rect 32240 -1990 32250 -1955
rect 32285 -1990 32295 -1955
rect 32330 -1990 32340 -1955
rect 32375 -1990 32385 -1955
rect 32420 -1990 32430 -1955
rect 32465 -1990 32475 -1955
rect 32510 -1990 32520 -1955
rect 32555 -1990 32565 -1955
rect 32600 -1990 32610 -1955
rect 32645 -1990 32655 -1955
rect 32690 -1990 32700 -1955
rect 32735 -1990 32745 -1955
rect 32780 -1990 32790 -1955
rect 32825 -1990 32835 -1955
rect 32870 -1990 32890 -1955
rect 31290 -2000 32890 -1990
rect 31290 -2035 31305 -2000
rect 31340 -2035 31350 -2000
rect 31385 -2035 31395 -2000
rect 31430 -2035 31440 -2000
rect 31475 -2035 31485 -2000
rect 31520 -2035 31530 -2000
rect 31565 -2035 31575 -2000
rect 31610 -2035 31620 -2000
rect 31655 -2035 31665 -2000
rect 31700 -2035 31710 -2000
rect 31745 -2035 31755 -2000
rect 31790 -2035 31800 -2000
rect 31835 -2035 31845 -2000
rect 31880 -2035 31890 -2000
rect 31925 -2035 31935 -2000
rect 31970 -2035 31980 -2000
rect 32015 -2035 32025 -2000
rect 32060 -2035 32070 -2000
rect 32105 -2035 32115 -2000
rect 32150 -2035 32160 -2000
rect 32195 -2035 32205 -2000
rect 32240 -2035 32250 -2000
rect 32285 -2035 32295 -2000
rect 32330 -2035 32340 -2000
rect 32375 -2035 32385 -2000
rect 32420 -2035 32430 -2000
rect 32465 -2035 32475 -2000
rect 32510 -2035 32520 -2000
rect 32555 -2035 32565 -2000
rect 32600 -2035 32610 -2000
rect 32645 -2035 32655 -2000
rect 32690 -2035 32700 -2000
rect 32735 -2035 32745 -2000
rect 32780 -2035 32790 -2000
rect 32825 -2035 32835 -2000
rect 32870 -2035 32890 -2000
rect 31290 -2045 32890 -2035
rect 31290 -2080 31305 -2045
rect 31340 -2080 31350 -2045
rect 31385 -2080 31395 -2045
rect 31430 -2080 31440 -2045
rect 31475 -2080 31485 -2045
rect 31520 -2080 31530 -2045
rect 31565 -2080 31575 -2045
rect 31610 -2080 31620 -2045
rect 31655 -2080 31665 -2045
rect 31700 -2080 31710 -2045
rect 31745 -2080 31755 -2045
rect 31790 -2080 31800 -2045
rect 31835 -2080 31845 -2045
rect 31880 -2080 31890 -2045
rect 31925 -2080 31935 -2045
rect 31970 -2080 31980 -2045
rect 32015 -2080 32025 -2045
rect 32060 -2080 32070 -2045
rect 32105 -2080 32115 -2045
rect 32150 -2080 32160 -2045
rect 32195 -2080 32205 -2045
rect 32240 -2080 32250 -2045
rect 32285 -2080 32295 -2045
rect 32330 -2080 32340 -2045
rect 32375 -2080 32385 -2045
rect 32420 -2080 32430 -2045
rect 32465 -2080 32475 -2045
rect 32510 -2080 32520 -2045
rect 32555 -2080 32565 -2045
rect 32600 -2080 32610 -2045
rect 32645 -2080 32655 -2045
rect 32690 -2080 32700 -2045
rect 32735 -2080 32745 -2045
rect 32780 -2080 32790 -2045
rect 32825 -2080 32835 -2045
rect 32870 -2080 32890 -2045
rect 31290 -2090 32890 -2080
rect 31290 -2125 31305 -2090
rect 31340 -2125 31350 -2090
rect 31385 -2125 31395 -2090
rect 31430 -2125 31440 -2090
rect 31475 -2125 31485 -2090
rect 31520 -2125 31530 -2090
rect 31565 -2125 31575 -2090
rect 31610 -2125 31620 -2090
rect 31655 -2125 31665 -2090
rect 31700 -2125 31710 -2090
rect 31745 -2125 31755 -2090
rect 31790 -2125 31800 -2090
rect 31835 -2125 31845 -2090
rect 31880 -2125 31890 -2090
rect 31925 -2125 31935 -2090
rect 31970 -2125 31980 -2090
rect 32015 -2125 32025 -2090
rect 32060 -2125 32070 -2090
rect 32105 -2125 32115 -2090
rect 32150 -2125 32160 -2090
rect 32195 -2125 32205 -2090
rect 32240 -2125 32250 -2090
rect 32285 -2125 32295 -2090
rect 32330 -2125 32340 -2090
rect 32375 -2125 32385 -2090
rect 32420 -2125 32430 -2090
rect 32465 -2125 32475 -2090
rect 32510 -2125 32520 -2090
rect 32555 -2125 32565 -2090
rect 32600 -2125 32610 -2090
rect 32645 -2125 32655 -2090
rect 32690 -2125 32700 -2090
rect 32735 -2125 32745 -2090
rect 32780 -2125 32790 -2090
rect 32825 -2125 32835 -2090
rect 32870 -2125 32890 -2090
rect 31290 -2135 32890 -2125
rect 31290 -2170 31305 -2135
rect 31340 -2170 31350 -2135
rect 31385 -2170 31395 -2135
rect 31430 -2170 31440 -2135
rect 31475 -2170 31485 -2135
rect 31520 -2170 31530 -2135
rect 31565 -2170 31575 -2135
rect 31610 -2170 31620 -2135
rect 31655 -2170 31665 -2135
rect 31700 -2170 31710 -2135
rect 31745 -2170 31755 -2135
rect 31790 -2170 31800 -2135
rect 31835 -2170 31845 -2135
rect 31880 -2170 31890 -2135
rect 31925 -2170 31935 -2135
rect 31970 -2170 31980 -2135
rect 32015 -2170 32025 -2135
rect 32060 -2170 32070 -2135
rect 32105 -2170 32115 -2135
rect 32150 -2170 32160 -2135
rect 32195 -2170 32205 -2135
rect 32240 -2170 32250 -2135
rect 32285 -2170 32295 -2135
rect 32330 -2170 32340 -2135
rect 32375 -2170 32385 -2135
rect 32420 -2170 32430 -2135
rect 32465 -2170 32475 -2135
rect 32510 -2170 32520 -2135
rect 32555 -2170 32565 -2135
rect 32600 -2170 32610 -2135
rect 32645 -2170 32655 -2135
rect 32690 -2170 32700 -2135
rect 32735 -2170 32745 -2135
rect 32780 -2170 32790 -2135
rect 32825 -2170 32835 -2135
rect 32870 -2170 32890 -2135
rect 31290 -2180 32890 -2170
rect 31290 -2215 31305 -2180
rect 31340 -2215 31350 -2180
rect 31385 -2215 31395 -2180
rect 31430 -2215 31440 -2180
rect 31475 -2215 31485 -2180
rect 31520 -2215 31530 -2180
rect 31565 -2215 31575 -2180
rect 31610 -2215 31620 -2180
rect 31655 -2215 31665 -2180
rect 31700 -2215 31710 -2180
rect 31745 -2215 31755 -2180
rect 31790 -2215 31800 -2180
rect 31835 -2215 31845 -2180
rect 31880 -2215 31890 -2180
rect 31925 -2215 31935 -2180
rect 31970 -2215 31980 -2180
rect 32015 -2215 32025 -2180
rect 32060 -2215 32070 -2180
rect 32105 -2215 32115 -2180
rect 32150 -2215 32160 -2180
rect 32195 -2215 32205 -2180
rect 32240 -2215 32250 -2180
rect 32285 -2215 32295 -2180
rect 32330 -2215 32340 -2180
rect 32375 -2215 32385 -2180
rect 32420 -2215 32430 -2180
rect 32465 -2215 32475 -2180
rect 32510 -2215 32520 -2180
rect 32555 -2215 32565 -2180
rect 32600 -2215 32610 -2180
rect 32645 -2215 32655 -2180
rect 32690 -2215 32700 -2180
rect 32735 -2215 32745 -2180
rect 32780 -2215 32790 -2180
rect 32825 -2215 32835 -2180
rect 32870 -2215 32890 -2180
rect 31290 -2225 32890 -2215
rect 31290 -2260 31305 -2225
rect 31340 -2260 31350 -2225
rect 31385 -2260 31395 -2225
rect 31430 -2260 31440 -2225
rect 31475 -2260 31485 -2225
rect 31520 -2260 31530 -2225
rect 31565 -2260 31575 -2225
rect 31610 -2260 31620 -2225
rect 31655 -2260 31665 -2225
rect 31700 -2260 31710 -2225
rect 31745 -2260 31755 -2225
rect 31790 -2260 31800 -2225
rect 31835 -2260 31845 -2225
rect 31880 -2260 31890 -2225
rect 31925 -2260 31935 -2225
rect 31970 -2260 31980 -2225
rect 32015 -2260 32025 -2225
rect 32060 -2260 32070 -2225
rect 32105 -2260 32115 -2225
rect 32150 -2260 32160 -2225
rect 32195 -2260 32205 -2225
rect 32240 -2260 32250 -2225
rect 32285 -2260 32295 -2225
rect 32330 -2260 32340 -2225
rect 32375 -2260 32385 -2225
rect 32420 -2260 32430 -2225
rect 32465 -2260 32475 -2225
rect 32510 -2260 32520 -2225
rect 32555 -2260 32565 -2225
rect 32600 -2260 32610 -2225
rect 32645 -2260 32655 -2225
rect 32690 -2260 32700 -2225
rect 32735 -2260 32745 -2225
rect 32780 -2260 32790 -2225
rect 32825 -2260 32835 -2225
rect 32870 -2260 32890 -2225
rect 31290 -2270 32890 -2260
rect 31290 -2305 31305 -2270
rect 31340 -2305 31350 -2270
rect 31385 -2305 31395 -2270
rect 31430 -2305 31440 -2270
rect 31475 -2305 31485 -2270
rect 31520 -2305 31530 -2270
rect 31565 -2305 31575 -2270
rect 31610 -2305 31620 -2270
rect 31655 -2305 31665 -2270
rect 31700 -2305 31710 -2270
rect 31745 -2305 31755 -2270
rect 31790 -2305 31800 -2270
rect 31835 -2305 31845 -2270
rect 31880 -2305 31890 -2270
rect 31925 -2305 31935 -2270
rect 31970 -2305 31980 -2270
rect 32015 -2305 32025 -2270
rect 32060 -2305 32070 -2270
rect 32105 -2305 32115 -2270
rect 32150 -2305 32160 -2270
rect 32195 -2305 32205 -2270
rect 32240 -2305 32250 -2270
rect 32285 -2305 32295 -2270
rect 32330 -2305 32340 -2270
rect 32375 -2305 32385 -2270
rect 32420 -2305 32430 -2270
rect 32465 -2305 32475 -2270
rect 32510 -2305 32520 -2270
rect 32555 -2305 32565 -2270
rect 32600 -2305 32610 -2270
rect 32645 -2305 32655 -2270
rect 32690 -2305 32700 -2270
rect 32735 -2305 32745 -2270
rect 32780 -2305 32790 -2270
rect 32825 -2305 32835 -2270
rect 32870 -2305 32890 -2270
rect 31290 -2315 32890 -2305
rect 31290 -2350 31305 -2315
rect 31340 -2350 31350 -2315
rect 31385 -2350 31395 -2315
rect 31430 -2350 31440 -2315
rect 31475 -2350 31485 -2315
rect 31520 -2350 31530 -2315
rect 31565 -2350 31575 -2315
rect 31610 -2350 31620 -2315
rect 31655 -2350 31665 -2315
rect 31700 -2350 31710 -2315
rect 31745 -2350 31755 -2315
rect 31790 -2350 31800 -2315
rect 31835 -2350 31845 -2315
rect 31880 -2350 31890 -2315
rect 31925 -2350 31935 -2315
rect 31970 -2350 31980 -2315
rect 32015 -2350 32025 -2315
rect 32060 -2350 32070 -2315
rect 32105 -2350 32115 -2315
rect 32150 -2350 32160 -2315
rect 32195 -2350 32205 -2315
rect 32240 -2350 32250 -2315
rect 32285 -2350 32295 -2315
rect 32330 -2350 32340 -2315
rect 32375 -2350 32385 -2315
rect 32420 -2350 32430 -2315
rect 32465 -2350 32475 -2315
rect 32510 -2350 32520 -2315
rect 32555 -2350 32565 -2315
rect 32600 -2350 32610 -2315
rect 32645 -2350 32655 -2315
rect 32690 -2350 32700 -2315
rect 32735 -2350 32745 -2315
rect 32780 -2350 32790 -2315
rect 32825 -2350 32835 -2315
rect 32870 -2350 32890 -2315
rect 31290 -2360 32890 -2350
rect 31290 -2395 31305 -2360
rect 31340 -2395 31350 -2360
rect 31385 -2395 31395 -2360
rect 31430 -2395 31440 -2360
rect 31475 -2395 31485 -2360
rect 31520 -2395 31530 -2360
rect 31565 -2395 31575 -2360
rect 31610 -2395 31620 -2360
rect 31655 -2395 31665 -2360
rect 31700 -2395 31710 -2360
rect 31745 -2395 31755 -2360
rect 31790 -2395 31800 -2360
rect 31835 -2395 31845 -2360
rect 31880 -2395 31890 -2360
rect 31925 -2395 31935 -2360
rect 31970 -2395 31980 -2360
rect 32015 -2395 32025 -2360
rect 32060 -2395 32070 -2360
rect 32105 -2395 32115 -2360
rect 32150 -2395 32160 -2360
rect 32195 -2395 32205 -2360
rect 32240 -2395 32250 -2360
rect 32285 -2395 32295 -2360
rect 32330 -2395 32340 -2360
rect 32375 -2395 32385 -2360
rect 32420 -2395 32430 -2360
rect 32465 -2395 32475 -2360
rect 32510 -2395 32520 -2360
rect 32555 -2395 32565 -2360
rect 32600 -2395 32610 -2360
rect 32645 -2395 32655 -2360
rect 32690 -2395 32700 -2360
rect 32735 -2395 32745 -2360
rect 32780 -2395 32790 -2360
rect 32825 -2395 32835 -2360
rect 32870 -2395 32890 -2360
rect 31290 -2405 32890 -2395
rect 31290 -2440 31305 -2405
rect 31340 -2440 31350 -2405
rect 31385 -2440 31395 -2405
rect 31430 -2440 31440 -2405
rect 31475 -2440 31485 -2405
rect 31520 -2440 31530 -2405
rect 31565 -2440 31575 -2405
rect 31610 -2440 31620 -2405
rect 31655 -2440 31665 -2405
rect 31700 -2440 31710 -2405
rect 31745 -2440 31755 -2405
rect 31790 -2440 31800 -2405
rect 31835 -2440 31845 -2405
rect 31880 -2440 31890 -2405
rect 31925 -2440 31935 -2405
rect 31970 -2440 31980 -2405
rect 32015 -2440 32025 -2405
rect 32060 -2440 32070 -2405
rect 32105 -2440 32115 -2405
rect 32150 -2440 32160 -2405
rect 32195 -2440 32205 -2405
rect 32240 -2440 32250 -2405
rect 32285 -2440 32295 -2405
rect 32330 -2440 32340 -2405
rect 32375 -2440 32385 -2405
rect 32420 -2440 32430 -2405
rect 32465 -2440 32475 -2405
rect 32510 -2440 32520 -2405
rect 32555 -2440 32565 -2405
rect 32600 -2440 32610 -2405
rect 32645 -2440 32655 -2405
rect 32690 -2440 32700 -2405
rect 32735 -2440 32745 -2405
rect 32780 -2440 32790 -2405
rect 32825 -2440 32835 -2405
rect 32870 -2440 32890 -2405
rect 31290 -2450 32890 -2440
rect 31290 -2485 31305 -2450
rect 31340 -2485 31350 -2450
rect 31385 -2485 31395 -2450
rect 31430 -2485 31440 -2450
rect 31475 -2485 31485 -2450
rect 31520 -2485 31530 -2450
rect 31565 -2485 31575 -2450
rect 31610 -2485 31620 -2450
rect 31655 -2485 31665 -2450
rect 31700 -2485 31710 -2450
rect 31745 -2485 31755 -2450
rect 31790 -2485 31800 -2450
rect 31835 -2485 31845 -2450
rect 31880 -2485 31890 -2450
rect 31925 -2485 31935 -2450
rect 31970 -2485 31980 -2450
rect 32015 -2485 32025 -2450
rect 32060 -2485 32070 -2450
rect 32105 -2485 32115 -2450
rect 32150 -2485 32160 -2450
rect 32195 -2485 32205 -2450
rect 32240 -2485 32250 -2450
rect 32285 -2485 32295 -2450
rect 32330 -2485 32340 -2450
rect 32375 -2485 32385 -2450
rect 32420 -2485 32430 -2450
rect 32465 -2485 32475 -2450
rect 32510 -2485 32520 -2450
rect 32555 -2485 32565 -2450
rect 32600 -2485 32610 -2450
rect 32645 -2485 32655 -2450
rect 32690 -2485 32700 -2450
rect 32735 -2485 32745 -2450
rect 32780 -2485 32790 -2450
rect 32825 -2485 32835 -2450
rect 32870 -2485 32890 -2450
rect 31290 -2495 32890 -2485
rect 31290 -2530 31305 -2495
rect 31340 -2530 31350 -2495
rect 31385 -2530 31395 -2495
rect 31430 -2530 31440 -2495
rect 31475 -2530 31485 -2495
rect 31520 -2530 31530 -2495
rect 31565 -2530 31575 -2495
rect 31610 -2530 31620 -2495
rect 31655 -2530 31665 -2495
rect 31700 -2530 31710 -2495
rect 31745 -2530 31755 -2495
rect 31790 -2530 31800 -2495
rect 31835 -2530 31845 -2495
rect 31880 -2530 31890 -2495
rect 31925 -2530 31935 -2495
rect 31970 -2530 31980 -2495
rect 32015 -2530 32025 -2495
rect 32060 -2530 32070 -2495
rect 32105 -2530 32115 -2495
rect 32150 -2530 32160 -2495
rect 32195 -2530 32205 -2495
rect 32240 -2530 32250 -2495
rect 32285 -2530 32295 -2495
rect 32330 -2530 32340 -2495
rect 32375 -2530 32385 -2495
rect 32420 -2530 32430 -2495
rect 32465 -2530 32475 -2495
rect 32510 -2530 32520 -2495
rect 32555 -2530 32565 -2495
rect 32600 -2530 32610 -2495
rect 32645 -2530 32655 -2495
rect 32690 -2530 32700 -2495
rect 32735 -2530 32745 -2495
rect 32780 -2530 32790 -2495
rect 32825 -2530 32835 -2495
rect 32870 -2530 32890 -2495
rect 31290 -2540 32890 -2530
rect 31290 -2575 31305 -2540
rect 31340 -2575 31350 -2540
rect 31385 -2575 31395 -2540
rect 31430 -2575 31440 -2540
rect 31475 -2575 31485 -2540
rect 31520 -2575 31530 -2540
rect 31565 -2575 31575 -2540
rect 31610 -2575 31620 -2540
rect 31655 -2575 31665 -2540
rect 31700 -2575 31710 -2540
rect 31745 -2575 31755 -2540
rect 31790 -2575 31800 -2540
rect 31835 -2575 31845 -2540
rect 31880 -2575 31890 -2540
rect 31925 -2575 31935 -2540
rect 31970 -2575 31980 -2540
rect 32015 -2575 32025 -2540
rect 32060 -2575 32070 -2540
rect 32105 -2575 32115 -2540
rect 32150 -2575 32160 -2540
rect 32195 -2575 32205 -2540
rect 32240 -2575 32250 -2540
rect 32285 -2575 32295 -2540
rect 32330 -2575 32340 -2540
rect 32375 -2575 32385 -2540
rect 32420 -2575 32430 -2540
rect 32465 -2575 32475 -2540
rect 32510 -2575 32520 -2540
rect 32555 -2575 32565 -2540
rect 32600 -2575 32610 -2540
rect 32645 -2575 32655 -2540
rect 32690 -2575 32700 -2540
rect 32735 -2575 32745 -2540
rect 32780 -2575 32790 -2540
rect 32825 -2575 32835 -2540
rect 32870 -2575 32890 -2540
rect 31290 -2585 32890 -2575
rect 31290 -2620 31305 -2585
rect 31340 -2620 31350 -2585
rect 31385 -2620 31395 -2585
rect 31430 -2620 31440 -2585
rect 31475 -2620 31485 -2585
rect 31520 -2620 31530 -2585
rect 31565 -2620 31575 -2585
rect 31610 -2620 31620 -2585
rect 31655 -2620 31665 -2585
rect 31700 -2620 31710 -2585
rect 31745 -2620 31755 -2585
rect 31790 -2620 31800 -2585
rect 31835 -2620 31845 -2585
rect 31880 -2620 31890 -2585
rect 31925 -2620 31935 -2585
rect 31970 -2620 31980 -2585
rect 32015 -2620 32025 -2585
rect 32060 -2620 32070 -2585
rect 32105 -2620 32115 -2585
rect 32150 -2620 32160 -2585
rect 32195 -2620 32205 -2585
rect 32240 -2620 32250 -2585
rect 32285 -2620 32295 -2585
rect 32330 -2620 32340 -2585
rect 32375 -2620 32385 -2585
rect 32420 -2620 32430 -2585
rect 32465 -2620 32475 -2585
rect 32510 -2620 32520 -2585
rect 32555 -2620 32565 -2585
rect 32600 -2620 32610 -2585
rect 32645 -2620 32655 -2585
rect 32690 -2620 32700 -2585
rect 32735 -2620 32745 -2585
rect 32780 -2620 32790 -2585
rect 32825 -2620 32835 -2585
rect 32870 -2620 32890 -2585
rect 31290 -2630 32890 -2620
rect 31290 -2665 31305 -2630
rect 31340 -2665 31350 -2630
rect 31385 -2665 31395 -2630
rect 31430 -2665 31440 -2630
rect 31475 -2665 31485 -2630
rect 31520 -2665 31530 -2630
rect 31565 -2665 31575 -2630
rect 31610 -2665 31620 -2630
rect 31655 -2665 31665 -2630
rect 31700 -2665 31710 -2630
rect 31745 -2665 31755 -2630
rect 31790 -2665 31800 -2630
rect 31835 -2665 31845 -2630
rect 31880 -2665 31890 -2630
rect 31925 -2665 31935 -2630
rect 31970 -2665 31980 -2630
rect 32015 -2665 32025 -2630
rect 32060 -2665 32070 -2630
rect 32105 -2665 32115 -2630
rect 32150 -2665 32160 -2630
rect 32195 -2665 32205 -2630
rect 32240 -2665 32250 -2630
rect 32285 -2665 32295 -2630
rect 32330 -2665 32340 -2630
rect 32375 -2665 32385 -2630
rect 32420 -2665 32430 -2630
rect 32465 -2665 32475 -2630
rect 32510 -2665 32520 -2630
rect 32555 -2665 32565 -2630
rect 32600 -2665 32610 -2630
rect 32645 -2665 32655 -2630
rect 32690 -2665 32700 -2630
rect 32735 -2665 32745 -2630
rect 32780 -2665 32790 -2630
rect 32825 -2665 32835 -2630
rect 32870 -2665 32890 -2630
rect 31290 -2675 32890 -2665
rect 31290 -2710 31305 -2675
rect 31340 -2710 31350 -2675
rect 31385 -2710 31395 -2675
rect 31430 -2710 31440 -2675
rect 31475 -2710 31485 -2675
rect 31520 -2710 31530 -2675
rect 31565 -2710 31575 -2675
rect 31610 -2710 31620 -2675
rect 31655 -2710 31665 -2675
rect 31700 -2710 31710 -2675
rect 31745 -2710 31755 -2675
rect 31790 -2710 31800 -2675
rect 31835 -2710 31845 -2675
rect 31880 -2710 31890 -2675
rect 31925 -2710 31935 -2675
rect 31970 -2710 31980 -2675
rect 32015 -2710 32025 -2675
rect 32060 -2710 32070 -2675
rect 32105 -2710 32115 -2675
rect 32150 -2710 32160 -2675
rect 32195 -2710 32205 -2675
rect 32240 -2710 32250 -2675
rect 32285 -2710 32295 -2675
rect 32330 -2710 32340 -2675
rect 32375 -2710 32385 -2675
rect 32420 -2710 32430 -2675
rect 32465 -2710 32475 -2675
rect 32510 -2710 32520 -2675
rect 32555 -2710 32565 -2675
rect 32600 -2710 32610 -2675
rect 32645 -2710 32655 -2675
rect 32690 -2710 32700 -2675
rect 32735 -2710 32745 -2675
rect 32780 -2710 32790 -2675
rect 32825 -2710 32835 -2675
rect 32870 -2710 32890 -2675
rect 31290 -2720 32890 -2710
rect 31290 -2755 31305 -2720
rect 31340 -2755 31350 -2720
rect 31385 -2755 31395 -2720
rect 31430 -2755 31440 -2720
rect 31475 -2755 31485 -2720
rect 31520 -2755 31530 -2720
rect 31565 -2755 31575 -2720
rect 31610 -2755 31620 -2720
rect 31655 -2755 31665 -2720
rect 31700 -2755 31710 -2720
rect 31745 -2755 31755 -2720
rect 31790 -2755 31800 -2720
rect 31835 -2755 31845 -2720
rect 31880 -2755 31890 -2720
rect 31925 -2755 31935 -2720
rect 31970 -2755 31980 -2720
rect 32015 -2755 32025 -2720
rect 32060 -2755 32070 -2720
rect 32105 -2755 32115 -2720
rect 32150 -2755 32160 -2720
rect 32195 -2755 32205 -2720
rect 32240 -2755 32250 -2720
rect 32285 -2755 32295 -2720
rect 32330 -2755 32340 -2720
rect 32375 -2755 32385 -2720
rect 32420 -2755 32430 -2720
rect 32465 -2755 32475 -2720
rect 32510 -2755 32520 -2720
rect 32555 -2755 32565 -2720
rect 32600 -2755 32610 -2720
rect 32645 -2755 32655 -2720
rect 32690 -2755 32700 -2720
rect 32735 -2755 32745 -2720
rect 32780 -2755 32790 -2720
rect 32825 -2755 32835 -2720
rect 32870 -2755 32890 -2720
rect 31290 -2765 32890 -2755
rect 31290 -2800 31305 -2765
rect 31340 -2800 31350 -2765
rect 31385 -2800 31395 -2765
rect 31430 -2800 31440 -2765
rect 31475 -2800 31485 -2765
rect 31520 -2800 31530 -2765
rect 31565 -2800 31575 -2765
rect 31610 -2800 31620 -2765
rect 31655 -2800 31665 -2765
rect 31700 -2800 31710 -2765
rect 31745 -2800 31755 -2765
rect 31790 -2800 31800 -2765
rect 31835 -2800 31845 -2765
rect 31880 -2800 31890 -2765
rect 31925 -2800 31935 -2765
rect 31970 -2800 31980 -2765
rect 32015 -2800 32025 -2765
rect 32060 -2800 32070 -2765
rect 32105 -2800 32115 -2765
rect 32150 -2800 32160 -2765
rect 32195 -2800 32205 -2765
rect 32240 -2800 32250 -2765
rect 32285 -2800 32295 -2765
rect 32330 -2800 32340 -2765
rect 32375 -2800 32385 -2765
rect 32420 -2800 32430 -2765
rect 32465 -2800 32475 -2765
rect 32510 -2800 32520 -2765
rect 32555 -2800 32565 -2765
rect 32600 -2800 32610 -2765
rect 32645 -2800 32655 -2765
rect 32690 -2800 32700 -2765
rect 32735 -2800 32745 -2765
rect 32780 -2800 32790 -2765
rect 32825 -2800 32835 -2765
rect 32870 -2800 32890 -2765
rect 31290 -2810 32890 -2800
rect 31290 -2845 31305 -2810
rect 31340 -2845 31350 -2810
rect 31385 -2845 31395 -2810
rect 31430 -2845 31440 -2810
rect 31475 -2845 31485 -2810
rect 31520 -2845 31530 -2810
rect 31565 -2845 31575 -2810
rect 31610 -2845 31620 -2810
rect 31655 -2845 31665 -2810
rect 31700 -2845 31710 -2810
rect 31745 -2845 31755 -2810
rect 31790 -2845 31800 -2810
rect 31835 -2845 31845 -2810
rect 31880 -2845 31890 -2810
rect 31925 -2845 31935 -2810
rect 31970 -2845 31980 -2810
rect 32015 -2845 32025 -2810
rect 32060 -2845 32070 -2810
rect 32105 -2845 32115 -2810
rect 32150 -2845 32160 -2810
rect 32195 -2845 32205 -2810
rect 32240 -2845 32250 -2810
rect 32285 -2845 32295 -2810
rect 32330 -2845 32340 -2810
rect 32375 -2845 32385 -2810
rect 32420 -2845 32430 -2810
rect 32465 -2845 32475 -2810
rect 32510 -2845 32520 -2810
rect 32555 -2845 32565 -2810
rect 32600 -2845 32610 -2810
rect 32645 -2845 32655 -2810
rect 32690 -2845 32700 -2810
rect 32735 -2845 32745 -2810
rect 32780 -2845 32790 -2810
rect 32825 -2845 32835 -2810
rect 32870 -2845 32890 -2810
rect 31290 -2855 32890 -2845
rect 31290 -2890 31305 -2855
rect 31340 -2890 31350 -2855
rect 31385 -2890 31395 -2855
rect 31430 -2890 31440 -2855
rect 31475 -2890 31485 -2855
rect 31520 -2890 31530 -2855
rect 31565 -2890 31575 -2855
rect 31610 -2890 31620 -2855
rect 31655 -2890 31665 -2855
rect 31700 -2890 31710 -2855
rect 31745 -2890 31755 -2855
rect 31790 -2890 31800 -2855
rect 31835 -2890 31845 -2855
rect 31880 -2890 31890 -2855
rect 31925 -2890 31935 -2855
rect 31970 -2890 31980 -2855
rect 32015 -2890 32025 -2855
rect 32060 -2890 32070 -2855
rect 32105 -2890 32115 -2855
rect 32150 -2890 32160 -2855
rect 32195 -2890 32205 -2855
rect 32240 -2890 32250 -2855
rect 32285 -2890 32295 -2855
rect 32330 -2890 32340 -2855
rect 32375 -2890 32385 -2855
rect 32420 -2890 32430 -2855
rect 32465 -2890 32475 -2855
rect 32510 -2890 32520 -2855
rect 32555 -2890 32565 -2855
rect 32600 -2890 32610 -2855
rect 32645 -2890 32655 -2855
rect 32690 -2890 32700 -2855
rect 32735 -2890 32745 -2855
rect 32780 -2890 32790 -2855
rect 32825 -2890 32835 -2855
rect 32870 -2890 32890 -2855
rect 31290 -2905 32890 -2890
rect 3410 -3015 3470 -3005
rect 3410 -3055 3420 -3015
rect 3460 -3055 3470 -3015
rect 3410 -3080 3470 -3055
rect 3410 -3120 3420 -3080
rect 3460 -3120 3470 -3080
rect 3410 -3150 3470 -3120
rect 3410 -3190 3420 -3150
rect 3460 -3190 3470 -3150
rect 3410 -3220 3470 -3190
rect 3410 -3260 3420 -3220
rect 3460 -3260 3470 -3220
rect 3410 -3290 3470 -3260
rect 3410 -3330 3420 -3290
rect 3460 -3330 3470 -3290
rect 3410 -3355 3470 -3330
rect 3410 -3395 3420 -3355
rect 3460 -3395 3470 -3355
rect 3410 -3415 3470 -3395
rect 3410 -3455 3420 -3415
rect 3460 -3455 3470 -3415
rect 3410 -3480 3470 -3455
rect 3410 -3520 3420 -3480
rect 3460 -3520 3470 -3480
rect 3410 -3550 3470 -3520
rect 3410 -3590 3420 -3550
rect 3460 -3590 3470 -3550
rect 3410 -3620 3470 -3590
rect 3410 -3660 3420 -3620
rect 3460 -3660 3470 -3620
rect 3410 -3690 3470 -3660
rect 3410 -3730 3420 -3690
rect 3460 -3730 3470 -3690
rect 3410 -3755 3470 -3730
rect 3410 -3795 3420 -3755
rect 3460 -3795 3470 -3755
rect 3410 -3815 3470 -3795
rect 3410 -3855 3420 -3815
rect 3460 -3855 3470 -3815
rect 3410 -3880 3470 -3855
rect 3410 -3920 3420 -3880
rect 3460 -3920 3470 -3880
rect 3410 -3950 3470 -3920
rect 3410 -3990 3420 -3950
rect 3460 -3990 3470 -3950
rect 3410 -4020 3470 -3990
rect 3410 -4060 3420 -4020
rect 3460 -4060 3470 -4020
rect 3410 -4090 3470 -4060
rect 3410 -4130 3420 -4090
rect 3460 -4130 3470 -4090
rect 3410 -4155 3470 -4130
rect 3410 -4195 3420 -4155
rect 3460 -4195 3470 -4155
rect 3410 -4215 3470 -4195
rect 3410 -4255 3420 -4215
rect 3460 -4255 3470 -4215
rect 3410 -4280 3470 -4255
rect 3410 -4320 3420 -4280
rect 3460 -4320 3470 -4280
rect 3410 -4350 3470 -4320
rect 3410 -4390 3420 -4350
rect 3460 -4390 3470 -4350
rect 3410 -4420 3470 -4390
rect 3410 -4460 3420 -4420
rect 3460 -4460 3470 -4420
rect 3410 -4490 3470 -4460
rect 3410 -4530 3420 -4490
rect 3460 -4530 3470 -4490
rect 3410 -4555 3470 -4530
rect 3410 -4595 3420 -4555
rect 3460 -4595 3470 -4555
rect 3410 -4605 3470 -4595
rect 3760 -3015 3820 -3005
rect 3760 -3055 3770 -3015
rect 3810 -3055 3820 -3015
rect 3760 -3080 3820 -3055
rect 3760 -3120 3770 -3080
rect 3810 -3120 3820 -3080
rect 3760 -3150 3820 -3120
rect 3760 -3190 3770 -3150
rect 3810 -3190 3820 -3150
rect 3760 -3220 3820 -3190
rect 3760 -3260 3770 -3220
rect 3810 -3260 3820 -3220
rect 3760 -3290 3820 -3260
rect 3760 -3330 3770 -3290
rect 3810 -3330 3820 -3290
rect 3760 -3355 3820 -3330
rect 3760 -3395 3770 -3355
rect 3810 -3395 3820 -3355
rect 3760 -3415 3820 -3395
rect 3760 -3455 3770 -3415
rect 3810 -3455 3820 -3415
rect 3760 -3480 3820 -3455
rect 3760 -3520 3770 -3480
rect 3810 -3520 3820 -3480
rect 3760 -3550 3820 -3520
rect 3760 -3590 3770 -3550
rect 3810 -3590 3820 -3550
rect 3760 -3620 3820 -3590
rect 3760 -3660 3770 -3620
rect 3810 -3660 3820 -3620
rect 3760 -3690 3820 -3660
rect 3760 -3730 3770 -3690
rect 3810 -3730 3820 -3690
rect 3760 -3755 3820 -3730
rect 3760 -3795 3770 -3755
rect 3810 -3795 3820 -3755
rect 3760 -3815 3820 -3795
rect 3760 -3855 3770 -3815
rect 3810 -3855 3820 -3815
rect 3760 -3880 3820 -3855
rect 3760 -3920 3770 -3880
rect 3810 -3920 3820 -3880
rect 3760 -3950 3820 -3920
rect 3760 -3990 3770 -3950
rect 3810 -3990 3820 -3950
rect 3760 -4020 3820 -3990
rect 3760 -4060 3770 -4020
rect 3810 -4060 3820 -4020
rect 3760 -4090 3820 -4060
rect 3760 -4130 3770 -4090
rect 3810 -4130 3820 -4090
rect 3760 -4155 3820 -4130
rect 3760 -4195 3770 -4155
rect 3810 -4195 3820 -4155
rect 3760 -4215 3820 -4195
rect 3760 -4255 3770 -4215
rect 3810 -4255 3820 -4215
rect 3760 -4280 3820 -4255
rect 3760 -4320 3770 -4280
rect 3810 -4320 3820 -4280
rect 3760 -4350 3820 -4320
rect 3760 -4390 3770 -4350
rect 3810 -4390 3820 -4350
rect 3760 -4420 3820 -4390
rect 3760 -4460 3770 -4420
rect 3810 -4460 3820 -4420
rect 3760 -4490 3820 -4460
rect 3760 -4530 3770 -4490
rect 3810 -4530 3820 -4490
rect 3760 -4555 3820 -4530
rect 3760 -4595 3770 -4555
rect 3810 -4595 3820 -4555
rect 3760 -4605 3820 -4595
rect 4110 -3015 4170 -3005
rect 4110 -3055 4120 -3015
rect 4160 -3055 4170 -3015
rect 4110 -3080 4170 -3055
rect 4110 -3120 4120 -3080
rect 4160 -3120 4170 -3080
rect 4110 -3150 4170 -3120
rect 4110 -3190 4120 -3150
rect 4160 -3190 4170 -3150
rect 4110 -3220 4170 -3190
rect 4110 -3260 4120 -3220
rect 4160 -3260 4170 -3220
rect 4110 -3290 4170 -3260
rect 4110 -3330 4120 -3290
rect 4160 -3330 4170 -3290
rect 4110 -3355 4170 -3330
rect 4110 -3395 4120 -3355
rect 4160 -3395 4170 -3355
rect 4110 -3415 4170 -3395
rect 4110 -3455 4120 -3415
rect 4160 -3455 4170 -3415
rect 4110 -3480 4170 -3455
rect 4110 -3520 4120 -3480
rect 4160 -3520 4170 -3480
rect 4110 -3550 4170 -3520
rect 4110 -3590 4120 -3550
rect 4160 -3590 4170 -3550
rect 4110 -3620 4170 -3590
rect 4110 -3660 4120 -3620
rect 4160 -3660 4170 -3620
rect 4110 -3690 4170 -3660
rect 4110 -3730 4120 -3690
rect 4160 -3730 4170 -3690
rect 4110 -3755 4170 -3730
rect 4110 -3795 4120 -3755
rect 4160 -3795 4170 -3755
rect 4110 -3815 4170 -3795
rect 4110 -3855 4120 -3815
rect 4160 -3855 4170 -3815
rect 4110 -3880 4170 -3855
rect 4110 -3920 4120 -3880
rect 4160 -3920 4170 -3880
rect 4110 -3950 4170 -3920
rect 4110 -3990 4120 -3950
rect 4160 -3990 4170 -3950
rect 4110 -4020 4170 -3990
rect 4110 -4060 4120 -4020
rect 4160 -4060 4170 -4020
rect 4110 -4090 4170 -4060
rect 4110 -4130 4120 -4090
rect 4160 -4130 4170 -4090
rect 4110 -4155 4170 -4130
rect 4110 -4195 4120 -4155
rect 4160 -4195 4170 -4155
rect 4110 -4215 4170 -4195
rect 4110 -4255 4120 -4215
rect 4160 -4255 4170 -4215
rect 4110 -4280 4170 -4255
rect 4110 -4320 4120 -4280
rect 4160 -4320 4170 -4280
rect 4110 -4350 4170 -4320
rect 4110 -4390 4120 -4350
rect 4160 -4390 4170 -4350
rect 4110 -4420 4170 -4390
rect 4110 -4460 4120 -4420
rect 4160 -4460 4170 -4420
rect 4110 -4490 4170 -4460
rect 4110 -4530 4120 -4490
rect 4160 -4530 4170 -4490
rect 4110 -4555 4170 -4530
rect 4110 -4595 4120 -4555
rect 4160 -4595 4170 -4555
rect 4110 -4605 4170 -4595
rect 4460 -3015 4520 -3005
rect 4460 -3055 4470 -3015
rect 4510 -3055 4520 -3015
rect 4460 -3080 4520 -3055
rect 4460 -3120 4470 -3080
rect 4510 -3120 4520 -3080
rect 4460 -3150 4520 -3120
rect 4460 -3190 4470 -3150
rect 4510 -3190 4520 -3150
rect 4460 -3220 4520 -3190
rect 4460 -3260 4470 -3220
rect 4510 -3260 4520 -3220
rect 4460 -3290 4520 -3260
rect 4460 -3330 4470 -3290
rect 4510 -3330 4520 -3290
rect 4460 -3355 4520 -3330
rect 4460 -3395 4470 -3355
rect 4510 -3395 4520 -3355
rect 4460 -3415 4520 -3395
rect 4460 -3455 4470 -3415
rect 4510 -3455 4520 -3415
rect 4460 -3480 4520 -3455
rect 4460 -3520 4470 -3480
rect 4510 -3520 4520 -3480
rect 4460 -3550 4520 -3520
rect 4460 -3590 4470 -3550
rect 4510 -3590 4520 -3550
rect 4460 -3620 4520 -3590
rect 4460 -3660 4470 -3620
rect 4510 -3660 4520 -3620
rect 4460 -3690 4520 -3660
rect 4460 -3730 4470 -3690
rect 4510 -3730 4520 -3690
rect 4460 -3755 4520 -3730
rect 4460 -3795 4470 -3755
rect 4510 -3795 4520 -3755
rect 4460 -3815 4520 -3795
rect 4460 -3855 4470 -3815
rect 4510 -3855 4520 -3815
rect 4460 -3880 4520 -3855
rect 4460 -3920 4470 -3880
rect 4510 -3920 4520 -3880
rect 4460 -3950 4520 -3920
rect 4460 -3990 4470 -3950
rect 4510 -3990 4520 -3950
rect 4460 -4020 4520 -3990
rect 4460 -4060 4470 -4020
rect 4510 -4060 4520 -4020
rect 4460 -4090 4520 -4060
rect 4460 -4130 4470 -4090
rect 4510 -4130 4520 -4090
rect 4460 -4155 4520 -4130
rect 4460 -4195 4470 -4155
rect 4510 -4195 4520 -4155
rect 4460 -4215 4520 -4195
rect 4460 -4255 4470 -4215
rect 4510 -4255 4520 -4215
rect 4460 -4280 4520 -4255
rect 4460 -4320 4470 -4280
rect 4510 -4320 4520 -4280
rect 4460 -4350 4520 -4320
rect 4460 -4390 4470 -4350
rect 4510 -4390 4520 -4350
rect 4460 -4420 4520 -4390
rect 4460 -4460 4470 -4420
rect 4510 -4460 4520 -4420
rect 4460 -4490 4520 -4460
rect 4460 -4530 4470 -4490
rect 4510 -4530 4520 -4490
rect 4460 -4555 4520 -4530
rect 4460 -4595 4470 -4555
rect 4510 -4595 4520 -4555
rect 4460 -4605 4520 -4595
rect 4810 -3015 4870 -3005
rect 4810 -3055 4820 -3015
rect 4860 -3055 4870 -3015
rect 4810 -3080 4870 -3055
rect 4810 -3120 4820 -3080
rect 4860 -3120 4870 -3080
rect 4810 -3150 4870 -3120
rect 4810 -3190 4820 -3150
rect 4860 -3190 4870 -3150
rect 4810 -3220 4870 -3190
rect 4810 -3260 4820 -3220
rect 4860 -3260 4870 -3220
rect 4810 -3290 4870 -3260
rect 4810 -3330 4820 -3290
rect 4860 -3330 4870 -3290
rect 4810 -3355 4870 -3330
rect 4810 -3395 4820 -3355
rect 4860 -3395 4870 -3355
rect 4810 -3415 4870 -3395
rect 4810 -3455 4820 -3415
rect 4860 -3455 4870 -3415
rect 4810 -3480 4870 -3455
rect 4810 -3520 4820 -3480
rect 4860 -3520 4870 -3480
rect 4810 -3550 4870 -3520
rect 4810 -3590 4820 -3550
rect 4860 -3590 4870 -3550
rect 4810 -3620 4870 -3590
rect 4810 -3660 4820 -3620
rect 4860 -3660 4870 -3620
rect 4810 -3690 4870 -3660
rect 4810 -3730 4820 -3690
rect 4860 -3730 4870 -3690
rect 4810 -3755 4870 -3730
rect 4810 -3795 4820 -3755
rect 4860 -3795 4870 -3755
rect 4810 -3815 4870 -3795
rect 4810 -3855 4820 -3815
rect 4860 -3855 4870 -3815
rect 4810 -3880 4870 -3855
rect 4810 -3920 4820 -3880
rect 4860 -3920 4870 -3880
rect 4810 -3950 4870 -3920
rect 4810 -3990 4820 -3950
rect 4860 -3990 4870 -3950
rect 4810 -4020 4870 -3990
rect 4810 -4060 4820 -4020
rect 4860 -4060 4870 -4020
rect 4810 -4090 4870 -4060
rect 4810 -4130 4820 -4090
rect 4860 -4130 4870 -4090
rect 4810 -4155 4870 -4130
rect 4810 -4195 4820 -4155
rect 4860 -4195 4870 -4155
rect 4810 -4215 4870 -4195
rect 4810 -4255 4820 -4215
rect 4860 -4255 4870 -4215
rect 4810 -4280 4870 -4255
rect 4810 -4320 4820 -4280
rect 4860 -4320 4870 -4280
rect 4810 -4350 4870 -4320
rect 4810 -4390 4820 -4350
rect 4860 -4390 4870 -4350
rect 4810 -4420 4870 -4390
rect 4810 -4460 4820 -4420
rect 4860 -4460 4870 -4420
rect 4810 -4490 4870 -4460
rect 4810 -4530 4820 -4490
rect 4860 -4530 4870 -4490
rect 4810 -4555 4870 -4530
rect 4810 -4595 4820 -4555
rect 4860 -4595 4870 -4555
rect 4810 -4605 4870 -4595
rect 5160 -3015 5220 -3005
rect 5160 -3055 5170 -3015
rect 5210 -3055 5220 -3015
rect 5160 -3080 5220 -3055
rect 5160 -3120 5170 -3080
rect 5210 -3120 5220 -3080
rect 5160 -3150 5220 -3120
rect 5160 -3190 5170 -3150
rect 5210 -3190 5220 -3150
rect 5160 -3220 5220 -3190
rect 5160 -3260 5170 -3220
rect 5210 -3260 5220 -3220
rect 5160 -3290 5220 -3260
rect 5160 -3330 5170 -3290
rect 5210 -3330 5220 -3290
rect 5160 -3355 5220 -3330
rect 5160 -3395 5170 -3355
rect 5210 -3395 5220 -3355
rect 5160 -3415 5220 -3395
rect 5160 -3455 5170 -3415
rect 5210 -3455 5220 -3415
rect 5160 -3480 5220 -3455
rect 5160 -3520 5170 -3480
rect 5210 -3520 5220 -3480
rect 5160 -3550 5220 -3520
rect 5160 -3590 5170 -3550
rect 5210 -3590 5220 -3550
rect 5160 -3620 5220 -3590
rect 5160 -3660 5170 -3620
rect 5210 -3660 5220 -3620
rect 5160 -3690 5220 -3660
rect 5160 -3730 5170 -3690
rect 5210 -3730 5220 -3690
rect 5160 -3755 5220 -3730
rect 5160 -3795 5170 -3755
rect 5210 -3795 5220 -3755
rect 5160 -3815 5220 -3795
rect 5160 -3855 5170 -3815
rect 5210 -3855 5220 -3815
rect 5160 -3880 5220 -3855
rect 5160 -3920 5170 -3880
rect 5210 -3920 5220 -3880
rect 5160 -3950 5220 -3920
rect 5160 -3990 5170 -3950
rect 5210 -3990 5220 -3950
rect 5160 -4020 5220 -3990
rect 5160 -4060 5170 -4020
rect 5210 -4060 5220 -4020
rect 5160 -4090 5220 -4060
rect 5160 -4130 5170 -4090
rect 5210 -4130 5220 -4090
rect 5160 -4155 5220 -4130
rect 5160 -4195 5170 -4155
rect 5210 -4195 5220 -4155
rect 5160 -4215 5220 -4195
rect 5160 -4255 5170 -4215
rect 5210 -4255 5220 -4215
rect 5160 -4280 5220 -4255
rect 5160 -4320 5170 -4280
rect 5210 -4320 5220 -4280
rect 5160 -4350 5220 -4320
rect 5160 -4390 5170 -4350
rect 5210 -4390 5220 -4350
rect 5160 -4420 5220 -4390
rect 5160 -4460 5170 -4420
rect 5210 -4460 5220 -4420
rect 5160 -4490 5220 -4460
rect 5160 -4530 5170 -4490
rect 5210 -4530 5220 -4490
rect 5160 -4555 5220 -4530
rect 5160 -4595 5170 -4555
rect 5210 -4595 5220 -4555
rect 5160 -4605 5220 -4595
rect 5510 -3015 5570 -3005
rect 5510 -3055 5520 -3015
rect 5560 -3055 5570 -3015
rect 5510 -3080 5570 -3055
rect 5510 -3120 5520 -3080
rect 5560 -3120 5570 -3080
rect 5510 -3150 5570 -3120
rect 5510 -3190 5520 -3150
rect 5560 -3190 5570 -3150
rect 5510 -3220 5570 -3190
rect 5510 -3260 5520 -3220
rect 5560 -3260 5570 -3220
rect 5510 -3290 5570 -3260
rect 5510 -3330 5520 -3290
rect 5560 -3330 5570 -3290
rect 5510 -3355 5570 -3330
rect 5510 -3395 5520 -3355
rect 5560 -3395 5570 -3355
rect 5510 -3415 5570 -3395
rect 5510 -3455 5520 -3415
rect 5560 -3455 5570 -3415
rect 5510 -3480 5570 -3455
rect 5510 -3520 5520 -3480
rect 5560 -3520 5570 -3480
rect 5510 -3550 5570 -3520
rect 5510 -3590 5520 -3550
rect 5560 -3590 5570 -3550
rect 5510 -3620 5570 -3590
rect 5510 -3660 5520 -3620
rect 5560 -3660 5570 -3620
rect 5510 -3690 5570 -3660
rect 5510 -3730 5520 -3690
rect 5560 -3730 5570 -3690
rect 5510 -3755 5570 -3730
rect 5510 -3795 5520 -3755
rect 5560 -3795 5570 -3755
rect 5510 -3815 5570 -3795
rect 5510 -3855 5520 -3815
rect 5560 -3855 5570 -3815
rect 5510 -3880 5570 -3855
rect 5510 -3920 5520 -3880
rect 5560 -3920 5570 -3880
rect 5510 -3950 5570 -3920
rect 5510 -3990 5520 -3950
rect 5560 -3990 5570 -3950
rect 5510 -4020 5570 -3990
rect 5510 -4060 5520 -4020
rect 5560 -4060 5570 -4020
rect 5510 -4090 5570 -4060
rect 5510 -4130 5520 -4090
rect 5560 -4130 5570 -4090
rect 5510 -4155 5570 -4130
rect 5510 -4195 5520 -4155
rect 5560 -4195 5570 -4155
rect 5510 -4215 5570 -4195
rect 5510 -4255 5520 -4215
rect 5560 -4255 5570 -4215
rect 5510 -4280 5570 -4255
rect 5510 -4320 5520 -4280
rect 5560 -4320 5570 -4280
rect 5510 -4350 5570 -4320
rect 5510 -4390 5520 -4350
rect 5560 -4390 5570 -4350
rect 5510 -4420 5570 -4390
rect 5510 -4460 5520 -4420
rect 5560 -4460 5570 -4420
rect 5510 -4490 5570 -4460
rect 5510 -4530 5520 -4490
rect 5560 -4530 5570 -4490
rect 5510 -4555 5570 -4530
rect 5510 -4595 5520 -4555
rect 5560 -4595 5570 -4555
rect 5510 -4605 5570 -4595
<< via3 >>
rect 2110 19310 2150 19315
rect 2110 19280 2115 19310
rect 2115 19280 2145 19310
rect 2145 19280 2150 19310
rect 2110 19275 2150 19280
rect 2110 19245 2150 19250
rect 2110 19215 2115 19245
rect 2115 19215 2145 19245
rect 2145 19215 2150 19245
rect 2110 19210 2150 19215
rect 2110 19175 2150 19180
rect 2110 19145 2115 19175
rect 2115 19145 2145 19175
rect 2145 19145 2150 19175
rect 2110 19140 2150 19145
rect 2110 19105 2150 19110
rect 2110 19075 2115 19105
rect 2115 19075 2145 19105
rect 2145 19075 2150 19105
rect 2110 19070 2150 19075
rect 2110 19035 2150 19040
rect 2110 19005 2115 19035
rect 2115 19005 2145 19035
rect 2145 19005 2150 19035
rect 2110 19000 2150 19005
rect 2110 18970 2150 18975
rect 2110 18940 2115 18970
rect 2115 18940 2145 18970
rect 2145 18940 2150 18970
rect 2110 18935 2150 18940
rect 2110 18910 2150 18915
rect 2110 18880 2115 18910
rect 2115 18880 2145 18910
rect 2145 18880 2150 18910
rect 2110 18875 2150 18880
rect 2110 18845 2150 18850
rect 2110 18815 2115 18845
rect 2115 18815 2145 18845
rect 2145 18815 2150 18845
rect 2110 18810 2150 18815
rect 2110 18775 2150 18780
rect 2110 18745 2115 18775
rect 2115 18745 2145 18775
rect 2145 18745 2150 18775
rect 2110 18740 2150 18745
rect 2110 18705 2150 18710
rect 2110 18675 2115 18705
rect 2115 18675 2145 18705
rect 2145 18675 2150 18705
rect 2110 18670 2150 18675
rect 2110 18635 2150 18640
rect 2110 18605 2115 18635
rect 2115 18605 2145 18635
rect 2145 18605 2150 18635
rect 2110 18600 2150 18605
rect 2110 18570 2150 18575
rect 2110 18540 2115 18570
rect 2115 18540 2145 18570
rect 2145 18540 2150 18570
rect 2110 18535 2150 18540
rect 2110 18510 2150 18515
rect 2110 18480 2115 18510
rect 2115 18480 2145 18510
rect 2145 18480 2150 18510
rect 2110 18475 2150 18480
rect 2110 18445 2150 18450
rect 2110 18415 2115 18445
rect 2115 18415 2145 18445
rect 2145 18415 2150 18445
rect 2110 18410 2150 18415
rect 2110 18375 2150 18380
rect 2110 18345 2115 18375
rect 2115 18345 2145 18375
rect 2145 18345 2150 18375
rect 2110 18340 2150 18345
rect 2110 18305 2150 18310
rect 2110 18275 2115 18305
rect 2115 18275 2145 18305
rect 2145 18275 2150 18305
rect 2110 18270 2150 18275
rect 2110 18235 2150 18240
rect 2110 18205 2115 18235
rect 2115 18205 2145 18235
rect 2145 18205 2150 18235
rect 2110 18200 2150 18205
rect 2110 18170 2150 18175
rect 2110 18140 2115 18170
rect 2115 18140 2145 18170
rect 2145 18140 2150 18170
rect 2110 18135 2150 18140
rect 2110 18110 2150 18115
rect 2110 18080 2115 18110
rect 2115 18080 2145 18110
rect 2145 18080 2150 18110
rect 2110 18075 2150 18080
rect 2110 18045 2150 18050
rect 2110 18015 2115 18045
rect 2115 18015 2145 18045
rect 2145 18015 2150 18045
rect 2110 18010 2150 18015
rect 2110 17975 2150 17980
rect 2110 17945 2115 17975
rect 2115 17945 2145 17975
rect 2145 17945 2150 17975
rect 2110 17940 2150 17945
rect 2110 17905 2150 17910
rect 2110 17875 2115 17905
rect 2115 17875 2145 17905
rect 2145 17875 2150 17905
rect 2110 17870 2150 17875
rect 2110 17835 2150 17840
rect 2110 17805 2115 17835
rect 2115 17805 2145 17835
rect 2145 17805 2150 17835
rect 2110 17800 2150 17805
rect 2110 17770 2150 17775
rect 2110 17740 2115 17770
rect 2115 17740 2145 17770
rect 2145 17740 2150 17770
rect 2110 17735 2150 17740
rect 6700 19310 6740 19315
rect 6700 19280 6705 19310
rect 6705 19280 6735 19310
rect 6735 19280 6740 19310
rect 6700 19275 6740 19280
rect 6700 19245 6740 19250
rect 6700 19215 6705 19245
rect 6705 19215 6735 19245
rect 6735 19215 6740 19245
rect 6700 19210 6740 19215
rect 6700 19175 6740 19180
rect 6700 19145 6705 19175
rect 6705 19145 6735 19175
rect 6735 19145 6740 19175
rect 6700 19140 6740 19145
rect 6700 19105 6740 19110
rect 6700 19075 6705 19105
rect 6705 19075 6735 19105
rect 6735 19075 6740 19105
rect 6700 19070 6740 19075
rect 6700 19035 6740 19040
rect 6700 19005 6705 19035
rect 6705 19005 6735 19035
rect 6735 19005 6740 19035
rect 6700 19000 6740 19005
rect 6700 18970 6740 18975
rect 6700 18940 6705 18970
rect 6705 18940 6735 18970
rect 6735 18940 6740 18970
rect 6700 18935 6740 18940
rect 6700 18910 6740 18915
rect 6700 18880 6705 18910
rect 6705 18880 6735 18910
rect 6735 18880 6740 18910
rect 6700 18875 6740 18880
rect 6700 18845 6740 18850
rect 6700 18815 6705 18845
rect 6705 18815 6735 18845
rect 6735 18815 6740 18845
rect 6700 18810 6740 18815
rect 6700 18775 6740 18780
rect 6700 18745 6705 18775
rect 6705 18745 6735 18775
rect 6735 18745 6740 18775
rect 6700 18740 6740 18745
rect 6700 18705 6740 18710
rect 6700 18675 6705 18705
rect 6705 18675 6735 18705
rect 6735 18675 6740 18705
rect 6700 18670 6740 18675
rect 6700 18635 6740 18640
rect 6700 18605 6705 18635
rect 6705 18605 6735 18635
rect 6735 18605 6740 18635
rect 6700 18600 6740 18605
rect 6700 18570 6740 18575
rect 6700 18540 6705 18570
rect 6705 18540 6735 18570
rect 6735 18540 6740 18570
rect 6700 18535 6740 18540
rect 6700 18510 6740 18515
rect 6700 18480 6705 18510
rect 6705 18480 6735 18510
rect 6735 18480 6740 18510
rect 6700 18475 6740 18480
rect 6700 18445 6740 18450
rect 6700 18415 6705 18445
rect 6705 18415 6735 18445
rect 6735 18415 6740 18445
rect 6700 18410 6740 18415
rect 6700 18375 6740 18380
rect 6700 18345 6705 18375
rect 6705 18345 6735 18375
rect 6735 18345 6740 18375
rect 6700 18340 6740 18345
rect 6700 18305 6740 18310
rect 6700 18275 6705 18305
rect 6705 18275 6735 18305
rect 6735 18275 6740 18305
rect 6700 18270 6740 18275
rect 6700 18235 6740 18240
rect 6700 18205 6705 18235
rect 6705 18205 6735 18235
rect 6735 18205 6740 18235
rect 6700 18200 6740 18205
rect 6700 18170 6740 18175
rect 6700 18140 6705 18170
rect 6705 18140 6735 18170
rect 6735 18140 6740 18170
rect 6700 18135 6740 18140
rect 6700 18110 6740 18115
rect 6700 18080 6705 18110
rect 6705 18080 6735 18110
rect 6735 18080 6740 18110
rect 6700 18075 6740 18080
rect 6700 18045 6740 18050
rect 6700 18015 6705 18045
rect 6705 18015 6735 18045
rect 6735 18015 6740 18045
rect 6700 18010 6740 18015
rect 6700 17975 6740 17980
rect 6700 17945 6705 17975
rect 6705 17945 6735 17975
rect 6735 17945 6740 17975
rect 6700 17940 6740 17945
rect 6700 17905 6740 17910
rect 6700 17875 6705 17905
rect 6705 17875 6735 17905
rect 6735 17875 6740 17905
rect 6700 17870 6740 17875
rect 6700 17835 6740 17840
rect 6700 17805 6705 17835
rect 6705 17805 6735 17835
rect 6735 17805 6740 17835
rect 6700 17800 6740 17805
rect 6700 17770 6740 17775
rect 6700 17740 6705 17770
rect 6705 17740 6735 17770
rect 6735 17740 6740 17770
rect 6700 17735 6740 17740
rect 31305 19270 31340 19305
rect 31350 19270 31385 19305
rect 31395 19270 31430 19305
rect 31440 19270 31475 19305
rect 31485 19270 31520 19305
rect 31530 19270 31565 19305
rect 31575 19270 31610 19305
rect 31620 19270 31655 19305
rect 31665 19270 31700 19305
rect 31710 19270 31745 19305
rect 31755 19270 31790 19305
rect 31800 19270 31835 19305
rect 31845 19270 31880 19305
rect 31890 19270 31925 19305
rect 31935 19270 31970 19305
rect 31980 19270 32015 19305
rect 32025 19270 32060 19305
rect 32070 19270 32105 19305
rect 32115 19270 32150 19305
rect 32160 19270 32195 19305
rect 32205 19270 32240 19305
rect 32250 19270 32285 19305
rect 32295 19270 32330 19305
rect 32340 19270 32375 19305
rect 32385 19270 32420 19305
rect 32430 19270 32465 19305
rect 32475 19270 32510 19305
rect 32520 19270 32555 19305
rect 32565 19270 32600 19305
rect 32610 19270 32645 19305
rect 32655 19270 32690 19305
rect 32700 19270 32735 19305
rect 32745 19270 32780 19305
rect 32790 19270 32825 19305
rect 32835 19270 32870 19305
rect 31305 19225 31340 19260
rect 31350 19225 31385 19260
rect 31395 19225 31430 19260
rect 31440 19225 31475 19260
rect 31485 19225 31520 19260
rect 31530 19225 31565 19260
rect 31575 19225 31610 19260
rect 31620 19225 31655 19260
rect 31665 19225 31700 19260
rect 31710 19225 31745 19260
rect 31755 19225 31790 19260
rect 31800 19225 31835 19260
rect 31845 19225 31880 19260
rect 31890 19225 31925 19260
rect 31935 19225 31970 19260
rect 31980 19225 32015 19260
rect 32025 19225 32060 19260
rect 32070 19225 32105 19260
rect 32115 19225 32150 19260
rect 32160 19225 32195 19260
rect 32205 19225 32240 19260
rect 32250 19225 32285 19260
rect 32295 19225 32330 19260
rect 32340 19225 32375 19260
rect 32385 19225 32420 19260
rect 32430 19225 32465 19260
rect 32475 19225 32510 19260
rect 32520 19225 32555 19260
rect 32565 19225 32600 19260
rect 32610 19225 32645 19260
rect 32655 19225 32690 19260
rect 32700 19225 32735 19260
rect 32745 19225 32780 19260
rect 32790 19225 32825 19260
rect 32835 19225 32870 19260
rect 31305 19180 31340 19215
rect 31350 19180 31385 19215
rect 31395 19180 31430 19215
rect 31440 19180 31475 19215
rect 31485 19180 31520 19215
rect 31530 19180 31565 19215
rect 31575 19180 31610 19215
rect 31620 19180 31655 19215
rect 31665 19180 31700 19215
rect 31710 19180 31745 19215
rect 31755 19180 31790 19215
rect 31800 19180 31835 19215
rect 31845 19180 31880 19215
rect 31890 19180 31925 19215
rect 31935 19180 31970 19215
rect 31980 19180 32015 19215
rect 32025 19180 32060 19215
rect 32070 19180 32105 19215
rect 32115 19180 32150 19215
rect 32160 19180 32195 19215
rect 32205 19180 32240 19215
rect 32250 19180 32285 19215
rect 32295 19180 32330 19215
rect 32340 19180 32375 19215
rect 32385 19180 32420 19215
rect 32430 19180 32465 19215
rect 32475 19180 32510 19215
rect 32520 19180 32555 19215
rect 32565 19180 32600 19215
rect 32610 19180 32645 19215
rect 32655 19180 32690 19215
rect 32700 19180 32735 19215
rect 32745 19180 32780 19215
rect 32790 19180 32825 19215
rect 32835 19180 32870 19215
rect 31305 19135 31340 19170
rect 31350 19135 31385 19170
rect 31395 19135 31430 19170
rect 31440 19135 31475 19170
rect 31485 19135 31520 19170
rect 31530 19135 31565 19170
rect 31575 19135 31610 19170
rect 31620 19135 31655 19170
rect 31665 19135 31700 19170
rect 31710 19135 31745 19170
rect 31755 19135 31790 19170
rect 31800 19135 31835 19170
rect 31845 19135 31880 19170
rect 31890 19135 31925 19170
rect 31935 19135 31970 19170
rect 31980 19135 32015 19170
rect 32025 19135 32060 19170
rect 32070 19135 32105 19170
rect 32115 19135 32150 19170
rect 32160 19135 32195 19170
rect 32205 19135 32240 19170
rect 32250 19135 32285 19170
rect 32295 19135 32330 19170
rect 32340 19135 32375 19170
rect 32385 19135 32420 19170
rect 32430 19135 32465 19170
rect 32475 19135 32510 19170
rect 32520 19135 32555 19170
rect 32565 19135 32600 19170
rect 32610 19135 32645 19170
rect 32655 19135 32690 19170
rect 32700 19135 32735 19170
rect 32745 19135 32780 19170
rect 32790 19135 32825 19170
rect 32835 19135 32870 19170
rect 31305 19090 31340 19125
rect 31350 19090 31385 19125
rect 31395 19090 31430 19125
rect 31440 19090 31475 19125
rect 31485 19090 31520 19125
rect 31530 19090 31565 19125
rect 31575 19090 31610 19125
rect 31620 19090 31655 19125
rect 31665 19090 31700 19125
rect 31710 19090 31745 19125
rect 31755 19090 31790 19125
rect 31800 19090 31835 19125
rect 31845 19090 31880 19125
rect 31890 19090 31925 19125
rect 31935 19090 31970 19125
rect 31980 19090 32015 19125
rect 32025 19090 32060 19125
rect 32070 19090 32105 19125
rect 32115 19090 32150 19125
rect 32160 19090 32195 19125
rect 32205 19090 32240 19125
rect 32250 19090 32285 19125
rect 32295 19090 32330 19125
rect 32340 19090 32375 19125
rect 32385 19090 32420 19125
rect 32430 19090 32465 19125
rect 32475 19090 32510 19125
rect 32520 19090 32555 19125
rect 32565 19090 32600 19125
rect 32610 19090 32645 19125
rect 32655 19090 32690 19125
rect 32700 19090 32735 19125
rect 32745 19090 32780 19125
rect 32790 19090 32825 19125
rect 32835 19090 32870 19125
rect 31305 19045 31340 19080
rect 31350 19045 31385 19080
rect 31395 19045 31430 19080
rect 31440 19045 31475 19080
rect 31485 19045 31520 19080
rect 31530 19045 31565 19080
rect 31575 19045 31610 19080
rect 31620 19045 31655 19080
rect 31665 19045 31700 19080
rect 31710 19045 31745 19080
rect 31755 19045 31790 19080
rect 31800 19045 31835 19080
rect 31845 19045 31880 19080
rect 31890 19045 31925 19080
rect 31935 19045 31970 19080
rect 31980 19045 32015 19080
rect 32025 19045 32060 19080
rect 32070 19045 32105 19080
rect 32115 19045 32150 19080
rect 32160 19045 32195 19080
rect 32205 19045 32240 19080
rect 32250 19045 32285 19080
rect 32295 19045 32330 19080
rect 32340 19045 32375 19080
rect 32385 19045 32420 19080
rect 32430 19045 32465 19080
rect 32475 19045 32510 19080
rect 32520 19045 32555 19080
rect 32565 19045 32600 19080
rect 32610 19045 32645 19080
rect 32655 19045 32690 19080
rect 32700 19045 32735 19080
rect 32745 19045 32780 19080
rect 32790 19045 32825 19080
rect 32835 19045 32870 19080
rect 31305 19000 31340 19035
rect 31350 19000 31385 19035
rect 31395 19000 31430 19035
rect 31440 19000 31475 19035
rect 31485 19000 31520 19035
rect 31530 19000 31565 19035
rect 31575 19000 31610 19035
rect 31620 19000 31655 19035
rect 31665 19000 31700 19035
rect 31710 19000 31745 19035
rect 31755 19000 31790 19035
rect 31800 19000 31835 19035
rect 31845 19000 31880 19035
rect 31890 19000 31925 19035
rect 31935 19000 31970 19035
rect 31980 19000 32015 19035
rect 32025 19000 32060 19035
rect 32070 19000 32105 19035
rect 32115 19000 32150 19035
rect 32160 19000 32195 19035
rect 32205 19000 32240 19035
rect 32250 19000 32285 19035
rect 32295 19000 32330 19035
rect 32340 19000 32375 19035
rect 32385 19000 32420 19035
rect 32430 19000 32465 19035
rect 32475 19000 32510 19035
rect 32520 19000 32555 19035
rect 32565 19000 32600 19035
rect 32610 19000 32645 19035
rect 32655 19000 32690 19035
rect 32700 19000 32735 19035
rect 32745 19000 32780 19035
rect 32790 19000 32825 19035
rect 32835 19000 32870 19035
rect 31305 18955 31340 18990
rect 31350 18955 31385 18990
rect 31395 18955 31430 18990
rect 31440 18955 31475 18990
rect 31485 18955 31520 18990
rect 31530 18955 31565 18990
rect 31575 18955 31610 18990
rect 31620 18955 31655 18990
rect 31665 18955 31700 18990
rect 31710 18955 31745 18990
rect 31755 18955 31790 18990
rect 31800 18955 31835 18990
rect 31845 18955 31880 18990
rect 31890 18955 31925 18990
rect 31935 18955 31970 18990
rect 31980 18955 32015 18990
rect 32025 18955 32060 18990
rect 32070 18955 32105 18990
rect 32115 18955 32150 18990
rect 32160 18955 32195 18990
rect 32205 18955 32240 18990
rect 32250 18955 32285 18990
rect 32295 18955 32330 18990
rect 32340 18955 32375 18990
rect 32385 18955 32420 18990
rect 32430 18955 32465 18990
rect 32475 18955 32510 18990
rect 32520 18955 32555 18990
rect 32565 18955 32600 18990
rect 32610 18955 32645 18990
rect 32655 18955 32690 18990
rect 32700 18955 32735 18990
rect 32745 18955 32780 18990
rect 32790 18955 32825 18990
rect 32835 18955 32870 18990
rect 31305 18910 31340 18945
rect 31350 18910 31385 18945
rect 31395 18910 31430 18945
rect 31440 18910 31475 18945
rect 31485 18910 31520 18945
rect 31530 18910 31565 18945
rect 31575 18910 31610 18945
rect 31620 18910 31655 18945
rect 31665 18910 31700 18945
rect 31710 18910 31745 18945
rect 31755 18910 31790 18945
rect 31800 18910 31835 18945
rect 31845 18910 31880 18945
rect 31890 18910 31925 18945
rect 31935 18910 31970 18945
rect 31980 18910 32015 18945
rect 32025 18910 32060 18945
rect 32070 18910 32105 18945
rect 32115 18910 32150 18945
rect 32160 18910 32195 18945
rect 32205 18910 32240 18945
rect 32250 18910 32285 18945
rect 32295 18910 32330 18945
rect 32340 18910 32375 18945
rect 32385 18910 32420 18945
rect 32430 18910 32465 18945
rect 32475 18910 32510 18945
rect 32520 18910 32555 18945
rect 32565 18910 32600 18945
rect 32610 18910 32645 18945
rect 32655 18910 32690 18945
rect 32700 18910 32735 18945
rect 32745 18910 32780 18945
rect 32790 18910 32825 18945
rect 32835 18910 32870 18945
rect 31305 18865 31340 18900
rect 31350 18865 31385 18900
rect 31395 18865 31430 18900
rect 31440 18865 31475 18900
rect 31485 18865 31520 18900
rect 31530 18865 31565 18900
rect 31575 18865 31610 18900
rect 31620 18865 31655 18900
rect 31665 18865 31700 18900
rect 31710 18865 31745 18900
rect 31755 18865 31790 18900
rect 31800 18865 31835 18900
rect 31845 18865 31880 18900
rect 31890 18865 31925 18900
rect 31935 18865 31970 18900
rect 31980 18865 32015 18900
rect 32025 18865 32060 18900
rect 32070 18865 32105 18900
rect 32115 18865 32150 18900
rect 32160 18865 32195 18900
rect 32205 18865 32240 18900
rect 32250 18865 32285 18900
rect 32295 18865 32330 18900
rect 32340 18865 32375 18900
rect 32385 18865 32420 18900
rect 32430 18865 32465 18900
rect 32475 18865 32510 18900
rect 32520 18865 32555 18900
rect 32565 18865 32600 18900
rect 32610 18865 32645 18900
rect 32655 18865 32690 18900
rect 32700 18865 32735 18900
rect 32745 18865 32780 18900
rect 32790 18865 32825 18900
rect 32835 18865 32870 18900
rect 31305 18820 31340 18855
rect 31350 18820 31385 18855
rect 31395 18820 31430 18855
rect 31440 18820 31475 18855
rect 31485 18820 31520 18855
rect 31530 18820 31565 18855
rect 31575 18820 31610 18855
rect 31620 18820 31655 18855
rect 31665 18820 31700 18855
rect 31710 18820 31745 18855
rect 31755 18820 31790 18855
rect 31800 18820 31835 18855
rect 31845 18820 31880 18855
rect 31890 18820 31925 18855
rect 31935 18820 31970 18855
rect 31980 18820 32015 18855
rect 32025 18820 32060 18855
rect 32070 18820 32105 18855
rect 32115 18820 32150 18855
rect 32160 18820 32195 18855
rect 32205 18820 32240 18855
rect 32250 18820 32285 18855
rect 32295 18820 32330 18855
rect 32340 18820 32375 18855
rect 32385 18820 32420 18855
rect 32430 18820 32465 18855
rect 32475 18820 32510 18855
rect 32520 18820 32555 18855
rect 32565 18820 32600 18855
rect 32610 18820 32645 18855
rect 32655 18820 32690 18855
rect 32700 18820 32735 18855
rect 32745 18820 32780 18855
rect 32790 18820 32825 18855
rect 32835 18820 32870 18855
rect 31305 18775 31340 18810
rect 31350 18775 31385 18810
rect 31395 18775 31430 18810
rect 31440 18775 31475 18810
rect 31485 18775 31520 18810
rect 31530 18775 31565 18810
rect 31575 18775 31610 18810
rect 31620 18775 31655 18810
rect 31665 18775 31700 18810
rect 31710 18775 31745 18810
rect 31755 18775 31790 18810
rect 31800 18775 31835 18810
rect 31845 18775 31880 18810
rect 31890 18775 31925 18810
rect 31935 18775 31970 18810
rect 31980 18775 32015 18810
rect 32025 18775 32060 18810
rect 32070 18775 32105 18810
rect 32115 18775 32150 18810
rect 32160 18775 32195 18810
rect 32205 18775 32240 18810
rect 32250 18775 32285 18810
rect 32295 18775 32330 18810
rect 32340 18775 32375 18810
rect 32385 18775 32420 18810
rect 32430 18775 32465 18810
rect 32475 18775 32510 18810
rect 32520 18775 32555 18810
rect 32565 18775 32600 18810
rect 32610 18775 32645 18810
rect 32655 18775 32690 18810
rect 32700 18775 32735 18810
rect 32745 18775 32780 18810
rect 32790 18775 32825 18810
rect 32835 18775 32870 18810
rect 31305 18730 31340 18765
rect 31350 18730 31385 18765
rect 31395 18730 31430 18765
rect 31440 18730 31475 18765
rect 31485 18730 31520 18765
rect 31530 18730 31565 18765
rect 31575 18730 31610 18765
rect 31620 18730 31655 18765
rect 31665 18730 31700 18765
rect 31710 18730 31745 18765
rect 31755 18730 31790 18765
rect 31800 18730 31835 18765
rect 31845 18730 31880 18765
rect 31890 18730 31925 18765
rect 31935 18730 31970 18765
rect 31980 18730 32015 18765
rect 32025 18730 32060 18765
rect 32070 18730 32105 18765
rect 32115 18730 32150 18765
rect 32160 18730 32195 18765
rect 32205 18730 32240 18765
rect 32250 18730 32285 18765
rect 32295 18730 32330 18765
rect 32340 18730 32375 18765
rect 32385 18730 32420 18765
rect 32430 18730 32465 18765
rect 32475 18730 32510 18765
rect 32520 18730 32555 18765
rect 32565 18730 32600 18765
rect 32610 18730 32645 18765
rect 32655 18730 32690 18765
rect 32700 18730 32735 18765
rect 32745 18730 32780 18765
rect 32790 18730 32825 18765
rect 32835 18730 32870 18765
rect 31305 18685 31340 18720
rect 31350 18685 31385 18720
rect 31395 18685 31430 18720
rect 31440 18685 31475 18720
rect 31485 18685 31520 18720
rect 31530 18685 31565 18720
rect 31575 18685 31610 18720
rect 31620 18685 31655 18720
rect 31665 18685 31700 18720
rect 31710 18685 31745 18720
rect 31755 18685 31790 18720
rect 31800 18685 31835 18720
rect 31845 18685 31880 18720
rect 31890 18685 31925 18720
rect 31935 18685 31970 18720
rect 31980 18685 32015 18720
rect 32025 18685 32060 18720
rect 32070 18685 32105 18720
rect 32115 18685 32150 18720
rect 32160 18685 32195 18720
rect 32205 18685 32240 18720
rect 32250 18685 32285 18720
rect 32295 18685 32330 18720
rect 32340 18685 32375 18720
rect 32385 18685 32420 18720
rect 32430 18685 32465 18720
rect 32475 18685 32510 18720
rect 32520 18685 32555 18720
rect 32565 18685 32600 18720
rect 32610 18685 32645 18720
rect 32655 18685 32690 18720
rect 32700 18685 32735 18720
rect 32745 18685 32780 18720
rect 32790 18685 32825 18720
rect 32835 18685 32870 18720
rect 31305 18640 31340 18675
rect 31350 18640 31385 18675
rect 31395 18640 31430 18675
rect 31440 18640 31475 18675
rect 31485 18640 31520 18675
rect 31530 18640 31565 18675
rect 31575 18640 31610 18675
rect 31620 18640 31655 18675
rect 31665 18640 31700 18675
rect 31710 18640 31745 18675
rect 31755 18640 31790 18675
rect 31800 18640 31835 18675
rect 31845 18640 31880 18675
rect 31890 18640 31925 18675
rect 31935 18640 31970 18675
rect 31980 18640 32015 18675
rect 32025 18640 32060 18675
rect 32070 18640 32105 18675
rect 32115 18640 32150 18675
rect 32160 18640 32195 18675
rect 32205 18640 32240 18675
rect 32250 18640 32285 18675
rect 32295 18640 32330 18675
rect 32340 18640 32375 18675
rect 32385 18640 32420 18675
rect 32430 18640 32465 18675
rect 32475 18640 32510 18675
rect 32520 18640 32555 18675
rect 32565 18640 32600 18675
rect 32610 18640 32645 18675
rect 32655 18640 32690 18675
rect 32700 18640 32735 18675
rect 32745 18640 32780 18675
rect 32790 18640 32825 18675
rect 32835 18640 32870 18675
rect 31305 18595 31340 18630
rect 31350 18595 31385 18630
rect 31395 18595 31430 18630
rect 31440 18595 31475 18630
rect 31485 18595 31520 18630
rect 31530 18595 31565 18630
rect 31575 18595 31610 18630
rect 31620 18595 31655 18630
rect 31665 18595 31700 18630
rect 31710 18595 31745 18630
rect 31755 18595 31790 18630
rect 31800 18595 31835 18630
rect 31845 18595 31880 18630
rect 31890 18595 31925 18630
rect 31935 18595 31970 18630
rect 31980 18595 32015 18630
rect 32025 18595 32060 18630
rect 32070 18595 32105 18630
rect 32115 18595 32150 18630
rect 32160 18595 32195 18630
rect 32205 18595 32240 18630
rect 32250 18595 32285 18630
rect 32295 18595 32330 18630
rect 32340 18595 32375 18630
rect 32385 18595 32420 18630
rect 32430 18595 32465 18630
rect 32475 18595 32510 18630
rect 32520 18595 32555 18630
rect 32565 18595 32600 18630
rect 32610 18595 32645 18630
rect 32655 18595 32690 18630
rect 32700 18595 32735 18630
rect 32745 18595 32780 18630
rect 32790 18595 32825 18630
rect 32835 18595 32870 18630
rect 31305 18550 31340 18585
rect 31350 18550 31385 18585
rect 31395 18550 31430 18585
rect 31440 18550 31475 18585
rect 31485 18550 31520 18585
rect 31530 18550 31565 18585
rect 31575 18550 31610 18585
rect 31620 18550 31655 18585
rect 31665 18550 31700 18585
rect 31710 18550 31745 18585
rect 31755 18550 31790 18585
rect 31800 18550 31835 18585
rect 31845 18550 31880 18585
rect 31890 18550 31925 18585
rect 31935 18550 31970 18585
rect 31980 18550 32015 18585
rect 32025 18550 32060 18585
rect 32070 18550 32105 18585
rect 32115 18550 32150 18585
rect 32160 18550 32195 18585
rect 32205 18550 32240 18585
rect 32250 18550 32285 18585
rect 32295 18550 32330 18585
rect 32340 18550 32375 18585
rect 32385 18550 32420 18585
rect 32430 18550 32465 18585
rect 32475 18550 32510 18585
rect 32520 18550 32555 18585
rect 32565 18550 32600 18585
rect 32610 18550 32645 18585
rect 32655 18550 32690 18585
rect 32700 18550 32735 18585
rect 32745 18550 32780 18585
rect 32790 18550 32825 18585
rect 32835 18550 32870 18585
rect 31305 18505 31340 18540
rect 31350 18505 31385 18540
rect 31395 18505 31430 18540
rect 31440 18505 31475 18540
rect 31485 18505 31520 18540
rect 31530 18505 31565 18540
rect 31575 18505 31610 18540
rect 31620 18505 31655 18540
rect 31665 18505 31700 18540
rect 31710 18505 31745 18540
rect 31755 18505 31790 18540
rect 31800 18505 31835 18540
rect 31845 18505 31880 18540
rect 31890 18505 31925 18540
rect 31935 18505 31970 18540
rect 31980 18505 32015 18540
rect 32025 18505 32060 18540
rect 32070 18505 32105 18540
rect 32115 18505 32150 18540
rect 32160 18505 32195 18540
rect 32205 18505 32240 18540
rect 32250 18505 32285 18540
rect 32295 18505 32330 18540
rect 32340 18505 32375 18540
rect 32385 18505 32420 18540
rect 32430 18505 32465 18540
rect 32475 18505 32510 18540
rect 32520 18505 32555 18540
rect 32565 18505 32600 18540
rect 32610 18505 32645 18540
rect 32655 18505 32690 18540
rect 32700 18505 32735 18540
rect 32745 18505 32780 18540
rect 32790 18505 32825 18540
rect 32835 18505 32870 18540
rect 31305 18460 31340 18495
rect 31350 18460 31385 18495
rect 31395 18460 31430 18495
rect 31440 18460 31475 18495
rect 31485 18460 31520 18495
rect 31530 18460 31565 18495
rect 31575 18460 31610 18495
rect 31620 18460 31655 18495
rect 31665 18460 31700 18495
rect 31710 18460 31745 18495
rect 31755 18460 31790 18495
rect 31800 18460 31835 18495
rect 31845 18460 31880 18495
rect 31890 18460 31925 18495
rect 31935 18460 31970 18495
rect 31980 18460 32015 18495
rect 32025 18460 32060 18495
rect 32070 18460 32105 18495
rect 32115 18460 32150 18495
rect 32160 18460 32195 18495
rect 32205 18460 32240 18495
rect 32250 18460 32285 18495
rect 32295 18460 32330 18495
rect 32340 18460 32375 18495
rect 32385 18460 32420 18495
rect 32430 18460 32465 18495
rect 32475 18460 32510 18495
rect 32520 18460 32555 18495
rect 32565 18460 32600 18495
rect 32610 18460 32645 18495
rect 32655 18460 32690 18495
rect 32700 18460 32735 18495
rect 32745 18460 32780 18495
rect 32790 18460 32825 18495
rect 32835 18460 32870 18495
rect 31305 18415 31340 18450
rect 31350 18415 31385 18450
rect 31395 18415 31430 18450
rect 31440 18415 31475 18450
rect 31485 18415 31520 18450
rect 31530 18415 31565 18450
rect 31575 18415 31610 18450
rect 31620 18415 31655 18450
rect 31665 18415 31700 18450
rect 31710 18415 31745 18450
rect 31755 18415 31790 18450
rect 31800 18415 31835 18450
rect 31845 18415 31880 18450
rect 31890 18415 31925 18450
rect 31935 18415 31970 18450
rect 31980 18415 32015 18450
rect 32025 18415 32060 18450
rect 32070 18415 32105 18450
rect 32115 18415 32150 18450
rect 32160 18415 32195 18450
rect 32205 18415 32240 18450
rect 32250 18415 32285 18450
rect 32295 18415 32330 18450
rect 32340 18415 32375 18450
rect 32385 18415 32420 18450
rect 32430 18415 32465 18450
rect 32475 18415 32510 18450
rect 32520 18415 32555 18450
rect 32565 18415 32600 18450
rect 32610 18415 32645 18450
rect 32655 18415 32690 18450
rect 32700 18415 32735 18450
rect 32745 18415 32780 18450
rect 32790 18415 32825 18450
rect 32835 18415 32870 18450
rect 31305 18370 31340 18405
rect 31350 18370 31385 18405
rect 31395 18370 31430 18405
rect 31440 18370 31475 18405
rect 31485 18370 31520 18405
rect 31530 18370 31565 18405
rect 31575 18370 31610 18405
rect 31620 18370 31655 18405
rect 31665 18370 31700 18405
rect 31710 18370 31745 18405
rect 31755 18370 31790 18405
rect 31800 18370 31835 18405
rect 31845 18370 31880 18405
rect 31890 18370 31925 18405
rect 31935 18370 31970 18405
rect 31980 18370 32015 18405
rect 32025 18370 32060 18405
rect 32070 18370 32105 18405
rect 32115 18370 32150 18405
rect 32160 18370 32195 18405
rect 32205 18370 32240 18405
rect 32250 18370 32285 18405
rect 32295 18370 32330 18405
rect 32340 18370 32375 18405
rect 32385 18370 32420 18405
rect 32430 18370 32465 18405
rect 32475 18370 32510 18405
rect 32520 18370 32555 18405
rect 32565 18370 32600 18405
rect 32610 18370 32645 18405
rect 32655 18370 32690 18405
rect 32700 18370 32735 18405
rect 32745 18370 32780 18405
rect 32790 18370 32825 18405
rect 32835 18370 32870 18405
rect 31305 18325 31340 18360
rect 31350 18325 31385 18360
rect 31395 18325 31430 18360
rect 31440 18325 31475 18360
rect 31485 18325 31520 18360
rect 31530 18325 31565 18360
rect 31575 18325 31610 18360
rect 31620 18325 31655 18360
rect 31665 18325 31700 18360
rect 31710 18325 31745 18360
rect 31755 18325 31790 18360
rect 31800 18325 31835 18360
rect 31845 18325 31880 18360
rect 31890 18325 31925 18360
rect 31935 18325 31970 18360
rect 31980 18325 32015 18360
rect 32025 18325 32060 18360
rect 32070 18325 32105 18360
rect 32115 18325 32150 18360
rect 32160 18325 32195 18360
rect 32205 18325 32240 18360
rect 32250 18325 32285 18360
rect 32295 18325 32330 18360
rect 32340 18325 32375 18360
rect 32385 18325 32420 18360
rect 32430 18325 32465 18360
rect 32475 18325 32510 18360
rect 32520 18325 32555 18360
rect 32565 18325 32600 18360
rect 32610 18325 32645 18360
rect 32655 18325 32690 18360
rect 32700 18325 32735 18360
rect 32745 18325 32780 18360
rect 32790 18325 32825 18360
rect 32835 18325 32870 18360
rect 31305 18280 31340 18315
rect 31350 18280 31385 18315
rect 31395 18280 31430 18315
rect 31440 18280 31475 18315
rect 31485 18280 31520 18315
rect 31530 18280 31565 18315
rect 31575 18280 31610 18315
rect 31620 18280 31655 18315
rect 31665 18280 31700 18315
rect 31710 18280 31745 18315
rect 31755 18280 31790 18315
rect 31800 18280 31835 18315
rect 31845 18280 31880 18315
rect 31890 18280 31925 18315
rect 31935 18280 31970 18315
rect 31980 18280 32015 18315
rect 32025 18280 32060 18315
rect 32070 18280 32105 18315
rect 32115 18280 32150 18315
rect 32160 18280 32195 18315
rect 32205 18280 32240 18315
rect 32250 18280 32285 18315
rect 32295 18280 32330 18315
rect 32340 18280 32375 18315
rect 32385 18280 32420 18315
rect 32430 18280 32465 18315
rect 32475 18280 32510 18315
rect 32520 18280 32555 18315
rect 32565 18280 32600 18315
rect 32610 18280 32645 18315
rect 32655 18280 32690 18315
rect 32700 18280 32735 18315
rect 32745 18280 32780 18315
rect 32790 18280 32825 18315
rect 32835 18280 32870 18315
rect 31305 18235 31340 18270
rect 31350 18235 31385 18270
rect 31395 18235 31430 18270
rect 31440 18235 31475 18270
rect 31485 18235 31520 18270
rect 31530 18235 31565 18270
rect 31575 18235 31610 18270
rect 31620 18235 31655 18270
rect 31665 18235 31700 18270
rect 31710 18235 31745 18270
rect 31755 18235 31790 18270
rect 31800 18235 31835 18270
rect 31845 18235 31880 18270
rect 31890 18235 31925 18270
rect 31935 18235 31970 18270
rect 31980 18235 32015 18270
rect 32025 18235 32060 18270
rect 32070 18235 32105 18270
rect 32115 18235 32150 18270
rect 32160 18235 32195 18270
rect 32205 18235 32240 18270
rect 32250 18235 32285 18270
rect 32295 18235 32330 18270
rect 32340 18235 32375 18270
rect 32385 18235 32420 18270
rect 32430 18235 32465 18270
rect 32475 18235 32510 18270
rect 32520 18235 32555 18270
rect 32565 18235 32600 18270
rect 32610 18235 32645 18270
rect 32655 18235 32690 18270
rect 32700 18235 32735 18270
rect 32745 18235 32780 18270
rect 32790 18235 32825 18270
rect 32835 18235 32870 18270
rect 31305 18190 31340 18225
rect 31350 18190 31385 18225
rect 31395 18190 31430 18225
rect 31440 18190 31475 18225
rect 31485 18190 31520 18225
rect 31530 18190 31565 18225
rect 31575 18190 31610 18225
rect 31620 18190 31655 18225
rect 31665 18190 31700 18225
rect 31710 18190 31745 18225
rect 31755 18190 31790 18225
rect 31800 18190 31835 18225
rect 31845 18190 31880 18225
rect 31890 18190 31925 18225
rect 31935 18190 31970 18225
rect 31980 18190 32015 18225
rect 32025 18190 32060 18225
rect 32070 18190 32105 18225
rect 32115 18190 32150 18225
rect 32160 18190 32195 18225
rect 32205 18190 32240 18225
rect 32250 18190 32285 18225
rect 32295 18190 32330 18225
rect 32340 18190 32375 18225
rect 32385 18190 32420 18225
rect 32430 18190 32465 18225
rect 32475 18190 32510 18225
rect 32520 18190 32555 18225
rect 32565 18190 32600 18225
rect 32610 18190 32645 18225
rect 32655 18190 32690 18225
rect 32700 18190 32735 18225
rect 32745 18190 32780 18225
rect 32790 18190 32825 18225
rect 32835 18190 32870 18225
rect 31305 18145 31340 18180
rect 31350 18145 31385 18180
rect 31395 18145 31430 18180
rect 31440 18145 31475 18180
rect 31485 18145 31520 18180
rect 31530 18145 31565 18180
rect 31575 18145 31610 18180
rect 31620 18145 31655 18180
rect 31665 18145 31700 18180
rect 31710 18145 31745 18180
rect 31755 18145 31790 18180
rect 31800 18145 31835 18180
rect 31845 18145 31880 18180
rect 31890 18145 31925 18180
rect 31935 18145 31970 18180
rect 31980 18145 32015 18180
rect 32025 18145 32060 18180
rect 32070 18145 32105 18180
rect 32115 18145 32150 18180
rect 32160 18145 32195 18180
rect 32205 18145 32240 18180
rect 32250 18145 32285 18180
rect 32295 18145 32330 18180
rect 32340 18145 32375 18180
rect 32385 18145 32420 18180
rect 32430 18145 32465 18180
rect 32475 18145 32510 18180
rect 32520 18145 32555 18180
rect 32565 18145 32600 18180
rect 32610 18145 32645 18180
rect 32655 18145 32690 18180
rect 32700 18145 32735 18180
rect 32745 18145 32780 18180
rect 32790 18145 32825 18180
rect 32835 18145 32870 18180
rect 31305 18100 31340 18135
rect 31350 18100 31385 18135
rect 31395 18100 31430 18135
rect 31440 18100 31475 18135
rect 31485 18100 31520 18135
rect 31530 18100 31565 18135
rect 31575 18100 31610 18135
rect 31620 18100 31655 18135
rect 31665 18100 31700 18135
rect 31710 18100 31745 18135
rect 31755 18100 31790 18135
rect 31800 18100 31835 18135
rect 31845 18100 31880 18135
rect 31890 18100 31925 18135
rect 31935 18100 31970 18135
rect 31980 18100 32015 18135
rect 32025 18100 32060 18135
rect 32070 18100 32105 18135
rect 32115 18100 32150 18135
rect 32160 18100 32195 18135
rect 32205 18100 32240 18135
rect 32250 18100 32285 18135
rect 32295 18100 32330 18135
rect 32340 18100 32375 18135
rect 32385 18100 32420 18135
rect 32430 18100 32465 18135
rect 32475 18100 32510 18135
rect 32520 18100 32555 18135
rect 32565 18100 32600 18135
rect 32610 18100 32645 18135
rect 32655 18100 32690 18135
rect 32700 18100 32735 18135
rect 32745 18100 32780 18135
rect 32790 18100 32825 18135
rect 32835 18100 32870 18135
rect 31305 18055 31340 18090
rect 31350 18055 31385 18090
rect 31395 18055 31430 18090
rect 31440 18055 31475 18090
rect 31485 18055 31520 18090
rect 31530 18055 31565 18090
rect 31575 18055 31610 18090
rect 31620 18055 31655 18090
rect 31665 18055 31700 18090
rect 31710 18055 31745 18090
rect 31755 18055 31790 18090
rect 31800 18055 31835 18090
rect 31845 18055 31880 18090
rect 31890 18055 31925 18090
rect 31935 18055 31970 18090
rect 31980 18055 32015 18090
rect 32025 18055 32060 18090
rect 32070 18055 32105 18090
rect 32115 18055 32150 18090
rect 32160 18055 32195 18090
rect 32205 18055 32240 18090
rect 32250 18055 32285 18090
rect 32295 18055 32330 18090
rect 32340 18055 32375 18090
rect 32385 18055 32420 18090
rect 32430 18055 32465 18090
rect 32475 18055 32510 18090
rect 32520 18055 32555 18090
rect 32565 18055 32600 18090
rect 32610 18055 32645 18090
rect 32655 18055 32690 18090
rect 32700 18055 32735 18090
rect 32745 18055 32780 18090
rect 32790 18055 32825 18090
rect 32835 18055 32870 18090
rect 31305 18010 31340 18045
rect 31350 18010 31385 18045
rect 31395 18010 31430 18045
rect 31440 18010 31475 18045
rect 31485 18010 31520 18045
rect 31530 18010 31565 18045
rect 31575 18010 31610 18045
rect 31620 18010 31655 18045
rect 31665 18010 31700 18045
rect 31710 18010 31745 18045
rect 31755 18010 31790 18045
rect 31800 18010 31835 18045
rect 31845 18010 31880 18045
rect 31890 18010 31925 18045
rect 31935 18010 31970 18045
rect 31980 18010 32015 18045
rect 32025 18010 32060 18045
rect 32070 18010 32105 18045
rect 32115 18010 32150 18045
rect 32160 18010 32195 18045
rect 32205 18010 32240 18045
rect 32250 18010 32285 18045
rect 32295 18010 32330 18045
rect 32340 18010 32375 18045
rect 32385 18010 32420 18045
rect 32430 18010 32465 18045
rect 32475 18010 32510 18045
rect 32520 18010 32555 18045
rect 32565 18010 32600 18045
rect 32610 18010 32645 18045
rect 32655 18010 32690 18045
rect 32700 18010 32735 18045
rect 32745 18010 32780 18045
rect 32790 18010 32825 18045
rect 32835 18010 32870 18045
rect 31305 17965 31340 18000
rect 31350 17965 31385 18000
rect 31395 17965 31430 18000
rect 31440 17965 31475 18000
rect 31485 17965 31520 18000
rect 31530 17965 31565 18000
rect 31575 17965 31610 18000
rect 31620 17965 31655 18000
rect 31665 17965 31700 18000
rect 31710 17965 31745 18000
rect 31755 17965 31790 18000
rect 31800 17965 31835 18000
rect 31845 17965 31880 18000
rect 31890 17965 31925 18000
rect 31935 17965 31970 18000
rect 31980 17965 32015 18000
rect 32025 17965 32060 18000
rect 32070 17965 32105 18000
rect 32115 17965 32150 18000
rect 32160 17965 32195 18000
rect 32205 17965 32240 18000
rect 32250 17965 32285 18000
rect 32295 17965 32330 18000
rect 32340 17965 32375 18000
rect 32385 17965 32420 18000
rect 32430 17965 32465 18000
rect 32475 17965 32510 18000
rect 32520 17965 32555 18000
rect 32565 17965 32600 18000
rect 32610 17965 32645 18000
rect 32655 17965 32690 18000
rect 32700 17965 32735 18000
rect 32745 17965 32780 18000
rect 32790 17965 32825 18000
rect 32835 17965 32870 18000
rect 31305 17920 31340 17955
rect 31350 17920 31385 17955
rect 31395 17920 31430 17955
rect 31440 17920 31475 17955
rect 31485 17920 31520 17955
rect 31530 17920 31565 17955
rect 31575 17920 31610 17955
rect 31620 17920 31655 17955
rect 31665 17920 31700 17955
rect 31710 17920 31745 17955
rect 31755 17920 31790 17955
rect 31800 17920 31835 17955
rect 31845 17920 31880 17955
rect 31890 17920 31925 17955
rect 31935 17920 31970 17955
rect 31980 17920 32015 17955
rect 32025 17920 32060 17955
rect 32070 17920 32105 17955
rect 32115 17920 32150 17955
rect 32160 17920 32195 17955
rect 32205 17920 32240 17955
rect 32250 17920 32285 17955
rect 32295 17920 32330 17955
rect 32340 17920 32375 17955
rect 32385 17920 32420 17955
rect 32430 17920 32465 17955
rect 32475 17920 32510 17955
rect 32520 17920 32555 17955
rect 32565 17920 32600 17955
rect 32610 17920 32645 17955
rect 32655 17920 32690 17955
rect 32700 17920 32735 17955
rect 32745 17920 32780 17955
rect 32790 17920 32825 17955
rect 32835 17920 32870 17955
rect 31305 17875 31340 17910
rect 31350 17875 31385 17910
rect 31395 17875 31430 17910
rect 31440 17875 31475 17910
rect 31485 17875 31520 17910
rect 31530 17875 31565 17910
rect 31575 17875 31610 17910
rect 31620 17875 31655 17910
rect 31665 17875 31700 17910
rect 31710 17875 31745 17910
rect 31755 17875 31790 17910
rect 31800 17875 31835 17910
rect 31845 17875 31880 17910
rect 31890 17875 31925 17910
rect 31935 17875 31970 17910
rect 31980 17875 32015 17910
rect 32025 17875 32060 17910
rect 32070 17875 32105 17910
rect 32115 17875 32150 17910
rect 32160 17875 32195 17910
rect 32205 17875 32240 17910
rect 32250 17875 32285 17910
rect 32295 17875 32330 17910
rect 32340 17875 32375 17910
rect 32385 17875 32420 17910
rect 32430 17875 32465 17910
rect 32475 17875 32510 17910
rect 32520 17875 32555 17910
rect 32565 17875 32600 17910
rect 32610 17875 32645 17910
rect 32655 17875 32690 17910
rect 32700 17875 32735 17910
rect 32745 17875 32780 17910
rect 32790 17875 32825 17910
rect 32835 17875 32870 17910
rect 31305 17830 31340 17865
rect 31350 17830 31385 17865
rect 31395 17830 31430 17865
rect 31440 17830 31475 17865
rect 31485 17830 31520 17865
rect 31530 17830 31565 17865
rect 31575 17830 31610 17865
rect 31620 17830 31655 17865
rect 31665 17830 31700 17865
rect 31710 17830 31745 17865
rect 31755 17830 31790 17865
rect 31800 17830 31835 17865
rect 31845 17830 31880 17865
rect 31890 17830 31925 17865
rect 31935 17830 31970 17865
rect 31980 17830 32015 17865
rect 32025 17830 32060 17865
rect 32070 17830 32105 17865
rect 32115 17830 32150 17865
rect 32160 17830 32195 17865
rect 32205 17830 32240 17865
rect 32250 17830 32285 17865
rect 32295 17830 32330 17865
rect 32340 17830 32375 17865
rect 32385 17830 32420 17865
rect 32430 17830 32465 17865
rect 32475 17830 32510 17865
rect 32520 17830 32555 17865
rect 32565 17830 32600 17865
rect 32610 17830 32645 17865
rect 32655 17830 32690 17865
rect 32700 17830 32735 17865
rect 32745 17830 32780 17865
rect 32790 17830 32825 17865
rect 32835 17830 32870 17865
rect 31305 17785 31340 17820
rect 31350 17785 31385 17820
rect 31395 17785 31430 17820
rect 31440 17785 31475 17820
rect 31485 17785 31520 17820
rect 31530 17785 31565 17820
rect 31575 17785 31610 17820
rect 31620 17785 31655 17820
rect 31665 17785 31700 17820
rect 31710 17785 31745 17820
rect 31755 17785 31790 17820
rect 31800 17785 31835 17820
rect 31845 17785 31880 17820
rect 31890 17785 31925 17820
rect 31935 17785 31970 17820
rect 31980 17785 32015 17820
rect 32025 17785 32060 17820
rect 32070 17785 32105 17820
rect 32115 17785 32150 17820
rect 32160 17785 32195 17820
rect 32205 17785 32240 17820
rect 32250 17785 32285 17820
rect 32295 17785 32330 17820
rect 32340 17785 32375 17820
rect 32385 17785 32420 17820
rect 32430 17785 32465 17820
rect 32475 17785 32510 17820
rect 32520 17785 32555 17820
rect 32565 17785 32600 17820
rect 32610 17785 32645 17820
rect 32655 17785 32690 17820
rect 32700 17785 32735 17820
rect 32745 17785 32780 17820
rect 32790 17785 32825 17820
rect 32835 17785 32870 17820
rect 31305 17740 31340 17775
rect 31350 17740 31385 17775
rect 31395 17740 31430 17775
rect 31440 17740 31475 17775
rect 31485 17740 31520 17775
rect 31530 17740 31565 17775
rect 31575 17740 31610 17775
rect 31620 17740 31655 17775
rect 31665 17740 31700 17775
rect 31710 17740 31745 17775
rect 31755 17740 31790 17775
rect 31800 17740 31835 17775
rect 31845 17740 31880 17775
rect 31890 17740 31925 17775
rect 31935 17740 31970 17775
rect 31980 17740 32015 17775
rect 32025 17740 32060 17775
rect 32070 17740 32105 17775
rect 32115 17740 32150 17775
rect 32160 17740 32195 17775
rect 32205 17740 32240 17775
rect 32250 17740 32285 17775
rect 32295 17740 32330 17775
rect 32340 17740 32375 17775
rect 32385 17740 32420 17775
rect 32430 17740 32465 17775
rect 32475 17740 32510 17775
rect 32520 17740 32555 17775
rect 32565 17740 32600 17775
rect 32610 17740 32645 17775
rect 32655 17740 32690 17775
rect 32700 17740 32735 17775
rect 32745 17740 32780 17775
rect 32790 17740 32825 17775
rect 32835 17740 32870 17775
rect -38755 9595 -38720 9630
rect -38710 9595 -38675 9630
rect -38665 9595 -38630 9630
rect -38620 9595 -38585 9630
rect -38575 9595 -38540 9630
rect -38530 9595 -38495 9630
rect -38485 9595 -38450 9630
rect -38440 9595 -38405 9630
rect -38395 9595 -38360 9630
rect -38350 9595 -38315 9630
rect -38305 9595 -38270 9630
rect -38260 9595 -38225 9630
rect -38215 9595 -38180 9630
rect -38170 9595 -38135 9630
rect -38125 9595 -38090 9630
rect -38080 9595 -38045 9630
rect -38035 9595 -38000 9630
rect -37990 9595 -37955 9630
rect -37945 9595 -37910 9630
rect -37900 9595 -37865 9630
rect -37855 9595 -37820 9630
rect -37810 9595 -37775 9630
rect -37765 9595 -37730 9630
rect -37720 9595 -37685 9630
rect -37675 9595 -37640 9630
rect -37630 9595 -37595 9630
rect -37585 9595 -37550 9630
rect -37540 9595 -37505 9630
rect -37495 9595 -37460 9630
rect -37450 9595 -37415 9630
rect -37405 9595 -37370 9630
rect -37360 9595 -37325 9630
rect -37315 9595 -37280 9630
rect -37270 9595 -37235 9630
rect -37225 9595 -37190 9630
rect -38755 9550 -38720 9585
rect -38710 9550 -38675 9585
rect -38665 9550 -38630 9585
rect -38620 9550 -38585 9585
rect -38575 9550 -38540 9585
rect -38530 9550 -38495 9585
rect -38485 9550 -38450 9585
rect -38440 9550 -38405 9585
rect -38395 9550 -38360 9585
rect -38350 9550 -38315 9585
rect -38305 9550 -38270 9585
rect -38260 9550 -38225 9585
rect -38215 9550 -38180 9585
rect -38170 9550 -38135 9585
rect -38125 9550 -38090 9585
rect -38080 9550 -38045 9585
rect -38035 9550 -38000 9585
rect -37990 9550 -37955 9585
rect -37945 9550 -37910 9585
rect -37900 9550 -37865 9585
rect -37855 9550 -37820 9585
rect -37810 9550 -37775 9585
rect -37765 9550 -37730 9585
rect -37720 9550 -37685 9585
rect -37675 9550 -37640 9585
rect -37630 9550 -37595 9585
rect -37585 9550 -37550 9585
rect -37540 9550 -37505 9585
rect -37495 9550 -37460 9585
rect -37450 9550 -37415 9585
rect -37405 9550 -37370 9585
rect -37360 9550 -37325 9585
rect -37315 9550 -37280 9585
rect -37270 9550 -37235 9585
rect -37225 9550 -37190 9585
rect -38755 9505 -38720 9540
rect -38710 9505 -38675 9540
rect -38665 9505 -38630 9540
rect -38620 9505 -38585 9540
rect -38575 9505 -38540 9540
rect -38530 9505 -38495 9540
rect -38485 9505 -38450 9540
rect -38440 9505 -38405 9540
rect -38395 9505 -38360 9540
rect -38350 9505 -38315 9540
rect -38305 9505 -38270 9540
rect -38260 9505 -38225 9540
rect -38215 9505 -38180 9540
rect -38170 9505 -38135 9540
rect -38125 9505 -38090 9540
rect -38080 9505 -38045 9540
rect -38035 9505 -38000 9540
rect -37990 9505 -37955 9540
rect -37945 9505 -37910 9540
rect -37900 9505 -37865 9540
rect -37855 9505 -37820 9540
rect -37810 9505 -37775 9540
rect -37765 9505 -37730 9540
rect -37720 9505 -37685 9540
rect -37675 9505 -37640 9540
rect -37630 9505 -37595 9540
rect -37585 9505 -37550 9540
rect -37540 9505 -37505 9540
rect -37495 9505 -37460 9540
rect -37450 9505 -37415 9540
rect -37405 9505 -37370 9540
rect -37360 9505 -37325 9540
rect -37315 9505 -37280 9540
rect -37270 9505 -37235 9540
rect -37225 9505 -37190 9540
rect -38755 9460 -38720 9495
rect -38710 9460 -38675 9495
rect -38665 9460 -38630 9495
rect -38620 9460 -38585 9495
rect -38575 9460 -38540 9495
rect -38530 9460 -38495 9495
rect -38485 9460 -38450 9495
rect -38440 9460 -38405 9495
rect -38395 9460 -38360 9495
rect -38350 9460 -38315 9495
rect -38305 9460 -38270 9495
rect -38260 9460 -38225 9495
rect -38215 9460 -38180 9495
rect -38170 9460 -38135 9495
rect -38125 9460 -38090 9495
rect -38080 9460 -38045 9495
rect -38035 9460 -38000 9495
rect -37990 9460 -37955 9495
rect -37945 9460 -37910 9495
rect -37900 9460 -37865 9495
rect -37855 9460 -37820 9495
rect -37810 9460 -37775 9495
rect -37765 9460 -37730 9495
rect -37720 9460 -37685 9495
rect -37675 9460 -37640 9495
rect -37630 9460 -37595 9495
rect -37585 9460 -37550 9495
rect -37540 9460 -37505 9495
rect -37495 9460 -37460 9495
rect -37450 9460 -37415 9495
rect -37405 9460 -37370 9495
rect -37360 9460 -37325 9495
rect -37315 9460 -37280 9495
rect -37270 9460 -37235 9495
rect -37225 9460 -37190 9495
rect -38755 9415 -38720 9450
rect -38710 9415 -38675 9450
rect -38665 9415 -38630 9450
rect -38620 9415 -38585 9450
rect -38575 9415 -38540 9450
rect -38530 9415 -38495 9450
rect -38485 9415 -38450 9450
rect -38440 9415 -38405 9450
rect -38395 9415 -38360 9450
rect -38350 9415 -38315 9450
rect -38305 9415 -38270 9450
rect -38260 9415 -38225 9450
rect -38215 9415 -38180 9450
rect -38170 9415 -38135 9450
rect -38125 9415 -38090 9450
rect -38080 9415 -38045 9450
rect -38035 9415 -38000 9450
rect -37990 9415 -37955 9450
rect -37945 9415 -37910 9450
rect -37900 9415 -37865 9450
rect -37855 9415 -37820 9450
rect -37810 9415 -37775 9450
rect -37765 9415 -37730 9450
rect -37720 9415 -37685 9450
rect -37675 9415 -37640 9450
rect -37630 9415 -37595 9450
rect -37585 9415 -37550 9450
rect -37540 9415 -37505 9450
rect -37495 9415 -37460 9450
rect -37450 9415 -37415 9450
rect -37405 9415 -37370 9450
rect -37360 9415 -37325 9450
rect -37315 9415 -37280 9450
rect -37270 9415 -37235 9450
rect -37225 9415 -37190 9450
rect -38755 9370 -38720 9405
rect -38710 9370 -38675 9405
rect -38665 9370 -38630 9405
rect -38620 9370 -38585 9405
rect -38575 9370 -38540 9405
rect -38530 9370 -38495 9405
rect -38485 9370 -38450 9405
rect -38440 9370 -38405 9405
rect -38395 9370 -38360 9405
rect -38350 9370 -38315 9405
rect -38305 9370 -38270 9405
rect -38260 9370 -38225 9405
rect -38215 9370 -38180 9405
rect -38170 9370 -38135 9405
rect -38125 9370 -38090 9405
rect -38080 9370 -38045 9405
rect -38035 9370 -38000 9405
rect -37990 9370 -37955 9405
rect -37945 9370 -37910 9405
rect -37900 9370 -37865 9405
rect -37855 9370 -37820 9405
rect -37810 9370 -37775 9405
rect -37765 9370 -37730 9405
rect -37720 9370 -37685 9405
rect -37675 9370 -37640 9405
rect -37630 9370 -37595 9405
rect -37585 9370 -37550 9405
rect -37540 9370 -37505 9405
rect -37495 9370 -37460 9405
rect -37450 9370 -37415 9405
rect -37405 9370 -37370 9405
rect -37360 9370 -37325 9405
rect -37315 9370 -37280 9405
rect -37270 9370 -37235 9405
rect -37225 9370 -37190 9405
rect -38755 9325 -38720 9360
rect -38710 9325 -38675 9360
rect -38665 9325 -38630 9360
rect -38620 9325 -38585 9360
rect -38575 9325 -38540 9360
rect -38530 9325 -38495 9360
rect -38485 9325 -38450 9360
rect -38440 9325 -38405 9360
rect -38395 9325 -38360 9360
rect -38350 9325 -38315 9360
rect -38305 9325 -38270 9360
rect -38260 9325 -38225 9360
rect -38215 9325 -38180 9360
rect -38170 9325 -38135 9360
rect -38125 9325 -38090 9360
rect -38080 9325 -38045 9360
rect -38035 9325 -38000 9360
rect -37990 9325 -37955 9360
rect -37945 9325 -37910 9360
rect -37900 9325 -37865 9360
rect -37855 9325 -37820 9360
rect -37810 9325 -37775 9360
rect -37765 9325 -37730 9360
rect -37720 9325 -37685 9360
rect -37675 9325 -37640 9360
rect -37630 9325 -37595 9360
rect -37585 9325 -37550 9360
rect -37540 9325 -37505 9360
rect -37495 9325 -37460 9360
rect -37450 9325 -37415 9360
rect -37405 9325 -37370 9360
rect -37360 9325 -37325 9360
rect -37315 9325 -37280 9360
rect -37270 9325 -37235 9360
rect -37225 9325 -37190 9360
rect -38755 9280 -38720 9315
rect -38710 9280 -38675 9315
rect -38665 9280 -38630 9315
rect -38620 9280 -38585 9315
rect -38575 9280 -38540 9315
rect -38530 9280 -38495 9315
rect -38485 9280 -38450 9315
rect -38440 9280 -38405 9315
rect -38395 9280 -38360 9315
rect -38350 9280 -38315 9315
rect -38305 9280 -38270 9315
rect -38260 9280 -38225 9315
rect -38215 9280 -38180 9315
rect -38170 9280 -38135 9315
rect -38125 9280 -38090 9315
rect -38080 9280 -38045 9315
rect -38035 9280 -38000 9315
rect -37990 9280 -37955 9315
rect -37945 9280 -37910 9315
rect -37900 9280 -37865 9315
rect -37855 9280 -37820 9315
rect -37810 9280 -37775 9315
rect -37765 9280 -37730 9315
rect -37720 9280 -37685 9315
rect -37675 9280 -37640 9315
rect -37630 9280 -37595 9315
rect -37585 9280 -37550 9315
rect -37540 9280 -37505 9315
rect -37495 9280 -37460 9315
rect -37450 9280 -37415 9315
rect -37405 9280 -37370 9315
rect -37360 9280 -37325 9315
rect -37315 9280 -37280 9315
rect -37270 9280 -37235 9315
rect -37225 9280 -37190 9315
rect -38755 9235 -38720 9270
rect -38710 9235 -38675 9270
rect -38665 9235 -38630 9270
rect -38620 9235 -38585 9270
rect -38575 9235 -38540 9270
rect -38530 9235 -38495 9270
rect -38485 9235 -38450 9270
rect -38440 9235 -38405 9270
rect -38395 9235 -38360 9270
rect -38350 9235 -38315 9270
rect -38305 9235 -38270 9270
rect -38260 9235 -38225 9270
rect -38215 9235 -38180 9270
rect -38170 9235 -38135 9270
rect -38125 9235 -38090 9270
rect -38080 9235 -38045 9270
rect -38035 9235 -38000 9270
rect -37990 9235 -37955 9270
rect -37945 9235 -37910 9270
rect -37900 9235 -37865 9270
rect -37855 9235 -37820 9270
rect -37810 9235 -37775 9270
rect -37765 9235 -37730 9270
rect -37720 9235 -37685 9270
rect -37675 9235 -37640 9270
rect -37630 9235 -37595 9270
rect -37585 9235 -37550 9270
rect -37540 9235 -37505 9270
rect -37495 9235 -37460 9270
rect -37450 9235 -37415 9270
rect -37405 9235 -37370 9270
rect -37360 9235 -37325 9270
rect -37315 9235 -37280 9270
rect -37270 9235 -37235 9270
rect -37225 9235 -37190 9270
rect -38755 9190 -38720 9225
rect -38710 9190 -38675 9225
rect -38665 9190 -38630 9225
rect -38620 9190 -38585 9225
rect -38575 9190 -38540 9225
rect -38530 9190 -38495 9225
rect -38485 9190 -38450 9225
rect -38440 9190 -38405 9225
rect -38395 9190 -38360 9225
rect -38350 9190 -38315 9225
rect -38305 9190 -38270 9225
rect -38260 9190 -38225 9225
rect -38215 9190 -38180 9225
rect -38170 9190 -38135 9225
rect -38125 9190 -38090 9225
rect -38080 9190 -38045 9225
rect -38035 9190 -38000 9225
rect -37990 9190 -37955 9225
rect -37945 9190 -37910 9225
rect -37900 9190 -37865 9225
rect -37855 9190 -37820 9225
rect -37810 9190 -37775 9225
rect -37765 9190 -37730 9225
rect -37720 9190 -37685 9225
rect -37675 9190 -37640 9225
rect -37630 9190 -37595 9225
rect -37585 9190 -37550 9225
rect -37540 9190 -37505 9225
rect -37495 9190 -37460 9225
rect -37450 9190 -37415 9225
rect -37405 9190 -37370 9225
rect -37360 9190 -37325 9225
rect -37315 9190 -37280 9225
rect -37270 9190 -37235 9225
rect -37225 9190 -37190 9225
rect -38755 9145 -38720 9180
rect -38710 9145 -38675 9180
rect -38665 9145 -38630 9180
rect -38620 9145 -38585 9180
rect -38575 9145 -38540 9180
rect -38530 9145 -38495 9180
rect -38485 9145 -38450 9180
rect -38440 9145 -38405 9180
rect -38395 9145 -38360 9180
rect -38350 9145 -38315 9180
rect -38305 9145 -38270 9180
rect -38260 9145 -38225 9180
rect -38215 9145 -38180 9180
rect -38170 9145 -38135 9180
rect -38125 9145 -38090 9180
rect -38080 9145 -38045 9180
rect -38035 9145 -38000 9180
rect -37990 9145 -37955 9180
rect -37945 9145 -37910 9180
rect -37900 9145 -37865 9180
rect -37855 9145 -37820 9180
rect -37810 9145 -37775 9180
rect -37765 9145 -37730 9180
rect -37720 9145 -37685 9180
rect -37675 9145 -37640 9180
rect -37630 9145 -37595 9180
rect -37585 9145 -37550 9180
rect -37540 9145 -37505 9180
rect -37495 9145 -37460 9180
rect -37450 9145 -37415 9180
rect -37405 9145 -37370 9180
rect -37360 9145 -37325 9180
rect -37315 9145 -37280 9180
rect -37270 9145 -37235 9180
rect -37225 9145 -37190 9180
rect -38755 9100 -38720 9135
rect -38710 9100 -38675 9135
rect -38665 9100 -38630 9135
rect -38620 9100 -38585 9135
rect -38575 9100 -38540 9135
rect -38530 9100 -38495 9135
rect -38485 9100 -38450 9135
rect -38440 9100 -38405 9135
rect -38395 9100 -38360 9135
rect -38350 9100 -38315 9135
rect -38305 9100 -38270 9135
rect -38260 9100 -38225 9135
rect -38215 9100 -38180 9135
rect -38170 9100 -38135 9135
rect -38125 9100 -38090 9135
rect -38080 9100 -38045 9135
rect -38035 9100 -38000 9135
rect -37990 9100 -37955 9135
rect -37945 9100 -37910 9135
rect -37900 9100 -37865 9135
rect -37855 9100 -37820 9135
rect -37810 9100 -37775 9135
rect -37765 9100 -37730 9135
rect -37720 9100 -37685 9135
rect -37675 9100 -37640 9135
rect -37630 9100 -37595 9135
rect -37585 9100 -37550 9135
rect -37540 9100 -37505 9135
rect -37495 9100 -37460 9135
rect -37450 9100 -37415 9135
rect -37405 9100 -37370 9135
rect -37360 9100 -37325 9135
rect -37315 9100 -37280 9135
rect -37270 9100 -37235 9135
rect -37225 9100 -37190 9135
rect -38755 9055 -38720 9090
rect -38710 9055 -38675 9090
rect -38665 9055 -38630 9090
rect -38620 9055 -38585 9090
rect -38575 9055 -38540 9090
rect -38530 9055 -38495 9090
rect -38485 9055 -38450 9090
rect -38440 9055 -38405 9090
rect -38395 9055 -38360 9090
rect -38350 9055 -38315 9090
rect -38305 9055 -38270 9090
rect -38260 9055 -38225 9090
rect -38215 9055 -38180 9090
rect -38170 9055 -38135 9090
rect -38125 9055 -38090 9090
rect -38080 9055 -38045 9090
rect -38035 9055 -38000 9090
rect -37990 9055 -37955 9090
rect -37945 9055 -37910 9090
rect -37900 9055 -37865 9090
rect -37855 9055 -37820 9090
rect -37810 9055 -37775 9090
rect -37765 9055 -37730 9090
rect -37720 9055 -37685 9090
rect -37675 9055 -37640 9090
rect -37630 9055 -37595 9090
rect -37585 9055 -37550 9090
rect -37540 9055 -37505 9090
rect -37495 9055 -37460 9090
rect -37450 9055 -37415 9090
rect -37405 9055 -37370 9090
rect -37360 9055 -37325 9090
rect -37315 9055 -37280 9090
rect -37270 9055 -37235 9090
rect -37225 9055 -37190 9090
rect -38755 9010 -38720 9045
rect -38710 9010 -38675 9045
rect -38665 9010 -38630 9045
rect -38620 9010 -38585 9045
rect -38575 9010 -38540 9045
rect -38530 9010 -38495 9045
rect -38485 9010 -38450 9045
rect -38440 9010 -38405 9045
rect -38395 9010 -38360 9045
rect -38350 9010 -38315 9045
rect -38305 9010 -38270 9045
rect -38260 9010 -38225 9045
rect -38215 9010 -38180 9045
rect -38170 9010 -38135 9045
rect -38125 9010 -38090 9045
rect -38080 9010 -38045 9045
rect -38035 9010 -38000 9045
rect -37990 9010 -37955 9045
rect -37945 9010 -37910 9045
rect -37900 9010 -37865 9045
rect -37855 9010 -37820 9045
rect -37810 9010 -37775 9045
rect -37765 9010 -37730 9045
rect -37720 9010 -37685 9045
rect -37675 9010 -37640 9045
rect -37630 9010 -37595 9045
rect -37585 9010 -37550 9045
rect -37540 9010 -37505 9045
rect -37495 9010 -37460 9045
rect -37450 9010 -37415 9045
rect -37405 9010 -37370 9045
rect -37360 9010 -37325 9045
rect -37315 9010 -37280 9045
rect -37270 9010 -37235 9045
rect -37225 9010 -37190 9045
rect -38755 8965 -38720 9000
rect -38710 8965 -38675 9000
rect -38665 8965 -38630 9000
rect -38620 8965 -38585 9000
rect -38575 8965 -38540 9000
rect -38530 8965 -38495 9000
rect -38485 8965 -38450 9000
rect -38440 8965 -38405 9000
rect -38395 8965 -38360 9000
rect -38350 8965 -38315 9000
rect -38305 8965 -38270 9000
rect -38260 8965 -38225 9000
rect -38215 8965 -38180 9000
rect -38170 8965 -38135 9000
rect -38125 8965 -38090 9000
rect -38080 8965 -38045 9000
rect -38035 8965 -38000 9000
rect -37990 8965 -37955 9000
rect -37945 8965 -37910 9000
rect -37900 8965 -37865 9000
rect -37855 8965 -37820 9000
rect -37810 8965 -37775 9000
rect -37765 8965 -37730 9000
rect -37720 8965 -37685 9000
rect -37675 8965 -37640 9000
rect -37630 8965 -37595 9000
rect -37585 8965 -37550 9000
rect -37540 8965 -37505 9000
rect -37495 8965 -37460 9000
rect -37450 8965 -37415 9000
rect -37405 8965 -37370 9000
rect -37360 8965 -37325 9000
rect -37315 8965 -37280 9000
rect -37270 8965 -37235 9000
rect -37225 8965 -37190 9000
rect -38755 8920 -38720 8955
rect -38710 8920 -38675 8955
rect -38665 8920 -38630 8955
rect -38620 8920 -38585 8955
rect -38575 8920 -38540 8955
rect -38530 8920 -38495 8955
rect -38485 8920 -38450 8955
rect -38440 8920 -38405 8955
rect -38395 8920 -38360 8955
rect -38350 8920 -38315 8955
rect -38305 8920 -38270 8955
rect -38260 8920 -38225 8955
rect -38215 8920 -38180 8955
rect -38170 8920 -38135 8955
rect -38125 8920 -38090 8955
rect -38080 8920 -38045 8955
rect -38035 8920 -38000 8955
rect -37990 8920 -37955 8955
rect -37945 8920 -37910 8955
rect -37900 8920 -37865 8955
rect -37855 8920 -37820 8955
rect -37810 8920 -37775 8955
rect -37765 8920 -37730 8955
rect -37720 8920 -37685 8955
rect -37675 8920 -37640 8955
rect -37630 8920 -37595 8955
rect -37585 8920 -37550 8955
rect -37540 8920 -37505 8955
rect -37495 8920 -37460 8955
rect -37450 8920 -37415 8955
rect -37405 8920 -37370 8955
rect -37360 8920 -37325 8955
rect -37315 8920 -37280 8955
rect -37270 8920 -37235 8955
rect -37225 8920 -37190 8955
rect -38755 8875 -38720 8910
rect -38710 8875 -38675 8910
rect -38665 8875 -38630 8910
rect -38620 8875 -38585 8910
rect -38575 8875 -38540 8910
rect -38530 8875 -38495 8910
rect -38485 8875 -38450 8910
rect -38440 8875 -38405 8910
rect -38395 8875 -38360 8910
rect -38350 8875 -38315 8910
rect -38305 8875 -38270 8910
rect -38260 8875 -38225 8910
rect -38215 8875 -38180 8910
rect -38170 8875 -38135 8910
rect -38125 8875 -38090 8910
rect -38080 8875 -38045 8910
rect -38035 8875 -38000 8910
rect -37990 8875 -37955 8910
rect -37945 8875 -37910 8910
rect -37900 8875 -37865 8910
rect -37855 8875 -37820 8910
rect -37810 8875 -37775 8910
rect -37765 8875 -37730 8910
rect -37720 8875 -37685 8910
rect -37675 8875 -37640 8910
rect -37630 8875 -37595 8910
rect -37585 8875 -37550 8910
rect -37540 8875 -37505 8910
rect -37495 8875 -37460 8910
rect -37450 8875 -37415 8910
rect -37405 8875 -37370 8910
rect -37360 8875 -37325 8910
rect -37315 8875 -37280 8910
rect -37270 8875 -37235 8910
rect -37225 8875 -37190 8910
rect -38755 8830 -38720 8865
rect -38710 8830 -38675 8865
rect -38665 8830 -38630 8865
rect -38620 8830 -38585 8865
rect -38575 8830 -38540 8865
rect -38530 8830 -38495 8865
rect -38485 8830 -38450 8865
rect -38440 8830 -38405 8865
rect -38395 8830 -38360 8865
rect -38350 8830 -38315 8865
rect -38305 8830 -38270 8865
rect -38260 8830 -38225 8865
rect -38215 8830 -38180 8865
rect -38170 8830 -38135 8865
rect -38125 8830 -38090 8865
rect -38080 8830 -38045 8865
rect -38035 8830 -38000 8865
rect -37990 8830 -37955 8865
rect -37945 8830 -37910 8865
rect -37900 8830 -37865 8865
rect -37855 8830 -37820 8865
rect -37810 8830 -37775 8865
rect -37765 8830 -37730 8865
rect -37720 8830 -37685 8865
rect -37675 8830 -37640 8865
rect -37630 8830 -37595 8865
rect -37585 8830 -37550 8865
rect -37540 8830 -37505 8865
rect -37495 8830 -37460 8865
rect -37450 8830 -37415 8865
rect -37405 8830 -37370 8865
rect -37360 8830 -37325 8865
rect -37315 8830 -37280 8865
rect -37270 8830 -37235 8865
rect -37225 8830 -37190 8865
rect -38755 8785 -38720 8820
rect -38710 8785 -38675 8820
rect -38665 8785 -38630 8820
rect -38620 8785 -38585 8820
rect -38575 8785 -38540 8820
rect -38530 8785 -38495 8820
rect -38485 8785 -38450 8820
rect -38440 8785 -38405 8820
rect -38395 8785 -38360 8820
rect -38350 8785 -38315 8820
rect -38305 8785 -38270 8820
rect -38260 8785 -38225 8820
rect -38215 8785 -38180 8820
rect -38170 8785 -38135 8820
rect -38125 8785 -38090 8820
rect -38080 8785 -38045 8820
rect -38035 8785 -38000 8820
rect -37990 8785 -37955 8820
rect -37945 8785 -37910 8820
rect -37900 8785 -37865 8820
rect -37855 8785 -37820 8820
rect -37810 8785 -37775 8820
rect -37765 8785 -37730 8820
rect -37720 8785 -37685 8820
rect -37675 8785 -37640 8820
rect -37630 8785 -37595 8820
rect -37585 8785 -37550 8820
rect -37540 8785 -37505 8820
rect -37495 8785 -37460 8820
rect -37450 8785 -37415 8820
rect -37405 8785 -37370 8820
rect -37360 8785 -37325 8820
rect -37315 8785 -37280 8820
rect -37270 8785 -37235 8820
rect -37225 8785 -37190 8820
rect -38755 8740 -38720 8775
rect -38710 8740 -38675 8775
rect -38665 8740 -38630 8775
rect -38620 8740 -38585 8775
rect -38575 8740 -38540 8775
rect -38530 8740 -38495 8775
rect -38485 8740 -38450 8775
rect -38440 8740 -38405 8775
rect -38395 8740 -38360 8775
rect -38350 8740 -38315 8775
rect -38305 8740 -38270 8775
rect -38260 8740 -38225 8775
rect -38215 8740 -38180 8775
rect -38170 8740 -38135 8775
rect -38125 8740 -38090 8775
rect -38080 8740 -38045 8775
rect -38035 8740 -38000 8775
rect -37990 8740 -37955 8775
rect -37945 8740 -37910 8775
rect -37900 8740 -37865 8775
rect -37855 8740 -37820 8775
rect -37810 8740 -37775 8775
rect -37765 8740 -37730 8775
rect -37720 8740 -37685 8775
rect -37675 8740 -37640 8775
rect -37630 8740 -37595 8775
rect -37585 8740 -37550 8775
rect -37540 8740 -37505 8775
rect -37495 8740 -37460 8775
rect -37450 8740 -37415 8775
rect -37405 8740 -37370 8775
rect -37360 8740 -37325 8775
rect -37315 8740 -37280 8775
rect -37270 8740 -37235 8775
rect -37225 8740 -37190 8775
rect -38755 8695 -38720 8730
rect -38710 8695 -38675 8730
rect -38665 8695 -38630 8730
rect -38620 8695 -38585 8730
rect -38575 8695 -38540 8730
rect -38530 8695 -38495 8730
rect -38485 8695 -38450 8730
rect -38440 8695 -38405 8730
rect -38395 8695 -38360 8730
rect -38350 8695 -38315 8730
rect -38305 8695 -38270 8730
rect -38260 8695 -38225 8730
rect -38215 8695 -38180 8730
rect -38170 8695 -38135 8730
rect -38125 8695 -38090 8730
rect -38080 8695 -38045 8730
rect -38035 8695 -38000 8730
rect -37990 8695 -37955 8730
rect -37945 8695 -37910 8730
rect -37900 8695 -37865 8730
rect -37855 8695 -37820 8730
rect -37810 8695 -37775 8730
rect -37765 8695 -37730 8730
rect -37720 8695 -37685 8730
rect -37675 8695 -37640 8730
rect -37630 8695 -37595 8730
rect -37585 8695 -37550 8730
rect -37540 8695 -37505 8730
rect -37495 8695 -37460 8730
rect -37450 8695 -37415 8730
rect -37405 8695 -37370 8730
rect -37360 8695 -37325 8730
rect -37315 8695 -37280 8730
rect -37270 8695 -37235 8730
rect -37225 8695 -37190 8730
rect -38755 8650 -38720 8685
rect -38710 8650 -38675 8685
rect -38665 8650 -38630 8685
rect -38620 8650 -38585 8685
rect -38575 8650 -38540 8685
rect -38530 8650 -38495 8685
rect -38485 8650 -38450 8685
rect -38440 8650 -38405 8685
rect -38395 8650 -38360 8685
rect -38350 8650 -38315 8685
rect -38305 8650 -38270 8685
rect -38260 8650 -38225 8685
rect -38215 8650 -38180 8685
rect -38170 8650 -38135 8685
rect -38125 8650 -38090 8685
rect -38080 8650 -38045 8685
rect -38035 8650 -38000 8685
rect -37990 8650 -37955 8685
rect -37945 8650 -37910 8685
rect -37900 8650 -37865 8685
rect -37855 8650 -37820 8685
rect -37810 8650 -37775 8685
rect -37765 8650 -37730 8685
rect -37720 8650 -37685 8685
rect -37675 8650 -37640 8685
rect -37630 8650 -37595 8685
rect -37585 8650 -37550 8685
rect -37540 8650 -37505 8685
rect -37495 8650 -37460 8685
rect -37450 8650 -37415 8685
rect -37405 8650 -37370 8685
rect -37360 8650 -37325 8685
rect -37315 8650 -37280 8685
rect -37270 8650 -37235 8685
rect -37225 8650 -37190 8685
rect -38755 8605 -38720 8640
rect -38710 8605 -38675 8640
rect -38665 8605 -38630 8640
rect -38620 8605 -38585 8640
rect -38575 8605 -38540 8640
rect -38530 8605 -38495 8640
rect -38485 8605 -38450 8640
rect -38440 8605 -38405 8640
rect -38395 8605 -38360 8640
rect -38350 8605 -38315 8640
rect -38305 8605 -38270 8640
rect -38260 8605 -38225 8640
rect -38215 8605 -38180 8640
rect -38170 8605 -38135 8640
rect -38125 8605 -38090 8640
rect -38080 8605 -38045 8640
rect -38035 8605 -38000 8640
rect -37990 8605 -37955 8640
rect -37945 8605 -37910 8640
rect -37900 8605 -37865 8640
rect -37855 8605 -37820 8640
rect -37810 8605 -37775 8640
rect -37765 8605 -37730 8640
rect -37720 8605 -37685 8640
rect -37675 8605 -37640 8640
rect -37630 8605 -37595 8640
rect -37585 8605 -37550 8640
rect -37540 8605 -37505 8640
rect -37495 8605 -37460 8640
rect -37450 8605 -37415 8640
rect -37405 8605 -37370 8640
rect -37360 8605 -37325 8640
rect -37315 8605 -37280 8640
rect -37270 8605 -37235 8640
rect -37225 8605 -37190 8640
rect -38755 8560 -38720 8595
rect -38710 8560 -38675 8595
rect -38665 8560 -38630 8595
rect -38620 8560 -38585 8595
rect -38575 8560 -38540 8595
rect -38530 8560 -38495 8595
rect -38485 8560 -38450 8595
rect -38440 8560 -38405 8595
rect -38395 8560 -38360 8595
rect -38350 8560 -38315 8595
rect -38305 8560 -38270 8595
rect -38260 8560 -38225 8595
rect -38215 8560 -38180 8595
rect -38170 8560 -38135 8595
rect -38125 8560 -38090 8595
rect -38080 8560 -38045 8595
rect -38035 8560 -38000 8595
rect -37990 8560 -37955 8595
rect -37945 8560 -37910 8595
rect -37900 8560 -37865 8595
rect -37855 8560 -37820 8595
rect -37810 8560 -37775 8595
rect -37765 8560 -37730 8595
rect -37720 8560 -37685 8595
rect -37675 8560 -37640 8595
rect -37630 8560 -37595 8595
rect -37585 8560 -37550 8595
rect -37540 8560 -37505 8595
rect -37495 8560 -37460 8595
rect -37450 8560 -37415 8595
rect -37405 8560 -37370 8595
rect -37360 8560 -37325 8595
rect -37315 8560 -37280 8595
rect -37270 8560 -37235 8595
rect -37225 8560 -37190 8595
rect -38755 8515 -38720 8550
rect -38710 8515 -38675 8550
rect -38665 8515 -38630 8550
rect -38620 8515 -38585 8550
rect -38575 8515 -38540 8550
rect -38530 8515 -38495 8550
rect -38485 8515 -38450 8550
rect -38440 8515 -38405 8550
rect -38395 8515 -38360 8550
rect -38350 8515 -38315 8550
rect -38305 8515 -38270 8550
rect -38260 8515 -38225 8550
rect -38215 8515 -38180 8550
rect -38170 8515 -38135 8550
rect -38125 8515 -38090 8550
rect -38080 8515 -38045 8550
rect -38035 8515 -38000 8550
rect -37990 8515 -37955 8550
rect -37945 8515 -37910 8550
rect -37900 8515 -37865 8550
rect -37855 8515 -37820 8550
rect -37810 8515 -37775 8550
rect -37765 8515 -37730 8550
rect -37720 8515 -37685 8550
rect -37675 8515 -37640 8550
rect -37630 8515 -37595 8550
rect -37585 8515 -37550 8550
rect -37540 8515 -37505 8550
rect -37495 8515 -37460 8550
rect -37450 8515 -37415 8550
rect -37405 8515 -37370 8550
rect -37360 8515 -37325 8550
rect -37315 8515 -37280 8550
rect -37270 8515 -37235 8550
rect -37225 8515 -37190 8550
rect -38755 8470 -38720 8505
rect -38710 8470 -38675 8505
rect -38665 8470 -38630 8505
rect -38620 8470 -38585 8505
rect -38575 8470 -38540 8505
rect -38530 8470 -38495 8505
rect -38485 8470 -38450 8505
rect -38440 8470 -38405 8505
rect -38395 8470 -38360 8505
rect -38350 8470 -38315 8505
rect -38305 8470 -38270 8505
rect -38260 8470 -38225 8505
rect -38215 8470 -38180 8505
rect -38170 8470 -38135 8505
rect -38125 8470 -38090 8505
rect -38080 8470 -38045 8505
rect -38035 8470 -38000 8505
rect -37990 8470 -37955 8505
rect -37945 8470 -37910 8505
rect -37900 8470 -37865 8505
rect -37855 8470 -37820 8505
rect -37810 8470 -37775 8505
rect -37765 8470 -37730 8505
rect -37720 8470 -37685 8505
rect -37675 8470 -37640 8505
rect -37630 8470 -37595 8505
rect -37585 8470 -37550 8505
rect -37540 8470 -37505 8505
rect -37495 8470 -37460 8505
rect -37450 8470 -37415 8505
rect -37405 8470 -37370 8505
rect -37360 8470 -37325 8505
rect -37315 8470 -37280 8505
rect -37270 8470 -37235 8505
rect -37225 8470 -37190 8505
rect -38755 8425 -38720 8460
rect -38710 8425 -38675 8460
rect -38665 8425 -38630 8460
rect -38620 8425 -38585 8460
rect -38575 8425 -38540 8460
rect -38530 8425 -38495 8460
rect -38485 8425 -38450 8460
rect -38440 8425 -38405 8460
rect -38395 8425 -38360 8460
rect -38350 8425 -38315 8460
rect -38305 8425 -38270 8460
rect -38260 8425 -38225 8460
rect -38215 8425 -38180 8460
rect -38170 8425 -38135 8460
rect -38125 8425 -38090 8460
rect -38080 8425 -38045 8460
rect -38035 8425 -38000 8460
rect -37990 8425 -37955 8460
rect -37945 8425 -37910 8460
rect -37900 8425 -37865 8460
rect -37855 8425 -37820 8460
rect -37810 8425 -37775 8460
rect -37765 8425 -37730 8460
rect -37720 8425 -37685 8460
rect -37675 8425 -37640 8460
rect -37630 8425 -37595 8460
rect -37585 8425 -37550 8460
rect -37540 8425 -37505 8460
rect -37495 8425 -37460 8460
rect -37450 8425 -37415 8460
rect -37405 8425 -37370 8460
rect -37360 8425 -37325 8460
rect -37315 8425 -37280 8460
rect -37270 8425 -37235 8460
rect -37225 8425 -37190 8460
rect -38755 8380 -38720 8415
rect -38710 8380 -38675 8415
rect -38665 8380 -38630 8415
rect -38620 8380 -38585 8415
rect -38575 8380 -38540 8415
rect -38530 8380 -38495 8415
rect -38485 8380 -38450 8415
rect -38440 8380 -38405 8415
rect -38395 8380 -38360 8415
rect -38350 8380 -38315 8415
rect -38305 8380 -38270 8415
rect -38260 8380 -38225 8415
rect -38215 8380 -38180 8415
rect -38170 8380 -38135 8415
rect -38125 8380 -38090 8415
rect -38080 8380 -38045 8415
rect -38035 8380 -38000 8415
rect -37990 8380 -37955 8415
rect -37945 8380 -37910 8415
rect -37900 8380 -37865 8415
rect -37855 8380 -37820 8415
rect -37810 8380 -37775 8415
rect -37765 8380 -37730 8415
rect -37720 8380 -37685 8415
rect -37675 8380 -37640 8415
rect -37630 8380 -37595 8415
rect -37585 8380 -37550 8415
rect -37540 8380 -37505 8415
rect -37495 8380 -37460 8415
rect -37450 8380 -37415 8415
rect -37405 8380 -37370 8415
rect -37360 8380 -37325 8415
rect -37315 8380 -37280 8415
rect -37270 8380 -37235 8415
rect -37225 8380 -37190 8415
rect -38755 8335 -38720 8370
rect -38710 8335 -38675 8370
rect -38665 8335 -38630 8370
rect -38620 8335 -38585 8370
rect -38575 8335 -38540 8370
rect -38530 8335 -38495 8370
rect -38485 8335 -38450 8370
rect -38440 8335 -38405 8370
rect -38395 8335 -38360 8370
rect -38350 8335 -38315 8370
rect -38305 8335 -38270 8370
rect -38260 8335 -38225 8370
rect -38215 8335 -38180 8370
rect -38170 8335 -38135 8370
rect -38125 8335 -38090 8370
rect -38080 8335 -38045 8370
rect -38035 8335 -38000 8370
rect -37990 8335 -37955 8370
rect -37945 8335 -37910 8370
rect -37900 8335 -37865 8370
rect -37855 8335 -37820 8370
rect -37810 8335 -37775 8370
rect -37765 8335 -37730 8370
rect -37720 8335 -37685 8370
rect -37675 8335 -37640 8370
rect -37630 8335 -37595 8370
rect -37585 8335 -37550 8370
rect -37540 8335 -37505 8370
rect -37495 8335 -37460 8370
rect -37450 8335 -37415 8370
rect -37405 8335 -37370 8370
rect -37360 8335 -37325 8370
rect -37315 8335 -37280 8370
rect -37270 8335 -37235 8370
rect -37225 8335 -37190 8370
rect -38755 8290 -38720 8325
rect -38710 8290 -38675 8325
rect -38665 8290 -38630 8325
rect -38620 8290 -38585 8325
rect -38575 8290 -38540 8325
rect -38530 8290 -38495 8325
rect -38485 8290 -38450 8325
rect -38440 8290 -38405 8325
rect -38395 8290 -38360 8325
rect -38350 8290 -38315 8325
rect -38305 8290 -38270 8325
rect -38260 8290 -38225 8325
rect -38215 8290 -38180 8325
rect -38170 8290 -38135 8325
rect -38125 8290 -38090 8325
rect -38080 8290 -38045 8325
rect -38035 8290 -38000 8325
rect -37990 8290 -37955 8325
rect -37945 8290 -37910 8325
rect -37900 8290 -37865 8325
rect -37855 8290 -37820 8325
rect -37810 8290 -37775 8325
rect -37765 8290 -37730 8325
rect -37720 8290 -37685 8325
rect -37675 8290 -37640 8325
rect -37630 8290 -37595 8325
rect -37585 8290 -37550 8325
rect -37540 8290 -37505 8325
rect -37495 8290 -37460 8325
rect -37450 8290 -37415 8325
rect -37405 8290 -37370 8325
rect -37360 8290 -37325 8325
rect -37315 8290 -37280 8325
rect -37270 8290 -37235 8325
rect -37225 8290 -37190 8325
rect -38755 8245 -38720 8280
rect -38710 8245 -38675 8280
rect -38665 8245 -38630 8280
rect -38620 8245 -38585 8280
rect -38575 8245 -38540 8280
rect -38530 8245 -38495 8280
rect -38485 8245 -38450 8280
rect -38440 8245 -38405 8280
rect -38395 8245 -38360 8280
rect -38350 8245 -38315 8280
rect -38305 8245 -38270 8280
rect -38260 8245 -38225 8280
rect -38215 8245 -38180 8280
rect -38170 8245 -38135 8280
rect -38125 8245 -38090 8280
rect -38080 8245 -38045 8280
rect -38035 8245 -38000 8280
rect -37990 8245 -37955 8280
rect -37945 8245 -37910 8280
rect -37900 8245 -37865 8280
rect -37855 8245 -37820 8280
rect -37810 8245 -37775 8280
rect -37765 8245 -37730 8280
rect -37720 8245 -37685 8280
rect -37675 8245 -37640 8280
rect -37630 8245 -37595 8280
rect -37585 8245 -37550 8280
rect -37540 8245 -37505 8280
rect -37495 8245 -37460 8280
rect -37450 8245 -37415 8280
rect -37405 8245 -37370 8280
rect -37360 8245 -37325 8280
rect -37315 8245 -37280 8280
rect -37270 8245 -37235 8280
rect -37225 8245 -37190 8280
rect -38755 8200 -38720 8235
rect -38710 8200 -38675 8235
rect -38665 8200 -38630 8235
rect -38620 8200 -38585 8235
rect -38575 8200 -38540 8235
rect -38530 8200 -38495 8235
rect -38485 8200 -38450 8235
rect -38440 8200 -38405 8235
rect -38395 8200 -38360 8235
rect -38350 8200 -38315 8235
rect -38305 8200 -38270 8235
rect -38260 8200 -38225 8235
rect -38215 8200 -38180 8235
rect -38170 8200 -38135 8235
rect -38125 8200 -38090 8235
rect -38080 8200 -38045 8235
rect -38035 8200 -38000 8235
rect -37990 8200 -37955 8235
rect -37945 8200 -37910 8235
rect -37900 8200 -37865 8235
rect -37855 8200 -37820 8235
rect -37810 8200 -37775 8235
rect -37765 8200 -37730 8235
rect -37720 8200 -37685 8235
rect -37675 8200 -37640 8235
rect -37630 8200 -37595 8235
rect -37585 8200 -37550 8235
rect -37540 8200 -37505 8235
rect -37495 8200 -37460 8235
rect -37450 8200 -37415 8235
rect -37405 8200 -37370 8235
rect -37360 8200 -37325 8235
rect -37315 8200 -37280 8235
rect -37270 8200 -37235 8235
rect -37225 8200 -37190 8235
rect -38755 8155 -38720 8190
rect -38710 8155 -38675 8190
rect -38665 8155 -38630 8190
rect -38620 8155 -38585 8190
rect -38575 8155 -38540 8190
rect -38530 8155 -38495 8190
rect -38485 8155 -38450 8190
rect -38440 8155 -38405 8190
rect -38395 8155 -38360 8190
rect -38350 8155 -38315 8190
rect -38305 8155 -38270 8190
rect -38260 8155 -38225 8190
rect -38215 8155 -38180 8190
rect -38170 8155 -38135 8190
rect -38125 8155 -38090 8190
rect -38080 8155 -38045 8190
rect -38035 8155 -38000 8190
rect -37990 8155 -37955 8190
rect -37945 8155 -37910 8190
rect -37900 8155 -37865 8190
rect -37855 8155 -37820 8190
rect -37810 8155 -37775 8190
rect -37765 8155 -37730 8190
rect -37720 8155 -37685 8190
rect -37675 8155 -37640 8190
rect -37630 8155 -37595 8190
rect -37585 8155 -37550 8190
rect -37540 8155 -37505 8190
rect -37495 8155 -37460 8190
rect -37450 8155 -37415 8190
rect -37405 8155 -37370 8190
rect -37360 8155 -37325 8190
rect -37315 8155 -37280 8190
rect -37270 8155 -37235 8190
rect -37225 8155 -37190 8190
rect -38755 8110 -38720 8145
rect -38710 8110 -38675 8145
rect -38665 8110 -38630 8145
rect -38620 8110 -38585 8145
rect -38575 8110 -38540 8145
rect -38530 8110 -38495 8145
rect -38485 8110 -38450 8145
rect -38440 8110 -38405 8145
rect -38395 8110 -38360 8145
rect -38350 8110 -38315 8145
rect -38305 8110 -38270 8145
rect -38260 8110 -38225 8145
rect -38215 8110 -38180 8145
rect -38170 8110 -38135 8145
rect -38125 8110 -38090 8145
rect -38080 8110 -38045 8145
rect -38035 8110 -38000 8145
rect -37990 8110 -37955 8145
rect -37945 8110 -37910 8145
rect -37900 8110 -37865 8145
rect -37855 8110 -37820 8145
rect -37810 8110 -37775 8145
rect -37765 8110 -37730 8145
rect -37720 8110 -37685 8145
rect -37675 8110 -37640 8145
rect -37630 8110 -37595 8145
rect -37585 8110 -37550 8145
rect -37540 8110 -37505 8145
rect -37495 8110 -37460 8145
rect -37450 8110 -37415 8145
rect -37405 8110 -37370 8145
rect -37360 8110 -37325 8145
rect -37315 8110 -37280 8145
rect -37270 8110 -37235 8145
rect -37225 8110 -37190 8145
rect 1320 9635 1360 9640
rect 1320 9605 1325 9635
rect 1325 9605 1355 9635
rect 1355 9605 1360 9635
rect 1320 9600 1360 9605
rect 1320 9570 1360 9575
rect 1320 9540 1325 9570
rect 1325 9540 1355 9570
rect 1355 9540 1360 9570
rect 1320 9535 1360 9540
rect 1320 9500 1360 9505
rect 1320 9470 1325 9500
rect 1325 9470 1355 9500
rect 1355 9470 1360 9500
rect 1320 9465 1360 9470
rect 1320 9430 1360 9435
rect 1320 9400 1325 9430
rect 1325 9400 1355 9430
rect 1355 9400 1360 9430
rect 1320 9395 1360 9400
rect 1320 9360 1360 9365
rect 1320 9330 1325 9360
rect 1325 9330 1355 9360
rect 1355 9330 1360 9360
rect 1320 9325 1360 9330
rect 1320 9295 1360 9300
rect 1320 9265 1325 9295
rect 1325 9265 1355 9295
rect 1355 9265 1360 9295
rect 1320 9260 1360 9265
rect 1320 9235 1360 9240
rect 1320 9205 1325 9235
rect 1325 9205 1355 9235
rect 1355 9205 1360 9235
rect 1320 9200 1360 9205
rect 1320 9170 1360 9175
rect 1320 9140 1325 9170
rect 1325 9140 1355 9170
rect 1355 9140 1360 9170
rect 1320 9135 1360 9140
rect 1320 9100 1360 9105
rect 1320 9070 1325 9100
rect 1325 9070 1355 9100
rect 1355 9070 1360 9100
rect 1320 9065 1360 9070
rect 1320 9030 1360 9035
rect 1320 9000 1325 9030
rect 1325 9000 1355 9030
rect 1355 9000 1360 9030
rect 1320 8995 1360 9000
rect 1320 8960 1360 8965
rect 1320 8930 1325 8960
rect 1325 8930 1355 8960
rect 1355 8930 1360 8960
rect 1320 8925 1360 8930
rect 1320 8895 1360 8900
rect 1320 8865 1325 8895
rect 1325 8865 1355 8895
rect 1355 8865 1360 8895
rect 1320 8860 1360 8865
rect 1320 8835 1360 8840
rect 1320 8805 1325 8835
rect 1325 8805 1355 8835
rect 1355 8805 1360 8835
rect 1320 8800 1360 8805
rect 1320 8770 1360 8775
rect 1320 8740 1325 8770
rect 1325 8740 1355 8770
rect 1355 8740 1360 8770
rect 1320 8735 1360 8740
rect 1320 8700 1360 8705
rect 1320 8670 1325 8700
rect 1325 8670 1355 8700
rect 1355 8670 1360 8700
rect 1320 8665 1360 8670
rect 1320 8630 1360 8635
rect 1320 8600 1325 8630
rect 1325 8600 1355 8630
rect 1355 8600 1360 8630
rect 1320 8595 1360 8600
rect 1320 8560 1360 8565
rect 1320 8530 1325 8560
rect 1325 8530 1355 8560
rect 1355 8530 1360 8560
rect 1320 8525 1360 8530
rect 1320 8495 1360 8500
rect 1320 8465 1325 8495
rect 1325 8465 1355 8495
rect 1355 8465 1360 8495
rect 1320 8460 1360 8465
rect 1320 8435 1360 8440
rect 1320 8405 1325 8435
rect 1325 8405 1355 8435
rect 1355 8405 1360 8435
rect 1320 8400 1360 8405
rect 1320 8370 1360 8375
rect 1320 8340 1325 8370
rect 1325 8340 1355 8370
rect 1355 8340 1360 8370
rect 1320 8335 1360 8340
rect 1320 8300 1360 8305
rect 1320 8270 1325 8300
rect 1325 8270 1355 8300
rect 1355 8270 1360 8300
rect 1320 8265 1360 8270
rect 1320 8230 1360 8235
rect 1320 8200 1325 8230
rect 1325 8200 1355 8230
rect 1355 8200 1360 8230
rect 1320 8195 1360 8200
rect 1320 8160 1360 8165
rect 1320 8130 1325 8160
rect 1325 8130 1355 8160
rect 1355 8130 1360 8160
rect 1320 8125 1360 8130
rect 2245 9635 2285 9640
rect 2245 9605 2250 9635
rect 2250 9605 2280 9635
rect 2280 9605 2285 9635
rect 2245 9600 2285 9605
rect 2245 9570 2285 9575
rect 2245 9540 2250 9570
rect 2250 9540 2280 9570
rect 2280 9540 2285 9570
rect 2245 9535 2285 9540
rect 2245 9500 2285 9505
rect 2245 9470 2250 9500
rect 2250 9470 2280 9500
rect 2280 9470 2285 9500
rect 2245 9465 2285 9470
rect 2245 9430 2285 9435
rect 2245 9400 2250 9430
rect 2250 9400 2280 9430
rect 2280 9400 2285 9430
rect 2245 9395 2285 9400
rect 2245 9360 2285 9365
rect 2245 9330 2250 9360
rect 2250 9330 2280 9360
rect 2280 9330 2285 9360
rect 2245 9325 2285 9330
rect 2245 9295 2285 9300
rect 2245 9265 2250 9295
rect 2250 9265 2280 9295
rect 2280 9265 2285 9295
rect 2245 9260 2285 9265
rect 2245 9235 2285 9240
rect 2245 9205 2250 9235
rect 2250 9205 2280 9235
rect 2280 9205 2285 9235
rect 2245 9200 2285 9205
rect 2245 9170 2285 9175
rect 2245 9140 2250 9170
rect 2250 9140 2280 9170
rect 2280 9140 2285 9170
rect 2245 9135 2285 9140
rect 2245 9100 2285 9105
rect 2245 9070 2250 9100
rect 2250 9070 2280 9100
rect 2280 9070 2285 9100
rect 2245 9065 2285 9070
rect 2245 9030 2285 9035
rect 2245 9000 2250 9030
rect 2250 9000 2280 9030
rect 2280 9000 2285 9030
rect 2245 8995 2285 9000
rect 2245 8960 2285 8965
rect 2245 8930 2250 8960
rect 2250 8930 2280 8960
rect 2280 8930 2285 8960
rect 2245 8925 2285 8930
rect 2245 8895 2285 8900
rect 2245 8865 2250 8895
rect 2250 8865 2280 8895
rect 2280 8865 2285 8895
rect 2245 8860 2285 8865
rect 2245 8835 2285 8840
rect 2245 8805 2250 8835
rect 2250 8805 2280 8835
rect 2280 8805 2285 8835
rect 2245 8800 2285 8805
rect 2245 8770 2285 8775
rect 2245 8740 2250 8770
rect 2250 8740 2280 8770
rect 2280 8740 2285 8770
rect 2245 8735 2285 8740
rect 2245 8700 2285 8705
rect 2245 8670 2250 8700
rect 2250 8670 2280 8700
rect 2280 8670 2285 8700
rect 2245 8665 2285 8670
rect 2245 8630 2285 8635
rect 2245 8600 2250 8630
rect 2250 8600 2280 8630
rect 2280 8600 2285 8630
rect 2245 8595 2285 8600
rect 2245 8560 2285 8565
rect 2245 8530 2250 8560
rect 2250 8530 2280 8560
rect 2280 8530 2285 8560
rect 2245 8525 2285 8530
rect 2245 8495 2285 8500
rect 2245 8465 2250 8495
rect 2250 8465 2280 8495
rect 2280 8465 2285 8495
rect 2245 8460 2285 8465
rect 2245 8435 2285 8440
rect 2245 8405 2250 8435
rect 2250 8405 2280 8435
rect 2280 8405 2285 8435
rect 2245 8400 2285 8405
rect 2245 8370 2285 8375
rect 2245 8340 2250 8370
rect 2250 8340 2280 8370
rect 2280 8340 2285 8370
rect 2245 8335 2285 8340
rect 2245 8300 2285 8305
rect 2245 8270 2250 8300
rect 2250 8270 2280 8300
rect 2280 8270 2285 8300
rect 2245 8265 2285 8270
rect 2245 8230 2285 8235
rect 2245 8200 2250 8230
rect 2250 8200 2280 8230
rect 2280 8200 2285 8230
rect 2245 8195 2285 8200
rect 2245 8160 2285 8165
rect 2245 8130 2250 8160
rect 2250 8130 2280 8160
rect 2280 8130 2285 8160
rect 2245 8125 2285 8130
rect 6700 9635 6740 9640
rect 6700 9605 6705 9635
rect 6705 9605 6735 9635
rect 6735 9605 6740 9635
rect 6700 9600 6740 9605
rect 6700 9570 6740 9575
rect 6700 9540 6705 9570
rect 6705 9540 6735 9570
rect 6735 9540 6740 9570
rect 6700 9535 6740 9540
rect 6700 9500 6740 9505
rect 6700 9470 6705 9500
rect 6705 9470 6735 9500
rect 6735 9470 6740 9500
rect 6700 9465 6740 9470
rect 6700 9430 6740 9435
rect 6700 9400 6705 9430
rect 6705 9400 6735 9430
rect 6735 9400 6740 9430
rect 6700 9395 6740 9400
rect 6700 9360 6740 9365
rect 6700 9330 6705 9360
rect 6705 9330 6735 9360
rect 6735 9330 6740 9360
rect 6700 9325 6740 9330
rect 6700 9295 6740 9300
rect 6700 9265 6705 9295
rect 6705 9265 6735 9295
rect 6735 9265 6740 9295
rect 6700 9260 6740 9265
rect 6700 9235 6740 9240
rect 6700 9205 6705 9235
rect 6705 9205 6735 9235
rect 6735 9205 6740 9235
rect 6700 9200 6740 9205
rect 6700 9170 6740 9175
rect 6700 9140 6705 9170
rect 6705 9140 6735 9170
rect 6735 9140 6740 9170
rect 6700 9135 6740 9140
rect 6700 9100 6740 9105
rect 6700 9070 6705 9100
rect 6705 9070 6735 9100
rect 6735 9070 6740 9100
rect 6700 9065 6740 9070
rect 6700 9030 6740 9035
rect 6700 9000 6705 9030
rect 6705 9000 6735 9030
rect 6735 9000 6740 9030
rect 6700 8995 6740 9000
rect 6700 8960 6740 8965
rect 6700 8930 6705 8960
rect 6705 8930 6735 8960
rect 6735 8930 6740 8960
rect 6700 8925 6740 8930
rect 6700 8895 6740 8900
rect 6700 8865 6705 8895
rect 6705 8865 6735 8895
rect 6735 8865 6740 8895
rect 6700 8860 6740 8865
rect 6700 8835 6740 8840
rect 6700 8805 6705 8835
rect 6705 8805 6735 8835
rect 6735 8805 6740 8835
rect 6700 8800 6740 8805
rect 6700 8770 6740 8775
rect 6700 8740 6705 8770
rect 6705 8740 6735 8770
rect 6735 8740 6740 8770
rect 6700 8735 6740 8740
rect 6700 8700 6740 8705
rect 6700 8670 6705 8700
rect 6705 8670 6735 8700
rect 6735 8670 6740 8700
rect 6700 8665 6740 8670
rect 6700 8630 6740 8635
rect 6700 8600 6705 8630
rect 6705 8600 6735 8630
rect 6735 8600 6740 8630
rect 6700 8595 6740 8600
rect 6700 8560 6740 8565
rect 6700 8530 6705 8560
rect 6705 8530 6735 8560
rect 6735 8530 6740 8560
rect 6700 8525 6740 8530
rect 6700 8495 6740 8500
rect 6700 8465 6705 8495
rect 6705 8465 6735 8495
rect 6735 8465 6740 8495
rect 6700 8460 6740 8465
rect 6700 8435 6740 8440
rect 6700 8405 6705 8435
rect 6705 8405 6735 8435
rect 6735 8405 6740 8435
rect 6700 8400 6740 8405
rect 6700 8370 6740 8375
rect 6700 8340 6705 8370
rect 6705 8340 6735 8370
rect 6735 8340 6740 8370
rect 6700 8335 6740 8340
rect 6700 8300 6740 8305
rect 6700 8270 6705 8300
rect 6705 8270 6735 8300
rect 6735 8270 6740 8300
rect 6700 8265 6740 8270
rect 6700 8230 6740 8235
rect 6700 8200 6705 8230
rect 6705 8200 6735 8230
rect 6735 8200 6740 8230
rect 6700 8195 6740 8200
rect 6700 8160 6740 8165
rect 6700 8130 6705 8160
rect 6705 8130 6735 8160
rect 6735 8130 6740 8160
rect 6700 8125 6740 8130
rect 7620 9635 7660 9640
rect 7620 9605 7625 9635
rect 7625 9605 7655 9635
rect 7655 9605 7660 9635
rect 7620 9600 7660 9605
rect 7620 9570 7660 9575
rect 7620 9540 7625 9570
rect 7625 9540 7655 9570
rect 7655 9540 7660 9570
rect 7620 9535 7660 9540
rect 7620 9500 7660 9505
rect 7620 9470 7625 9500
rect 7625 9470 7655 9500
rect 7655 9470 7660 9500
rect 7620 9465 7660 9470
rect 7620 9430 7660 9435
rect 7620 9400 7625 9430
rect 7625 9400 7655 9430
rect 7655 9400 7660 9430
rect 7620 9395 7660 9400
rect 7620 9360 7660 9365
rect 7620 9330 7625 9360
rect 7625 9330 7655 9360
rect 7655 9330 7660 9360
rect 7620 9325 7660 9330
rect 7620 9295 7660 9300
rect 7620 9265 7625 9295
rect 7625 9265 7655 9295
rect 7655 9265 7660 9295
rect 7620 9260 7660 9265
rect 7620 9235 7660 9240
rect 7620 9205 7625 9235
rect 7625 9205 7655 9235
rect 7655 9205 7660 9235
rect 7620 9200 7660 9205
rect 7620 9170 7660 9175
rect 7620 9140 7625 9170
rect 7625 9140 7655 9170
rect 7655 9140 7660 9170
rect 7620 9135 7660 9140
rect 7620 9100 7660 9105
rect 7620 9070 7625 9100
rect 7625 9070 7655 9100
rect 7655 9070 7660 9100
rect 7620 9065 7660 9070
rect 7620 9030 7660 9035
rect 7620 9000 7625 9030
rect 7625 9000 7655 9030
rect 7655 9000 7660 9030
rect 7620 8995 7660 9000
rect 7620 8960 7660 8965
rect 7620 8930 7625 8960
rect 7625 8930 7655 8960
rect 7655 8930 7660 8960
rect 7620 8925 7660 8930
rect 7620 8895 7660 8900
rect 7620 8865 7625 8895
rect 7625 8865 7655 8895
rect 7655 8865 7660 8895
rect 7620 8860 7660 8865
rect 7620 8835 7660 8840
rect 7620 8805 7625 8835
rect 7625 8805 7655 8835
rect 7655 8805 7660 8835
rect 7620 8800 7660 8805
rect 7620 8770 7660 8775
rect 7620 8740 7625 8770
rect 7625 8740 7655 8770
rect 7655 8740 7660 8770
rect 7620 8735 7660 8740
rect 7620 8700 7660 8705
rect 7620 8670 7625 8700
rect 7625 8670 7655 8700
rect 7655 8670 7660 8700
rect 7620 8665 7660 8670
rect 7620 8630 7660 8635
rect 7620 8600 7625 8630
rect 7625 8600 7655 8630
rect 7655 8600 7660 8630
rect 7620 8595 7660 8600
rect 7620 8560 7660 8565
rect 7620 8530 7625 8560
rect 7625 8530 7655 8560
rect 7655 8530 7660 8560
rect 7620 8525 7660 8530
rect 7620 8495 7660 8500
rect 7620 8465 7625 8495
rect 7625 8465 7655 8495
rect 7655 8465 7660 8495
rect 7620 8460 7660 8465
rect 7620 8435 7660 8440
rect 7620 8405 7625 8435
rect 7625 8405 7655 8435
rect 7655 8405 7660 8435
rect 7620 8400 7660 8405
rect 7620 8370 7660 8375
rect 7620 8340 7625 8370
rect 7625 8340 7655 8370
rect 7655 8340 7660 8370
rect 7620 8335 7660 8340
rect 7620 8300 7660 8305
rect 7620 8270 7625 8300
rect 7625 8270 7655 8300
rect 7655 8270 7660 8300
rect 7620 8265 7660 8270
rect 7620 8230 7660 8235
rect 7620 8200 7625 8230
rect 7625 8200 7655 8230
rect 7655 8200 7660 8230
rect 7620 8195 7660 8200
rect 7620 8160 7660 8165
rect 7620 8130 7625 8160
rect 7625 8130 7655 8160
rect 7655 8130 7660 8160
rect 7620 8125 7660 8130
rect 31305 7995 31340 8030
rect 31350 7995 31385 8030
rect 31395 7995 31430 8030
rect 31440 7995 31475 8030
rect 31485 7995 31520 8030
rect 31530 7995 31565 8030
rect 31575 7995 31610 8030
rect 31620 7995 31655 8030
rect 31665 7995 31700 8030
rect 31710 7995 31745 8030
rect 31755 7995 31790 8030
rect 31800 7995 31835 8030
rect 31845 7995 31880 8030
rect 31890 7995 31925 8030
rect 31935 7995 31970 8030
rect 31980 7995 32015 8030
rect 32025 7995 32060 8030
rect 32070 7995 32105 8030
rect 32115 7995 32150 8030
rect 32160 7995 32195 8030
rect 32205 7995 32240 8030
rect 32250 7995 32285 8030
rect 32295 7995 32330 8030
rect 32340 7995 32375 8030
rect 32385 7995 32420 8030
rect 32430 7995 32465 8030
rect 32475 7995 32510 8030
rect 32520 7995 32555 8030
rect 32565 7995 32600 8030
rect 32610 7995 32645 8030
rect 32655 7995 32690 8030
rect 32700 7995 32735 8030
rect 32745 7995 32780 8030
rect 32790 7995 32825 8030
rect 32835 7995 32870 8030
rect -38755 7935 -38720 7970
rect -38710 7935 -38675 7970
rect -38665 7935 -38630 7970
rect -38620 7935 -38585 7970
rect -38575 7935 -38540 7970
rect -38530 7935 -38495 7970
rect -38485 7935 -38450 7970
rect -38440 7935 -38405 7970
rect -38395 7935 -38360 7970
rect -38350 7935 -38315 7970
rect -38305 7935 -38270 7970
rect -38260 7935 -38225 7970
rect -38215 7935 -38180 7970
rect -38170 7935 -38135 7970
rect -38125 7935 -38090 7970
rect -38080 7935 -38045 7970
rect -38035 7935 -38000 7970
rect -37990 7935 -37955 7970
rect -37945 7935 -37910 7970
rect -37900 7935 -37865 7970
rect -37855 7935 -37820 7970
rect -37810 7935 -37775 7970
rect -37765 7935 -37730 7970
rect -37720 7935 -37685 7970
rect -37675 7935 -37640 7970
rect -37630 7935 -37595 7970
rect -37585 7935 -37550 7970
rect -37540 7935 -37505 7970
rect -37495 7935 -37460 7970
rect -37450 7935 -37415 7970
rect -37405 7935 -37370 7970
rect -37360 7935 -37325 7970
rect -37315 7935 -37280 7970
rect -37270 7935 -37235 7970
rect -37225 7935 -37190 7970
rect -38755 7890 -38720 7925
rect -38710 7890 -38675 7925
rect -38665 7890 -38630 7925
rect -38620 7890 -38585 7925
rect -38575 7890 -38540 7925
rect -38530 7890 -38495 7925
rect -38485 7890 -38450 7925
rect -38440 7890 -38405 7925
rect -38395 7890 -38360 7925
rect -38350 7890 -38315 7925
rect -38305 7890 -38270 7925
rect -38260 7890 -38225 7925
rect -38215 7890 -38180 7925
rect -38170 7890 -38135 7925
rect -38125 7890 -38090 7925
rect -38080 7890 -38045 7925
rect -38035 7890 -38000 7925
rect -37990 7890 -37955 7925
rect -37945 7890 -37910 7925
rect -37900 7890 -37865 7925
rect -37855 7890 -37820 7925
rect -37810 7890 -37775 7925
rect -37765 7890 -37730 7925
rect -37720 7890 -37685 7925
rect -37675 7890 -37640 7925
rect -37630 7890 -37595 7925
rect -37585 7890 -37550 7925
rect -37540 7890 -37505 7925
rect -37495 7890 -37460 7925
rect -37450 7890 -37415 7925
rect -37405 7890 -37370 7925
rect -37360 7890 -37325 7925
rect -37315 7890 -37280 7925
rect -37270 7890 -37235 7925
rect -37225 7890 -37190 7925
rect -38755 7845 -38720 7880
rect -38710 7845 -38675 7880
rect -38665 7845 -38630 7880
rect -38620 7845 -38585 7880
rect -38575 7845 -38540 7880
rect -38530 7845 -38495 7880
rect -38485 7845 -38450 7880
rect -38440 7845 -38405 7880
rect -38395 7845 -38360 7880
rect -38350 7845 -38315 7880
rect -38305 7845 -38270 7880
rect -38260 7845 -38225 7880
rect -38215 7845 -38180 7880
rect -38170 7845 -38135 7880
rect -38125 7845 -38090 7880
rect -38080 7845 -38045 7880
rect -38035 7845 -38000 7880
rect -37990 7845 -37955 7880
rect -37945 7845 -37910 7880
rect -37900 7845 -37865 7880
rect -37855 7845 -37820 7880
rect -37810 7845 -37775 7880
rect -37765 7845 -37730 7880
rect -37720 7845 -37685 7880
rect -37675 7845 -37640 7880
rect -37630 7845 -37595 7880
rect -37585 7845 -37550 7880
rect -37540 7845 -37505 7880
rect -37495 7845 -37460 7880
rect -37450 7845 -37415 7880
rect -37405 7845 -37370 7880
rect -37360 7845 -37325 7880
rect -37315 7845 -37280 7880
rect -37270 7845 -37235 7880
rect -37225 7845 -37190 7880
rect -38755 7800 -38720 7835
rect -38710 7800 -38675 7835
rect -38665 7800 -38630 7835
rect -38620 7800 -38585 7835
rect -38575 7800 -38540 7835
rect -38530 7800 -38495 7835
rect -38485 7800 -38450 7835
rect -38440 7800 -38405 7835
rect -38395 7800 -38360 7835
rect -38350 7800 -38315 7835
rect -38305 7800 -38270 7835
rect -38260 7800 -38225 7835
rect -38215 7800 -38180 7835
rect -38170 7800 -38135 7835
rect -38125 7800 -38090 7835
rect -38080 7800 -38045 7835
rect -38035 7800 -38000 7835
rect -37990 7800 -37955 7835
rect -37945 7800 -37910 7835
rect -37900 7800 -37865 7835
rect -37855 7800 -37820 7835
rect -37810 7800 -37775 7835
rect -37765 7800 -37730 7835
rect -37720 7800 -37685 7835
rect -37675 7800 -37640 7835
rect -37630 7800 -37595 7835
rect -37585 7800 -37550 7835
rect -37540 7800 -37505 7835
rect -37495 7800 -37460 7835
rect -37450 7800 -37415 7835
rect -37405 7800 -37370 7835
rect -37360 7800 -37325 7835
rect -37315 7800 -37280 7835
rect -37270 7800 -37235 7835
rect -37225 7800 -37190 7835
rect -38755 7755 -38720 7790
rect -38710 7755 -38675 7790
rect -38665 7755 -38630 7790
rect -38620 7755 -38585 7790
rect -38575 7755 -38540 7790
rect -38530 7755 -38495 7790
rect -38485 7755 -38450 7790
rect -38440 7755 -38405 7790
rect -38395 7755 -38360 7790
rect -38350 7755 -38315 7790
rect -38305 7755 -38270 7790
rect -38260 7755 -38225 7790
rect -38215 7755 -38180 7790
rect -38170 7755 -38135 7790
rect -38125 7755 -38090 7790
rect -38080 7755 -38045 7790
rect -38035 7755 -38000 7790
rect -37990 7755 -37955 7790
rect -37945 7755 -37910 7790
rect -37900 7755 -37865 7790
rect -37855 7755 -37820 7790
rect -37810 7755 -37775 7790
rect -37765 7755 -37730 7790
rect -37720 7755 -37685 7790
rect -37675 7755 -37640 7790
rect -37630 7755 -37595 7790
rect -37585 7755 -37550 7790
rect -37540 7755 -37505 7790
rect -37495 7755 -37460 7790
rect -37450 7755 -37415 7790
rect -37405 7755 -37370 7790
rect -37360 7755 -37325 7790
rect -37315 7755 -37280 7790
rect -37270 7755 -37235 7790
rect -37225 7755 -37190 7790
rect -38755 7710 -38720 7745
rect -38710 7710 -38675 7745
rect -38665 7710 -38630 7745
rect -38620 7710 -38585 7745
rect -38575 7710 -38540 7745
rect -38530 7710 -38495 7745
rect -38485 7710 -38450 7745
rect -38440 7710 -38405 7745
rect -38395 7710 -38360 7745
rect -38350 7710 -38315 7745
rect -38305 7710 -38270 7745
rect -38260 7710 -38225 7745
rect -38215 7710 -38180 7745
rect -38170 7710 -38135 7745
rect -38125 7710 -38090 7745
rect -38080 7710 -38045 7745
rect -38035 7710 -38000 7745
rect -37990 7710 -37955 7745
rect -37945 7710 -37910 7745
rect -37900 7710 -37865 7745
rect -37855 7710 -37820 7745
rect -37810 7710 -37775 7745
rect -37765 7710 -37730 7745
rect -37720 7710 -37685 7745
rect -37675 7710 -37640 7745
rect -37630 7710 -37595 7745
rect -37585 7710 -37550 7745
rect -37540 7710 -37505 7745
rect -37495 7710 -37460 7745
rect -37450 7710 -37415 7745
rect -37405 7710 -37370 7745
rect -37360 7710 -37325 7745
rect -37315 7710 -37280 7745
rect -37270 7710 -37235 7745
rect -37225 7710 -37190 7745
rect -38755 7665 -38720 7700
rect -38710 7665 -38675 7700
rect -38665 7665 -38630 7700
rect -38620 7665 -38585 7700
rect -38575 7665 -38540 7700
rect -38530 7665 -38495 7700
rect -38485 7665 -38450 7700
rect -38440 7665 -38405 7700
rect -38395 7665 -38360 7700
rect -38350 7665 -38315 7700
rect -38305 7665 -38270 7700
rect -38260 7665 -38225 7700
rect -38215 7665 -38180 7700
rect -38170 7665 -38135 7700
rect -38125 7665 -38090 7700
rect -38080 7665 -38045 7700
rect -38035 7665 -38000 7700
rect -37990 7665 -37955 7700
rect -37945 7665 -37910 7700
rect -37900 7665 -37865 7700
rect -37855 7665 -37820 7700
rect -37810 7665 -37775 7700
rect -37765 7665 -37730 7700
rect -37720 7665 -37685 7700
rect -37675 7665 -37640 7700
rect -37630 7665 -37595 7700
rect -37585 7665 -37550 7700
rect -37540 7665 -37505 7700
rect -37495 7665 -37460 7700
rect -37450 7665 -37415 7700
rect -37405 7665 -37370 7700
rect -37360 7665 -37325 7700
rect -37315 7665 -37280 7700
rect -37270 7665 -37235 7700
rect -37225 7665 -37190 7700
rect -38755 7620 -38720 7655
rect -38710 7620 -38675 7655
rect -38665 7620 -38630 7655
rect -38620 7620 -38585 7655
rect -38575 7620 -38540 7655
rect -38530 7620 -38495 7655
rect -38485 7620 -38450 7655
rect -38440 7620 -38405 7655
rect -38395 7620 -38360 7655
rect -38350 7620 -38315 7655
rect -38305 7620 -38270 7655
rect -38260 7620 -38225 7655
rect -38215 7620 -38180 7655
rect -38170 7620 -38135 7655
rect -38125 7620 -38090 7655
rect -38080 7620 -38045 7655
rect -38035 7620 -38000 7655
rect -37990 7620 -37955 7655
rect -37945 7620 -37910 7655
rect -37900 7620 -37865 7655
rect -37855 7620 -37820 7655
rect -37810 7620 -37775 7655
rect -37765 7620 -37730 7655
rect -37720 7620 -37685 7655
rect -37675 7620 -37640 7655
rect -37630 7620 -37595 7655
rect -37585 7620 -37550 7655
rect -37540 7620 -37505 7655
rect -37495 7620 -37460 7655
rect -37450 7620 -37415 7655
rect -37405 7620 -37370 7655
rect -37360 7620 -37325 7655
rect -37315 7620 -37280 7655
rect -37270 7620 -37235 7655
rect -37225 7620 -37190 7655
rect -38755 7575 -38720 7610
rect -38710 7575 -38675 7610
rect -38665 7575 -38630 7610
rect -38620 7575 -38585 7610
rect -38575 7575 -38540 7610
rect -38530 7575 -38495 7610
rect -38485 7575 -38450 7610
rect -38440 7575 -38405 7610
rect -38395 7575 -38360 7610
rect -38350 7575 -38315 7610
rect -38305 7575 -38270 7610
rect -38260 7575 -38225 7610
rect -38215 7575 -38180 7610
rect -38170 7575 -38135 7610
rect -38125 7575 -38090 7610
rect -38080 7575 -38045 7610
rect -38035 7575 -38000 7610
rect -37990 7575 -37955 7610
rect -37945 7575 -37910 7610
rect -37900 7575 -37865 7610
rect -37855 7575 -37820 7610
rect -37810 7575 -37775 7610
rect -37765 7575 -37730 7610
rect -37720 7575 -37685 7610
rect -37675 7575 -37640 7610
rect -37630 7575 -37595 7610
rect -37585 7575 -37550 7610
rect -37540 7575 -37505 7610
rect -37495 7575 -37460 7610
rect -37450 7575 -37415 7610
rect -37405 7575 -37370 7610
rect -37360 7575 -37325 7610
rect -37315 7575 -37280 7610
rect -37270 7575 -37235 7610
rect -37225 7575 -37190 7610
rect -38755 7530 -38720 7565
rect -38710 7530 -38675 7565
rect -38665 7530 -38630 7565
rect -38620 7530 -38585 7565
rect -38575 7530 -38540 7565
rect -38530 7530 -38495 7565
rect -38485 7530 -38450 7565
rect -38440 7530 -38405 7565
rect -38395 7530 -38360 7565
rect -38350 7530 -38315 7565
rect -38305 7530 -38270 7565
rect -38260 7530 -38225 7565
rect -38215 7530 -38180 7565
rect -38170 7530 -38135 7565
rect -38125 7530 -38090 7565
rect -38080 7530 -38045 7565
rect -38035 7530 -38000 7565
rect -37990 7530 -37955 7565
rect -37945 7530 -37910 7565
rect -37900 7530 -37865 7565
rect -37855 7530 -37820 7565
rect -37810 7530 -37775 7565
rect -37765 7530 -37730 7565
rect -37720 7530 -37685 7565
rect -37675 7530 -37640 7565
rect -37630 7530 -37595 7565
rect -37585 7530 -37550 7565
rect -37540 7530 -37505 7565
rect -37495 7530 -37460 7565
rect -37450 7530 -37415 7565
rect -37405 7530 -37370 7565
rect -37360 7530 -37325 7565
rect -37315 7530 -37280 7565
rect -37270 7530 -37235 7565
rect -37225 7530 -37190 7565
rect -38755 7485 -38720 7520
rect -38710 7485 -38675 7520
rect -38665 7485 -38630 7520
rect -38620 7485 -38585 7520
rect -38575 7485 -38540 7520
rect -38530 7485 -38495 7520
rect -38485 7485 -38450 7520
rect -38440 7485 -38405 7520
rect -38395 7485 -38360 7520
rect -38350 7485 -38315 7520
rect -38305 7485 -38270 7520
rect -38260 7485 -38225 7520
rect -38215 7485 -38180 7520
rect -38170 7485 -38135 7520
rect -38125 7485 -38090 7520
rect -38080 7485 -38045 7520
rect -38035 7485 -38000 7520
rect -37990 7485 -37955 7520
rect -37945 7485 -37910 7520
rect -37900 7485 -37865 7520
rect -37855 7485 -37820 7520
rect -37810 7485 -37775 7520
rect -37765 7485 -37730 7520
rect -37720 7485 -37685 7520
rect -37675 7485 -37640 7520
rect -37630 7485 -37595 7520
rect -37585 7485 -37550 7520
rect -37540 7485 -37505 7520
rect -37495 7485 -37460 7520
rect -37450 7485 -37415 7520
rect -37405 7485 -37370 7520
rect -37360 7485 -37325 7520
rect -37315 7485 -37280 7520
rect -37270 7485 -37235 7520
rect -37225 7485 -37190 7520
rect -38755 7440 -38720 7475
rect -38710 7440 -38675 7475
rect -38665 7440 -38630 7475
rect -38620 7440 -38585 7475
rect -38575 7440 -38540 7475
rect -38530 7440 -38495 7475
rect -38485 7440 -38450 7475
rect -38440 7440 -38405 7475
rect -38395 7440 -38360 7475
rect -38350 7440 -38315 7475
rect -38305 7440 -38270 7475
rect -38260 7440 -38225 7475
rect -38215 7440 -38180 7475
rect -38170 7440 -38135 7475
rect -38125 7440 -38090 7475
rect -38080 7440 -38045 7475
rect -38035 7440 -38000 7475
rect -37990 7440 -37955 7475
rect -37945 7440 -37910 7475
rect -37900 7440 -37865 7475
rect -37855 7440 -37820 7475
rect -37810 7440 -37775 7475
rect -37765 7440 -37730 7475
rect -37720 7440 -37685 7475
rect -37675 7440 -37640 7475
rect -37630 7440 -37595 7475
rect -37585 7440 -37550 7475
rect -37540 7440 -37505 7475
rect -37495 7440 -37460 7475
rect -37450 7440 -37415 7475
rect -37405 7440 -37370 7475
rect -37360 7440 -37325 7475
rect -37315 7440 -37280 7475
rect -37270 7440 -37235 7475
rect -37225 7440 -37190 7475
rect -38755 7395 -38720 7430
rect -38710 7395 -38675 7430
rect -38665 7395 -38630 7430
rect -38620 7395 -38585 7430
rect -38575 7395 -38540 7430
rect -38530 7395 -38495 7430
rect -38485 7395 -38450 7430
rect -38440 7395 -38405 7430
rect -38395 7395 -38360 7430
rect -38350 7395 -38315 7430
rect -38305 7395 -38270 7430
rect -38260 7395 -38225 7430
rect -38215 7395 -38180 7430
rect -38170 7395 -38135 7430
rect -38125 7395 -38090 7430
rect -38080 7395 -38045 7430
rect -38035 7395 -38000 7430
rect -37990 7395 -37955 7430
rect -37945 7395 -37910 7430
rect -37900 7395 -37865 7430
rect -37855 7395 -37820 7430
rect -37810 7395 -37775 7430
rect -37765 7395 -37730 7430
rect -37720 7395 -37685 7430
rect -37675 7395 -37640 7430
rect -37630 7395 -37595 7430
rect -37585 7395 -37550 7430
rect -37540 7395 -37505 7430
rect -37495 7395 -37460 7430
rect -37450 7395 -37415 7430
rect -37405 7395 -37370 7430
rect -37360 7395 -37325 7430
rect -37315 7395 -37280 7430
rect -37270 7395 -37235 7430
rect -37225 7395 -37190 7430
rect -38755 7350 -38720 7385
rect -38710 7350 -38675 7385
rect -38665 7350 -38630 7385
rect -38620 7350 -38585 7385
rect -38575 7350 -38540 7385
rect -38530 7350 -38495 7385
rect -38485 7350 -38450 7385
rect -38440 7350 -38405 7385
rect -38395 7350 -38360 7385
rect -38350 7350 -38315 7385
rect -38305 7350 -38270 7385
rect -38260 7350 -38225 7385
rect -38215 7350 -38180 7385
rect -38170 7350 -38135 7385
rect -38125 7350 -38090 7385
rect -38080 7350 -38045 7385
rect -38035 7350 -38000 7385
rect -37990 7350 -37955 7385
rect -37945 7350 -37910 7385
rect -37900 7350 -37865 7385
rect -37855 7350 -37820 7385
rect -37810 7350 -37775 7385
rect -37765 7350 -37730 7385
rect -37720 7350 -37685 7385
rect -37675 7350 -37640 7385
rect -37630 7350 -37595 7385
rect -37585 7350 -37550 7385
rect -37540 7350 -37505 7385
rect -37495 7350 -37460 7385
rect -37450 7350 -37415 7385
rect -37405 7350 -37370 7385
rect -37360 7350 -37325 7385
rect -37315 7350 -37280 7385
rect -37270 7350 -37235 7385
rect -37225 7350 -37190 7385
rect -38755 7305 -38720 7340
rect -38710 7305 -38675 7340
rect -38665 7305 -38630 7340
rect -38620 7305 -38585 7340
rect -38575 7305 -38540 7340
rect -38530 7305 -38495 7340
rect -38485 7305 -38450 7340
rect -38440 7305 -38405 7340
rect -38395 7305 -38360 7340
rect -38350 7305 -38315 7340
rect -38305 7305 -38270 7340
rect -38260 7305 -38225 7340
rect -38215 7305 -38180 7340
rect -38170 7305 -38135 7340
rect -38125 7305 -38090 7340
rect -38080 7305 -38045 7340
rect -38035 7305 -38000 7340
rect -37990 7305 -37955 7340
rect -37945 7305 -37910 7340
rect -37900 7305 -37865 7340
rect -37855 7305 -37820 7340
rect -37810 7305 -37775 7340
rect -37765 7305 -37730 7340
rect -37720 7305 -37685 7340
rect -37675 7305 -37640 7340
rect -37630 7305 -37595 7340
rect -37585 7305 -37550 7340
rect -37540 7305 -37505 7340
rect -37495 7305 -37460 7340
rect -37450 7305 -37415 7340
rect -37405 7305 -37370 7340
rect -37360 7305 -37325 7340
rect -37315 7305 -37280 7340
rect -37270 7305 -37235 7340
rect -37225 7305 -37190 7340
rect -38755 7260 -38720 7295
rect -38710 7260 -38675 7295
rect -38665 7260 -38630 7295
rect -38620 7260 -38585 7295
rect -38575 7260 -38540 7295
rect -38530 7260 -38495 7295
rect -38485 7260 -38450 7295
rect -38440 7260 -38405 7295
rect -38395 7260 -38360 7295
rect -38350 7260 -38315 7295
rect -38305 7260 -38270 7295
rect -38260 7260 -38225 7295
rect -38215 7260 -38180 7295
rect -38170 7260 -38135 7295
rect -38125 7260 -38090 7295
rect -38080 7260 -38045 7295
rect -38035 7260 -38000 7295
rect -37990 7260 -37955 7295
rect -37945 7260 -37910 7295
rect -37900 7260 -37865 7295
rect -37855 7260 -37820 7295
rect -37810 7260 -37775 7295
rect -37765 7260 -37730 7295
rect -37720 7260 -37685 7295
rect -37675 7260 -37640 7295
rect -37630 7260 -37595 7295
rect -37585 7260 -37550 7295
rect -37540 7260 -37505 7295
rect -37495 7260 -37460 7295
rect -37450 7260 -37415 7295
rect -37405 7260 -37370 7295
rect -37360 7260 -37325 7295
rect -37315 7260 -37280 7295
rect -37270 7260 -37235 7295
rect -37225 7260 -37190 7295
rect -38755 7215 -38720 7250
rect -38710 7215 -38675 7250
rect -38665 7215 -38630 7250
rect -38620 7215 -38585 7250
rect -38575 7215 -38540 7250
rect -38530 7215 -38495 7250
rect -38485 7215 -38450 7250
rect -38440 7215 -38405 7250
rect -38395 7215 -38360 7250
rect -38350 7215 -38315 7250
rect -38305 7215 -38270 7250
rect -38260 7215 -38225 7250
rect -38215 7215 -38180 7250
rect -38170 7215 -38135 7250
rect -38125 7215 -38090 7250
rect -38080 7215 -38045 7250
rect -38035 7215 -38000 7250
rect -37990 7215 -37955 7250
rect -37945 7215 -37910 7250
rect -37900 7215 -37865 7250
rect -37855 7215 -37820 7250
rect -37810 7215 -37775 7250
rect -37765 7215 -37730 7250
rect -37720 7215 -37685 7250
rect -37675 7215 -37640 7250
rect -37630 7215 -37595 7250
rect -37585 7215 -37550 7250
rect -37540 7215 -37505 7250
rect -37495 7215 -37460 7250
rect -37450 7215 -37415 7250
rect -37405 7215 -37370 7250
rect -37360 7215 -37325 7250
rect -37315 7215 -37280 7250
rect -37270 7215 -37235 7250
rect -37225 7215 -37190 7250
rect -38755 7170 -38720 7205
rect -38710 7170 -38675 7205
rect -38665 7170 -38630 7205
rect -38620 7170 -38585 7205
rect -38575 7170 -38540 7205
rect -38530 7170 -38495 7205
rect -38485 7170 -38450 7205
rect -38440 7170 -38405 7205
rect -38395 7170 -38360 7205
rect -38350 7170 -38315 7205
rect -38305 7170 -38270 7205
rect -38260 7170 -38225 7205
rect -38215 7170 -38180 7205
rect -38170 7170 -38135 7205
rect -38125 7170 -38090 7205
rect -38080 7170 -38045 7205
rect -38035 7170 -38000 7205
rect -37990 7170 -37955 7205
rect -37945 7170 -37910 7205
rect -37900 7170 -37865 7205
rect -37855 7170 -37820 7205
rect -37810 7170 -37775 7205
rect -37765 7170 -37730 7205
rect -37720 7170 -37685 7205
rect -37675 7170 -37640 7205
rect -37630 7170 -37595 7205
rect -37585 7170 -37550 7205
rect -37540 7170 -37505 7205
rect -37495 7170 -37460 7205
rect -37450 7170 -37415 7205
rect -37405 7170 -37370 7205
rect -37360 7170 -37325 7205
rect -37315 7170 -37280 7205
rect -37270 7170 -37235 7205
rect -37225 7170 -37190 7205
rect -38755 7125 -38720 7160
rect -38710 7125 -38675 7160
rect -38665 7125 -38630 7160
rect -38620 7125 -38585 7160
rect -38575 7125 -38540 7160
rect -38530 7125 -38495 7160
rect -38485 7125 -38450 7160
rect -38440 7125 -38405 7160
rect -38395 7125 -38360 7160
rect -38350 7125 -38315 7160
rect -38305 7125 -38270 7160
rect -38260 7125 -38225 7160
rect -38215 7125 -38180 7160
rect -38170 7125 -38135 7160
rect -38125 7125 -38090 7160
rect -38080 7125 -38045 7160
rect -38035 7125 -38000 7160
rect -37990 7125 -37955 7160
rect -37945 7125 -37910 7160
rect -37900 7125 -37865 7160
rect -37855 7125 -37820 7160
rect -37810 7125 -37775 7160
rect -37765 7125 -37730 7160
rect -37720 7125 -37685 7160
rect -37675 7125 -37640 7160
rect -37630 7125 -37595 7160
rect -37585 7125 -37550 7160
rect -37540 7125 -37505 7160
rect -37495 7125 -37460 7160
rect -37450 7125 -37415 7160
rect -37405 7125 -37370 7160
rect -37360 7125 -37325 7160
rect -37315 7125 -37280 7160
rect -37270 7125 -37235 7160
rect -37225 7125 -37190 7160
rect -38755 7080 -38720 7115
rect -38710 7080 -38675 7115
rect -38665 7080 -38630 7115
rect -38620 7080 -38585 7115
rect -38575 7080 -38540 7115
rect -38530 7080 -38495 7115
rect -38485 7080 -38450 7115
rect -38440 7080 -38405 7115
rect -38395 7080 -38360 7115
rect -38350 7080 -38315 7115
rect -38305 7080 -38270 7115
rect -38260 7080 -38225 7115
rect -38215 7080 -38180 7115
rect -38170 7080 -38135 7115
rect -38125 7080 -38090 7115
rect -38080 7080 -38045 7115
rect -38035 7080 -38000 7115
rect -37990 7080 -37955 7115
rect -37945 7080 -37910 7115
rect -37900 7080 -37865 7115
rect -37855 7080 -37820 7115
rect -37810 7080 -37775 7115
rect -37765 7080 -37730 7115
rect -37720 7080 -37685 7115
rect -37675 7080 -37640 7115
rect -37630 7080 -37595 7115
rect -37585 7080 -37550 7115
rect -37540 7080 -37505 7115
rect -37495 7080 -37460 7115
rect -37450 7080 -37415 7115
rect -37405 7080 -37370 7115
rect -37360 7080 -37325 7115
rect -37315 7080 -37280 7115
rect -37270 7080 -37235 7115
rect -37225 7080 -37190 7115
rect -38755 7035 -38720 7070
rect -38710 7035 -38675 7070
rect -38665 7035 -38630 7070
rect -38620 7035 -38585 7070
rect -38575 7035 -38540 7070
rect -38530 7035 -38495 7070
rect -38485 7035 -38450 7070
rect -38440 7035 -38405 7070
rect -38395 7035 -38360 7070
rect -38350 7035 -38315 7070
rect -38305 7035 -38270 7070
rect -38260 7035 -38225 7070
rect -38215 7035 -38180 7070
rect -38170 7035 -38135 7070
rect -38125 7035 -38090 7070
rect -38080 7035 -38045 7070
rect -38035 7035 -38000 7070
rect -37990 7035 -37955 7070
rect -37945 7035 -37910 7070
rect -37900 7035 -37865 7070
rect -37855 7035 -37820 7070
rect -37810 7035 -37775 7070
rect -37765 7035 -37730 7070
rect -37720 7035 -37685 7070
rect -37675 7035 -37640 7070
rect -37630 7035 -37595 7070
rect -37585 7035 -37550 7070
rect -37540 7035 -37505 7070
rect -37495 7035 -37460 7070
rect -37450 7035 -37415 7070
rect -37405 7035 -37370 7070
rect -37360 7035 -37325 7070
rect -37315 7035 -37280 7070
rect -37270 7035 -37235 7070
rect -37225 7035 -37190 7070
rect -38755 6990 -38720 7025
rect -38710 6990 -38675 7025
rect -38665 6990 -38630 7025
rect -38620 6990 -38585 7025
rect -38575 6990 -38540 7025
rect -38530 6990 -38495 7025
rect -38485 6990 -38450 7025
rect -38440 6990 -38405 7025
rect -38395 6990 -38360 7025
rect -38350 6990 -38315 7025
rect -38305 6990 -38270 7025
rect -38260 6990 -38225 7025
rect -38215 6990 -38180 7025
rect -38170 6990 -38135 7025
rect -38125 6990 -38090 7025
rect -38080 6990 -38045 7025
rect -38035 6990 -38000 7025
rect -37990 6990 -37955 7025
rect -37945 6990 -37910 7025
rect -37900 6990 -37865 7025
rect -37855 6990 -37820 7025
rect -37810 6990 -37775 7025
rect -37765 6990 -37730 7025
rect -37720 6990 -37685 7025
rect -37675 6990 -37640 7025
rect -37630 6990 -37595 7025
rect -37585 6990 -37550 7025
rect -37540 6990 -37505 7025
rect -37495 6990 -37460 7025
rect -37450 6990 -37415 7025
rect -37405 6990 -37370 7025
rect -37360 6990 -37325 7025
rect -37315 6990 -37280 7025
rect -37270 6990 -37235 7025
rect -37225 6990 -37190 7025
rect -38755 6945 -38720 6980
rect -38710 6945 -38675 6980
rect -38665 6945 -38630 6980
rect -38620 6945 -38585 6980
rect -38575 6945 -38540 6980
rect -38530 6945 -38495 6980
rect -38485 6945 -38450 6980
rect -38440 6945 -38405 6980
rect -38395 6945 -38360 6980
rect -38350 6945 -38315 6980
rect -38305 6945 -38270 6980
rect -38260 6945 -38225 6980
rect -38215 6945 -38180 6980
rect -38170 6945 -38135 6980
rect -38125 6945 -38090 6980
rect -38080 6945 -38045 6980
rect -38035 6945 -38000 6980
rect -37990 6945 -37955 6980
rect -37945 6945 -37910 6980
rect -37900 6945 -37865 6980
rect -37855 6945 -37820 6980
rect -37810 6945 -37775 6980
rect -37765 6945 -37730 6980
rect -37720 6945 -37685 6980
rect -37675 6945 -37640 6980
rect -37630 6945 -37595 6980
rect -37585 6945 -37550 6980
rect -37540 6945 -37505 6980
rect -37495 6945 -37460 6980
rect -37450 6945 -37415 6980
rect -37405 6945 -37370 6980
rect -37360 6945 -37325 6980
rect -37315 6945 -37280 6980
rect -37270 6945 -37235 6980
rect -37225 6945 -37190 6980
rect -38755 6900 -38720 6935
rect -38710 6900 -38675 6935
rect -38665 6900 -38630 6935
rect -38620 6900 -38585 6935
rect -38575 6900 -38540 6935
rect -38530 6900 -38495 6935
rect -38485 6900 -38450 6935
rect -38440 6900 -38405 6935
rect -38395 6900 -38360 6935
rect -38350 6900 -38315 6935
rect -38305 6900 -38270 6935
rect -38260 6900 -38225 6935
rect -38215 6900 -38180 6935
rect -38170 6900 -38135 6935
rect -38125 6900 -38090 6935
rect -38080 6900 -38045 6935
rect -38035 6900 -38000 6935
rect -37990 6900 -37955 6935
rect -37945 6900 -37910 6935
rect -37900 6900 -37865 6935
rect -37855 6900 -37820 6935
rect -37810 6900 -37775 6935
rect -37765 6900 -37730 6935
rect -37720 6900 -37685 6935
rect -37675 6900 -37640 6935
rect -37630 6900 -37595 6935
rect -37585 6900 -37550 6935
rect -37540 6900 -37505 6935
rect -37495 6900 -37460 6935
rect -37450 6900 -37415 6935
rect -37405 6900 -37370 6935
rect -37360 6900 -37325 6935
rect -37315 6900 -37280 6935
rect -37270 6900 -37235 6935
rect -37225 6900 -37190 6935
rect -38755 6855 -38720 6890
rect -38710 6855 -38675 6890
rect -38665 6855 -38630 6890
rect -38620 6855 -38585 6890
rect -38575 6855 -38540 6890
rect -38530 6855 -38495 6890
rect -38485 6855 -38450 6890
rect -38440 6855 -38405 6890
rect -38395 6855 -38360 6890
rect -38350 6855 -38315 6890
rect -38305 6855 -38270 6890
rect -38260 6855 -38225 6890
rect -38215 6855 -38180 6890
rect -38170 6855 -38135 6890
rect -38125 6855 -38090 6890
rect -38080 6855 -38045 6890
rect -38035 6855 -38000 6890
rect -37990 6855 -37955 6890
rect -37945 6855 -37910 6890
rect -37900 6855 -37865 6890
rect -37855 6855 -37820 6890
rect -37810 6855 -37775 6890
rect -37765 6855 -37730 6890
rect -37720 6855 -37685 6890
rect -37675 6855 -37640 6890
rect -37630 6855 -37595 6890
rect -37585 6855 -37550 6890
rect -37540 6855 -37505 6890
rect -37495 6855 -37460 6890
rect -37450 6855 -37415 6890
rect -37405 6855 -37370 6890
rect -37360 6855 -37325 6890
rect -37315 6855 -37280 6890
rect -37270 6855 -37235 6890
rect -37225 6855 -37190 6890
rect -38755 6810 -38720 6845
rect -38710 6810 -38675 6845
rect -38665 6810 -38630 6845
rect -38620 6810 -38585 6845
rect -38575 6810 -38540 6845
rect -38530 6810 -38495 6845
rect -38485 6810 -38450 6845
rect -38440 6810 -38405 6845
rect -38395 6810 -38360 6845
rect -38350 6810 -38315 6845
rect -38305 6810 -38270 6845
rect -38260 6810 -38225 6845
rect -38215 6810 -38180 6845
rect -38170 6810 -38135 6845
rect -38125 6810 -38090 6845
rect -38080 6810 -38045 6845
rect -38035 6810 -38000 6845
rect -37990 6810 -37955 6845
rect -37945 6810 -37910 6845
rect -37900 6810 -37865 6845
rect -37855 6810 -37820 6845
rect -37810 6810 -37775 6845
rect -37765 6810 -37730 6845
rect -37720 6810 -37685 6845
rect -37675 6810 -37640 6845
rect -37630 6810 -37595 6845
rect -37585 6810 -37550 6845
rect -37540 6810 -37505 6845
rect -37495 6810 -37460 6845
rect -37450 6810 -37415 6845
rect -37405 6810 -37370 6845
rect -37360 6810 -37325 6845
rect -37315 6810 -37280 6845
rect -37270 6810 -37235 6845
rect -37225 6810 -37190 6845
rect -38755 6765 -38720 6800
rect -38710 6765 -38675 6800
rect -38665 6765 -38630 6800
rect -38620 6765 -38585 6800
rect -38575 6765 -38540 6800
rect -38530 6765 -38495 6800
rect -38485 6765 -38450 6800
rect -38440 6765 -38405 6800
rect -38395 6765 -38360 6800
rect -38350 6765 -38315 6800
rect -38305 6765 -38270 6800
rect -38260 6765 -38225 6800
rect -38215 6765 -38180 6800
rect -38170 6765 -38135 6800
rect -38125 6765 -38090 6800
rect -38080 6765 -38045 6800
rect -38035 6765 -38000 6800
rect -37990 6765 -37955 6800
rect -37945 6765 -37910 6800
rect -37900 6765 -37865 6800
rect -37855 6765 -37820 6800
rect -37810 6765 -37775 6800
rect -37765 6765 -37730 6800
rect -37720 6765 -37685 6800
rect -37675 6765 -37640 6800
rect -37630 6765 -37595 6800
rect -37585 6765 -37550 6800
rect -37540 6765 -37505 6800
rect -37495 6765 -37460 6800
rect -37450 6765 -37415 6800
rect -37405 6765 -37370 6800
rect -37360 6765 -37325 6800
rect -37315 6765 -37280 6800
rect -37270 6765 -37235 6800
rect -37225 6765 -37190 6800
rect -38755 6720 -38720 6755
rect -38710 6720 -38675 6755
rect -38665 6720 -38630 6755
rect -38620 6720 -38585 6755
rect -38575 6720 -38540 6755
rect -38530 6720 -38495 6755
rect -38485 6720 -38450 6755
rect -38440 6720 -38405 6755
rect -38395 6720 -38360 6755
rect -38350 6720 -38315 6755
rect -38305 6720 -38270 6755
rect -38260 6720 -38225 6755
rect -38215 6720 -38180 6755
rect -38170 6720 -38135 6755
rect -38125 6720 -38090 6755
rect -38080 6720 -38045 6755
rect -38035 6720 -38000 6755
rect -37990 6720 -37955 6755
rect -37945 6720 -37910 6755
rect -37900 6720 -37865 6755
rect -37855 6720 -37820 6755
rect -37810 6720 -37775 6755
rect -37765 6720 -37730 6755
rect -37720 6720 -37685 6755
rect -37675 6720 -37640 6755
rect -37630 6720 -37595 6755
rect -37585 6720 -37550 6755
rect -37540 6720 -37505 6755
rect -37495 6720 -37460 6755
rect -37450 6720 -37415 6755
rect -37405 6720 -37370 6755
rect -37360 6720 -37325 6755
rect -37315 6720 -37280 6755
rect -37270 6720 -37235 6755
rect -37225 6720 -37190 6755
rect -38755 6675 -38720 6710
rect -38710 6675 -38675 6710
rect -38665 6675 -38630 6710
rect -38620 6675 -38585 6710
rect -38575 6675 -38540 6710
rect -38530 6675 -38495 6710
rect -38485 6675 -38450 6710
rect -38440 6675 -38405 6710
rect -38395 6675 -38360 6710
rect -38350 6675 -38315 6710
rect -38305 6675 -38270 6710
rect -38260 6675 -38225 6710
rect -38215 6675 -38180 6710
rect -38170 6675 -38135 6710
rect -38125 6675 -38090 6710
rect -38080 6675 -38045 6710
rect -38035 6675 -38000 6710
rect -37990 6675 -37955 6710
rect -37945 6675 -37910 6710
rect -37900 6675 -37865 6710
rect -37855 6675 -37820 6710
rect -37810 6675 -37775 6710
rect -37765 6675 -37730 6710
rect -37720 6675 -37685 6710
rect -37675 6675 -37640 6710
rect -37630 6675 -37595 6710
rect -37585 6675 -37550 6710
rect -37540 6675 -37505 6710
rect -37495 6675 -37460 6710
rect -37450 6675 -37415 6710
rect -37405 6675 -37370 6710
rect -37360 6675 -37325 6710
rect -37315 6675 -37280 6710
rect -37270 6675 -37235 6710
rect -37225 6675 -37190 6710
rect -38755 6630 -38720 6665
rect -38710 6630 -38675 6665
rect -38665 6630 -38630 6665
rect -38620 6630 -38585 6665
rect -38575 6630 -38540 6665
rect -38530 6630 -38495 6665
rect -38485 6630 -38450 6665
rect -38440 6630 -38405 6665
rect -38395 6630 -38360 6665
rect -38350 6630 -38315 6665
rect -38305 6630 -38270 6665
rect -38260 6630 -38225 6665
rect -38215 6630 -38180 6665
rect -38170 6630 -38135 6665
rect -38125 6630 -38090 6665
rect -38080 6630 -38045 6665
rect -38035 6630 -38000 6665
rect -37990 6630 -37955 6665
rect -37945 6630 -37910 6665
rect -37900 6630 -37865 6665
rect -37855 6630 -37820 6665
rect -37810 6630 -37775 6665
rect -37765 6630 -37730 6665
rect -37720 6630 -37685 6665
rect -37675 6630 -37640 6665
rect -37630 6630 -37595 6665
rect -37585 6630 -37550 6665
rect -37540 6630 -37505 6665
rect -37495 6630 -37460 6665
rect -37450 6630 -37415 6665
rect -37405 6630 -37370 6665
rect -37360 6630 -37325 6665
rect -37315 6630 -37280 6665
rect -37270 6630 -37235 6665
rect -37225 6630 -37190 6665
rect -38755 6585 -38720 6620
rect -38710 6585 -38675 6620
rect -38665 6585 -38630 6620
rect -38620 6585 -38585 6620
rect -38575 6585 -38540 6620
rect -38530 6585 -38495 6620
rect -38485 6585 -38450 6620
rect -38440 6585 -38405 6620
rect -38395 6585 -38360 6620
rect -38350 6585 -38315 6620
rect -38305 6585 -38270 6620
rect -38260 6585 -38225 6620
rect -38215 6585 -38180 6620
rect -38170 6585 -38135 6620
rect -38125 6585 -38090 6620
rect -38080 6585 -38045 6620
rect -38035 6585 -38000 6620
rect -37990 6585 -37955 6620
rect -37945 6585 -37910 6620
rect -37900 6585 -37865 6620
rect -37855 6585 -37820 6620
rect -37810 6585 -37775 6620
rect -37765 6585 -37730 6620
rect -37720 6585 -37685 6620
rect -37675 6585 -37640 6620
rect -37630 6585 -37595 6620
rect -37585 6585 -37550 6620
rect -37540 6585 -37505 6620
rect -37495 6585 -37460 6620
rect -37450 6585 -37415 6620
rect -37405 6585 -37370 6620
rect -37360 6585 -37325 6620
rect -37315 6585 -37280 6620
rect -37270 6585 -37235 6620
rect -37225 6585 -37190 6620
rect -38755 6540 -38720 6575
rect -38710 6540 -38675 6575
rect -38665 6540 -38630 6575
rect -38620 6540 -38585 6575
rect -38575 6540 -38540 6575
rect -38530 6540 -38495 6575
rect -38485 6540 -38450 6575
rect -38440 6540 -38405 6575
rect -38395 6540 -38360 6575
rect -38350 6540 -38315 6575
rect -38305 6540 -38270 6575
rect -38260 6540 -38225 6575
rect -38215 6540 -38180 6575
rect -38170 6540 -38135 6575
rect -38125 6540 -38090 6575
rect -38080 6540 -38045 6575
rect -38035 6540 -38000 6575
rect -37990 6540 -37955 6575
rect -37945 6540 -37910 6575
rect -37900 6540 -37865 6575
rect -37855 6540 -37820 6575
rect -37810 6540 -37775 6575
rect -37765 6540 -37730 6575
rect -37720 6540 -37685 6575
rect -37675 6540 -37640 6575
rect -37630 6540 -37595 6575
rect -37585 6540 -37550 6575
rect -37540 6540 -37505 6575
rect -37495 6540 -37460 6575
rect -37450 6540 -37415 6575
rect -37405 6540 -37370 6575
rect -37360 6540 -37325 6575
rect -37315 6540 -37280 6575
rect -37270 6540 -37235 6575
rect -37225 6540 -37190 6575
rect -38755 6495 -38720 6530
rect -38710 6495 -38675 6530
rect -38665 6495 -38630 6530
rect -38620 6495 -38585 6530
rect -38575 6495 -38540 6530
rect -38530 6495 -38495 6530
rect -38485 6495 -38450 6530
rect -38440 6495 -38405 6530
rect -38395 6495 -38360 6530
rect -38350 6495 -38315 6530
rect -38305 6495 -38270 6530
rect -38260 6495 -38225 6530
rect -38215 6495 -38180 6530
rect -38170 6495 -38135 6530
rect -38125 6495 -38090 6530
rect -38080 6495 -38045 6530
rect -38035 6495 -38000 6530
rect -37990 6495 -37955 6530
rect -37945 6495 -37910 6530
rect -37900 6495 -37865 6530
rect -37855 6495 -37820 6530
rect -37810 6495 -37775 6530
rect -37765 6495 -37730 6530
rect -37720 6495 -37685 6530
rect -37675 6495 -37640 6530
rect -37630 6495 -37595 6530
rect -37585 6495 -37550 6530
rect -37540 6495 -37505 6530
rect -37495 6495 -37460 6530
rect -37450 6495 -37415 6530
rect -37405 6495 -37370 6530
rect -37360 6495 -37325 6530
rect -37315 6495 -37280 6530
rect -37270 6495 -37235 6530
rect -37225 6495 -37190 6530
rect -38755 6450 -38720 6485
rect -38710 6450 -38675 6485
rect -38665 6450 -38630 6485
rect -38620 6450 -38585 6485
rect -38575 6450 -38540 6485
rect -38530 6450 -38495 6485
rect -38485 6450 -38450 6485
rect -38440 6450 -38405 6485
rect -38395 6450 -38360 6485
rect -38350 6450 -38315 6485
rect -38305 6450 -38270 6485
rect -38260 6450 -38225 6485
rect -38215 6450 -38180 6485
rect -38170 6450 -38135 6485
rect -38125 6450 -38090 6485
rect -38080 6450 -38045 6485
rect -38035 6450 -38000 6485
rect -37990 6450 -37955 6485
rect -37945 6450 -37910 6485
rect -37900 6450 -37865 6485
rect -37855 6450 -37820 6485
rect -37810 6450 -37775 6485
rect -37765 6450 -37730 6485
rect -37720 6450 -37685 6485
rect -37675 6450 -37640 6485
rect -37630 6450 -37595 6485
rect -37585 6450 -37550 6485
rect -37540 6450 -37505 6485
rect -37495 6450 -37460 6485
rect -37450 6450 -37415 6485
rect -37405 6450 -37370 6485
rect -37360 6450 -37325 6485
rect -37315 6450 -37280 6485
rect -37270 6450 -37235 6485
rect -37225 6450 -37190 6485
rect 3175 7955 3215 7960
rect 3175 7925 3180 7955
rect 3180 7925 3210 7955
rect 3210 7925 3215 7955
rect 3175 7920 3215 7925
rect 3235 7955 3275 7960
rect 3235 7925 3240 7955
rect 3240 7925 3270 7955
rect 3270 7925 3275 7955
rect 3235 7920 3275 7925
rect 3175 7885 3215 7890
rect 3175 7855 3180 7885
rect 3180 7855 3210 7885
rect 3210 7855 3215 7885
rect 3175 7850 3215 7855
rect 3235 7885 3275 7890
rect 3235 7855 3240 7885
rect 3240 7855 3270 7885
rect 3270 7855 3275 7885
rect 3235 7850 3275 7855
rect 3175 7815 3215 7820
rect 3175 7785 3180 7815
rect 3180 7785 3210 7815
rect 3210 7785 3215 7815
rect 3175 7780 3215 7785
rect 3235 7815 3275 7820
rect 3235 7785 3240 7815
rect 3240 7785 3270 7815
rect 3270 7785 3275 7815
rect 3235 7780 3275 7785
rect 3175 7745 3215 7750
rect 3175 7715 3180 7745
rect 3180 7715 3210 7745
rect 3210 7715 3215 7745
rect 3175 7710 3215 7715
rect 3235 7745 3275 7750
rect 3235 7715 3240 7745
rect 3240 7715 3270 7745
rect 3270 7715 3275 7745
rect 3235 7710 3275 7715
rect 3175 7680 3215 7685
rect 3175 7650 3180 7680
rect 3180 7650 3210 7680
rect 3210 7650 3215 7680
rect 3175 7645 3215 7650
rect 3235 7680 3275 7685
rect 3235 7650 3240 7680
rect 3240 7650 3270 7680
rect 3270 7650 3275 7680
rect 3235 7645 3275 7650
rect 3175 7620 3215 7625
rect 3175 7590 3180 7620
rect 3180 7590 3210 7620
rect 3210 7590 3215 7620
rect 3175 7585 3215 7590
rect 3235 7620 3275 7625
rect 3235 7590 3240 7620
rect 3240 7590 3270 7620
rect 3270 7590 3275 7620
rect 3235 7585 3275 7590
rect 3175 7555 3215 7560
rect 3175 7525 3180 7555
rect 3180 7525 3210 7555
rect 3210 7525 3215 7555
rect 3175 7520 3215 7525
rect 3235 7555 3275 7560
rect 3235 7525 3240 7555
rect 3240 7525 3270 7555
rect 3270 7525 3275 7555
rect 3235 7520 3275 7525
rect 3175 7485 3215 7490
rect 3175 7455 3180 7485
rect 3180 7455 3210 7485
rect 3210 7455 3215 7485
rect 3175 7450 3215 7455
rect 3235 7485 3275 7490
rect 3235 7455 3240 7485
rect 3240 7455 3270 7485
rect 3270 7455 3275 7485
rect 3235 7450 3275 7455
rect 3175 7415 3215 7420
rect 3175 7385 3180 7415
rect 3180 7385 3210 7415
rect 3210 7385 3215 7415
rect 3175 7380 3215 7385
rect 3235 7415 3275 7420
rect 3235 7385 3240 7415
rect 3240 7385 3270 7415
rect 3270 7385 3275 7415
rect 3235 7380 3275 7385
rect 3175 7345 3215 7350
rect 3175 7315 3180 7345
rect 3180 7315 3210 7345
rect 3210 7315 3215 7345
rect 3175 7310 3215 7315
rect 3235 7345 3275 7350
rect 3235 7315 3240 7345
rect 3240 7315 3270 7345
rect 3270 7315 3275 7345
rect 3235 7310 3275 7315
rect 3175 7280 3215 7285
rect 3175 7250 3180 7280
rect 3180 7250 3210 7280
rect 3210 7250 3215 7280
rect 3175 7245 3215 7250
rect 3235 7280 3275 7285
rect 3235 7250 3240 7280
rect 3240 7250 3270 7280
rect 3270 7250 3275 7280
rect 3235 7245 3275 7250
rect 3175 7220 3215 7225
rect 3175 7190 3180 7220
rect 3180 7190 3210 7220
rect 3210 7190 3215 7220
rect 3175 7185 3215 7190
rect 3235 7220 3275 7225
rect 3235 7190 3240 7220
rect 3240 7190 3270 7220
rect 3270 7190 3275 7220
rect 3235 7185 3275 7190
rect 3175 7155 3215 7160
rect 3175 7125 3180 7155
rect 3180 7125 3210 7155
rect 3210 7125 3215 7155
rect 3175 7120 3215 7125
rect 3235 7155 3275 7160
rect 3235 7125 3240 7155
rect 3240 7125 3270 7155
rect 3270 7125 3275 7155
rect 3235 7120 3275 7125
rect 3175 7085 3215 7090
rect 3175 7055 3180 7085
rect 3180 7055 3210 7085
rect 3210 7055 3215 7085
rect 3175 7050 3215 7055
rect 3235 7085 3275 7090
rect 3235 7055 3240 7085
rect 3240 7055 3270 7085
rect 3270 7055 3275 7085
rect 3235 7050 3275 7055
rect 3175 7015 3215 7020
rect 3175 6985 3180 7015
rect 3180 6985 3210 7015
rect 3210 6985 3215 7015
rect 3175 6980 3215 6985
rect 3235 7015 3275 7020
rect 3235 6985 3240 7015
rect 3240 6985 3270 7015
rect 3270 6985 3275 7015
rect 3235 6980 3275 6985
rect 3175 6945 3215 6950
rect 3175 6915 3180 6945
rect 3180 6915 3210 6945
rect 3210 6915 3215 6945
rect 3175 6910 3215 6915
rect 3235 6945 3275 6950
rect 3235 6915 3240 6945
rect 3240 6915 3270 6945
rect 3270 6915 3275 6945
rect 3235 6910 3275 6915
rect 3175 6880 3215 6885
rect 3175 6850 3180 6880
rect 3180 6850 3210 6880
rect 3210 6850 3215 6880
rect 3175 6845 3215 6850
rect 3235 6880 3275 6885
rect 3235 6850 3240 6880
rect 3240 6850 3270 6880
rect 3270 6850 3275 6880
rect 3235 6845 3275 6850
rect 3175 6820 3215 6825
rect 3175 6790 3180 6820
rect 3180 6790 3210 6820
rect 3210 6790 3215 6820
rect 3175 6785 3215 6790
rect 3235 6820 3275 6825
rect 3235 6790 3240 6820
rect 3240 6790 3270 6820
rect 3270 6790 3275 6820
rect 3235 6785 3275 6790
rect 3175 6755 3215 6760
rect 3175 6725 3180 6755
rect 3180 6725 3210 6755
rect 3210 6725 3215 6755
rect 3175 6720 3215 6725
rect 3235 6755 3275 6760
rect 3235 6725 3240 6755
rect 3240 6725 3270 6755
rect 3270 6725 3275 6755
rect 3235 6720 3275 6725
rect 3175 6685 3215 6690
rect 3175 6655 3180 6685
rect 3180 6655 3210 6685
rect 3210 6655 3215 6685
rect 3175 6650 3215 6655
rect 3235 6685 3275 6690
rect 3235 6655 3240 6685
rect 3240 6655 3270 6685
rect 3270 6655 3275 6685
rect 3235 6650 3275 6655
rect 3175 6615 3215 6620
rect 3175 6585 3180 6615
rect 3180 6585 3210 6615
rect 3210 6585 3215 6615
rect 3175 6580 3215 6585
rect 3235 6615 3275 6620
rect 3235 6585 3240 6615
rect 3240 6585 3270 6615
rect 3270 6585 3275 6615
rect 3235 6580 3275 6585
rect 3175 6545 3215 6550
rect 3175 6515 3180 6545
rect 3180 6515 3210 6545
rect 3210 6515 3215 6545
rect 3175 6510 3215 6515
rect 3235 6545 3275 6550
rect 3235 6515 3240 6545
rect 3240 6515 3270 6545
rect 3270 6515 3275 6545
rect 3235 6510 3275 6515
rect 3175 6480 3215 6485
rect 3175 6450 3180 6480
rect 3180 6450 3210 6480
rect 3210 6450 3215 6480
rect 3175 6445 3215 6450
rect 3235 6480 3275 6485
rect 3235 6450 3240 6480
rect 3240 6450 3270 6480
rect 3270 6450 3275 6480
rect 3235 6445 3275 6450
rect 3345 7955 3385 7960
rect 3345 7925 3350 7955
rect 3350 7925 3380 7955
rect 3380 7925 3385 7955
rect 3345 7920 3385 7925
rect 3345 7885 3385 7890
rect 3345 7855 3350 7885
rect 3350 7855 3380 7885
rect 3380 7855 3385 7885
rect 3345 7850 3385 7855
rect 3345 7815 3385 7820
rect 3345 7785 3350 7815
rect 3350 7785 3380 7815
rect 3380 7785 3385 7815
rect 3345 7780 3385 7785
rect 3345 7745 3385 7750
rect 3345 7715 3350 7745
rect 3350 7715 3380 7745
rect 3380 7715 3385 7745
rect 3345 7710 3385 7715
rect 3345 7680 3385 7685
rect 3345 7650 3350 7680
rect 3350 7650 3380 7680
rect 3380 7650 3385 7680
rect 3345 7645 3385 7650
rect 3345 7620 3385 7625
rect 3345 7590 3350 7620
rect 3350 7590 3380 7620
rect 3380 7590 3385 7620
rect 3345 7585 3385 7590
rect 3345 7555 3385 7560
rect 3345 7525 3350 7555
rect 3350 7525 3380 7555
rect 3380 7525 3385 7555
rect 3345 7520 3385 7525
rect 3345 7485 3385 7490
rect 3345 7455 3350 7485
rect 3350 7455 3380 7485
rect 3380 7455 3385 7485
rect 3345 7450 3385 7455
rect 3345 7415 3385 7420
rect 3345 7385 3350 7415
rect 3350 7385 3380 7415
rect 3380 7385 3385 7415
rect 3345 7380 3385 7385
rect 3345 7345 3385 7350
rect 3345 7315 3350 7345
rect 3350 7315 3380 7345
rect 3380 7315 3385 7345
rect 3345 7310 3385 7315
rect 3345 7280 3385 7285
rect 3345 7250 3350 7280
rect 3350 7250 3380 7280
rect 3380 7250 3385 7280
rect 3345 7245 3385 7250
rect 3345 7220 3385 7225
rect 3345 7190 3350 7220
rect 3350 7190 3380 7220
rect 3380 7190 3385 7220
rect 3345 7185 3385 7190
rect 3345 7155 3385 7160
rect 3345 7125 3350 7155
rect 3350 7125 3380 7155
rect 3380 7125 3385 7155
rect 3345 7120 3385 7125
rect 3345 7085 3385 7090
rect 3345 7055 3350 7085
rect 3350 7055 3380 7085
rect 3380 7055 3385 7085
rect 3345 7050 3385 7055
rect 3345 7015 3385 7020
rect 3345 6985 3350 7015
rect 3350 6985 3380 7015
rect 3380 6985 3385 7015
rect 3345 6980 3385 6985
rect 3345 6945 3385 6950
rect 3345 6915 3350 6945
rect 3350 6915 3380 6945
rect 3380 6915 3385 6945
rect 3345 6910 3385 6915
rect 3345 6880 3385 6885
rect 3345 6850 3350 6880
rect 3350 6850 3380 6880
rect 3380 6850 3385 6880
rect 3345 6845 3385 6850
rect 3345 6820 3385 6825
rect 3345 6790 3350 6820
rect 3350 6790 3380 6820
rect 3380 6790 3385 6820
rect 3345 6785 3385 6790
rect 3345 6755 3385 6760
rect 3345 6725 3350 6755
rect 3350 6725 3380 6755
rect 3380 6725 3385 6755
rect 3345 6720 3385 6725
rect 3345 6685 3385 6690
rect 3345 6655 3350 6685
rect 3350 6655 3380 6685
rect 3380 6655 3385 6685
rect 3345 6650 3385 6655
rect 3345 6615 3385 6620
rect 3345 6585 3350 6615
rect 3350 6585 3380 6615
rect 3380 6585 3385 6615
rect 3345 6580 3385 6585
rect 3345 6545 3385 6550
rect 3345 6515 3350 6545
rect 3350 6515 3380 6545
rect 3380 6515 3385 6545
rect 3345 6510 3385 6515
rect 3345 6480 3385 6485
rect 3345 6450 3350 6480
rect 3350 6450 3380 6480
rect 3380 6450 3385 6480
rect 3345 6445 3385 6450
rect 31305 7950 31340 7985
rect 31350 7950 31385 7985
rect 31395 7950 31430 7985
rect 31440 7950 31475 7985
rect 31485 7950 31520 7985
rect 31530 7950 31565 7985
rect 31575 7950 31610 7985
rect 31620 7950 31655 7985
rect 31665 7950 31700 7985
rect 31710 7950 31745 7985
rect 31755 7950 31790 7985
rect 31800 7950 31835 7985
rect 31845 7950 31880 7985
rect 31890 7950 31925 7985
rect 31935 7950 31970 7985
rect 31980 7950 32015 7985
rect 32025 7950 32060 7985
rect 32070 7950 32105 7985
rect 32115 7950 32150 7985
rect 32160 7950 32195 7985
rect 32205 7950 32240 7985
rect 32250 7950 32285 7985
rect 32295 7950 32330 7985
rect 32340 7950 32375 7985
rect 32385 7950 32420 7985
rect 32430 7950 32465 7985
rect 32475 7950 32510 7985
rect 32520 7950 32555 7985
rect 32565 7950 32600 7985
rect 32610 7950 32645 7985
rect 32655 7950 32690 7985
rect 32700 7950 32735 7985
rect 32745 7950 32780 7985
rect 32790 7950 32825 7985
rect 32835 7950 32870 7985
rect 31305 7905 31340 7940
rect 31350 7905 31385 7940
rect 31395 7905 31430 7940
rect 31440 7905 31475 7940
rect 31485 7905 31520 7940
rect 31530 7905 31565 7940
rect 31575 7905 31610 7940
rect 31620 7905 31655 7940
rect 31665 7905 31700 7940
rect 31710 7905 31745 7940
rect 31755 7905 31790 7940
rect 31800 7905 31835 7940
rect 31845 7905 31880 7940
rect 31890 7905 31925 7940
rect 31935 7905 31970 7940
rect 31980 7905 32015 7940
rect 32025 7905 32060 7940
rect 32070 7905 32105 7940
rect 32115 7905 32150 7940
rect 32160 7905 32195 7940
rect 32205 7905 32240 7940
rect 32250 7905 32285 7940
rect 32295 7905 32330 7940
rect 32340 7905 32375 7940
rect 32385 7905 32420 7940
rect 32430 7905 32465 7940
rect 32475 7905 32510 7940
rect 32520 7905 32555 7940
rect 32565 7905 32600 7940
rect 32610 7905 32645 7940
rect 32655 7905 32690 7940
rect 32700 7905 32735 7940
rect 32745 7905 32780 7940
rect 32790 7905 32825 7940
rect 32835 7905 32870 7940
rect 31305 7860 31340 7895
rect 31350 7860 31385 7895
rect 31395 7860 31430 7895
rect 31440 7860 31475 7895
rect 31485 7860 31520 7895
rect 31530 7860 31565 7895
rect 31575 7860 31610 7895
rect 31620 7860 31655 7895
rect 31665 7860 31700 7895
rect 31710 7860 31745 7895
rect 31755 7860 31790 7895
rect 31800 7860 31835 7895
rect 31845 7860 31880 7895
rect 31890 7860 31925 7895
rect 31935 7860 31970 7895
rect 31980 7860 32015 7895
rect 32025 7860 32060 7895
rect 32070 7860 32105 7895
rect 32115 7860 32150 7895
rect 32160 7860 32195 7895
rect 32205 7860 32240 7895
rect 32250 7860 32285 7895
rect 32295 7860 32330 7895
rect 32340 7860 32375 7895
rect 32385 7860 32420 7895
rect 32430 7860 32465 7895
rect 32475 7860 32510 7895
rect 32520 7860 32555 7895
rect 32565 7860 32600 7895
rect 32610 7860 32645 7895
rect 32655 7860 32690 7895
rect 32700 7860 32735 7895
rect 32745 7860 32780 7895
rect 32790 7860 32825 7895
rect 32835 7860 32870 7895
rect 31305 7815 31340 7850
rect 31350 7815 31385 7850
rect 31395 7815 31430 7850
rect 31440 7815 31475 7850
rect 31485 7815 31520 7850
rect 31530 7815 31565 7850
rect 31575 7815 31610 7850
rect 31620 7815 31655 7850
rect 31665 7815 31700 7850
rect 31710 7815 31745 7850
rect 31755 7815 31790 7850
rect 31800 7815 31835 7850
rect 31845 7815 31880 7850
rect 31890 7815 31925 7850
rect 31935 7815 31970 7850
rect 31980 7815 32015 7850
rect 32025 7815 32060 7850
rect 32070 7815 32105 7850
rect 32115 7815 32150 7850
rect 32160 7815 32195 7850
rect 32205 7815 32240 7850
rect 32250 7815 32285 7850
rect 32295 7815 32330 7850
rect 32340 7815 32375 7850
rect 32385 7815 32420 7850
rect 32430 7815 32465 7850
rect 32475 7815 32510 7850
rect 32520 7815 32555 7850
rect 32565 7815 32600 7850
rect 32610 7815 32645 7850
rect 32655 7815 32690 7850
rect 32700 7815 32735 7850
rect 32745 7815 32780 7850
rect 32790 7815 32825 7850
rect 32835 7815 32870 7850
rect 31305 7770 31340 7805
rect 31350 7770 31385 7805
rect 31395 7770 31430 7805
rect 31440 7770 31475 7805
rect 31485 7770 31520 7805
rect 31530 7770 31565 7805
rect 31575 7770 31610 7805
rect 31620 7770 31655 7805
rect 31665 7770 31700 7805
rect 31710 7770 31745 7805
rect 31755 7770 31790 7805
rect 31800 7770 31835 7805
rect 31845 7770 31880 7805
rect 31890 7770 31925 7805
rect 31935 7770 31970 7805
rect 31980 7770 32015 7805
rect 32025 7770 32060 7805
rect 32070 7770 32105 7805
rect 32115 7770 32150 7805
rect 32160 7770 32195 7805
rect 32205 7770 32240 7805
rect 32250 7770 32285 7805
rect 32295 7770 32330 7805
rect 32340 7770 32375 7805
rect 32385 7770 32420 7805
rect 32430 7770 32465 7805
rect 32475 7770 32510 7805
rect 32520 7770 32555 7805
rect 32565 7770 32600 7805
rect 32610 7770 32645 7805
rect 32655 7770 32690 7805
rect 32700 7770 32735 7805
rect 32745 7770 32780 7805
rect 32790 7770 32825 7805
rect 32835 7770 32870 7805
rect 31305 7725 31340 7760
rect 31350 7725 31385 7760
rect 31395 7725 31430 7760
rect 31440 7725 31475 7760
rect 31485 7725 31520 7760
rect 31530 7725 31565 7760
rect 31575 7725 31610 7760
rect 31620 7725 31655 7760
rect 31665 7725 31700 7760
rect 31710 7725 31745 7760
rect 31755 7725 31790 7760
rect 31800 7725 31835 7760
rect 31845 7725 31880 7760
rect 31890 7725 31925 7760
rect 31935 7725 31970 7760
rect 31980 7725 32015 7760
rect 32025 7725 32060 7760
rect 32070 7725 32105 7760
rect 32115 7725 32150 7760
rect 32160 7725 32195 7760
rect 32205 7725 32240 7760
rect 32250 7725 32285 7760
rect 32295 7725 32330 7760
rect 32340 7725 32375 7760
rect 32385 7725 32420 7760
rect 32430 7725 32465 7760
rect 32475 7725 32510 7760
rect 32520 7725 32555 7760
rect 32565 7725 32600 7760
rect 32610 7725 32645 7760
rect 32655 7725 32690 7760
rect 32700 7725 32735 7760
rect 32745 7725 32780 7760
rect 32790 7725 32825 7760
rect 32835 7725 32870 7760
rect 31305 7680 31340 7715
rect 31350 7680 31385 7715
rect 31395 7680 31430 7715
rect 31440 7680 31475 7715
rect 31485 7680 31520 7715
rect 31530 7680 31565 7715
rect 31575 7680 31610 7715
rect 31620 7680 31655 7715
rect 31665 7680 31700 7715
rect 31710 7680 31745 7715
rect 31755 7680 31790 7715
rect 31800 7680 31835 7715
rect 31845 7680 31880 7715
rect 31890 7680 31925 7715
rect 31935 7680 31970 7715
rect 31980 7680 32015 7715
rect 32025 7680 32060 7715
rect 32070 7680 32105 7715
rect 32115 7680 32150 7715
rect 32160 7680 32195 7715
rect 32205 7680 32240 7715
rect 32250 7680 32285 7715
rect 32295 7680 32330 7715
rect 32340 7680 32375 7715
rect 32385 7680 32420 7715
rect 32430 7680 32465 7715
rect 32475 7680 32510 7715
rect 32520 7680 32555 7715
rect 32565 7680 32600 7715
rect 32610 7680 32645 7715
rect 32655 7680 32690 7715
rect 32700 7680 32735 7715
rect 32745 7680 32780 7715
rect 32790 7680 32825 7715
rect 32835 7680 32870 7715
rect 31305 7635 31340 7670
rect 31350 7635 31385 7670
rect 31395 7635 31430 7670
rect 31440 7635 31475 7670
rect 31485 7635 31520 7670
rect 31530 7635 31565 7670
rect 31575 7635 31610 7670
rect 31620 7635 31655 7670
rect 31665 7635 31700 7670
rect 31710 7635 31745 7670
rect 31755 7635 31790 7670
rect 31800 7635 31835 7670
rect 31845 7635 31880 7670
rect 31890 7635 31925 7670
rect 31935 7635 31970 7670
rect 31980 7635 32015 7670
rect 32025 7635 32060 7670
rect 32070 7635 32105 7670
rect 32115 7635 32150 7670
rect 32160 7635 32195 7670
rect 32205 7635 32240 7670
rect 32250 7635 32285 7670
rect 32295 7635 32330 7670
rect 32340 7635 32375 7670
rect 32385 7635 32420 7670
rect 32430 7635 32465 7670
rect 32475 7635 32510 7670
rect 32520 7635 32555 7670
rect 32565 7635 32600 7670
rect 32610 7635 32645 7670
rect 32655 7635 32690 7670
rect 32700 7635 32735 7670
rect 32745 7635 32780 7670
rect 32790 7635 32825 7670
rect 32835 7635 32870 7670
rect 31305 7590 31340 7625
rect 31350 7590 31385 7625
rect 31395 7590 31430 7625
rect 31440 7590 31475 7625
rect 31485 7590 31520 7625
rect 31530 7590 31565 7625
rect 31575 7590 31610 7625
rect 31620 7590 31655 7625
rect 31665 7590 31700 7625
rect 31710 7590 31745 7625
rect 31755 7590 31790 7625
rect 31800 7590 31835 7625
rect 31845 7590 31880 7625
rect 31890 7590 31925 7625
rect 31935 7590 31970 7625
rect 31980 7590 32015 7625
rect 32025 7590 32060 7625
rect 32070 7590 32105 7625
rect 32115 7590 32150 7625
rect 32160 7590 32195 7625
rect 32205 7590 32240 7625
rect 32250 7590 32285 7625
rect 32295 7590 32330 7625
rect 32340 7590 32375 7625
rect 32385 7590 32420 7625
rect 32430 7590 32465 7625
rect 32475 7590 32510 7625
rect 32520 7590 32555 7625
rect 32565 7590 32600 7625
rect 32610 7590 32645 7625
rect 32655 7590 32690 7625
rect 32700 7590 32735 7625
rect 32745 7590 32780 7625
rect 32790 7590 32825 7625
rect 32835 7590 32870 7625
rect 31305 7545 31340 7580
rect 31350 7545 31385 7580
rect 31395 7545 31430 7580
rect 31440 7545 31475 7580
rect 31485 7545 31520 7580
rect 31530 7545 31565 7580
rect 31575 7545 31610 7580
rect 31620 7545 31655 7580
rect 31665 7545 31700 7580
rect 31710 7545 31745 7580
rect 31755 7545 31790 7580
rect 31800 7545 31835 7580
rect 31845 7545 31880 7580
rect 31890 7545 31925 7580
rect 31935 7545 31970 7580
rect 31980 7545 32015 7580
rect 32025 7545 32060 7580
rect 32070 7545 32105 7580
rect 32115 7545 32150 7580
rect 32160 7545 32195 7580
rect 32205 7545 32240 7580
rect 32250 7545 32285 7580
rect 32295 7545 32330 7580
rect 32340 7545 32375 7580
rect 32385 7545 32420 7580
rect 32430 7545 32465 7580
rect 32475 7545 32510 7580
rect 32520 7545 32555 7580
rect 32565 7545 32600 7580
rect 32610 7545 32645 7580
rect 32655 7545 32690 7580
rect 32700 7545 32735 7580
rect 32745 7545 32780 7580
rect 32790 7545 32825 7580
rect 32835 7545 32870 7580
rect 31305 7500 31340 7535
rect 31350 7500 31385 7535
rect 31395 7500 31430 7535
rect 31440 7500 31475 7535
rect 31485 7500 31520 7535
rect 31530 7500 31565 7535
rect 31575 7500 31610 7535
rect 31620 7500 31655 7535
rect 31665 7500 31700 7535
rect 31710 7500 31745 7535
rect 31755 7500 31790 7535
rect 31800 7500 31835 7535
rect 31845 7500 31880 7535
rect 31890 7500 31925 7535
rect 31935 7500 31970 7535
rect 31980 7500 32015 7535
rect 32025 7500 32060 7535
rect 32070 7500 32105 7535
rect 32115 7500 32150 7535
rect 32160 7500 32195 7535
rect 32205 7500 32240 7535
rect 32250 7500 32285 7535
rect 32295 7500 32330 7535
rect 32340 7500 32375 7535
rect 32385 7500 32420 7535
rect 32430 7500 32465 7535
rect 32475 7500 32510 7535
rect 32520 7500 32555 7535
rect 32565 7500 32600 7535
rect 32610 7500 32645 7535
rect 32655 7500 32690 7535
rect 32700 7500 32735 7535
rect 32745 7500 32780 7535
rect 32790 7500 32825 7535
rect 32835 7500 32870 7535
rect 31305 7455 31340 7490
rect 31350 7455 31385 7490
rect 31395 7455 31430 7490
rect 31440 7455 31475 7490
rect 31485 7455 31520 7490
rect 31530 7455 31565 7490
rect 31575 7455 31610 7490
rect 31620 7455 31655 7490
rect 31665 7455 31700 7490
rect 31710 7455 31745 7490
rect 31755 7455 31790 7490
rect 31800 7455 31835 7490
rect 31845 7455 31880 7490
rect 31890 7455 31925 7490
rect 31935 7455 31970 7490
rect 31980 7455 32015 7490
rect 32025 7455 32060 7490
rect 32070 7455 32105 7490
rect 32115 7455 32150 7490
rect 32160 7455 32195 7490
rect 32205 7455 32240 7490
rect 32250 7455 32285 7490
rect 32295 7455 32330 7490
rect 32340 7455 32375 7490
rect 32385 7455 32420 7490
rect 32430 7455 32465 7490
rect 32475 7455 32510 7490
rect 32520 7455 32555 7490
rect 32565 7455 32600 7490
rect 32610 7455 32645 7490
rect 32655 7455 32690 7490
rect 32700 7455 32735 7490
rect 32745 7455 32780 7490
rect 32790 7455 32825 7490
rect 32835 7455 32870 7490
rect 31305 7410 31340 7445
rect 31350 7410 31385 7445
rect 31395 7410 31430 7445
rect 31440 7410 31475 7445
rect 31485 7410 31520 7445
rect 31530 7410 31565 7445
rect 31575 7410 31610 7445
rect 31620 7410 31655 7445
rect 31665 7410 31700 7445
rect 31710 7410 31745 7445
rect 31755 7410 31790 7445
rect 31800 7410 31835 7445
rect 31845 7410 31880 7445
rect 31890 7410 31925 7445
rect 31935 7410 31970 7445
rect 31980 7410 32015 7445
rect 32025 7410 32060 7445
rect 32070 7410 32105 7445
rect 32115 7410 32150 7445
rect 32160 7410 32195 7445
rect 32205 7410 32240 7445
rect 32250 7410 32285 7445
rect 32295 7410 32330 7445
rect 32340 7410 32375 7445
rect 32385 7410 32420 7445
rect 32430 7410 32465 7445
rect 32475 7410 32510 7445
rect 32520 7410 32555 7445
rect 32565 7410 32600 7445
rect 32610 7410 32645 7445
rect 32655 7410 32690 7445
rect 32700 7410 32735 7445
rect 32745 7410 32780 7445
rect 32790 7410 32825 7445
rect 32835 7410 32870 7445
rect 31305 7365 31340 7400
rect 31350 7365 31385 7400
rect 31395 7365 31430 7400
rect 31440 7365 31475 7400
rect 31485 7365 31520 7400
rect 31530 7365 31565 7400
rect 31575 7365 31610 7400
rect 31620 7365 31655 7400
rect 31665 7365 31700 7400
rect 31710 7365 31745 7400
rect 31755 7365 31790 7400
rect 31800 7365 31835 7400
rect 31845 7365 31880 7400
rect 31890 7365 31925 7400
rect 31935 7365 31970 7400
rect 31980 7365 32015 7400
rect 32025 7365 32060 7400
rect 32070 7365 32105 7400
rect 32115 7365 32150 7400
rect 32160 7365 32195 7400
rect 32205 7365 32240 7400
rect 32250 7365 32285 7400
rect 32295 7365 32330 7400
rect 32340 7365 32375 7400
rect 32385 7365 32420 7400
rect 32430 7365 32465 7400
rect 32475 7365 32510 7400
rect 32520 7365 32555 7400
rect 32565 7365 32600 7400
rect 32610 7365 32645 7400
rect 32655 7365 32690 7400
rect 32700 7365 32735 7400
rect 32745 7365 32780 7400
rect 32790 7365 32825 7400
rect 32835 7365 32870 7400
rect 31305 7320 31340 7355
rect 31350 7320 31385 7355
rect 31395 7320 31430 7355
rect 31440 7320 31475 7355
rect 31485 7320 31520 7355
rect 31530 7320 31565 7355
rect 31575 7320 31610 7355
rect 31620 7320 31655 7355
rect 31665 7320 31700 7355
rect 31710 7320 31745 7355
rect 31755 7320 31790 7355
rect 31800 7320 31835 7355
rect 31845 7320 31880 7355
rect 31890 7320 31925 7355
rect 31935 7320 31970 7355
rect 31980 7320 32015 7355
rect 32025 7320 32060 7355
rect 32070 7320 32105 7355
rect 32115 7320 32150 7355
rect 32160 7320 32195 7355
rect 32205 7320 32240 7355
rect 32250 7320 32285 7355
rect 32295 7320 32330 7355
rect 32340 7320 32375 7355
rect 32385 7320 32420 7355
rect 32430 7320 32465 7355
rect 32475 7320 32510 7355
rect 32520 7320 32555 7355
rect 32565 7320 32600 7355
rect 32610 7320 32645 7355
rect 32655 7320 32690 7355
rect 32700 7320 32735 7355
rect 32745 7320 32780 7355
rect 32790 7320 32825 7355
rect 32835 7320 32870 7355
rect 31305 7275 31340 7310
rect 31350 7275 31385 7310
rect 31395 7275 31430 7310
rect 31440 7275 31475 7310
rect 31485 7275 31520 7310
rect 31530 7275 31565 7310
rect 31575 7275 31610 7310
rect 31620 7275 31655 7310
rect 31665 7275 31700 7310
rect 31710 7275 31745 7310
rect 31755 7275 31790 7310
rect 31800 7275 31835 7310
rect 31845 7275 31880 7310
rect 31890 7275 31925 7310
rect 31935 7275 31970 7310
rect 31980 7275 32015 7310
rect 32025 7275 32060 7310
rect 32070 7275 32105 7310
rect 32115 7275 32150 7310
rect 32160 7275 32195 7310
rect 32205 7275 32240 7310
rect 32250 7275 32285 7310
rect 32295 7275 32330 7310
rect 32340 7275 32375 7310
rect 32385 7275 32420 7310
rect 32430 7275 32465 7310
rect 32475 7275 32510 7310
rect 32520 7275 32555 7310
rect 32565 7275 32600 7310
rect 32610 7275 32645 7310
rect 32655 7275 32690 7310
rect 32700 7275 32735 7310
rect 32745 7275 32780 7310
rect 32790 7275 32825 7310
rect 32835 7275 32870 7310
rect 31305 7230 31340 7265
rect 31350 7230 31385 7265
rect 31395 7230 31430 7265
rect 31440 7230 31475 7265
rect 31485 7230 31520 7265
rect 31530 7230 31565 7265
rect 31575 7230 31610 7265
rect 31620 7230 31655 7265
rect 31665 7230 31700 7265
rect 31710 7230 31745 7265
rect 31755 7230 31790 7265
rect 31800 7230 31835 7265
rect 31845 7230 31880 7265
rect 31890 7230 31925 7265
rect 31935 7230 31970 7265
rect 31980 7230 32015 7265
rect 32025 7230 32060 7265
rect 32070 7230 32105 7265
rect 32115 7230 32150 7265
rect 32160 7230 32195 7265
rect 32205 7230 32240 7265
rect 32250 7230 32285 7265
rect 32295 7230 32330 7265
rect 32340 7230 32375 7265
rect 32385 7230 32420 7265
rect 32430 7230 32465 7265
rect 32475 7230 32510 7265
rect 32520 7230 32555 7265
rect 32565 7230 32600 7265
rect 32610 7230 32645 7265
rect 32655 7230 32690 7265
rect 32700 7230 32735 7265
rect 32745 7230 32780 7265
rect 32790 7230 32825 7265
rect 32835 7230 32870 7265
rect 31305 7185 31340 7220
rect 31350 7185 31385 7220
rect 31395 7185 31430 7220
rect 31440 7185 31475 7220
rect 31485 7185 31520 7220
rect 31530 7185 31565 7220
rect 31575 7185 31610 7220
rect 31620 7185 31655 7220
rect 31665 7185 31700 7220
rect 31710 7185 31745 7220
rect 31755 7185 31790 7220
rect 31800 7185 31835 7220
rect 31845 7185 31880 7220
rect 31890 7185 31925 7220
rect 31935 7185 31970 7220
rect 31980 7185 32015 7220
rect 32025 7185 32060 7220
rect 32070 7185 32105 7220
rect 32115 7185 32150 7220
rect 32160 7185 32195 7220
rect 32205 7185 32240 7220
rect 32250 7185 32285 7220
rect 32295 7185 32330 7220
rect 32340 7185 32375 7220
rect 32385 7185 32420 7220
rect 32430 7185 32465 7220
rect 32475 7185 32510 7220
rect 32520 7185 32555 7220
rect 32565 7185 32600 7220
rect 32610 7185 32645 7220
rect 32655 7185 32690 7220
rect 32700 7185 32735 7220
rect 32745 7185 32780 7220
rect 32790 7185 32825 7220
rect 32835 7185 32870 7220
rect 31305 7140 31340 7175
rect 31350 7140 31385 7175
rect 31395 7140 31430 7175
rect 31440 7140 31475 7175
rect 31485 7140 31520 7175
rect 31530 7140 31565 7175
rect 31575 7140 31610 7175
rect 31620 7140 31655 7175
rect 31665 7140 31700 7175
rect 31710 7140 31745 7175
rect 31755 7140 31790 7175
rect 31800 7140 31835 7175
rect 31845 7140 31880 7175
rect 31890 7140 31925 7175
rect 31935 7140 31970 7175
rect 31980 7140 32015 7175
rect 32025 7140 32060 7175
rect 32070 7140 32105 7175
rect 32115 7140 32150 7175
rect 32160 7140 32195 7175
rect 32205 7140 32240 7175
rect 32250 7140 32285 7175
rect 32295 7140 32330 7175
rect 32340 7140 32375 7175
rect 32385 7140 32420 7175
rect 32430 7140 32465 7175
rect 32475 7140 32510 7175
rect 32520 7140 32555 7175
rect 32565 7140 32600 7175
rect 32610 7140 32645 7175
rect 32655 7140 32690 7175
rect 32700 7140 32735 7175
rect 32745 7140 32780 7175
rect 32790 7140 32825 7175
rect 32835 7140 32870 7175
rect 31305 7095 31340 7130
rect 31350 7095 31385 7130
rect 31395 7095 31430 7130
rect 31440 7095 31475 7130
rect 31485 7095 31520 7130
rect 31530 7095 31565 7130
rect 31575 7095 31610 7130
rect 31620 7095 31655 7130
rect 31665 7095 31700 7130
rect 31710 7095 31745 7130
rect 31755 7095 31790 7130
rect 31800 7095 31835 7130
rect 31845 7095 31880 7130
rect 31890 7095 31925 7130
rect 31935 7095 31970 7130
rect 31980 7095 32015 7130
rect 32025 7095 32060 7130
rect 32070 7095 32105 7130
rect 32115 7095 32150 7130
rect 32160 7095 32195 7130
rect 32205 7095 32240 7130
rect 32250 7095 32285 7130
rect 32295 7095 32330 7130
rect 32340 7095 32375 7130
rect 32385 7095 32420 7130
rect 32430 7095 32465 7130
rect 32475 7095 32510 7130
rect 32520 7095 32555 7130
rect 32565 7095 32600 7130
rect 32610 7095 32645 7130
rect 32655 7095 32690 7130
rect 32700 7095 32735 7130
rect 32745 7095 32780 7130
rect 32790 7095 32825 7130
rect 32835 7095 32870 7130
rect 31305 7050 31340 7085
rect 31350 7050 31385 7085
rect 31395 7050 31430 7085
rect 31440 7050 31475 7085
rect 31485 7050 31520 7085
rect 31530 7050 31565 7085
rect 31575 7050 31610 7085
rect 31620 7050 31655 7085
rect 31665 7050 31700 7085
rect 31710 7050 31745 7085
rect 31755 7050 31790 7085
rect 31800 7050 31835 7085
rect 31845 7050 31880 7085
rect 31890 7050 31925 7085
rect 31935 7050 31970 7085
rect 31980 7050 32015 7085
rect 32025 7050 32060 7085
rect 32070 7050 32105 7085
rect 32115 7050 32150 7085
rect 32160 7050 32195 7085
rect 32205 7050 32240 7085
rect 32250 7050 32285 7085
rect 32295 7050 32330 7085
rect 32340 7050 32375 7085
rect 32385 7050 32420 7085
rect 32430 7050 32465 7085
rect 32475 7050 32510 7085
rect 32520 7050 32555 7085
rect 32565 7050 32600 7085
rect 32610 7050 32645 7085
rect 32655 7050 32690 7085
rect 32700 7050 32735 7085
rect 32745 7050 32780 7085
rect 32790 7050 32825 7085
rect 32835 7050 32870 7085
rect 31305 7005 31340 7040
rect 31350 7005 31385 7040
rect 31395 7005 31430 7040
rect 31440 7005 31475 7040
rect 31485 7005 31520 7040
rect 31530 7005 31565 7040
rect 31575 7005 31610 7040
rect 31620 7005 31655 7040
rect 31665 7005 31700 7040
rect 31710 7005 31745 7040
rect 31755 7005 31790 7040
rect 31800 7005 31835 7040
rect 31845 7005 31880 7040
rect 31890 7005 31925 7040
rect 31935 7005 31970 7040
rect 31980 7005 32015 7040
rect 32025 7005 32060 7040
rect 32070 7005 32105 7040
rect 32115 7005 32150 7040
rect 32160 7005 32195 7040
rect 32205 7005 32240 7040
rect 32250 7005 32285 7040
rect 32295 7005 32330 7040
rect 32340 7005 32375 7040
rect 32385 7005 32420 7040
rect 32430 7005 32465 7040
rect 32475 7005 32510 7040
rect 32520 7005 32555 7040
rect 32565 7005 32600 7040
rect 32610 7005 32645 7040
rect 32655 7005 32690 7040
rect 32700 7005 32735 7040
rect 32745 7005 32780 7040
rect 32790 7005 32825 7040
rect 32835 7005 32870 7040
rect 31305 6960 31340 6995
rect 31350 6960 31385 6995
rect 31395 6960 31430 6995
rect 31440 6960 31475 6995
rect 31485 6960 31520 6995
rect 31530 6960 31565 6995
rect 31575 6960 31610 6995
rect 31620 6960 31655 6995
rect 31665 6960 31700 6995
rect 31710 6960 31745 6995
rect 31755 6960 31790 6995
rect 31800 6960 31835 6995
rect 31845 6960 31880 6995
rect 31890 6960 31925 6995
rect 31935 6960 31970 6995
rect 31980 6960 32015 6995
rect 32025 6960 32060 6995
rect 32070 6960 32105 6995
rect 32115 6960 32150 6995
rect 32160 6960 32195 6995
rect 32205 6960 32240 6995
rect 32250 6960 32285 6995
rect 32295 6960 32330 6995
rect 32340 6960 32375 6995
rect 32385 6960 32420 6995
rect 32430 6960 32465 6995
rect 32475 6960 32510 6995
rect 32520 6960 32555 6995
rect 32565 6960 32600 6995
rect 32610 6960 32645 6995
rect 32655 6960 32690 6995
rect 32700 6960 32735 6995
rect 32745 6960 32780 6995
rect 32790 6960 32825 6995
rect 32835 6960 32870 6995
rect 31305 6915 31340 6950
rect 31350 6915 31385 6950
rect 31395 6915 31430 6950
rect 31440 6915 31475 6950
rect 31485 6915 31520 6950
rect 31530 6915 31565 6950
rect 31575 6915 31610 6950
rect 31620 6915 31655 6950
rect 31665 6915 31700 6950
rect 31710 6915 31745 6950
rect 31755 6915 31790 6950
rect 31800 6915 31835 6950
rect 31845 6915 31880 6950
rect 31890 6915 31925 6950
rect 31935 6915 31970 6950
rect 31980 6915 32015 6950
rect 32025 6915 32060 6950
rect 32070 6915 32105 6950
rect 32115 6915 32150 6950
rect 32160 6915 32195 6950
rect 32205 6915 32240 6950
rect 32250 6915 32285 6950
rect 32295 6915 32330 6950
rect 32340 6915 32375 6950
rect 32385 6915 32420 6950
rect 32430 6915 32465 6950
rect 32475 6915 32510 6950
rect 32520 6915 32555 6950
rect 32565 6915 32600 6950
rect 32610 6915 32645 6950
rect 32655 6915 32690 6950
rect 32700 6915 32735 6950
rect 32745 6915 32780 6950
rect 32790 6915 32825 6950
rect 32835 6915 32870 6950
rect 31305 6870 31340 6905
rect 31350 6870 31385 6905
rect 31395 6870 31430 6905
rect 31440 6870 31475 6905
rect 31485 6870 31520 6905
rect 31530 6870 31565 6905
rect 31575 6870 31610 6905
rect 31620 6870 31655 6905
rect 31665 6870 31700 6905
rect 31710 6870 31745 6905
rect 31755 6870 31790 6905
rect 31800 6870 31835 6905
rect 31845 6870 31880 6905
rect 31890 6870 31925 6905
rect 31935 6870 31970 6905
rect 31980 6870 32015 6905
rect 32025 6870 32060 6905
rect 32070 6870 32105 6905
rect 32115 6870 32150 6905
rect 32160 6870 32195 6905
rect 32205 6870 32240 6905
rect 32250 6870 32285 6905
rect 32295 6870 32330 6905
rect 32340 6870 32375 6905
rect 32385 6870 32420 6905
rect 32430 6870 32465 6905
rect 32475 6870 32510 6905
rect 32520 6870 32555 6905
rect 32565 6870 32600 6905
rect 32610 6870 32645 6905
rect 32655 6870 32690 6905
rect 32700 6870 32735 6905
rect 32745 6870 32780 6905
rect 32790 6870 32825 6905
rect 32835 6870 32870 6905
rect 31305 6825 31340 6860
rect 31350 6825 31385 6860
rect 31395 6825 31430 6860
rect 31440 6825 31475 6860
rect 31485 6825 31520 6860
rect 31530 6825 31565 6860
rect 31575 6825 31610 6860
rect 31620 6825 31655 6860
rect 31665 6825 31700 6860
rect 31710 6825 31745 6860
rect 31755 6825 31790 6860
rect 31800 6825 31835 6860
rect 31845 6825 31880 6860
rect 31890 6825 31925 6860
rect 31935 6825 31970 6860
rect 31980 6825 32015 6860
rect 32025 6825 32060 6860
rect 32070 6825 32105 6860
rect 32115 6825 32150 6860
rect 32160 6825 32195 6860
rect 32205 6825 32240 6860
rect 32250 6825 32285 6860
rect 32295 6825 32330 6860
rect 32340 6825 32375 6860
rect 32385 6825 32420 6860
rect 32430 6825 32465 6860
rect 32475 6825 32510 6860
rect 32520 6825 32555 6860
rect 32565 6825 32600 6860
rect 32610 6825 32645 6860
rect 32655 6825 32690 6860
rect 32700 6825 32735 6860
rect 32745 6825 32780 6860
rect 32790 6825 32825 6860
rect 32835 6825 32870 6860
rect 31305 6780 31340 6815
rect 31350 6780 31385 6815
rect 31395 6780 31430 6815
rect 31440 6780 31475 6815
rect 31485 6780 31520 6815
rect 31530 6780 31565 6815
rect 31575 6780 31610 6815
rect 31620 6780 31655 6815
rect 31665 6780 31700 6815
rect 31710 6780 31745 6815
rect 31755 6780 31790 6815
rect 31800 6780 31835 6815
rect 31845 6780 31880 6815
rect 31890 6780 31925 6815
rect 31935 6780 31970 6815
rect 31980 6780 32015 6815
rect 32025 6780 32060 6815
rect 32070 6780 32105 6815
rect 32115 6780 32150 6815
rect 32160 6780 32195 6815
rect 32205 6780 32240 6815
rect 32250 6780 32285 6815
rect 32295 6780 32330 6815
rect 32340 6780 32375 6815
rect 32385 6780 32420 6815
rect 32430 6780 32465 6815
rect 32475 6780 32510 6815
rect 32520 6780 32555 6815
rect 32565 6780 32600 6815
rect 32610 6780 32645 6815
rect 32655 6780 32690 6815
rect 32700 6780 32735 6815
rect 32745 6780 32780 6815
rect 32790 6780 32825 6815
rect 32835 6780 32870 6815
rect 31305 6735 31340 6770
rect 31350 6735 31385 6770
rect 31395 6735 31430 6770
rect 31440 6735 31475 6770
rect 31485 6735 31520 6770
rect 31530 6735 31565 6770
rect 31575 6735 31610 6770
rect 31620 6735 31655 6770
rect 31665 6735 31700 6770
rect 31710 6735 31745 6770
rect 31755 6735 31790 6770
rect 31800 6735 31835 6770
rect 31845 6735 31880 6770
rect 31890 6735 31925 6770
rect 31935 6735 31970 6770
rect 31980 6735 32015 6770
rect 32025 6735 32060 6770
rect 32070 6735 32105 6770
rect 32115 6735 32150 6770
rect 32160 6735 32195 6770
rect 32205 6735 32240 6770
rect 32250 6735 32285 6770
rect 32295 6735 32330 6770
rect 32340 6735 32375 6770
rect 32385 6735 32420 6770
rect 32430 6735 32465 6770
rect 32475 6735 32510 6770
rect 32520 6735 32555 6770
rect 32565 6735 32600 6770
rect 32610 6735 32645 6770
rect 32655 6735 32690 6770
rect 32700 6735 32735 6770
rect 32745 6735 32780 6770
rect 32790 6735 32825 6770
rect 32835 6735 32870 6770
rect 31305 6690 31340 6725
rect 31350 6690 31385 6725
rect 31395 6690 31430 6725
rect 31440 6690 31475 6725
rect 31485 6690 31520 6725
rect 31530 6690 31565 6725
rect 31575 6690 31610 6725
rect 31620 6690 31655 6725
rect 31665 6690 31700 6725
rect 31710 6690 31745 6725
rect 31755 6690 31790 6725
rect 31800 6690 31835 6725
rect 31845 6690 31880 6725
rect 31890 6690 31925 6725
rect 31935 6690 31970 6725
rect 31980 6690 32015 6725
rect 32025 6690 32060 6725
rect 32070 6690 32105 6725
rect 32115 6690 32150 6725
rect 32160 6690 32195 6725
rect 32205 6690 32240 6725
rect 32250 6690 32285 6725
rect 32295 6690 32330 6725
rect 32340 6690 32375 6725
rect 32385 6690 32420 6725
rect 32430 6690 32465 6725
rect 32475 6690 32510 6725
rect 32520 6690 32555 6725
rect 32565 6690 32600 6725
rect 32610 6690 32645 6725
rect 32655 6690 32690 6725
rect 32700 6690 32735 6725
rect 32745 6690 32780 6725
rect 32790 6690 32825 6725
rect 32835 6690 32870 6725
rect 31305 6645 31340 6680
rect 31350 6645 31385 6680
rect 31395 6645 31430 6680
rect 31440 6645 31475 6680
rect 31485 6645 31520 6680
rect 31530 6645 31565 6680
rect 31575 6645 31610 6680
rect 31620 6645 31655 6680
rect 31665 6645 31700 6680
rect 31710 6645 31745 6680
rect 31755 6645 31790 6680
rect 31800 6645 31835 6680
rect 31845 6645 31880 6680
rect 31890 6645 31925 6680
rect 31935 6645 31970 6680
rect 31980 6645 32015 6680
rect 32025 6645 32060 6680
rect 32070 6645 32105 6680
rect 32115 6645 32150 6680
rect 32160 6645 32195 6680
rect 32205 6645 32240 6680
rect 32250 6645 32285 6680
rect 32295 6645 32330 6680
rect 32340 6645 32375 6680
rect 32385 6645 32420 6680
rect 32430 6645 32465 6680
rect 32475 6645 32510 6680
rect 32520 6645 32555 6680
rect 32565 6645 32600 6680
rect 32610 6645 32645 6680
rect 32655 6645 32690 6680
rect 32700 6645 32735 6680
rect 32745 6645 32780 6680
rect 32790 6645 32825 6680
rect 32835 6645 32870 6680
rect 31305 6600 31340 6635
rect 31350 6600 31385 6635
rect 31395 6600 31430 6635
rect 31440 6600 31475 6635
rect 31485 6600 31520 6635
rect 31530 6600 31565 6635
rect 31575 6600 31610 6635
rect 31620 6600 31655 6635
rect 31665 6600 31700 6635
rect 31710 6600 31745 6635
rect 31755 6600 31790 6635
rect 31800 6600 31835 6635
rect 31845 6600 31880 6635
rect 31890 6600 31925 6635
rect 31935 6600 31970 6635
rect 31980 6600 32015 6635
rect 32025 6600 32060 6635
rect 32070 6600 32105 6635
rect 32115 6600 32150 6635
rect 32160 6600 32195 6635
rect 32205 6600 32240 6635
rect 32250 6600 32285 6635
rect 32295 6600 32330 6635
rect 32340 6600 32375 6635
rect 32385 6600 32420 6635
rect 32430 6600 32465 6635
rect 32475 6600 32510 6635
rect 32520 6600 32555 6635
rect 32565 6600 32600 6635
rect 32610 6600 32645 6635
rect 32655 6600 32690 6635
rect 32700 6600 32735 6635
rect 32745 6600 32780 6635
rect 32790 6600 32825 6635
rect 32835 6600 32870 6635
rect 31305 6555 31340 6590
rect 31350 6555 31385 6590
rect 31395 6555 31430 6590
rect 31440 6555 31475 6590
rect 31485 6555 31520 6590
rect 31530 6555 31565 6590
rect 31575 6555 31610 6590
rect 31620 6555 31655 6590
rect 31665 6555 31700 6590
rect 31710 6555 31745 6590
rect 31755 6555 31790 6590
rect 31800 6555 31835 6590
rect 31845 6555 31880 6590
rect 31890 6555 31925 6590
rect 31935 6555 31970 6590
rect 31980 6555 32015 6590
rect 32025 6555 32060 6590
rect 32070 6555 32105 6590
rect 32115 6555 32150 6590
rect 32160 6555 32195 6590
rect 32205 6555 32240 6590
rect 32250 6555 32285 6590
rect 32295 6555 32330 6590
rect 32340 6555 32375 6590
rect 32385 6555 32420 6590
rect 32430 6555 32465 6590
rect 32475 6555 32510 6590
rect 32520 6555 32555 6590
rect 32565 6555 32600 6590
rect 32610 6555 32645 6590
rect 32655 6555 32690 6590
rect 32700 6555 32735 6590
rect 32745 6555 32780 6590
rect 32790 6555 32825 6590
rect 32835 6555 32870 6590
rect 31305 6510 31340 6545
rect 31350 6510 31385 6545
rect 31395 6510 31430 6545
rect 31440 6510 31475 6545
rect 31485 6510 31520 6545
rect 31530 6510 31565 6545
rect 31575 6510 31610 6545
rect 31620 6510 31655 6545
rect 31665 6510 31700 6545
rect 31710 6510 31745 6545
rect 31755 6510 31790 6545
rect 31800 6510 31835 6545
rect 31845 6510 31880 6545
rect 31890 6510 31925 6545
rect 31935 6510 31970 6545
rect 31980 6510 32015 6545
rect 32025 6510 32060 6545
rect 32070 6510 32105 6545
rect 32115 6510 32150 6545
rect 32160 6510 32195 6545
rect 32205 6510 32240 6545
rect 32250 6510 32285 6545
rect 32295 6510 32330 6545
rect 32340 6510 32375 6545
rect 32385 6510 32420 6545
rect 32430 6510 32465 6545
rect 32475 6510 32510 6545
rect 32520 6510 32555 6545
rect 32565 6510 32600 6545
rect 32610 6510 32645 6545
rect 32655 6510 32690 6545
rect 32700 6510 32735 6545
rect 32745 6510 32780 6545
rect 32790 6510 32825 6545
rect 32835 6510 32870 6545
rect 31305 6465 31340 6500
rect 31350 6465 31385 6500
rect 31395 6465 31430 6500
rect 31440 6465 31475 6500
rect 31485 6465 31520 6500
rect 31530 6465 31565 6500
rect 31575 6465 31610 6500
rect 31620 6465 31655 6500
rect 31665 6465 31700 6500
rect 31710 6465 31745 6500
rect 31755 6465 31790 6500
rect 31800 6465 31835 6500
rect 31845 6465 31880 6500
rect 31890 6465 31925 6500
rect 31935 6465 31970 6500
rect 31980 6465 32015 6500
rect 32025 6465 32060 6500
rect 32070 6465 32105 6500
rect 32115 6465 32150 6500
rect 32160 6465 32195 6500
rect 32205 6465 32240 6500
rect 32250 6465 32285 6500
rect 32295 6465 32330 6500
rect 32340 6465 32375 6500
rect 32385 6465 32420 6500
rect 32430 6465 32465 6500
rect 32475 6465 32510 6500
rect 32520 6465 32555 6500
rect 32565 6465 32600 6500
rect 32610 6465 32645 6500
rect 32655 6465 32690 6500
rect 32700 6465 32735 6500
rect 32745 6465 32780 6500
rect 32790 6465 32825 6500
rect 32835 6465 32870 6500
rect -80 -1320 -40 -1315
rect -80 -1350 -75 -1320
rect -75 -1350 -45 -1320
rect -45 -1350 -40 -1320
rect -80 -1355 -40 -1350
rect -80 -1385 -40 -1380
rect -80 -1415 -75 -1385
rect -75 -1415 -45 -1385
rect -45 -1415 -40 -1385
rect -80 -1420 -40 -1415
rect -80 -1455 -40 -1450
rect -80 -1485 -75 -1455
rect -75 -1485 -45 -1455
rect -45 -1485 -40 -1455
rect -80 -1490 -40 -1485
rect -80 -1525 -40 -1520
rect -80 -1555 -75 -1525
rect -75 -1555 -45 -1525
rect -45 -1555 -40 -1525
rect -80 -1560 -40 -1555
rect -80 -1595 -40 -1590
rect -80 -1625 -75 -1595
rect -75 -1625 -45 -1595
rect -45 -1625 -40 -1595
rect -80 -1630 -40 -1625
rect -80 -1660 -40 -1655
rect -80 -1690 -75 -1660
rect -75 -1690 -45 -1660
rect -45 -1690 -40 -1660
rect -80 -1695 -40 -1690
rect -80 -1720 -40 -1715
rect -80 -1750 -75 -1720
rect -75 -1750 -45 -1720
rect -45 -1750 -40 -1720
rect -80 -1755 -40 -1750
rect -80 -1785 -40 -1780
rect -80 -1815 -75 -1785
rect -75 -1815 -45 -1785
rect -45 -1815 -40 -1785
rect -80 -1820 -40 -1815
rect -80 -1855 -40 -1850
rect -80 -1885 -75 -1855
rect -75 -1885 -45 -1855
rect -45 -1885 -40 -1855
rect -80 -1890 -40 -1885
rect -80 -1925 -40 -1920
rect -80 -1955 -75 -1925
rect -75 -1955 -45 -1925
rect -45 -1955 -40 -1925
rect -80 -1960 -40 -1955
rect -80 -1995 -40 -1990
rect -80 -2025 -75 -1995
rect -75 -2025 -45 -1995
rect -45 -2025 -40 -1995
rect -80 -2030 -40 -2025
rect -80 -2060 -40 -2055
rect -80 -2090 -75 -2060
rect -75 -2090 -45 -2060
rect -45 -2090 -40 -2060
rect -80 -2095 -40 -2090
rect -80 -2120 -40 -2115
rect -80 -2150 -75 -2120
rect -75 -2150 -45 -2120
rect -45 -2150 -40 -2120
rect -80 -2155 -40 -2150
rect -80 -2185 -40 -2180
rect -80 -2215 -75 -2185
rect -75 -2215 -45 -2185
rect -45 -2215 -40 -2185
rect -80 -2220 -40 -2215
rect -80 -2255 -40 -2250
rect -80 -2285 -75 -2255
rect -75 -2285 -45 -2255
rect -45 -2285 -40 -2255
rect -80 -2290 -40 -2285
rect -80 -2325 -40 -2320
rect -80 -2355 -75 -2325
rect -75 -2355 -45 -2325
rect -45 -2355 -40 -2325
rect -80 -2360 -40 -2355
rect -80 -2395 -40 -2390
rect -80 -2425 -75 -2395
rect -75 -2425 -45 -2395
rect -45 -2425 -40 -2395
rect -80 -2430 -40 -2425
rect -80 -2460 -40 -2455
rect -80 -2490 -75 -2460
rect -75 -2490 -45 -2460
rect -45 -2490 -40 -2460
rect -80 -2495 -40 -2490
rect -80 -2520 -40 -2515
rect -80 -2550 -75 -2520
rect -75 -2550 -45 -2520
rect -45 -2550 -40 -2520
rect -80 -2555 -40 -2550
rect -80 -2585 -40 -2580
rect -80 -2615 -75 -2585
rect -75 -2615 -45 -2585
rect -45 -2615 -40 -2585
rect -80 -2620 -40 -2615
rect -80 -2655 -40 -2650
rect -80 -2685 -75 -2655
rect -75 -2685 -45 -2655
rect -45 -2685 -40 -2655
rect -80 -2690 -40 -2685
rect -80 -2725 -40 -2720
rect -80 -2755 -75 -2725
rect -75 -2755 -45 -2725
rect -45 -2755 -40 -2725
rect -80 -2760 -40 -2755
rect -80 -2795 -40 -2790
rect -80 -2825 -75 -2795
rect -75 -2825 -45 -2795
rect -45 -2825 -40 -2795
rect -80 -2830 -40 -2825
rect -80 -2860 -40 -2855
rect -80 -2890 -75 -2860
rect -75 -2890 -45 -2860
rect -45 -2890 -40 -2860
rect -80 -2895 -40 -2890
rect 270 -1320 310 -1315
rect 270 -1350 275 -1320
rect 275 -1350 305 -1320
rect 305 -1350 310 -1320
rect 270 -1355 310 -1350
rect 270 -1385 310 -1380
rect 270 -1415 275 -1385
rect 275 -1415 305 -1385
rect 305 -1415 310 -1385
rect 270 -1420 310 -1415
rect 270 -1455 310 -1450
rect 270 -1485 275 -1455
rect 275 -1485 305 -1455
rect 305 -1485 310 -1455
rect 270 -1490 310 -1485
rect 270 -1525 310 -1520
rect 270 -1555 275 -1525
rect 275 -1555 305 -1525
rect 305 -1555 310 -1525
rect 270 -1560 310 -1555
rect 270 -1595 310 -1590
rect 270 -1625 275 -1595
rect 275 -1625 305 -1595
rect 305 -1625 310 -1595
rect 270 -1630 310 -1625
rect 270 -1660 310 -1655
rect 270 -1690 275 -1660
rect 275 -1690 305 -1660
rect 305 -1690 310 -1660
rect 270 -1695 310 -1690
rect 270 -1720 310 -1715
rect 270 -1750 275 -1720
rect 275 -1750 305 -1720
rect 305 -1750 310 -1720
rect 270 -1755 310 -1750
rect 270 -1785 310 -1780
rect 270 -1815 275 -1785
rect 275 -1815 305 -1785
rect 305 -1815 310 -1785
rect 270 -1820 310 -1815
rect 270 -1855 310 -1850
rect 270 -1885 275 -1855
rect 275 -1885 305 -1855
rect 305 -1885 310 -1855
rect 270 -1890 310 -1885
rect 270 -1925 310 -1920
rect 270 -1955 275 -1925
rect 275 -1955 305 -1925
rect 305 -1955 310 -1925
rect 270 -1960 310 -1955
rect 270 -1995 310 -1990
rect 270 -2025 275 -1995
rect 275 -2025 305 -1995
rect 305 -2025 310 -1995
rect 270 -2030 310 -2025
rect 270 -2060 310 -2055
rect 270 -2090 275 -2060
rect 275 -2090 305 -2060
rect 305 -2090 310 -2060
rect 270 -2095 310 -2090
rect 270 -2120 310 -2115
rect 270 -2150 275 -2120
rect 275 -2150 305 -2120
rect 305 -2150 310 -2120
rect 270 -2155 310 -2150
rect 270 -2185 310 -2180
rect 270 -2215 275 -2185
rect 275 -2215 305 -2185
rect 305 -2215 310 -2185
rect 270 -2220 310 -2215
rect 270 -2255 310 -2250
rect 270 -2285 275 -2255
rect 275 -2285 305 -2255
rect 305 -2285 310 -2255
rect 270 -2290 310 -2285
rect 270 -2325 310 -2320
rect 270 -2355 275 -2325
rect 275 -2355 305 -2325
rect 305 -2355 310 -2325
rect 270 -2360 310 -2355
rect 270 -2395 310 -2390
rect 270 -2425 275 -2395
rect 275 -2425 305 -2395
rect 305 -2425 310 -2395
rect 270 -2430 310 -2425
rect 270 -2460 310 -2455
rect 270 -2490 275 -2460
rect 275 -2490 305 -2460
rect 305 -2490 310 -2460
rect 270 -2495 310 -2490
rect 270 -2520 310 -2515
rect 270 -2550 275 -2520
rect 275 -2550 305 -2520
rect 305 -2550 310 -2520
rect 270 -2555 310 -2550
rect 270 -2585 310 -2580
rect 270 -2615 275 -2585
rect 275 -2615 305 -2585
rect 305 -2615 310 -2585
rect 270 -2620 310 -2615
rect 270 -2655 310 -2650
rect 270 -2685 275 -2655
rect 275 -2685 305 -2655
rect 305 -2685 310 -2655
rect 270 -2690 310 -2685
rect 270 -2725 310 -2720
rect 270 -2755 275 -2725
rect 275 -2755 305 -2725
rect 305 -2755 310 -2725
rect 270 -2760 310 -2755
rect 270 -2795 310 -2790
rect 270 -2825 275 -2795
rect 275 -2825 305 -2795
rect 305 -2825 310 -2795
rect 270 -2830 310 -2825
rect 270 -2860 310 -2855
rect 270 -2890 275 -2860
rect 275 -2890 305 -2860
rect 305 -2890 310 -2860
rect 270 -2895 310 -2890
rect 620 -1320 660 -1315
rect 620 -1350 625 -1320
rect 625 -1350 655 -1320
rect 655 -1350 660 -1320
rect 620 -1355 660 -1350
rect 620 -1385 660 -1380
rect 620 -1415 625 -1385
rect 625 -1415 655 -1385
rect 655 -1415 660 -1385
rect 620 -1420 660 -1415
rect 620 -1455 660 -1450
rect 620 -1485 625 -1455
rect 625 -1485 655 -1455
rect 655 -1485 660 -1455
rect 620 -1490 660 -1485
rect 620 -1525 660 -1520
rect 620 -1555 625 -1525
rect 625 -1555 655 -1525
rect 655 -1555 660 -1525
rect 620 -1560 660 -1555
rect 620 -1595 660 -1590
rect 620 -1625 625 -1595
rect 625 -1625 655 -1595
rect 655 -1625 660 -1595
rect 620 -1630 660 -1625
rect 620 -1660 660 -1655
rect 620 -1690 625 -1660
rect 625 -1690 655 -1660
rect 655 -1690 660 -1660
rect 620 -1695 660 -1690
rect 620 -1720 660 -1715
rect 620 -1750 625 -1720
rect 625 -1750 655 -1720
rect 655 -1750 660 -1720
rect 620 -1755 660 -1750
rect 620 -1785 660 -1780
rect 620 -1815 625 -1785
rect 625 -1815 655 -1785
rect 655 -1815 660 -1785
rect 620 -1820 660 -1815
rect 620 -1855 660 -1850
rect 620 -1885 625 -1855
rect 625 -1885 655 -1855
rect 655 -1885 660 -1855
rect 620 -1890 660 -1885
rect 620 -1925 660 -1920
rect 620 -1955 625 -1925
rect 625 -1955 655 -1925
rect 655 -1955 660 -1925
rect 620 -1960 660 -1955
rect 620 -1995 660 -1990
rect 620 -2025 625 -1995
rect 625 -2025 655 -1995
rect 655 -2025 660 -1995
rect 620 -2030 660 -2025
rect 620 -2060 660 -2055
rect 620 -2090 625 -2060
rect 625 -2090 655 -2060
rect 655 -2090 660 -2060
rect 620 -2095 660 -2090
rect 620 -2120 660 -2115
rect 620 -2150 625 -2120
rect 625 -2150 655 -2120
rect 655 -2150 660 -2120
rect 620 -2155 660 -2150
rect 620 -2185 660 -2180
rect 620 -2215 625 -2185
rect 625 -2215 655 -2185
rect 655 -2215 660 -2185
rect 620 -2220 660 -2215
rect 620 -2255 660 -2250
rect 620 -2285 625 -2255
rect 625 -2285 655 -2255
rect 655 -2285 660 -2255
rect 620 -2290 660 -2285
rect 620 -2325 660 -2320
rect 620 -2355 625 -2325
rect 625 -2355 655 -2325
rect 655 -2355 660 -2325
rect 620 -2360 660 -2355
rect 620 -2395 660 -2390
rect 620 -2425 625 -2395
rect 625 -2425 655 -2395
rect 655 -2425 660 -2395
rect 620 -2430 660 -2425
rect 620 -2460 660 -2455
rect 620 -2490 625 -2460
rect 625 -2490 655 -2460
rect 655 -2490 660 -2460
rect 620 -2495 660 -2490
rect 620 -2520 660 -2515
rect 620 -2550 625 -2520
rect 625 -2550 655 -2520
rect 655 -2550 660 -2520
rect 620 -2555 660 -2550
rect 620 -2585 660 -2580
rect 620 -2615 625 -2585
rect 625 -2615 655 -2585
rect 655 -2615 660 -2585
rect 620 -2620 660 -2615
rect 620 -2655 660 -2650
rect 620 -2685 625 -2655
rect 625 -2685 655 -2655
rect 655 -2685 660 -2655
rect 620 -2690 660 -2685
rect 620 -2725 660 -2720
rect 620 -2755 625 -2725
rect 625 -2755 655 -2725
rect 655 -2755 660 -2725
rect 620 -2760 660 -2755
rect 620 -2795 660 -2790
rect 620 -2825 625 -2795
rect 625 -2825 655 -2795
rect 655 -2825 660 -2795
rect 620 -2830 660 -2825
rect 620 -2860 660 -2855
rect 620 -2890 625 -2860
rect 625 -2890 655 -2860
rect 655 -2890 660 -2860
rect 620 -2895 660 -2890
rect 970 -1320 1010 -1315
rect 970 -1350 975 -1320
rect 975 -1350 1005 -1320
rect 1005 -1350 1010 -1320
rect 970 -1355 1010 -1350
rect 970 -1385 1010 -1380
rect 970 -1415 975 -1385
rect 975 -1415 1005 -1385
rect 1005 -1415 1010 -1385
rect 970 -1420 1010 -1415
rect 970 -1455 1010 -1450
rect 970 -1485 975 -1455
rect 975 -1485 1005 -1455
rect 1005 -1485 1010 -1455
rect 970 -1490 1010 -1485
rect 970 -1525 1010 -1520
rect 970 -1555 975 -1525
rect 975 -1555 1005 -1525
rect 1005 -1555 1010 -1525
rect 970 -1560 1010 -1555
rect 970 -1595 1010 -1590
rect 970 -1625 975 -1595
rect 975 -1625 1005 -1595
rect 1005 -1625 1010 -1595
rect 970 -1630 1010 -1625
rect 970 -1660 1010 -1655
rect 970 -1690 975 -1660
rect 975 -1690 1005 -1660
rect 1005 -1690 1010 -1660
rect 970 -1695 1010 -1690
rect 970 -1720 1010 -1715
rect 970 -1750 975 -1720
rect 975 -1750 1005 -1720
rect 1005 -1750 1010 -1720
rect 970 -1755 1010 -1750
rect 970 -1785 1010 -1780
rect 970 -1815 975 -1785
rect 975 -1815 1005 -1785
rect 1005 -1815 1010 -1785
rect 970 -1820 1010 -1815
rect 970 -1855 1010 -1850
rect 970 -1885 975 -1855
rect 975 -1885 1005 -1855
rect 1005 -1885 1010 -1855
rect 970 -1890 1010 -1885
rect 970 -1925 1010 -1920
rect 970 -1955 975 -1925
rect 975 -1955 1005 -1925
rect 1005 -1955 1010 -1925
rect 970 -1960 1010 -1955
rect 970 -1995 1010 -1990
rect 970 -2025 975 -1995
rect 975 -2025 1005 -1995
rect 1005 -2025 1010 -1995
rect 970 -2030 1010 -2025
rect 970 -2060 1010 -2055
rect 970 -2090 975 -2060
rect 975 -2090 1005 -2060
rect 1005 -2090 1010 -2060
rect 970 -2095 1010 -2090
rect 970 -2120 1010 -2115
rect 970 -2150 975 -2120
rect 975 -2150 1005 -2120
rect 1005 -2150 1010 -2120
rect 970 -2155 1010 -2150
rect 970 -2185 1010 -2180
rect 970 -2215 975 -2185
rect 975 -2215 1005 -2185
rect 1005 -2215 1010 -2185
rect 970 -2220 1010 -2215
rect 970 -2255 1010 -2250
rect 970 -2285 975 -2255
rect 975 -2285 1005 -2255
rect 1005 -2285 1010 -2255
rect 970 -2290 1010 -2285
rect 970 -2325 1010 -2320
rect 970 -2355 975 -2325
rect 975 -2355 1005 -2325
rect 1005 -2355 1010 -2325
rect 970 -2360 1010 -2355
rect 970 -2395 1010 -2390
rect 970 -2425 975 -2395
rect 975 -2425 1005 -2395
rect 1005 -2425 1010 -2395
rect 970 -2430 1010 -2425
rect 970 -2460 1010 -2455
rect 970 -2490 975 -2460
rect 975 -2490 1005 -2460
rect 1005 -2490 1010 -2460
rect 970 -2495 1010 -2490
rect 970 -2520 1010 -2515
rect 970 -2550 975 -2520
rect 975 -2550 1005 -2520
rect 1005 -2550 1010 -2520
rect 970 -2555 1010 -2550
rect 970 -2585 1010 -2580
rect 970 -2615 975 -2585
rect 975 -2615 1005 -2585
rect 1005 -2615 1010 -2585
rect 970 -2620 1010 -2615
rect 970 -2655 1010 -2650
rect 970 -2685 975 -2655
rect 975 -2685 1005 -2655
rect 1005 -2685 1010 -2655
rect 970 -2690 1010 -2685
rect 970 -2725 1010 -2720
rect 970 -2755 975 -2725
rect 975 -2755 1005 -2725
rect 1005 -2755 1010 -2725
rect 970 -2760 1010 -2755
rect 970 -2795 1010 -2790
rect 970 -2825 975 -2795
rect 975 -2825 1005 -2795
rect 1005 -2825 1010 -2795
rect 970 -2830 1010 -2825
rect 970 -2860 1010 -2855
rect 970 -2890 975 -2860
rect 975 -2890 1005 -2860
rect 1005 -2890 1010 -2860
rect 970 -2895 1010 -2890
rect 1320 -1320 1360 -1315
rect 1320 -1350 1325 -1320
rect 1325 -1350 1355 -1320
rect 1355 -1350 1360 -1320
rect 1320 -1355 1360 -1350
rect 1320 -1385 1360 -1380
rect 1320 -1415 1325 -1385
rect 1325 -1415 1355 -1385
rect 1355 -1415 1360 -1385
rect 1320 -1420 1360 -1415
rect 1320 -1455 1360 -1450
rect 1320 -1485 1325 -1455
rect 1325 -1485 1355 -1455
rect 1355 -1485 1360 -1455
rect 1320 -1490 1360 -1485
rect 1320 -1525 1360 -1520
rect 1320 -1555 1325 -1525
rect 1325 -1555 1355 -1525
rect 1355 -1555 1360 -1525
rect 1320 -1560 1360 -1555
rect 1320 -1595 1360 -1590
rect 1320 -1625 1325 -1595
rect 1325 -1625 1355 -1595
rect 1355 -1625 1360 -1595
rect 1320 -1630 1360 -1625
rect 1320 -1660 1360 -1655
rect 1320 -1690 1325 -1660
rect 1325 -1690 1355 -1660
rect 1355 -1690 1360 -1660
rect 1320 -1695 1360 -1690
rect 1320 -1720 1360 -1715
rect 1320 -1750 1325 -1720
rect 1325 -1750 1355 -1720
rect 1355 -1750 1360 -1720
rect 1320 -1755 1360 -1750
rect 1320 -1785 1360 -1780
rect 1320 -1815 1325 -1785
rect 1325 -1815 1355 -1785
rect 1355 -1815 1360 -1785
rect 1320 -1820 1360 -1815
rect 1320 -1855 1360 -1850
rect 1320 -1885 1325 -1855
rect 1325 -1885 1355 -1855
rect 1355 -1885 1360 -1855
rect 1320 -1890 1360 -1885
rect 1320 -1925 1360 -1920
rect 1320 -1955 1325 -1925
rect 1325 -1955 1355 -1925
rect 1355 -1955 1360 -1925
rect 1320 -1960 1360 -1955
rect 1320 -1995 1360 -1990
rect 1320 -2025 1325 -1995
rect 1325 -2025 1355 -1995
rect 1355 -2025 1360 -1995
rect 1320 -2030 1360 -2025
rect 1320 -2060 1360 -2055
rect 1320 -2090 1325 -2060
rect 1325 -2090 1355 -2060
rect 1355 -2090 1360 -2060
rect 1320 -2095 1360 -2090
rect 1320 -2120 1360 -2115
rect 1320 -2150 1325 -2120
rect 1325 -2150 1355 -2120
rect 1355 -2150 1360 -2120
rect 1320 -2155 1360 -2150
rect 1320 -2185 1360 -2180
rect 1320 -2215 1325 -2185
rect 1325 -2215 1355 -2185
rect 1355 -2215 1360 -2185
rect 1320 -2220 1360 -2215
rect 1320 -2255 1360 -2250
rect 1320 -2285 1325 -2255
rect 1325 -2285 1355 -2255
rect 1355 -2285 1360 -2255
rect 1320 -2290 1360 -2285
rect 1320 -2325 1360 -2320
rect 1320 -2355 1325 -2325
rect 1325 -2355 1355 -2325
rect 1355 -2355 1360 -2325
rect 1320 -2360 1360 -2355
rect 1320 -2395 1360 -2390
rect 1320 -2425 1325 -2395
rect 1325 -2425 1355 -2395
rect 1355 -2425 1360 -2395
rect 1320 -2430 1360 -2425
rect 1320 -2460 1360 -2455
rect 1320 -2490 1325 -2460
rect 1325 -2490 1355 -2460
rect 1355 -2490 1360 -2460
rect 1320 -2495 1360 -2490
rect 1320 -2520 1360 -2515
rect 1320 -2550 1325 -2520
rect 1325 -2550 1355 -2520
rect 1355 -2550 1360 -2520
rect 1320 -2555 1360 -2550
rect 1320 -2585 1360 -2580
rect 1320 -2615 1325 -2585
rect 1325 -2615 1355 -2585
rect 1355 -2615 1360 -2585
rect 1320 -2620 1360 -2615
rect 1320 -2655 1360 -2650
rect 1320 -2685 1325 -2655
rect 1325 -2685 1355 -2655
rect 1355 -2685 1360 -2655
rect 1320 -2690 1360 -2685
rect 1320 -2725 1360 -2720
rect 1320 -2755 1325 -2725
rect 1325 -2755 1355 -2725
rect 1355 -2755 1360 -2725
rect 1320 -2760 1360 -2755
rect 1320 -2795 1360 -2790
rect 1320 -2825 1325 -2795
rect 1325 -2825 1355 -2795
rect 1355 -2825 1360 -2795
rect 1320 -2830 1360 -2825
rect 1320 -2860 1360 -2855
rect 1320 -2890 1325 -2860
rect 1325 -2890 1355 -2860
rect 1355 -2890 1360 -2860
rect 1320 -2895 1360 -2890
rect 1670 -1320 1710 -1315
rect 1670 -1350 1675 -1320
rect 1675 -1350 1705 -1320
rect 1705 -1350 1710 -1320
rect 1670 -1355 1710 -1350
rect 1670 -1385 1710 -1380
rect 1670 -1415 1675 -1385
rect 1675 -1415 1705 -1385
rect 1705 -1415 1710 -1385
rect 1670 -1420 1710 -1415
rect 1670 -1455 1710 -1450
rect 1670 -1485 1675 -1455
rect 1675 -1485 1705 -1455
rect 1705 -1485 1710 -1455
rect 1670 -1490 1710 -1485
rect 1670 -1525 1710 -1520
rect 1670 -1555 1675 -1525
rect 1675 -1555 1705 -1525
rect 1705 -1555 1710 -1525
rect 1670 -1560 1710 -1555
rect 1670 -1595 1710 -1590
rect 1670 -1625 1675 -1595
rect 1675 -1625 1705 -1595
rect 1705 -1625 1710 -1595
rect 1670 -1630 1710 -1625
rect 1670 -1660 1710 -1655
rect 1670 -1690 1675 -1660
rect 1675 -1690 1705 -1660
rect 1705 -1690 1710 -1660
rect 1670 -1695 1710 -1690
rect 1670 -1720 1710 -1715
rect 1670 -1750 1675 -1720
rect 1675 -1750 1705 -1720
rect 1705 -1750 1710 -1720
rect 1670 -1755 1710 -1750
rect 1670 -1785 1710 -1780
rect 1670 -1815 1675 -1785
rect 1675 -1815 1705 -1785
rect 1705 -1815 1710 -1785
rect 1670 -1820 1710 -1815
rect 1670 -1855 1710 -1850
rect 1670 -1885 1675 -1855
rect 1675 -1885 1705 -1855
rect 1705 -1885 1710 -1855
rect 1670 -1890 1710 -1885
rect 1670 -1925 1710 -1920
rect 1670 -1955 1675 -1925
rect 1675 -1955 1705 -1925
rect 1705 -1955 1710 -1925
rect 1670 -1960 1710 -1955
rect 1670 -1995 1710 -1990
rect 1670 -2025 1675 -1995
rect 1675 -2025 1705 -1995
rect 1705 -2025 1710 -1995
rect 1670 -2030 1710 -2025
rect 1670 -2060 1710 -2055
rect 1670 -2090 1675 -2060
rect 1675 -2090 1705 -2060
rect 1705 -2090 1710 -2060
rect 1670 -2095 1710 -2090
rect 1670 -2120 1710 -2115
rect 1670 -2150 1675 -2120
rect 1675 -2150 1705 -2120
rect 1705 -2150 1710 -2120
rect 1670 -2155 1710 -2150
rect 1670 -2185 1710 -2180
rect 1670 -2215 1675 -2185
rect 1675 -2215 1705 -2185
rect 1705 -2215 1710 -2185
rect 1670 -2220 1710 -2215
rect 1670 -2255 1710 -2250
rect 1670 -2285 1675 -2255
rect 1675 -2285 1705 -2255
rect 1705 -2285 1710 -2255
rect 1670 -2290 1710 -2285
rect 1670 -2325 1710 -2320
rect 1670 -2355 1675 -2325
rect 1675 -2355 1705 -2325
rect 1705 -2355 1710 -2325
rect 1670 -2360 1710 -2355
rect 1670 -2395 1710 -2390
rect 1670 -2425 1675 -2395
rect 1675 -2425 1705 -2395
rect 1705 -2425 1710 -2395
rect 1670 -2430 1710 -2425
rect 1670 -2460 1710 -2455
rect 1670 -2490 1675 -2460
rect 1675 -2490 1705 -2460
rect 1705 -2490 1710 -2460
rect 1670 -2495 1710 -2490
rect 1670 -2520 1710 -2515
rect 1670 -2550 1675 -2520
rect 1675 -2550 1705 -2520
rect 1705 -2550 1710 -2520
rect 1670 -2555 1710 -2550
rect 1670 -2585 1710 -2580
rect 1670 -2615 1675 -2585
rect 1675 -2615 1705 -2585
rect 1705 -2615 1710 -2585
rect 1670 -2620 1710 -2615
rect 1670 -2655 1710 -2650
rect 1670 -2685 1675 -2655
rect 1675 -2685 1705 -2655
rect 1705 -2685 1710 -2655
rect 1670 -2690 1710 -2685
rect 1670 -2725 1710 -2720
rect 1670 -2755 1675 -2725
rect 1675 -2755 1705 -2725
rect 1705 -2755 1710 -2725
rect 1670 -2760 1710 -2755
rect 1670 -2795 1710 -2790
rect 1670 -2825 1675 -2795
rect 1675 -2825 1705 -2795
rect 1705 -2825 1710 -2795
rect 1670 -2830 1710 -2825
rect 1670 -2860 1710 -2855
rect 1670 -2890 1675 -2860
rect 1675 -2890 1705 -2860
rect 1705 -2890 1710 -2860
rect 1670 -2895 1710 -2890
rect 2020 -1320 2060 -1315
rect 2020 -1350 2025 -1320
rect 2025 -1350 2055 -1320
rect 2055 -1350 2060 -1320
rect 2020 -1355 2060 -1350
rect 2020 -1385 2060 -1380
rect 2020 -1415 2025 -1385
rect 2025 -1415 2055 -1385
rect 2055 -1415 2060 -1385
rect 2020 -1420 2060 -1415
rect 2020 -1455 2060 -1450
rect 2020 -1485 2025 -1455
rect 2025 -1485 2055 -1455
rect 2055 -1485 2060 -1455
rect 2020 -1490 2060 -1485
rect 2020 -1525 2060 -1520
rect 2020 -1555 2025 -1525
rect 2025 -1555 2055 -1525
rect 2055 -1555 2060 -1525
rect 2020 -1560 2060 -1555
rect 2020 -1595 2060 -1590
rect 2020 -1625 2025 -1595
rect 2025 -1625 2055 -1595
rect 2055 -1625 2060 -1595
rect 2020 -1630 2060 -1625
rect 2020 -1660 2060 -1655
rect 2020 -1690 2025 -1660
rect 2025 -1690 2055 -1660
rect 2055 -1690 2060 -1660
rect 2020 -1695 2060 -1690
rect 2020 -1720 2060 -1715
rect 2020 -1750 2025 -1720
rect 2025 -1750 2055 -1720
rect 2055 -1750 2060 -1720
rect 2020 -1755 2060 -1750
rect 2020 -1785 2060 -1780
rect 2020 -1815 2025 -1785
rect 2025 -1815 2055 -1785
rect 2055 -1815 2060 -1785
rect 2020 -1820 2060 -1815
rect 2020 -1855 2060 -1850
rect 2020 -1885 2025 -1855
rect 2025 -1885 2055 -1855
rect 2055 -1885 2060 -1855
rect 2020 -1890 2060 -1885
rect 2020 -1925 2060 -1920
rect 2020 -1955 2025 -1925
rect 2025 -1955 2055 -1925
rect 2055 -1955 2060 -1925
rect 2020 -1960 2060 -1955
rect 2020 -1995 2060 -1990
rect 2020 -2025 2025 -1995
rect 2025 -2025 2055 -1995
rect 2055 -2025 2060 -1995
rect 2020 -2030 2060 -2025
rect 2020 -2060 2060 -2055
rect 2020 -2090 2025 -2060
rect 2025 -2090 2055 -2060
rect 2055 -2090 2060 -2060
rect 2020 -2095 2060 -2090
rect 2020 -2120 2060 -2115
rect 2020 -2150 2025 -2120
rect 2025 -2150 2055 -2120
rect 2055 -2150 2060 -2120
rect 2020 -2155 2060 -2150
rect 2020 -2185 2060 -2180
rect 2020 -2215 2025 -2185
rect 2025 -2215 2055 -2185
rect 2055 -2215 2060 -2185
rect 2020 -2220 2060 -2215
rect 2020 -2255 2060 -2250
rect 2020 -2285 2025 -2255
rect 2025 -2285 2055 -2255
rect 2055 -2285 2060 -2255
rect 2020 -2290 2060 -2285
rect 2020 -2325 2060 -2320
rect 2020 -2355 2025 -2325
rect 2025 -2355 2055 -2325
rect 2055 -2355 2060 -2325
rect 2020 -2360 2060 -2355
rect 2020 -2395 2060 -2390
rect 2020 -2425 2025 -2395
rect 2025 -2425 2055 -2395
rect 2055 -2425 2060 -2395
rect 2020 -2430 2060 -2425
rect 2020 -2460 2060 -2455
rect 2020 -2490 2025 -2460
rect 2025 -2490 2055 -2460
rect 2055 -2490 2060 -2460
rect 2020 -2495 2060 -2490
rect 2020 -2520 2060 -2515
rect 2020 -2550 2025 -2520
rect 2025 -2550 2055 -2520
rect 2055 -2550 2060 -2520
rect 2020 -2555 2060 -2550
rect 2020 -2585 2060 -2580
rect 2020 -2615 2025 -2585
rect 2025 -2615 2055 -2585
rect 2055 -2615 2060 -2585
rect 2020 -2620 2060 -2615
rect 2020 -2655 2060 -2650
rect 2020 -2685 2025 -2655
rect 2025 -2685 2055 -2655
rect 2055 -2685 2060 -2655
rect 2020 -2690 2060 -2685
rect 2020 -2725 2060 -2720
rect 2020 -2755 2025 -2725
rect 2025 -2755 2055 -2725
rect 2055 -2755 2060 -2725
rect 2020 -2760 2060 -2755
rect 2020 -2795 2060 -2790
rect 2020 -2825 2025 -2795
rect 2025 -2825 2055 -2795
rect 2055 -2825 2060 -2795
rect 2020 -2830 2060 -2825
rect 2020 -2860 2060 -2855
rect 2020 -2890 2025 -2860
rect 2025 -2890 2055 -2860
rect 2055 -2890 2060 -2860
rect 2020 -2895 2060 -2890
rect 2370 -1320 2410 -1315
rect 2370 -1350 2375 -1320
rect 2375 -1350 2405 -1320
rect 2405 -1350 2410 -1320
rect 2370 -1355 2410 -1350
rect 2370 -1385 2410 -1380
rect 2370 -1415 2375 -1385
rect 2375 -1415 2405 -1385
rect 2405 -1415 2410 -1385
rect 2370 -1420 2410 -1415
rect 2370 -1455 2410 -1450
rect 2370 -1485 2375 -1455
rect 2375 -1485 2405 -1455
rect 2405 -1485 2410 -1455
rect 2370 -1490 2410 -1485
rect 2370 -1525 2410 -1520
rect 2370 -1555 2375 -1525
rect 2375 -1555 2405 -1525
rect 2405 -1555 2410 -1525
rect 2370 -1560 2410 -1555
rect 2370 -1595 2410 -1590
rect 2370 -1625 2375 -1595
rect 2375 -1625 2405 -1595
rect 2405 -1625 2410 -1595
rect 2370 -1630 2410 -1625
rect 2370 -1660 2410 -1655
rect 2370 -1690 2375 -1660
rect 2375 -1690 2405 -1660
rect 2405 -1690 2410 -1660
rect 2370 -1695 2410 -1690
rect 2370 -1720 2410 -1715
rect 2370 -1750 2375 -1720
rect 2375 -1750 2405 -1720
rect 2405 -1750 2410 -1720
rect 2370 -1755 2410 -1750
rect 2370 -1785 2410 -1780
rect 2370 -1815 2375 -1785
rect 2375 -1815 2405 -1785
rect 2405 -1815 2410 -1785
rect 2370 -1820 2410 -1815
rect 2370 -1855 2410 -1850
rect 2370 -1885 2375 -1855
rect 2375 -1885 2405 -1855
rect 2405 -1885 2410 -1855
rect 2370 -1890 2410 -1885
rect 2370 -1925 2410 -1920
rect 2370 -1955 2375 -1925
rect 2375 -1955 2405 -1925
rect 2405 -1955 2410 -1925
rect 2370 -1960 2410 -1955
rect 2370 -1995 2410 -1990
rect 2370 -2025 2375 -1995
rect 2375 -2025 2405 -1995
rect 2405 -2025 2410 -1995
rect 2370 -2030 2410 -2025
rect 2370 -2060 2410 -2055
rect 2370 -2090 2375 -2060
rect 2375 -2090 2405 -2060
rect 2405 -2090 2410 -2060
rect 2370 -2095 2410 -2090
rect 2370 -2120 2410 -2115
rect 2370 -2150 2375 -2120
rect 2375 -2150 2405 -2120
rect 2405 -2150 2410 -2120
rect 2370 -2155 2410 -2150
rect 2370 -2185 2410 -2180
rect 2370 -2215 2375 -2185
rect 2375 -2215 2405 -2185
rect 2405 -2215 2410 -2185
rect 2370 -2220 2410 -2215
rect 2370 -2255 2410 -2250
rect 2370 -2285 2375 -2255
rect 2375 -2285 2405 -2255
rect 2405 -2285 2410 -2255
rect 2370 -2290 2410 -2285
rect 2370 -2325 2410 -2320
rect 2370 -2355 2375 -2325
rect 2375 -2355 2405 -2325
rect 2405 -2355 2410 -2325
rect 2370 -2360 2410 -2355
rect 2370 -2395 2410 -2390
rect 2370 -2425 2375 -2395
rect 2375 -2425 2405 -2395
rect 2405 -2425 2410 -2395
rect 2370 -2430 2410 -2425
rect 2370 -2460 2410 -2455
rect 2370 -2490 2375 -2460
rect 2375 -2490 2405 -2460
rect 2405 -2490 2410 -2460
rect 2370 -2495 2410 -2490
rect 2370 -2520 2410 -2515
rect 2370 -2550 2375 -2520
rect 2375 -2550 2405 -2520
rect 2405 -2550 2410 -2520
rect 2370 -2555 2410 -2550
rect 2370 -2585 2410 -2580
rect 2370 -2615 2375 -2585
rect 2375 -2615 2405 -2585
rect 2405 -2615 2410 -2585
rect 2370 -2620 2410 -2615
rect 2370 -2655 2410 -2650
rect 2370 -2685 2375 -2655
rect 2375 -2685 2405 -2655
rect 2405 -2685 2410 -2655
rect 2370 -2690 2410 -2685
rect 2370 -2725 2410 -2720
rect 2370 -2755 2375 -2725
rect 2375 -2755 2405 -2725
rect 2405 -2755 2410 -2725
rect 2370 -2760 2410 -2755
rect 2370 -2795 2410 -2790
rect 2370 -2825 2375 -2795
rect 2375 -2825 2405 -2795
rect 2405 -2825 2410 -2795
rect 2370 -2830 2410 -2825
rect 2370 -2860 2410 -2855
rect 2370 -2890 2375 -2860
rect 2375 -2890 2405 -2860
rect 2405 -2890 2410 -2860
rect 2370 -2895 2410 -2890
rect 2720 -1320 2760 -1315
rect 2720 -1350 2725 -1320
rect 2725 -1350 2755 -1320
rect 2755 -1350 2760 -1320
rect 2720 -1355 2760 -1350
rect 2720 -1385 2760 -1380
rect 2720 -1415 2725 -1385
rect 2725 -1415 2755 -1385
rect 2755 -1415 2760 -1385
rect 2720 -1420 2760 -1415
rect 2720 -1455 2760 -1450
rect 2720 -1485 2725 -1455
rect 2725 -1485 2755 -1455
rect 2755 -1485 2760 -1455
rect 2720 -1490 2760 -1485
rect 2720 -1525 2760 -1520
rect 2720 -1555 2725 -1525
rect 2725 -1555 2755 -1525
rect 2755 -1555 2760 -1525
rect 2720 -1560 2760 -1555
rect 2720 -1595 2760 -1590
rect 2720 -1625 2725 -1595
rect 2725 -1625 2755 -1595
rect 2755 -1625 2760 -1595
rect 2720 -1630 2760 -1625
rect 2720 -1660 2760 -1655
rect 2720 -1690 2725 -1660
rect 2725 -1690 2755 -1660
rect 2755 -1690 2760 -1660
rect 2720 -1695 2760 -1690
rect 2720 -1720 2760 -1715
rect 2720 -1750 2725 -1720
rect 2725 -1750 2755 -1720
rect 2755 -1750 2760 -1720
rect 2720 -1755 2760 -1750
rect 2720 -1785 2760 -1780
rect 2720 -1815 2725 -1785
rect 2725 -1815 2755 -1785
rect 2755 -1815 2760 -1785
rect 2720 -1820 2760 -1815
rect 2720 -1855 2760 -1850
rect 2720 -1885 2725 -1855
rect 2725 -1885 2755 -1855
rect 2755 -1885 2760 -1855
rect 2720 -1890 2760 -1885
rect 2720 -1925 2760 -1920
rect 2720 -1955 2725 -1925
rect 2725 -1955 2755 -1925
rect 2755 -1955 2760 -1925
rect 2720 -1960 2760 -1955
rect 2720 -1995 2760 -1990
rect 2720 -2025 2725 -1995
rect 2725 -2025 2755 -1995
rect 2755 -2025 2760 -1995
rect 2720 -2030 2760 -2025
rect 2720 -2060 2760 -2055
rect 2720 -2090 2725 -2060
rect 2725 -2090 2755 -2060
rect 2755 -2090 2760 -2060
rect 2720 -2095 2760 -2090
rect 2720 -2120 2760 -2115
rect 2720 -2150 2725 -2120
rect 2725 -2150 2755 -2120
rect 2755 -2150 2760 -2120
rect 2720 -2155 2760 -2150
rect 2720 -2185 2760 -2180
rect 2720 -2215 2725 -2185
rect 2725 -2215 2755 -2185
rect 2755 -2215 2760 -2185
rect 2720 -2220 2760 -2215
rect 2720 -2255 2760 -2250
rect 2720 -2285 2725 -2255
rect 2725 -2285 2755 -2255
rect 2755 -2285 2760 -2255
rect 2720 -2290 2760 -2285
rect 2720 -2325 2760 -2320
rect 2720 -2355 2725 -2325
rect 2725 -2355 2755 -2325
rect 2755 -2355 2760 -2325
rect 2720 -2360 2760 -2355
rect 2720 -2395 2760 -2390
rect 2720 -2425 2725 -2395
rect 2725 -2425 2755 -2395
rect 2755 -2425 2760 -2395
rect 2720 -2430 2760 -2425
rect 2720 -2460 2760 -2455
rect 2720 -2490 2725 -2460
rect 2725 -2490 2755 -2460
rect 2755 -2490 2760 -2460
rect 2720 -2495 2760 -2490
rect 2720 -2520 2760 -2515
rect 2720 -2550 2725 -2520
rect 2725 -2550 2755 -2520
rect 2755 -2550 2760 -2520
rect 2720 -2555 2760 -2550
rect 2720 -2585 2760 -2580
rect 2720 -2615 2725 -2585
rect 2725 -2615 2755 -2585
rect 2755 -2615 2760 -2585
rect 2720 -2620 2760 -2615
rect 2720 -2655 2760 -2650
rect 2720 -2685 2725 -2655
rect 2725 -2685 2755 -2655
rect 2755 -2685 2760 -2655
rect 2720 -2690 2760 -2685
rect 2720 -2725 2760 -2720
rect 2720 -2755 2725 -2725
rect 2725 -2755 2755 -2725
rect 2755 -2755 2760 -2725
rect 2720 -2760 2760 -2755
rect 2720 -2795 2760 -2790
rect 2720 -2825 2725 -2795
rect 2725 -2825 2755 -2795
rect 2755 -2825 2760 -2795
rect 2720 -2830 2760 -2825
rect 2720 -2860 2760 -2855
rect 2720 -2890 2725 -2860
rect 2725 -2890 2755 -2860
rect 2755 -2890 2760 -2860
rect 2720 -2895 2760 -2890
rect 3070 -1320 3110 -1315
rect 3070 -1350 3075 -1320
rect 3075 -1350 3105 -1320
rect 3105 -1350 3110 -1320
rect 3070 -1355 3110 -1350
rect 3070 -1385 3110 -1380
rect 3070 -1415 3075 -1385
rect 3075 -1415 3105 -1385
rect 3105 -1415 3110 -1385
rect 3070 -1420 3110 -1415
rect 3070 -1455 3110 -1450
rect 3070 -1485 3075 -1455
rect 3075 -1485 3105 -1455
rect 3105 -1485 3110 -1455
rect 3070 -1490 3110 -1485
rect 3070 -1525 3110 -1520
rect 3070 -1555 3075 -1525
rect 3075 -1555 3105 -1525
rect 3105 -1555 3110 -1525
rect 3070 -1560 3110 -1555
rect 3070 -1595 3110 -1590
rect 3070 -1625 3075 -1595
rect 3075 -1625 3105 -1595
rect 3105 -1625 3110 -1595
rect 3070 -1630 3110 -1625
rect 3070 -1660 3110 -1655
rect 3070 -1690 3075 -1660
rect 3075 -1690 3105 -1660
rect 3105 -1690 3110 -1660
rect 3070 -1695 3110 -1690
rect 3070 -1720 3110 -1715
rect 3070 -1750 3075 -1720
rect 3075 -1750 3105 -1720
rect 3105 -1750 3110 -1720
rect 3070 -1755 3110 -1750
rect 3070 -1785 3110 -1780
rect 3070 -1815 3075 -1785
rect 3075 -1815 3105 -1785
rect 3105 -1815 3110 -1785
rect 3070 -1820 3110 -1815
rect 3070 -1855 3110 -1850
rect 3070 -1885 3075 -1855
rect 3075 -1885 3105 -1855
rect 3105 -1885 3110 -1855
rect 3070 -1890 3110 -1885
rect 3070 -1925 3110 -1920
rect 3070 -1955 3075 -1925
rect 3075 -1955 3105 -1925
rect 3105 -1955 3110 -1925
rect 3070 -1960 3110 -1955
rect 3070 -1995 3110 -1990
rect 3070 -2025 3075 -1995
rect 3075 -2025 3105 -1995
rect 3105 -2025 3110 -1995
rect 3070 -2030 3110 -2025
rect 3070 -2060 3110 -2055
rect 3070 -2090 3075 -2060
rect 3075 -2090 3105 -2060
rect 3105 -2090 3110 -2060
rect 3070 -2095 3110 -2090
rect 3070 -2120 3110 -2115
rect 3070 -2150 3075 -2120
rect 3075 -2150 3105 -2120
rect 3105 -2150 3110 -2120
rect 3070 -2155 3110 -2150
rect 3070 -2185 3110 -2180
rect 3070 -2215 3075 -2185
rect 3075 -2215 3105 -2185
rect 3105 -2215 3110 -2185
rect 3070 -2220 3110 -2215
rect 3070 -2255 3110 -2250
rect 3070 -2285 3075 -2255
rect 3075 -2285 3105 -2255
rect 3105 -2285 3110 -2255
rect 3070 -2290 3110 -2285
rect 3070 -2325 3110 -2320
rect 3070 -2355 3075 -2325
rect 3075 -2355 3105 -2325
rect 3105 -2355 3110 -2325
rect 3070 -2360 3110 -2355
rect 3070 -2395 3110 -2390
rect 3070 -2425 3075 -2395
rect 3075 -2425 3105 -2395
rect 3105 -2425 3110 -2395
rect 3070 -2430 3110 -2425
rect 3070 -2460 3110 -2455
rect 3070 -2490 3075 -2460
rect 3075 -2490 3105 -2460
rect 3105 -2490 3110 -2460
rect 3070 -2495 3110 -2490
rect 3070 -2520 3110 -2515
rect 3070 -2550 3075 -2520
rect 3075 -2550 3105 -2520
rect 3105 -2550 3110 -2520
rect 3070 -2555 3110 -2550
rect 3070 -2585 3110 -2580
rect 3070 -2615 3075 -2585
rect 3075 -2615 3105 -2585
rect 3105 -2615 3110 -2585
rect 3070 -2620 3110 -2615
rect 3070 -2655 3110 -2650
rect 3070 -2685 3075 -2655
rect 3075 -2685 3105 -2655
rect 3105 -2685 3110 -2655
rect 3070 -2690 3110 -2685
rect 3070 -2725 3110 -2720
rect 3070 -2755 3075 -2725
rect 3075 -2755 3105 -2725
rect 3105 -2755 3110 -2725
rect 3070 -2760 3110 -2755
rect 3070 -2795 3110 -2790
rect 3070 -2825 3075 -2795
rect 3075 -2825 3105 -2795
rect 3105 -2825 3110 -2795
rect 3070 -2830 3110 -2825
rect 3070 -2860 3110 -2855
rect 3070 -2890 3075 -2860
rect 3075 -2890 3105 -2860
rect 3105 -2890 3110 -2860
rect 3070 -2895 3110 -2890
rect 5870 -1320 5910 -1315
rect 5870 -1350 5875 -1320
rect 5875 -1350 5905 -1320
rect 5905 -1350 5910 -1320
rect 5870 -1355 5910 -1350
rect 5870 -1385 5910 -1380
rect 5870 -1415 5875 -1385
rect 5875 -1415 5905 -1385
rect 5905 -1415 5910 -1385
rect 5870 -1420 5910 -1415
rect 5870 -1455 5910 -1450
rect 5870 -1485 5875 -1455
rect 5875 -1485 5905 -1455
rect 5905 -1485 5910 -1455
rect 5870 -1490 5910 -1485
rect 5870 -1525 5910 -1520
rect 5870 -1555 5875 -1525
rect 5875 -1555 5905 -1525
rect 5905 -1555 5910 -1525
rect 5870 -1560 5910 -1555
rect 5870 -1595 5910 -1590
rect 5870 -1625 5875 -1595
rect 5875 -1625 5905 -1595
rect 5905 -1625 5910 -1595
rect 5870 -1630 5910 -1625
rect 5870 -1660 5910 -1655
rect 5870 -1690 5875 -1660
rect 5875 -1690 5905 -1660
rect 5905 -1690 5910 -1660
rect 5870 -1695 5910 -1690
rect 5870 -1720 5910 -1715
rect 5870 -1750 5875 -1720
rect 5875 -1750 5905 -1720
rect 5905 -1750 5910 -1720
rect 5870 -1755 5910 -1750
rect 5870 -1785 5910 -1780
rect 5870 -1815 5875 -1785
rect 5875 -1815 5905 -1785
rect 5905 -1815 5910 -1785
rect 5870 -1820 5910 -1815
rect 5870 -1855 5910 -1850
rect 5870 -1885 5875 -1855
rect 5875 -1885 5905 -1855
rect 5905 -1885 5910 -1855
rect 5870 -1890 5910 -1885
rect 5870 -1925 5910 -1920
rect 5870 -1955 5875 -1925
rect 5875 -1955 5905 -1925
rect 5905 -1955 5910 -1925
rect 5870 -1960 5910 -1955
rect 5870 -1995 5910 -1990
rect 5870 -2025 5875 -1995
rect 5875 -2025 5905 -1995
rect 5905 -2025 5910 -1995
rect 5870 -2030 5910 -2025
rect 5870 -2060 5910 -2055
rect 5870 -2090 5875 -2060
rect 5875 -2090 5905 -2060
rect 5905 -2090 5910 -2060
rect 5870 -2095 5910 -2090
rect 5870 -2120 5910 -2115
rect 5870 -2150 5875 -2120
rect 5875 -2150 5905 -2120
rect 5905 -2150 5910 -2120
rect 5870 -2155 5910 -2150
rect 5870 -2185 5910 -2180
rect 5870 -2215 5875 -2185
rect 5875 -2215 5905 -2185
rect 5905 -2215 5910 -2185
rect 5870 -2220 5910 -2215
rect 5870 -2255 5910 -2250
rect 5870 -2285 5875 -2255
rect 5875 -2285 5905 -2255
rect 5905 -2285 5910 -2255
rect 5870 -2290 5910 -2285
rect 5870 -2325 5910 -2320
rect 5870 -2355 5875 -2325
rect 5875 -2355 5905 -2325
rect 5905 -2355 5910 -2325
rect 5870 -2360 5910 -2355
rect 5870 -2395 5910 -2390
rect 5870 -2425 5875 -2395
rect 5875 -2425 5905 -2395
rect 5905 -2425 5910 -2395
rect 5870 -2430 5910 -2425
rect 5870 -2460 5910 -2455
rect 5870 -2490 5875 -2460
rect 5875 -2490 5905 -2460
rect 5905 -2490 5910 -2460
rect 5870 -2495 5910 -2490
rect 5870 -2520 5910 -2515
rect 5870 -2550 5875 -2520
rect 5875 -2550 5905 -2520
rect 5905 -2550 5910 -2520
rect 5870 -2555 5910 -2550
rect 5870 -2585 5910 -2580
rect 5870 -2615 5875 -2585
rect 5875 -2615 5905 -2585
rect 5905 -2615 5910 -2585
rect 5870 -2620 5910 -2615
rect 5870 -2655 5910 -2650
rect 5870 -2685 5875 -2655
rect 5875 -2685 5905 -2655
rect 5905 -2685 5910 -2655
rect 5870 -2690 5910 -2685
rect 5870 -2725 5910 -2720
rect 5870 -2755 5875 -2725
rect 5875 -2755 5905 -2725
rect 5905 -2755 5910 -2725
rect 5870 -2760 5910 -2755
rect 5870 -2795 5910 -2790
rect 5870 -2825 5875 -2795
rect 5875 -2825 5905 -2795
rect 5905 -2825 5910 -2795
rect 5870 -2830 5910 -2825
rect 5870 -2860 5910 -2855
rect 5870 -2890 5875 -2860
rect 5875 -2890 5905 -2860
rect 5905 -2890 5910 -2860
rect 5870 -2895 5910 -2890
rect 6220 -1320 6260 -1315
rect 6220 -1350 6225 -1320
rect 6225 -1350 6255 -1320
rect 6255 -1350 6260 -1320
rect 6220 -1355 6260 -1350
rect 6220 -1385 6260 -1380
rect 6220 -1415 6225 -1385
rect 6225 -1415 6255 -1385
rect 6255 -1415 6260 -1385
rect 6220 -1420 6260 -1415
rect 6220 -1455 6260 -1450
rect 6220 -1485 6225 -1455
rect 6225 -1485 6255 -1455
rect 6255 -1485 6260 -1455
rect 6220 -1490 6260 -1485
rect 6220 -1525 6260 -1520
rect 6220 -1555 6225 -1525
rect 6225 -1555 6255 -1525
rect 6255 -1555 6260 -1525
rect 6220 -1560 6260 -1555
rect 6220 -1595 6260 -1590
rect 6220 -1625 6225 -1595
rect 6225 -1625 6255 -1595
rect 6255 -1625 6260 -1595
rect 6220 -1630 6260 -1625
rect 6220 -1660 6260 -1655
rect 6220 -1690 6225 -1660
rect 6225 -1690 6255 -1660
rect 6255 -1690 6260 -1660
rect 6220 -1695 6260 -1690
rect 6220 -1720 6260 -1715
rect 6220 -1750 6225 -1720
rect 6225 -1750 6255 -1720
rect 6255 -1750 6260 -1720
rect 6220 -1755 6260 -1750
rect 6220 -1785 6260 -1780
rect 6220 -1815 6225 -1785
rect 6225 -1815 6255 -1785
rect 6255 -1815 6260 -1785
rect 6220 -1820 6260 -1815
rect 6220 -1855 6260 -1850
rect 6220 -1885 6225 -1855
rect 6225 -1885 6255 -1855
rect 6255 -1885 6260 -1855
rect 6220 -1890 6260 -1885
rect 6220 -1925 6260 -1920
rect 6220 -1955 6225 -1925
rect 6225 -1955 6255 -1925
rect 6255 -1955 6260 -1925
rect 6220 -1960 6260 -1955
rect 6220 -1995 6260 -1990
rect 6220 -2025 6225 -1995
rect 6225 -2025 6255 -1995
rect 6255 -2025 6260 -1995
rect 6220 -2030 6260 -2025
rect 6220 -2060 6260 -2055
rect 6220 -2090 6225 -2060
rect 6225 -2090 6255 -2060
rect 6255 -2090 6260 -2060
rect 6220 -2095 6260 -2090
rect 6220 -2120 6260 -2115
rect 6220 -2150 6225 -2120
rect 6225 -2150 6255 -2120
rect 6255 -2150 6260 -2120
rect 6220 -2155 6260 -2150
rect 6220 -2185 6260 -2180
rect 6220 -2215 6225 -2185
rect 6225 -2215 6255 -2185
rect 6255 -2215 6260 -2185
rect 6220 -2220 6260 -2215
rect 6220 -2255 6260 -2250
rect 6220 -2285 6225 -2255
rect 6225 -2285 6255 -2255
rect 6255 -2285 6260 -2255
rect 6220 -2290 6260 -2285
rect 6220 -2325 6260 -2320
rect 6220 -2355 6225 -2325
rect 6225 -2355 6255 -2325
rect 6255 -2355 6260 -2325
rect 6220 -2360 6260 -2355
rect 6220 -2395 6260 -2390
rect 6220 -2425 6225 -2395
rect 6225 -2425 6255 -2395
rect 6255 -2425 6260 -2395
rect 6220 -2430 6260 -2425
rect 6220 -2460 6260 -2455
rect 6220 -2490 6225 -2460
rect 6225 -2490 6255 -2460
rect 6255 -2490 6260 -2460
rect 6220 -2495 6260 -2490
rect 6220 -2520 6260 -2515
rect 6220 -2550 6225 -2520
rect 6225 -2550 6255 -2520
rect 6255 -2550 6260 -2520
rect 6220 -2555 6260 -2550
rect 6220 -2585 6260 -2580
rect 6220 -2615 6225 -2585
rect 6225 -2615 6255 -2585
rect 6255 -2615 6260 -2585
rect 6220 -2620 6260 -2615
rect 6220 -2655 6260 -2650
rect 6220 -2685 6225 -2655
rect 6225 -2685 6255 -2655
rect 6255 -2685 6260 -2655
rect 6220 -2690 6260 -2685
rect 6220 -2725 6260 -2720
rect 6220 -2755 6225 -2725
rect 6225 -2755 6255 -2725
rect 6255 -2755 6260 -2725
rect 6220 -2760 6260 -2755
rect 6220 -2795 6260 -2790
rect 6220 -2825 6225 -2795
rect 6225 -2825 6255 -2795
rect 6255 -2825 6260 -2795
rect 6220 -2830 6260 -2825
rect 6220 -2860 6260 -2855
rect 6220 -2890 6225 -2860
rect 6225 -2890 6255 -2860
rect 6255 -2890 6260 -2860
rect 6220 -2895 6260 -2890
rect 6570 -1320 6610 -1315
rect 6570 -1350 6575 -1320
rect 6575 -1350 6605 -1320
rect 6605 -1350 6610 -1320
rect 6570 -1355 6610 -1350
rect 6570 -1385 6610 -1380
rect 6570 -1415 6575 -1385
rect 6575 -1415 6605 -1385
rect 6605 -1415 6610 -1385
rect 6570 -1420 6610 -1415
rect 6570 -1455 6610 -1450
rect 6570 -1485 6575 -1455
rect 6575 -1485 6605 -1455
rect 6605 -1485 6610 -1455
rect 6570 -1490 6610 -1485
rect 6570 -1525 6610 -1520
rect 6570 -1555 6575 -1525
rect 6575 -1555 6605 -1525
rect 6605 -1555 6610 -1525
rect 6570 -1560 6610 -1555
rect 6570 -1595 6610 -1590
rect 6570 -1625 6575 -1595
rect 6575 -1625 6605 -1595
rect 6605 -1625 6610 -1595
rect 6570 -1630 6610 -1625
rect 6570 -1660 6610 -1655
rect 6570 -1690 6575 -1660
rect 6575 -1690 6605 -1660
rect 6605 -1690 6610 -1660
rect 6570 -1695 6610 -1690
rect 6570 -1720 6610 -1715
rect 6570 -1750 6575 -1720
rect 6575 -1750 6605 -1720
rect 6605 -1750 6610 -1720
rect 6570 -1755 6610 -1750
rect 6570 -1785 6610 -1780
rect 6570 -1815 6575 -1785
rect 6575 -1815 6605 -1785
rect 6605 -1815 6610 -1785
rect 6570 -1820 6610 -1815
rect 6570 -1855 6610 -1850
rect 6570 -1885 6575 -1855
rect 6575 -1885 6605 -1855
rect 6605 -1885 6610 -1855
rect 6570 -1890 6610 -1885
rect 6570 -1925 6610 -1920
rect 6570 -1955 6575 -1925
rect 6575 -1955 6605 -1925
rect 6605 -1955 6610 -1925
rect 6570 -1960 6610 -1955
rect 6570 -1995 6610 -1990
rect 6570 -2025 6575 -1995
rect 6575 -2025 6605 -1995
rect 6605 -2025 6610 -1995
rect 6570 -2030 6610 -2025
rect 6570 -2060 6610 -2055
rect 6570 -2090 6575 -2060
rect 6575 -2090 6605 -2060
rect 6605 -2090 6610 -2060
rect 6570 -2095 6610 -2090
rect 6570 -2120 6610 -2115
rect 6570 -2150 6575 -2120
rect 6575 -2150 6605 -2120
rect 6605 -2150 6610 -2120
rect 6570 -2155 6610 -2150
rect 6570 -2185 6610 -2180
rect 6570 -2215 6575 -2185
rect 6575 -2215 6605 -2185
rect 6605 -2215 6610 -2185
rect 6570 -2220 6610 -2215
rect 6570 -2255 6610 -2250
rect 6570 -2285 6575 -2255
rect 6575 -2285 6605 -2255
rect 6605 -2285 6610 -2255
rect 6570 -2290 6610 -2285
rect 6570 -2325 6610 -2320
rect 6570 -2355 6575 -2325
rect 6575 -2355 6605 -2325
rect 6605 -2355 6610 -2325
rect 6570 -2360 6610 -2355
rect 6570 -2395 6610 -2390
rect 6570 -2425 6575 -2395
rect 6575 -2425 6605 -2395
rect 6605 -2425 6610 -2395
rect 6570 -2430 6610 -2425
rect 6570 -2460 6610 -2455
rect 6570 -2490 6575 -2460
rect 6575 -2490 6605 -2460
rect 6605 -2490 6610 -2460
rect 6570 -2495 6610 -2490
rect 6570 -2520 6610 -2515
rect 6570 -2550 6575 -2520
rect 6575 -2550 6605 -2520
rect 6605 -2550 6610 -2520
rect 6570 -2555 6610 -2550
rect 6570 -2585 6610 -2580
rect 6570 -2615 6575 -2585
rect 6575 -2615 6605 -2585
rect 6605 -2615 6610 -2585
rect 6570 -2620 6610 -2615
rect 6570 -2655 6610 -2650
rect 6570 -2685 6575 -2655
rect 6575 -2685 6605 -2655
rect 6605 -2685 6610 -2655
rect 6570 -2690 6610 -2685
rect 6570 -2725 6610 -2720
rect 6570 -2755 6575 -2725
rect 6575 -2755 6605 -2725
rect 6605 -2755 6610 -2725
rect 6570 -2760 6610 -2755
rect 6570 -2795 6610 -2790
rect 6570 -2825 6575 -2795
rect 6575 -2825 6605 -2795
rect 6605 -2825 6610 -2795
rect 6570 -2830 6610 -2825
rect 6570 -2860 6610 -2855
rect 6570 -2890 6575 -2860
rect 6575 -2890 6605 -2860
rect 6605 -2890 6610 -2860
rect 6570 -2895 6610 -2890
rect 6920 -1320 6960 -1315
rect 6920 -1350 6925 -1320
rect 6925 -1350 6955 -1320
rect 6955 -1350 6960 -1320
rect 6920 -1355 6960 -1350
rect 6920 -1385 6960 -1380
rect 6920 -1415 6925 -1385
rect 6925 -1415 6955 -1385
rect 6955 -1415 6960 -1385
rect 6920 -1420 6960 -1415
rect 6920 -1455 6960 -1450
rect 6920 -1485 6925 -1455
rect 6925 -1485 6955 -1455
rect 6955 -1485 6960 -1455
rect 6920 -1490 6960 -1485
rect 6920 -1525 6960 -1520
rect 6920 -1555 6925 -1525
rect 6925 -1555 6955 -1525
rect 6955 -1555 6960 -1525
rect 6920 -1560 6960 -1555
rect 6920 -1595 6960 -1590
rect 6920 -1625 6925 -1595
rect 6925 -1625 6955 -1595
rect 6955 -1625 6960 -1595
rect 6920 -1630 6960 -1625
rect 6920 -1660 6960 -1655
rect 6920 -1690 6925 -1660
rect 6925 -1690 6955 -1660
rect 6955 -1690 6960 -1660
rect 6920 -1695 6960 -1690
rect 6920 -1720 6960 -1715
rect 6920 -1750 6925 -1720
rect 6925 -1750 6955 -1720
rect 6955 -1750 6960 -1720
rect 6920 -1755 6960 -1750
rect 6920 -1785 6960 -1780
rect 6920 -1815 6925 -1785
rect 6925 -1815 6955 -1785
rect 6955 -1815 6960 -1785
rect 6920 -1820 6960 -1815
rect 6920 -1855 6960 -1850
rect 6920 -1885 6925 -1855
rect 6925 -1885 6955 -1855
rect 6955 -1885 6960 -1855
rect 6920 -1890 6960 -1885
rect 6920 -1925 6960 -1920
rect 6920 -1955 6925 -1925
rect 6925 -1955 6955 -1925
rect 6955 -1955 6960 -1925
rect 6920 -1960 6960 -1955
rect 6920 -1995 6960 -1990
rect 6920 -2025 6925 -1995
rect 6925 -2025 6955 -1995
rect 6955 -2025 6960 -1995
rect 6920 -2030 6960 -2025
rect 6920 -2060 6960 -2055
rect 6920 -2090 6925 -2060
rect 6925 -2090 6955 -2060
rect 6955 -2090 6960 -2060
rect 6920 -2095 6960 -2090
rect 6920 -2120 6960 -2115
rect 6920 -2150 6925 -2120
rect 6925 -2150 6955 -2120
rect 6955 -2150 6960 -2120
rect 6920 -2155 6960 -2150
rect 6920 -2185 6960 -2180
rect 6920 -2215 6925 -2185
rect 6925 -2215 6955 -2185
rect 6955 -2215 6960 -2185
rect 6920 -2220 6960 -2215
rect 6920 -2255 6960 -2250
rect 6920 -2285 6925 -2255
rect 6925 -2285 6955 -2255
rect 6955 -2285 6960 -2255
rect 6920 -2290 6960 -2285
rect 6920 -2325 6960 -2320
rect 6920 -2355 6925 -2325
rect 6925 -2355 6955 -2325
rect 6955 -2355 6960 -2325
rect 6920 -2360 6960 -2355
rect 6920 -2395 6960 -2390
rect 6920 -2425 6925 -2395
rect 6925 -2425 6955 -2395
rect 6955 -2425 6960 -2395
rect 6920 -2430 6960 -2425
rect 6920 -2460 6960 -2455
rect 6920 -2490 6925 -2460
rect 6925 -2490 6955 -2460
rect 6955 -2490 6960 -2460
rect 6920 -2495 6960 -2490
rect 6920 -2520 6960 -2515
rect 6920 -2550 6925 -2520
rect 6925 -2550 6955 -2520
rect 6955 -2550 6960 -2520
rect 6920 -2555 6960 -2550
rect 6920 -2585 6960 -2580
rect 6920 -2615 6925 -2585
rect 6925 -2615 6955 -2585
rect 6955 -2615 6960 -2585
rect 6920 -2620 6960 -2615
rect 6920 -2655 6960 -2650
rect 6920 -2685 6925 -2655
rect 6925 -2685 6955 -2655
rect 6955 -2685 6960 -2655
rect 6920 -2690 6960 -2685
rect 6920 -2725 6960 -2720
rect 6920 -2755 6925 -2725
rect 6925 -2755 6955 -2725
rect 6955 -2755 6960 -2725
rect 6920 -2760 6960 -2755
rect 6920 -2795 6960 -2790
rect 6920 -2825 6925 -2795
rect 6925 -2825 6955 -2795
rect 6955 -2825 6960 -2795
rect 6920 -2830 6960 -2825
rect 6920 -2860 6960 -2855
rect 6920 -2890 6925 -2860
rect 6925 -2890 6955 -2860
rect 6955 -2890 6960 -2860
rect 6920 -2895 6960 -2890
rect 7270 -1320 7310 -1315
rect 7270 -1350 7275 -1320
rect 7275 -1350 7305 -1320
rect 7305 -1350 7310 -1320
rect 7270 -1355 7310 -1350
rect 7270 -1385 7310 -1380
rect 7270 -1415 7275 -1385
rect 7275 -1415 7305 -1385
rect 7305 -1415 7310 -1385
rect 7270 -1420 7310 -1415
rect 7270 -1455 7310 -1450
rect 7270 -1485 7275 -1455
rect 7275 -1485 7305 -1455
rect 7305 -1485 7310 -1455
rect 7270 -1490 7310 -1485
rect 7270 -1525 7310 -1520
rect 7270 -1555 7275 -1525
rect 7275 -1555 7305 -1525
rect 7305 -1555 7310 -1525
rect 7270 -1560 7310 -1555
rect 7270 -1595 7310 -1590
rect 7270 -1625 7275 -1595
rect 7275 -1625 7305 -1595
rect 7305 -1625 7310 -1595
rect 7270 -1630 7310 -1625
rect 7270 -1660 7310 -1655
rect 7270 -1690 7275 -1660
rect 7275 -1690 7305 -1660
rect 7305 -1690 7310 -1660
rect 7270 -1695 7310 -1690
rect 7270 -1720 7310 -1715
rect 7270 -1750 7275 -1720
rect 7275 -1750 7305 -1720
rect 7305 -1750 7310 -1720
rect 7270 -1755 7310 -1750
rect 7270 -1785 7310 -1780
rect 7270 -1815 7275 -1785
rect 7275 -1815 7305 -1785
rect 7305 -1815 7310 -1785
rect 7270 -1820 7310 -1815
rect 7270 -1855 7310 -1850
rect 7270 -1885 7275 -1855
rect 7275 -1885 7305 -1855
rect 7305 -1885 7310 -1855
rect 7270 -1890 7310 -1885
rect 7270 -1925 7310 -1920
rect 7270 -1955 7275 -1925
rect 7275 -1955 7305 -1925
rect 7305 -1955 7310 -1925
rect 7270 -1960 7310 -1955
rect 7270 -1995 7310 -1990
rect 7270 -2025 7275 -1995
rect 7275 -2025 7305 -1995
rect 7305 -2025 7310 -1995
rect 7270 -2030 7310 -2025
rect 7270 -2060 7310 -2055
rect 7270 -2090 7275 -2060
rect 7275 -2090 7305 -2060
rect 7305 -2090 7310 -2060
rect 7270 -2095 7310 -2090
rect 7270 -2120 7310 -2115
rect 7270 -2150 7275 -2120
rect 7275 -2150 7305 -2120
rect 7305 -2150 7310 -2120
rect 7270 -2155 7310 -2150
rect 7270 -2185 7310 -2180
rect 7270 -2215 7275 -2185
rect 7275 -2215 7305 -2185
rect 7305 -2215 7310 -2185
rect 7270 -2220 7310 -2215
rect 7270 -2255 7310 -2250
rect 7270 -2285 7275 -2255
rect 7275 -2285 7305 -2255
rect 7305 -2285 7310 -2255
rect 7270 -2290 7310 -2285
rect 7270 -2325 7310 -2320
rect 7270 -2355 7275 -2325
rect 7275 -2355 7305 -2325
rect 7305 -2355 7310 -2325
rect 7270 -2360 7310 -2355
rect 7270 -2395 7310 -2390
rect 7270 -2425 7275 -2395
rect 7275 -2425 7305 -2395
rect 7305 -2425 7310 -2395
rect 7270 -2430 7310 -2425
rect 7270 -2460 7310 -2455
rect 7270 -2490 7275 -2460
rect 7275 -2490 7305 -2460
rect 7305 -2490 7310 -2460
rect 7270 -2495 7310 -2490
rect 7270 -2520 7310 -2515
rect 7270 -2550 7275 -2520
rect 7275 -2550 7305 -2520
rect 7305 -2550 7310 -2520
rect 7270 -2555 7310 -2550
rect 7270 -2585 7310 -2580
rect 7270 -2615 7275 -2585
rect 7275 -2615 7305 -2585
rect 7305 -2615 7310 -2585
rect 7270 -2620 7310 -2615
rect 7270 -2655 7310 -2650
rect 7270 -2685 7275 -2655
rect 7275 -2685 7305 -2655
rect 7305 -2685 7310 -2655
rect 7270 -2690 7310 -2685
rect 7270 -2725 7310 -2720
rect 7270 -2755 7275 -2725
rect 7275 -2755 7305 -2725
rect 7305 -2755 7310 -2725
rect 7270 -2760 7310 -2755
rect 7270 -2795 7310 -2790
rect 7270 -2825 7275 -2795
rect 7275 -2825 7305 -2795
rect 7305 -2825 7310 -2795
rect 7270 -2830 7310 -2825
rect 7270 -2860 7310 -2855
rect 7270 -2890 7275 -2860
rect 7275 -2890 7305 -2860
rect 7305 -2890 7310 -2860
rect 7270 -2895 7310 -2890
rect 7620 -1320 7660 -1315
rect 7620 -1350 7625 -1320
rect 7625 -1350 7655 -1320
rect 7655 -1350 7660 -1320
rect 7620 -1355 7660 -1350
rect 7620 -1385 7660 -1380
rect 7620 -1415 7625 -1385
rect 7625 -1415 7655 -1385
rect 7655 -1415 7660 -1385
rect 7620 -1420 7660 -1415
rect 7620 -1455 7660 -1450
rect 7620 -1485 7625 -1455
rect 7625 -1485 7655 -1455
rect 7655 -1485 7660 -1455
rect 7620 -1490 7660 -1485
rect 7620 -1525 7660 -1520
rect 7620 -1555 7625 -1525
rect 7625 -1555 7655 -1525
rect 7655 -1555 7660 -1525
rect 7620 -1560 7660 -1555
rect 7620 -1595 7660 -1590
rect 7620 -1625 7625 -1595
rect 7625 -1625 7655 -1595
rect 7655 -1625 7660 -1595
rect 7620 -1630 7660 -1625
rect 7620 -1660 7660 -1655
rect 7620 -1690 7625 -1660
rect 7625 -1690 7655 -1660
rect 7655 -1690 7660 -1660
rect 7620 -1695 7660 -1690
rect 7620 -1720 7660 -1715
rect 7620 -1750 7625 -1720
rect 7625 -1750 7655 -1720
rect 7655 -1750 7660 -1720
rect 7620 -1755 7660 -1750
rect 7620 -1785 7660 -1780
rect 7620 -1815 7625 -1785
rect 7625 -1815 7655 -1785
rect 7655 -1815 7660 -1785
rect 7620 -1820 7660 -1815
rect 7620 -1855 7660 -1850
rect 7620 -1885 7625 -1855
rect 7625 -1885 7655 -1855
rect 7655 -1885 7660 -1855
rect 7620 -1890 7660 -1885
rect 7620 -1925 7660 -1920
rect 7620 -1955 7625 -1925
rect 7625 -1955 7655 -1925
rect 7655 -1955 7660 -1925
rect 7620 -1960 7660 -1955
rect 7620 -1995 7660 -1990
rect 7620 -2025 7625 -1995
rect 7625 -2025 7655 -1995
rect 7655 -2025 7660 -1995
rect 7620 -2030 7660 -2025
rect 7620 -2060 7660 -2055
rect 7620 -2090 7625 -2060
rect 7625 -2090 7655 -2060
rect 7655 -2090 7660 -2060
rect 7620 -2095 7660 -2090
rect 7620 -2120 7660 -2115
rect 7620 -2150 7625 -2120
rect 7625 -2150 7655 -2120
rect 7655 -2150 7660 -2120
rect 7620 -2155 7660 -2150
rect 7620 -2185 7660 -2180
rect 7620 -2215 7625 -2185
rect 7625 -2215 7655 -2185
rect 7655 -2215 7660 -2185
rect 7620 -2220 7660 -2215
rect 7620 -2255 7660 -2250
rect 7620 -2285 7625 -2255
rect 7625 -2285 7655 -2255
rect 7655 -2285 7660 -2255
rect 7620 -2290 7660 -2285
rect 7620 -2325 7660 -2320
rect 7620 -2355 7625 -2325
rect 7625 -2355 7655 -2325
rect 7655 -2355 7660 -2325
rect 7620 -2360 7660 -2355
rect 7620 -2395 7660 -2390
rect 7620 -2425 7625 -2395
rect 7625 -2425 7655 -2395
rect 7655 -2425 7660 -2395
rect 7620 -2430 7660 -2425
rect 7620 -2460 7660 -2455
rect 7620 -2490 7625 -2460
rect 7625 -2490 7655 -2460
rect 7655 -2490 7660 -2460
rect 7620 -2495 7660 -2490
rect 7620 -2520 7660 -2515
rect 7620 -2550 7625 -2520
rect 7625 -2550 7655 -2520
rect 7655 -2550 7660 -2520
rect 7620 -2555 7660 -2550
rect 7620 -2585 7660 -2580
rect 7620 -2615 7625 -2585
rect 7625 -2615 7655 -2585
rect 7655 -2615 7660 -2585
rect 7620 -2620 7660 -2615
rect 7620 -2655 7660 -2650
rect 7620 -2685 7625 -2655
rect 7625 -2685 7655 -2655
rect 7655 -2685 7660 -2655
rect 7620 -2690 7660 -2685
rect 7620 -2725 7660 -2720
rect 7620 -2755 7625 -2725
rect 7625 -2755 7655 -2725
rect 7655 -2755 7660 -2725
rect 7620 -2760 7660 -2755
rect 7620 -2795 7660 -2790
rect 7620 -2825 7625 -2795
rect 7625 -2825 7655 -2795
rect 7655 -2825 7660 -2795
rect 7620 -2830 7660 -2825
rect 7620 -2860 7660 -2855
rect 7620 -2890 7625 -2860
rect 7625 -2890 7655 -2860
rect 7655 -2890 7660 -2860
rect 7620 -2895 7660 -2890
rect 7970 -1320 8010 -1315
rect 7970 -1350 7975 -1320
rect 7975 -1350 8005 -1320
rect 8005 -1350 8010 -1320
rect 7970 -1355 8010 -1350
rect 7970 -1385 8010 -1380
rect 7970 -1415 7975 -1385
rect 7975 -1415 8005 -1385
rect 8005 -1415 8010 -1385
rect 7970 -1420 8010 -1415
rect 7970 -1455 8010 -1450
rect 7970 -1485 7975 -1455
rect 7975 -1485 8005 -1455
rect 8005 -1485 8010 -1455
rect 7970 -1490 8010 -1485
rect 7970 -1525 8010 -1520
rect 7970 -1555 7975 -1525
rect 7975 -1555 8005 -1525
rect 8005 -1555 8010 -1525
rect 7970 -1560 8010 -1555
rect 7970 -1595 8010 -1590
rect 7970 -1625 7975 -1595
rect 7975 -1625 8005 -1595
rect 8005 -1625 8010 -1595
rect 7970 -1630 8010 -1625
rect 7970 -1660 8010 -1655
rect 7970 -1690 7975 -1660
rect 7975 -1690 8005 -1660
rect 8005 -1690 8010 -1660
rect 7970 -1695 8010 -1690
rect 7970 -1720 8010 -1715
rect 7970 -1750 7975 -1720
rect 7975 -1750 8005 -1720
rect 8005 -1750 8010 -1720
rect 7970 -1755 8010 -1750
rect 7970 -1785 8010 -1780
rect 7970 -1815 7975 -1785
rect 7975 -1815 8005 -1785
rect 8005 -1815 8010 -1785
rect 7970 -1820 8010 -1815
rect 7970 -1855 8010 -1850
rect 7970 -1885 7975 -1855
rect 7975 -1885 8005 -1855
rect 8005 -1885 8010 -1855
rect 7970 -1890 8010 -1885
rect 7970 -1925 8010 -1920
rect 7970 -1955 7975 -1925
rect 7975 -1955 8005 -1925
rect 8005 -1955 8010 -1925
rect 7970 -1960 8010 -1955
rect 7970 -1995 8010 -1990
rect 7970 -2025 7975 -1995
rect 7975 -2025 8005 -1995
rect 8005 -2025 8010 -1995
rect 7970 -2030 8010 -2025
rect 7970 -2060 8010 -2055
rect 7970 -2090 7975 -2060
rect 7975 -2090 8005 -2060
rect 8005 -2090 8010 -2060
rect 7970 -2095 8010 -2090
rect 7970 -2120 8010 -2115
rect 7970 -2150 7975 -2120
rect 7975 -2150 8005 -2120
rect 8005 -2150 8010 -2120
rect 7970 -2155 8010 -2150
rect 7970 -2185 8010 -2180
rect 7970 -2215 7975 -2185
rect 7975 -2215 8005 -2185
rect 8005 -2215 8010 -2185
rect 7970 -2220 8010 -2215
rect 7970 -2255 8010 -2250
rect 7970 -2285 7975 -2255
rect 7975 -2285 8005 -2255
rect 8005 -2285 8010 -2255
rect 7970 -2290 8010 -2285
rect 7970 -2325 8010 -2320
rect 7970 -2355 7975 -2325
rect 7975 -2355 8005 -2325
rect 8005 -2355 8010 -2325
rect 7970 -2360 8010 -2355
rect 7970 -2395 8010 -2390
rect 7970 -2425 7975 -2395
rect 7975 -2425 8005 -2395
rect 8005 -2425 8010 -2395
rect 7970 -2430 8010 -2425
rect 7970 -2460 8010 -2455
rect 7970 -2490 7975 -2460
rect 7975 -2490 8005 -2460
rect 8005 -2490 8010 -2460
rect 7970 -2495 8010 -2490
rect 7970 -2520 8010 -2515
rect 7970 -2550 7975 -2520
rect 7975 -2550 8005 -2520
rect 8005 -2550 8010 -2520
rect 7970 -2555 8010 -2550
rect 7970 -2585 8010 -2580
rect 7970 -2615 7975 -2585
rect 7975 -2615 8005 -2585
rect 8005 -2615 8010 -2585
rect 7970 -2620 8010 -2615
rect 7970 -2655 8010 -2650
rect 7970 -2685 7975 -2655
rect 7975 -2685 8005 -2655
rect 8005 -2685 8010 -2655
rect 7970 -2690 8010 -2685
rect 7970 -2725 8010 -2720
rect 7970 -2755 7975 -2725
rect 7975 -2755 8005 -2725
rect 8005 -2755 8010 -2725
rect 7970 -2760 8010 -2755
rect 7970 -2795 8010 -2790
rect 7970 -2825 7975 -2795
rect 7975 -2825 8005 -2795
rect 8005 -2825 8010 -2795
rect 7970 -2830 8010 -2825
rect 7970 -2860 8010 -2855
rect 7970 -2890 7975 -2860
rect 7975 -2890 8005 -2860
rect 8005 -2890 8010 -2860
rect 7970 -2895 8010 -2890
rect 8320 -1320 8360 -1315
rect 8320 -1350 8325 -1320
rect 8325 -1350 8355 -1320
rect 8355 -1350 8360 -1320
rect 8320 -1355 8360 -1350
rect 8320 -1385 8360 -1380
rect 8320 -1415 8325 -1385
rect 8325 -1415 8355 -1385
rect 8355 -1415 8360 -1385
rect 8320 -1420 8360 -1415
rect 8320 -1455 8360 -1450
rect 8320 -1485 8325 -1455
rect 8325 -1485 8355 -1455
rect 8355 -1485 8360 -1455
rect 8320 -1490 8360 -1485
rect 8320 -1525 8360 -1520
rect 8320 -1555 8325 -1525
rect 8325 -1555 8355 -1525
rect 8355 -1555 8360 -1525
rect 8320 -1560 8360 -1555
rect 8320 -1595 8360 -1590
rect 8320 -1625 8325 -1595
rect 8325 -1625 8355 -1595
rect 8355 -1625 8360 -1595
rect 8320 -1630 8360 -1625
rect 8320 -1660 8360 -1655
rect 8320 -1690 8325 -1660
rect 8325 -1690 8355 -1660
rect 8355 -1690 8360 -1660
rect 8320 -1695 8360 -1690
rect 8320 -1720 8360 -1715
rect 8320 -1750 8325 -1720
rect 8325 -1750 8355 -1720
rect 8355 -1750 8360 -1720
rect 8320 -1755 8360 -1750
rect 8320 -1785 8360 -1780
rect 8320 -1815 8325 -1785
rect 8325 -1815 8355 -1785
rect 8355 -1815 8360 -1785
rect 8320 -1820 8360 -1815
rect 8320 -1855 8360 -1850
rect 8320 -1885 8325 -1855
rect 8325 -1885 8355 -1855
rect 8355 -1885 8360 -1855
rect 8320 -1890 8360 -1885
rect 8320 -1925 8360 -1920
rect 8320 -1955 8325 -1925
rect 8325 -1955 8355 -1925
rect 8355 -1955 8360 -1925
rect 8320 -1960 8360 -1955
rect 8320 -1995 8360 -1990
rect 8320 -2025 8325 -1995
rect 8325 -2025 8355 -1995
rect 8355 -2025 8360 -1995
rect 8320 -2030 8360 -2025
rect 8320 -2060 8360 -2055
rect 8320 -2090 8325 -2060
rect 8325 -2090 8355 -2060
rect 8355 -2090 8360 -2060
rect 8320 -2095 8360 -2090
rect 8320 -2120 8360 -2115
rect 8320 -2150 8325 -2120
rect 8325 -2150 8355 -2120
rect 8355 -2150 8360 -2120
rect 8320 -2155 8360 -2150
rect 8320 -2185 8360 -2180
rect 8320 -2215 8325 -2185
rect 8325 -2215 8355 -2185
rect 8355 -2215 8360 -2185
rect 8320 -2220 8360 -2215
rect 8320 -2255 8360 -2250
rect 8320 -2285 8325 -2255
rect 8325 -2285 8355 -2255
rect 8355 -2285 8360 -2255
rect 8320 -2290 8360 -2285
rect 8320 -2325 8360 -2320
rect 8320 -2355 8325 -2325
rect 8325 -2355 8355 -2325
rect 8355 -2355 8360 -2325
rect 8320 -2360 8360 -2355
rect 8320 -2395 8360 -2390
rect 8320 -2425 8325 -2395
rect 8325 -2425 8355 -2395
rect 8355 -2425 8360 -2395
rect 8320 -2430 8360 -2425
rect 8320 -2460 8360 -2455
rect 8320 -2490 8325 -2460
rect 8325 -2490 8355 -2460
rect 8355 -2490 8360 -2460
rect 8320 -2495 8360 -2490
rect 8320 -2520 8360 -2515
rect 8320 -2550 8325 -2520
rect 8325 -2550 8355 -2520
rect 8355 -2550 8360 -2520
rect 8320 -2555 8360 -2550
rect 8320 -2585 8360 -2580
rect 8320 -2615 8325 -2585
rect 8325 -2615 8355 -2585
rect 8355 -2615 8360 -2585
rect 8320 -2620 8360 -2615
rect 8320 -2655 8360 -2650
rect 8320 -2685 8325 -2655
rect 8325 -2685 8355 -2655
rect 8355 -2685 8360 -2655
rect 8320 -2690 8360 -2685
rect 8320 -2725 8360 -2720
rect 8320 -2755 8325 -2725
rect 8325 -2755 8355 -2725
rect 8355 -2755 8360 -2725
rect 8320 -2760 8360 -2755
rect 8320 -2795 8360 -2790
rect 8320 -2825 8325 -2795
rect 8325 -2825 8355 -2795
rect 8355 -2825 8360 -2795
rect 8320 -2830 8360 -2825
rect 8320 -2860 8360 -2855
rect 8320 -2890 8325 -2860
rect 8325 -2890 8355 -2860
rect 8355 -2890 8360 -2860
rect 8320 -2895 8360 -2890
rect 8670 -1320 8710 -1315
rect 8670 -1350 8675 -1320
rect 8675 -1350 8705 -1320
rect 8705 -1350 8710 -1320
rect 8670 -1355 8710 -1350
rect 8670 -1385 8710 -1380
rect 8670 -1415 8675 -1385
rect 8675 -1415 8705 -1385
rect 8705 -1415 8710 -1385
rect 8670 -1420 8710 -1415
rect 8670 -1455 8710 -1450
rect 8670 -1485 8675 -1455
rect 8675 -1485 8705 -1455
rect 8705 -1485 8710 -1455
rect 8670 -1490 8710 -1485
rect 8670 -1525 8710 -1520
rect 8670 -1555 8675 -1525
rect 8675 -1555 8705 -1525
rect 8705 -1555 8710 -1525
rect 8670 -1560 8710 -1555
rect 8670 -1595 8710 -1590
rect 8670 -1625 8675 -1595
rect 8675 -1625 8705 -1595
rect 8705 -1625 8710 -1595
rect 8670 -1630 8710 -1625
rect 8670 -1660 8710 -1655
rect 8670 -1690 8675 -1660
rect 8675 -1690 8705 -1660
rect 8705 -1690 8710 -1660
rect 8670 -1695 8710 -1690
rect 8670 -1720 8710 -1715
rect 8670 -1750 8675 -1720
rect 8675 -1750 8705 -1720
rect 8705 -1750 8710 -1720
rect 8670 -1755 8710 -1750
rect 8670 -1785 8710 -1780
rect 8670 -1815 8675 -1785
rect 8675 -1815 8705 -1785
rect 8705 -1815 8710 -1785
rect 8670 -1820 8710 -1815
rect 8670 -1855 8710 -1850
rect 8670 -1885 8675 -1855
rect 8675 -1885 8705 -1855
rect 8705 -1885 8710 -1855
rect 8670 -1890 8710 -1885
rect 8670 -1925 8710 -1920
rect 8670 -1955 8675 -1925
rect 8675 -1955 8705 -1925
rect 8705 -1955 8710 -1925
rect 8670 -1960 8710 -1955
rect 8670 -1995 8710 -1990
rect 8670 -2025 8675 -1995
rect 8675 -2025 8705 -1995
rect 8705 -2025 8710 -1995
rect 8670 -2030 8710 -2025
rect 8670 -2060 8710 -2055
rect 8670 -2090 8675 -2060
rect 8675 -2090 8705 -2060
rect 8705 -2090 8710 -2060
rect 8670 -2095 8710 -2090
rect 8670 -2120 8710 -2115
rect 8670 -2150 8675 -2120
rect 8675 -2150 8705 -2120
rect 8705 -2150 8710 -2120
rect 8670 -2155 8710 -2150
rect 8670 -2185 8710 -2180
rect 8670 -2215 8675 -2185
rect 8675 -2215 8705 -2185
rect 8705 -2215 8710 -2185
rect 8670 -2220 8710 -2215
rect 8670 -2255 8710 -2250
rect 8670 -2285 8675 -2255
rect 8675 -2285 8705 -2255
rect 8705 -2285 8710 -2255
rect 8670 -2290 8710 -2285
rect 8670 -2325 8710 -2320
rect 8670 -2355 8675 -2325
rect 8675 -2355 8705 -2325
rect 8705 -2355 8710 -2325
rect 8670 -2360 8710 -2355
rect 8670 -2395 8710 -2390
rect 8670 -2425 8675 -2395
rect 8675 -2425 8705 -2395
rect 8705 -2425 8710 -2395
rect 8670 -2430 8710 -2425
rect 8670 -2460 8710 -2455
rect 8670 -2490 8675 -2460
rect 8675 -2490 8705 -2460
rect 8705 -2490 8710 -2460
rect 8670 -2495 8710 -2490
rect 8670 -2520 8710 -2515
rect 8670 -2550 8675 -2520
rect 8675 -2550 8705 -2520
rect 8705 -2550 8710 -2520
rect 8670 -2555 8710 -2550
rect 8670 -2585 8710 -2580
rect 8670 -2615 8675 -2585
rect 8675 -2615 8705 -2585
rect 8705 -2615 8710 -2585
rect 8670 -2620 8710 -2615
rect 8670 -2655 8710 -2650
rect 8670 -2685 8675 -2655
rect 8675 -2685 8705 -2655
rect 8705 -2685 8710 -2655
rect 8670 -2690 8710 -2685
rect 8670 -2725 8710 -2720
rect 8670 -2755 8675 -2725
rect 8675 -2755 8705 -2725
rect 8705 -2755 8710 -2725
rect 8670 -2760 8710 -2755
rect 8670 -2795 8710 -2790
rect 8670 -2825 8675 -2795
rect 8675 -2825 8705 -2795
rect 8705 -2825 8710 -2795
rect 8670 -2830 8710 -2825
rect 8670 -2860 8710 -2855
rect 8670 -2890 8675 -2860
rect 8675 -2890 8705 -2860
rect 8705 -2890 8710 -2860
rect 8670 -2895 8710 -2890
rect 9020 -1320 9060 -1315
rect 9020 -1350 9025 -1320
rect 9025 -1350 9055 -1320
rect 9055 -1350 9060 -1320
rect 9020 -1355 9060 -1350
rect 9020 -1385 9060 -1380
rect 9020 -1415 9025 -1385
rect 9025 -1415 9055 -1385
rect 9055 -1415 9060 -1385
rect 9020 -1420 9060 -1415
rect 9020 -1455 9060 -1450
rect 9020 -1485 9025 -1455
rect 9025 -1485 9055 -1455
rect 9055 -1485 9060 -1455
rect 9020 -1490 9060 -1485
rect 9020 -1525 9060 -1520
rect 9020 -1555 9025 -1525
rect 9025 -1555 9055 -1525
rect 9055 -1555 9060 -1525
rect 9020 -1560 9060 -1555
rect 9020 -1595 9060 -1590
rect 9020 -1625 9025 -1595
rect 9025 -1625 9055 -1595
rect 9055 -1625 9060 -1595
rect 9020 -1630 9060 -1625
rect 9020 -1660 9060 -1655
rect 9020 -1690 9025 -1660
rect 9025 -1690 9055 -1660
rect 9055 -1690 9060 -1660
rect 9020 -1695 9060 -1690
rect 9020 -1720 9060 -1715
rect 9020 -1750 9025 -1720
rect 9025 -1750 9055 -1720
rect 9055 -1750 9060 -1720
rect 9020 -1755 9060 -1750
rect 9020 -1785 9060 -1780
rect 9020 -1815 9025 -1785
rect 9025 -1815 9055 -1785
rect 9055 -1815 9060 -1785
rect 9020 -1820 9060 -1815
rect 9020 -1855 9060 -1850
rect 9020 -1885 9025 -1855
rect 9025 -1885 9055 -1855
rect 9055 -1885 9060 -1855
rect 9020 -1890 9060 -1885
rect 9020 -1925 9060 -1920
rect 9020 -1955 9025 -1925
rect 9025 -1955 9055 -1925
rect 9055 -1955 9060 -1925
rect 9020 -1960 9060 -1955
rect 9020 -1995 9060 -1990
rect 9020 -2025 9025 -1995
rect 9025 -2025 9055 -1995
rect 9055 -2025 9060 -1995
rect 9020 -2030 9060 -2025
rect 9020 -2060 9060 -2055
rect 9020 -2090 9025 -2060
rect 9025 -2090 9055 -2060
rect 9055 -2090 9060 -2060
rect 9020 -2095 9060 -2090
rect 9020 -2120 9060 -2115
rect 9020 -2150 9025 -2120
rect 9025 -2150 9055 -2120
rect 9055 -2150 9060 -2120
rect 9020 -2155 9060 -2150
rect 9020 -2185 9060 -2180
rect 9020 -2215 9025 -2185
rect 9025 -2215 9055 -2185
rect 9055 -2215 9060 -2185
rect 9020 -2220 9060 -2215
rect 9020 -2255 9060 -2250
rect 9020 -2285 9025 -2255
rect 9025 -2285 9055 -2255
rect 9055 -2285 9060 -2255
rect 9020 -2290 9060 -2285
rect 9020 -2325 9060 -2320
rect 9020 -2355 9025 -2325
rect 9025 -2355 9055 -2325
rect 9055 -2355 9060 -2325
rect 9020 -2360 9060 -2355
rect 9020 -2395 9060 -2390
rect 9020 -2425 9025 -2395
rect 9025 -2425 9055 -2395
rect 9055 -2425 9060 -2395
rect 9020 -2430 9060 -2425
rect 9020 -2460 9060 -2455
rect 9020 -2490 9025 -2460
rect 9025 -2490 9055 -2460
rect 9055 -2490 9060 -2460
rect 9020 -2495 9060 -2490
rect 9020 -2520 9060 -2515
rect 9020 -2550 9025 -2520
rect 9025 -2550 9055 -2520
rect 9055 -2550 9060 -2520
rect 9020 -2555 9060 -2550
rect 9020 -2585 9060 -2580
rect 9020 -2615 9025 -2585
rect 9025 -2615 9055 -2585
rect 9055 -2615 9060 -2585
rect 9020 -2620 9060 -2615
rect 9020 -2655 9060 -2650
rect 9020 -2685 9025 -2655
rect 9025 -2685 9055 -2655
rect 9055 -2685 9060 -2655
rect 9020 -2690 9060 -2685
rect 9020 -2725 9060 -2720
rect 9020 -2755 9025 -2725
rect 9025 -2755 9055 -2725
rect 9055 -2755 9060 -2725
rect 9020 -2760 9060 -2755
rect 9020 -2795 9060 -2790
rect 9020 -2825 9025 -2795
rect 9025 -2825 9055 -2795
rect 9055 -2825 9060 -2795
rect 9020 -2830 9060 -2825
rect 9020 -2860 9060 -2855
rect 9020 -2890 9025 -2860
rect 9025 -2890 9055 -2860
rect 9055 -2890 9060 -2860
rect 9020 -2895 9060 -2890
rect 31305 -1360 31340 -1325
rect 31350 -1360 31385 -1325
rect 31395 -1360 31430 -1325
rect 31440 -1360 31475 -1325
rect 31485 -1360 31520 -1325
rect 31530 -1360 31565 -1325
rect 31575 -1360 31610 -1325
rect 31620 -1360 31655 -1325
rect 31665 -1360 31700 -1325
rect 31710 -1360 31745 -1325
rect 31755 -1360 31790 -1325
rect 31800 -1360 31835 -1325
rect 31845 -1360 31880 -1325
rect 31890 -1360 31925 -1325
rect 31935 -1360 31970 -1325
rect 31980 -1360 32015 -1325
rect 32025 -1360 32060 -1325
rect 32070 -1360 32105 -1325
rect 32115 -1360 32150 -1325
rect 32160 -1360 32195 -1325
rect 32205 -1360 32240 -1325
rect 32250 -1360 32285 -1325
rect 32295 -1360 32330 -1325
rect 32340 -1360 32375 -1325
rect 32385 -1360 32420 -1325
rect 32430 -1360 32465 -1325
rect 32475 -1360 32510 -1325
rect 32520 -1360 32555 -1325
rect 32565 -1360 32600 -1325
rect 32610 -1360 32645 -1325
rect 32655 -1360 32690 -1325
rect 32700 -1360 32735 -1325
rect 32745 -1360 32780 -1325
rect 32790 -1360 32825 -1325
rect 32835 -1360 32870 -1325
rect 31305 -1405 31340 -1370
rect 31350 -1405 31385 -1370
rect 31395 -1405 31430 -1370
rect 31440 -1405 31475 -1370
rect 31485 -1405 31520 -1370
rect 31530 -1405 31565 -1370
rect 31575 -1405 31610 -1370
rect 31620 -1405 31655 -1370
rect 31665 -1405 31700 -1370
rect 31710 -1405 31745 -1370
rect 31755 -1405 31790 -1370
rect 31800 -1405 31835 -1370
rect 31845 -1405 31880 -1370
rect 31890 -1405 31925 -1370
rect 31935 -1405 31970 -1370
rect 31980 -1405 32015 -1370
rect 32025 -1405 32060 -1370
rect 32070 -1405 32105 -1370
rect 32115 -1405 32150 -1370
rect 32160 -1405 32195 -1370
rect 32205 -1405 32240 -1370
rect 32250 -1405 32285 -1370
rect 32295 -1405 32330 -1370
rect 32340 -1405 32375 -1370
rect 32385 -1405 32420 -1370
rect 32430 -1405 32465 -1370
rect 32475 -1405 32510 -1370
rect 32520 -1405 32555 -1370
rect 32565 -1405 32600 -1370
rect 32610 -1405 32645 -1370
rect 32655 -1405 32690 -1370
rect 32700 -1405 32735 -1370
rect 32745 -1405 32780 -1370
rect 32790 -1405 32825 -1370
rect 32835 -1405 32870 -1370
rect 31305 -1450 31340 -1415
rect 31350 -1450 31385 -1415
rect 31395 -1450 31430 -1415
rect 31440 -1450 31475 -1415
rect 31485 -1450 31520 -1415
rect 31530 -1450 31565 -1415
rect 31575 -1450 31610 -1415
rect 31620 -1450 31655 -1415
rect 31665 -1450 31700 -1415
rect 31710 -1450 31745 -1415
rect 31755 -1450 31790 -1415
rect 31800 -1450 31835 -1415
rect 31845 -1450 31880 -1415
rect 31890 -1450 31925 -1415
rect 31935 -1450 31970 -1415
rect 31980 -1450 32015 -1415
rect 32025 -1450 32060 -1415
rect 32070 -1450 32105 -1415
rect 32115 -1450 32150 -1415
rect 32160 -1450 32195 -1415
rect 32205 -1450 32240 -1415
rect 32250 -1450 32285 -1415
rect 32295 -1450 32330 -1415
rect 32340 -1450 32375 -1415
rect 32385 -1450 32420 -1415
rect 32430 -1450 32465 -1415
rect 32475 -1450 32510 -1415
rect 32520 -1450 32555 -1415
rect 32565 -1450 32600 -1415
rect 32610 -1450 32645 -1415
rect 32655 -1450 32690 -1415
rect 32700 -1450 32735 -1415
rect 32745 -1450 32780 -1415
rect 32790 -1450 32825 -1415
rect 32835 -1450 32870 -1415
rect 31305 -1495 31340 -1460
rect 31350 -1495 31385 -1460
rect 31395 -1495 31430 -1460
rect 31440 -1495 31475 -1460
rect 31485 -1495 31520 -1460
rect 31530 -1495 31565 -1460
rect 31575 -1495 31610 -1460
rect 31620 -1495 31655 -1460
rect 31665 -1495 31700 -1460
rect 31710 -1495 31745 -1460
rect 31755 -1495 31790 -1460
rect 31800 -1495 31835 -1460
rect 31845 -1495 31880 -1460
rect 31890 -1495 31925 -1460
rect 31935 -1495 31970 -1460
rect 31980 -1495 32015 -1460
rect 32025 -1495 32060 -1460
rect 32070 -1495 32105 -1460
rect 32115 -1495 32150 -1460
rect 32160 -1495 32195 -1460
rect 32205 -1495 32240 -1460
rect 32250 -1495 32285 -1460
rect 32295 -1495 32330 -1460
rect 32340 -1495 32375 -1460
rect 32385 -1495 32420 -1460
rect 32430 -1495 32465 -1460
rect 32475 -1495 32510 -1460
rect 32520 -1495 32555 -1460
rect 32565 -1495 32600 -1460
rect 32610 -1495 32645 -1460
rect 32655 -1495 32690 -1460
rect 32700 -1495 32735 -1460
rect 32745 -1495 32780 -1460
rect 32790 -1495 32825 -1460
rect 32835 -1495 32870 -1460
rect 31305 -1540 31340 -1505
rect 31350 -1540 31385 -1505
rect 31395 -1540 31430 -1505
rect 31440 -1540 31475 -1505
rect 31485 -1540 31520 -1505
rect 31530 -1540 31565 -1505
rect 31575 -1540 31610 -1505
rect 31620 -1540 31655 -1505
rect 31665 -1540 31700 -1505
rect 31710 -1540 31745 -1505
rect 31755 -1540 31790 -1505
rect 31800 -1540 31835 -1505
rect 31845 -1540 31880 -1505
rect 31890 -1540 31925 -1505
rect 31935 -1540 31970 -1505
rect 31980 -1540 32015 -1505
rect 32025 -1540 32060 -1505
rect 32070 -1540 32105 -1505
rect 32115 -1540 32150 -1505
rect 32160 -1540 32195 -1505
rect 32205 -1540 32240 -1505
rect 32250 -1540 32285 -1505
rect 32295 -1540 32330 -1505
rect 32340 -1540 32375 -1505
rect 32385 -1540 32420 -1505
rect 32430 -1540 32465 -1505
rect 32475 -1540 32510 -1505
rect 32520 -1540 32555 -1505
rect 32565 -1540 32600 -1505
rect 32610 -1540 32645 -1505
rect 32655 -1540 32690 -1505
rect 32700 -1540 32735 -1505
rect 32745 -1540 32780 -1505
rect 32790 -1540 32825 -1505
rect 32835 -1540 32870 -1505
rect 31305 -1585 31340 -1550
rect 31350 -1585 31385 -1550
rect 31395 -1585 31430 -1550
rect 31440 -1585 31475 -1550
rect 31485 -1585 31520 -1550
rect 31530 -1585 31565 -1550
rect 31575 -1585 31610 -1550
rect 31620 -1585 31655 -1550
rect 31665 -1585 31700 -1550
rect 31710 -1585 31745 -1550
rect 31755 -1585 31790 -1550
rect 31800 -1585 31835 -1550
rect 31845 -1585 31880 -1550
rect 31890 -1585 31925 -1550
rect 31935 -1585 31970 -1550
rect 31980 -1585 32015 -1550
rect 32025 -1585 32060 -1550
rect 32070 -1585 32105 -1550
rect 32115 -1585 32150 -1550
rect 32160 -1585 32195 -1550
rect 32205 -1585 32240 -1550
rect 32250 -1585 32285 -1550
rect 32295 -1585 32330 -1550
rect 32340 -1585 32375 -1550
rect 32385 -1585 32420 -1550
rect 32430 -1585 32465 -1550
rect 32475 -1585 32510 -1550
rect 32520 -1585 32555 -1550
rect 32565 -1585 32600 -1550
rect 32610 -1585 32645 -1550
rect 32655 -1585 32690 -1550
rect 32700 -1585 32735 -1550
rect 32745 -1585 32780 -1550
rect 32790 -1585 32825 -1550
rect 32835 -1585 32870 -1550
rect 31305 -1630 31340 -1595
rect 31350 -1630 31385 -1595
rect 31395 -1630 31430 -1595
rect 31440 -1630 31475 -1595
rect 31485 -1630 31520 -1595
rect 31530 -1630 31565 -1595
rect 31575 -1630 31610 -1595
rect 31620 -1630 31655 -1595
rect 31665 -1630 31700 -1595
rect 31710 -1630 31745 -1595
rect 31755 -1630 31790 -1595
rect 31800 -1630 31835 -1595
rect 31845 -1630 31880 -1595
rect 31890 -1630 31925 -1595
rect 31935 -1630 31970 -1595
rect 31980 -1630 32015 -1595
rect 32025 -1630 32060 -1595
rect 32070 -1630 32105 -1595
rect 32115 -1630 32150 -1595
rect 32160 -1630 32195 -1595
rect 32205 -1630 32240 -1595
rect 32250 -1630 32285 -1595
rect 32295 -1630 32330 -1595
rect 32340 -1630 32375 -1595
rect 32385 -1630 32420 -1595
rect 32430 -1630 32465 -1595
rect 32475 -1630 32510 -1595
rect 32520 -1630 32555 -1595
rect 32565 -1630 32600 -1595
rect 32610 -1630 32645 -1595
rect 32655 -1630 32690 -1595
rect 32700 -1630 32735 -1595
rect 32745 -1630 32780 -1595
rect 32790 -1630 32825 -1595
rect 32835 -1630 32870 -1595
rect 31305 -1675 31340 -1640
rect 31350 -1675 31385 -1640
rect 31395 -1675 31430 -1640
rect 31440 -1675 31475 -1640
rect 31485 -1675 31520 -1640
rect 31530 -1675 31565 -1640
rect 31575 -1675 31610 -1640
rect 31620 -1675 31655 -1640
rect 31665 -1675 31700 -1640
rect 31710 -1675 31745 -1640
rect 31755 -1675 31790 -1640
rect 31800 -1675 31835 -1640
rect 31845 -1675 31880 -1640
rect 31890 -1675 31925 -1640
rect 31935 -1675 31970 -1640
rect 31980 -1675 32015 -1640
rect 32025 -1675 32060 -1640
rect 32070 -1675 32105 -1640
rect 32115 -1675 32150 -1640
rect 32160 -1675 32195 -1640
rect 32205 -1675 32240 -1640
rect 32250 -1675 32285 -1640
rect 32295 -1675 32330 -1640
rect 32340 -1675 32375 -1640
rect 32385 -1675 32420 -1640
rect 32430 -1675 32465 -1640
rect 32475 -1675 32510 -1640
rect 32520 -1675 32555 -1640
rect 32565 -1675 32600 -1640
rect 32610 -1675 32645 -1640
rect 32655 -1675 32690 -1640
rect 32700 -1675 32735 -1640
rect 32745 -1675 32780 -1640
rect 32790 -1675 32825 -1640
rect 32835 -1675 32870 -1640
rect 31305 -1720 31340 -1685
rect 31350 -1720 31385 -1685
rect 31395 -1720 31430 -1685
rect 31440 -1720 31475 -1685
rect 31485 -1720 31520 -1685
rect 31530 -1720 31565 -1685
rect 31575 -1720 31610 -1685
rect 31620 -1720 31655 -1685
rect 31665 -1720 31700 -1685
rect 31710 -1720 31745 -1685
rect 31755 -1720 31790 -1685
rect 31800 -1720 31835 -1685
rect 31845 -1720 31880 -1685
rect 31890 -1720 31925 -1685
rect 31935 -1720 31970 -1685
rect 31980 -1720 32015 -1685
rect 32025 -1720 32060 -1685
rect 32070 -1720 32105 -1685
rect 32115 -1720 32150 -1685
rect 32160 -1720 32195 -1685
rect 32205 -1720 32240 -1685
rect 32250 -1720 32285 -1685
rect 32295 -1720 32330 -1685
rect 32340 -1720 32375 -1685
rect 32385 -1720 32420 -1685
rect 32430 -1720 32465 -1685
rect 32475 -1720 32510 -1685
rect 32520 -1720 32555 -1685
rect 32565 -1720 32600 -1685
rect 32610 -1720 32645 -1685
rect 32655 -1720 32690 -1685
rect 32700 -1720 32735 -1685
rect 32745 -1720 32780 -1685
rect 32790 -1720 32825 -1685
rect 32835 -1720 32870 -1685
rect 31305 -1765 31340 -1730
rect 31350 -1765 31385 -1730
rect 31395 -1765 31430 -1730
rect 31440 -1765 31475 -1730
rect 31485 -1765 31520 -1730
rect 31530 -1765 31565 -1730
rect 31575 -1765 31610 -1730
rect 31620 -1765 31655 -1730
rect 31665 -1765 31700 -1730
rect 31710 -1765 31745 -1730
rect 31755 -1765 31790 -1730
rect 31800 -1765 31835 -1730
rect 31845 -1765 31880 -1730
rect 31890 -1765 31925 -1730
rect 31935 -1765 31970 -1730
rect 31980 -1765 32015 -1730
rect 32025 -1765 32060 -1730
rect 32070 -1765 32105 -1730
rect 32115 -1765 32150 -1730
rect 32160 -1765 32195 -1730
rect 32205 -1765 32240 -1730
rect 32250 -1765 32285 -1730
rect 32295 -1765 32330 -1730
rect 32340 -1765 32375 -1730
rect 32385 -1765 32420 -1730
rect 32430 -1765 32465 -1730
rect 32475 -1765 32510 -1730
rect 32520 -1765 32555 -1730
rect 32565 -1765 32600 -1730
rect 32610 -1765 32645 -1730
rect 32655 -1765 32690 -1730
rect 32700 -1765 32735 -1730
rect 32745 -1765 32780 -1730
rect 32790 -1765 32825 -1730
rect 32835 -1765 32870 -1730
rect 31305 -1810 31340 -1775
rect 31350 -1810 31385 -1775
rect 31395 -1810 31430 -1775
rect 31440 -1810 31475 -1775
rect 31485 -1810 31520 -1775
rect 31530 -1810 31565 -1775
rect 31575 -1810 31610 -1775
rect 31620 -1810 31655 -1775
rect 31665 -1810 31700 -1775
rect 31710 -1810 31745 -1775
rect 31755 -1810 31790 -1775
rect 31800 -1810 31835 -1775
rect 31845 -1810 31880 -1775
rect 31890 -1810 31925 -1775
rect 31935 -1810 31970 -1775
rect 31980 -1810 32015 -1775
rect 32025 -1810 32060 -1775
rect 32070 -1810 32105 -1775
rect 32115 -1810 32150 -1775
rect 32160 -1810 32195 -1775
rect 32205 -1810 32240 -1775
rect 32250 -1810 32285 -1775
rect 32295 -1810 32330 -1775
rect 32340 -1810 32375 -1775
rect 32385 -1810 32420 -1775
rect 32430 -1810 32465 -1775
rect 32475 -1810 32510 -1775
rect 32520 -1810 32555 -1775
rect 32565 -1810 32600 -1775
rect 32610 -1810 32645 -1775
rect 32655 -1810 32690 -1775
rect 32700 -1810 32735 -1775
rect 32745 -1810 32780 -1775
rect 32790 -1810 32825 -1775
rect 32835 -1810 32870 -1775
rect 31305 -1855 31340 -1820
rect 31350 -1855 31385 -1820
rect 31395 -1855 31430 -1820
rect 31440 -1855 31475 -1820
rect 31485 -1855 31520 -1820
rect 31530 -1855 31565 -1820
rect 31575 -1855 31610 -1820
rect 31620 -1855 31655 -1820
rect 31665 -1855 31700 -1820
rect 31710 -1855 31745 -1820
rect 31755 -1855 31790 -1820
rect 31800 -1855 31835 -1820
rect 31845 -1855 31880 -1820
rect 31890 -1855 31925 -1820
rect 31935 -1855 31970 -1820
rect 31980 -1855 32015 -1820
rect 32025 -1855 32060 -1820
rect 32070 -1855 32105 -1820
rect 32115 -1855 32150 -1820
rect 32160 -1855 32195 -1820
rect 32205 -1855 32240 -1820
rect 32250 -1855 32285 -1820
rect 32295 -1855 32330 -1820
rect 32340 -1855 32375 -1820
rect 32385 -1855 32420 -1820
rect 32430 -1855 32465 -1820
rect 32475 -1855 32510 -1820
rect 32520 -1855 32555 -1820
rect 32565 -1855 32600 -1820
rect 32610 -1855 32645 -1820
rect 32655 -1855 32690 -1820
rect 32700 -1855 32735 -1820
rect 32745 -1855 32780 -1820
rect 32790 -1855 32825 -1820
rect 32835 -1855 32870 -1820
rect 31305 -1900 31340 -1865
rect 31350 -1900 31385 -1865
rect 31395 -1900 31430 -1865
rect 31440 -1900 31475 -1865
rect 31485 -1900 31520 -1865
rect 31530 -1900 31565 -1865
rect 31575 -1900 31610 -1865
rect 31620 -1900 31655 -1865
rect 31665 -1900 31700 -1865
rect 31710 -1900 31745 -1865
rect 31755 -1900 31790 -1865
rect 31800 -1900 31835 -1865
rect 31845 -1900 31880 -1865
rect 31890 -1900 31925 -1865
rect 31935 -1900 31970 -1865
rect 31980 -1900 32015 -1865
rect 32025 -1900 32060 -1865
rect 32070 -1900 32105 -1865
rect 32115 -1900 32150 -1865
rect 32160 -1900 32195 -1865
rect 32205 -1900 32240 -1865
rect 32250 -1900 32285 -1865
rect 32295 -1900 32330 -1865
rect 32340 -1900 32375 -1865
rect 32385 -1900 32420 -1865
rect 32430 -1900 32465 -1865
rect 32475 -1900 32510 -1865
rect 32520 -1900 32555 -1865
rect 32565 -1900 32600 -1865
rect 32610 -1900 32645 -1865
rect 32655 -1900 32690 -1865
rect 32700 -1900 32735 -1865
rect 32745 -1900 32780 -1865
rect 32790 -1900 32825 -1865
rect 32835 -1900 32870 -1865
rect 31305 -1945 31340 -1910
rect 31350 -1945 31385 -1910
rect 31395 -1945 31430 -1910
rect 31440 -1945 31475 -1910
rect 31485 -1945 31520 -1910
rect 31530 -1945 31565 -1910
rect 31575 -1945 31610 -1910
rect 31620 -1945 31655 -1910
rect 31665 -1945 31700 -1910
rect 31710 -1945 31745 -1910
rect 31755 -1945 31790 -1910
rect 31800 -1945 31835 -1910
rect 31845 -1945 31880 -1910
rect 31890 -1945 31925 -1910
rect 31935 -1945 31970 -1910
rect 31980 -1945 32015 -1910
rect 32025 -1945 32060 -1910
rect 32070 -1945 32105 -1910
rect 32115 -1945 32150 -1910
rect 32160 -1945 32195 -1910
rect 32205 -1945 32240 -1910
rect 32250 -1945 32285 -1910
rect 32295 -1945 32330 -1910
rect 32340 -1945 32375 -1910
rect 32385 -1945 32420 -1910
rect 32430 -1945 32465 -1910
rect 32475 -1945 32510 -1910
rect 32520 -1945 32555 -1910
rect 32565 -1945 32600 -1910
rect 32610 -1945 32645 -1910
rect 32655 -1945 32690 -1910
rect 32700 -1945 32735 -1910
rect 32745 -1945 32780 -1910
rect 32790 -1945 32825 -1910
rect 32835 -1945 32870 -1910
rect 31305 -1990 31340 -1955
rect 31350 -1990 31385 -1955
rect 31395 -1990 31430 -1955
rect 31440 -1990 31475 -1955
rect 31485 -1990 31520 -1955
rect 31530 -1990 31565 -1955
rect 31575 -1990 31610 -1955
rect 31620 -1990 31655 -1955
rect 31665 -1990 31700 -1955
rect 31710 -1990 31745 -1955
rect 31755 -1990 31790 -1955
rect 31800 -1990 31835 -1955
rect 31845 -1990 31880 -1955
rect 31890 -1990 31925 -1955
rect 31935 -1990 31970 -1955
rect 31980 -1990 32015 -1955
rect 32025 -1990 32060 -1955
rect 32070 -1990 32105 -1955
rect 32115 -1990 32150 -1955
rect 32160 -1990 32195 -1955
rect 32205 -1990 32240 -1955
rect 32250 -1990 32285 -1955
rect 32295 -1990 32330 -1955
rect 32340 -1990 32375 -1955
rect 32385 -1990 32420 -1955
rect 32430 -1990 32465 -1955
rect 32475 -1990 32510 -1955
rect 32520 -1990 32555 -1955
rect 32565 -1990 32600 -1955
rect 32610 -1990 32645 -1955
rect 32655 -1990 32690 -1955
rect 32700 -1990 32735 -1955
rect 32745 -1990 32780 -1955
rect 32790 -1990 32825 -1955
rect 32835 -1990 32870 -1955
rect 31305 -2035 31340 -2000
rect 31350 -2035 31385 -2000
rect 31395 -2035 31430 -2000
rect 31440 -2035 31475 -2000
rect 31485 -2035 31520 -2000
rect 31530 -2035 31565 -2000
rect 31575 -2035 31610 -2000
rect 31620 -2035 31655 -2000
rect 31665 -2035 31700 -2000
rect 31710 -2035 31745 -2000
rect 31755 -2035 31790 -2000
rect 31800 -2035 31835 -2000
rect 31845 -2035 31880 -2000
rect 31890 -2035 31925 -2000
rect 31935 -2035 31970 -2000
rect 31980 -2035 32015 -2000
rect 32025 -2035 32060 -2000
rect 32070 -2035 32105 -2000
rect 32115 -2035 32150 -2000
rect 32160 -2035 32195 -2000
rect 32205 -2035 32240 -2000
rect 32250 -2035 32285 -2000
rect 32295 -2035 32330 -2000
rect 32340 -2035 32375 -2000
rect 32385 -2035 32420 -2000
rect 32430 -2035 32465 -2000
rect 32475 -2035 32510 -2000
rect 32520 -2035 32555 -2000
rect 32565 -2035 32600 -2000
rect 32610 -2035 32645 -2000
rect 32655 -2035 32690 -2000
rect 32700 -2035 32735 -2000
rect 32745 -2035 32780 -2000
rect 32790 -2035 32825 -2000
rect 32835 -2035 32870 -2000
rect 31305 -2080 31340 -2045
rect 31350 -2080 31385 -2045
rect 31395 -2080 31430 -2045
rect 31440 -2080 31475 -2045
rect 31485 -2080 31520 -2045
rect 31530 -2080 31565 -2045
rect 31575 -2080 31610 -2045
rect 31620 -2080 31655 -2045
rect 31665 -2080 31700 -2045
rect 31710 -2080 31745 -2045
rect 31755 -2080 31790 -2045
rect 31800 -2080 31835 -2045
rect 31845 -2080 31880 -2045
rect 31890 -2080 31925 -2045
rect 31935 -2080 31970 -2045
rect 31980 -2080 32015 -2045
rect 32025 -2080 32060 -2045
rect 32070 -2080 32105 -2045
rect 32115 -2080 32150 -2045
rect 32160 -2080 32195 -2045
rect 32205 -2080 32240 -2045
rect 32250 -2080 32285 -2045
rect 32295 -2080 32330 -2045
rect 32340 -2080 32375 -2045
rect 32385 -2080 32420 -2045
rect 32430 -2080 32465 -2045
rect 32475 -2080 32510 -2045
rect 32520 -2080 32555 -2045
rect 32565 -2080 32600 -2045
rect 32610 -2080 32645 -2045
rect 32655 -2080 32690 -2045
rect 32700 -2080 32735 -2045
rect 32745 -2080 32780 -2045
rect 32790 -2080 32825 -2045
rect 32835 -2080 32870 -2045
rect 31305 -2125 31340 -2090
rect 31350 -2125 31385 -2090
rect 31395 -2125 31430 -2090
rect 31440 -2125 31475 -2090
rect 31485 -2125 31520 -2090
rect 31530 -2125 31565 -2090
rect 31575 -2125 31610 -2090
rect 31620 -2125 31655 -2090
rect 31665 -2125 31700 -2090
rect 31710 -2125 31745 -2090
rect 31755 -2125 31790 -2090
rect 31800 -2125 31835 -2090
rect 31845 -2125 31880 -2090
rect 31890 -2125 31925 -2090
rect 31935 -2125 31970 -2090
rect 31980 -2125 32015 -2090
rect 32025 -2125 32060 -2090
rect 32070 -2125 32105 -2090
rect 32115 -2125 32150 -2090
rect 32160 -2125 32195 -2090
rect 32205 -2125 32240 -2090
rect 32250 -2125 32285 -2090
rect 32295 -2125 32330 -2090
rect 32340 -2125 32375 -2090
rect 32385 -2125 32420 -2090
rect 32430 -2125 32465 -2090
rect 32475 -2125 32510 -2090
rect 32520 -2125 32555 -2090
rect 32565 -2125 32600 -2090
rect 32610 -2125 32645 -2090
rect 32655 -2125 32690 -2090
rect 32700 -2125 32735 -2090
rect 32745 -2125 32780 -2090
rect 32790 -2125 32825 -2090
rect 32835 -2125 32870 -2090
rect 31305 -2170 31340 -2135
rect 31350 -2170 31385 -2135
rect 31395 -2170 31430 -2135
rect 31440 -2170 31475 -2135
rect 31485 -2170 31520 -2135
rect 31530 -2170 31565 -2135
rect 31575 -2170 31610 -2135
rect 31620 -2170 31655 -2135
rect 31665 -2170 31700 -2135
rect 31710 -2170 31745 -2135
rect 31755 -2170 31790 -2135
rect 31800 -2170 31835 -2135
rect 31845 -2170 31880 -2135
rect 31890 -2170 31925 -2135
rect 31935 -2170 31970 -2135
rect 31980 -2170 32015 -2135
rect 32025 -2170 32060 -2135
rect 32070 -2170 32105 -2135
rect 32115 -2170 32150 -2135
rect 32160 -2170 32195 -2135
rect 32205 -2170 32240 -2135
rect 32250 -2170 32285 -2135
rect 32295 -2170 32330 -2135
rect 32340 -2170 32375 -2135
rect 32385 -2170 32420 -2135
rect 32430 -2170 32465 -2135
rect 32475 -2170 32510 -2135
rect 32520 -2170 32555 -2135
rect 32565 -2170 32600 -2135
rect 32610 -2170 32645 -2135
rect 32655 -2170 32690 -2135
rect 32700 -2170 32735 -2135
rect 32745 -2170 32780 -2135
rect 32790 -2170 32825 -2135
rect 32835 -2170 32870 -2135
rect 31305 -2215 31340 -2180
rect 31350 -2215 31385 -2180
rect 31395 -2215 31430 -2180
rect 31440 -2215 31475 -2180
rect 31485 -2215 31520 -2180
rect 31530 -2215 31565 -2180
rect 31575 -2215 31610 -2180
rect 31620 -2215 31655 -2180
rect 31665 -2215 31700 -2180
rect 31710 -2215 31745 -2180
rect 31755 -2215 31790 -2180
rect 31800 -2215 31835 -2180
rect 31845 -2215 31880 -2180
rect 31890 -2215 31925 -2180
rect 31935 -2215 31970 -2180
rect 31980 -2215 32015 -2180
rect 32025 -2215 32060 -2180
rect 32070 -2215 32105 -2180
rect 32115 -2215 32150 -2180
rect 32160 -2215 32195 -2180
rect 32205 -2215 32240 -2180
rect 32250 -2215 32285 -2180
rect 32295 -2215 32330 -2180
rect 32340 -2215 32375 -2180
rect 32385 -2215 32420 -2180
rect 32430 -2215 32465 -2180
rect 32475 -2215 32510 -2180
rect 32520 -2215 32555 -2180
rect 32565 -2215 32600 -2180
rect 32610 -2215 32645 -2180
rect 32655 -2215 32690 -2180
rect 32700 -2215 32735 -2180
rect 32745 -2215 32780 -2180
rect 32790 -2215 32825 -2180
rect 32835 -2215 32870 -2180
rect 31305 -2260 31340 -2225
rect 31350 -2260 31385 -2225
rect 31395 -2260 31430 -2225
rect 31440 -2260 31475 -2225
rect 31485 -2260 31520 -2225
rect 31530 -2260 31565 -2225
rect 31575 -2260 31610 -2225
rect 31620 -2260 31655 -2225
rect 31665 -2260 31700 -2225
rect 31710 -2260 31745 -2225
rect 31755 -2260 31790 -2225
rect 31800 -2260 31835 -2225
rect 31845 -2260 31880 -2225
rect 31890 -2260 31925 -2225
rect 31935 -2260 31970 -2225
rect 31980 -2260 32015 -2225
rect 32025 -2260 32060 -2225
rect 32070 -2260 32105 -2225
rect 32115 -2260 32150 -2225
rect 32160 -2260 32195 -2225
rect 32205 -2260 32240 -2225
rect 32250 -2260 32285 -2225
rect 32295 -2260 32330 -2225
rect 32340 -2260 32375 -2225
rect 32385 -2260 32420 -2225
rect 32430 -2260 32465 -2225
rect 32475 -2260 32510 -2225
rect 32520 -2260 32555 -2225
rect 32565 -2260 32600 -2225
rect 32610 -2260 32645 -2225
rect 32655 -2260 32690 -2225
rect 32700 -2260 32735 -2225
rect 32745 -2260 32780 -2225
rect 32790 -2260 32825 -2225
rect 32835 -2260 32870 -2225
rect 31305 -2305 31340 -2270
rect 31350 -2305 31385 -2270
rect 31395 -2305 31430 -2270
rect 31440 -2305 31475 -2270
rect 31485 -2305 31520 -2270
rect 31530 -2305 31565 -2270
rect 31575 -2305 31610 -2270
rect 31620 -2305 31655 -2270
rect 31665 -2305 31700 -2270
rect 31710 -2305 31745 -2270
rect 31755 -2305 31790 -2270
rect 31800 -2305 31835 -2270
rect 31845 -2305 31880 -2270
rect 31890 -2305 31925 -2270
rect 31935 -2305 31970 -2270
rect 31980 -2305 32015 -2270
rect 32025 -2305 32060 -2270
rect 32070 -2305 32105 -2270
rect 32115 -2305 32150 -2270
rect 32160 -2305 32195 -2270
rect 32205 -2305 32240 -2270
rect 32250 -2305 32285 -2270
rect 32295 -2305 32330 -2270
rect 32340 -2305 32375 -2270
rect 32385 -2305 32420 -2270
rect 32430 -2305 32465 -2270
rect 32475 -2305 32510 -2270
rect 32520 -2305 32555 -2270
rect 32565 -2305 32600 -2270
rect 32610 -2305 32645 -2270
rect 32655 -2305 32690 -2270
rect 32700 -2305 32735 -2270
rect 32745 -2305 32780 -2270
rect 32790 -2305 32825 -2270
rect 32835 -2305 32870 -2270
rect 31305 -2350 31340 -2315
rect 31350 -2350 31385 -2315
rect 31395 -2350 31430 -2315
rect 31440 -2350 31475 -2315
rect 31485 -2350 31520 -2315
rect 31530 -2350 31565 -2315
rect 31575 -2350 31610 -2315
rect 31620 -2350 31655 -2315
rect 31665 -2350 31700 -2315
rect 31710 -2350 31745 -2315
rect 31755 -2350 31790 -2315
rect 31800 -2350 31835 -2315
rect 31845 -2350 31880 -2315
rect 31890 -2350 31925 -2315
rect 31935 -2350 31970 -2315
rect 31980 -2350 32015 -2315
rect 32025 -2350 32060 -2315
rect 32070 -2350 32105 -2315
rect 32115 -2350 32150 -2315
rect 32160 -2350 32195 -2315
rect 32205 -2350 32240 -2315
rect 32250 -2350 32285 -2315
rect 32295 -2350 32330 -2315
rect 32340 -2350 32375 -2315
rect 32385 -2350 32420 -2315
rect 32430 -2350 32465 -2315
rect 32475 -2350 32510 -2315
rect 32520 -2350 32555 -2315
rect 32565 -2350 32600 -2315
rect 32610 -2350 32645 -2315
rect 32655 -2350 32690 -2315
rect 32700 -2350 32735 -2315
rect 32745 -2350 32780 -2315
rect 32790 -2350 32825 -2315
rect 32835 -2350 32870 -2315
rect 31305 -2395 31340 -2360
rect 31350 -2395 31385 -2360
rect 31395 -2395 31430 -2360
rect 31440 -2395 31475 -2360
rect 31485 -2395 31520 -2360
rect 31530 -2395 31565 -2360
rect 31575 -2395 31610 -2360
rect 31620 -2395 31655 -2360
rect 31665 -2395 31700 -2360
rect 31710 -2395 31745 -2360
rect 31755 -2395 31790 -2360
rect 31800 -2395 31835 -2360
rect 31845 -2395 31880 -2360
rect 31890 -2395 31925 -2360
rect 31935 -2395 31970 -2360
rect 31980 -2395 32015 -2360
rect 32025 -2395 32060 -2360
rect 32070 -2395 32105 -2360
rect 32115 -2395 32150 -2360
rect 32160 -2395 32195 -2360
rect 32205 -2395 32240 -2360
rect 32250 -2395 32285 -2360
rect 32295 -2395 32330 -2360
rect 32340 -2395 32375 -2360
rect 32385 -2395 32420 -2360
rect 32430 -2395 32465 -2360
rect 32475 -2395 32510 -2360
rect 32520 -2395 32555 -2360
rect 32565 -2395 32600 -2360
rect 32610 -2395 32645 -2360
rect 32655 -2395 32690 -2360
rect 32700 -2395 32735 -2360
rect 32745 -2395 32780 -2360
rect 32790 -2395 32825 -2360
rect 32835 -2395 32870 -2360
rect 31305 -2440 31340 -2405
rect 31350 -2440 31385 -2405
rect 31395 -2440 31430 -2405
rect 31440 -2440 31475 -2405
rect 31485 -2440 31520 -2405
rect 31530 -2440 31565 -2405
rect 31575 -2440 31610 -2405
rect 31620 -2440 31655 -2405
rect 31665 -2440 31700 -2405
rect 31710 -2440 31745 -2405
rect 31755 -2440 31790 -2405
rect 31800 -2440 31835 -2405
rect 31845 -2440 31880 -2405
rect 31890 -2440 31925 -2405
rect 31935 -2440 31970 -2405
rect 31980 -2440 32015 -2405
rect 32025 -2440 32060 -2405
rect 32070 -2440 32105 -2405
rect 32115 -2440 32150 -2405
rect 32160 -2440 32195 -2405
rect 32205 -2440 32240 -2405
rect 32250 -2440 32285 -2405
rect 32295 -2440 32330 -2405
rect 32340 -2440 32375 -2405
rect 32385 -2440 32420 -2405
rect 32430 -2440 32465 -2405
rect 32475 -2440 32510 -2405
rect 32520 -2440 32555 -2405
rect 32565 -2440 32600 -2405
rect 32610 -2440 32645 -2405
rect 32655 -2440 32690 -2405
rect 32700 -2440 32735 -2405
rect 32745 -2440 32780 -2405
rect 32790 -2440 32825 -2405
rect 32835 -2440 32870 -2405
rect 31305 -2485 31340 -2450
rect 31350 -2485 31385 -2450
rect 31395 -2485 31430 -2450
rect 31440 -2485 31475 -2450
rect 31485 -2485 31520 -2450
rect 31530 -2485 31565 -2450
rect 31575 -2485 31610 -2450
rect 31620 -2485 31655 -2450
rect 31665 -2485 31700 -2450
rect 31710 -2485 31745 -2450
rect 31755 -2485 31790 -2450
rect 31800 -2485 31835 -2450
rect 31845 -2485 31880 -2450
rect 31890 -2485 31925 -2450
rect 31935 -2485 31970 -2450
rect 31980 -2485 32015 -2450
rect 32025 -2485 32060 -2450
rect 32070 -2485 32105 -2450
rect 32115 -2485 32150 -2450
rect 32160 -2485 32195 -2450
rect 32205 -2485 32240 -2450
rect 32250 -2485 32285 -2450
rect 32295 -2485 32330 -2450
rect 32340 -2485 32375 -2450
rect 32385 -2485 32420 -2450
rect 32430 -2485 32465 -2450
rect 32475 -2485 32510 -2450
rect 32520 -2485 32555 -2450
rect 32565 -2485 32600 -2450
rect 32610 -2485 32645 -2450
rect 32655 -2485 32690 -2450
rect 32700 -2485 32735 -2450
rect 32745 -2485 32780 -2450
rect 32790 -2485 32825 -2450
rect 32835 -2485 32870 -2450
rect 31305 -2530 31340 -2495
rect 31350 -2530 31385 -2495
rect 31395 -2530 31430 -2495
rect 31440 -2530 31475 -2495
rect 31485 -2530 31520 -2495
rect 31530 -2530 31565 -2495
rect 31575 -2530 31610 -2495
rect 31620 -2530 31655 -2495
rect 31665 -2530 31700 -2495
rect 31710 -2530 31745 -2495
rect 31755 -2530 31790 -2495
rect 31800 -2530 31835 -2495
rect 31845 -2530 31880 -2495
rect 31890 -2530 31925 -2495
rect 31935 -2530 31970 -2495
rect 31980 -2530 32015 -2495
rect 32025 -2530 32060 -2495
rect 32070 -2530 32105 -2495
rect 32115 -2530 32150 -2495
rect 32160 -2530 32195 -2495
rect 32205 -2530 32240 -2495
rect 32250 -2530 32285 -2495
rect 32295 -2530 32330 -2495
rect 32340 -2530 32375 -2495
rect 32385 -2530 32420 -2495
rect 32430 -2530 32465 -2495
rect 32475 -2530 32510 -2495
rect 32520 -2530 32555 -2495
rect 32565 -2530 32600 -2495
rect 32610 -2530 32645 -2495
rect 32655 -2530 32690 -2495
rect 32700 -2530 32735 -2495
rect 32745 -2530 32780 -2495
rect 32790 -2530 32825 -2495
rect 32835 -2530 32870 -2495
rect 31305 -2575 31340 -2540
rect 31350 -2575 31385 -2540
rect 31395 -2575 31430 -2540
rect 31440 -2575 31475 -2540
rect 31485 -2575 31520 -2540
rect 31530 -2575 31565 -2540
rect 31575 -2575 31610 -2540
rect 31620 -2575 31655 -2540
rect 31665 -2575 31700 -2540
rect 31710 -2575 31745 -2540
rect 31755 -2575 31790 -2540
rect 31800 -2575 31835 -2540
rect 31845 -2575 31880 -2540
rect 31890 -2575 31925 -2540
rect 31935 -2575 31970 -2540
rect 31980 -2575 32015 -2540
rect 32025 -2575 32060 -2540
rect 32070 -2575 32105 -2540
rect 32115 -2575 32150 -2540
rect 32160 -2575 32195 -2540
rect 32205 -2575 32240 -2540
rect 32250 -2575 32285 -2540
rect 32295 -2575 32330 -2540
rect 32340 -2575 32375 -2540
rect 32385 -2575 32420 -2540
rect 32430 -2575 32465 -2540
rect 32475 -2575 32510 -2540
rect 32520 -2575 32555 -2540
rect 32565 -2575 32600 -2540
rect 32610 -2575 32645 -2540
rect 32655 -2575 32690 -2540
rect 32700 -2575 32735 -2540
rect 32745 -2575 32780 -2540
rect 32790 -2575 32825 -2540
rect 32835 -2575 32870 -2540
rect 31305 -2620 31340 -2585
rect 31350 -2620 31385 -2585
rect 31395 -2620 31430 -2585
rect 31440 -2620 31475 -2585
rect 31485 -2620 31520 -2585
rect 31530 -2620 31565 -2585
rect 31575 -2620 31610 -2585
rect 31620 -2620 31655 -2585
rect 31665 -2620 31700 -2585
rect 31710 -2620 31745 -2585
rect 31755 -2620 31790 -2585
rect 31800 -2620 31835 -2585
rect 31845 -2620 31880 -2585
rect 31890 -2620 31925 -2585
rect 31935 -2620 31970 -2585
rect 31980 -2620 32015 -2585
rect 32025 -2620 32060 -2585
rect 32070 -2620 32105 -2585
rect 32115 -2620 32150 -2585
rect 32160 -2620 32195 -2585
rect 32205 -2620 32240 -2585
rect 32250 -2620 32285 -2585
rect 32295 -2620 32330 -2585
rect 32340 -2620 32375 -2585
rect 32385 -2620 32420 -2585
rect 32430 -2620 32465 -2585
rect 32475 -2620 32510 -2585
rect 32520 -2620 32555 -2585
rect 32565 -2620 32600 -2585
rect 32610 -2620 32645 -2585
rect 32655 -2620 32690 -2585
rect 32700 -2620 32735 -2585
rect 32745 -2620 32780 -2585
rect 32790 -2620 32825 -2585
rect 32835 -2620 32870 -2585
rect 31305 -2665 31340 -2630
rect 31350 -2665 31385 -2630
rect 31395 -2665 31430 -2630
rect 31440 -2665 31475 -2630
rect 31485 -2665 31520 -2630
rect 31530 -2665 31565 -2630
rect 31575 -2665 31610 -2630
rect 31620 -2665 31655 -2630
rect 31665 -2665 31700 -2630
rect 31710 -2665 31745 -2630
rect 31755 -2665 31790 -2630
rect 31800 -2665 31835 -2630
rect 31845 -2665 31880 -2630
rect 31890 -2665 31925 -2630
rect 31935 -2665 31970 -2630
rect 31980 -2665 32015 -2630
rect 32025 -2665 32060 -2630
rect 32070 -2665 32105 -2630
rect 32115 -2665 32150 -2630
rect 32160 -2665 32195 -2630
rect 32205 -2665 32240 -2630
rect 32250 -2665 32285 -2630
rect 32295 -2665 32330 -2630
rect 32340 -2665 32375 -2630
rect 32385 -2665 32420 -2630
rect 32430 -2665 32465 -2630
rect 32475 -2665 32510 -2630
rect 32520 -2665 32555 -2630
rect 32565 -2665 32600 -2630
rect 32610 -2665 32645 -2630
rect 32655 -2665 32690 -2630
rect 32700 -2665 32735 -2630
rect 32745 -2665 32780 -2630
rect 32790 -2665 32825 -2630
rect 32835 -2665 32870 -2630
rect 31305 -2710 31340 -2675
rect 31350 -2710 31385 -2675
rect 31395 -2710 31430 -2675
rect 31440 -2710 31475 -2675
rect 31485 -2710 31520 -2675
rect 31530 -2710 31565 -2675
rect 31575 -2710 31610 -2675
rect 31620 -2710 31655 -2675
rect 31665 -2710 31700 -2675
rect 31710 -2710 31745 -2675
rect 31755 -2710 31790 -2675
rect 31800 -2710 31835 -2675
rect 31845 -2710 31880 -2675
rect 31890 -2710 31925 -2675
rect 31935 -2710 31970 -2675
rect 31980 -2710 32015 -2675
rect 32025 -2710 32060 -2675
rect 32070 -2710 32105 -2675
rect 32115 -2710 32150 -2675
rect 32160 -2710 32195 -2675
rect 32205 -2710 32240 -2675
rect 32250 -2710 32285 -2675
rect 32295 -2710 32330 -2675
rect 32340 -2710 32375 -2675
rect 32385 -2710 32420 -2675
rect 32430 -2710 32465 -2675
rect 32475 -2710 32510 -2675
rect 32520 -2710 32555 -2675
rect 32565 -2710 32600 -2675
rect 32610 -2710 32645 -2675
rect 32655 -2710 32690 -2675
rect 32700 -2710 32735 -2675
rect 32745 -2710 32780 -2675
rect 32790 -2710 32825 -2675
rect 32835 -2710 32870 -2675
rect 31305 -2755 31340 -2720
rect 31350 -2755 31385 -2720
rect 31395 -2755 31430 -2720
rect 31440 -2755 31475 -2720
rect 31485 -2755 31520 -2720
rect 31530 -2755 31565 -2720
rect 31575 -2755 31610 -2720
rect 31620 -2755 31655 -2720
rect 31665 -2755 31700 -2720
rect 31710 -2755 31745 -2720
rect 31755 -2755 31790 -2720
rect 31800 -2755 31835 -2720
rect 31845 -2755 31880 -2720
rect 31890 -2755 31925 -2720
rect 31935 -2755 31970 -2720
rect 31980 -2755 32015 -2720
rect 32025 -2755 32060 -2720
rect 32070 -2755 32105 -2720
rect 32115 -2755 32150 -2720
rect 32160 -2755 32195 -2720
rect 32205 -2755 32240 -2720
rect 32250 -2755 32285 -2720
rect 32295 -2755 32330 -2720
rect 32340 -2755 32375 -2720
rect 32385 -2755 32420 -2720
rect 32430 -2755 32465 -2720
rect 32475 -2755 32510 -2720
rect 32520 -2755 32555 -2720
rect 32565 -2755 32600 -2720
rect 32610 -2755 32645 -2720
rect 32655 -2755 32690 -2720
rect 32700 -2755 32735 -2720
rect 32745 -2755 32780 -2720
rect 32790 -2755 32825 -2720
rect 32835 -2755 32870 -2720
rect 31305 -2800 31340 -2765
rect 31350 -2800 31385 -2765
rect 31395 -2800 31430 -2765
rect 31440 -2800 31475 -2765
rect 31485 -2800 31520 -2765
rect 31530 -2800 31565 -2765
rect 31575 -2800 31610 -2765
rect 31620 -2800 31655 -2765
rect 31665 -2800 31700 -2765
rect 31710 -2800 31745 -2765
rect 31755 -2800 31790 -2765
rect 31800 -2800 31835 -2765
rect 31845 -2800 31880 -2765
rect 31890 -2800 31925 -2765
rect 31935 -2800 31970 -2765
rect 31980 -2800 32015 -2765
rect 32025 -2800 32060 -2765
rect 32070 -2800 32105 -2765
rect 32115 -2800 32150 -2765
rect 32160 -2800 32195 -2765
rect 32205 -2800 32240 -2765
rect 32250 -2800 32285 -2765
rect 32295 -2800 32330 -2765
rect 32340 -2800 32375 -2765
rect 32385 -2800 32420 -2765
rect 32430 -2800 32465 -2765
rect 32475 -2800 32510 -2765
rect 32520 -2800 32555 -2765
rect 32565 -2800 32600 -2765
rect 32610 -2800 32645 -2765
rect 32655 -2800 32690 -2765
rect 32700 -2800 32735 -2765
rect 32745 -2800 32780 -2765
rect 32790 -2800 32825 -2765
rect 32835 -2800 32870 -2765
rect 31305 -2845 31340 -2810
rect 31350 -2845 31385 -2810
rect 31395 -2845 31430 -2810
rect 31440 -2845 31475 -2810
rect 31485 -2845 31520 -2810
rect 31530 -2845 31565 -2810
rect 31575 -2845 31610 -2810
rect 31620 -2845 31655 -2810
rect 31665 -2845 31700 -2810
rect 31710 -2845 31745 -2810
rect 31755 -2845 31790 -2810
rect 31800 -2845 31835 -2810
rect 31845 -2845 31880 -2810
rect 31890 -2845 31925 -2810
rect 31935 -2845 31970 -2810
rect 31980 -2845 32015 -2810
rect 32025 -2845 32060 -2810
rect 32070 -2845 32105 -2810
rect 32115 -2845 32150 -2810
rect 32160 -2845 32195 -2810
rect 32205 -2845 32240 -2810
rect 32250 -2845 32285 -2810
rect 32295 -2845 32330 -2810
rect 32340 -2845 32375 -2810
rect 32385 -2845 32420 -2810
rect 32430 -2845 32465 -2810
rect 32475 -2845 32510 -2810
rect 32520 -2845 32555 -2810
rect 32565 -2845 32600 -2810
rect 32610 -2845 32645 -2810
rect 32655 -2845 32690 -2810
rect 32700 -2845 32735 -2810
rect 32745 -2845 32780 -2810
rect 32790 -2845 32825 -2810
rect 32835 -2845 32870 -2810
rect 31305 -2890 31340 -2855
rect 31350 -2890 31385 -2855
rect 31395 -2890 31430 -2855
rect 31440 -2890 31475 -2855
rect 31485 -2890 31520 -2855
rect 31530 -2890 31565 -2855
rect 31575 -2890 31610 -2855
rect 31620 -2890 31655 -2855
rect 31665 -2890 31700 -2855
rect 31710 -2890 31745 -2855
rect 31755 -2890 31790 -2855
rect 31800 -2890 31835 -2855
rect 31845 -2890 31880 -2855
rect 31890 -2890 31925 -2855
rect 31935 -2890 31970 -2855
rect 31980 -2890 32015 -2855
rect 32025 -2890 32060 -2855
rect 32070 -2890 32105 -2855
rect 32115 -2890 32150 -2855
rect 32160 -2890 32195 -2855
rect 32205 -2890 32240 -2855
rect 32250 -2890 32285 -2855
rect 32295 -2890 32330 -2855
rect 32340 -2890 32375 -2855
rect 32385 -2890 32420 -2855
rect 32430 -2890 32465 -2855
rect 32475 -2890 32510 -2855
rect 32520 -2890 32555 -2855
rect 32565 -2890 32600 -2855
rect 32610 -2890 32645 -2855
rect 32655 -2890 32690 -2855
rect 32700 -2890 32735 -2855
rect 32745 -2890 32780 -2855
rect 32790 -2890 32825 -2855
rect 32835 -2890 32870 -2855
rect 3420 -3020 3460 -3015
rect 3420 -3050 3425 -3020
rect 3425 -3050 3455 -3020
rect 3455 -3050 3460 -3020
rect 3420 -3055 3460 -3050
rect 3420 -3085 3460 -3080
rect 3420 -3115 3425 -3085
rect 3425 -3115 3455 -3085
rect 3455 -3115 3460 -3085
rect 3420 -3120 3460 -3115
rect 3420 -3155 3460 -3150
rect 3420 -3185 3425 -3155
rect 3425 -3185 3455 -3155
rect 3455 -3185 3460 -3155
rect 3420 -3190 3460 -3185
rect 3420 -3225 3460 -3220
rect 3420 -3255 3425 -3225
rect 3425 -3255 3455 -3225
rect 3455 -3255 3460 -3225
rect 3420 -3260 3460 -3255
rect 3420 -3295 3460 -3290
rect 3420 -3325 3425 -3295
rect 3425 -3325 3455 -3295
rect 3455 -3325 3460 -3295
rect 3420 -3330 3460 -3325
rect 3420 -3360 3460 -3355
rect 3420 -3390 3425 -3360
rect 3425 -3390 3455 -3360
rect 3455 -3390 3460 -3360
rect 3420 -3395 3460 -3390
rect 3420 -3420 3460 -3415
rect 3420 -3450 3425 -3420
rect 3425 -3450 3455 -3420
rect 3455 -3450 3460 -3420
rect 3420 -3455 3460 -3450
rect 3420 -3485 3460 -3480
rect 3420 -3515 3425 -3485
rect 3425 -3515 3455 -3485
rect 3455 -3515 3460 -3485
rect 3420 -3520 3460 -3515
rect 3420 -3555 3460 -3550
rect 3420 -3585 3425 -3555
rect 3425 -3585 3455 -3555
rect 3455 -3585 3460 -3555
rect 3420 -3590 3460 -3585
rect 3420 -3625 3460 -3620
rect 3420 -3655 3425 -3625
rect 3425 -3655 3455 -3625
rect 3455 -3655 3460 -3625
rect 3420 -3660 3460 -3655
rect 3420 -3695 3460 -3690
rect 3420 -3725 3425 -3695
rect 3425 -3725 3455 -3695
rect 3455 -3725 3460 -3695
rect 3420 -3730 3460 -3725
rect 3420 -3760 3460 -3755
rect 3420 -3790 3425 -3760
rect 3425 -3790 3455 -3760
rect 3455 -3790 3460 -3760
rect 3420 -3795 3460 -3790
rect 3420 -3820 3460 -3815
rect 3420 -3850 3425 -3820
rect 3425 -3850 3455 -3820
rect 3455 -3850 3460 -3820
rect 3420 -3855 3460 -3850
rect 3420 -3885 3460 -3880
rect 3420 -3915 3425 -3885
rect 3425 -3915 3455 -3885
rect 3455 -3915 3460 -3885
rect 3420 -3920 3460 -3915
rect 3420 -3955 3460 -3950
rect 3420 -3985 3425 -3955
rect 3425 -3985 3455 -3955
rect 3455 -3985 3460 -3955
rect 3420 -3990 3460 -3985
rect 3420 -4025 3460 -4020
rect 3420 -4055 3425 -4025
rect 3425 -4055 3455 -4025
rect 3455 -4055 3460 -4025
rect 3420 -4060 3460 -4055
rect 3420 -4095 3460 -4090
rect 3420 -4125 3425 -4095
rect 3425 -4125 3455 -4095
rect 3455 -4125 3460 -4095
rect 3420 -4130 3460 -4125
rect 3420 -4160 3460 -4155
rect 3420 -4190 3425 -4160
rect 3425 -4190 3455 -4160
rect 3455 -4190 3460 -4160
rect 3420 -4195 3460 -4190
rect 3420 -4220 3460 -4215
rect 3420 -4250 3425 -4220
rect 3425 -4250 3455 -4220
rect 3455 -4250 3460 -4220
rect 3420 -4255 3460 -4250
rect 3420 -4285 3460 -4280
rect 3420 -4315 3425 -4285
rect 3425 -4315 3455 -4285
rect 3455 -4315 3460 -4285
rect 3420 -4320 3460 -4315
rect 3420 -4355 3460 -4350
rect 3420 -4385 3425 -4355
rect 3425 -4385 3455 -4355
rect 3455 -4385 3460 -4355
rect 3420 -4390 3460 -4385
rect 3420 -4425 3460 -4420
rect 3420 -4455 3425 -4425
rect 3425 -4455 3455 -4425
rect 3455 -4455 3460 -4425
rect 3420 -4460 3460 -4455
rect 3420 -4495 3460 -4490
rect 3420 -4525 3425 -4495
rect 3425 -4525 3455 -4495
rect 3455 -4525 3460 -4495
rect 3420 -4530 3460 -4525
rect 3420 -4560 3460 -4555
rect 3420 -4590 3425 -4560
rect 3425 -4590 3455 -4560
rect 3455 -4590 3460 -4560
rect 3420 -4595 3460 -4590
rect 3770 -3020 3810 -3015
rect 3770 -3050 3775 -3020
rect 3775 -3050 3805 -3020
rect 3805 -3050 3810 -3020
rect 3770 -3055 3810 -3050
rect 3770 -3085 3810 -3080
rect 3770 -3115 3775 -3085
rect 3775 -3115 3805 -3085
rect 3805 -3115 3810 -3085
rect 3770 -3120 3810 -3115
rect 3770 -3155 3810 -3150
rect 3770 -3185 3775 -3155
rect 3775 -3185 3805 -3155
rect 3805 -3185 3810 -3155
rect 3770 -3190 3810 -3185
rect 3770 -3225 3810 -3220
rect 3770 -3255 3775 -3225
rect 3775 -3255 3805 -3225
rect 3805 -3255 3810 -3225
rect 3770 -3260 3810 -3255
rect 3770 -3295 3810 -3290
rect 3770 -3325 3775 -3295
rect 3775 -3325 3805 -3295
rect 3805 -3325 3810 -3295
rect 3770 -3330 3810 -3325
rect 3770 -3360 3810 -3355
rect 3770 -3390 3775 -3360
rect 3775 -3390 3805 -3360
rect 3805 -3390 3810 -3360
rect 3770 -3395 3810 -3390
rect 3770 -3420 3810 -3415
rect 3770 -3450 3775 -3420
rect 3775 -3450 3805 -3420
rect 3805 -3450 3810 -3420
rect 3770 -3455 3810 -3450
rect 3770 -3485 3810 -3480
rect 3770 -3515 3775 -3485
rect 3775 -3515 3805 -3485
rect 3805 -3515 3810 -3485
rect 3770 -3520 3810 -3515
rect 3770 -3555 3810 -3550
rect 3770 -3585 3775 -3555
rect 3775 -3585 3805 -3555
rect 3805 -3585 3810 -3555
rect 3770 -3590 3810 -3585
rect 3770 -3625 3810 -3620
rect 3770 -3655 3775 -3625
rect 3775 -3655 3805 -3625
rect 3805 -3655 3810 -3625
rect 3770 -3660 3810 -3655
rect 3770 -3695 3810 -3690
rect 3770 -3725 3775 -3695
rect 3775 -3725 3805 -3695
rect 3805 -3725 3810 -3695
rect 3770 -3730 3810 -3725
rect 3770 -3760 3810 -3755
rect 3770 -3790 3775 -3760
rect 3775 -3790 3805 -3760
rect 3805 -3790 3810 -3760
rect 3770 -3795 3810 -3790
rect 3770 -3820 3810 -3815
rect 3770 -3850 3775 -3820
rect 3775 -3850 3805 -3820
rect 3805 -3850 3810 -3820
rect 3770 -3855 3810 -3850
rect 3770 -3885 3810 -3880
rect 3770 -3915 3775 -3885
rect 3775 -3915 3805 -3885
rect 3805 -3915 3810 -3885
rect 3770 -3920 3810 -3915
rect 3770 -3955 3810 -3950
rect 3770 -3985 3775 -3955
rect 3775 -3985 3805 -3955
rect 3805 -3985 3810 -3955
rect 3770 -3990 3810 -3985
rect 3770 -4025 3810 -4020
rect 3770 -4055 3775 -4025
rect 3775 -4055 3805 -4025
rect 3805 -4055 3810 -4025
rect 3770 -4060 3810 -4055
rect 3770 -4095 3810 -4090
rect 3770 -4125 3775 -4095
rect 3775 -4125 3805 -4095
rect 3805 -4125 3810 -4095
rect 3770 -4130 3810 -4125
rect 3770 -4160 3810 -4155
rect 3770 -4190 3775 -4160
rect 3775 -4190 3805 -4160
rect 3805 -4190 3810 -4160
rect 3770 -4195 3810 -4190
rect 3770 -4220 3810 -4215
rect 3770 -4250 3775 -4220
rect 3775 -4250 3805 -4220
rect 3805 -4250 3810 -4220
rect 3770 -4255 3810 -4250
rect 3770 -4285 3810 -4280
rect 3770 -4315 3775 -4285
rect 3775 -4315 3805 -4285
rect 3805 -4315 3810 -4285
rect 3770 -4320 3810 -4315
rect 3770 -4355 3810 -4350
rect 3770 -4385 3775 -4355
rect 3775 -4385 3805 -4355
rect 3805 -4385 3810 -4355
rect 3770 -4390 3810 -4385
rect 3770 -4425 3810 -4420
rect 3770 -4455 3775 -4425
rect 3775 -4455 3805 -4425
rect 3805 -4455 3810 -4425
rect 3770 -4460 3810 -4455
rect 3770 -4495 3810 -4490
rect 3770 -4525 3775 -4495
rect 3775 -4525 3805 -4495
rect 3805 -4525 3810 -4495
rect 3770 -4530 3810 -4525
rect 3770 -4560 3810 -4555
rect 3770 -4590 3775 -4560
rect 3775 -4590 3805 -4560
rect 3805 -4590 3810 -4560
rect 3770 -4595 3810 -4590
rect 4120 -3020 4160 -3015
rect 4120 -3050 4125 -3020
rect 4125 -3050 4155 -3020
rect 4155 -3050 4160 -3020
rect 4120 -3055 4160 -3050
rect 4120 -3085 4160 -3080
rect 4120 -3115 4125 -3085
rect 4125 -3115 4155 -3085
rect 4155 -3115 4160 -3085
rect 4120 -3120 4160 -3115
rect 4120 -3155 4160 -3150
rect 4120 -3185 4125 -3155
rect 4125 -3185 4155 -3155
rect 4155 -3185 4160 -3155
rect 4120 -3190 4160 -3185
rect 4120 -3225 4160 -3220
rect 4120 -3255 4125 -3225
rect 4125 -3255 4155 -3225
rect 4155 -3255 4160 -3225
rect 4120 -3260 4160 -3255
rect 4120 -3295 4160 -3290
rect 4120 -3325 4125 -3295
rect 4125 -3325 4155 -3295
rect 4155 -3325 4160 -3295
rect 4120 -3330 4160 -3325
rect 4120 -3360 4160 -3355
rect 4120 -3390 4125 -3360
rect 4125 -3390 4155 -3360
rect 4155 -3390 4160 -3360
rect 4120 -3395 4160 -3390
rect 4120 -3420 4160 -3415
rect 4120 -3450 4125 -3420
rect 4125 -3450 4155 -3420
rect 4155 -3450 4160 -3420
rect 4120 -3455 4160 -3450
rect 4120 -3485 4160 -3480
rect 4120 -3515 4125 -3485
rect 4125 -3515 4155 -3485
rect 4155 -3515 4160 -3485
rect 4120 -3520 4160 -3515
rect 4120 -3555 4160 -3550
rect 4120 -3585 4125 -3555
rect 4125 -3585 4155 -3555
rect 4155 -3585 4160 -3555
rect 4120 -3590 4160 -3585
rect 4120 -3625 4160 -3620
rect 4120 -3655 4125 -3625
rect 4125 -3655 4155 -3625
rect 4155 -3655 4160 -3625
rect 4120 -3660 4160 -3655
rect 4120 -3695 4160 -3690
rect 4120 -3725 4125 -3695
rect 4125 -3725 4155 -3695
rect 4155 -3725 4160 -3695
rect 4120 -3730 4160 -3725
rect 4120 -3760 4160 -3755
rect 4120 -3790 4125 -3760
rect 4125 -3790 4155 -3760
rect 4155 -3790 4160 -3760
rect 4120 -3795 4160 -3790
rect 4120 -3820 4160 -3815
rect 4120 -3850 4125 -3820
rect 4125 -3850 4155 -3820
rect 4155 -3850 4160 -3820
rect 4120 -3855 4160 -3850
rect 4120 -3885 4160 -3880
rect 4120 -3915 4125 -3885
rect 4125 -3915 4155 -3885
rect 4155 -3915 4160 -3885
rect 4120 -3920 4160 -3915
rect 4120 -3955 4160 -3950
rect 4120 -3985 4125 -3955
rect 4125 -3985 4155 -3955
rect 4155 -3985 4160 -3955
rect 4120 -3990 4160 -3985
rect 4120 -4025 4160 -4020
rect 4120 -4055 4125 -4025
rect 4125 -4055 4155 -4025
rect 4155 -4055 4160 -4025
rect 4120 -4060 4160 -4055
rect 4120 -4095 4160 -4090
rect 4120 -4125 4125 -4095
rect 4125 -4125 4155 -4095
rect 4155 -4125 4160 -4095
rect 4120 -4130 4160 -4125
rect 4120 -4160 4160 -4155
rect 4120 -4190 4125 -4160
rect 4125 -4190 4155 -4160
rect 4155 -4190 4160 -4160
rect 4120 -4195 4160 -4190
rect 4120 -4220 4160 -4215
rect 4120 -4250 4125 -4220
rect 4125 -4250 4155 -4220
rect 4155 -4250 4160 -4220
rect 4120 -4255 4160 -4250
rect 4120 -4285 4160 -4280
rect 4120 -4315 4125 -4285
rect 4125 -4315 4155 -4285
rect 4155 -4315 4160 -4285
rect 4120 -4320 4160 -4315
rect 4120 -4355 4160 -4350
rect 4120 -4385 4125 -4355
rect 4125 -4385 4155 -4355
rect 4155 -4385 4160 -4355
rect 4120 -4390 4160 -4385
rect 4120 -4425 4160 -4420
rect 4120 -4455 4125 -4425
rect 4125 -4455 4155 -4425
rect 4155 -4455 4160 -4425
rect 4120 -4460 4160 -4455
rect 4120 -4495 4160 -4490
rect 4120 -4525 4125 -4495
rect 4125 -4525 4155 -4495
rect 4155 -4525 4160 -4495
rect 4120 -4530 4160 -4525
rect 4120 -4560 4160 -4555
rect 4120 -4590 4125 -4560
rect 4125 -4590 4155 -4560
rect 4155 -4590 4160 -4560
rect 4120 -4595 4160 -4590
rect 4470 -3020 4510 -3015
rect 4470 -3050 4475 -3020
rect 4475 -3050 4505 -3020
rect 4505 -3050 4510 -3020
rect 4470 -3055 4510 -3050
rect 4470 -3085 4510 -3080
rect 4470 -3115 4475 -3085
rect 4475 -3115 4505 -3085
rect 4505 -3115 4510 -3085
rect 4470 -3120 4510 -3115
rect 4470 -3155 4510 -3150
rect 4470 -3185 4475 -3155
rect 4475 -3185 4505 -3155
rect 4505 -3185 4510 -3155
rect 4470 -3190 4510 -3185
rect 4470 -3225 4510 -3220
rect 4470 -3255 4475 -3225
rect 4475 -3255 4505 -3225
rect 4505 -3255 4510 -3225
rect 4470 -3260 4510 -3255
rect 4470 -3295 4510 -3290
rect 4470 -3325 4475 -3295
rect 4475 -3325 4505 -3295
rect 4505 -3325 4510 -3295
rect 4470 -3330 4510 -3325
rect 4470 -3360 4510 -3355
rect 4470 -3390 4475 -3360
rect 4475 -3390 4505 -3360
rect 4505 -3390 4510 -3360
rect 4470 -3395 4510 -3390
rect 4470 -3420 4510 -3415
rect 4470 -3450 4475 -3420
rect 4475 -3450 4505 -3420
rect 4505 -3450 4510 -3420
rect 4470 -3455 4510 -3450
rect 4470 -3485 4510 -3480
rect 4470 -3515 4475 -3485
rect 4475 -3515 4505 -3485
rect 4505 -3515 4510 -3485
rect 4470 -3520 4510 -3515
rect 4470 -3555 4510 -3550
rect 4470 -3585 4475 -3555
rect 4475 -3585 4505 -3555
rect 4505 -3585 4510 -3555
rect 4470 -3590 4510 -3585
rect 4470 -3625 4510 -3620
rect 4470 -3655 4475 -3625
rect 4475 -3655 4505 -3625
rect 4505 -3655 4510 -3625
rect 4470 -3660 4510 -3655
rect 4470 -3695 4510 -3690
rect 4470 -3725 4475 -3695
rect 4475 -3725 4505 -3695
rect 4505 -3725 4510 -3695
rect 4470 -3730 4510 -3725
rect 4470 -3760 4510 -3755
rect 4470 -3790 4475 -3760
rect 4475 -3790 4505 -3760
rect 4505 -3790 4510 -3760
rect 4470 -3795 4510 -3790
rect 4470 -3820 4510 -3815
rect 4470 -3850 4475 -3820
rect 4475 -3850 4505 -3820
rect 4505 -3850 4510 -3820
rect 4470 -3855 4510 -3850
rect 4470 -3885 4510 -3880
rect 4470 -3915 4475 -3885
rect 4475 -3915 4505 -3885
rect 4505 -3915 4510 -3885
rect 4470 -3920 4510 -3915
rect 4470 -3955 4510 -3950
rect 4470 -3985 4475 -3955
rect 4475 -3985 4505 -3955
rect 4505 -3985 4510 -3955
rect 4470 -3990 4510 -3985
rect 4470 -4025 4510 -4020
rect 4470 -4055 4475 -4025
rect 4475 -4055 4505 -4025
rect 4505 -4055 4510 -4025
rect 4470 -4060 4510 -4055
rect 4470 -4095 4510 -4090
rect 4470 -4125 4475 -4095
rect 4475 -4125 4505 -4095
rect 4505 -4125 4510 -4095
rect 4470 -4130 4510 -4125
rect 4470 -4160 4510 -4155
rect 4470 -4190 4475 -4160
rect 4475 -4190 4505 -4160
rect 4505 -4190 4510 -4160
rect 4470 -4195 4510 -4190
rect 4470 -4220 4510 -4215
rect 4470 -4250 4475 -4220
rect 4475 -4250 4505 -4220
rect 4505 -4250 4510 -4220
rect 4470 -4255 4510 -4250
rect 4470 -4285 4510 -4280
rect 4470 -4315 4475 -4285
rect 4475 -4315 4505 -4285
rect 4505 -4315 4510 -4285
rect 4470 -4320 4510 -4315
rect 4470 -4355 4510 -4350
rect 4470 -4385 4475 -4355
rect 4475 -4385 4505 -4355
rect 4505 -4385 4510 -4355
rect 4470 -4390 4510 -4385
rect 4470 -4425 4510 -4420
rect 4470 -4455 4475 -4425
rect 4475 -4455 4505 -4425
rect 4505 -4455 4510 -4425
rect 4470 -4460 4510 -4455
rect 4470 -4495 4510 -4490
rect 4470 -4525 4475 -4495
rect 4475 -4525 4505 -4495
rect 4505 -4525 4510 -4495
rect 4470 -4530 4510 -4525
rect 4470 -4560 4510 -4555
rect 4470 -4590 4475 -4560
rect 4475 -4590 4505 -4560
rect 4505 -4590 4510 -4560
rect 4470 -4595 4510 -4590
rect 4820 -3020 4860 -3015
rect 4820 -3050 4825 -3020
rect 4825 -3050 4855 -3020
rect 4855 -3050 4860 -3020
rect 4820 -3055 4860 -3050
rect 4820 -3085 4860 -3080
rect 4820 -3115 4825 -3085
rect 4825 -3115 4855 -3085
rect 4855 -3115 4860 -3085
rect 4820 -3120 4860 -3115
rect 4820 -3155 4860 -3150
rect 4820 -3185 4825 -3155
rect 4825 -3185 4855 -3155
rect 4855 -3185 4860 -3155
rect 4820 -3190 4860 -3185
rect 4820 -3225 4860 -3220
rect 4820 -3255 4825 -3225
rect 4825 -3255 4855 -3225
rect 4855 -3255 4860 -3225
rect 4820 -3260 4860 -3255
rect 4820 -3295 4860 -3290
rect 4820 -3325 4825 -3295
rect 4825 -3325 4855 -3295
rect 4855 -3325 4860 -3295
rect 4820 -3330 4860 -3325
rect 4820 -3360 4860 -3355
rect 4820 -3390 4825 -3360
rect 4825 -3390 4855 -3360
rect 4855 -3390 4860 -3360
rect 4820 -3395 4860 -3390
rect 4820 -3420 4860 -3415
rect 4820 -3450 4825 -3420
rect 4825 -3450 4855 -3420
rect 4855 -3450 4860 -3420
rect 4820 -3455 4860 -3450
rect 4820 -3485 4860 -3480
rect 4820 -3515 4825 -3485
rect 4825 -3515 4855 -3485
rect 4855 -3515 4860 -3485
rect 4820 -3520 4860 -3515
rect 4820 -3555 4860 -3550
rect 4820 -3585 4825 -3555
rect 4825 -3585 4855 -3555
rect 4855 -3585 4860 -3555
rect 4820 -3590 4860 -3585
rect 4820 -3625 4860 -3620
rect 4820 -3655 4825 -3625
rect 4825 -3655 4855 -3625
rect 4855 -3655 4860 -3625
rect 4820 -3660 4860 -3655
rect 4820 -3695 4860 -3690
rect 4820 -3725 4825 -3695
rect 4825 -3725 4855 -3695
rect 4855 -3725 4860 -3695
rect 4820 -3730 4860 -3725
rect 4820 -3760 4860 -3755
rect 4820 -3790 4825 -3760
rect 4825 -3790 4855 -3760
rect 4855 -3790 4860 -3760
rect 4820 -3795 4860 -3790
rect 4820 -3820 4860 -3815
rect 4820 -3850 4825 -3820
rect 4825 -3850 4855 -3820
rect 4855 -3850 4860 -3820
rect 4820 -3855 4860 -3850
rect 4820 -3885 4860 -3880
rect 4820 -3915 4825 -3885
rect 4825 -3915 4855 -3885
rect 4855 -3915 4860 -3885
rect 4820 -3920 4860 -3915
rect 4820 -3955 4860 -3950
rect 4820 -3985 4825 -3955
rect 4825 -3985 4855 -3955
rect 4855 -3985 4860 -3955
rect 4820 -3990 4860 -3985
rect 4820 -4025 4860 -4020
rect 4820 -4055 4825 -4025
rect 4825 -4055 4855 -4025
rect 4855 -4055 4860 -4025
rect 4820 -4060 4860 -4055
rect 4820 -4095 4860 -4090
rect 4820 -4125 4825 -4095
rect 4825 -4125 4855 -4095
rect 4855 -4125 4860 -4095
rect 4820 -4130 4860 -4125
rect 4820 -4160 4860 -4155
rect 4820 -4190 4825 -4160
rect 4825 -4190 4855 -4160
rect 4855 -4190 4860 -4160
rect 4820 -4195 4860 -4190
rect 4820 -4220 4860 -4215
rect 4820 -4250 4825 -4220
rect 4825 -4250 4855 -4220
rect 4855 -4250 4860 -4220
rect 4820 -4255 4860 -4250
rect 4820 -4285 4860 -4280
rect 4820 -4315 4825 -4285
rect 4825 -4315 4855 -4285
rect 4855 -4315 4860 -4285
rect 4820 -4320 4860 -4315
rect 4820 -4355 4860 -4350
rect 4820 -4385 4825 -4355
rect 4825 -4385 4855 -4355
rect 4855 -4385 4860 -4355
rect 4820 -4390 4860 -4385
rect 4820 -4425 4860 -4420
rect 4820 -4455 4825 -4425
rect 4825 -4455 4855 -4425
rect 4855 -4455 4860 -4425
rect 4820 -4460 4860 -4455
rect 4820 -4495 4860 -4490
rect 4820 -4525 4825 -4495
rect 4825 -4525 4855 -4495
rect 4855 -4525 4860 -4495
rect 4820 -4530 4860 -4525
rect 4820 -4560 4860 -4555
rect 4820 -4590 4825 -4560
rect 4825 -4590 4855 -4560
rect 4855 -4590 4860 -4560
rect 4820 -4595 4860 -4590
rect 5170 -3020 5210 -3015
rect 5170 -3050 5175 -3020
rect 5175 -3050 5205 -3020
rect 5205 -3050 5210 -3020
rect 5170 -3055 5210 -3050
rect 5170 -3085 5210 -3080
rect 5170 -3115 5175 -3085
rect 5175 -3115 5205 -3085
rect 5205 -3115 5210 -3085
rect 5170 -3120 5210 -3115
rect 5170 -3155 5210 -3150
rect 5170 -3185 5175 -3155
rect 5175 -3185 5205 -3155
rect 5205 -3185 5210 -3155
rect 5170 -3190 5210 -3185
rect 5170 -3225 5210 -3220
rect 5170 -3255 5175 -3225
rect 5175 -3255 5205 -3225
rect 5205 -3255 5210 -3225
rect 5170 -3260 5210 -3255
rect 5170 -3295 5210 -3290
rect 5170 -3325 5175 -3295
rect 5175 -3325 5205 -3295
rect 5205 -3325 5210 -3295
rect 5170 -3330 5210 -3325
rect 5170 -3360 5210 -3355
rect 5170 -3390 5175 -3360
rect 5175 -3390 5205 -3360
rect 5205 -3390 5210 -3360
rect 5170 -3395 5210 -3390
rect 5170 -3420 5210 -3415
rect 5170 -3450 5175 -3420
rect 5175 -3450 5205 -3420
rect 5205 -3450 5210 -3420
rect 5170 -3455 5210 -3450
rect 5170 -3485 5210 -3480
rect 5170 -3515 5175 -3485
rect 5175 -3515 5205 -3485
rect 5205 -3515 5210 -3485
rect 5170 -3520 5210 -3515
rect 5170 -3555 5210 -3550
rect 5170 -3585 5175 -3555
rect 5175 -3585 5205 -3555
rect 5205 -3585 5210 -3555
rect 5170 -3590 5210 -3585
rect 5170 -3625 5210 -3620
rect 5170 -3655 5175 -3625
rect 5175 -3655 5205 -3625
rect 5205 -3655 5210 -3625
rect 5170 -3660 5210 -3655
rect 5170 -3695 5210 -3690
rect 5170 -3725 5175 -3695
rect 5175 -3725 5205 -3695
rect 5205 -3725 5210 -3695
rect 5170 -3730 5210 -3725
rect 5170 -3760 5210 -3755
rect 5170 -3790 5175 -3760
rect 5175 -3790 5205 -3760
rect 5205 -3790 5210 -3760
rect 5170 -3795 5210 -3790
rect 5170 -3820 5210 -3815
rect 5170 -3850 5175 -3820
rect 5175 -3850 5205 -3820
rect 5205 -3850 5210 -3820
rect 5170 -3855 5210 -3850
rect 5170 -3885 5210 -3880
rect 5170 -3915 5175 -3885
rect 5175 -3915 5205 -3885
rect 5205 -3915 5210 -3885
rect 5170 -3920 5210 -3915
rect 5170 -3955 5210 -3950
rect 5170 -3985 5175 -3955
rect 5175 -3985 5205 -3955
rect 5205 -3985 5210 -3955
rect 5170 -3990 5210 -3985
rect 5170 -4025 5210 -4020
rect 5170 -4055 5175 -4025
rect 5175 -4055 5205 -4025
rect 5205 -4055 5210 -4025
rect 5170 -4060 5210 -4055
rect 5170 -4095 5210 -4090
rect 5170 -4125 5175 -4095
rect 5175 -4125 5205 -4095
rect 5205 -4125 5210 -4095
rect 5170 -4130 5210 -4125
rect 5170 -4160 5210 -4155
rect 5170 -4190 5175 -4160
rect 5175 -4190 5205 -4160
rect 5205 -4190 5210 -4160
rect 5170 -4195 5210 -4190
rect 5170 -4220 5210 -4215
rect 5170 -4250 5175 -4220
rect 5175 -4250 5205 -4220
rect 5205 -4250 5210 -4220
rect 5170 -4255 5210 -4250
rect 5170 -4285 5210 -4280
rect 5170 -4315 5175 -4285
rect 5175 -4315 5205 -4285
rect 5205 -4315 5210 -4285
rect 5170 -4320 5210 -4315
rect 5170 -4355 5210 -4350
rect 5170 -4385 5175 -4355
rect 5175 -4385 5205 -4355
rect 5205 -4385 5210 -4355
rect 5170 -4390 5210 -4385
rect 5170 -4425 5210 -4420
rect 5170 -4455 5175 -4425
rect 5175 -4455 5205 -4425
rect 5205 -4455 5210 -4425
rect 5170 -4460 5210 -4455
rect 5170 -4495 5210 -4490
rect 5170 -4525 5175 -4495
rect 5175 -4525 5205 -4495
rect 5205 -4525 5210 -4495
rect 5170 -4530 5210 -4525
rect 5170 -4560 5210 -4555
rect 5170 -4590 5175 -4560
rect 5175 -4590 5205 -4560
rect 5205 -4590 5210 -4560
rect 5170 -4595 5210 -4590
rect 5520 -3020 5560 -3015
rect 5520 -3050 5525 -3020
rect 5525 -3050 5555 -3020
rect 5555 -3050 5560 -3020
rect 5520 -3055 5560 -3050
rect 5520 -3085 5560 -3080
rect 5520 -3115 5525 -3085
rect 5525 -3115 5555 -3085
rect 5555 -3115 5560 -3085
rect 5520 -3120 5560 -3115
rect 5520 -3155 5560 -3150
rect 5520 -3185 5525 -3155
rect 5525 -3185 5555 -3155
rect 5555 -3185 5560 -3155
rect 5520 -3190 5560 -3185
rect 5520 -3225 5560 -3220
rect 5520 -3255 5525 -3225
rect 5525 -3255 5555 -3225
rect 5555 -3255 5560 -3225
rect 5520 -3260 5560 -3255
rect 5520 -3295 5560 -3290
rect 5520 -3325 5525 -3295
rect 5525 -3325 5555 -3295
rect 5555 -3325 5560 -3295
rect 5520 -3330 5560 -3325
rect 5520 -3360 5560 -3355
rect 5520 -3390 5525 -3360
rect 5525 -3390 5555 -3360
rect 5555 -3390 5560 -3360
rect 5520 -3395 5560 -3390
rect 5520 -3420 5560 -3415
rect 5520 -3450 5525 -3420
rect 5525 -3450 5555 -3420
rect 5555 -3450 5560 -3420
rect 5520 -3455 5560 -3450
rect 5520 -3485 5560 -3480
rect 5520 -3515 5525 -3485
rect 5525 -3515 5555 -3485
rect 5555 -3515 5560 -3485
rect 5520 -3520 5560 -3515
rect 5520 -3555 5560 -3550
rect 5520 -3585 5525 -3555
rect 5525 -3585 5555 -3555
rect 5555 -3585 5560 -3555
rect 5520 -3590 5560 -3585
rect 5520 -3625 5560 -3620
rect 5520 -3655 5525 -3625
rect 5525 -3655 5555 -3625
rect 5555 -3655 5560 -3625
rect 5520 -3660 5560 -3655
rect 5520 -3695 5560 -3690
rect 5520 -3725 5525 -3695
rect 5525 -3725 5555 -3695
rect 5555 -3725 5560 -3695
rect 5520 -3730 5560 -3725
rect 5520 -3760 5560 -3755
rect 5520 -3790 5525 -3760
rect 5525 -3790 5555 -3760
rect 5555 -3790 5560 -3760
rect 5520 -3795 5560 -3790
rect 5520 -3820 5560 -3815
rect 5520 -3850 5525 -3820
rect 5525 -3850 5555 -3820
rect 5555 -3850 5560 -3820
rect 5520 -3855 5560 -3850
rect 5520 -3885 5560 -3880
rect 5520 -3915 5525 -3885
rect 5525 -3915 5555 -3885
rect 5555 -3915 5560 -3885
rect 5520 -3920 5560 -3915
rect 5520 -3955 5560 -3950
rect 5520 -3985 5525 -3955
rect 5525 -3985 5555 -3955
rect 5555 -3985 5560 -3955
rect 5520 -3990 5560 -3985
rect 5520 -4025 5560 -4020
rect 5520 -4055 5525 -4025
rect 5525 -4055 5555 -4025
rect 5555 -4055 5560 -4025
rect 5520 -4060 5560 -4055
rect 5520 -4095 5560 -4090
rect 5520 -4125 5525 -4095
rect 5525 -4125 5555 -4095
rect 5555 -4125 5560 -4095
rect 5520 -4130 5560 -4125
rect 5520 -4160 5560 -4155
rect 5520 -4190 5525 -4160
rect 5525 -4190 5555 -4160
rect 5555 -4190 5560 -4160
rect 5520 -4195 5560 -4190
rect 5520 -4220 5560 -4215
rect 5520 -4250 5525 -4220
rect 5525 -4250 5555 -4220
rect 5555 -4250 5560 -4220
rect 5520 -4255 5560 -4250
rect 5520 -4285 5560 -4280
rect 5520 -4315 5525 -4285
rect 5525 -4315 5555 -4285
rect 5555 -4315 5560 -4285
rect 5520 -4320 5560 -4315
rect 5520 -4355 5560 -4350
rect 5520 -4385 5525 -4355
rect 5525 -4385 5555 -4355
rect 5555 -4385 5560 -4355
rect 5520 -4390 5560 -4385
rect 5520 -4425 5560 -4420
rect 5520 -4455 5525 -4425
rect 5525 -4455 5555 -4425
rect 5555 -4455 5560 -4425
rect 5520 -4460 5560 -4455
rect 5520 -4495 5560 -4490
rect 5520 -4525 5525 -4495
rect 5525 -4525 5555 -4495
rect 5555 -4525 5560 -4495
rect 5520 -4530 5560 -4525
rect 5520 -4560 5560 -4555
rect 5520 -4590 5525 -4560
rect 5525 -4590 5555 -4560
rect 5555 -4590 5560 -4560
rect 5520 -4595 5560 -4590
<< metal4 >>
rect 2070 19315 32890 19325
rect 2070 19275 2110 19315
rect 2150 19275 6700 19315
rect 6740 19305 32890 19315
rect 6740 19275 31305 19305
rect 2070 19270 31305 19275
rect 31340 19270 31350 19305
rect 31385 19270 31395 19305
rect 31430 19270 31440 19305
rect 31475 19270 31485 19305
rect 31520 19270 31530 19305
rect 31565 19270 31575 19305
rect 31610 19270 31620 19305
rect 31655 19270 31665 19305
rect 31700 19270 31710 19305
rect 31745 19270 31755 19305
rect 31790 19270 31800 19305
rect 31835 19270 31845 19305
rect 31880 19270 31890 19305
rect 31925 19270 31935 19305
rect 31970 19270 31980 19305
rect 32015 19270 32025 19305
rect 32060 19270 32070 19305
rect 32105 19270 32115 19305
rect 32150 19270 32160 19305
rect 32195 19270 32205 19305
rect 32240 19270 32250 19305
rect 32285 19270 32295 19305
rect 32330 19270 32340 19305
rect 32375 19270 32385 19305
rect 32420 19270 32430 19305
rect 32465 19270 32475 19305
rect 32510 19270 32520 19305
rect 32555 19270 32565 19305
rect 32600 19270 32610 19305
rect 32645 19270 32655 19305
rect 32690 19270 32700 19305
rect 32735 19270 32745 19305
rect 32780 19270 32790 19305
rect 32825 19270 32835 19305
rect 32870 19270 32890 19305
rect 2070 19260 32890 19270
rect 2070 19250 31305 19260
rect 2070 19210 2110 19250
rect 2150 19210 6700 19250
rect 6740 19225 31305 19250
rect 31340 19225 31350 19260
rect 31385 19225 31395 19260
rect 31430 19225 31440 19260
rect 31475 19225 31485 19260
rect 31520 19225 31530 19260
rect 31565 19225 31575 19260
rect 31610 19225 31620 19260
rect 31655 19225 31665 19260
rect 31700 19225 31710 19260
rect 31745 19225 31755 19260
rect 31790 19225 31800 19260
rect 31835 19225 31845 19260
rect 31880 19225 31890 19260
rect 31925 19225 31935 19260
rect 31970 19225 31980 19260
rect 32015 19225 32025 19260
rect 32060 19225 32070 19260
rect 32105 19225 32115 19260
rect 32150 19225 32160 19260
rect 32195 19225 32205 19260
rect 32240 19225 32250 19260
rect 32285 19225 32295 19260
rect 32330 19225 32340 19260
rect 32375 19225 32385 19260
rect 32420 19225 32430 19260
rect 32465 19225 32475 19260
rect 32510 19225 32520 19260
rect 32555 19225 32565 19260
rect 32600 19225 32610 19260
rect 32645 19225 32655 19260
rect 32690 19225 32700 19260
rect 32735 19225 32745 19260
rect 32780 19225 32790 19260
rect 32825 19225 32835 19260
rect 32870 19225 32890 19260
rect 6740 19215 32890 19225
rect 6740 19210 31305 19215
rect 2070 19180 31305 19210
rect 31340 19180 31350 19215
rect 31385 19180 31395 19215
rect 31430 19180 31440 19215
rect 31475 19180 31485 19215
rect 31520 19180 31530 19215
rect 31565 19180 31575 19215
rect 31610 19180 31620 19215
rect 31655 19180 31665 19215
rect 31700 19180 31710 19215
rect 31745 19180 31755 19215
rect 31790 19180 31800 19215
rect 31835 19180 31845 19215
rect 31880 19180 31890 19215
rect 31925 19180 31935 19215
rect 31970 19180 31980 19215
rect 32015 19180 32025 19215
rect 32060 19180 32070 19215
rect 32105 19180 32115 19215
rect 32150 19180 32160 19215
rect 32195 19180 32205 19215
rect 32240 19180 32250 19215
rect 32285 19180 32295 19215
rect 32330 19180 32340 19215
rect 32375 19180 32385 19215
rect 32420 19180 32430 19215
rect 32465 19180 32475 19215
rect 32510 19180 32520 19215
rect 32555 19180 32565 19215
rect 32600 19180 32610 19215
rect 32645 19180 32655 19215
rect 32690 19180 32700 19215
rect 32735 19180 32745 19215
rect 32780 19180 32790 19215
rect 32825 19180 32835 19215
rect 32870 19180 32890 19215
rect 2070 19140 2110 19180
rect 2150 19140 6700 19180
rect 6740 19170 32890 19180
rect 6740 19140 31305 19170
rect 2070 19135 31305 19140
rect 31340 19135 31350 19170
rect 31385 19135 31395 19170
rect 31430 19135 31440 19170
rect 31475 19135 31485 19170
rect 31520 19135 31530 19170
rect 31565 19135 31575 19170
rect 31610 19135 31620 19170
rect 31655 19135 31665 19170
rect 31700 19135 31710 19170
rect 31745 19135 31755 19170
rect 31790 19135 31800 19170
rect 31835 19135 31845 19170
rect 31880 19135 31890 19170
rect 31925 19135 31935 19170
rect 31970 19135 31980 19170
rect 32015 19135 32025 19170
rect 32060 19135 32070 19170
rect 32105 19135 32115 19170
rect 32150 19135 32160 19170
rect 32195 19135 32205 19170
rect 32240 19135 32250 19170
rect 32285 19135 32295 19170
rect 32330 19135 32340 19170
rect 32375 19135 32385 19170
rect 32420 19135 32430 19170
rect 32465 19135 32475 19170
rect 32510 19135 32520 19170
rect 32555 19135 32565 19170
rect 32600 19135 32610 19170
rect 32645 19135 32655 19170
rect 32690 19135 32700 19170
rect 32735 19135 32745 19170
rect 32780 19135 32790 19170
rect 32825 19135 32835 19170
rect 32870 19135 32890 19170
rect 2070 19125 32890 19135
rect 2070 19110 31305 19125
rect 2070 19070 2110 19110
rect 2150 19070 6700 19110
rect 6740 19090 31305 19110
rect 31340 19090 31350 19125
rect 31385 19090 31395 19125
rect 31430 19090 31440 19125
rect 31475 19090 31485 19125
rect 31520 19090 31530 19125
rect 31565 19090 31575 19125
rect 31610 19090 31620 19125
rect 31655 19090 31665 19125
rect 31700 19090 31710 19125
rect 31745 19090 31755 19125
rect 31790 19090 31800 19125
rect 31835 19090 31845 19125
rect 31880 19090 31890 19125
rect 31925 19090 31935 19125
rect 31970 19090 31980 19125
rect 32015 19090 32025 19125
rect 32060 19090 32070 19125
rect 32105 19090 32115 19125
rect 32150 19090 32160 19125
rect 32195 19090 32205 19125
rect 32240 19090 32250 19125
rect 32285 19090 32295 19125
rect 32330 19090 32340 19125
rect 32375 19090 32385 19125
rect 32420 19090 32430 19125
rect 32465 19090 32475 19125
rect 32510 19090 32520 19125
rect 32555 19090 32565 19125
rect 32600 19090 32610 19125
rect 32645 19090 32655 19125
rect 32690 19090 32700 19125
rect 32735 19090 32745 19125
rect 32780 19090 32790 19125
rect 32825 19090 32835 19125
rect 32870 19090 32890 19125
rect 6740 19080 32890 19090
rect 6740 19070 31305 19080
rect 2070 19045 31305 19070
rect 31340 19045 31350 19080
rect 31385 19045 31395 19080
rect 31430 19045 31440 19080
rect 31475 19045 31485 19080
rect 31520 19045 31530 19080
rect 31565 19045 31575 19080
rect 31610 19045 31620 19080
rect 31655 19045 31665 19080
rect 31700 19045 31710 19080
rect 31745 19045 31755 19080
rect 31790 19045 31800 19080
rect 31835 19045 31845 19080
rect 31880 19045 31890 19080
rect 31925 19045 31935 19080
rect 31970 19045 31980 19080
rect 32015 19045 32025 19080
rect 32060 19045 32070 19080
rect 32105 19045 32115 19080
rect 32150 19045 32160 19080
rect 32195 19045 32205 19080
rect 32240 19045 32250 19080
rect 32285 19045 32295 19080
rect 32330 19045 32340 19080
rect 32375 19045 32385 19080
rect 32420 19045 32430 19080
rect 32465 19045 32475 19080
rect 32510 19045 32520 19080
rect 32555 19045 32565 19080
rect 32600 19045 32610 19080
rect 32645 19045 32655 19080
rect 32690 19045 32700 19080
rect 32735 19045 32745 19080
rect 32780 19045 32790 19080
rect 32825 19045 32835 19080
rect 32870 19045 32890 19080
rect 2070 19040 32890 19045
rect 2070 19000 2110 19040
rect 2150 19000 6700 19040
rect 6740 19035 32890 19040
rect 6740 19000 31305 19035
rect 31340 19000 31350 19035
rect 31385 19000 31395 19035
rect 31430 19000 31440 19035
rect 31475 19000 31485 19035
rect 31520 19000 31530 19035
rect 31565 19000 31575 19035
rect 31610 19000 31620 19035
rect 31655 19000 31665 19035
rect 31700 19000 31710 19035
rect 31745 19000 31755 19035
rect 31790 19000 31800 19035
rect 31835 19000 31845 19035
rect 31880 19000 31890 19035
rect 31925 19000 31935 19035
rect 31970 19000 31980 19035
rect 32015 19000 32025 19035
rect 32060 19000 32070 19035
rect 32105 19000 32115 19035
rect 32150 19000 32160 19035
rect 32195 19000 32205 19035
rect 32240 19000 32250 19035
rect 32285 19000 32295 19035
rect 32330 19000 32340 19035
rect 32375 19000 32385 19035
rect 32420 19000 32430 19035
rect 32465 19000 32475 19035
rect 32510 19000 32520 19035
rect 32555 19000 32565 19035
rect 32600 19000 32610 19035
rect 32645 19000 32655 19035
rect 32690 19000 32700 19035
rect 32735 19000 32745 19035
rect 32780 19000 32790 19035
rect 32825 19000 32835 19035
rect 32870 19000 32890 19035
rect 2070 18990 32890 19000
rect 2070 18975 31305 18990
rect 2070 18935 2110 18975
rect 2150 18935 6700 18975
rect 6740 18955 31305 18975
rect 31340 18955 31350 18990
rect 31385 18955 31395 18990
rect 31430 18955 31440 18990
rect 31475 18955 31485 18990
rect 31520 18955 31530 18990
rect 31565 18955 31575 18990
rect 31610 18955 31620 18990
rect 31655 18955 31665 18990
rect 31700 18955 31710 18990
rect 31745 18955 31755 18990
rect 31790 18955 31800 18990
rect 31835 18955 31845 18990
rect 31880 18955 31890 18990
rect 31925 18955 31935 18990
rect 31970 18955 31980 18990
rect 32015 18955 32025 18990
rect 32060 18955 32070 18990
rect 32105 18955 32115 18990
rect 32150 18955 32160 18990
rect 32195 18955 32205 18990
rect 32240 18955 32250 18990
rect 32285 18955 32295 18990
rect 32330 18955 32340 18990
rect 32375 18955 32385 18990
rect 32420 18955 32430 18990
rect 32465 18955 32475 18990
rect 32510 18955 32520 18990
rect 32555 18955 32565 18990
rect 32600 18955 32610 18990
rect 32645 18955 32655 18990
rect 32690 18955 32700 18990
rect 32735 18955 32745 18990
rect 32780 18955 32790 18990
rect 32825 18955 32835 18990
rect 32870 18955 32890 18990
rect 6740 18945 32890 18955
rect 6740 18935 31305 18945
rect 2070 18915 31305 18935
rect 2070 18875 2110 18915
rect 2150 18875 6700 18915
rect 6740 18910 31305 18915
rect 31340 18910 31350 18945
rect 31385 18910 31395 18945
rect 31430 18910 31440 18945
rect 31475 18910 31485 18945
rect 31520 18910 31530 18945
rect 31565 18910 31575 18945
rect 31610 18910 31620 18945
rect 31655 18910 31665 18945
rect 31700 18910 31710 18945
rect 31745 18910 31755 18945
rect 31790 18910 31800 18945
rect 31835 18910 31845 18945
rect 31880 18910 31890 18945
rect 31925 18910 31935 18945
rect 31970 18910 31980 18945
rect 32015 18910 32025 18945
rect 32060 18910 32070 18945
rect 32105 18910 32115 18945
rect 32150 18910 32160 18945
rect 32195 18910 32205 18945
rect 32240 18910 32250 18945
rect 32285 18910 32295 18945
rect 32330 18910 32340 18945
rect 32375 18910 32385 18945
rect 32420 18910 32430 18945
rect 32465 18910 32475 18945
rect 32510 18910 32520 18945
rect 32555 18910 32565 18945
rect 32600 18910 32610 18945
rect 32645 18910 32655 18945
rect 32690 18910 32700 18945
rect 32735 18910 32745 18945
rect 32780 18910 32790 18945
rect 32825 18910 32835 18945
rect 32870 18910 32890 18945
rect 6740 18900 32890 18910
rect 6740 18875 31305 18900
rect 2070 18865 31305 18875
rect 31340 18865 31350 18900
rect 31385 18865 31395 18900
rect 31430 18865 31440 18900
rect 31475 18865 31485 18900
rect 31520 18865 31530 18900
rect 31565 18865 31575 18900
rect 31610 18865 31620 18900
rect 31655 18865 31665 18900
rect 31700 18865 31710 18900
rect 31745 18865 31755 18900
rect 31790 18865 31800 18900
rect 31835 18865 31845 18900
rect 31880 18865 31890 18900
rect 31925 18865 31935 18900
rect 31970 18865 31980 18900
rect 32015 18865 32025 18900
rect 32060 18865 32070 18900
rect 32105 18865 32115 18900
rect 32150 18865 32160 18900
rect 32195 18865 32205 18900
rect 32240 18865 32250 18900
rect 32285 18865 32295 18900
rect 32330 18865 32340 18900
rect 32375 18865 32385 18900
rect 32420 18865 32430 18900
rect 32465 18865 32475 18900
rect 32510 18865 32520 18900
rect 32555 18865 32565 18900
rect 32600 18865 32610 18900
rect 32645 18865 32655 18900
rect 32690 18865 32700 18900
rect 32735 18865 32745 18900
rect 32780 18865 32790 18900
rect 32825 18865 32835 18900
rect 32870 18865 32890 18900
rect 2070 18855 32890 18865
rect 2070 18850 31305 18855
rect 2070 18810 2110 18850
rect 2150 18810 6700 18850
rect 6740 18820 31305 18850
rect 31340 18820 31350 18855
rect 31385 18820 31395 18855
rect 31430 18820 31440 18855
rect 31475 18820 31485 18855
rect 31520 18820 31530 18855
rect 31565 18820 31575 18855
rect 31610 18820 31620 18855
rect 31655 18820 31665 18855
rect 31700 18820 31710 18855
rect 31745 18820 31755 18855
rect 31790 18820 31800 18855
rect 31835 18820 31845 18855
rect 31880 18820 31890 18855
rect 31925 18820 31935 18855
rect 31970 18820 31980 18855
rect 32015 18820 32025 18855
rect 32060 18820 32070 18855
rect 32105 18820 32115 18855
rect 32150 18820 32160 18855
rect 32195 18820 32205 18855
rect 32240 18820 32250 18855
rect 32285 18820 32295 18855
rect 32330 18820 32340 18855
rect 32375 18820 32385 18855
rect 32420 18820 32430 18855
rect 32465 18820 32475 18855
rect 32510 18820 32520 18855
rect 32555 18820 32565 18855
rect 32600 18820 32610 18855
rect 32645 18820 32655 18855
rect 32690 18820 32700 18855
rect 32735 18820 32745 18855
rect 32780 18820 32790 18855
rect 32825 18820 32835 18855
rect 32870 18820 32890 18855
rect 6740 18810 32890 18820
rect 2070 18780 31305 18810
rect 2070 18740 2110 18780
rect 2150 18740 6700 18780
rect 6740 18775 31305 18780
rect 31340 18775 31350 18810
rect 31385 18775 31395 18810
rect 31430 18775 31440 18810
rect 31475 18775 31485 18810
rect 31520 18775 31530 18810
rect 31565 18775 31575 18810
rect 31610 18775 31620 18810
rect 31655 18775 31665 18810
rect 31700 18775 31710 18810
rect 31745 18775 31755 18810
rect 31790 18775 31800 18810
rect 31835 18775 31845 18810
rect 31880 18775 31890 18810
rect 31925 18775 31935 18810
rect 31970 18775 31980 18810
rect 32015 18775 32025 18810
rect 32060 18775 32070 18810
rect 32105 18775 32115 18810
rect 32150 18775 32160 18810
rect 32195 18775 32205 18810
rect 32240 18775 32250 18810
rect 32285 18775 32295 18810
rect 32330 18775 32340 18810
rect 32375 18775 32385 18810
rect 32420 18775 32430 18810
rect 32465 18775 32475 18810
rect 32510 18775 32520 18810
rect 32555 18775 32565 18810
rect 32600 18775 32610 18810
rect 32645 18775 32655 18810
rect 32690 18775 32700 18810
rect 32735 18775 32745 18810
rect 32780 18775 32790 18810
rect 32825 18775 32835 18810
rect 32870 18775 32890 18810
rect 6740 18765 32890 18775
rect 6740 18740 31305 18765
rect 2070 18730 31305 18740
rect 31340 18730 31350 18765
rect 31385 18730 31395 18765
rect 31430 18730 31440 18765
rect 31475 18730 31485 18765
rect 31520 18730 31530 18765
rect 31565 18730 31575 18765
rect 31610 18730 31620 18765
rect 31655 18730 31665 18765
rect 31700 18730 31710 18765
rect 31745 18730 31755 18765
rect 31790 18730 31800 18765
rect 31835 18730 31845 18765
rect 31880 18730 31890 18765
rect 31925 18730 31935 18765
rect 31970 18730 31980 18765
rect 32015 18730 32025 18765
rect 32060 18730 32070 18765
rect 32105 18730 32115 18765
rect 32150 18730 32160 18765
rect 32195 18730 32205 18765
rect 32240 18730 32250 18765
rect 32285 18730 32295 18765
rect 32330 18730 32340 18765
rect 32375 18730 32385 18765
rect 32420 18730 32430 18765
rect 32465 18730 32475 18765
rect 32510 18730 32520 18765
rect 32555 18730 32565 18765
rect 32600 18730 32610 18765
rect 32645 18730 32655 18765
rect 32690 18730 32700 18765
rect 32735 18730 32745 18765
rect 32780 18730 32790 18765
rect 32825 18730 32835 18765
rect 32870 18730 32890 18765
rect 2070 18720 32890 18730
rect 2070 18710 31305 18720
rect 2070 18670 2110 18710
rect 2150 18670 6700 18710
rect 6740 18685 31305 18710
rect 31340 18685 31350 18720
rect 31385 18685 31395 18720
rect 31430 18685 31440 18720
rect 31475 18685 31485 18720
rect 31520 18685 31530 18720
rect 31565 18685 31575 18720
rect 31610 18685 31620 18720
rect 31655 18685 31665 18720
rect 31700 18685 31710 18720
rect 31745 18685 31755 18720
rect 31790 18685 31800 18720
rect 31835 18685 31845 18720
rect 31880 18685 31890 18720
rect 31925 18685 31935 18720
rect 31970 18685 31980 18720
rect 32015 18685 32025 18720
rect 32060 18685 32070 18720
rect 32105 18685 32115 18720
rect 32150 18685 32160 18720
rect 32195 18685 32205 18720
rect 32240 18685 32250 18720
rect 32285 18685 32295 18720
rect 32330 18685 32340 18720
rect 32375 18685 32385 18720
rect 32420 18685 32430 18720
rect 32465 18685 32475 18720
rect 32510 18685 32520 18720
rect 32555 18685 32565 18720
rect 32600 18685 32610 18720
rect 32645 18685 32655 18720
rect 32690 18685 32700 18720
rect 32735 18685 32745 18720
rect 32780 18685 32790 18720
rect 32825 18685 32835 18720
rect 32870 18685 32890 18720
rect 6740 18675 32890 18685
rect 6740 18670 31305 18675
rect 2070 18640 31305 18670
rect 31340 18640 31350 18675
rect 31385 18640 31395 18675
rect 31430 18640 31440 18675
rect 31475 18640 31485 18675
rect 31520 18640 31530 18675
rect 31565 18640 31575 18675
rect 31610 18640 31620 18675
rect 31655 18640 31665 18675
rect 31700 18640 31710 18675
rect 31745 18640 31755 18675
rect 31790 18640 31800 18675
rect 31835 18640 31845 18675
rect 31880 18640 31890 18675
rect 31925 18640 31935 18675
rect 31970 18640 31980 18675
rect 32015 18640 32025 18675
rect 32060 18640 32070 18675
rect 32105 18640 32115 18675
rect 32150 18640 32160 18675
rect 32195 18640 32205 18675
rect 32240 18640 32250 18675
rect 32285 18640 32295 18675
rect 32330 18640 32340 18675
rect 32375 18640 32385 18675
rect 32420 18640 32430 18675
rect 32465 18640 32475 18675
rect 32510 18640 32520 18675
rect 32555 18640 32565 18675
rect 32600 18640 32610 18675
rect 32645 18640 32655 18675
rect 32690 18640 32700 18675
rect 32735 18640 32745 18675
rect 32780 18640 32790 18675
rect 32825 18640 32835 18675
rect 32870 18640 32890 18675
rect 2070 18600 2110 18640
rect 2150 18600 6700 18640
rect 6740 18630 32890 18640
rect 6740 18600 31305 18630
rect 2070 18595 31305 18600
rect 31340 18595 31350 18630
rect 31385 18595 31395 18630
rect 31430 18595 31440 18630
rect 31475 18595 31485 18630
rect 31520 18595 31530 18630
rect 31565 18595 31575 18630
rect 31610 18595 31620 18630
rect 31655 18595 31665 18630
rect 31700 18595 31710 18630
rect 31745 18595 31755 18630
rect 31790 18595 31800 18630
rect 31835 18595 31845 18630
rect 31880 18595 31890 18630
rect 31925 18595 31935 18630
rect 31970 18595 31980 18630
rect 32015 18595 32025 18630
rect 32060 18595 32070 18630
rect 32105 18595 32115 18630
rect 32150 18595 32160 18630
rect 32195 18595 32205 18630
rect 32240 18595 32250 18630
rect 32285 18595 32295 18630
rect 32330 18595 32340 18630
rect 32375 18595 32385 18630
rect 32420 18595 32430 18630
rect 32465 18595 32475 18630
rect 32510 18595 32520 18630
rect 32555 18595 32565 18630
rect 32600 18595 32610 18630
rect 32645 18595 32655 18630
rect 32690 18595 32700 18630
rect 32735 18595 32745 18630
rect 32780 18595 32790 18630
rect 32825 18595 32835 18630
rect 32870 18595 32890 18630
rect 2070 18585 32890 18595
rect 2070 18575 31305 18585
rect 2070 18535 2110 18575
rect 2150 18535 6700 18575
rect 6740 18550 31305 18575
rect 31340 18550 31350 18585
rect 31385 18550 31395 18585
rect 31430 18550 31440 18585
rect 31475 18550 31485 18585
rect 31520 18550 31530 18585
rect 31565 18550 31575 18585
rect 31610 18550 31620 18585
rect 31655 18550 31665 18585
rect 31700 18550 31710 18585
rect 31745 18550 31755 18585
rect 31790 18550 31800 18585
rect 31835 18550 31845 18585
rect 31880 18550 31890 18585
rect 31925 18550 31935 18585
rect 31970 18550 31980 18585
rect 32015 18550 32025 18585
rect 32060 18550 32070 18585
rect 32105 18550 32115 18585
rect 32150 18550 32160 18585
rect 32195 18550 32205 18585
rect 32240 18550 32250 18585
rect 32285 18550 32295 18585
rect 32330 18550 32340 18585
rect 32375 18550 32385 18585
rect 32420 18550 32430 18585
rect 32465 18550 32475 18585
rect 32510 18550 32520 18585
rect 32555 18550 32565 18585
rect 32600 18550 32610 18585
rect 32645 18550 32655 18585
rect 32690 18550 32700 18585
rect 32735 18550 32745 18585
rect 32780 18550 32790 18585
rect 32825 18550 32835 18585
rect 32870 18550 32890 18585
rect 6740 18540 32890 18550
rect 6740 18535 31305 18540
rect 2070 18515 31305 18535
rect 2070 18475 2110 18515
rect 2150 18475 6700 18515
rect 6740 18505 31305 18515
rect 31340 18505 31350 18540
rect 31385 18505 31395 18540
rect 31430 18505 31440 18540
rect 31475 18505 31485 18540
rect 31520 18505 31530 18540
rect 31565 18505 31575 18540
rect 31610 18505 31620 18540
rect 31655 18505 31665 18540
rect 31700 18505 31710 18540
rect 31745 18505 31755 18540
rect 31790 18505 31800 18540
rect 31835 18505 31845 18540
rect 31880 18505 31890 18540
rect 31925 18505 31935 18540
rect 31970 18505 31980 18540
rect 32015 18505 32025 18540
rect 32060 18505 32070 18540
rect 32105 18505 32115 18540
rect 32150 18505 32160 18540
rect 32195 18505 32205 18540
rect 32240 18505 32250 18540
rect 32285 18505 32295 18540
rect 32330 18505 32340 18540
rect 32375 18505 32385 18540
rect 32420 18505 32430 18540
rect 32465 18505 32475 18540
rect 32510 18505 32520 18540
rect 32555 18505 32565 18540
rect 32600 18505 32610 18540
rect 32645 18505 32655 18540
rect 32690 18505 32700 18540
rect 32735 18505 32745 18540
rect 32780 18505 32790 18540
rect 32825 18505 32835 18540
rect 32870 18505 32890 18540
rect 6740 18495 32890 18505
rect 6740 18475 31305 18495
rect 2070 18460 31305 18475
rect 31340 18460 31350 18495
rect 31385 18460 31395 18495
rect 31430 18460 31440 18495
rect 31475 18460 31485 18495
rect 31520 18460 31530 18495
rect 31565 18460 31575 18495
rect 31610 18460 31620 18495
rect 31655 18460 31665 18495
rect 31700 18460 31710 18495
rect 31745 18460 31755 18495
rect 31790 18460 31800 18495
rect 31835 18460 31845 18495
rect 31880 18460 31890 18495
rect 31925 18460 31935 18495
rect 31970 18460 31980 18495
rect 32015 18460 32025 18495
rect 32060 18460 32070 18495
rect 32105 18460 32115 18495
rect 32150 18460 32160 18495
rect 32195 18460 32205 18495
rect 32240 18460 32250 18495
rect 32285 18460 32295 18495
rect 32330 18460 32340 18495
rect 32375 18460 32385 18495
rect 32420 18460 32430 18495
rect 32465 18460 32475 18495
rect 32510 18460 32520 18495
rect 32555 18460 32565 18495
rect 32600 18460 32610 18495
rect 32645 18460 32655 18495
rect 32690 18460 32700 18495
rect 32735 18460 32745 18495
rect 32780 18460 32790 18495
rect 32825 18460 32835 18495
rect 32870 18460 32890 18495
rect 2070 18450 32890 18460
rect 2070 18410 2110 18450
rect 2150 18410 6700 18450
rect 6740 18415 31305 18450
rect 31340 18415 31350 18450
rect 31385 18415 31395 18450
rect 31430 18415 31440 18450
rect 31475 18415 31485 18450
rect 31520 18415 31530 18450
rect 31565 18415 31575 18450
rect 31610 18415 31620 18450
rect 31655 18415 31665 18450
rect 31700 18415 31710 18450
rect 31745 18415 31755 18450
rect 31790 18415 31800 18450
rect 31835 18415 31845 18450
rect 31880 18415 31890 18450
rect 31925 18415 31935 18450
rect 31970 18415 31980 18450
rect 32015 18415 32025 18450
rect 32060 18415 32070 18450
rect 32105 18415 32115 18450
rect 32150 18415 32160 18450
rect 32195 18415 32205 18450
rect 32240 18415 32250 18450
rect 32285 18415 32295 18450
rect 32330 18415 32340 18450
rect 32375 18415 32385 18450
rect 32420 18415 32430 18450
rect 32465 18415 32475 18450
rect 32510 18415 32520 18450
rect 32555 18415 32565 18450
rect 32600 18415 32610 18450
rect 32645 18415 32655 18450
rect 32690 18415 32700 18450
rect 32735 18415 32745 18450
rect 32780 18415 32790 18450
rect 32825 18415 32835 18450
rect 32870 18415 32890 18450
rect 6740 18410 32890 18415
rect 2070 18405 32890 18410
rect 2070 18380 31305 18405
rect 2070 18340 2110 18380
rect 2150 18340 6700 18380
rect 6740 18370 31305 18380
rect 31340 18370 31350 18405
rect 31385 18370 31395 18405
rect 31430 18370 31440 18405
rect 31475 18370 31485 18405
rect 31520 18370 31530 18405
rect 31565 18370 31575 18405
rect 31610 18370 31620 18405
rect 31655 18370 31665 18405
rect 31700 18370 31710 18405
rect 31745 18370 31755 18405
rect 31790 18370 31800 18405
rect 31835 18370 31845 18405
rect 31880 18370 31890 18405
rect 31925 18370 31935 18405
rect 31970 18370 31980 18405
rect 32015 18370 32025 18405
rect 32060 18370 32070 18405
rect 32105 18370 32115 18405
rect 32150 18370 32160 18405
rect 32195 18370 32205 18405
rect 32240 18370 32250 18405
rect 32285 18370 32295 18405
rect 32330 18370 32340 18405
rect 32375 18370 32385 18405
rect 32420 18370 32430 18405
rect 32465 18370 32475 18405
rect 32510 18370 32520 18405
rect 32555 18370 32565 18405
rect 32600 18370 32610 18405
rect 32645 18370 32655 18405
rect 32690 18370 32700 18405
rect 32735 18370 32745 18405
rect 32780 18370 32790 18405
rect 32825 18370 32835 18405
rect 32870 18370 32890 18405
rect 6740 18360 32890 18370
rect 6740 18340 31305 18360
rect 2070 18325 31305 18340
rect 31340 18325 31350 18360
rect 31385 18325 31395 18360
rect 31430 18325 31440 18360
rect 31475 18325 31485 18360
rect 31520 18325 31530 18360
rect 31565 18325 31575 18360
rect 31610 18325 31620 18360
rect 31655 18325 31665 18360
rect 31700 18325 31710 18360
rect 31745 18325 31755 18360
rect 31790 18325 31800 18360
rect 31835 18325 31845 18360
rect 31880 18325 31890 18360
rect 31925 18325 31935 18360
rect 31970 18325 31980 18360
rect 32015 18325 32025 18360
rect 32060 18325 32070 18360
rect 32105 18325 32115 18360
rect 32150 18325 32160 18360
rect 32195 18325 32205 18360
rect 32240 18325 32250 18360
rect 32285 18325 32295 18360
rect 32330 18325 32340 18360
rect 32375 18325 32385 18360
rect 32420 18325 32430 18360
rect 32465 18325 32475 18360
rect 32510 18325 32520 18360
rect 32555 18325 32565 18360
rect 32600 18325 32610 18360
rect 32645 18325 32655 18360
rect 32690 18325 32700 18360
rect 32735 18325 32745 18360
rect 32780 18325 32790 18360
rect 32825 18325 32835 18360
rect 32870 18325 32890 18360
rect 2070 18315 32890 18325
rect 2070 18310 31305 18315
rect 2070 18270 2110 18310
rect 2150 18270 6700 18310
rect 6740 18280 31305 18310
rect 31340 18280 31350 18315
rect 31385 18280 31395 18315
rect 31430 18280 31440 18315
rect 31475 18280 31485 18315
rect 31520 18280 31530 18315
rect 31565 18280 31575 18315
rect 31610 18280 31620 18315
rect 31655 18280 31665 18315
rect 31700 18280 31710 18315
rect 31745 18280 31755 18315
rect 31790 18280 31800 18315
rect 31835 18280 31845 18315
rect 31880 18280 31890 18315
rect 31925 18280 31935 18315
rect 31970 18280 31980 18315
rect 32015 18280 32025 18315
rect 32060 18280 32070 18315
rect 32105 18280 32115 18315
rect 32150 18280 32160 18315
rect 32195 18280 32205 18315
rect 32240 18280 32250 18315
rect 32285 18280 32295 18315
rect 32330 18280 32340 18315
rect 32375 18280 32385 18315
rect 32420 18280 32430 18315
rect 32465 18280 32475 18315
rect 32510 18280 32520 18315
rect 32555 18280 32565 18315
rect 32600 18280 32610 18315
rect 32645 18280 32655 18315
rect 32690 18280 32700 18315
rect 32735 18280 32745 18315
rect 32780 18280 32790 18315
rect 32825 18280 32835 18315
rect 32870 18280 32890 18315
rect 6740 18270 32890 18280
rect 2070 18240 31305 18270
rect 2070 18200 2110 18240
rect 2150 18200 6700 18240
rect 6740 18235 31305 18240
rect 31340 18235 31350 18270
rect 31385 18235 31395 18270
rect 31430 18235 31440 18270
rect 31475 18235 31485 18270
rect 31520 18235 31530 18270
rect 31565 18235 31575 18270
rect 31610 18235 31620 18270
rect 31655 18235 31665 18270
rect 31700 18235 31710 18270
rect 31745 18235 31755 18270
rect 31790 18235 31800 18270
rect 31835 18235 31845 18270
rect 31880 18235 31890 18270
rect 31925 18235 31935 18270
rect 31970 18235 31980 18270
rect 32015 18235 32025 18270
rect 32060 18235 32070 18270
rect 32105 18235 32115 18270
rect 32150 18235 32160 18270
rect 32195 18235 32205 18270
rect 32240 18235 32250 18270
rect 32285 18235 32295 18270
rect 32330 18235 32340 18270
rect 32375 18235 32385 18270
rect 32420 18235 32430 18270
rect 32465 18235 32475 18270
rect 32510 18235 32520 18270
rect 32555 18235 32565 18270
rect 32600 18235 32610 18270
rect 32645 18235 32655 18270
rect 32690 18235 32700 18270
rect 32735 18235 32745 18270
rect 32780 18235 32790 18270
rect 32825 18235 32835 18270
rect 32870 18235 32890 18270
rect 6740 18225 32890 18235
rect 6740 18200 31305 18225
rect 2070 18190 31305 18200
rect 31340 18190 31350 18225
rect 31385 18190 31395 18225
rect 31430 18190 31440 18225
rect 31475 18190 31485 18225
rect 31520 18190 31530 18225
rect 31565 18190 31575 18225
rect 31610 18190 31620 18225
rect 31655 18190 31665 18225
rect 31700 18190 31710 18225
rect 31745 18190 31755 18225
rect 31790 18190 31800 18225
rect 31835 18190 31845 18225
rect 31880 18190 31890 18225
rect 31925 18190 31935 18225
rect 31970 18190 31980 18225
rect 32015 18190 32025 18225
rect 32060 18190 32070 18225
rect 32105 18190 32115 18225
rect 32150 18190 32160 18225
rect 32195 18190 32205 18225
rect 32240 18190 32250 18225
rect 32285 18190 32295 18225
rect 32330 18190 32340 18225
rect 32375 18190 32385 18225
rect 32420 18190 32430 18225
rect 32465 18190 32475 18225
rect 32510 18190 32520 18225
rect 32555 18190 32565 18225
rect 32600 18190 32610 18225
rect 32645 18190 32655 18225
rect 32690 18190 32700 18225
rect 32735 18190 32745 18225
rect 32780 18190 32790 18225
rect 32825 18190 32835 18225
rect 32870 18190 32890 18225
rect 2070 18180 32890 18190
rect 2070 18175 31305 18180
rect 2070 18135 2110 18175
rect 2150 18135 6700 18175
rect 6740 18145 31305 18175
rect 31340 18145 31350 18180
rect 31385 18145 31395 18180
rect 31430 18145 31440 18180
rect 31475 18145 31485 18180
rect 31520 18145 31530 18180
rect 31565 18145 31575 18180
rect 31610 18145 31620 18180
rect 31655 18145 31665 18180
rect 31700 18145 31710 18180
rect 31745 18145 31755 18180
rect 31790 18145 31800 18180
rect 31835 18145 31845 18180
rect 31880 18145 31890 18180
rect 31925 18145 31935 18180
rect 31970 18145 31980 18180
rect 32015 18145 32025 18180
rect 32060 18145 32070 18180
rect 32105 18145 32115 18180
rect 32150 18145 32160 18180
rect 32195 18145 32205 18180
rect 32240 18145 32250 18180
rect 32285 18145 32295 18180
rect 32330 18145 32340 18180
rect 32375 18145 32385 18180
rect 32420 18145 32430 18180
rect 32465 18145 32475 18180
rect 32510 18145 32520 18180
rect 32555 18145 32565 18180
rect 32600 18145 32610 18180
rect 32645 18145 32655 18180
rect 32690 18145 32700 18180
rect 32735 18145 32745 18180
rect 32780 18145 32790 18180
rect 32825 18145 32835 18180
rect 32870 18145 32890 18180
rect 6740 18135 32890 18145
rect 2070 18115 31305 18135
rect 2070 18075 2110 18115
rect 2150 18075 6700 18115
rect 6740 18100 31305 18115
rect 31340 18100 31350 18135
rect 31385 18100 31395 18135
rect 31430 18100 31440 18135
rect 31475 18100 31485 18135
rect 31520 18100 31530 18135
rect 31565 18100 31575 18135
rect 31610 18100 31620 18135
rect 31655 18100 31665 18135
rect 31700 18100 31710 18135
rect 31745 18100 31755 18135
rect 31790 18100 31800 18135
rect 31835 18100 31845 18135
rect 31880 18100 31890 18135
rect 31925 18100 31935 18135
rect 31970 18100 31980 18135
rect 32015 18100 32025 18135
rect 32060 18100 32070 18135
rect 32105 18100 32115 18135
rect 32150 18100 32160 18135
rect 32195 18100 32205 18135
rect 32240 18100 32250 18135
rect 32285 18100 32295 18135
rect 32330 18100 32340 18135
rect 32375 18100 32385 18135
rect 32420 18100 32430 18135
rect 32465 18100 32475 18135
rect 32510 18100 32520 18135
rect 32555 18100 32565 18135
rect 32600 18100 32610 18135
rect 32645 18100 32655 18135
rect 32690 18100 32700 18135
rect 32735 18100 32745 18135
rect 32780 18100 32790 18135
rect 32825 18100 32835 18135
rect 32870 18100 32890 18135
rect 6740 18090 32890 18100
rect 6740 18075 31305 18090
rect 2070 18055 31305 18075
rect 31340 18055 31350 18090
rect 31385 18055 31395 18090
rect 31430 18055 31440 18090
rect 31475 18055 31485 18090
rect 31520 18055 31530 18090
rect 31565 18055 31575 18090
rect 31610 18055 31620 18090
rect 31655 18055 31665 18090
rect 31700 18055 31710 18090
rect 31745 18055 31755 18090
rect 31790 18055 31800 18090
rect 31835 18055 31845 18090
rect 31880 18055 31890 18090
rect 31925 18055 31935 18090
rect 31970 18055 31980 18090
rect 32015 18055 32025 18090
rect 32060 18055 32070 18090
rect 32105 18055 32115 18090
rect 32150 18055 32160 18090
rect 32195 18055 32205 18090
rect 32240 18055 32250 18090
rect 32285 18055 32295 18090
rect 32330 18055 32340 18090
rect 32375 18055 32385 18090
rect 32420 18055 32430 18090
rect 32465 18055 32475 18090
rect 32510 18055 32520 18090
rect 32555 18055 32565 18090
rect 32600 18055 32610 18090
rect 32645 18055 32655 18090
rect 32690 18055 32700 18090
rect 32735 18055 32745 18090
rect 32780 18055 32790 18090
rect 32825 18055 32835 18090
rect 32870 18055 32890 18090
rect 2070 18050 32890 18055
rect 2070 18010 2110 18050
rect 2150 18010 6700 18050
rect 6740 18045 32890 18050
rect 6740 18010 31305 18045
rect 31340 18010 31350 18045
rect 31385 18010 31395 18045
rect 31430 18010 31440 18045
rect 31475 18010 31485 18045
rect 31520 18010 31530 18045
rect 31565 18010 31575 18045
rect 31610 18010 31620 18045
rect 31655 18010 31665 18045
rect 31700 18010 31710 18045
rect 31745 18010 31755 18045
rect 31790 18010 31800 18045
rect 31835 18010 31845 18045
rect 31880 18010 31890 18045
rect 31925 18010 31935 18045
rect 31970 18010 31980 18045
rect 32015 18010 32025 18045
rect 32060 18010 32070 18045
rect 32105 18010 32115 18045
rect 32150 18010 32160 18045
rect 32195 18010 32205 18045
rect 32240 18010 32250 18045
rect 32285 18010 32295 18045
rect 32330 18010 32340 18045
rect 32375 18010 32385 18045
rect 32420 18010 32430 18045
rect 32465 18010 32475 18045
rect 32510 18010 32520 18045
rect 32555 18010 32565 18045
rect 32600 18010 32610 18045
rect 32645 18010 32655 18045
rect 32690 18010 32700 18045
rect 32735 18010 32745 18045
rect 32780 18010 32790 18045
rect 32825 18010 32835 18045
rect 32870 18010 32890 18045
rect 2070 18000 32890 18010
rect 2070 17980 31305 18000
rect 2070 17940 2110 17980
rect 2150 17940 6700 17980
rect 6740 17965 31305 17980
rect 31340 17965 31350 18000
rect 31385 17965 31395 18000
rect 31430 17965 31440 18000
rect 31475 17965 31485 18000
rect 31520 17965 31530 18000
rect 31565 17965 31575 18000
rect 31610 17965 31620 18000
rect 31655 17965 31665 18000
rect 31700 17965 31710 18000
rect 31745 17965 31755 18000
rect 31790 17965 31800 18000
rect 31835 17965 31845 18000
rect 31880 17965 31890 18000
rect 31925 17965 31935 18000
rect 31970 17965 31980 18000
rect 32015 17965 32025 18000
rect 32060 17965 32070 18000
rect 32105 17965 32115 18000
rect 32150 17965 32160 18000
rect 32195 17965 32205 18000
rect 32240 17965 32250 18000
rect 32285 17965 32295 18000
rect 32330 17965 32340 18000
rect 32375 17965 32385 18000
rect 32420 17965 32430 18000
rect 32465 17965 32475 18000
rect 32510 17965 32520 18000
rect 32555 17965 32565 18000
rect 32600 17965 32610 18000
rect 32645 17965 32655 18000
rect 32690 17965 32700 18000
rect 32735 17965 32745 18000
rect 32780 17965 32790 18000
rect 32825 17965 32835 18000
rect 32870 17965 32890 18000
rect 6740 17955 32890 17965
rect 6740 17940 31305 17955
rect 2070 17920 31305 17940
rect 31340 17920 31350 17955
rect 31385 17920 31395 17955
rect 31430 17920 31440 17955
rect 31475 17920 31485 17955
rect 31520 17920 31530 17955
rect 31565 17920 31575 17955
rect 31610 17920 31620 17955
rect 31655 17920 31665 17955
rect 31700 17920 31710 17955
rect 31745 17920 31755 17955
rect 31790 17920 31800 17955
rect 31835 17920 31845 17955
rect 31880 17920 31890 17955
rect 31925 17920 31935 17955
rect 31970 17920 31980 17955
rect 32015 17920 32025 17955
rect 32060 17920 32070 17955
rect 32105 17920 32115 17955
rect 32150 17920 32160 17955
rect 32195 17920 32205 17955
rect 32240 17920 32250 17955
rect 32285 17920 32295 17955
rect 32330 17920 32340 17955
rect 32375 17920 32385 17955
rect 32420 17920 32430 17955
rect 32465 17920 32475 17955
rect 32510 17920 32520 17955
rect 32555 17920 32565 17955
rect 32600 17920 32610 17955
rect 32645 17920 32655 17955
rect 32690 17920 32700 17955
rect 32735 17920 32745 17955
rect 32780 17920 32790 17955
rect 32825 17920 32835 17955
rect 32870 17920 32890 17955
rect 2070 17910 32890 17920
rect 2070 17870 2110 17910
rect 2150 17870 6700 17910
rect 6740 17875 31305 17910
rect 31340 17875 31350 17910
rect 31385 17875 31395 17910
rect 31430 17875 31440 17910
rect 31475 17875 31485 17910
rect 31520 17875 31530 17910
rect 31565 17875 31575 17910
rect 31610 17875 31620 17910
rect 31655 17875 31665 17910
rect 31700 17875 31710 17910
rect 31745 17875 31755 17910
rect 31790 17875 31800 17910
rect 31835 17875 31845 17910
rect 31880 17875 31890 17910
rect 31925 17875 31935 17910
rect 31970 17875 31980 17910
rect 32015 17875 32025 17910
rect 32060 17875 32070 17910
rect 32105 17875 32115 17910
rect 32150 17875 32160 17910
rect 32195 17875 32205 17910
rect 32240 17875 32250 17910
rect 32285 17875 32295 17910
rect 32330 17875 32340 17910
rect 32375 17875 32385 17910
rect 32420 17875 32430 17910
rect 32465 17875 32475 17910
rect 32510 17875 32520 17910
rect 32555 17875 32565 17910
rect 32600 17875 32610 17910
rect 32645 17875 32655 17910
rect 32690 17875 32700 17910
rect 32735 17875 32745 17910
rect 32780 17875 32790 17910
rect 32825 17875 32835 17910
rect 32870 17875 32890 17910
rect 6740 17870 32890 17875
rect 2070 17865 32890 17870
rect 2070 17840 31305 17865
rect 2070 17800 2110 17840
rect 2150 17800 6700 17840
rect 6740 17830 31305 17840
rect 31340 17830 31350 17865
rect 31385 17830 31395 17865
rect 31430 17830 31440 17865
rect 31475 17830 31485 17865
rect 31520 17830 31530 17865
rect 31565 17830 31575 17865
rect 31610 17830 31620 17865
rect 31655 17830 31665 17865
rect 31700 17830 31710 17865
rect 31745 17830 31755 17865
rect 31790 17830 31800 17865
rect 31835 17830 31845 17865
rect 31880 17830 31890 17865
rect 31925 17830 31935 17865
rect 31970 17830 31980 17865
rect 32015 17830 32025 17865
rect 32060 17830 32070 17865
rect 32105 17830 32115 17865
rect 32150 17830 32160 17865
rect 32195 17830 32205 17865
rect 32240 17830 32250 17865
rect 32285 17830 32295 17865
rect 32330 17830 32340 17865
rect 32375 17830 32385 17865
rect 32420 17830 32430 17865
rect 32465 17830 32475 17865
rect 32510 17830 32520 17865
rect 32555 17830 32565 17865
rect 32600 17830 32610 17865
rect 32645 17830 32655 17865
rect 32690 17830 32700 17865
rect 32735 17830 32745 17865
rect 32780 17830 32790 17865
rect 32825 17830 32835 17865
rect 32870 17830 32890 17865
rect 6740 17820 32890 17830
rect 6740 17800 31305 17820
rect 2070 17785 31305 17800
rect 31340 17785 31350 17820
rect 31385 17785 31395 17820
rect 31430 17785 31440 17820
rect 31475 17785 31485 17820
rect 31520 17785 31530 17820
rect 31565 17785 31575 17820
rect 31610 17785 31620 17820
rect 31655 17785 31665 17820
rect 31700 17785 31710 17820
rect 31745 17785 31755 17820
rect 31790 17785 31800 17820
rect 31835 17785 31845 17820
rect 31880 17785 31890 17820
rect 31925 17785 31935 17820
rect 31970 17785 31980 17820
rect 32015 17785 32025 17820
rect 32060 17785 32070 17820
rect 32105 17785 32115 17820
rect 32150 17785 32160 17820
rect 32195 17785 32205 17820
rect 32240 17785 32250 17820
rect 32285 17785 32295 17820
rect 32330 17785 32340 17820
rect 32375 17785 32385 17820
rect 32420 17785 32430 17820
rect 32465 17785 32475 17820
rect 32510 17785 32520 17820
rect 32555 17785 32565 17820
rect 32600 17785 32610 17820
rect 32645 17785 32655 17820
rect 32690 17785 32700 17820
rect 32735 17785 32745 17820
rect 32780 17785 32790 17820
rect 32825 17785 32835 17820
rect 32870 17785 32890 17820
rect 2070 17775 32890 17785
rect 2070 17735 2110 17775
rect 2150 17735 6700 17775
rect 6740 17740 31305 17775
rect 31340 17740 31350 17775
rect 31385 17740 31395 17775
rect 31430 17740 31440 17775
rect 31475 17740 31485 17775
rect 31520 17740 31530 17775
rect 31565 17740 31575 17775
rect 31610 17740 31620 17775
rect 31655 17740 31665 17775
rect 31700 17740 31710 17775
rect 31745 17740 31755 17775
rect 31790 17740 31800 17775
rect 31835 17740 31845 17775
rect 31880 17740 31890 17775
rect 31925 17740 31935 17775
rect 31970 17740 31980 17775
rect 32015 17740 32025 17775
rect 32060 17740 32070 17775
rect 32105 17740 32115 17775
rect 32150 17740 32160 17775
rect 32195 17740 32205 17775
rect 32240 17740 32250 17775
rect 32285 17740 32295 17775
rect 32330 17740 32340 17775
rect 32375 17740 32385 17775
rect 32420 17740 32430 17775
rect 32465 17740 32475 17775
rect 32510 17740 32520 17775
rect 32555 17740 32565 17775
rect 32600 17740 32610 17775
rect 32645 17740 32655 17775
rect 32690 17740 32700 17775
rect 32735 17740 32745 17775
rect 32780 17740 32790 17775
rect 32825 17740 32835 17775
rect 32870 17740 32890 17775
rect 6740 17735 32890 17740
rect 2070 17725 32890 17735
rect -38770 9640 7700 9650
rect -38770 9630 1320 9640
rect -38770 9595 -38755 9630
rect -38720 9595 -38710 9630
rect -38675 9595 -38665 9630
rect -38630 9595 -38620 9630
rect -38585 9595 -38575 9630
rect -38540 9595 -38530 9630
rect -38495 9595 -38485 9630
rect -38450 9595 -38440 9630
rect -38405 9595 -38395 9630
rect -38360 9595 -38350 9630
rect -38315 9595 -38305 9630
rect -38270 9595 -38260 9630
rect -38225 9595 -38215 9630
rect -38180 9595 -38170 9630
rect -38135 9595 -38125 9630
rect -38090 9595 -38080 9630
rect -38045 9595 -38035 9630
rect -38000 9595 -37990 9630
rect -37955 9595 -37945 9630
rect -37910 9595 -37900 9630
rect -37865 9595 -37855 9630
rect -37820 9595 -37810 9630
rect -37775 9595 -37765 9630
rect -37730 9595 -37720 9630
rect -37685 9595 -37675 9630
rect -37640 9595 -37630 9630
rect -37595 9595 -37585 9630
rect -37550 9595 -37540 9630
rect -37505 9595 -37495 9630
rect -37460 9595 -37450 9630
rect -37415 9595 -37405 9630
rect -37370 9595 -37360 9630
rect -37325 9595 -37315 9630
rect -37280 9595 -37270 9630
rect -37235 9595 -37225 9630
rect -37190 9600 1320 9630
rect 1360 9600 2245 9640
rect 2285 9600 6700 9640
rect 6740 9600 7620 9640
rect 7660 9600 7700 9640
rect -37190 9595 7700 9600
rect -38770 9585 7700 9595
rect -38770 9550 -38755 9585
rect -38720 9550 -38710 9585
rect -38675 9550 -38665 9585
rect -38630 9550 -38620 9585
rect -38585 9550 -38575 9585
rect -38540 9550 -38530 9585
rect -38495 9550 -38485 9585
rect -38450 9550 -38440 9585
rect -38405 9550 -38395 9585
rect -38360 9550 -38350 9585
rect -38315 9550 -38305 9585
rect -38270 9550 -38260 9585
rect -38225 9550 -38215 9585
rect -38180 9550 -38170 9585
rect -38135 9550 -38125 9585
rect -38090 9550 -38080 9585
rect -38045 9550 -38035 9585
rect -38000 9550 -37990 9585
rect -37955 9550 -37945 9585
rect -37910 9550 -37900 9585
rect -37865 9550 -37855 9585
rect -37820 9550 -37810 9585
rect -37775 9550 -37765 9585
rect -37730 9550 -37720 9585
rect -37685 9550 -37675 9585
rect -37640 9550 -37630 9585
rect -37595 9550 -37585 9585
rect -37550 9550 -37540 9585
rect -37505 9550 -37495 9585
rect -37460 9550 -37450 9585
rect -37415 9550 -37405 9585
rect -37370 9550 -37360 9585
rect -37325 9550 -37315 9585
rect -37280 9550 -37270 9585
rect -37235 9550 -37225 9585
rect -37190 9575 7700 9585
rect -37190 9550 1320 9575
rect -38770 9540 1320 9550
rect -38770 9505 -38755 9540
rect -38720 9505 -38710 9540
rect -38675 9505 -38665 9540
rect -38630 9505 -38620 9540
rect -38585 9505 -38575 9540
rect -38540 9505 -38530 9540
rect -38495 9505 -38485 9540
rect -38450 9505 -38440 9540
rect -38405 9505 -38395 9540
rect -38360 9505 -38350 9540
rect -38315 9505 -38305 9540
rect -38270 9505 -38260 9540
rect -38225 9505 -38215 9540
rect -38180 9505 -38170 9540
rect -38135 9505 -38125 9540
rect -38090 9505 -38080 9540
rect -38045 9505 -38035 9540
rect -38000 9505 -37990 9540
rect -37955 9505 -37945 9540
rect -37910 9505 -37900 9540
rect -37865 9505 -37855 9540
rect -37820 9505 -37810 9540
rect -37775 9505 -37765 9540
rect -37730 9505 -37720 9540
rect -37685 9505 -37675 9540
rect -37640 9505 -37630 9540
rect -37595 9505 -37585 9540
rect -37550 9505 -37540 9540
rect -37505 9505 -37495 9540
rect -37460 9505 -37450 9540
rect -37415 9505 -37405 9540
rect -37370 9505 -37360 9540
rect -37325 9505 -37315 9540
rect -37280 9505 -37270 9540
rect -37235 9505 -37225 9540
rect -37190 9535 1320 9540
rect 1360 9535 2245 9575
rect 2285 9535 6700 9575
rect 6740 9535 7620 9575
rect 7660 9535 7700 9575
rect -37190 9505 7700 9535
rect -38770 9495 1320 9505
rect -38770 9460 -38755 9495
rect -38720 9460 -38710 9495
rect -38675 9460 -38665 9495
rect -38630 9460 -38620 9495
rect -38585 9460 -38575 9495
rect -38540 9460 -38530 9495
rect -38495 9460 -38485 9495
rect -38450 9460 -38440 9495
rect -38405 9460 -38395 9495
rect -38360 9460 -38350 9495
rect -38315 9460 -38305 9495
rect -38270 9460 -38260 9495
rect -38225 9460 -38215 9495
rect -38180 9460 -38170 9495
rect -38135 9460 -38125 9495
rect -38090 9460 -38080 9495
rect -38045 9460 -38035 9495
rect -38000 9460 -37990 9495
rect -37955 9460 -37945 9495
rect -37910 9460 -37900 9495
rect -37865 9460 -37855 9495
rect -37820 9460 -37810 9495
rect -37775 9460 -37765 9495
rect -37730 9460 -37720 9495
rect -37685 9460 -37675 9495
rect -37640 9460 -37630 9495
rect -37595 9460 -37585 9495
rect -37550 9460 -37540 9495
rect -37505 9460 -37495 9495
rect -37460 9460 -37450 9495
rect -37415 9460 -37405 9495
rect -37370 9460 -37360 9495
rect -37325 9460 -37315 9495
rect -37280 9460 -37270 9495
rect -37235 9460 -37225 9495
rect -37190 9465 1320 9495
rect 1360 9465 2245 9505
rect 2285 9465 6700 9505
rect 6740 9465 7620 9505
rect 7660 9465 7700 9505
rect -37190 9460 7700 9465
rect -38770 9450 7700 9460
rect -38770 9415 -38755 9450
rect -38720 9415 -38710 9450
rect -38675 9415 -38665 9450
rect -38630 9415 -38620 9450
rect -38585 9415 -38575 9450
rect -38540 9415 -38530 9450
rect -38495 9415 -38485 9450
rect -38450 9415 -38440 9450
rect -38405 9415 -38395 9450
rect -38360 9415 -38350 9450
rect -38315 9415 -38305 9450
rect -38270 9415 -38260 9450
rect -38225 9415 -38215 9450
rect -38180 9415 -38170 9450
rect -38135 9415 -38125 9450
rect -38090 9415 -38080 9450
rect -38045 9415 -38035 9450
rect -38000 9415 -37990 9450
rect -37955 9415 -37945 9450
rect -37910 9415 -37900 9450
rect -37865 9415 -37855 9450
rect -37820 9415 -37810 9450
rect -37775 9415 -37765 9450
rect -37730 9415 -37720 9450
rect -37685 9415 -37675 9450
rect -37640 9415 -37630 9450
rect -37595 9415 -37585 9450
rect -37550 9415 -37540 9450
rect -37505 9415 -37495 9450
rect -37460 9415 -37450 9450
rect -37415 9415 -37405 9450
rect -37370 9415 -37360 9450
rect -37325 9415 -37315 9450
rect -37280 9415 -37270 9450
rect -37235 9415 -37225 9450
rect -37190 9435 7700 9450
rect -37190 9415 1320 9435
rect -38770 9405 1320 9415
rect -38770 9370 -38755 9405
rect -38720 9370 -38710 9405
rect -38675 9370 -38665 9405
rect -38630 9370 -38620 9405
rect -38585 9370 -38575 9405
rect -38540 9370 -38530 9405
rect -38495 9370 -38485 9405
rect -38450 9370 -38440 9405
rect -38405 9370 -38395 9405
rect -38360 9370 -38350 9405
rect -38315 9370 -38305 9405
rect -38270 9370 -38260 9405
rect -38225 9370 -38215 9405
rect -38180 9370 -38170 9405
rect -38135 9370 -38125 9405
rect -38090 9370 -38080 9405
rect -38045 9370 -38035 9405
rect -38000 9370 -37990 9405
rect -37955 9370 -37945 9405
rect -37910 9370 -37900 9405
rect -37865 9370 -37855 9405
rect -37820 9370 -37810 9405
rect -37775 9370 -37765 9405
rect -37730 9370 -37720 9405
rect -37685 9370 -37675 9405
rect -37640 9370 -37630 9405
rect -37595 9370 -37585 9405
rect -37550 9370 -37540 9405
rect -37505 9370 -37495 9405
rect -37460 9370 -37450 9405
rect -37415 9370 -37405 9405
rect -37370 9370 -37360 9405
rect -37325 9370 -37315 9405
rect -37280 9370 -37270 9405
rect -37235 9370 -37225 9405
rect -37190 9395 1320 9405
rect 1360 9395 2245 9435
rect 2285 9395 6700 9435
rect 6740 9395 7620 9435
rect 7660 9395 7700 9435
rect -37190 9370 7700 9395
rect -38770 9365 7700 9370
rect -38770 9360 1320 9365
rect -38770 9325 -38755 9360
rect -38720 9325 -38710 9360
rect -38675 9325 -38665 9360
rect -38630 9325 -38620 9360
rect -38585 9325 -38575 9360
rect -38540 9325 -38530 9360
rect -38495 9325 -38485 9360
rect -38450 9325 -38440 9360
rect -38405 9325 -38395 9360
rect -38360 9325 -38350 9360
rect -38315 9325 -38305 9360
rect -38270 9325 -38260 9360
rect -38225 9325 -38215 9360
rect -38180 9325 -38170 9360
rect -38135 9325 -38125 9360
rect -38090 9325 -38080 9360
rect -38045 9325 -38035 9360
rect -38000 9325 -37990 9360
rect -37955 9325 -37945 9360
rect -37910 9325 -37900 9360
rect -37865 9325 -37855 9360
rect -37820 9325 -37810 9360
rect -37775 9325 -37765 9360
rect -37730 9325 -37720 9360
rect -37685 9325 -37675 9360
rect -37640 9325 -37630 9360
rect -37595 9325 -37585 9360
rect -37550 9325 -37540 9360
rect -37505 9325 -37495 9360
rect -37460 9325 -37450 9360
rect -37415 9325 -37405 9360
rect -37370 9325 -37360 9360
rect -37325 9325 -37315 9360
rect -37280 9325 -37270 9360
rect -37235 9325 -37225 9360
rect -37190 9325 1320 9360
rect 1360 9325 2245 9365
rect 2285 9325 6700 9365
rect 6740 9325 7620 9365
rect 7660 9325 7700 9365
rect -38770 9315 7700 9325
rect -38770 9280 -38755 9315
rect -38720 9280 -38710 9315
rect -38675 9280 -38665 9315
rect -38630 9280 -38620 9315
rect -38585 9280 -38575 9315
rect -38540 9280 -38530 9315
rect -38495 9280 -38485 9315
rect -38450 9280 -38440 9315
rect -38405 9280 -38395 9315
rect -38360 9280 -38350 9315
rect -38315 9280 -38305 9315
rect -38270 9280 -38260 9315
rect -38225 9280 -38215 9315
rect -38180 9280 -38170 9315
rect -38135 9280 -38125 9315
rect -38090 9280 -38080 9315
rect -38045 9280 -38035 9315
rect -38000 9280 -37990 9315
rect -37955 9280 -37945 9315
rect -37910 9280 -37900 9315
rect -37865 9280 -37855 9315
rect -37820 9280 -37810 9315
rect -37775 9280 -37765 9315
rect -37730 9280 -37720 9315
rect -37685 9280 -37675 9315
rect -37640 9280 -37630 9315
rect -37595 9280 -37585 9315
rect -37550 9280 -37540 9315
rect -37505 9280 -37495 9315
rect -37460 9280 -37450 9315
rect -37415 9280 -37405 9315
rect -37370 9280 -37360 9315
rect -37325 9280 -37315 9315
rect -37280 9280 -37270 9315
rect -37235 9280 -37225 9315
rect -37190 9300 7700 9315
rect -37190 9280 1320 9300
rect -38770 9270 1320 9280
rect -38770 9235 -38755 9270
rect -38720 9235 -38710 9270
rect -38675 9235 -38665 9270
rect -38630 9235 -38620 9270
rect -38585 9235 -38575 9270
rect -38540 9235 -38530 9270
rect -38495 9235 -38485 9270
rect -38450 9235 -38440 9270
rect -38405 9235 -38395 9270
rect -38360 9235 -38350 9270
rect -38315 9235 -38305 9270
rect -38270 9235 -38260 9270
rect -38225 9235 -38215 9270
rect -38180 9235 -38170 9270
rect -38135 9235 -38125 9270
rect -38090 9235 -38080 9270
rect -38045 9235 -38035 9270
rect -38000 9235 -37990 9270
rect -37955 9235 -37945 9270
rect -37910 9235 -37900 9270
rect -37865 9235 -37855 9270
rect -37820 9235 -37810 9270
rect -37775 9235 -37765 9270
rect -37730 9235 -37720 9270
rect -37685 9235 -37675 9270
rect -37640 9235 -37630 9270
rect -37595 9235 -37585 9270
rect -37550 9235 -37540 9270
rect -37505 9235 -37495 9270
rect -37460 9235 -37450 9270
rect -37415 9235 -37405 9270
rect -37370 9235 -37360 9270
rect -37325 9235 -37315 9270
rect -37280 9235 -37270 9270
rect -37235 9235 -37225 9270
rect -37190 9260 1320 9270
rect 1360 9260 2245 9300
rect 2285 9260 6700 9300
rect 6740 9260 7620 9300
rect 7660 9260 7700 9300
rect -37190 9240 7700 9260
rect -37190 9235 1320 9240
rect -38770 9225 1320 9235
rect -38770 9190 -38755 9225
rect -38720 9190 -38710 9225
rect -38675 9190 -38665 9225
rect -38630 9190 -38620 9225
rect -38585 9190 -38575 9225
rect -38540 9190 -38530 9225
rect -38495 9190 -38485 9225
rect -38450 9190 -38440 9225
rect -38405 9190 -38395 9225
rect -38360 9190 -38350 9225
rect -38315 9190 -38305 9225
rect -38270 9190 -38260 9225
rect -38225 9190 -38215 9225
rect -38180 9190 -38170 9225
rect -38135 9190 -38125 9225
rect -38090 9190 -38080 9225
rect -38045 9190 -38035 9225
rect -38000 9190 -37990 9225
rect -37955 9190 -37945 9225
rect -37910 9190 -37900 9225
rect -37865 9190 -37855 9225
rect -37820 9190 -37810 9225
rect -37775 9190 -37765 9225
rect -37730 9190 -37720 9225
rect -37685 9190 -37675 9225
rect -37640 9190 -37630 9225
rect -37595 9190 -37585 9225
rect -37550 9190 -37540 9225
rect -37505 9190 -37495 9225
rect -37460 9190 -37450 9225
rect -37415 9190 -37405 9225
rect -37370 9190 -37360 9225
rect -37325 9190 -37315 9225
rect -37280 9190 -37270 9225
rect -37235 9190 -37225 9225
rect -37190 9200 1320 9225
rect 1360 9200 2245 9240
rect 2285 9200 6700 9240
rect 6740 9200 7620 9240
rect 7660 9200 7700 9240
rect -37190 9190 7700 9200
rect -38770 9180 7700 9190
rect -38770 9145 -38755 9180
rect -38720 9145 -38710 9180
rect -38675 9145 -38665 9180
rect -38630 9145 -38620 9180
rect -38585 9145 -38575 9180
rect -38540 9145 -38530 9180
rect -38495 9145 -38485 9180
rect -38450 9145 -38440 9180
rect -38405 9145 -38395 9180
rect -38360 9145 -38350 9180
rect -38315 9145 -38305 9180
rect -38270 9145 -38260 9180
rect -38225 9145 -38215 9180
rect -38180 9145 -38170 9180
rect -38135 9145 -38125 9180
rect -38090 9145 -38080 9180
rect -38045 9145 -38035 9180
rect -38000 9145 -37990 9180
rect -37955 9145 -37945 9180
rect -37910 9145 -37900 9180
rect -37865 9145 -37855 9180
rect -37820 9145 -37810 9180
rect -37775 9145 -37765 9180
rect -37730 9145 -37720 9180
rect -37685 9145 -37675 9180
rect -37640 9145 -37630 9180
rect -37595 9145 -37585 9180
rect -37550 9145 -37540 9180
rect -37505 9145 -37495 9180
rect -37460 9145 -37450 9180
rect -37415 9145 -37405 9180
rect -37370 9145 -37360 9180
rect -37325 9145 -37315 9180
rect -37280 9145 -37270 9180
rect -37235 9145 -37225 9180
rect -37190 9175 7700 9180
rect -37190 9145 1320 9175
rect -38770 9135 1320 9145
rect 1360 9135 2245 9175
rect 2285 9135 6700 9175
rect 6740 9135 7620 9175
rect 7660 9135 7700 9175
rect -38770 9100 -38755 9135
rect -38720 9100 -38710 9135
rect -38675 9100 -38665 9135
rect -38630 9100 -38620 9135
rect -38585 9100 -38575 9135
rect -38540 9100 -38530 9135
rect -38495 9100 -38485 9135
rect -38450 9100 -38440 9135
rect -38405 9100 -38395 9135
rect -38360 9100 -38350 9135
rect -38315 9100 -38305 9135
rect -38270 9100 -38260 9135
rect -38225 9100 -38215 9135
rect -38180 9100 -38170 9135
rect -38135 9100 -38125 9135
rect -38090 9100 -38080 9135
rect -38045 9100 -38035 9135
rect -38000 9100 -37990 9135
rect -37955 9100 -37945 9135
rect -37910 9100 -37900 9135
rect -37865 9100 -37855 9135
rect -37820 9100 -37810 9135
rect -37775 9100 -37765 9135
rect -37730 9100 -37720 9135
rect -37685 9100 -37675 9135
rect -37640 9100 -37630 9135
rect -37595 9100 -37585 9135
rect -37550 9100 -37540 9135
rect -37505 9100 -37495 9135
rect -37460 9100 -37450 9135
rect -37415 9100 -37405 9135
rect -37370 9100 -37360 9135
rect -37325 9100 -37315 9135
rect -37280 9100 -37270 9135
rect -37235 9100 -37225 9135
rect -37190 9105 7700 9135
rect -37190 9100 1320 9105
rect -38770 9090 1320 9100
rect -38770 9055 -38755 9090
rect -38720 9055 -38710 9090
rect -38675 9055 -38665 9090
rect -38630 9055 -38620 9090
rect -38585 9055 -38575 9090
rect -38540 9055 -38530 9090
rect -38495 9055 -38485 9090
rect -38450 9055 -38440 9090
rect -38405 9055 -38395 9090
rect -38360 9055 -38350 9090
rect -38315 9055 -38305 9090
rect -38270 9055 -38260 9090
rect -38225 9055 -38215 9090
rect -38180 9055 -38170 9090
rect -38135 9055 -38125 9090
rect -38090 9055 -38080 9090
rect -38045 9055 -38035 9090
rect -38000 9055 -37990 9090
rect -37955 9055 -37945 9090
rect -37910 9055 -37900 9090
rect -37865 9055 -37855 9090
rect -37820 9055 -37810 9090
rect -37775 9055 -37765 9090
rect -37730 9055 -37720 9090
rect -37685 9055 -37675 9090
rect -37640 9055 -37630 9090
rect -37595 9055 -37585 9090
rect -37550 9055 -37540 9090
rect -37505 9055 -37495 9090
rect -37460 9055 -37450 9090
rect -37415 9055 -37405 9090
rect -37370 9055 -37360 9090
rect -37325 9055 -37315 9090
rect -37280 9055 -37270 9090
rect -37235 9055 -37225 9090
rect -37190 9065 1320 9090
rect 1360 9065 2245 9105
rect 2285 9065 6700 9105
rect 6740 9065 7620 9105
rect 7660 9065 7700 9105
rect -37190 9055 7700 9065
rect -38770 9045 7700 9055
rect -38770 9010 -38755 9045
rect -38720 9010 -38710 9045
rect -38675 9010 -38665 9045
rect -38630 9010 -38620 9045
rect -38585 9010 -38575 9045
rect -38540 9010 -38530 9045
rect -38495 9010 -38485 9045
rect -38450 9010 -38440 9045
rect -38405 9010 -38395 9045
rect -38360 9010 -38350 9045
rect -38315 9010 -38305 9045
rect -38270 9010 -38260 9045
rect -38225 9010 -38215 9045
rect -38180 9010 -38170 9045
rect -38135 9010 -38125 9045
rect -38090 9010 -38080 9045
rect -38045 9010 -38035 9045
rect -38000 9010 -37990 9045
rect -37955 9010 -37945 9045
rect -37910 9010 -37900 9045
rect -37865 9010 -37855 9045
rect -37820 9010 -37810 9045
rect -37775 9010 -37765 9045
rect -37730 9010 -37720 9045
rect -37685 9010 -37675 9045
rect -37640 9010 -37630 9045
rect -37595 9010 -37585 9045
rect -37550 9010 -37540 9045
rect -37505 9010 -37495 9045
rect -37460 9010 -37450 9045
rect -37415 9010 -37405 9045
rect -37370 9010 -37360 9045
rect -37325 9010 -37315 9045
rect -37280 9010 -37270 9045
rect -37235 9010 -37225 9045
rect -37190 9035 7700 9045
rect -37190 9010 1320 9035
rect -38770 9000 1320 9010
rect -38770 8965 -38755 9000
rect -38720 8965 -38710 9000
rect -38675 8965 -38665 9000
rect -38630 8965 -38620 9000
rect -38585 8965 -38575 9000
rect -38540 8965 -38530 9000
rect -38495 8965 -38485 9000
rect -38450 8965 -38440 9000
rect -38405 8965 -38395 9000
rect -38360 8965 -38350 9000
rect -38315 8965 -38305 9000
rect -38270 8965 -38260 9000
rect -38225 8965 -38215 9000
rect -38180 8965 -38170 9000
rect -38135 8965 -38125 9000
rect -38090 8965 -38080 9000
rect -38045 8965 -38035 9000
rect -38000 8965 -37990 9000
rect -37955 8965 -37945 9000
rect -37910 8965 -37900 9000
rect -37865 8965 -37855 9000
rect -37820 8965 -37810 9000
rect -37775 8965 -37765 9000
rect -37730 8965 -37720 9000
rect -37685 8965 -37675 9000
rect -37640 8965 -37630 9000
rect -37595 8965 -37585 9000
rect -37550 8965 -37540 9000
rect -37505 8965 -37495 9000
rect -37460 8965 -37450 9000
rect -37415 8965 -37405 9000
rect -37370 8965 -37360 9000
rect -37325 8965 -37315 9000
rect -37280 8965 -37270 9000
rect -37235 8965 -37225 9000
rect -37190 8995 1320 9000
rect 1360 8995 2245 9035
rect 2285 8995 6700 9035
rect 6740 8995 7620 9035
rect 7660 8995 7700 9035
rect -37190 8965 7700 8995
rect -38770 8955 1320 8965
rect -38770 8920 -38755 8955
rect -38720 8920 -38710 8955
rect -38675 8920 -38665 8955
rect -38630 8920 -38620 8955
rect -38585 8920 -38575 8955
rect -38540 8920 -38530 8955
rect -38495 8920 -38485 8955
rect -38450 8920 -38440 8955
rect -38405 8920 -38395 8955
rect -38360 8920 -38350 8955
rect -38315 8920 -38305 8955
rect -38270 8920 -38260 8955
rect -38225 8920 -38215 8955
rect -38180 8920 -38170 8955
rect -38135 8920 -38125 8955
rect -38090 8920 -38080 8955
rect -38045 8920 -38035 8955
rect -38000 8920 -37990 8955
rect -37955 8920 -37945 8955
rect -37910 8920 -37900 8955
rect -37865 8920 -37855 8955
rect -37820 8920 -37810 8955
rect -37775 8920 -37765 8955
rect -37730 8920 -37720 8955
rect -37685 8920 -37675 8955
rect -37640 8920 -37630 8955
rect -37595 8920 -37585 8955
rect -37550 8920 -37540 8955
rect -37505 8920 -37495 8955
rect -37460 8920 -37450 8955
rect -37415 8920 -37405 8955
rect -37370 8920 -37360 8955
rect -37325 8920 -37315 8955
rect -37280 8920 -37270 8955
rect -37235 8920 -37225 8955
rect -37190 8925 1320 8955
rect 1360 8925 2245 8965
rect 2285 8925 6700 8965
rect 6740 8925 7620 8965
rect 7660 8925 7700 8965
rect -37190 8920 7700 8925
rect -38770 8910 7700 8920
rect -38770 8875 -38755 8910
rect -38720 8875 -38710 8910
rect -38675 8875 -38665 8910
rect -38630 8875 -38620 8910
rect -38585 8875 -38575 8910
rect -38540 8875 -38530 8910
rect -38495 8875 -38485 8910
rect -38450 8875 -38440 8910
rect -38405 8875 -38395 8910
rect -38360 8875 -38350 8910
rect -38315 8875 -38305 8910
rect -38270 8875 -38260 8910
rect -38225 8875 -38215 8910
rect -38180 8875 -38170 8910
rect -38135 8875 -38125 8910
rect -38090 8875 -38080 8910
rect -38045 8875 -38035 8910
rect -38000 8875 -37990 8910
rect -37955 8875 -37945 8910
rect -37910 8875 -37900 8910
rect -37865 8875 -37855 8910
rect -37820 8875 -37810 8910
rect -37775 8875 -37765 8910
rect -37730 8875 -37720 8910
rect -37685 8875 -37675 8910
rect -37640 8875 -37630 8910
rect -37595 8875 -37585 8910
rect -37550 8875 -37540 8910
rect -37505 8875 -37495 8910
rect -37460 8875 -37450 8910
rect -37415 8875 -37405 8910
rect -37370 8875 -37360 8910
rect -37325 8875 -37315 8910
rect -37280 8875 -37270 8910
rect -37235 8875 -37225 8910
rect -37190 8900 7700 8910
rect -37190 8875 1320 8900
rect -38770 8865 1320 8875
rect -38770 8830 -38755 8865
rect -38720 8830 -38710 8865
rect -38675 8830 -38665 8865
rect -38630 8830 -38620 8865
rect -38585 8830 -38575 8865
rect -38540 8830 -38530 8865
rect -38495 8830 -38485 8865
rect -38450 8830 -38440 8865
rect -38405 8830 -38395 8865
rect -38360 8830 -38350 8865
rect -38315 8830 -38305 8865
rect -38270 8830 -38260 8865
rect -38225 8830 -38215 8865
rect -38180 8830 -38170 8865
rect -38135 8830 -38125 8865
rect -38090 8830 -38080 8865
rect -38045 8830 -38035 8865
rect -38000 8830 -37990 8865
rect -37955 8830 -37945 8865
rect -37910 8830 -37900 8865
rect -37865 8830 -37855 8865
rect -37820 8830 -37810 8865
rect -37775 8830 -37765 8865
rect -37730 8830 -37720 8865
rect -37685 8830 -37675 8865
rect -37640 8830 -37630 8865
rect -37595 8830 -37585 8865
rect -37550 8830 -37540 8865
rect -37505 8830 -37495 8865
rect -37460 8830 -37450 8865
rect -37415 8830 -37405 8865
rect -37370 8830 -37360 8865
rect -37325 8830 -37315 8865
rect -37280 8830 -37270 8865
rect -37235 8830 -37225 8865
rect -37190 8860 1320 8865
rect 1360 8860 2245 8900
rect 2285 8860 6700 8900
rect 6740 8860 7620 8900
rect 7660 8860 7700 8900
rect -37190 8840 7700 8860
rect -37190 8830 1320 8840
rect -38770 8820 1320 8830
rect -38770 8785 -38755 8820
rect -38720 8785 -38710 8820
rect -38675 8785 -38665 8820
rect -38630 8785 -38620 8820
rect -38585 8785 -38575 8820
rect -38540 8785 -38530 8820
rect -38495 8785 -38485 8820
rect -38450 8785 -38440 8820
rect -38405 8785 -38395 8820
rect -38360 8785 -38350 8820
rect -38315 8785 -38305 8820
rect -38270 8785 -38260 8820
rect -38225 8785 -38215 8820
rect -38180 8785 -38170 8820
rect -38135 8785 -38125 8820
rect -38090 8785 -38080 8820
rect -38045 8785 -38035 8820
rect -38000 8785 -37990 8820
rect -37955 8785 -37945 8820
rect -37910 8785 -37900 8820
rect -37865 8785 -37855 8820
rect -37820 8785 -37810 8820
rect -37775 8785 -37765 8820
rect -37730 8785 -37720 8820
rect -37685 8785 -37675 8820
rect -37640 8785 -37630 8820
rect -37595 8785 -37585 8820
rect -37550 8785 -37540 8820
rect -37505 8785 -37495 8820
rect -37460 8785 -37450 8820
rect -37415 8785 -37405 8820
rect -37370 8785 -37360 8820
rect -37325 8785 -37315 8820
rect -37280 8785 -37270 8820
rect -37235 8785 -37225 8820
rect -37190 8800 1320 8820
rect 1360 8800 2245 8840
rect 2285 8800 6700 8840
rect 6740 8800 7620 8840
rect 7660 8800 7700 8840
rect -37190 8785 7700 8800
rect -38770 8775 7700 8785
rect -38770 8740 -38755 8775
rect -38720 8740 -38710 8775
rect -38675 8740 -38665 8775
rect -38630 8740 -38620 8775
rect -38585 8740 -38575 8775
rect -38540 8740 -38530 8775
rect -38495 8740 -38485 8775
rect -38450 8740 -38440 8775
rect -38405 8740 -38395 8775
rect -38360 8740 -38350 8775
rect -38315 8740 -38305 8775
rect -38270 8740 -38260 8775
rect -38225 8740 -38215 8775
rect -38180 8740 -38170 8775
rect -38135 8740 -38125 8775
rect -38090 8740 -38080 8775
rect -38045 8740 -38035 8775
rect -38000 8740 -37990 8775
rect -37955 8740 -37945 8775
rect -37910 8740 -37900 8775
rect -37865 8740 -37855 8775
rect -37820 8740 -37810 8775
rect -37775 8740 -37765 8775
rect -37730 8740 -37720 8775
rect -37685 8740 -37675 8775
rect -37640 8740 -37630 8775
rect -37595 8740 -37585 8775
rect -37550 8740 -37540 8775
rect -37505 8740 -37495 8775
rect -37460 8740 -37450 8775
rect -37415 8740 -37405 8775
rect -37370 8740 -37360 8775
rect -37325 8740 -37315 8775
rect -37280 8740 -37270 8775
rect -37235 8740 -37225 8775
rect -37190 8740 1320 8775
rect -38770 8735 1320 8740
rect 1360 8735 2245 8775
rect 2285 8735 6700 8775
rect 6740 8735 7620 8775
rect 7660 8735 7700 8775
rect -38770 8730 7700 8735
rect -38770 8695 -38755 8730
rect -38720 8695 -38710 8730
rect -38675 8695 -38665 8730
rect -38630 8695 -38620 8730
rect -38585 8695 -38575 8730
rect -38540 8695 -38530 8730
rect -38495 8695 -38485 8730
rect -38450 8695 -38440 8730
rect -38405 8695 -38395 8730
rect -38360 8695 -38350 8730
rect -38315 8695 -38305 8730
rect -38270 8695 -38260 8730
rect -38225 8695 -38215 8730
rect -38180 8695 -38170 8730
rect -38135 8695 -38125 8730
rect -38090 8695 -38080 8730
rect -38045 8695 -38035 8730
rect -38000 8695 -37990 8730
rect -37955 8695 -37945 8730
rect -37910 8695 -37900 8730
rect -37865 8695 -37855 8730
rect -37820 8695 -37810 8730
rect -37775 8695 -37765 8730
rect -37730 8695 -37720 8730
rect -37685 8695 -37675 8730
rect -37640 8695 -37630 8730
rect -37595 8695 -37585 8730
rect -37550 8695 -37540 8730
rect -37505 8695 -37495 8730
rect -37460 8695 -37450 8730
rect -37415 8695 -37405 8730
rect -37370 8695 -37360 8730
rect -37325 8695 -37315 8730
rect -37280 8695 -37270 8730
rect -37235 8695 -37225 8730
rect -37190 8705 7700 8730
rect -37190 8695 1320 8705
rect -38770 8685 1320 8695
rect -38770 8650 -38755 8685
rect -38720 8650 -38710 8685
rect -38675 8650 -38665 8685
rect -38630 8650 -38620 8685
rect -38585 8650 -38575 8685
rect -38540 8650 -38530 8685
rect -38495 8650 -38485 8685
rect -38450 8650 -38440 8685
rect -38405 8650 -38395 8685
rect -38360 8650 -38350 8685
rect -38315 8650 -38305 8685
rect -38270 8650 -38260 8685
rect -38225 8650 -38215 8685
rect -38180 8650 -38170 8685
rect -38135 8650 -38125 8685
rect -38090 8650 -38080 8685
rect -38045 8650 -38035 8685
rect -38000 8650 -37990 8685
rect -37955 8650 -37945 8685
rect -37910 8650 -37900 8685
rect -37865 8650 -37855 8685
rect -37820 8650 -37810 8685
rect -37775 8650 -37765 8685
rect -37730 8650 -37720 8685
rect -37685 8650 -37675 8685
rect -37640 8650 -37630 8685
rect -37595 8650 -37585 8685
rect -37550 8650 -37540 8685
rect -37505 8650 -37495 8685
rect -37460 8650 -37450 8685
rect -37415 8650 -37405 8685
rect -37370 8650 -37360 8685
rect -37325 8650 -37315 8685
rect -37280 8650 -37270 8685
rect -37235 8650 -37225 8685
rect -37190 8665 1320 8685
rect 1360 8665 2245 8705
rect 2285 8665 6700 8705
rect 6740 8665 7620 8705
rect 7660 8665 7700 8705
rect -37190 8650 7700 8665
rect -38770 8640 7700 8650
rect -38770 8605 -38755 8640
rect -38720 8605 -38710 8640
rect -38675 8605 -38665 8640
rect -38630 8605 -38620 8640
rect -38585 8605 -38575 8640
rect -38540 8605 -38530 8640
rect -38495 8605 -38485 8640
rect -38450 8605 -38440 8640
rect -38405 8605 -38395 8640
rect -38360 8605 -38350 8640
rect -38315 8605 -38305 8640
rect -38270 8605 -38260 8640
rect -38225 8605 -38215 8640
rect -38180 8605 -38170 8640
rect -38135 8605 -38125 8640
rect -38090 8605 -38080 8640
rect -38045 8605 -38035 8640
rect -38000 8605 -37990 8640
rect -37955 8605 -37945 8640
rect -37910 8605 -37900 8640
rect -37865 8605 -37855 8640
rect -37820 8605 -37810 8640
rect -37775 8605 -37765 8640
rect -37730 8605 -37720 8640
rect -37685 8605 -37675 8640
rect -37640 8605 -37630 8640
rect -37595 8605 -37585 8640
rect -37550 8605 -37540 8640
rect -37505 8605 -37495 8640
rect -37460 8605 -37450 8640
rect -37415 8605 -37405 8640
rect -37370 8605 -37360 8640
rect -37325 8605 -37315 8640
rect -37280 8605 -37270 8640
rect -37235 8605 -37225 8640
rect -37190 8635 7700 8640
rect -37190 8605 1320 8635
rect -38770 8595 1320 8605
rect 1360 8595 2245 8635
rect 2285 8595 6700 8635
rect 6740 8595 7620 8635
rect 7660 8595 7700 8635
rect -38770 8560 -38755 8595
rect -38720 8560 -38710 8595
rect -38675 8560 -38665 8595
rect -38630 8560 -38620 8595
rect -38585 8560 -38575 8595
rect -38540 8560 -38530 8595
rect -38495 8560 -38485 8595
rect -38450 8560 -38440 8595
rect -38405 8560 -38395 8595
rect -38360 8560 -38350 8595
rect -38315 8560 -38305 8595
rect -38270 8560 -38260 8595
rect -38225 8560 -38215 8595
rect -38180 8560 -38170 8595
rect -38135 8560 -38125 8595
rect -38090 8560 -38080 8595
rect -38045 8560 -38035 8595
rect -38000 8560 -37990 8595
rect -37955 8560 -37945 8595
rect -37910 8560 -37900 8595
rect -37865 8560 -37855 8595
rect -37820 8560 -37810 8595
rect -37775 8560 -37765 8595
rect -37730 8560 -37720 8595
rect -37685 8560 -37675 8595
rect -37640 8560 -37630 8595
rect -37595 8560 -37585 8595
rect -37550 8560 -37540 8595
rect -37505 8560 -37495 8595
rect -37460 8560 -37450 8595
rect -37415 8560 -37405 8595
rect -37370 8560 -37360 8595
rect -37325 8560 -37315 8595
rect -37280 8560 -37270 8595
rect -37235 8560 -37225 8595
rect -37190 8565 7700 8595
rect -37190 8560 1320 8565
rect -38770 8550 1320 8560
rect -38770 8515 -38755 8550
rect -38720 8515 -38710 8550
rect -38675 8515 -38665 8550
rect -38630 8515 -38620 8550
rect -38585 8515 -38575 8550
rect -38540 8515 -38530 8550
rect -38495 8515 -38485 8550
rect -38450 8515 -38440 8550
rect -38405 8515 -38395 8550
rect -38360 8515 -38350 8550
rect -38315 8515 -38305 8550
rect -38270 8515 -38260 8550
rect -38225 8515 -38215 8550
rect -38180 8515 -38170 8550
rect -38135 8515 -38125 8550
rect -38090 8515 -38080 8550
rect -38045 8515 -38035 8550
rect -38000 8515 -37990 8550
rect -37955 8515 -37945 8550
rect -37910 8515 -37900 8550
rect -37865 8515 -37855 8550
rect -37820 8515 -37810 8550
rect -37775 8515 -37765 8550
rect -37730 8515 -37720 8550
rect -37685 8515 -37675 8550
rect -37640 8515 -37630 8550
rect -37595 8515 -37585 8550
rect -37550 8515 -37540 8550
rect -37505 8515 -37495 8550
rect -37460 8515 -37450 8550
rect -37415 8515 -37405 8550
rect -37370 8515 -37360 8550
rect -37325 8515 -37315 8550
rect -37280 8515 -37270 8550
rect -37235 8515 -37225 8550
rect -37190 8525 1320 8550
rect 1360 8525 2245 8565
rect 2285 8525 6700 8565
rect 6740 8525 7620 8565
rect 7660 8525 7700 8565
rect -37190 8515 7700 8525
rect -38770 8505 7700 8515
rect -38770 8470 -38755 8505
rect -38720 8470 -38710 8505
rect -38675 8470 -38665 8505
rect -38630 8470 -38620 8505
rect -38585 8470 -38575 8505
rect -38540 8470 -38530 8505
rect -38495 8470 -38485 8505
rect -38450 8470 -38440 8505
rect -38405 8470 -38395 8505
rect -38360 8470 -38350 8505
rect -38315 8470 -38305 8505
rect -38270 8470 -38260 8505
rect -38225 8470 -38215 8505
rect -38180 8470 -38170 8505
rect -38135 8470 -38125 8505
rect -38090 8470 -38080 8505
rect -38045 8470 -38035 8505
rect -38000 8470 -37990 8505
rect -37955 8470 -37945 8505
rect -37910 8470 -37900 8505
rect -37865 8470 -37855 8505
rect -37820 8470 -37810 8505
rect -37775 8470 -37765 8505
rect -37730 8470 -37720 8505
rect -37685 8470 -37675 8505
rect -37640 8470 -37630 8505
rect -37595 8470 -37585 8505
rect -37550 8470 -37540 8505
rect -37505 8470 -37495 8505
rect -37460 8470 -37450 8505
rect -37415 8470 -37405 8505
rect -37370 8470 -37360 8505
rect -37325 8470 -37315 8505
rect -37280 8470 -37270 8505
rect -37235 8470 -37225 8505
rect -37190 8500 7700 8505
rect -37190 8470 1320 8500
rect -38770 8460 1320 8470
rect 1360 8460 2245 8500
rect 2285 8460 6700 8500
rect 6740 8460 7620 8500
rect 7660 8460 7700 8500
rect -38770 8425 -38755 8460
rect -38720 8425 -38710 8460
rect -38675 8425 -38665 8460
rect -38630 8425 -38620 8460
rect -38585 8425 -38575 8460
rect -38540 8425 -38530 8460
rect -38495 8425 -38485 8460
rect -38450 8425 -38440 8460
rect -38405 8425 -38395 8460
rect -38360 8425 -38350 8460
rect -38315 8425 -38305 8460
rect -38270 8425 -38260 8460
rect -38225 8425 -38215 8460
rect -38180 8425 -38170 8460
rect -38135 8425 -38125 8460
rect -38090 8425 -38080 8460
rect -38045 8425 -38035 8460
rect -38000 8425 -37990 8460
rect -37955 8425 -37945 8460
rect -37910 8425 -37900 8460
rect -37865 8425 -37855 8460
rect -37820 8425 -37810 8460
rect -37775 8425 -37765 8460
rect -37730 8425 -37720 8460
rect -37685 8425 -37675 8460
rect -37640 8425 -37630 8460
rect -37595 8425 -37585 8460
rect -37550 8425 -37540 8460
rect -37505 8425 -37495 8460
rect -37460 8425 -37450 8460
rect -37415 8425 -37405 8460
rect -37370 8425 -37360 8460
rect -37325 8425 -37315 8460
rect -37280 8425 -37270 8460
rect -37235 8425 -37225 8460
rect -37190 8440 7700 8460
rect -37190 8425 1320 8440
rect -38770 8415 1320 8425
rect -38770 8380 -38755 8415
rect -38720 8380 -38710 8415
rect -38675 8380 -38665 8415
rect -38630 8380 -38620 8415
rect -38585 8380 -38575 8415
rect -38540 8380 -38530 8415
rect -38495 8380 -38485 8415
rect -38450 8380 -38440 8415
rect -38405 8380 -38395 8415
rect -38360 8380 -38350 8415
rect -38315 8380 -38305 8415
rect -38270 8380 -38260 8415
rect -38225 8380 -38215 8415
rect -38180 8380 -38170 8415
rect -38135 8380 -38125 8415
rect -38090 8380 -38080 8415
rect -38045 8380 -38035 8415
rect -38000 8380 -37990 8415
rect -37955 8380 -37945 8415
rect -37910 8380 -37900 8415
rect -37865 8380 -37855 8415
rect -37820 8380 -37810 8415
rect -37775 8380 -37765 8415
rect -37730 8380 -37720 8415
rect -37685 8380 -37675 8415
rect -37640 8380 -37630 8415
rect -37595 8380 -37585 8415
rect -37550 8380 -37540 8415
rect -37505 8380 -37495 8415
rect -37460 8380 -37450 8415
rect -37415 8380 -37405 8415
rect -37370 8380 -37360 8415
rect -37325 8380 -37315 8415
rect -37280 8380 -37270 8415
rect -37235 8380 -37225 8415
rect -37190 8400 1320 8415
rect 1360 8400 2245 8440
rect 2285 8400 6700 8440
rect 6740 8400 7620 8440
rect 7660 8400 7700 8440
rect -37190 8380 7700 8400
rect -38770 8375 7700 8380
rect -38770 8370 1320 8375
rect -38770 8335 -38755 8370
rect -38720 8335 -38710 8370
rect -38675 8335 -38665 8370
rect -38630 8335 -38620 8370
rect -38585 8335 -38575 8370
rect -38540 8335 -38530 8370
rect -38495 8335 -38485 8370
rect -38450 8335 -38440 8370
rect -38405 8335 -38395 8370
rect -38360 8335 -38350 8370
rect -38315 8335 -38305 8370
rect -38270 8335 -38260 8370
rect -38225 8335 -38215 8370
rect -38180 8335 -38170 8370
rect -38135 8335 -38125 8370
rect -38090 8335 -38080 8370
rect -38045 8335 -38035 8370
rect -38000 8335 -37990 8370
rect -37955 8335 -37945 8370
rect -37910 8335 -37900 8370
rect -37865 8335 -37855 8370
rect -37820 8335 -37810 8370
rect -37775 8335 -37765 8370
rect -37730 8335 -37720 8370
rect -37685 8335 -37675 8370
rect -37640 8335 -37630 8370
rect -37595 8335 -37585 8370
rect -37550 8335 -37540 8370
rect -37505 8335 -37495 8370
rect -37460 8335 -37450 8370
rect -37415 8335 -37405 8370
rect -37370 8335 -37360 8370
rect -37325 8335 -37315 8370
rect -37280 8335 -37270 8370
rect -37235 8335 -37225 8370
rect -37190 8335 1320 8370
rect 1360 8335 2245 8375
rect 2285 8335 6700 8375
rect 6740 8335 7620 8375
rect 7660 8335 7700 8375
rect -38770 8325 7700 8335
rect -38770 8290 -38755 8325
rect -38720 8290 -38710 8325
rect -38675 8290 -38665 8325
rect -38630 8290 -38620 8325
rect -38585 8290 -38575 8325
rect -38540 8290 -38530 8325
rect -38495 8290 -38485 8325
rect -38450 8290 -38440 8325
rect -38405 8290 -38395 8325
rect -38360 8290 -38350 8325
rect -38315 8290 -38305 8325
rect -38270 8290 -38260 8325
rect -38225 8290 -38215 8325
rect -38180 8290 -38170 8325
rect -38135 8290 -38125 8325
rect -38090 8290 -38080 8325
rect -38045 8290 -38035 8325
rect -38000 8290 -37990 8325
rect -37955 8290 -37945 8325
rect -37910 8290 -37900 8325
rect -37865 8290 -37855 8325
rect -37820 8290 -37810 8325
rect -37775 8290 -37765 8325
rect -37730 8290 -37720 8325
rect -37685 8290 -37675 8325
rect -37640 8290 -37630 8325
rect -37595 8290 -37585 8325
rect -37550 8290 -37540 8325
rect -37505 8290 -37495 8325
rect -37460 8290 -37450 8325
rect -37415 8290 -37405 8325
rect -37370 8290 -37360 8325
rect -37325 8290 -37315 8325
rect -37280 8290 -37270 8325
rect -37235 8290 -37225 8325
rect -37190 8305 7700 8325
rect -37190 8290 1320 8305
rect -38770 8280 1320 8290
rect -38770 8245 -38755 8280
rect -38720 8245 -38710 8280
rect -38675 8245 -38665 8280
rect -38630 8245 -38620 8280
rect -38585 8245 -38575 8280
rect -38540 8245 -38530 8280
rect -38495 8245 -38485 8280
rect -38450 8245 -38440 8280
rect -38405 8245 -38395 8280
rect -38360 8245 -38350 8280
rect -38315 8245 -38305 8280
rect -38270 8245 -38260 8280
rect -38225 8245 -38215 8280
rect -38180 8245 -38170 8280
rect -38135 8245 -38125 8280
rect -38090 8245 -38080 8280
rect -38045 8245 -38035 8280
rect -38000 8245 -37990 8280
rect -37955 8245 -37945 8280
rect -37910 8245 -37900 8280
rect -37865 8245 -37855 8280
rect -37820 8245 -37810 8280
rect -37775 8245 -37765 8280
rect -37730 8245 -37720 8280
rect -37685 8245 -37675 8280
rect -37640 8245 -37630 8280
rect -37595 8245 -37585 8280
rect -37550 8245 -37540 8280
rect -37505 8245 -37495 8280
rect -37460 8245 -37450 8280
rect -37415 8245 -37405 8280
rect -37370 8245 -37360 8280
rect -37325 8245 -37315 8280
rect -37280 8245 -37270 8280
rect -37235 8245 -37225 8280
rect -37190 8265 1320 8280
rect 1360 8265 2245 8305
rect 2285 8265 6700 8305
rect 6740 8265 7620 8305
rect 7660 8265 7700 8305
rect -37190 8245 7700 8265
rect -38770 8235 7700 8245
rect -38770 8200 -38755 8235
rect -38720 8200 -38710 8235
rect -38675 8200 -38665 8235
rect -38630 8200 -38620 8235
rect -38585 8200 -38575 8235
rect -38540 8200 -38530 8235
rect -38495 8200 -38485 8235
rect -38450 8200 -38440 8235
rect -38405 8200 -38395 8235
rect -38360 8200 -38350 8235
rect -38315 8200 -38305 8235
rect -38270 8200 -38260 8235
rect -38225 8200 -38215 8235
rect -38180 8200 -38170 8235
rect -38135 8200 -38125 8235
rect -38090 8200 -38080 8235
rect -38045 8200 -38035 8235
rect -38000 8200 -37990 8235
rect -37955 8200 -37945 8235
rect -37910 8200 -37900 8235
rect -37865 8200 -37855 8235
rect -37820 8200 -37810 8235
rect -37775 8200 -37765 8235
rect -37730 8200 -37720 8235
rect -37685 8200 -37675 8235
rect -37640 8200 -37630 8235
rect -37595 8200 -37585 8235
rect -37550 8200 -37540 8235
rect -37505 8200 -37495 8235
rect -37460 8200 -37450 8235
rect -37415 8200 -37405 8235
rect -37370 8200 -37360 8235
rect -37325 8200 -37315 8235
rect -37280 8200 -37270 8235
rect -37235 8200 -37225 8235
rect -37190 8200 1320 8235
rect -38770 8195 1320 8200
rect 1360 8195 2245 8235
rect 2285 8195 6700 8235
rect 6740 8195 7620 8235
rect 7660 8195 7700 8235
rect -38770 8190 7700 8195
rect -38770 8155 -38755 8190
rect -38720 8155 -38710 8190
rect -38675 8155 -38665 8190
rect -38630 8155 -38620 8190
rect -38585 8155 -38575 8190
rect -38540 8155 -38530 8190
rect -38495 8155 -38485 8190
rect -38450 8155 -38440 8190
rect -38405 8155 -38395 8190
rect -38360 8155 -38350 8190
rect -38315 8155 -38305 8190
rect -38270 8155 -38260 8190
rect -38225 8155 -38215 8190
rect -38180 8155 -38170 8190
rect -38135 8155 -38125 8190
rect -38090 8155 -38080 8190
rect -38045 8155 -38035 8190
rect -38000 8155 -37990 8190
rect -37955 8155 -37945 8190
rect -37910 8155 -37900 8190
rect -37865 8155 -37855 8190
rect -37820 8155 -37810 8190
rect -37775 8155 -37765 8190
rect -37730 8155 -37720 8190
rect -37685 8155 -37675 8190
rect -37640 8155 -37630 8190
rect -37595 8155 -37585 8190
rect -37550 8155 -37540 8190
rect -37505 8155 -37495 8190
rect -37460 8155 -37450 8190
rect -37415 8155 -37405 8190
rect -37370 8155 -37360 8190
rect -37325 8155 -37315 8190
rect -37280 8155 -37270 8190
rect -37235 8155 -37225 8190
rect -37190 8165 7700 8190
rect -37190 8155 1320 8165
rect -38770 8145 1320 8155
rect -38770 8110 -38755 8145
rect -38720 8110 -38710 8145
rect -38675 8110 -38665 8145
rect -38630 8110 -38620 8145
rect -38585 8110 -38575 8145
rect -38540 8110 -38530 8145
rect -38495 8110 -38485 8145
rect -38450 8110 -38440 8145
rect -38405 8110 -38395 8145
rect -38360 8110 -38350 8145
rect -38315 8110 -38305 8145
rect -38270 8110 -38260 8145
rect -38225 8110 -38215 8145
rect -38180 8110 -38170 8145
rect -38135 8110 -38125 8145
rect -38090 8110 -38080 8145
rect -38045 8110 -38035 8145
rect -38000 8110 -37990 8145
rect -37955 8110 -37945 8145
rect -37910 8110 -37900 8145
rect -37865 8110 -37855 8145
rect -37820 8110 -37810 8145
rect -37775 8110 -37765 8145
rect -37730 8110 -37720 8145
rect -37685 8110 -37675 8145
rect -37640 8110 -37630 8145
rect -37595 8110 -37585 8145
rect -37550 8110 -37540 8145
rect -37505 8110 -37495 8145
rect -37460 8110 -37450 8145
rect -37415 8110 -37405 8145
rect -37370 8110 -37360 8145
rect -37325 8110 -37315 8145
rect -37280 8110 -37270 8145
rect -37235 8110 -37225 8145
rect -37190 8125 1320 8145
rect 1360 8125 2245 8165
rect 2285 8125 6700 8165
rect 6740 8125 7620 8165
rect 7660 8125 7700 8165
rect -37190 8110 7700 8125
rect -38770 8105 7700 8110
rect 31290 8030 35620 8050
rect 31290 7995 31305 8030
rect 31340 7995 31350 8030
rect 31385 7995 31395 8030
rect 31430 7995 31440 8030
rect 31475 7995 31485 8030
rect 31520 7995 31530 8030
rect 31565 7995 31575 8030
rect 31610 7995 31620 8030
rect 31655 7995 31665 8030
rect 31700 7995 31710 8030
rect 31745 7995 31755 8030
rect 31790 7995 31800 8030
rect 31835 7995 31845 8030
rect 31880 7995 31890 8030
rect 31925 7995 31935 8030
rect 31970 7995 31980 8030
rect 32015 7995 32025 8030
rect 32060 7995 32070 8030
rect 32105 7995 32115 8030
rect 32150 7995 32160 8030
rect 32195 7995 32205 8030
rect 32240 7995 32250 8030
rect 32285 7995 32295 8030
rect 32330 7995 32340 8030
rect 32375 7995 32385 8030
rect 32420 7995 32430 8030
rect 32465 7995 32475 8030
rect 32510 7995 32520 8030
rect 32555 7995 32565 8030
rect 32600 7995 32610 8030
rect 32645 7995 32655 8030
rect 32690 7995 32700 8030
rect 32735 7995 32745 8030
rect 32780 7995 32790 8030
rect 32825 7995 32835 8030
rect 32870 7995 35620 8030
rect 31290 7985 35620 7995
rect -38770 7970 3390 7980
rect -38770 7935 -38755 7970
rect -38720 7935 -38710 7970
rect -38675 7935 -38665 7970
rect -38630 7935 -38620 7970
rect -38585 7935 -38575 7970
rect -38540 7935 -38530 7970
rect -38495 7935 -38485 7970
rect -38450 7935 -38440 7970
rect -38405 7935 -38395 7970
rect -38360 7935 -38350 7970
rect -38315 7935 -38305 7970
rect -38270 7935 -38260 7970
rect -38225 7935 -38215 7970
rect -38180 7935 -38170 7970
rect -38135 7935 -38125 7970
rect -38090 7935 -38080 7970
rect -38045 7935 -38035 7970
rect -38000 7935 -37990 7970
rect -37955 7935 -37945 7970
rect -37910 7935 -37900 7970
rect -37865 7935 -37855 7970
rect -37820 7935 -37810 7970
rect -37775 7935 -37765 7970
rect -37730 7935 -37720 7970
rect -37685 7935 -37675 7970
rect -37640 7935 -37630 7970
rect -37595 7935 -37585 7970
rect -37550 7935 -37540 7970
rect -37505 7935 -37495 7970
rect -37460 7935 -37450 7970
rect -37415 7935 -37405 7970
rect -37370 7935 -37360 7970
rect -37325 7935 -37315 7970
rect -37280 7935 -37270 7970
rect -37235 7935 -37225 7970
rect -37190 7960 3390 7970
rect -37190 7935 3175 7960
rect -38770 7925 3175 7935
rect -38770 7890 -38755 7925
rect -38720 7890 -38710 7925
rect -38675 7890 -38665 7925
rect -38630 7890 -38620 7925
rect -38585 7890 -38575 7925
rect -38540 7890 -38530 7925
rect -38495 7890 -38485 7925
rect -38450 7890 -38440 7925
rect -38405 7890 -38395 7925
rect -38360 7890 -38350 7925
rect -38315 7890 -38305 7925
rect -38270 7890 -38260 7925
rect -38225 7890 -38215 7925
rect -38180 7890 -38170 7925
rect -38135 7890 -38125 7925
rect -38090 7890 -38080 7925
rect -38045 7890 -38035 7925
rect -38000 7890 -37990 7925
rect -37955 7890 -37945 7925
rect -37910 7890 -37900 7925
rect -37865 7890 -37855 7925
rect -37820 7890 -37810 7925
rect -37775 7890 -37765 7925
rect -37730 7890 -37720 7925
rect -37685 7890 -37675 7925
rect -37640 7890 -37630 7925
rect -37595 7890 -37585 7925
rect -37550 7890 -37540 7925
rect -37505 7890 -37495 7925
rect -37460 7890 -37450 7925
rect -37415 7890 -37405 7925
rect -37370 7890 -37360 7925
rect -37325 7890 -37315 7925
rect -37280 7890 -37270 7925
rect -37235 7890 -37225 7925
rect -37190 7920 3175 7925
rect 3215 7920 3235 7960
rect 3275 7920 3345 7960
rect 3385 7920 3390 7960
rect -37190 7890 3390 7920
rect -38770 7880 3175 7890
rect -38770 7845 -38755 7880
rect -38720 7845 -38710 7880
rect -38675 7845 -38665 7880
rect -38630 7845 -38620 7880
rect -38585 7845 -38575 7880
rect -38540 7845 -38530 7880
rect -38495 7845 -38485 7880
rect -38450 7845 -38440 7880
rect -38405 7845 -38395 7880
rect -38360 7845 -38350 7880
rect -38315 7845 -38305 7880
rect -38270 7845 -38260 7880
rect -38225 7845 -38215 7880
rect -38180 7845 -38170 7880
rect -38135 7845 -38125 7880
rect -38090 7845 -38080 7880
rect -38045 7845 -38035 7880
rect -38000 7845 -37990 7880
rect -37955 7845 -37945 7880
rect -37910 7845 -37900 7880
rect -37865 7845 -37855 7880
rect -37820 7845 -37810 7880
rect -37775 7845 -37765 7880
rect -37730 7845 -37720 7880
rect -37685 7845 -37675 7880
rect -37640 7845 -37630 7880
rect -37595 7845 -37585 7880
rect -37550 7845 -37540 7880
rect -37505 7845 -37495 7880
rect -37460 7845 -37450 7880
rect -37415 7845 -37405 7880
rect -37370 7845 -37360 7880
rect -37325 7845 -37315 7880
rect -37280 7845 -37270 7880
rect -37235 7845 -37225 7880
rect -37190 7850 3175 7880
rect 3215 7850 3235 7890
rect 3275 7850 3345 7890
rect 3385 7850 3390 7890
rect -37190 7845 3390 7850
rect -38770 7835 3390 7845
rect -38770 7800 -38755 7835
rect -38720 7800 -38710 7835
rect -38675 7800 -38665 7835
rect -38630 7800 -38620 7835
rect -38585 7800 -38575 7835
rect -38540 7800 -38530 7835
rect -38495 7800 -38485 7835
rect -38450 7800 -38440 7835
rect -38405 7800 -38395 7835
rect -38360 7800 -38350 7835
rect -38315 7800 -38305 7835
rect -38270 7800 -38260 7835
rect -38225 7800 -38215 7835
rect -38180 7800 -38170 7835
rect -38135 7800 -38125 7835
rect -38090 7800 -38080 7835
rect -38045 7800 -38035 7835
rect -38000 7800 -37990 7835
rect -37955 7800 -37945 7835
rect -37910 7800 -37900 7835
rect -37865 7800 -37855 7835
rect -37820 7800 -37810 7835
rect -37775 7800 -37765 7835
rect -37730 7800 -37720 7835
rect -37685 7800 -37675 7835
rect -37640 7800 -37630 7835
rect -37595 7800 -37585 7835
rect -37550 7800 -37540 7835
rect -37505 7800 -37495 7835
rect -37460 7800 -37450 7835
rect -37415 7800 -37405 7835
rect -37370 7800 -37360 7835
rect -37325 7800 -37315 7835
rect -37280 7800 -37270 7835
rect -37235 7800 -37225 7835
rect -37190 7820 3390 7835
rect -37190 7800 3175 7820
rect -38770 7790 3175 7800
rect -38770 7755 -38755 7790
rect -38720 7755 -38710 7790
rect -38675 7755 -38665 7790
rect -38630 7755 -38620 7790
rect -38585 7755 -38575 7790
rect -38540 7755 -38530 7790
rect -38495 7755 -38485 7790
rect -38450 7755 -38440 7790
rect -38405 7755 -38395 7790
rect -38360 7755 -38350 7790
rect -38315 7755 -38305 7790
rect -38270 7755 -38260 7790
rect -38225 7755 -38215 7790
rect -38180 7755 -38170 7790
rect -38135 7755 -38125 7790
rect -38090 7755 -38080 7790
rect -38045 7755 -38035 7790
rect -38000 7755 -37990 7790
rect -37955 7755 -37945 7790
rect -37910 7755 -37900 7790
rect -37865 7755 -37855 7790
rect -37820 7755 -37810 7790
rect -37775 7755 -37765 7790
rect -37730 7755 -37720 7790
rect -37685 7755 -37675 7790
rect -37640 7755 -37630 7790
rect -37595 7755 -37585 7790
rect -37550 7755 -37540 7790
rect -37505 7755 -37495 7790
rect -37460 7755 -37450 7790
rect -37415 7755 -37405 7790
rect -37370 7755 -37360 7790
rect -37325 7755 -37315 7790
rect -37280 7755 -37270 7790
rect -37235 7755 -37225 7790
rect -37190 7780 3175 7790
rect 3215 7780 3235 7820
rect 3275 7780 3345 7820
rect 3385 7780 3390 7820
rect -37190 7755 3390 7780
rect -38770 7750 3390 7755
rect -38770 7745 3175 7750
rect -38770 7710 -38755 7745
rect -38720 7710 -38710 7745
rect -38675 7710 -38665 7745
rect -38630 7710 -38620 7745
rect -38585 7710 -38575 7745
rect -38540 7710 -38530 7745
rect -38495 7710 -38485 7745
rect -38450 7710 -38440 7745
rect -38405 7710 -38395 7745
rect -38360 7710 -38350 7745
rect -38315 7710 -38305 7745
rect -38270 7710 -38260 7745
rect -38225 7710 -38215 7745
rect -38180 7710 -38170 7745
rect -38135 7710 -38125 7745
rect -38090 7710 -38080 7745
rect -38045 7710 -38035 7745
rect -38000 7710 -37990 7745
rect -37955 7710 -37945 7745
rect -37910 7710 -37900 7745
rect -37865 7710 -37855 7745
rect -37820 7710 -37810 7745
rect -37775 7710 -37765 7745
rect -37730 7710 -37720 7745
rect -37685 7710 -37675 7745
rect -37640 7710 -37630 7745
rect -37595 7710 -37585 7745
rect -37550 7710 -37540 7745
rect -37505 7710 -37495 7745
rect -37460 7710 -37450 7745
rect -37415 7710 -37405 7745
rect -37370 7710 -37360 7745
rect -37325 7710 -37315 7745
rect -37280 7710 -37270 7745
rect -37235 7710 -37225 7745
rect -37190 7710 3175 7745
rect 3215 7710 3235 7750
rect 3275 7710 3345 7750
rect 3385 7710 3390 7750
rect -38770 7700 3390 7710
rect -38770 7665 -38755 7700
rect -38720 7665 -38710 7700
rect -38675 7665 -38665 7700
rect -38630 7665 -38620 7700
rect -38585 7665 -38575 7700
rect -38540 7665 -38530 7700
rect -38495 7665 -38485 7700
rect -38450 7665 -38440 7700
rect -38405 7665 -38395 7700
rect -38360 7665 -38350 7700
rect -38315 7665 -38305 7700
rect -38270 7665 -38260 7700
rect -38225 7665 -38215 7700
rect -38180 7665 -38170 7700
rect -38135 7665 -38125 7700
rect -38090 7665 -38080 7700
rect -38045 7665 -38035 7700
rect -38000 7665 -37990 7700
rect -37955 7665 -37945 7700
rect -37910 7665 -37900 7700
rect -37865 7665 -37855 7700
rect -37820 7665 -37810 7700
rect -37775 7665 -37765 7700
rect -37730 7665 -37720 7700
rect -37685 7665 -37675 7700
rect -37640 7665 -37630 7700
rect -37595 7665 -37585 7700
rect -37550 7665 -37540 7700
rect -37505 7665 -37495 7700
rect -37460 7665 -37450 7700
rect -37415 7665 -37405 7700
rect -37370 7665 -37360 7700
rect -37325 7665 -37315 7700
rect -37280 7665 -37270 7700
rect -37235 7665 -37225 7700
rect -37190 7685 3390 7700
rect -37190 7665 3175 7685
rect -38770 7655 3175 7665
rect -38770 7620 -38755 7655
rect -38720 7620 -38710 7655
rect -38675 7620 -38665 7655
rect -38630 7620 -38620 7655
rect -38585 7620 -38575 7655
rect -38540 7620 -38530 7655
rect -38495 7620 -38485 7655
rect -38450 7620 -38440 7655
rect -38405 7620 -38395 7655
rect -38360 7620 -38350 7655
rect -38315 7620 -38305 7655
rect -38270 7620 -38260 7655
rect -38225 7620 -38215 7655
rect -38180 7620 -38170 7655
rect -38135 7620 -38125 7655
rect -38090 7620 -38080 7655
rect -38045 7620 -38035 7655
rect -38000 7620 -37990 7655
rect -37955 7620 -37945 7655
rect -37910 7620 -37900 7655
rect -37865 7620 -37855 7655
rect -37820 7620 -37810 7655
rect -37775 7620 -37765 7655
rect -37730 7620 -37720 7655
rect -37685 7620 -37675 7655
rect -37640 7620 -37630 7655
rect -37595 7620 -37585 7655
rect -37550 7620 -37540 7655
rect -37505 7620 -37495 7655
rect -37460 7620 -37450 7655
rect -37415 7620 -37405 7655
rect -37370 7620 -37360 7655
rect -37325 7620 -37315 7655
rect -37280 7620 -37270 7655
rect -37235 7620 -37225 7655
rect -37190 7645 3175 7655
rect 3215 7645 3235 7685
rect 3275 7645 3345 7685
rect 3385 7645 3390 7685
rect -37190 7625 3390 7645
rect -37190 7620 3175 7625
rect -38770 7610 3175 7620
rect -38770 7575 -38755 7610
rect -38720 7575 -38710 7610
rect -38675 7575 -38665 7610
rect -38630 7575 -38620 7610
rect -38585 7575 -38575 7610
rect -38540 7575 -38530 7610
rect -38495 7575 -38485 7610
rect -38450 7575 -38440 7610
rect -38405 7575 -38395 7610
rect -38360 7575 -38350 7610
rect -38315 7575 -38305 7610
rect -38270 7575 -38260 7610
rect -38225 7575 -38215 7610
rect -38180 7575 -38170 7610
rect -38135 7575 -38125 7610
rect -38090 7575 -38080 7610
rect -38045 7575 -38035 7610
rect -38000 7575 -37990 7610
rect -37955 7575 -37945 7610
rect -37910 7575 -37900 7610
rect -37865 7575 -37855 7610
rect -37820 7575 -37810 7610
rect -37775 7575 -37765 7610
rect -37730 7575 -37720 7610
rect -37685 7575 -37675 7610
rect -37640 7575 -37630 7610
rect -37595 7575 -37585 7610
rect -37550 7575 -37540 7610
rect -37505 7575 -37495 7610
rect -37460 7575 -37450 7610
rect -37415 7575 -37405 7610
rect -37370 7575 -37360 7610
rect -37325 7575 -37315 7610
rect -37280 7575 -37270 7610
rect -37235 7575 -37225 7610
rect -37190 7585 3175 7610
rect 3215 7585 3235 7625
rect 3275 7585 3345 7625
rect 3385 7585 3390 7625
rect -37190 7575 3390 7585
rect -38770 7565 3390 7575
rect -38770 7530 -38755 7565
rect -38720 7530 -38710 7565
rect -38675 7530 -38665 7565
rect -38630 7530 -38620 7565
rect -38585 7530 -38575 7565
rect -38540 7530 -38530 7565
rect -38495 7530 -38485 7565
rect -38450 7530 -38440 7565
rect -38405 7530 -38395 7565
rect -38360 7530 -38350 7565
rect -38315 7530 -38305 7565
rect -38270 7530 -38260 7565
rect -38225 7530 -38215 7565
rect -38180 7530 -38170 7565
rect -38135 7530 -38125 7565
rect -38090 7530 -38080 7565
rect -38045 7530 -38035 7565
rect -38000 7530 -37990 7565
rect -37955 7530 -37945 7565
rect -37910 7530 -37900 7565
rect -37865 7530 -37855 7565
rect -37820 7530 -37810 7565
rect -37775 7530 -37765 7565
rect -37730 7530 -37720 7565
rect -37685 7530 -37675 7565
rect -37640 7530 -37630 7565
rect -37595 7530 -37585 7565
rect -37550 7530 -37540 7565
rect -37505 7530 -37495 7565
rect -37460 7530 -37450 7565
rect -37415 7530 -37405 7565
rect -37370 7530 -37360 7565
rect -37325 7530 -37315 7565
rect -37280 7530 -37270 7565
rect -37235 7530 -37225 7565
rect -37190 7560 3390 7565
rect -37190 7530 3175 7560
rect -38770 7520 3175 7530
rect 3215 7520 3235 7560
rect 3275 7520 3345 7560
rect 3385 7520 3390 7560
rect -38770 7485 -38755 7520
rect -38720 7485 -38710 7520
rect -38675 7485 -38665 7520
rect -38630 7485 -38620 7520
rect -38585 7485 -38575 7520
rect -38540 7485 -38530 7520
rect -38495 7485 -38485 7520
rect -38450 7485 -38440 7520
rect -38405 7485 -38395 7520
rect -38360 7485 -38350 7520
rect -38315 7485 -38305 7520
rect -38270 7485 -38260 7520
rect -38225 7485 -38215 7520
rect -38180 7485 -38170 7520
rect -38135 7485 -38125 7520
rect -38090 7485 -38080 7520
rect -38045 7485 -38035 7520
rect -38000 7485 -37990 7520
rect -37955 7485 -37945 7520
rect -37910 7485 -37900 7520
rect -37865 7485 -37855 7520
rect -37820 7485 -37810 7520
rect -37775 7485 -37765 7520
rect -37730 7485 -37720 7520
rect -37685 7485 -37675 7520
rect -37640 7485 -37630 7520
rect -37595 7485 -37585 7520
rect -37550 7485 -37540 7520
rect -37505 7485 -37495 7520
rect -37460 7485 -37450 7520
rect -37415 7485 -37405 7520
rect -37370 7485 -37360 7520
rect -37325 7485 -37315 7520
rect -37280 7485 -37270 7520
rect -37235 7485 -37225 7520
rect -37190 7490 3390 7520
rect -37190 7485 3175 7490
rect -38770 7475 3175 7485
rect -38770 7440 -38755 7475
rect -38720 7440 -38710 7475
rect -38675 7440 -38665 7475
rect -38630 7440 -38620 7475
rect -38585 7440 -38575 7475
rect -38540 7440 -38530 7475
rect -38495 7440 -38485 7475
rect -38450 7440 -38440 7475
rect -38405 7440 -38395 7475
rect -38360 7440 -38350 7475
rect -38315 7440 -38305 7475
rect -38270 7440 -38260 7475
rect -38225 7440 -38215 7475
rect -38180 7440 -38170 7475
rect -38135 7440 -38125 7475
rect -38090 7440 -38080 7475
rect -38045 7440 -38035 7475
rect -38000 7440 -37990 7475
rect -37955 7440 -37945 7475
rect -37910 7440 -37900 7475
rect -37865 7440 -37855 7475
rect -37820 7440 -37810 7475
rect -37775 7440 -37765 7475
rect -37730 7440 -37720 7475
rect -37685 7440 -37675 7475
rect -37640 7440 -37630 7475
rect -37595 7440 -37585 7475
rect -37550 7440 -37540 7475
rect -37505 7440 -37495 7475
rect -37460 7440 -37450 7475
rect -37415 7440 -37405 7475
rect -37370 7440 -37360 7475
rect -37325 7440 -37315 7475
rect -37280 7440 -37270 7475
rect -37235 7440 -37225 7475
rect -37190 7450 3175 7475
rect 3215 7450 3235 7490
rect 3275 7450 3345 7490
rect 3385 7450 3390 7490
rect -37190 7440 3390 7450
rect -38770 7430 3390 7440
rect -38770 7395 -38755 7430
rect -38720 7395 -38710 7430
rect -38675 7395 -38665 7430
rect -38630 7395 -38620 7430
rect -38585 7395 -38575 7430
rect -38540 7395 -38530 7430
rect -38495 7395 -38485 7430
rect -38450 7395 -38440 7430
rect -38405 7395 -38395 7430
rect -38360 7395 -38350 7430
rect -38315 7395 -38305 7430
rect -38270 7395 -38260 7430
rect -38225 7395 -38215 7430
rect -38180 7395 -38170 7430
rect -38135 7395 -38125 7430
rect -38090 7395 -38080 7430
rect -38045 7395 -38035 7430
rect -38000 7395 -37990 7430
rect -37955 7395 -37945 7430
rect -37910 7395 -37900 7430
rect -37865 7395 -37855 7430
rect -37820 7395 -37810 7430
rect -37775 7395 -37765 7430
rect -37730 7395 -37720 7430
rect -37685 7395 -37675 7430
rect -37640 7395 -37630 7430
rect -37595 7395 -37585 7430
rect -37550 7395 -37540 7430
rect -37505 7395 -37495 7430
rect -37460 7395 -37450 7430
rect -37415 7395 -37405 7430
rect -37370 7395 -37360 7430
rect -37325 7395 -37315 7430
rect -37280 7395 -37270 7430
rect -37235 7395 -37225 7430
rect -37190 7420 3390 7430
rect -37190 7395 3175 7420
rect -38770 7385 3175 7395
rect -38770 7350 -38755 7385
rect -38720 7350 -38710 7385
rect -38675 7350 -38665 7385
rect -38630 7350 -38620 7385
rect -38585 7350 -38575 7385
rect -38540 7350 -38530 7385
rect -38495 7350 -38485 7385
rect -38450 7350 -38440 7385
rect -38405 7350 -38395 7385
rect -38360 7350 -38350 7385
rect -38315 7350 -38305 7385
rect -38270 7350 -38260 7385
rect -38225 7350 -38215 7385
rect -38180 7350 -38170 7385
rect -38135 7350 -38125 7385
rect -38090 7350 -38080 7385
rect -38045 7350 -38035 7385
rect -38000 7350 -37990 7385
rect -37955 7350 -37945 7385
rect -37910 7350 -37900 7385
rect -37865 7350 -37855 7385
rect -37820 7350 -37810 7385
rect -37775 7350 -37765 7385
rect -37730 7350 -37720 7385
rect -37685 7350 -37675 7385
rect -37640 7350 -37630 7385
rect -37595 7350 -37585 7385
rect -37550 7350 -37540 7385
rect -37505 7350 -37495 7385
rect -37460 7350 -37450 7385
rect -37415 7350 -37405 7385
rect -37370 7350 -37360 7385
rect -37325 7350 -37315 7385
rect -37280 7350 -37270 7385
rect -37235 7350 -37225 7385
rect -37190 7380 3175 7385
rect 3215 7380 3235 7420
rect 3275 7380 3345 7420
rect 3385 7380 3390 7420
rect -37190 7350 3390 7380
rect -38770 7340 3175 7350
rect -38770 7305 -38755 7340
rect -38720 7305 -38710 7340
rect -38675 7305 -38665 7340
rect -38630 7305 -38620 7340
rect -38585 7305 -38575 7340
rect -38540 7305 -38530 7340
rect -38495 7305 -38485 7340
rect -38450 7305 -38440 7340
rect -38405 7305 -38395 7340
rect -38360 7305 -38350 7340
rect -38315 7305 -38305 7340
rect -38270 7305 -38260 7340
rect -38225 7305 -38215 7340
rect -38180 7305 -38170 7340
rect -38135 7305 -38125 7340
rect -38090 7305 -38080 7340
rect -38045 7305 -38035 7340
rect -38000 7305 -37990 7340
rect -37955 7305 -37945 7340
rect -37910 7305 -37900 7340
rect -37865 7305 -37855 7340
rect -37820 7305 -37810 7340
rect -37775 7305 -37765 7340
rect -37730 7305 -37720 7340
rect -37685 7305 -37675 7340
rect -37640 7305 -37630 7340
rect -37595 7305 -37585 7340
rect -37550 7305 -37540 7340
rect -37505 7305 -37495 7340
rect -37460 7305 -37450 7340
rect -37415 7305 -37405 7340
rect -37370 7305 -37360 7340
rect -37325 7305 -37315 7340
rect -37280 7305 -37270 7340
rect -37235 7305 -37225 7340
rect -37190 7310 3175 7340
rect 3215 7310 3235 7350
rect 3275 7310 3345 7350
rect 3385 7310 3390 7350
rect -37190 7305 3390 7310
rect -38770 7295 3390 7305
rect -38770 7260 -38755 7295
rect -38720 7260 -38710 7295
rect -38675 7260 -38665 7295
rect -38630 7260 -38620 7295
rect -38585 7260 -38575 7295
rect -38540 7260 -38530 7295
rect -38495 7260 -38485 7295
rect -38450 7260 -38440 7295
rect -38405 7260 -38395 7295
rect -38360 7260 -38350 7295
rect -38315 7260 -38305 7295
rect -38270 7260 -38260 7295
rect -38225 7260 -38215 7295
rect -38180 7260 -38170 7295
rect -38135 7260 -38125 7295
rect -38090 7260 -38080 7295
rect -38045 7260 -38035 7295
rect -38000 7260 -37990 7295
rect -37955 7260 -37945 7295
rect -37910 7260 -37900 7295
rect -37865 7260 -37855 7295
rect -37820 7260 -37810 7295
rect -37775 7260 -37765 7295
rect -37730 7260 -37720 7295
rect -37685 7260 -37675 7295
rect -37640 7260 -37630 7295
rect -37595 7260 -37585 7295
rect -37550 7260 -37540 7295
rect -37505 7260 -37495 7295
rect -37460 7260 -37450 7295
rect -37415 7260 -37405 7295
rect -37370 7260 -37360 7295
rect -37325 7260 -37315 7295
rect -37280 7260 -37270 7295
rect -37235 7260 -37225 7295
rect -37190 7285 3390 7295
rect -37190 7260 3175 7285
rect -38770 7250 3175 7260
rect -38770 7215 -38755 7250
rect -38720 7215 -38710 7250
rect -38675 7215 -38665 7250
rect -38630 7215 -38620 7250
rect -38585 7215 -38575 7250
rect -38540 7215 -38530 7250
rect -38495 7215 -38485 7250
rect -38450 7215 -38440 7250
rect -38405 7215 -38395 7250
rect -38360 7215 -38350 7250
rect -38315 7215 -38305 7250
rect -38270 7215 -38260 7250
rect -38225 7215 -38215 7250
rect -38180 7215 -38170 7250
rect -38135 7215 -38125 7250
rect -38090 7215 -38080 7250
rect -38045 7215 -38035 7250
rect -38000 7215 -37990 7250
rect -37955 7215 -37945 7250
rect -37910 7215 -37900 7250
rect -37865 7215 -37855 7250
rect -37820 7215 -37810 7250
rect -37775 7215 -37765 7250
rect -37730 7215 -37720 7250
rect -37685 7215 -37675 7250
rect -37640 7215 -37630 7250
rect -37595 7215 -37585 7250
rect -37550 7215 -37540 7250
rect -37505 7215 -37495 7250
rect -37460 7215 -37450 7250
rect -37415 7215 -37405 7250
rect -37370 7215 -37360 7250
rect -37325 7215 -37315 7250
rect -37280 7215 -37270 7250
rect -37235 7215 -37225 7250
rect -37190 7245 3175 7250
rect 3215 7245 3235 7285
rect 3275 7245 3345 7285
rect 3385 7245 3390 7285
rect -37190 7225 3390 7245
rect -37190 7215 3175 7225
rect -38770 7205 3175 7215
rect -38770 7170 -38755 7205
rect -38720 7170 -38710 7205
rect -38675 7170 -38665 7205
rect -38630 7170 -38620 7205
rect -38585 7170 -38575 7205
rect -38540 7170 -38530 7205
rect -38495 7170 -38485 7205
rect -38450 7170 -38440 7205
rect -38405 7170 -38395 7205
rect -38360 7170 -38350 7205
rect -38315 7170 -38305 7205
rect -38270 7170 -38260 7205
rect -38225 7170 -38215 7205
rect -38180 7170 -38170 7205
rect -38135 7170 -38125 7205
rect -38090 7170 -38080 7205
rect -38045 7170 -38035 7205
rect -38000 7170 -37990 7205
rect -37955 7170 -37945 7205
rect -37910 7170 -37900 7205
rect -37865 7170 -37855 7205
rect -37820 7170 -37810 7205
rect -37775 7170 -37765 7205
rect -37730 7170 -37720 7205
rect -37685 7170 -37675 7205
rect -37640 7170 -37630 7205
rect -37595 7170 -37585 7205
rect -37550 7170 -37540 7205
rect -37505 7170 -37495 7205
rect -37460 7170 -37450 7205
rect -37415 7170 -37405 7205
rect -37370 7170 -37360 7205
rect -37325 7170 -37315 7205
rect -37280 7170 -37270 7205
rect -37235 7170 -37225 7205
rect -37190 7185 3175 7205
rect 3215 7185 3235 7225
rect 3275 7185 3345 7225
rect 3385 7185 3390 7225
rect -37190 7170 3390 7185
rect -38770 7160 3390 7170
rect -38770 7125 -38755 7160
rect -38720 7125 -38710 7160
rect -38675 7125 -38665 7160
rect -38630 7125 -38620 7160
rect -38585 7125 -38575 7160
rect -38540 7125 -38530 7160
rect -38495 7125 -38485 7160
rect -38450 7125 -38440 7160
rect -38405 7125 -38395 7160
rect -38360 7125 -38350 7160
rect -38315 7125 -38305 7160
rect -38270 7125 -38260 7160
rect -38225 7125 -38215 7160
rect -38180 7125 -38170 7160
rect -38135 7125 -38125 7160
rect -38090 7125 -38080 7160
rect -38045 7125 -38035 7160
rect -38000 7125 -37990 7160
rect -37955 7125 -37945 7160
rect -37910 7125 -37900 7160
rect -37865 7125 -37855 7160
rect -37820 7125 -37810 7160
rect -37775 7125 -37765 7160
rect -37730 7125 -37720 7160
rect -37685 7125 -37675 7160
rect -37640 7125 -37630 7160
rect -37595 7125 -37585 7160
rect -37550 7125 -37540 7160
rect -37505 7125 -37495 7160
rect -37460 7125 -37450 7160
rect -37415 7125 -37405 7160
rect -37370 7125 -37360 7160
rect -37325 7125 -37315 7160
rect -37280 7125 -37270 7160
rect -37235 7125 -37225 7160
rect -37190 7125 3175 7160
rect -38770 7120 3175 7125
rect 3215 7120 3235 7160
rect 3275 7120 3345 7160
rect 3385 7120 3390 7160
rect -38770 7115 3390 7120
rect -38770 7080 -38755 7115
rect -38720 7080 -38710 7115
rect -38675 7080 -38665 7115
rect -38630 7080 -38620 7115
rect -38585 7080 -38575 7115
rect -38540 7080 -38530 7115
rect -38495 7080 -38485 7115
rect -38450 7080 -38440 7115
rect -38405 7080 -38395 7115
rect -38360 7080 -38350 7115
rect -38315 7080 -38305 7115
rect -38270 7080 -38260 7115
rect -38225 7080 -38215 7115
rect -38180 7080 -38170 7115
rect -38135 7080 -38125 7115
rect -38090 7080 -38080 7115
rect -38045 7080 -38035 7115
rect -38000 7080 -37990 7115
rect -37955 7080 -37945 7115
rect -37910 7080 -37900 7115
rect -37865 7080 -37855 7115
rect -37820 7080 -37810 7115
rect -37775 7080 -37765 7115
rect -37730 7080 -37720 7115
rect -37685 7080 -37675 7115
rect -37640 7080 -37630 7115
rect -37595 7080 -37585 7115
rect -37550 7080 -37540 7115
rect -37505 7080 -37495 7115
rect -37460 7080 -37450 7115
rect -37415 7080 -37405 7115
rect -37370 7080 -37360 7115
rect -37325 7080 -37315 7115
rect -37280 7080 -37270 7115
rect -37235 7080 -37225 7115
rect -37190 7090 3390 7115
rect -37190 7080 3175 7090
rect -38770 7070 3175 7080
rect -38770 7035 -38755 7070
rect -38720 7035 -38710 7070
rect -38675 7035 -38665 7070
rect -38630 7035 -38620 7070
rect -38585 7035 -38575 7070
rect -38540 7035 -38530 7070
rect -38495 7035 -38485 7070
rect -38450 7035 -38440 7070
rect -38405 7035 -38395 7070
rect -38360 7035 -38350 7070
rect -38315 7035 -38305 7070
rect -38270 7035 -38260 7070
rect -38225 7035 -38215 7070
rect -38180 7035 -38170 7070
rect -38135 7035 -38125 7070
rect -38090 7035 -38080 7070
rect -38045 7035 -38035 7070
rect -38000 7035 -37990 7070
rect -37955 7035 -37945 7070
rect -37910 7035 -37900 7070
rect -37865 7035 -37855 7070
rect -37820 7035 -37810 7070
rect -37775 7035 -37765 7070
rect -37730 7035 -37720 7070
rect -37685 7035 -37675 7070
rect -37640 7035 -37630 7070
rect -37595 7035 -37585 7070
rect -37550 7035 -37540 7070
rect -37505 7035 -37495 7070
rect -37460 7035 -37450 7070
rect -37415 7035 -37405 7070
rect -37370 7035 -37360 7070
rect -37325 7035 -37315 7070
rect -37280 7035 -37270 7070
rect -37235 7035 -37225 7070
rect -37190 7050 3175 7070
rect 3215 7050 3235 7090
rect 3275 7050 3345 7090
rect 3385 7050 3390 7090
rect -37190 7035 3390 7050
rect -38770 7025 3390 7035
rect -38770 6990 -38755 7025
rect -38720 6990 -38710 7025
rect -38675 6990 -38665 7025
rect -38630 6990 -38620 7025
rect -38585 6990 -38575 7025
rect -38540 6990 -38530 7025
rect -38495 6990 -38485 7025
rect -38450 6990 -38440 7025
rect -38405 6990 -38395 7025
rect -38360 6990 -38350 7025
rect -38315 6990 -38305 7025
rect -38270 6990 -38260 7025
rect -38225 6990 -38215 7025
rect -38180 6990 -38170 7025
rect -38135 6990 -38125 7025
rect -38090 6990 -38080 7025
rect -38045 6990 -38035 7025
rect -38000 6990 -37990 7025
rect -37955 6990 -37945 7025
rect -37910 6990 -37900 7025
rect -37865 6990 -37855 7025
rect -37820 6990 -37810 7025
rect -37775 6990 -37765 7025
rect -37730 6990 -37720 7025
rect -37685 6990 -37675 7025
rect -37640 6990 -37630 7025
rect -37595 6990 -37585 7025
rect -37550 6990 -37540 7025
rect -37505 6990 -37495 7025
rect -37460 6990 -37450 7025
rect -37415 6990 -37405 7025
rect -37370 6990 -37360 7025
rect -37325 6990 -37315 7025
rect -37280 6990 -37270 7025
rect -37235 6990 -37225 7025
rect -37190 7020 3390 7025
rect -37190 6990 3175 7020
rect -38770 6980 3175 6990
rect 3215 6980 3235 7020
rect 3275 6980 3345 7020
rect 3385 6980 3390 7020
rect -38770 6945 -38755 6980
rect -38720 6945 -38710 6980
rect -38675 6945 -38665 6980
rect -38630 6945 -38620 6980
rect -38585 6945 -38575 6980
rect -38540 6945 -38530 6980
rect -38495 6945 -38485 6980
rect -38450 6945 -38440 6980
rect -38405 6945 -38395 6980
rect -38360 6945 -38350 6980
rect -38315 6945 -38305 6980
rect -38270 6945 -38260 6980
rect -38225 6945 -38215 6980
rect -38180 6945 -38170 6980
rect -38135 6945 -38125 6980
rect -38090 6945 -38080 6980
rect -38045 6945 -38035 6980
rect -38000 6945 -37990 6980
rect -37955 6945 -37945 6980
rect -37910 6945 -37900 6980
rect -37865 6945 -37855 6980
rect -37820 6945 -37810 6980
rect -37775 6945 -37765 6980
rect -37730 6945 -37720 6980
rect -37685 6945 -37675 6980
rect -37640 6945 -37630 6980
rect -37595 6945 -37585 6980
rect -37550 6945 -37540 6980
rect -37505 6945 -37495 6980
rect -37460 6945 -37450 6980
rect -37415 6945 -37405 6980
rect -37370 6945 -37360 6980
rect -37325 6945 -37315 6980
rect -37280 6945 -37270 6980
rect -37235 6945 -37225 6980
rect -37190 6950 3390 6980
rect -37190 6945 3175 6950
rect -38770 6935 3175 6945
rect -38770 6900 -38755 6935
rect -38720 6900 -38710 6935
rect -38675 6900 -38665 6935
rect -38630 6900 -38620 6935
rect -38585 6900 -38575 6935
rect -38540 6900 -38530 6935
rect -38495 6900 -38485 6935
rect -38450 6900 -38440 6935
rect -38405 6900 -38395 6935
rect -38360 6900 -38350 6935
rect -38315 6900 -38305 6935
rect -38270 6900 -38260 6935
rect -38225 6900 -38215 6935
rect -38180 6900 -38170 6935
rect -38135 6900 -38125 6935
rect -38090 6900 -38080 6935
rect -38045 6900 -38035 6935
rect -38000 6900 -37990 6935
rect -37955 6900 -37945 6935
rect -37910 6900 -37900 6935
rect -37865 6900 -37855 6935
rect -37820 6900 -37810 6935
rect -37775 6900 -37765 6935
rect -37730 6900 -37720 6935
rect -37685 6900 -37675 6935
rect -37640 6900 -37630 6935
rect -37595 6900 -37585 6935
rect -37550 6900 -37540 6935
rect -37505 6900 -37495 6935
rect -37460 6900 -37450 6935
rect -37415 6900 -37405 6935
rect -37370 6900 -37360 6935
rect -37325 6900 -37315 6935
rect -37280 6900 -37270 6935
rect -37235 6900 -37225 6935
rect -37190 6910 3175 6935
rect 3215 6910 3235 6950
rect 3275 6910 3345 6950
rect 3385 6910 3390 6950
rect -37190 6900 3390 6910
rect -38770 6890 3390 6900
rect -38770 6855 -38755 6890
rect -38720 6855 -38710 6890
rect -38675 6855 -38665 6890
rect -38630 6855 -38620 6890
rect -38585 6855 -38575 6890
rect -38540 6855 -38530 6890
rect -38495 6855 -38485 6890
rect -38450 6855 -38440 6890
rect -38405 6855 -38395 6890
rect -38360 6855 -38350 6890
rect -38315 6855 -38305 6890
rect -38270 6855 -38260 6890
rect -38225 6855 -38215 6890
rect -38180 6855 -38170 6890
rect -38135 6855 -38125 6890
rect -38090 6855 -38080 6890
rect -38045 6855 -38035 6890
rect -38000 6855 -37990 6890
rect -37955 6855 -37945 6890
rect -37910 6855 -37900 6890
rect -37865 6855 -37855 6890
rect -37820 6855 -37810 6890
rect -37775 6855 -37765 6890
rect -37730 6855 -37720 6890
rect -37685 6855 -37675 6890
rect -37640 6855 -37630 6890
rect -37595 6855 -37585 6890
rect -37550 6855 -37540 6890
rect -37505 6855 -37495 6890
rect -37460 6855 -37450 6890
rect -37415 6855 -37405 6890
rect -37370 6855 -37360 6890
rect -37325 6855 -37315 6890
rect -37280 6855 -37270 6890
rect -37235 6855 -37225 6890
rect -37190 6885 3390 6890
rect -37190 6855 3175 6885
rect -38770 6845 3175 6855
rect 3215 6845 3235 6885
rect 3275 6845 3345 6885
rect 3385 6845 3390 6885
rect -38770 6810 -38755 6845
rect -38720 6810 -38710 6845
rect -38675 6810 -38665 6845
rect -38630 6810 -38620 6845
rect -38585 6810 -38575 6845
rect -38540 6810 -38530 6845
rect -38495 6810 -38485 6845
rect -38450 6810 -38440 6845
rect -38405 6810 -38395 6845
rect -38360 6810 -38350 6845
rect -38315 6810 -38305 6845
rect -38270 6810 -38260 6845
rect -38225 6810 -38215 6845
rect -38180 6810 -38170 6845
rect -38135 6810 -38125 6845
rect -38090 6810 -38080 6845
rect -38045 6810 -38035 6845
rect -38000 6810 -37990 6845
rect -37955 6810 -37945 6845
rect -37910 6810 -37900 6845
rect -37865 6810 -37855 6845
rect -37820 6810 -37810 6845
rect -37775 6810 -37765 6845
rect -37730 6810 -37720 6845
rect -37685 6810 -37675 6845
rect -37640 6810 -37630 6845
rect -37595 6810 -37585 6845
rect -37550 6810 -37540 6845
rect -37505 6810 -37495 6845
rect -37460 6810 -37450 6845
rect -37415 6810 -37405 6845
rect -37370 6810 -37360 6845
rect -37325 6810 -37315 6845
rect -37280 6810 -37270 6845
rect -37235 6810 -37225 6845
rect -37190 6825 3390 6845
rect -37190 6810 3175 6825
rect -38770 6800 3175 6810
rect -38770 6765 -38755 6800
rect -38720 6765 -38710 6800
rect -38675 6765 -38665 6800
rect -38630 6765 -38620 6800
rect -38585 6765 -38575 6800
rect -38540 6765 -38530 6800
rect -38495 6765 -38485 6800
rect -38450 6765 -38440 6800
rect -38405 6765 -38395 6800
rect -38360 6765 -38350 6800
rect -38315 6765 -38305 6800
rect -38270 6765 -38260 6800
rect -38225 6765 -38215 6800
rect -38180 6765 -38170 6800
rect -38135 6765 -38125 6800
rect -38090 6765 -38080 6800
rect -38045 6765 -38035 6800
rect -38000 6765 -37990 6800
rect -37955 6765 -37945 6800
rect -37910 6765 -37900 6800
rect -37865 6765 -37855 6800
rect -37820 6765 -37810 6800
rect -37775 6765 -37765 6800
rect -37730 6765 -37720 6800
rect -37685 6765 -37675 6800
rect -37640 6765 -37630 6800
rect -37595 6765 -37585 6800
rect -37550 6765 -37540 6800
rect -37505 6765 -37495 6800
rect -37460 6765 -37450 6800
rect -37415 6765 -37405 6800
rect -37370 6765 -37360 6800
rect -37325 6765 -37315 6800
rect -37280 6765 -37270 6800
rect -37235 6765 -37225 6800
rect -37190 6785 3175 6800
rect 3215 6785 3235 6825
rect 3275 6785 3345 6825
rect 3385 6785 3390 6825
rect -37190 6765 3390 6785
rect -38770 6760 3390 6765
rect -38770 6755 3175 6760
rect -38770 6720 -38755 6755
rect -38720 6720 -38710 6755
rect -38675 6720 -38665 6755
rect -38630 6720 -38620 6755
rect -38585 6720 -38575 6755
rect -38540 6720 -38530 6755
rect -38495 6720 -38485 6755
rect -38450 6720 -38440 6755
rect -38405 6720 -38395 6755
rect -38360 6720 -38350 6755
rect -38315 6720 -38305 6755
rect -38270 6720 -38260 6755
rect -38225 6720 -38215 6755
rect -38180 6720 -38170 6755
rect -38135 6720 -38125 6755
rect -38090 6720 -38080 6755
rect -38045 6720 -38035 6755
rect -38000 6720 -37990 6755
rect -37955 6720 -37945 6755
rect -37910 6720 -37900 6755
rect -37865 6720 -37855 6755
rect -37820 6720 -37810 6755
rect -37775 6720 -37765 6755
rect -37730 6720 -37720 6755
rect -37685 6720 -37675 6755
rect -37640 6720 -37630 6755
rect -37595 6720 -37585 6755
rect -37550 6720 -37540 6755
rect -37505 6720 -37495 6755
rect -37460 6720 -37450 6755
rect -37415 6720 -37405 6755
rect -37370 6720 -37360 6755
rect -37325 6720 -37315 6755
rect -37280 6720 -37270 6755
rect -37235 6720 -37225 6755
rect -37190 6720 3175 6755
rect 3215 6720 3235 6760
rect 3275 6720 3345 6760
rect 3385 6720 3390 6760
rect -38770 6710 3390 6720
rect -38770 6675 -38755 6710
rect -38720 6675 -38710 6710
rect -38675 6675 -38665 6710
rect -38630 6675 -38620 6710
rect -38585 6675 -38575 6710
rect -38540 6675 -38530 6710
rect -38495 6675 -38485 6710
rect -38450 6675 -38440 6710
rect -38405 6675 -38395 6710
rect -38360 6675 -38350 6710
rect -38315 6675 -38305 6710
rect -38270 6675 -38260 6710
rect -38225 6675 -38215 6710
rect -38180 6675 -38170 6710
rect -38135 6675 -38125 6710
rect -38090 6675 -38080 6710
rect -38045 6675 -38035 6710
rect -38000 6675 -37990 6710
rect -37955 6675 -37945 6710
rect -37910 6675 -37900 6710
rect -37865 6675 -37855 6710
rect -37820 6675 -37810 6710
rect -37775 6675 -37765 6710
rect -37730 6675 -37720 6710
rect -37685 6675 -37675 6710
rect -37640 6675 -37630 6710
rect -37595 6675 -37585 6710
rect -37550 6675 -37540 6710
rect -37505 6675 -37495 6710
rect -37460 6675 -37450 6710
rect -37415 6675 -37405 6710
rect -37370 6675 -37360 6710
rect -37325 6675 -37315 6710
rect -37280 6675 -37270 6710
rect -37235 6675 -37225 6710
rect -37190 6690 3390 6710
rect -37190 6675 3175 6690
rect -38770 6665 3175 6675
rect -38770 6630 -38755 6665
rect -38720 6630 -38710 6665
rect -38675 6630 -38665 6665
rect -38630 6630 -38620 6665
rect -38585 6630 -38575 6665
rect -38540 6630 -38530 6665
rect -38495 6630 -38485 6665
rect -38450 6630 -38440 6665
rect -38405 6630 -38395 6665
rect -38360 6630 -38350 6665
rect -38315 6630 -38305 6665
rect -38270 6630 -38260 6665
rect -38225 6630 -38215 6665
rect -38180 6630 -38170 6665
rect -38135 6630 -38125 6665
rect -38090 6630 -38080 6665
rect -38045 6630 -38035 6665
rect -38000 6630 -37990 6665
rect -37955 6630 -37945 6665
rect -37910 6630 -37900 6665
rect -37865 6630 -37855 6665
rect -37820 6630 -37810 6665
rect -37775 6630 -37765 6665
rect -37730 6630 -37720 6665
rect -37685 6630 -37675 6665
rect -37640 6630 -37630 6665
rect -37595 6630 -37585 6665
rect -37550 6630 -37540 6665
rect -37505 6630 -37495 6665
rect -37460 6630 -37450 6665
rect -37415 6630 -37405 6665
rect -37370 6630 -37360 6665
rect -37325 6630 -37315 6665
rect -37280 6630 -37270 6665
rect -37235 6630 -37225 6665
rect -37190 6650 3175 6665
rect 3215 6650 3235 6690
rect 3275 6650 3345 6690
rect 3385 6650 3390 6690
rect -37190 6630 3390 6650
rect -38770 6620 3390 6630
rect -38770 6585 -38755 6620
rect -38720 6585 -38710 6620
rect -38675 6585 -38665 6620
rect -38630 6585 -38620 6620
rect -38585 6585 -38575 6620
rect -38540 6585 -38530 6620
rect -38495 6585 -38485 6620
rect -38450 6585 -38440 6620
rect -38405 6585 -38395 6620
rect -38360 6585 -38350 6620
rect -38315 6585 -38305 6620
rect -38270 6585 -38260 6620
rect -38225 6585 -38215 6620
rect -38180 6585 -38170 6620
rect -38135 6585 -38125 6620
rect -38090 6585 -38080 6620
rect -38045 6585 -38035 6620
rect -38000 6585 -37990 6620
rect -37955 6585 -37945 6620
rect -37910 6585 -37900 6620
rect -37865 6585 -37855 6620
rect -37820 6585 -37810 6620
rect -37775 6585 -37765 6620
rect -37730 6585 -37720 6620
rect -37685 6585 -37675 6620
rect -37640 6585 -37630 6620
rect -37595 6585 -37585 6620
rect -37550 6585 -37540 6620
rect -37505 6585 -37495 6620
rect -37460 6585 -37450 6620
rect -37415 6585 -37405 6620
rect -37370 6585 -37360 6620
rect -37325 6585 -37315 6620
rect -37280 6585 -37270 6620
rect -37235 6585 -37225 6620
rect -37190 6585 3175 6620
rect -38770 6580 3175 6585
rect 3215 6580 3235 6620
rect 3275 6580 3345 6620
rect 3385 6580 3390 6620
rect -38770 6575 3390 6580
rect -38770 6540 -38755 6575
rect -38720 6540 -38710 6575
rect -38675 6540 -38665 6575
rect -38630 6540 -38620 6575
rect -38585 6540 -38575 6575
rect -38540 6540 -38530 6575
rect -38495 6540 -38485 6575
rect -38450 6540 -38440 6575
rect -38405 6540 -38395 6575
rect -38360 6540 -38350 6575
rect -38315 6540 -38305 6575
rect -38270 6540 -38260 6575
rect -38225 6540 -38215 6575
rect -38180 6540 -38170 6575
rect -38135 6540 -38125 6575
rect -38090 6540 -38080 6575
rect -38045 6540 -38035 6575
rect -38000 6540 -37990 6575
rect -37955 6540 -37945 6575
rect -37910 6540 -37900 6575
rect -37865 6540 -37855 6575
rect -37820 6540 -37810 6575
rect -37775 6540 -37765 6575
rect -37730 6540 -37720 6575
rect -37685 6540 -37675 6575
rect -37640 6540 -37630 6575
rect -37595 6540 -37585 6575
rect -37550 6540 -37540 6575
rect -37505 6540 -37495 6575
rect -37460 6540 -37450 6575
rect -37415 6540 -37405 6575
rect -37370 6540 -37360 6575
rect -37325 6540 -37315 6575
rect -37280 6540 -37270 6575
rect -37235 6540 -37225 6575
rect -37190 6550 3390 6575
rect -37190 6540 3175 6550
rect -38770 6530 3175 6540
rect -38770 6495 -38755 6530
rect -38720 6495 -38710 6530
rect -38675 6495 -38665 6530
rect -38630 6495 -38620 6530
rect -38585 6495 -38575 6530
rect -38540 6495 -38530 6530
rect -38495 6495 -38485 6530
rect -38450 6495 -38440 6530
rect -38405 6495 -38395 6530
rect -38360 6495 -38350 6530
rect -38315 6495 -38305 6530
rect -38270 6495 -38260 6530
rect -38225 6495 -38215 6530
rect -38180 6495 -38170 6530
rect -38135 6495 -38125 6530
rect -38090 6495 -38080 6530
rect -38045 6495 -38035 6530
rect -38000 6495 -37990 6530
rect -37955 6495 -37945 6530
rect -37910 6495 -37900 6530
rect -37865 6495 -37855 6530
rect -37820 6495 -37810 6530
rect -37775 6495 -37765 6530
rect -37730 6495 -37720 6530
rect -37685 6495 -37675 6530
rect -37640 6495 -37630 6530
rect -37595 6495 -37585 6530
rect -37550 6495 -37540 6530
rect -37505 6495 -37495 6530
rect -37460 6495 -37450 6530
rect -37415 6495 -37405 6530
rect -37370 6495 -37360 6530
rect -37325 6495 -37315 6530
rect -37280 6495 -37270 6530
rect -37235 6495 -37225 6530
rect -37190 6510 3175 6530
rect 3215 6510 3235 6550
rect 3275 6510 3345 6550
rect 3385 6510 3390 6550
rect -37190 6495 3390 6510
rect -38770 6485 3390 6495
rect -38770 6450 -38755 6485
rect -38720 6450 -38710 6485
rect -38675 6450 -38665 6485
rect -38630 6450 -38620 6485
rect -38585 6450 -38575 6485
rect -38540 6450 -38530 6485
rect -38495 6450 -38485 6485
rect -38450 6450 -38440 6485
rect -38405 6450 -38395 6485
rect -38360 6450 -38350 6485
rect -38315 6450 -38305 6485
rect -38270 6450 -38260 6485
rect -38225 6450 -38215 6485
rect -38180 6450 -38170 6485
rect -38135 6450 -38125 6485
rect -38090 6450 -38080 6485
rect -38045 6450 -38035 6485
rect -38000 6450 -37990 6485
rect -37955 6450 -37945 6485
rect -37910 6450 -37900 6485
rect -37865 6450 -37855 6485
rect -37820 6450 -37810 6485
rect -37775 6450 -37765 6485
rect -37730 6450 -37720 6485
rect -37685 6450 -37675 6485
rect -37640 6450 -37630 6485
rect -37595 6450 -37585 6485
rect -37550 6450 -37540 6485
rect -37505 6450 -37495 6485
rect -37460 6450 -37450 6485
rect -37415 6450 -37405 6485
rect -37370 6450 -37360 6485
rect -37325 6450 -37315 6485
rect -37280 6450 -37270 6485
rect -37235 6450 -37225 6485
rect -37190 6450 3175 6485
rect -38770 6445 3175 6450
rect 3215 6445 3235 6485
rect 3275 6445 3345 6485
rect 3385 6445 3390 6485
rect 31290 7950 31305 7985
rect 31340 7950 31350 7985
rect 31385 7950 31395 7985
rect 31430 7950 31440 7985
rect 31475 7950 31485 7985
rect 31520 7950 31530 7985
rect 31565 7950 31575 7985
rect 31610 7950 31620 7985
rect 31655 7950 31665 7985
rect 31700 7950 31710 7985
rect 31745 7950 31755 7985
rect 31790 7950 31800 7985
rect 31835 7950 31845 7985
rect 31880 7950 31890 7985
rect 31925 7950 31935 7985
rect 31970 7950 31980 7985
rect 32015 7950 32025 7985
rect 32060 7950 32070 7985
rect 32105 7950 32115 7985
rect 32150 7950 32160 7985
rect 32195 7950 32205 7985
rect 32240 7950 32250 7985
rect 32285 7950 32295 7985
rect 32330 7950 32340 7985
rect 32375 7950 32385 7985
rect 32420 7950 32430 7985
rect 32465 7950 32475 7985
rect 32510 7950 32520 7985
rect 32555 7950 32565 7985
rect 32600 7950 32610 7985
rect 32645 7950 32655 7985
rect 32690 7950 32700 7985
rect 32735 7950 32745 7985
rect 32780 7950 32790 7985
rect 32825 7950 32835 7985
rect 32870 7950 35620 7985
rect 31290 7940 35620 7950
rect 31290 7905 31305 7940
rect 31340 7905 31350 7940
rect 31385 7905 31395 7940
rect 31430 7905 31440 7940
rect 31475 7905 31485 7940
rect 31520 7905 31530 7940
rect 31565 7905 31575 7940
rect 31610 7905 31620 7940
rect 31655 7905 31665 7940
rect 31700 7905 31710 7940
rect 31745 7905 31755 7940
rect 31790 7905 31800 7940
rect 31835 7905 31845 7940
rect 31880 7905 31890 7940
rect 31925 7905 31935 7940
rect 31970 7905 31980 7940
rect 32015 7905 32025 7940
rect 32060 7905 32070 7940
rect 32105 7905 32115 7940
rect 32150 7905 32160 7940
rect 32195 7905 32205 7940
rect 32240 7905 32250 7940
rect 32285 7905 32295 7940
rect 32330 7905 32340 7940
rect 32375 7905 32385 7940
rect 32420 7905 32430 7940
rect 32465 7905 32475 7940
rect 32510 7905 32520 7940
rect 32555 7905 32565 7940
rect 32600 7905 32610 7940
rect 32645 7905 32655 7940
rect 32690 7905 32700 7940
rect 32735 7905 32745 7940
rect 32780 7905 32790 7940
rect 32825 7905 32835 7940
rect 32870 7905 35620 7940
rect 31290 7895 35620 7905
rect 31290 7860 31305 7895
rect 31340 7860 31350 7895
rect 31385 7860 31395 7895
rect 31430 7860 31440 7895
rect 31475 7860 31485 7895
rect 31520 7860 31530 7895
rect 31565 7860 31575 7895
rect 31610 7860 31620 7895
rect 31655 7860 31665 7895
rect 31700 7860 31710 7895
rect 31745 7860 31755 7895
rect 31790 7860 31800 7895
rect 31835 7860 31845 7895
rect 31880 7860 31890 7895
rect 31925 7860 31935 7895
rect 31970 7860 31980 7895
rect 32015 7860 32025 7895
rect 32060 7860 32070 7895
rect 32105 7860 32115 7895
rect 32150 7860 32160 7895
rect 32195 7860 32205 7895
rect 32240 7860 32250 7895
rect 32285 7860 32295 7895
rect 32330 7860 32340 7895
rect 32375 7860 32385 7895
rect 32420 7860 32430 7895
rect 32465 7860 32475 7895
rect 32510 7860 32520 7895
rect 32555 7860 32565 7895
rect 32600 7860 32610 7895
rect 32645 7860 32655 7895
rect 32690 7860 32700 7895
rect 32735 7860 32745 7895
rect 32780 7860 32790 7895
rect 32825 7860 32835 7895
rect 32870 7860 35620 7895
rect 31290 7850 35620 7860
rect 31290 7815 31305 7850
rect 31340 7815 31350 7850
rect 31385 7815 31395 7850
rect 31430 7815 31440 7850
rect 31475 7815 31485 7850
rect 31520 7815 31530 7850
rect 31565 7815 31575 7850
rect 31610 7815 31620 7850
rect 31655 7815 31665 7850
rect 31700 7815 31710 7850
rect 31745 7815 31755 7850
rect 31790 7815 31800 7850
rect 31835 7815 31845 7850
rect 31880 7815 31890 7850
rect 31925 7815 31935 7850
rect 31970 7815 31980 7850
rect 32015 7815 32025 7850
rect 32060 7815 32070 7850
rect 32105 7815 32115 7850
rect 32150 7815 32160 7850
rect 32195 7815 32205 7850
rect 32240 7815 32250 7850
rect 32285 7815 32295 7850
rect 32330 7815 32340 7850
rect 32375 7815 32385 7850
rect 32420 7815 32430 7850
rect 32465 7815 32475 7850
rect 32510 7815 32520 7850
rect 32555 7815 32565 7850
rect 32600 7815 32610 7850
rect 32645 7815 32655 7850
rect 32690 7815 32700 7850
rect 32735 7815 32745 7850
rect 32780 7815 32790 7850
rect 32825 7815 32835 7850
rect 32870 7815 35620 7850
rect 31290 7805 35620 7815
rect 31290 7770 31305 7805
rect 31340 7770 31350 7805
rect 31385 7770 31395 7805
rect 31430 7770 31440 7805
rect 31475 7770 31485 7805
rect 31520 7770 31530 7805
rect 31565 7770 31575 7805
rect 31610 7770 31620 7805
rect 31655 7770 31665 7805
rect 31700 7770 31710 7805
rect 31745 7770 31755 7805
rect 31790 7770 31800 7805
rect 31835 7770 31845 7805
rect 31880 7770 31890 7805
rect 31925 7770 31935 7805
rect 31970 7770 31980 7805
rect 32015 7770 32025 7805
rect 32060 7770 32070 7805
rect 32105 7770 32115 7805
rect 32150 7770 32160 7805
rect 32195 7770 32205 7805
rect 32240 7770 32250 7805
rect 32285 7770 32295 7805
rect 32330 7770 32340 7805
rect 32375 7770 32385 7805
rect 32420 7770 32430 7805
rect 32465 7770 32475 7805
rect 32510 7770 32520 7805
rect 32555 7770 32565 7805
rect 32600 7770 32610 7805
rect 32645 7770 32655 7805
rect 32690 7770 32700 7805
rect 32735 7770 32745 7805
rect 32780 7770 32790 7805
rect 32825 7770 32835 7805
rect 32870 7770 35620 7805
rect 31290 7760 35620 7770
rect 31290 7725 31305 7760
rect 31340 7725 31350 7760
rect 31385 7725 31395 7760
rect 31430 7725 31440 7760
rect 31475 7725 31485 7760
rect 31520 7725 31530 7760
rect 31565 7725 31575 7760
rect 31610 7725 31620 7760
rect 31655 7725 31665 7760
rect 31700 7725 31710 7760
rect 31745 7725 31755 7760
rect 31790 7725 31800 7760
rect 31835 7725 31845 7760
rect 31880 7725 31890 7760
rect 31925 7725 31935 7760
rect 31970 7725 31980 7760
rect 32015 7725 32025 7760
rect 32060 7725 32070 7760
rect 32105 7725 32115 7760
rect 32150 7725 32160 7760
rect 32195 7725 32205 7760
rect 32240 7725 32250 7760
rect 32285 7725 32295 7760
rect 32330 7725 32340 7760
rect 32375 7725 32385 7760
rect 32420 7725 32430 7760
rect 32465 7725 32475 7760
rect 32510 7725 32520 7760
rect 32555 7725 32565 7760
rect 32600 7725 32610 7760
rect 32645 7725 32655 7760
rect 32690 7725 32700 7760
rect 32735 7725 32745 7760
rect 32780 7725 32790 7760
rect 32825 7725 32835 7760
rect 32870 7725 35620 7760
rect 31290 7715 35620 7725
rect 31290 7680 31305 7715
rect 31340 7680 31350 7715
rect 31385 7680 31395 7715
rect 31430 7680 31440 7715
rect 31475 7680 31485 7715
rect 31520 7680 31530 7715
rect 31565 7680 31575 7715
rect 31610 7680 31620 7715
rect 31655 7680 31665 7715
rect 31700 7680 31710 7715
rect 31745 7680 31755 7715
rect 31790 7680 31800 7715
rect 31835 7680 31845 7715
rect 31880 7680 31890 7715
rect 31925 7680 31935 7715
rect 31970 7680 31980 7715
rect 32015 7680 32025 7715
rect 32060 7680 32070 7715
rect 32105 7680 32115 7715
rect 32150 7680 32160 7715
rect 32195 7680 32205 7715
rect 32240 7680 32250 7715
rect 32285 7680 32295 7715
rect 32330 7680 32340 7715
rect 32375 7680 32385 7715
rect 32420 7680 32430 7715
rect 32465 7680 32475 7715
rect 32510 7680 32520 7715
rect 32555 7680 32565 7715
rect 32600 7680 32610 7715
rect 32645 7680 32655 7715
rect 32690 7680 32700 7715
rect 32735 7680 32745 7715
rect 32780 7680 32790 7715
rect 32825 7680 32835 7715
rect 32870 7680 35620 7715
rect 31290 7670 35620 7680
rect 31290 7635 31305 7670
rect 31340 7635 31350 7670
rect 31385 7635 31395 7670
rect 31430 7635 31440 7670
rect 31475 7635 31485 7670
rect 31520 7635 31530 7670
rect 31565 7635 31575 7670
rect 31610 7635 31620 7670
rect 31655 7635 31665 7670
rect 31700 7635 31710 7670
rect 31745 7635 31755 7670
rect 31790 7635 31800 7670
rect 31835 7635 31845 7670
rect 31880 7635 31890 7670
rect 31925 7635 31935 7670
rect 31970 7635 31980 7670
rect 32015 7635 32025 7670
rect 32060 7635 32070 7670
rect 32105 7635 32115 7670
rect 32150 7635 32160 7670
rect 32195 7635 32205 7670
rect 32240 7635 32250 7670
rect 32285 7635 32295 7670
rect 32330 7635 32340 7670
rect 32375 7635 32385 7670
rect 32420 7635 32430 7670
rect 32465 7635 32475 7670
rect 32510 7635 32520 7670
rect 32555 7635 32565 7670
rect 32600 7635 32610 7670
rect 32645 7635 32655 7670
rect 32690 7635 32700 7670
rect 32735 7635 32745 7670
rect 32780 7635 32790 7670
rect 32825 7635 32835 7670
rect 32870 7635 35620 7670
rect 31290 7625 35620 7635
rect 31290 7590 31305 7625
rect 31340 7590 31350 7625
rect 31385 7590 31395 7625
rect 31430 7590 31440 7625
rect 31475 7590 31485 7625
rect 31520 7590 31530 7625
rect 31565 7590 31575 7625
rect 31610 7590 31620 7625
rect 31655 7590 31665 7625
rect 31700 7590 31710 7625
rect 31745 7590 31755 7625
rect 31790 7590 31800 7625
rect 31835 7590 31845 7625
rect 31880 7590 31890 7625
rect 31925 7590 31935 7625
rect 31970 7590 31980 7625
rect 32015 7590 32025 7625
rect 32060 7590 32070 7625
rect 32105 7590 32115 7625
rect 32150 7590 32160 7625
rect 32195 7590 32205 7625
rect 32240 7590 32250 7625
rect 32285 7590 32295 7625
rect 32330 7590 32340 7625
rect 32375 7590 32385 7625
rect 32420 7590 32430 7625
rect 32465 7590 32475 7625
rect 32510 7590 32520 7625
rect 32555 7590 32565 7625
rect 32600 7590 32610 7625
rect 32645 7590 32655 7625
rect 32690 7590 32700 7625
rect 32735 7590 32745 7625
rect 32780 7590 32790 7625
rect 32825 7590 32835 7625
rect 32870 7590 35620 7625
rect 31290 7580 35620 7590
rect 31290 7545 31305 7580
rect 31340 7545 31350 7580
rect 31385 7545 31395 7580
rect 31430 7545 31440 7580
rect 31475 7545 31485 7580
rect 31520 7545 31530 7580
rect 31565 7545 31575 7580
rect 31610 7545 31620 7580
rect 31655 7545 31665 7580
rect 31700 7545 31710 7580
rect 31745 7545 31755 7580
rect 31790 7545 31800 7580
rect 31835 7545 31845 7580
rect 31880 7545 31890 7580
rect 31925 7545 31935 7580
rect 31970 7545 31980 7580
rect 32015 7545 32025 7580
rect 32060 7545 32070 7580
rect 32105 7545 32115 7580
rect 32150 7545 32160 7580
rect 32195 7545 32205 7580
rect 32240 7545 32250 7580
rect 32285 7545 32295 7580
rect 32330 7545 32340 7580
rect 32375 7545 32385 7580
rect 32420 7545 32430 7580
rect 32465 7545 32475 7580
rect 32510 7545 32520 7580
rect 32555 7545 32565 7580
rect 32600 7545 32610 7580
rect 32645 7545 32655 7580
rect 32690 7545 32700 7580
rect 32735 7545 32745 7580
rect 32780 7545 32790 7580
rect 32825 7545 32835 7580
rect 32870 7545 35620 7580
rect 31290 7535 35620 7545
rect 31290 7500 31305 7535
rect 31340 7500 31350 7535
rect 31385 7500 31395 7535
rect 31430 7500 31440 7535
rect 31475 7500 31485 7535
rect 31520 7500 31530 7535
rect 31565 7500 31575 7535
rect 31610 7500 31620 7535
rect 31655 7500 31665 7535
rect 31700 7500 31710 7535
rect 31745 7500 31755 7535
rect 31790 7500 31800 7535
rect 31835 7500 31845 7535
rect 31880 7500 31890 7535
rect 31925 7500 31935 7535
rect 31970 7500 31980 7535
rect 32015 7500 32025 7535
rect 32060 7500 32070 7535
rect 32105 7500 32115 7535
rect 32150 7500 32160 7535
rect 32195 7500 32205 7535
rect 32240 7500 32250 7535
rect 32285 7500 32295 7535
rect 32330 7500 32340 7535
rect 32375 7500 32385 7535
rect 32420 7500 32430 7535
rect 32465 7500 32475 7535
rect 32510 7500 32520 7535
rect 32555 7500 32565 7535
rect 32600 7500 32610 7535
rect 32645 7500 32655 7535
rect 32690 7500 32700 7535
rect 32735 7500 32745 7535
rect 32780 7500 32790 7535
rect 32825 7500 32835 7535
rect 32870 7500 35620 7535
rect 31290 7490 35620 7500
rect 31290 7455 31305 7490
rect 31340 7455 31350 7490
rect 31385 7455 31395 7490
rect 31430 7455 31440 7490
rect 31475 7455 31485 7490
rect 31520 7455 31530 7490
rect 31565 7455 31575 7490
rect 31610 7455 31620 7490
rect 31655 7455 31665 7490
rect 31700 7455 31710 7490
rect 31745 7455 31755 7490
rect 31790 7455 31800 7490
rect 31835 7455 31845 7490
rect 31880 7455 31890 7490
rect 31925 7455 31935 7490
rect 31970 7455 31980 7490
rect 32015 7455 32025 7490
rect 32060 7455 32070 7490
rect 32105 7455 32115 7490
rect 32150 7455 32160 7490
rect 32195 7455 32205 7490
rect 32240 7455 32250 7490
rect 32285 7455 32295 7490
rect 32330 7455 32340 7490
rect 32375 7455 32385 7490
rect 32420 7455 32430 7490
rect 32465 7455 32475 7490
rect 32510 7455 32520 7490
rect 32555 7455 32565 7490
rect 32600 7455 32610 7490
rect 32645 7455 32655 7490
rect 32690 7455 32700 7490
rect 32735 7455 32745 7490
rect 32780 7455 32790 7490
rect 32825 7455 32835 7490
rect 32870 7455 35620 7490
rect 31290 7445 35620 7455
rect 31290 7410 31305 7445
rect 31340 7410 31350 7445
rect 31385 7410 31395 7445
rect 31430 7410 31440 7445
rect 31475 7410 31485 7445
rect 31520 7410 31530 7445
rect 31565 7410 31575 7445
rect 31610 7410 31620 7445
rect 31655 7410 31665 7445
rect 31700 7410 31710 7445
rect 31745 7410 31755 7445
rect 31790 7410 31800 7445
rect 31835 7410 31845 7445
rect 31880 7410 31890 7445
rect 31925 7410 31935 7445
rect 31970 7410 31980 7445
rect 32015 7410 32025 7445
rect 32060 7410 32070 7445
rect 32105 7410 32115 7445
rect 32150 7410 32160 7445
rect 32195 7410 32205 7445
rect 32240 7410 32250 7445
rect 32285 7410 32295 7445
rect 32330 7410 32340 7445
rect 32375 7410 32385 7445
rect 32420 7410 32430 7445
rect 32465 7410 32475 7445
rect 32510 7410 32520 7445
rect 32555 7410 32565 7445
rect 32600 7410 32610 7445
rect 32645 7410 32655 7445
rect 32690 7410 32700 7445
rect 32735 7410 32745 7445
rect 32780 7410 32790 7445
rect 32825 7410 32835 7445
rect 32870 7410 35620 7445
rect 31290 7400 35620 7410
rect 31290 7365 31305 7400
rect 31340 7365 31350 7400
rect 31385 7365 31395 7400
rect 31430 7365 31440 7400
rect 31475 7365 31485 7400
rect 31520 7365 31530 7400
rect 31565 7365 31575 7400
rect 31610 7365 31620 7400
rect 31655 7365 31665 7400
rect 31700 7365 31710 7400
rect 31745 7365 31755 7400
rect 31790 7365 31800 7400
rect 31835 7365 31845 7400
rect 31880 7365 31890 7400
rect 31925 7365 31935 7400
rect 31970 7365 31980 7400
rect 32015 7365 32025 7400
rect 32060 7365 32070 7400
rect 32105 7365 32115 7400
rect 32150 7365 32160 7400
rect 32195 7365 32205 7400
rect 32240 7365 32250 7400
rect 32285 7365 32295 7400
rect 32330 7365 32340 7400
rect 32375 7365 32385 7400
rect 32420 7365 32430 7400
rect 32465 7365 32475 7400
rect 32510 7365 32520 7400
rect 32555 7365 32565 7400
rect 32600 7365 32610 7400
rect 32645 7365 32655 7400
rect 32690 7365 32700 7400
rect 32735 7365 32745 7400
rect 32780 7365 32790 7400
rect 32825 7365 32835 7400
rect 32870 7365 35620 7400
rect 31290 7355 35620 7365
rect 31290 7320 31305 7355
rect 31340 7320 31350 7355
rect 31385 7320 31395 7355
rect 31430 7320 31440 7355
rect 31475 7320 31485 7355
rect 31520 7320 31530 7355
rect 31565 7320 31575 7355
rect 31610 7320 31620 7355
rect 31655 7320 31665 7355
rect 31700 7320 31710 7355
rect 31745 7320 31755 7355
rect 31790 7320 31800 7355
rect 31835 7320 31845 7355
rect 31880 7320 31890 7355
rect 31925 7320 31935 7355
rect 31970 7320 31980 7355
rect 32015 7320 32025 7355
rect 32060 7320 32070 7355
rect 32105 7320 32115 7355
rect 32150 7320 32160 7355
rect 32195 7320 32205 7355
rect 32240 7320 32250 7355
rect 32285 7320 32295 7355
rect 32330 7320 32340 7355
rect 32375 7320 32385 7355
rect 32420 7320 32430 7355
rect 32465 7320 32475 7355
rect 32510 7320 32520 7355
rect 32555 7320 32565 7355
rect 32600 7320 32610 7355
rect 32645 7320 32655 7355
rect 32690 7320 32700 7355
rect 32735 7320 32745 7355
rect 32780 7320 32790 7355
rect 32825 7320 32835 7355
rect 32870 7320 35620 7355
rect 31290 7310 35620 7320
rect 31290 7275 31305 7310
rect 31340 7275 31350 7310
rect 31385 7275 31395 7310
rect 31430 7275 31440 7310
rect 31475 7275 31485 7310
rect 31520 7275 31530 7310
rect 31565 7275 31575 7310
rect 31610 7275 31620 7310
rect 31655 7275 31665 7310
rect 31700 7275 31710 7310
rect 31745 7275 31755 7310
rect 31790 7275 31800 7310
rect 31835 7275 31845 7310
rect 31880 7275 31890 7310
rect 31925 7275 31935 7310
rect 31970 7275 31980 7310
rect 32015 7275 32025 7310
rect 32060 7275 32070 7310
rect 32105 7275 32115 7310
rect 32150 7275 32160 7310
rect 32195 7275 32205 7310
rect 32240 7275 32250 7310
rect 32285 7275 32295 7310
rect 32330 7275 32340 7310
rect 32375 7275 32385 7310
rect 32420 7275 32430 7310
rect 32465 7275 32475 7310
rect 32510 7275 32520 7310
rect 32555 7275 32565 7310
rect 32600 7275 32610 7310
rect 32645 7275 32655 7310
rect 32690 7275 32700 7310
rect 32735 7275 32745 7310
rect 32780 7275 32790 7310
rect 32825 7275 32835 7310
rect 32870 7275 35620 7310
rect 31290 7265 35620 7275
rect 31290 7230 31305 7265
rect 31340 7230 31350 7265
rect 31385 7230 31395 7265
rect 31430 7230 31440 7265
rect 31475 7230 31485 7265
rect 31520 7230 31530 7265
rect 31565 7230 31575 7265
rect 31610 7230 31620 7265
rect 31655 7230 31665 7265
rect 31700 7230 31710 7265
rect 31745 7230 31755 7265
rect 31790 7230 31800 7265
rect 31835 7230 31845 7265
rect 31880 7230 31890 7265
rect 31925 7230 31935 7265
rect 31970 7230 31980 7265
rect 32015 7230 32025 7265
rect 32060 7230 32070 7265
rect 32105 7230 32115 7265
rect 32150 7230 32160 7265
rect 32195 7230 32205 7265
rect 32240 7230 32250 7265
rect 32285 7230 32295 7265
rect 32330 7230 32340 7265
rect 32375 7230 32385 7265
rect 32420 7230 32430 7265
rect 32465 7230 32475 7265
rect 32510 7230 32520 7265
rect 32555 7230 32565 7265
rect 32600 7230 32610 7265
rect 32645 7230 32655 7265
rect 32690 7230 32700 7265
rect 32735 7230 32745 7265
rect 32780 7230 32790 7265
rect 32825 7230 32835 7265
rect 32870 7230 35620 7265
rect 31290 7220 35620 7230
rect 31290 7185 31305 7220
rect 31340 7185 31350 7220
rect 31385 7185 31395 7220
rect 31430 7185 31440 7220
rect 31475 7185 31485 7220
rect 31520 7185 31530 7220
rect 31565 7185 31575 7220
rect 31610 7185 31620 7220
rect 31655 7185 31665 7220
rect 31700 7185 31710 7220
rect 31745 7185 31755 7220
rect 31790 7185 31800 7220
rect 31835 7185 31845 7220
rect 31880 7185 31890 7220
rect 31925 7185 31935 7220
rect 31970 7185 31980 7220
rect 32015 7185 32025 7220
rect 32060 7185 32070 7220
rect 32105 7185 32115 7220
rect 32150 7185 32160 7220
rect 32195 7185 32205 7220
rect 32240 7185 32250 7220
rect 32285 7185 32295 7220
rect 32330 7185 32340 7220
rect 32375 7185 32385 7220
rect 32420 7185 32430 7220
rect 32465 7185 32475 7220
rect 32510 7185 32520 7220
rect 32555 7185 32565 7220
rect 32600 7185 32610 7220
rect 32645 7185 32655 7220
rect 32690 7185 32700 7220
rect 32735 7185 32745 7220
rect 32780 7185 32790 7220
rect 32825 7185 32835 7220
rect 32870 7185 35620 7220
rect 31290 7175 35620 7185
rect 31290 7140 31305 7175
rect 31340 7140 31350 7175
rect 31385 7140 31395 7175
rect 31430 7140 31440 7175
rect 31475 7140 31485 7175
rect 31520 7140 31530 7175
rect 31565 7140 31575 7175
rect 31610 7140 31620 7175
rect 31655 7140 31665 7175
rect 31700 7140 31710 7175
rect 31745 7140 31755 7175
rect 31790 7140 31800 7175
rect 31835 7140 31845 7175
rect 31880 7140 31890 7175
rect 31925 7140 31935 7175
rect 31970 7140 31980 7175
rect 32015 7140 32025 7175
rect 32060 7140 32070 7175
rect 32105 7140 32115 7175
rect 32150 7140 32160 7175
rect 32195 7140 32205 7175
rect 32240 7140 32250 7175
rect 32285 7140 32295 7175
rect 32330 7140 32340 7175
rect 32375 7140 32385 7175
rect 32420 7140 32430 7175
rect 32465 7140 32475 7175
rect 32510 7140 32520 7175
rect 32555 7140 32565 7175
rect 32600 7140 32610 7175
rect 32645 7140 32655 7175
rect 32690 7140 32700 7175
rect 32735 7140 32745 7175
rect 32780 7140 32790 7175
rect 32825 7140 32835 7175
rect 32870 7140 35620 7175
rect 31290 7130 35620 7140
rect 31290 7095 31305 7130
rect 31340 7095 31350 7130
rect 31385 7095 31395 7130
rect 31430 7095 31440 7130
rect 31475 7095 31485 7130
rect 31520 7095 31530 7130
rect 31565 7095 31575 7130
rect 31610 7095 31620 7130
rect 31655 7095 31665 7130
rect 31700 7095 31710 7130
rect 31745 7095 31755 7130
rect 31790 7095 31800 7130
rect 31835 7095 31845 7130
rect 31880 7095 31890 7130
rect 31925 7095 31935 7130
rect 31970 7095 31980 7130
rect 32015 7095 32025 7130
rect 32060 7095 32070 7130
rect 32105 7095 32115 7130
rect 32150 7095 32160 7130
rect 32195 7095 32205 7130
rect 32240 7095 32250 7130
rect 32285 7095 32295 7130
rect 32330 7095 32340 7130
rect 32375 7095 32385 7130
rect 32420 7095 32430 7130
rect 32465 7095 32475 7130
rect 32510 7095 32520 7130
rect 32555 7095 32565 7130
rect 32600 7095 32610 7130
rect 32645 7095 32655 7130
rect 32690 7095 32700 7130
rect 32735 7095 32745 7130
rect 32780 7095 32790 7130
rect 32825 7095 32835 7130
rect 32870 7095 35620 7130
rect 31290 7085 35620 7095
rect 31290 7050 31305 7085
rect 31340 7050 31350 7085
rect 31385 7050 31395 7085
rect 31430 7050 31440 7085
rect 31475 7050 31485 7085
rect 31520 7050 31530 7085
rect 31565 7050 31575 7085
rect 31610 7050 31620 7085
rect 31655 7050 31665 7085
rect 31700 7050 31710 7085
rect 31745 7050 31755 7085
rect 31790 7050 31800 7085
rect 31835 7050 31845 7085
rect 31880 7050 31890 7085
rect 31925 7050 31935 7085
rect 31970 7050 31980 7085
rect 32015 7050 32025 7085
rect 32060 7050 32070 7085
rect 32105 7050 32115 7085
rect 32150 7050 32160 7085
rect 32195 7050 32205 7085
rect 32240 7050 32250 7085
rect 32285 7050 32295 7085
rect 32330 7050 32340 7085
rect 32375 7050 32385 7085
rect 32420 7050 32430 7085
rect 32465 7050 32475 7085
rect 32510 7050 32520 7085
rect 32555 7050 32565 7085
rect 32600 7050 32610 7085
rect 32645 7050 32655 7085
rect 32690 7050 32700 7085
rect 32735 7050 32745 7085
rect 32780 7050 32790 7085
rect 32825 7050 32835 7085
rect 32870 7050 35620 7085
rect 31290 7040 35620 7050
rect 31290 7005 31305 7040
rect 31340 7005 31350 7040
rect 31385 7005 31395 7040
rect 31430 7005 31440 7040
rect 31475 7005 31485 7040
rect 31520 7005 31530 7040
rect 31565 7005 31575 7040
rect 31610 7005 31620 7040
rect 31655 7005 31665 7040
rect 31700 7005 31710 7040
rect 31745 7005 31755 7040
rect 31790 7005 31800 7040
rect 31835 7005 31845 7040
rect 31880 7005 31890 7040
rect 31925 7005 31935 7040
rect 31970 7005 31980 7040
rect 32015 7005 32025 7040
rect 32060 7005 32070 7040
rect 32105 7005 32115 7040
rect 32150 7005 32160 7040
rect 32195 7005 32205 7040
rect 32240 7005 32250 7040
rect 32285 7005 32295 7040
rect 32330 7005 32340 7040
rect 32375 7005 32385 7040
rect 32420 7005 32430 7040
rect 32465 7005 32475 7040
rect 32510 7005 32520 7040
rect 32555 7005 32565 7040
rect 32600 7005 32610 7040
rect 32645 7005 32655 7040
rect 32690 7005 32700 7040
rect 32735 7005 32745 7040
rect 32780 7005 32790 7040
rect 32825 7005 32835 7040
rect 32870 7005 35620 7040
rect 31290 6995 35620 7005
rect 31290 6960 31305 6995
rect 31340 6960 31350 6995
rect 31385 6960 31395 6995
rect 31430 6960 31440 6995
rect 31475 6960 31485 6995
rect 31520 6960 31530 6995
rect 31565 6960 31575 6995
rect 31610 6960 31620 6995
rect 31655 6960 31665 6995
rect 31700 6960 31710 6995
rect 31745 6960 31755 6995
rect 31790 6960 31800 6995
rect 31835 6960 31845 6995
rect 31880 6960 31890 6995
rect 31925 6960 31935 6995
rect 31970 6960 31980 6995
rect 32015 6960 32025 6995
rect 32060 6960 32070 6995
rect 32105 6960 32115 6995
rect 32150 6960 32160 6995
rect 32195 6960 32205 6995
rect 32240 6960 32250 6995
rect 32285 6960 32295 6995
rect 32330 6960 32340 6995
rect 32375 6960 32385 6995
rect 32420 6960 32430 6995
rect 32465 6960 32475 6995
rect 32510 6960 32520 6995
rect 32555 6960 32565 6995
rect 32600 6960 32610 6995
rect 32645 6960 32655 6995
rect 32690 6960 32700 6995
rect 32735 6960 32745 6995
rect 32780 6960 32790 6995
rect 32825 6960 32835 6995
rect 32870 6960 35620 6995
rect 31290 6950 35620 6960
rect 31290 6915 31305 6950
rect 31340 6915 31350 6950
rect 31385 6915 31395 6950
rect 31430 6915 31440 6950
rect 31475 6915 31485 6950
rect 31520 6915 31530 6950
rect 31565 6915 31575 6950
rect 31610 6915 31620 6950
rect 31655 6915 31665 6950
rect 31700 6915 31710 6950
rect 31745 6915 31755 6950
rect 31790 6915 31800 6950
rect 31835 6915 31845 6950
rect 31880 6915 31890 6950
rect 31925 6915 31935 6950
rect 31970 6915 31980 6950
rect 32015 6915 32025 6950
rect 32060 6915 32070 6950
rect 32105 6915 32115 6950
rect 32150 6915 32160 6950
rect 32195 6915 32205 6950
rect 32240 6915 32250 6950
rect 32285 6915 32295 6950
rect 32330 6915 32340 6950
rect 32375 6915 32385 6950
rect 32420 6915 32430 6950
rect 32465 6915 32475 6950
rect 32510 6915 32520 6950
rect 32555 6915 32565 6950
rect 32600 6915 32610 6950
rect 32645 6915 32655 6950
rect 32690 6915 32700 6950
rect 32735 6915 32745 6950
rect 32780 6915 32790 6950
rect 32825 6915 32835 6950
rect 32870 6915 35620 6950
rect 31290 6905 35620 6915
rect 31290 6870 31305 6905
rect 31340 6870 31350 6905
rect 31385 6870 31395 6905
rect 31430 6870 31440 6905
rect 31475 6870 31485 6905
rect 31520 6870 31530 6905
rect 31565 6870 31575 6905
rect 31610 6870 31620 6905
rect 31655 6870 31665 6905
rect 31700 6870 31710 6905
rect 31745 6870 31755 6905
rect 31790 6870 31800 6905
rect 31835 6870 31845 6905
rect 31880 6870 31890 6905
rect 31925 6870 31935 6905
rect 31970 6870 31980 6905
rect 32015 6870 32025 6905
rect 32060 6870 32070 6905
rect 32105 6870 32115 6905
rect 32150 6870 32160 6905
rect 32195 6870 32205 6905
rect 32240 6870 32250 6905
rect 32285 6870 32295 6905
rect 32330 6870 32340 6905
rect 32375 6870 32385 6905
rect 32420 6870 32430 6905
rect 32465 6870 32475 6905
rect 32510 6870 32520 6905
rect 32555 6870 32565 6905
rect 32600 6870 32610 6905
rect 32645 6870 32655 6905
rect 32690 6870 32700 6905
rect 32735 6870 32745 6905
rect 32780 6870 32790 6905
rect 32825 6870 32835 6905
rect 32870 6870 35620 6905
rect 31290 6860 35620 6870
rect 31290 6825 31305 6860
rect 31340 6825 31350 6860
rect 31385 6825 31395 6860
rect 31430 6825 31440 6860
rect 31475 6825 31485 6860
rect 31520 6825 31530 6860
rect 31565 6825 31575 6860
rect 31610 6825 31620 6860
rect 31655 6825 31665 6860
rect 31700 6825 31710 6860
rect 31745 6825 31755 6860
rect 31790 6825 31800 6860
rect 31835 6825 31845 6860
rect 31880 6825 31890 6860
rect 31925 6825 31935 6860
rect 31970 6825 31980 6860
rect 32015 6825 32025 6860
rect 32060 6825 32070 6860
rect 32105 6825 32115 6860
rect 32150 6825 32160 6860
rect 32195 6825 32205 6860
rect 32240 6825 32250 6860
rect 32285 6825 32295 6860
rect 32330 6825 32340 6860
rect 32375 6825 32385 6860
rect 32420 6825 32430 6860
rect 32465 6825 32475 6860
rect 32510 6825 32520 6860
rect 32555 6825 32565 6860
rect 32600 6825 32610 6860
rect 32645 6825 32655 6860
rect 32690 6825 32700 6860
rect 32735 6825 32745 6860
rect 32780 6825 32790 6860
rect 32825 6825 32835 6860
rect 32870 6825 35620 6860
rect 31290 6815 35620 6825
rect 31290 6780 31305 6815
rect 31340 6780 31350 6815
rect 31385 6780 31395 6815
rect 31430 6780 31440 6815
rect 31475 6780 31485 6815
rect 31520 6780 31530 6815
rect 31565 6780 31575 6815
rect 31610 6780 31620 6815
rect 31655 6780 31665 6815
rect 31700 6780 31710 6815
rect 31745 6780 31755 6815
rect 31790 6780 31800 6815
rect 31835 6780 31845 6815
rect 31880 6780 31890 6815
rect 31925 6780 31935 6815
rect 31970 6780 31980 6815
rect 32015 6780 32025 6815
rect 32060 6780 32070 6815
rect 32105 6780 32115 6815
rect 32150 6780 32160 6815
rect 32195 6780 32205 6815
rect 32240 6780 32250 6815
rect 32285 6780 32295 6815
rect 32330 6780 32340 6815
rect 32375 6780 32385 6815
rect 32420 6780 32430 6815
rect 32465 6780 32475 6815
rect 32510 6780 32520 6815
rect 32555 6780 32565 6815
rect 32600 6780 32610 6815
rect 32645 6780 32655 6815
rect 32690 6780 32700 6815
rect 32735 6780 32745 6815
rect 32780 6780 32790 6815
rect 32825 6780 32835 6815
rect 32870 6780 35620 6815
rect 31290 6770 35620 6780
rect 31290 6735 31305 6770
rect 31340 6735 31350 6770
rect 31385 6735 31395 6770
rect 31430 6735 31440 6770
rect 31475 6735 31485 6770
rect 31520 6735 31530 6770
rect 31565 6735 31575 6770
rect 31610 6735 31620 6770
rect 31655 6735 31665 6770
rect 31700 6735 31710 6770
rect 31745 6735 31755 6770
rect 31790 6735 31800 6770
rect 31835 6735 31845 6770
rect 31880 6735 31890 6770
rect 31925 6735 31935 6770
rect 31970 6735 31980 6770
rect 32015 6735 32025 6770
rect 32060 6735 32070 6770
rect 32105 6735 32115 6770
rect 32150 6735 32160 6770
rect 32195 6735 32205 6770
rect 32240 6735 32250 6770
rect 32285 6735 32295 6770
rect 32330 6735 32340 6770
rect 32375 6735 32385 6770
rect 32420 6735 32430 6770
rect 32465 6735 32475 6770
rect 32510 6735 32520 6770
rect 32555 6735 32565 6770
rect 32600 6735 32610 6770
rect 32645 6735 32655 6770
rect 32690 6735 32700 6770
rect 32735 6735 32745 6770
rect 32780 6735 32790 6770
rect 32825 6735 32835 6770
rect 32870 6735 35620 6770
rect 31290 6725 35620 6735
rect 31290 6690 31305 6725
rect 31340 6690 31350 6725
rect 31385 6690 31395 6725
rect 31430 6690 31440 6725
rect 31475 6690 31485 6725
rect 31520 6690 31530 6725
rect 31565 6690 31575 6725
rect 31610 6690 31620 6725
rect 31655 6690 31665 6725
rect 31700 6690 31710 6725
rect 31745 6690 31755 6725
rect 31790 6690 31800 6725
rect 31835 6690 31845 6725
rect 31880 6690 31890 6725
rect 31925 6690 31935 6725
rect 31970 6690 31980 6725
rect 32015 6690 32025 6725
rect 32060 6690 32070 6725
rect 32105 6690 32115 6725
rect 32150 6690 32160 6725
rect 32195 6690 32205 6725
rect 32240 6690 32250 6725
rect 32285 6690 32295 6725
rect 32330 6690 32340 6725
rect 32375 6690 32385 6725
rect 32420 6690 32430 6725
rect 32465 6690 32475 6725
rect 32510 6690 32520 6725
rect 32555 6690 32565 6725
rect 32600 6690 32610 6725
rect 32645 6690 32655 6725
rect 32690 6690 32700 6725
rect 32735 6690 32745 6725
rect 32780 6690 32790 6725
rect 32825 6690 32835 6725
rect 32870 6690 35620 6725
rect 31290 6680 35620 6690
rect 31290 6645 31305 6680
rect 31340 6645 31350 6680
rect 31385 6645 31395 6680
rect 31430 6645 31440 6680
rect 31475 6645 31485 6680
rect 31520 6645 31530 6680
rect 31565 6645 31575 6680
rect 31610 6645 31620 6680
rect 31655 6645 31665 6680
rect 31700 6645 31710 6680
rect 31745 6645 31755 6680
rect 31790 6645 31800 6680
rect 31835 6645 31845 6680
rect 31880 6645 31890 6680
rect 31925 6645 31935 6680
rect 31970 6645 31980 6680
rect 32015 6645 32025 6680
rect 32060 6645 32070 6680
rect 32105 6645 32115 6680
rect 32150 6645 32160 6680
rect 32195 6645 32205 6680
rect 32240 6645 32250 6680
rect 32285 6645 32295 6680
rect 32330 6645 32340 6680
rect 32375 6645 32385 6680
rect 32420 6645 32430 6680
rect 32465 6645 32475 6680
rect 32510 6645 32520 6680
rect 32555 6645 32565 6680
rect 32600 6645 32610 6680
rect 32645 6645 32655 6680
rect 32690 6645 32700 6680
rect 32735 6645 32745 6680
rect 32780 6645 32790 6680
rect 32825 6645 32835 6680
rect 32870 6645 35620 6680
rect 31290 6635 35620 6645
rect 31290 6600 31305 6635
rect 31340 6600 31350 6635
rect 31385 6600 31395 6635
rect 31430 6600 31440 6635
rect 31475 6600 31485 6635
rect 31520 6600 31530 6635
rect 31565 6600 31575 6635
rect 31610 6600 31620 6635
rect 31655 6600 31665 6635
rect 31700 6600 31710 6635
rect 31745 6600 31755 6635
rect 31790 6600 31800 6635
rect 31835 6600 31845 6635
rect 31880 6600 31890 6635
rect 31925 6600 31935 6635
rect 31970 6600 31980 6635
rect 32015 6600 32025 6635
rect 32060 6600 32070 6635
rect 32105 6600 32115 6635
rect 32150 6600 32160 6635
rect 32195 6600 32205 6635
rect 32240 6600 32250 6635
rect 32285 6600 32295 6635
rect 32330 6600 32340 6635
rect 32375 6600 32385 6635
rect 32420 6600 32430 6635
rect 32465 6600 32475 6635
rect 32510 6600 32520 6635
rect 32555 6600 32565 6635
rect 32600 6600 32610 6635
rect 32645 6600 32655 6635
rect 32690 6600 32700 6635
rect 32735 6600 32745 6635
rect 32780 6600 32790 6635
rect 32825 6600 32835 6635
rect 32870 6600 35620 6635
rect 31290 6590 35620 6600
rect 31290 6555 31305 6590
rect 31340 6555 31350 6590
rect 31385 6555 31395 6590
rect 31430 6555 31440 6590
rect 31475 6555 31485 6590
rect 31520 6555 31530 6590
rect 31565 6555 31575 6590
rect 31610 6555 31620 6590
rect 31655 6555 31665 6590
rect 31700 6555 31710 6590
rect 31745 6555 31755 6590
rect 31790 6555 31800 6590
rect 31835 6555 31845 6590
rect 31880 6555 31890 6590
rect 31925 6555 31935 6590
rect 31970 6555 31980 6590
rect 32015 6555 32025 6590
rect 32060 6555 32070 6590
rect 32105 6555 32115 6590
rect 32150 6555 32160 6590
rect 32195 6555 32205 6590
rect 32240 6555 32250 6590
rect 32285 6555 32295 6590
rect 32330 6555 32340 6590
rect 32375 6555 32385 6590
rect 32420 6555 32430 6590
rect 32465 6555 32475 6590
rect 32510 6555 32520 6590
rect 32555 6555 32565 6590
rect 32600 6555 32610 6590
rect 32645 6555 32655 6590
rect 32690 6555 32700 6590
rect 32735 6555 32745 6590
rect 32780 6555 32790 6590
rect 32825 6555 32835 6590
rect 32870 6555 35620 6590
rect 31290 6545 35620 6555
rect 31290 6510 31305 6545
rect 31340 6510 31350 6545
rect 31385 6510 31395 6545
rect 31430 6510 31440 6545
rect 31475 6510 31485 6545
rect 31520 6510 31530 6545
rect 31565 6510 31575 6545
rect 31610 6510 31620 6545
rect 31655 6510 31665 6545
rect 31700 6510 31710 6545
rect 31745 6510 31755 6545
rect 31790 6510 31800 6545
rect 31835 6510 31845 6545
rect 31880 6510 31890 6545
rect 31925 6510 31935 6545
rect 31970 6510 31980 6545
rect 32015 6510 32025 6545
rect 32060 6510 32070 6545
rect 32105 6510 32115 6545
rect 32150 6510 32160 6545
rect 32195 6510 32205 6545
rect 32240 6510 32250 6545
rect 32285 6510 32295 6545
rect 32330 6510 32340 6545
rect 32375 6510 32385 6545
rect 32420 6510 32430 6545
rect 32465 6510 32475 6545
rect 32510 6510 32520 6545
rect 32555 6510 32565 6545
rect 32600 6510 32610 6545
rect 32645 6510 32655 6545
rect 32690 6510 32700 6545
rect 32735 6510 32745 6545
rect 32780 6510 32790 6545
rect 32825 6510 32835 6545
rect 32870 6510 35620 6545
rect 31290 6500 35620 6510
rect 31290 6465 31305 6500
rect 31340 6465 31350 6500
rect 31385 6465 31395 6500
rect 31430 6465 31440 6500
rect 31475 6465 31485 6500
rect 31520 6465 31530 6500
rect 31565 6465 31575 6500
rect 31610 6465 31620 6500
rect 31655 6465 31665 6500
rect 31700 6465 31710 6500
rect 31745 6465 31755 6500
rect 31790 6465 31800 6500
rect 31835 6465 31845 6500
rect 31880 6465 31890 6500
rect 31925 6465 31935 6500
rect 31970 6465 31980 6500
rect 32015 6465 32025 6500
rect 32060 6465 32070 6500
rect 32105 6465 32115 6500
rect 32150 6465 32160 6500
rect 32195 6465 32205 6500
rect 32240 6465 32250 6500
rect 32285 6465 32295 6500
rect 32330 6465 32340 6500
rect 32375 6465 32385 6500
rect 32420 6465 32430 6500
rect 32465 6465 32475 6500
rect 32510 6465 32520 6500
rect 32555 6465 32565 6500
rect 32600 6465 32610 6500
rect 32645 6465 32655 6500
rect 32690 6465 32700 6500
rect 32735 6465 32745 6500
rect 32780 6465 32790 6500
rect 32825 6465 32835 6500
rect 32870 6465 35620 6500
rect 31290 6450 35620 6465
rect -38770 6435 3390 6445
rect -120 -1315 32890 -1305
rect -120 -1355 -80 -1315
rect -40 -1355 270 -1315
rect 310 -1355 620 -1315
rect 660 -1355 970 -1315
rect 1010 -1355 1320 -1315
rect 1360 -1355 1670 -1315
rect 1710 -1355 2020 -1315
rect 2060 -1355 2370 -1315
rect 2410 -1355 2720 -1315
rect 2760 -1355 3070 -1315
rect 3110 -1355 5870 -1315
rect 5910 -1355 6220 -1315
rect 6260 -1355 6570 -1315
rect 6610 -1355 6920 -1315
rect 6960 -1355 7270 -1315
rect 7310 -1355 7620 -1315
rect 7660 -1355 7970 -1315
rect 8010 -1355 8320 -1315
rect 8360 -1355 8670 -1315
rect 8710 -1355 9020 -1315
rect 9060 -1325 32890 -1315
rect 9060 -1355 31305 -1325
rect -120 -1360 31305 -1355
rect 31340 -1360 31350 -1325
rect 31385 -1360 31395 -1325
rect 31430 -1360 31440 -1325
rect 31475 -1360 31485 -1325
rect 31520 -1360 31530 -1325
rect 31565 -1360 31575 -1325
rect 31610 -1360 31620 -1325
rect 31655 -1360 31665 -1325
rect 31700 -1360 31710 -1325
rect 31745 -1360 31755 -1325
rect 31790 -1360 31800 -1325
rect 31835 -1360 31845 -1325
rect 31880 -1360 31890 -1325
rect 31925 -1360 31935 -1325
rect 31970 -1360 31980 -1325
rect 32015 -1360 32025 -1325
rect 32060 -1360 32070 -1325
rect 32105 -1360 32115 -1325
rect 32150 -1360 32160 -1325
rect 32195 -1360 32205 -1325
rect 32240 -1360 32250 -1325
rect 32285 -1360 32295 -1325
rect 32330 -1360 32340 -1325
rect 32375 -1360 32385 -1325
rect 32420 -1360 32430 -1325
rect 32465 -1360 32475 -1325
rect 32510 -1360 32520 -1325
rect 32555 -1360 32565 -1325
rect 32600 -1360 32610 -1325
rect 32645 -1360 32655 -1325
rect 32690 -1360 32700 -1325
rect 32735 -1360 32745 -1325
rect 32780 -1360 32790 -1325
rect 32825 -1360 32835 -1325
rect 32870 -1360 32890 -1325
rect -120 -1370 32890 -1360
rect -120 -1380 31305 -1370
rect -120 -1420 -80 -1380
rect -40 -1420 270 -1380
rect 310 -1420 620 -1380
rect 660 -1420 970 -1380
rect 1010 -1420 1320 -1380
rect 1360 -1420 1670 -1380
rect 1710 -1420 2020 -1380
rect 2060 -1420 2370 -1380
rect 2410 -1420 2720 -1380
rect 2760 -1420 3070 -1380
rect 3110 -1420 5870 -1380
rect 5910 -1420 6220 -1380
rect 6260 -1420 6570 -1380
rect 6610 -1420 6920 -1380
rect 6960 -1420 7270 -1380
rect 7310 -1420 7620 -1380
rect 7660 -1420 7970 -1380
rect 8010 -1420 8320 -1380
rect 8360 -1420 8670 -1380
rect 8710 -1420 9020 -1380
rect 9060 -1405 31305 -1380
rect 31340 -1405 31350 -1370
rect 31385 -1405 31395 -1370
rect 31430 -1405 31440 -1370
rect 31475 -1405 31485 -1370
rect 31520 -1405 31530 -1370
rect 31565 -1405 31575 -1370
rect 31610 -1405 31620 -1370
rect 31655 -1405 31665 -1370
rect 31700 -1405 31710 -1370
rect 31745 -1405 31755 -1370
rect 31790 -1405 31800 -1370
rect 31835 -1405 31845 -1370
rect 31880 -1405 31890 -1370
rect 31925 -1405 31935 -1370
rect 31970 -1405 31980 -1370
rect 32015 -1405 32025 -1370
rect 32060 -1405 32070 -1370
rect 32105 -1405 32115 -1370
rect 32150 -1405 32160 -1370
rect 32195 -1405 32205 -1370
rect 32240 -1405 32250 -1370
rect 32285 -1405 32295 -1370
rect 32330 -1405 32340 -1370
rect 32375 -1405 32385 -1370
rect 32420 -1405 32430 -1370
rect 32465 -1405 32475 -1370
rect 32510 -1405 32520 -1370
rect 32555 -1405 32565 -1370
rect 32600 -1405 32610 -1370
rect 32645 -1405 32655 -1370
rect 32690 -1405 32700 -1370
rect 32735 -1405 32745 -1370
rect 32780 -1405 32790 -1370
rect 32825 -1405 32835 -1370
rect 32870 -1405 32890 -1370
rect 9060 -1415 32890 -1405
rect 9060 -1420 31305 -1415
rect -120 -1450 31305 -1420
rect 31340 -1450 31350 -1415
rect 31385 -1450 31395 -1415
rect 31430 -1450 31440 -1415
rect 31475 -1450 31485 -1415
rect 31520 -1450 31530 -1415
rect 31565 -1450 31575 -1415
rect 31610 -1450 31620 -1415
rect 31655 -1450 31665 -1415
rect 31700 -1450 31710 -1415
rect 31745 -1450 31755 -1415
rect 31790 -1450 31800 -1415
rect 31835 -1450 31845 -1415
rect 31880 -1450 31890 -1415
rect 31925 -1450 31935 -1415
rect 31970 -1450 31980 -1415
rect 32015 -1450 32025 -1415
rect 32060 -1450 32070 -1415
rect 32105 -1450 32115 -1415
rect 32150 -1450 32160 -1415
rect 32195 -1450 32205 -1415
rect 32240 -1450 32250 -1415
rect 32285 -1450 32295 -1415
rect 32330 -1450 32340 -1415
rect 32375 -1450 32385 -1415
rect 32420 -1450 32430 -1415
rect 32465 -1450 32475 -1415
rect 32510 -1450 32520 -1415
rect 32555 -1450 32565 -1415
rect 32600 -1450 32610 -1415
rect 32645 -1450 32655 -1415
rect 32690 -1450 32700 -1415
rect 32735 -1450 32745 -1415
rect 32780 -1450 32790 -1415
rect 32825 -1450 32835 -1415
rect 32870 -1450 32890 -1415
rect -120 -1490 -80 -1450
rect -40 -1490 270 -1450
rect 310 -1490 620 -1450
rect 660 -1490 970 -1450
rect 1010 -1490 1320 -1450
rect 1360 -1490 1670 -1450
rect 1710 -1490 2020 -1450
rect 2060 -1490 2370 -1450
rect 2410 -1490 2720 -1450
rect 2760 -1490 3070 -1450
rect 3110 -1490 5870 -1450
rect 5910 -1490 6220 -1450
rect 6260 -1490 6570 -1450
rect 6610 -1490 6920 -1450
rect 6960 -1490 7270 -1450
rect 7310 -1490 7620 -1450
rect 7660 -1490 7970 -1450
rect 8010 -1490 8320 -1450
rect 8360 -1490 8670 -1450
rect 8710 -1490 9020 -1450
rect 9060 -1460 32890 -1450
rect 9060 -1490 31305 -1460
rect -120 -1495 31305 -1490
rect 31340 -1495 31350 -1460
rect 31385 -1495 31395 -1460
rect 31430 -1495 31440 -1460
rect 31475 -1495 31485 -1460
rect 31520 -1495 31530 -1460
rect 31565 -1495 31575 -1460
rect 31610 -1495 31620 -1460
rect 31655 -1495 31665 -1460
rect 31700 -1495 31710 -1460
rect 31745 -1495 31755 -1460
rect 31790 -1495 31800 -1460
rect 31835 -1495 31845 -1460
rect 31880 -1495 31890 -1460
rect 31925 -1495 31935 -1460
rect 31970 -1495 31980 -1460
rect 32015 -1495 32025 -1460
rect 32060 -1495 32070 -1460
rect 32105 -1495 32115 -1460
rect 32150 -1495 32160 -1460
rect 32195 -1495 32205 -1460
rect 32240 -1495 32250 -1460
rect 32285 -1495 32295 -1460
rect 32330 -1495 32340 -1460
rect 32375 -1495 32385 -1460
rect 32420 -1495 32430 -1460
rect 32465 -1495 32475 -1460
rect 32510 -1495 32520 -1460
rect 32555 -1495 32565 -1460
rect 32600 -1495 32610 -1460
rect 32645 -1495 32655 -1460
rect 32690 -1495 32700 -1460
rect 32735 -1495 32745 -1460
rect 32780 -1495 32790 -1460
rect 32825 -1495 32835 -1460
rect 32870 -1495 32890 -1460
rect -120 -1505 32890 -1495
rect -120 -1520 31305 -1505
rect -120 -1560 -80 -1520
rect -40 -1560 270 -1520
rect 310 -1560 620 -1520
rect 660 -1560 970 -1520
rect 1010 -1560 1320 -1520
rect 1360 -1560 1670 -1520
rect 1710 -1560 2020 -1520
rect 2060 -1560 2370 -1520
rect 2410 -1560 2720 -1520
rect 2760 -1560 3070 -1520
rect 3110 -1560 5870 -1520
rect 5910 -1560 6220 -1520
rect 6260 -1560 6570 -1520
rect 6610 -1560 6920 -1520
rect 6960 -1560 7270 -1520
rect 7310 -1560 7620 -1520
rect 7660 -1560 7970 -1520
rect 8010 -1560 8320 -1520
rect 8360 -1560 8670 -1520
rect 8710 -1560 9020 -1520
rect 9060 -1540 31305 -1520
rect 31340 -1540 31350 -1505
rect 31385 -1540 31395 -1505
rect 31430 -1540 31440 -1505
rect 31475 -1540 31485 -1505
rect 31520 -1540 31530 -1505
rect 31565 -1540 31575 -1505
rect 31610 -1540 31620 -1505
rect 31655 -1540 31665 -1505
rect 31700 -1540 31710 -1505
rect 31745 -1540 31755 -1505
rect 31790 -1540 31800 -1505
rect 31835 -1540 31845 -1505
rect 31880 -1540 31890 -1505
rect 31925 -1540 31935 -1505
rect 31970 -1540 31980 -1505
rect 32015 -1540 32025 -1505
rect 32060 -1540 32070 -1505
rect 32105 -1540 32115 -1505
rect 32150 -1540 32160 -1505
rect 32195 -1540 32205 -1505
rect 32240 -1540 32250 -1505
rect 32285 -1540 32295 -1505
rect 32330 -1540 32340 -1505
rect 32375 -1540 32385 -1505
rect 32420 -1540 32430 -1505
rect 32465 -1540 32475 -1505
rect 32510 -1540 32520 -1505
rect 32555 -1540 32565 -1505
rect 32600 -1540 32610 -1505
rect 32645 -1540 32655 -1505
rect 32690 -1540 32700 -1505
rect 32735 -1540 32745 -1505
rect 32780 -1540 32790 -1505
rect 32825 -1540 32835 -1505
rect 32870 -1540 32890 -1505
rect 9060 -1550 32890 -1540
rect 9060 -1560 31305 -1550
rect -120 -1585 31305 -1560
rect 31340 -1585 31350 -1550
rect 31385 -1585 31395 -1550
rect 31430 -1585 31440 -1550
rect 31475 -1585 31485 -1550
rect 31520 -1585 31530 -1550
rect 31565 -1585 31575 -1550
rect 31610 -1585 31620 -1550
rect 31655 -1585 31665 -1550
rect 31700 -1585 31710 -1550
rect 31745 -1585 31755 -1550
rect 31790 -1585 31800 -1550
rect 31835 -1585 31845 -1550
rect 31880 -1585 31890 -1550
rect 31925 -1585 31935 -1550
rect 31970 -1585 31980 -1550
rect 32015 -1585 32025 -1550
rect 32060 -1585 32070 -1550
rect 32105 -1585 32115 -1550
rect 32150 -1585 32160 -1550
rect 32195 -1585 32205 -1550
rect 32240 -1585 32250 -1550
rect 32285 -1585 32295 -1550
rect 32330 -1585 32340 -1550
rect 32375 -1585 32385 -1550
rect 32420 -1585 32430 -1550
rect 32465 -1585 32475 -1550
rect 32510 -1585 32520 -1550
rect 32555 -1585 32565 -1550
rect 32600 -1585 32610 -1550
rect 32645 -1585 32655 -1550
rect 32690 -1585 32700 -1550
rect 32735 -1585 32745 -1550
rect 32780 -1585 32790 -1550
rect 32825 -1585 32835 -1550
rect 32870 -1585 32890 -1550
rect -120 -1590 32890 -1585
rect -120 -1630 -80 -1590
rect -40 -1630 270 -1590
rect 310 -1630 620 -1590
rect 660 -1630 970 -1590
rect 1010 -1630 1320 -1590
rect 1360 -1630 1670 -1590
rect 1710 -1630 2020 -1590
rect 2060 -1630 2370 -1590
rect 2410 -1630 2720 -1590
rect 2760 -1630 3070 -1590
rect 3110 -1630 5870 -1590
rect 5910 -1630 6220 -1590
rect 6260 -1630 6570 -1590
rect 6610 -1630 6920 -1590
rect 6960 -1630 7270 -1590
rect 7310 -1630 7620 -1590
rect 7660 -1630 7970 -1590
rect 8010 -1630 8320 -1590
rect 8360 -1630 8670 -1590
rect 8710 -1630 9020 -1590
rect 9060 -1595 32890 -1590
rect 9060 -1630 31305 -1595
rect 31340 -1630 31350 -1595
rect 31385 -1630 31395 -1595
rect 31430 -1630 31440 -1595
rect 31475 -1630 31485 -1595
rect 31520 -1630 31530 -1595
rect 31565 -1630 31575 -1595
rect 31610 -1630 31620 -1595
rect 31655 -1630 31665 -1595
rect 31700 -1630 31710 -1595
rect 31745 -1630 31755 -1595
rect 31790 -1630 31800 -1595
rect 31835 -1630 31845 -1595
rect 31880 -1630 31890 -1595
rect 31925 -1630 31935 -1595
rect 31970 -1630 31980 -1595
rect 32015 -1630 32025 -1595
rect 32060 -1630 32070 -1595
rect 32105 -1630 32115 -1595
rect 32150 -1630 32160 -1595
rect 32195 -1630 32205 -1595
rect 32240 -1630 32250 -1595
rect 32285 -1630 32295 -1595
rect 32330 -1630 32340 -1595
rect 32375 -1630 32385 -1595
rect 32420 -1630 32430 -1595
rect 32465 -1630 32475 -1595
rect 32510 -1630 32520 -1595
rect 32555 -1630 32565 -1595
rect 32600 -1630 32610 -1595
rect 32645 -1630 32655 -1595
rect 32690 -1630 32700 -1595
rect 32735 -1630 32745 -1595
rect 32780 -1630 32790 -1595
rect 32825 -1630 32835 -1595
rect 32870 -1630 32890 -1595
rect -120 -1640 32890 -1630
rect -120 -1655 31305 -1640
rect -120 -1695 -80 -1655
rect -40 -1695 270 -1655
rect 310 -1695 620 -1655
rect 660 -1695 970 -1655
rect 1010 -1695 1320 -1655
rect 1360 -1695 1670 -1655
rect 1710 -1695 2020 -1655
rect 2060 -1695 2370 -1655
rect 2410 -1695 2720 -1655
rect 2760 -1695 3070 -1655
rect 3110 -1695 5870 -1655
rect 5910 -1695 6220 -1655
rect 6260 -1695 6570 -1655
rect 6610 -1695 6920 -1655
rect 6960 -1695 7270 -1655
rect 7310 -1695 7620 -1655
rect 7660 -1695 7970 -1655
rect 8010 -1695 8320 -1655
rect 8360 -1695 8670 -1655
rect 8710 -1695 9020 -1655
rect 9060 -1675 31305 -1655
rect 31340 -1675 31350 -1640
rect 31385 -1675 31395 -1640
rect 31430 -1675 31440 -1640
rect 31475 -1675 31485 -1640
rect 31520 -1675 31530 -1640
rect 31565 -1675 31575 -1640
rect 31610 -1675 31620 -1640
rect 31655 -1675 31665 -1640
rect 31700 -1675 31710 -1640
rect 31745 -1675 31755 -1640
rect 31790 -1675 31800 -1640
rect 31835 -1675 31845 -1640
rect 31880 -1675 31890 -1640
rect 31925 -1675 31935 -1640
rect 31970 -1675 31980 -1640
rect 32015 -1675 32025 -1640
rect 32060 -1675 32070 -1640
rect 32105 -1675 32115 -1640
rect 32150 -1675 32160 -1640
rect 32195 -1675 32205 -1640
rect 32240 -1675 32250 -1640
rect 32285 -1675 32295 -1640
rect 32330 -1675 32340 -1640
rect 32375 -1675 32385 -1640
rect 32420 -1675 32430 -1640
rect 32465 -1675 32475 -1640
rect 32510 -1675 32520 -1640
rect 32555 -1675 32565 -1640
rect 32600 -1675 32610 -1640
rect 32645 -1675 32655 -1640
rect 32690 -1675 32700 -1640
rect 32735 -1675 32745 -1640
rect 32780 -1675 32790 -1640
rect 32825 -1675 32835 -1640
rect 32870 -1675 32890 -1640
rect 9060 -1685 32890 -1675
rect 9060 -1695 31305 -1685
rect -120 -1715 31305 -1695
rect -120 -1755 -80 -1715
rect -40 -1755 270 -1715
rect 310 -1755 620 -1715
rect 660 -1755 970 -1715
rect 1010 -1755 1320 -1715
rect 1360 -1755 1670 -1715
rect 1710 -1755 2020 -1715
rect 2060 -1755 2370 -1715
rect 2410 -1755 2720 -1715
rect 2760 -1755 3070 -1715
rect 3110 -1755 5870 -1715
rect 5910 -1755 6220 -1715
rect 6260 -1755 6570 -1715
rect 6610 -1755 6920 -1715
rect 6960 -1755 7270 -1715
rect 7310 -1755 7620 -1715
rect 7660 -1755 7970 -1715
rect 8010 -1755 8320 -1715
rect 8360 -1755 8670 -1715
rect 8710 -1755 9020 -1715
rect 9060 -1720 31305 -1715
rect 31340 -1720 31350 -1685
rect 31385 -1720 31395 -1685
rect 31430 -1720 31440 -1685
rect 31475 -1720 31485 -1685
rect 31520 -1720 31530 -1685
rect 31565 -1720 31575 -1685
rect 31610 -1720 31620 -1685
rect 31655 -1720 31665 -1685
rect 31700 -1720 31710 -1685
rect 31745 -1720 31755 -1685
rect 31790 -1720 31800 -1685
rect 31835 -1720 31845 -1685
rect 31880 -1720 31890 -1685
rect 31925 -1720 31935 -1685
rect 31970 -1720 31980 -1685
rect 32015 -1720 32025 -1685
rect 32060 -1720 32070 -1685
rect 32105 -1720 32115 -1685
rect 32150 -1720 32160 -1685
rect 32195 -1720 32205 -1685
rect 32240 -1720 32250 -1685
rect 32285 -1720 32295 -1685
rect 32330 -1720 32340 -1685
rect 32375 -1720 32385 -1685
rect 32420 -1720 32430 -1685
rect 32465 -1720 32475 -1685
rect 32510 -1720 32520 -1685
rect 32555 -1720 32565 -1685
rect 32600 -1720 32610 -1685
rect 32645 -1720 32655 -1685
rect 32690 -1720 32700 -1685
rect 32735 -1720 32745 -1685
rect 32780 -1720 32790 -1685
rect 32825 -1720 32835 -1685
rect 32870 -1720 32890 -1685
rect 9060 -1730 32890 -1720
rect 9060 -1755 31305 -1730
rect -120 -1765 31305 -1755
rect 31340 -1765 31350 -1730
rect 31385 -1765 31395 -1730
rect 31430 -1765 31440 -1730
rect 31475 -1765 31485 -1730
rect 31520 -1765 31530 -1730
rect 31565 -1765 31575 -1730
rect 31610 -1765 31620 -1730
rect 31655 -1765 31665 -1730
rect 31700 -1765 31710 -1730
rect 31745 -1765 31755 -1730
rect 31790 -1765 31800 -1730
rect 31835 -1765 31845 -1730
rect 31880 -1765 31890 -1730
rect 31925 -1765 31935 -1730
rect 31970 -1765 31980 -1730
rect 32015 -1765 32025 -1730
rect 32060 -1765 32070 -1730
rect 32105 -1765 32115 -1730
rect 32150 -1765 32160 -1730
rect 32195 -1765 32205 -1730
rect 32240 -1765 32250 -1730
rect 32285 -1765 32295 -1730
rect 32330 -1765 32340 -1730
rect 32375 -1765 32385 -1730
rect 32420 -1765 32430 -1730
rect 32465 -1765 32475 -1730
rect 32510 -1765 32520 -1730
rect 32555 -1765 32565 -1730
rect 32600 -1765 32610 -1730
rect 32645 -1765 32655 -1730
rect 32690 -1765 32700 -1730
rect 32735 -1765 32745 -1730
rect 32780 -1765 32790 -1730
rect 32825 -1765 32835 -1730
rect 32870 -1765 32890 -1730
rect -120 -1775 32890 -1765
rect -120 -1780 31305 -1775
rect -120 -1820 -80 -1780
rect -40 -1820 270 -1780
rect 310 -1820 620 -1780
rect 660 -1820 970 -1780
rect 1010 -1820 1320 -1780
rect 1360 -1820 1670 -1780
rect 1710 -1820 2020 -1780
rect 2060 -1820 2370 -1780
rect 2410 -1820 2720 -1780
rect 2760 -1820 3070 -1780
rect 3110 -1820 5870 -1780
rect 5910 -1820 6220 -1780
rect 6260 -1820 6570 -1780
rect 6610 -1820 6920 -1780
rect 6960 -1820 7270 -1780
rect 7310 -1820 7620 -1780
rect 7660 -1820 7970 -1780
rect 8010 -1820 8320 -1780
rect 8360 -1820 8670 -1780
rect 8710 -1820 9020 -1780
rect 9060 -1810 31305 -1780
rect 31340 -1810 31350 -1775
rect 31385 -1810 31395 -1775
rect 31430 -1810 31440 -1775
rect 31475 -1810 31485 -1775
rect 31520 -1810 31530 -1775
rect 31565 -1810 31575 -1775
rect 31610 -1810 31620 -1775
rect 31655 -1810 31665 -1775
rect 31700 -1810 31710 -1775
rect 31745 -1810 31755 -1775
rect 31790 -1810 31800 -1775
rect 31835 -1810 31845 -1775
rect 31880 -1810 31890 -1775
rect 31925 -1810 31935 -1775
rect 31970 -1810 31980 -1775
rect 32015 -1810 32025 -1775
rect 32060 -1810 32070 -1775
rect 32105 -1810 32115 -1775
rect 32150 -1810 32160 -1775
rect 32195 -1810 32205 -1775
rect 32240 -1810 32250 -1775
rect 32285 -1810 32295 -1775
rect 32330 -1810 32340 -1775
rect 32375 -1810 32385 -1775
rect 32420 -1810 32430 -1775
rect 32465 -1810 32475 -1775
rect 32510 -1810 32520 -1775
rect 32555 -1810 32565 -1775
rect 32600 -1810 32610 -1775
rect 32645 -1810 32655 -1775
rect 32690 -1810 32700 -1775
rect 32735 -1810 32745 -1775
rect 32780 -1810 32790 -1775
rect 32825 -1810 32835 -1775
rect 32870 -1810 32890 -1775
rect 9060 -1820 32890 -1810
rect -120 -1850 31305 -1820
rect -120 -1890 -80 -1850
rect -40 -1890 270 -1850
rect 310 -1890 620 -1850
rect 660 -1890 970 -1850
rect 1010 -1890 1320 -1850
rect 1360 -1890 1670 -1850
rect 1710 -1890 2020 -1850
rect 2060 -1890 2370 -1850
rect 2410 -1890 2720 -1850
rect 2760 -1890 3070 -1850
rect 3110 -1890 5870 -1850
rect 5910 -1890 6220 -1850
rect 6260 -1890 6570 -1850
rect 6610 -1890 6920 -1850
rect 6960 -1890 7270 -1850
rect 7310 -1890 7620 -1850
rect 7660 -1890 7970 -1850
rect 8010 -1890 8320 -1850
rect 8360 -1890 8670 -1850
rect 8710 -1890 9020 -1850
rect 9060 -1855 31305 -1850
rect 31340 -1855 31350 -1820
rect 31385 -1855 31395 -1820
rect 31430 -1855 31440 -1820
rect 31475 -1855 31485 -1820
rect 31520 -1855 31530 -1820
rect 31565 -1855 31575 -1820
rect 31610 -1855 31620 -1820
rect 31655 -1855 31665 -1820
rect 31700 -1855 31710 -1820
rect 31745 -1855 31755 -1820
rect 31790 -1855 31800 -1820
rect 31835 -1855 31845 -1820
rect 31880 -1855 31890 -1820
rect 31925 -1855 31935 -1820
rect 31970 -1855 31980 -1820
rect 32015 -1855 32025 -1820
rect 32060 -1855 32070 -1820
rect 32105 -1855 32115 -1820
rect 32150 -1855 32160 -1820
rect 32195 -1855 32205 -1820
rect 32240 -1855 32250 -1820
rect 32285 -1855 32295 -1820
rect 32330 -1855 32340 -1820
rect 32375 -1855 32385 -1820
rect 32420 -1855 32430 -1820
rect 32465 -1855 32475 -1820
rect 32510 -1855 32520 -1820
rect 32555 -1855 32565 -1820
rect 32600 -1855 32610 -1820
rect 32645 -1855 32655 -1820
rect 32690 -1855 32700 -1820
rect 32735 -1855 32745 -1820
rect 32780 -1855 32790 -1820
rect 32825 -1855 32835 -1820
rect 32870 -1855 32890 -1820
rect 9060 -1865 32890 -1855
rect 9060 -1890 31305 -1865
rect -120 -1900 31305 -1890
rect 31340 -1900 31350 -1865
rect 31385 -1900 31395 -1865
rect 31430 -1900 31440 -1865
rect 31475 -1900 31485 -1865
rect 31520 -1900 31530 -1865
rect 31565 -1900 31575 -1865
rect 31610 -1900 31620 -1865
rect 31655 -1900 31665 -1865
rect 31700 -1900 31710 -1865
rect 31745 -1900 31755 -1865
rect 31790 -1900 31800 -1865
rect 31835 -1900 31845 -1865
rect 31880 -1900 31890 -1865
rect 31925 -1900 31935 -1865
rect 31970 -1900 31980 -1865
rect 32015 -1900 32025 -1865
rect 32060 -1900 32070 -1865
rect 32105 -1900 32115 -1865
rect 32150 -1900 32160 -1865
rect 32195 -1900 32205 -1865
rect 32240 -1900 32250 -1865
rect 32285 -1900 32295 -1865
rect 32330 -1900 32340 -1865
rect 32375 -1900 32385 -1865
rect 32420 -1900 32430 -1865
rect 32465 -1900 32475 -1865
rect 32510 -1900 32520 -1865
rect 32555 -1900 32565 -1865
rect 32600 -1900 32610 -1865
rect 32645 -1900 32655 -1865
rect 32690 -1900 32700 -1865
rect 32735 -1900 32745 -1865
rect 32780 -1900 32790 -1865
rect 32825 -1900 32835 -1865
rect 32870 -1900 32890 -1865
rect -120 -1910 32890 -1900
rect -120 -1920 31305 -1910
rect -120 -1960 -80 -1920
rect -40 -1960 270 -1920
rect 310 -1960 620 -1920
rect 660 -1960 970 -1920
rect 1010 -1960 1320 -1920
rect 1360 -1960 1670 -1920
rect 1710 -1960 2020 -1920
rect 2060 -1960 2370 -1920
rect 2410 -1960 2720 -1920
rect 2760 -1960 3070 -1920
rect 3110 -1960 5870 -1920
rect 5910 -1960 6220 -1920
rect 6260 -1960 6570 -1920
rect 6610 -1960 6920 -1920
rect 6960 -1960 7270 -1920
rect 7310 -1960 7620 -1920
rect 7660 -1960 7970 -1920
rect 8010 -1960 8320 -1920
rect 8360 -1960 8670 -1920
rect 8710 -1960 9020 -1920
rect 9060 -1945 31305 -1920
rect 31340 -1945 31350 -1910
rect 31385 -1945 31395 -1910
rect 31430 -1945 31440 -1910
rect 31475 -1945 31485 -1910
rect 31520 -1945 31530 -1910
rect 31565 -1945 31575 -1910
rect 31610 -1945 31620 -1910
rect 31655 -1945 31665 -1910
rect 31700 -1945 31710 -1910
rect 31745 -1945 31755 -1910
rect 31790 -1945 31800 -1910
rect 31835 -1945 31845 -1910
rect 31880 -1945 31890 -1910
rect 31925 -1945 31935 -1910
rect 31970 -1945 31980 -1910
rect 32015 -1945 32025 -1910
rect 32060 -1945 32070 -1910
rect 32105 -1945 32115 -1910
rect 32150 -1945 32160 -1910
rect 32195 -1945 32205 -1910
rect 32240 -1945 32250 -1910
rect 32285 -1945 32295 -1910
rect 32330 -1945 32340 -1910
rect 32375 -1945 32385 -1910
rect 32420 -1945 32430 -1910
rect 32465 -1945 32475 -1910
rect 32510 -1945 32520 -1910
rect 32555 -1945 32565 -1910
rect 32600 -1945 32610 -1910
rect 32645 -1945 32655 -1910
rect 32690 -1945 32700 -1910
rect 32735 -1945 32745 -1910
rect 32780 -1945 32790 -1910
rect 32825 -1945 32835 -1910
rect 32870 -1945 32890 -1910
rect 9060 -1955 32890 -1945
rect 9060 -1960 31305 -1955
rect -120 -1990 31305 -1960
rect 31340 -1990 31350 -1955
rect 31385 -1990 31395 -1955
rect 31430 -1990 31440 -1955
rect 31475 -1990 31485 -1955
rect 31520 -1990 31530 -1955
rect 31565 -1990 31575 -1955
rect 31610 -1990 31620 -1955
rect 31655 -1990 31665 -1955
rect 31700 -1990 31710 -1955
rect 31745 -1990 31755 -1955
rect 31790 -1990 31800 -1955
rect 31835 -1990 31845 -1955
rect 31880 -1990 31890 -1955
rect 31925 -1990 31935 -1955
rect 31970 -1990 31980 -1955
rect 32015 -1990 32025 -1955
rect 32060 -1990 32070 -1955
rect 32105 -1990 32115 -1955
rect 32150 -1990 32160 -1955
rect 32195 -1990 32205 -1955
rect 32240 -1990 32250 -1955
rect 32285 -1990 32295 -1955
rect 32330 -1990 32340 -1955
rect 32375 -1990 32385 -1955
rect 32420 -1990 32430 -1955
rect 32465 -1990 32475 -1955
rect 32510 -1990 32520 -1955
rect 32555 -1990 32565 -1955
rect 32600 -1990 32610 -1955
rect 32645 -1990 32655 -1955
rect 32690 -1990 32700 -1955
rect 32735 -1990 32745 -1955
rect 32780 -1990 32790 -1955
rect 32825 -1990 32835 -1955
rect 32870 -1990 32890 -1955
rect -120 -2030 -80 -1990
rect -40 -2030 270 -1990
rect 310 -2030 620 -1990
rect 660 -2030 970 -1990
rect 1010 -2030 1320 -1990
rect 1360 -2030 1670 -1990
rect 1710 -2030 2020 -1990
rect 2060 -2030 2370 -1990
rect 2410 -2030 2720 -1990
rect 2760 -2030 3070 -1990
rect 3110 -2030 5870 -1990
rect 5910 -2030 6220 -1990
rect 6260 -2030 6570 -1990
rect 6610 -2030 6920 -1990
rect 6960 -2030 7270 -1990
rect 7310 -2030 7620 -1990
rect 7660 -2030 7970 -1990
rect 8010 -2030 8320 -1990
rect 8360 -2030 8670 -1990
rect 8710 -2030 9020 -1990
rect 9060 -2000 32890 -1990
rect 9060 -2030 31305 -2000
rect -120 -2035 31305 -2030
rect 31340 -2035 31350 -2000
rect 31385 -2035 31395 -2000
rect 31430 -2035 31440 -2000
rect 31475 -2035 31485 -2000
rect 31520 -2035 31530 -2000
rect 31565 -2035 31575 -2000
rect 31610 -2035 31620 -2000
rect 31655 -2035 31665 -2000
rect 31700 -2035 31710 -2000
rect 31745 -2035 31755 -2000
rect 31790 -2035 31800 -2000
rect 31835 -2035 31845 -2000
rect 31880 -2035 31890 -2000
rect 31925 -2035 31935 -2000
rect 31970 -2035 31980 -2000
rect 32015 -2035 32025 -2000
rect 32060 -2035 32070 -2000
rect 32105 -2035 32115 -2000
rect 32150 -2035 32160 -2000
rect 32195 -2035 32205 -2000
rect 32240 -2035 32250 -2000
rect 32285 -2035 32295 -2000
rect 32330 -2035 32340 -2000
rect 32375 -2035 32385 -2000
rect 32420 -2035 32430 -2000
rect 32465 -2035 32475 -2000
rect 32510 -2035 32520 -2000
rect 32555 -2035 32565 -2000
rect 32600 -2035 32610 -2000
rect 32645 -2035 32655 -2000
rect 32690 -2035 32700 -2000
rect 32735 -2035 32745 -2000
rect 32780 -2035 32790 -2000
rect 32825 -2035 32835 -2000
rect 32870 -2035 32890 -2000
rect -120 -2045 32890 -2035
rect -120 -2055 31305 -2045
rect -120 -2095 -80 -2055
rect -40 -2095 270 -2055
rect 310 -2095 620 -2055
rect 660 -2095 970 -2055
rect 1010 -2095 1320 -2055
rect 1360 -2095 1670 -2055
rect 1710 -2095 2020 -2055
rect 2060 -2095 2370 -2055
rect 2410 -2095 2720 -2055
rect 2760 -2095 3070 -2055
rect 3110 -2095 5870 -2055
rect 5910 -2095 6220 -2055
rect 6260 -2095 6570 -2055
rect 6610 -2095 6920 -2055
rect 6960 -2095 7270 -2055
rect 7310 -2095 7620 -2055
rect 7660 -2095 7970 -2055
rect 8010 -2095 8320 -2055
rect 8360 -2095 8670 -2055
rect 8710 -2095 9020 -2055
rect 9060 -2080 31305 -2055
rect 31340 -2080 31350 -2045
rect 31385 -2080 31395 -2045
rect 31430 -2080 31440 -2045
rect 31475 -2080 31485 -2045
rect 31520 -2080 31530 -2045
rect 31565 -2080 31575 -2045
rect 31610 -2080 31620 -2045
rect 31655 -2080 31665 -2045
rect 31700 -2080 31710 -2045
rect 31745 -2080 31755 -2045
rect 31790 -2080 31800 -2045
rect 31835 -2080 31845 -2045
rect 31880 -2080 31890 -2045
rect 31925 -2080 31935 -2045
rect 31970 -2080 31980 -2045
rect 32015 -2080 32025 -2045
rect 32060 -2080 32070 -2045
rect 32105 -2080 32115 -2045
rect 32150 -2080 32160 -2045
rect 32195 -2080 32205 -2045
rect 32240 -2080 32250 -2045
rect 32285 -2080 32295 -2045
rect 32330 -2080 32340 -2045
rect 32375 -2080 32385 -2045
rect 32420 -2080 32430 -2045
rect 32465 -2080 32475 -2045
rect 32510 -2080 32520 -2045
rect 32555 -2080 32565 -2045
rect 32600 -2080 32610 -2045
rect 32645 -2080 32655 -2045
rect 32690 -2080 32700 -2045
rect 32735 -2080 32745 -2045
rect 32780 -2080 32790 -2045
rect 32825 -2080 32835 -2045
rect 32870 -2080 32890 -2045
rect 9060 -2090 32890 -2080
rect 9060 -2095 31305 -2090
rect -120 -2115 31305 -2095
rect -120 -2155 -80 -2115
rect -40 -2155 270 -2115
rect 310 -2155 620 -2115
rect 660 -2155 970 -2115
rect 1010 -2155 1320 -2115
rect 1360 -2155 1670 -2115
rect 1710 -2155 2020 -2115
rect 2060 -2155 2370 -2115
rect 2410 -2155 2720 -2115
rect 2760 -2155 3070 -2115
rect 3110 -2155 5870 -2115
rect 5910 -2155 6220 -2115
rect 6260 -2155 6570 -2115
rect 6610 -2155 6920 -2115
rect 6960 -2155 7270 -2115
rect 7310 -2155 7620 -2115
rect 7660 -2155 7970 -2115
rect 8010 -2155 8320 -2115
rect 8360 -2155 8670 -2115
rect 8710 -2155 9020 -2115
rect 9060 -2125 31305 -2115
rect 31340 -2125 31350 -2090
rect 31385 -2125 31395 -2090
rect 31430 -2125 31440 -2090
rect 31475 -2125 31485 -2090
rect 31520 -2125 31530 -2090
rect 31565 -2125 31575 -2090
rect 31610 -2125 31620 -2090
rect 31655 -2125 31665 -2090
rect 31700 -2125 31710 -2090
rect 31745 -2125 31755 -2090
rect 31790 -2125 31800 -2090
rect 31835 -2125 31845 -2090
rect 31880 -2125 31890 -2090
rect 31925 -2125 31935 -2090
rect 31970 -2125 31980 -2090
rect 32015 -2125 32025 -2090
rect 32060 -2125 32070 -2090
rect 32105 -2125 32115 -2090
rect 32150 -2125 32160 -2090
rect 32195 -2125 32205 -2090
rect 32240 -2125 32250 -2090
rect 32285 -2125 32295 -2090
rect 32330 -2125 32340 -2090
rect 32375 -2125 32385 -2090
rect 32420 -2125 32430 -2090
rect 32465 -2125 32475 -2090
rect 32510 -2125 32520 -2090
rect 32555 -2125 32565 -2090
rect 32600 -2125 32610 -2090
rect 32645 -2125 32655 -2090
rect 32690 -2125 32700 -2090
rect 32735 -2125 32745 -2090
rect 32780 -2125 32790 -2090
rect 32825 -2125 32835 -2090
rect 32870 -2125 32890 -2090
rect 9060 -2135 32890 -2125
rect 9060 -2155 31305 -2135
rect -120 -2170 31305 -2155
rect 31340 -2170 31350 -2135
rect 31385 -2170 31395 -2135
rect 31430 -2170 31440 -2135
rect 31475 -2170 31485 -2135
rect 31520 -2170 31530 -2135
rect 31565 -2170 31575 -2135
rect 31610 -2170 31620 -2135
rect 31655 -2170 31665 -2135
rect 31700 -2170 31710 -2135
rect 31745 -2170 31755 -2135
rect 31790 -2170 31800 -2135
rect 31835 -2170 31845 -2135
rect 31880 -2170 31890 -2135
rect 31925 -2170 31935 -2135
rect 31970 -2170 31980 -2135
rect 32015 -2170 32025 -2135
rect 32060 -2170 32070 -2135
rect 32105 -2170 32115 -2135
rect 32150 -2170 32160 -2135
rect 32195 -2170 32205 -2135
rect 32240 -2170 32250 -2135
rect 32285 -2170 32295 -2135
rect 32330 -2170 32340 -2135
rect 32375 -2170 32385 -2135
rect 32420 -2170 32430 -2135
rect 32465 -2170 32475 -2135
rect 32510 -2170 32520 -2135
rect 32555 -2170 32565 -2135
rect 32600 -2170 32610 -2135
rect 32645 -2170 32655 -2135
rect 32690 -2170 32700 -2135
rect 32735 -2170 32745 -2135
rect 32780 -2170 32790 -2135
rect 32825 -2170 32835 -2135
rect 32870 -2170 32890 -2135
rect -120 -2180 32890 -2170
rect -120 -2220 -80 -2180
rect -40 -2220 270 -2180
rect 310 -2220 620 -2180
rect 660 -2220 970 -2180
rect 1010 -2220 1320 -2180
rect 1360 -2220 1670 -2180
rect 1710 -2220 2020 -2180
rect 2060 -2220 2370 -2180
rect 2410 -2220 2720 -2180
rect 2760 -2220 3070 -2180
rect 3110 -2220 5870 -2180
rect 5910 -2220 6220 -2180
rect 6260 -2220 6570 -2180
rect 6610 -2220 6920 -2180
rect 6960 -2220 7270 -2180
rect 7310 -2220 7620 -2180
rect 7660 -2220 7970 -2180
rect 8010 -2220 8320 -2180
rect 8360 -2220 8670 -2180
rect 8710 -2220 9020 -2180
rect 9060 -2215 31305 -2180
rect 31340 -2215 31350 -2180
rect 31385 -2215 31395 -2180
rect 31430 -2215 31440 -2180
rect 31475 -2215 31485 -2180
rect 31520 -2215 31530 -2180
rect 31565 -2215 31575 -2180
rect 31610 -2215 31620 -2180
rect 31655 -2215 31665 -2180
rect 31700 -2215 31710 -2180
rect 31745 -2215 31755 -2180
rect 31790 -2215 31800 -2180
rect 31835 -2215 31845 -2180
rect 31880 -2215 31890 -2180
rect 31925 -2215 31935 -2180
rect 31970 -2215 31980 -2180
rect 32015 -2215 32025 -2180
rect 32060 -2215 32070 -2180
rect 32105 -2215 32115 -2180
rect 32150 -2215 32160 -2180
rect 32195 -2215 32205 -2180
rect 32240 -2215 32250 -2180
rect 32285 -2215 32295 -2180
rect 32330 -2215 32340 -2180
rect 32375 -2215 32385 -2180
rect 32420 -2215 32430 -2180
rect 32465 -2215 32475 -2180
rect 32510 -2215 32520 -2180
rect 32555 -2215 32565 -2180
rect 32600 -2215 32610 -2180
rect 32645 -2215 32655 -2180
rect 32690 -2215 32700 -2180
rect 32735 -2215 32745 -2180
rect 32780 -2215 32790 -2180
rect 32825 -2215 32835 -2180
rect 32870 -2215 32890 -2180
rect 9060 -2220 32890 -2215
rect -120 -2225 32890 -2220
rect -120 -2250 31305 -2225
rect -120 -2290 -80 -2250
rect -40 -2290 270 -2250
rect 310 -2290 620 -2250
rect 660 -2290 970 -2250
rect 1010 -2290 1320 -2250
rect 1360 -2290 1670 -2250
rect 1710 -2290 2020 -2250
rect 2060 -2290 2370 -2250
rect 2410 -2290 2720 -2250
rect 2760 -2290 3070 -2250
rect 3110 -2290 5870 -2250
rect 5910 -2290 6220 -2250
rect 6260 -2290 6570 -2250
rect 6610 -2290 6920 -2250
rect 6960 -2290 7270 -2250
rect 7310 -2290 7620 -2250
rect 7660 -2290 7970 -2250
rect 8010 -2290 8320 -2250
rect 8360 -2290 8670 -2250
rect 8710 -2290 9020 -2250
rect 9060 -2260 31305 -2250
rect 31340 -2260 31350 -2225
rect 31385 -2260 31395 -2225
rect 31430 -2260 31440 -2225
rect 31475 -2260 31485 -2225
rect 31520 -2260 31530 -2225
rect 31565 -2260 31575 -2225
rect 31610 -2260 31620 -2225
rect 31655 -2260 31665 -2225
rect 31700 -2260 31710 -2225
rect 31745 -2260 31755 -2225
rect 31790 -2260 31800 -2225
rect 31835 -2260 31845 -2225
rect 31880 -2260 31890 -2225
rect 31925 -2260 31935 -2225
rect 31970 -2260 31980 -2225
rect 32015 -2260 32025 -2225
rect 32060 -2260 32070 -2225
rect 32105 -2260 32115 -2225
rect 32150 -2260 32160 -2225
rect 32195 -2260 32205 -2225
rect 32240 -2260 32250 -2225
rect 32285 -2260 32295 -2225
rect 32330 -2260 32340 -2225
rect 32375 -2260 32385 -2225
rect 32420 -2260 32430 -2225
rect 32465 -2260 32475 -2225
rect 32510 -2260 32520 -2225
rect 32555 -2260 32565 -2225
rect 32600 -2260 32610 -2225
rect 32645 -2260 32655 -2225
rect 32690 -2260 32700 -2225
rect 32735 -2260 32745 -2225
rect 32780 -2260 32790 -2225
rect 32825 -2260 32835 -2225
rect 32870 -2260 32890 -2225
rect 9060 -2270 32890 -2260
rect 9060 -2290 31305 -2270
rect -120 -2305 31305 -2290
rect 31340 -2305 31350 -2270
rect 31385 -2305 31395 -2270
rect 31430 -2305 31440 -2270
rect 31475 -2305 31485 -2270
rect 31520 -2305 31530 -2270
rect 31565 -2305 31575 -2270
rect 31610 -2305 31620 -2270
rect 31655 -2305 31665 -2270
rect 31700 -2305 31710 -2270
rect 31745 -2305 31755 -2270
rect 31790 -2305 31800 -2270
rect 31835 -2305 31845 -2270
rect 31880 -2305 31890 -2270
rect 31925 -2305 31935 -2270
rect 31970 -2305 31980 -2270
rect 32015 -2305 32025 -2270
rect 32060 -2305 32070 -2270
rect 32105 -2305 32115 -2270
rect 32150 -2305 32160 -2270
rect 32195 -2305 32205 -2270
rect 32240 -2305 32250 -2270
rect 32285 -2305 32295 -2270
rect 32330 -2305 32340 -2270
rect 32375 -2305 32385 -2270
rect 32420 -2305 32430 -2270
rect 32465 -2305 32475 -2270
rect 32510 -2305 32520 -2270
rect 32555 -2305 32565 -2270
rect 32600 -2305 32610 -2270
rect 32645 -2305 32655 -2270
rect 32690 -2305 32700 -2270
rect 32735 -2305 32745 -2270
rect 32780 -2305 32790 -2270
rect 32825 -2305 32835 -2270
rect 32870 -2305 32890 -2270
rect -120 -2315 32890 -2305
rect -120 -2320 31305 -2315
rect -120 -2360 -80 -2320
rect -40 -2360 270 -2320
rect 310 -2360 620 -2320
rect 660 -2360 970 -2320
rect 1010 -2360 1320 -2320
rect 1360 -2360 1670 -2320
rect 1710 -2360 2020 -2320
rect 2060 -2360 2370 -2320
rect 2410 -2360 2720 -2320
rect 2760 -2360 3070 -2320
rect 3110 -2360 5870 -2320
rect 5910 -2360 6220 -2320
rect 6260 -2360 6570 -2320
rect 6610 -2360 6920 -2320
rect 6960 -2360 7270 -2320
rect 7310 -2360 7620 -2320
rect 7660 -2360 7970 -2320
rect 8010 -2360 8320 -2320
rect 8360 -2360 8670 -2320
rect 8710 -2360 9020 -2320
rect 9060 -2350 31305 -2320
rect 31340 -2350 31350 -2315
rect 31385 -2350 31395 -2315
rect 31430 -2350 31440 -2315
rect 31475 -2350 31485 -2315
rect 31520 -2350 31530 -2315
rect 31565 -2350 31575 -2315
rect 31610 -2350 31620 -2315
rect 31655 -2350 31665 -2315
rect 31700 -2350 31710 -2315
rect 31745 -2350 31755 -2315
rect 31790 -2350 31800 -2315
rect 31835 -2350 31845 -2315
rect 31880 -2350 31890 -2315
rect 31925 -2350 31935 -2315
rect 31970 -2350 31980 -2315
rect 32015 -2350 32025 -2315
rect 32060 -2350 32070 -2315
rect 32105 -2350 32115 -2315
rect 32150 -2350 32160 -2315
rect 32195 -2350 32205 -2315
rect 32240 -2350 32250 -2315
rect 32285 -2350 32295 -2315
rect 32330 -2350 32340 -2315
rect 32375 -2350 32385 -2315
rect 32420 -2350 32430 -2315
rect 32465 -2350 32475 -2315
rect 32510 -2350 32520 -2315
rect 32555 -2350 32565 -2315
rect 32600 -2350 32610 -2315
rect 32645 -2350 32655 -2315
rect 32690 -2350 32700 -2315
rect 32735 -2350 32745 -2315
rect 32780 -2350 32790 -2315
rect 32825 -2350 32835 -2315
rect 32870 -2350 32890 -2315
rect 9060 -2360 32890 -2350
rect -120 -2390 31305 -2360
rect -120 -2430 -80 -2390
rect -40 -2430 270 -2390
rect 310 -2430 620 -2390
rect 660 -2430 970 -2390
rect 1010 -2430 1320 -2390
rect 1360 -2430 1670 -2390
rect 1710 -2430 2020 -2390
rect 2060 -2430 2370 -2390
rect 2410 -2430 2720 -2390
rect 2760 -2430 3070 -2390
rect 3110 -2430 5870 -2390
rect 5910 -2430 6220 -2390
rect 6260 -2430 6570 -2390
rect 6610 -2430 6920 -2390
rect 6960 -2430 7270 -2390
rect 7310 -2430 7620 -2390
rect 7660 -2430 7970 -2390
rect 8010 -2430 8320 -2390
rect 8360 -2430 8670 -2390
rect 8710 -2430 9020 -2390
rect 9060 -2395 31305 -2390
rect 31340 -2395 31350 -2360
rect 31385 -2395 31395 -2360
rect 31430 -2395 31440 -2360
rect 31475 -2395 31485 -2360
rect 31520 -2395 31530 -2360
rect 31565 -2395 31575 -2360
rect 31610 -2395 31620 -2360
rect 31655 -2395 31665 -2360
rect 31700 -2395 31710 -2360
rect 31745 -2395 31755 -2360
rect 31790 -2395 31800 -2360
rect 31835 -2395 31845 -2360
rect 31880 -2395 31890 -2360
rect 31925 -2395 31935 -2360
rect 31970 -2395 31980 -2360
rect 32015 -2395 32025 -2360
rect 32060 -2395 32070 -2360
rect 32105 -2395 32115 -2360
rect 32150 -2395 32160 -2360
rect 32195 -2395 32205 -2360
rect 32240 -2395 32250 -2360
rect 32285 -2395 32295 -2360
rect 32330 -2395 32340 -2360
rect 32375 -2395 32385 -2360
rect 32420 -2395 32430 -2360
rect 32465 -2395 32475 -2360
rect 32510 -2395 32520 -2360
rect 32555 -2395 32565 -2360
rect 32600 -2395 32610 -2360
rect 32645 -2395 32655 -2360
rect 32690 -2395 32700 -2360
rect 32735 -2395 32745 -2360
rect 32780 -2395 32790 -2360
rect 32825 -2395 32835 -2360
rect 32870 -2395 32890 -2360
rect 9060 -2405 32890 -2395
rect 9060 -2430 31305 -2405
rect -120 -2440 31305 -2430
rect 31340 -2440 31350 -2405
rect 31385 -2440 31395 -2405
rect 31430 -2440 31440 -2405
rect 31475 -2440 31485 -2405
rect 31520 -2440 31530 -2405
rect 31565 -2440 31575 -2405
rect 31610 -2440 31620 -2405
rect 31655 -2440 31665 -2405
rect 31700 -2440 31710 -2405
rect 31745 -2440 31755 -2405
rect 31790 -2440 31800 -2405
rect 31835 -2440 31845 -2405
rect 31880 -2440 31890 -2405
rect 31925 -2440 31935 -2405
rect 31970 -2440 31980 -2405
rect 32015 -2440 32025 -2405
rect 32060 -2440 32070 -2405
rect 32105 -2440 32115 -2405
rect 32150 -2440 32160 -2405
rect 32195 -2440 32205 -2405
rect 32240 -2440 32250 -2405
rect 32285 -2440 32295 -2405
rect 32330 -2440 32340 -2405
rect 32375 -2440 32385 -2405
rect 32420 -2440 32430 -2405
rect 32465 -2440 32475 -2405
rect 32510 -2440 32520 -2405
rect 32555 -2440 32565 -2405
rect 32600 -2440 32610 -2405
rect 32645 -2440 32655 -2405
rect 32690 -2440 32700 -2405
rect 32735 -2440 32745 -2405
rect 32780 -2440 32790 -2405
rect 32825 -2440 32835 -2405
rect 32870 -2440 32890 -2405
rect -120 -2450 32890 -2440
rect -120 -2455 31305 -2450
rect -120 -2495 -80 -2455
rect -40 -2495 270 -2455
rect 310 -2495 620 -2455
rect 660 -2495 970 -2455
rect 1010 -2495 1320 -2455
rect 1360 -2495 1670 -2455
rect 1710 -2495 2020 -2455
rect 2060 -2495 2370 -2455
rect 2410 -2495 2720 -2455
rect 2760 -2495 3070 -2455
rect 3110 -2495 5870 -2455
rect 5910 -2495 6220 -2455
rect 6260 -2495 6570 -2455
rect 6610 -2495 6920 -2455
rect 6960 -2495 7270 -2455
rect 7310 -2495 7620 -2455
rect 7660 -2495 7970 -2455
rect 8010 -2495 8320 -2455
rect 8360 -2495 8670 -2455
rect 8710 -2495 9020 -2455
rect 9060 -2485 31305 -2455
rect 31340 -2485 31350 -2450
rect 31385 -2485 31395 -2450
rect 31430 -2485 31440 -2450
rect 31475 -2485 31485 -2450
rect 31520 -2485 31530 -2450
rect 31565 -2485 31575 -2450
rect 31610 -2485 31620 -2450
rect 31655 -2485 31665 -2450
rect 31700 -2485 31710 -2450
rect 31745 -2485 31755 -2450
rect 31790 -2485 31800 -2450
rect 31835 -2485 31845 -2450
rect 31880 -2485 31890 -2450
rect 31925 -2485 31935 -2450
rect 31970 -2485 31980 -2450
rect 32015 -2485 32025 -2450
rect 32060 -2485 32070 -2450
rect 32105 -2485 32115 -2450
rect 32150 -2485 32160 -2450
rect 32195 -2485 32205 -2450
rect 32240 -2485 32250 -2450
rect 32285 -2485 32295 -2450
rect 32330 -2485 32340 -2450
rect 32375 -2485 32385 -2450
rect 32420 -2485 32430 -2450
rect 32465 -2485 32475 -2450
rect 32510 -2485 32520 -2450
rect 32555 -2485 32565 -2450
rect 32600 -2485 32610 -2450
rect 32645 -2485 32655 -2450
rect 32690 -2485 32700 -2450
rect 32735 -2485 32745 -2450
rect 32780 -2485 32790 -2450
rect 32825 -2485 32835 -2450
rect 32870 -2485 32890 -2450
rect 9060 -2495 32890 -2485
rect -120 -2515 31305 -2495
rect -120 -2555 -80 -2515
rect -40 -2555 270 -2515
rect 310 -2555 620 -2515
rect 660 -2555 970 -2515
rect 1010 -2555 1320 -2515
rect 1360 -2555 1670 -2515
rect 1710 -2555 2020 -2515
rect 2060 -2555 2370 -2515
rect 2410 -2555 2720 -2515
rect 2760 -2555 3070 -2515
rect 3110 -2555 5870 -2515
rect 5910 -2555 6220 -2515
rect 6260 -2555 6570 -2515
rect 6610 -2555 6920 -2515
rect 6960 -2555 7270 -2515
rect 7310 -2555 7620 -2515
rect 7660 -2555 7970 -2515
rect 8010 -2555 8320 -2515
rect 8360 -2555 8670 -2515
rect 8710 -2555 9020 -2515
rect 9060 -2530 31305 -2515
rect 31340 -2530 31350 -2495
rect 31385 -2530 31395 -2495
rect 31430 -2530 31440 -2495
rect 31475 -2530 31485 -2495
rect 31520 -2530 31530 -2495
rect 31565 -2530 31575 -2495
rect 31610 -2530 31620 -2495
rect 31655 -2530 31665 -2495
rect 31700 -2530 31710 -2495
rect 31745 -2530 31755 -2495
rect 31790 -2530 31800 -2495
rect 31835 -2530 31845 -2495
rect 31880 -2530 31890 -2495
rect 31925 -2530 31935 -2495
rect 31970 -2530 31980 -2495
rect 32015 -2530 32025 -2495
rect 32060 -2530 32070 -2495
rect 32105 -2530 32115 -2495
rect 32150 -2530 32160 -2495
rect 32195 -2530 32205 -2495
rect 32240 -2530 32250 -2495
rect 32285 -2530 32295 -2495
rect 32330 -2530 32340 -2495
rect 32375 -2530 32385 -2495
rect 32420 -2530 32430 -2495
rect 32465 -2530 32475 -2495
rect 32510 -2530 32520 -2495
rect 32555 -2530 32565 -2495
rect 32600 -2530 32610 -2495
rect 32645 -2530 32655 -2495
rect 32690 -2530 32700 -2495
rect 32735 -2530 32745 -2495
rect 32780 -2530 32790 -2495
rect 32825 -2530 32835 -2495
rect 32870 -2530 32890 -2495
rect 9060 -2540 32890 -2530
rect 9060 -2555 31305 -2540
rect -120 -2575 31305 -2555
rect 31340 -2575 31350 -2540
rect 31385 -2575 31395 -2540
rect 31430 -2575 31440 -2540
rect 31475 -2575 31485 -2540
rect 31520 -2575 31530 -2540
rect 31565 -2575 31575 -2540
rect 31610 -2575 31620 -2540
rect 31655 -2575 31665 -2540
rect 31700 -2575 31710 -2540
rect 31745 -2575 31755 -2540
rect 31790 -2575 31800 -2540
rect 31835 -2575 31845 -2540
rect 31880 -2575 31890 -2540
rect 31925 -2575 31935 -2540
rect 31970 -2575 31980 -2540
rect 32015 -2575 32025 -2540
rect 32060 -2575 32070 -2540
rect 32105 -2575 32115 -2540
rect 32150 -2575 32160 -2540
rect 32195 -2575 32205 -2540
rect 32240 -2575 32250 -2540
rect 32285 -2575 32295 -2540
rect 32330 -2575 32340 -2540
rect 32375 -2575 32385 -2540
rect 32420 -2575 32430 -2540
rect 32465 -2575 32475 -2540
rect 32510 -2575 32520 -2540
rect 32555 -2575 32565 -2540
rect 32600 -2575 32610 -2540
rect 32645 -2575 32655 -2540
rect 32690 -2575 32700 -2540
rect 32735 -2575 32745 -2540
rect 32780 -2575 32790 -2540
rect 32825 -2575 32835 -2540
rect 32870 -2575 32890 -2540
rect -120 -2580 32890 -2575
rect -120 -2620 -80 -2580
rect -40 -2620 270 -2580
rect 310 -2620 620 -2580
rect 660 -2620 970 -2580
rect 1010 -2620 1320 -2580
rect 1360 -2620 1670 -2580
rect 1710 -2620 2020 -2580
rect 2060 -2620 2370 -2580
rect 2410 -2620 2720 -2580
rect 2760 -2620 3070 -2580
rect 3110 -2620 5870 -2580
rect 5910 -2620 6220 -2580
rect 6260 -2620 6570 -2580
rect 6610 -2620 6920 -2580
rect 6960 -2620 7270 -2580
rect 7310 -2620 7620 -2580
rect 7660 -2620 7970 -2580
rect 8010 -2620 8320 -2580
rect 8360 -2620 8670 -2580
rect 8710 -2620 9020 -2580
rect 9060 -2585 32890 -2580
rect 9060 -2620 31305 -2585
rect 31340 -2620 31350 -2585
rect 31385 -2620 31395 -2585
rect 31430 -2620 31440 -2585
rect 31475 -2620 31485 -2585
rect 31520 -2620 31530 -2585
rect 31565 -2620 31575 -2585
rect 31610 -2620 31620 -2585
rect 31655 -2620 31665 -2585
rect 31700 -2620 31710 -2585
rect 31745 -2620 31755 -2585
rect 31790 -2620 31800 -2585
rect 31835 -2620 31845 -2585
rect 31880 -2620 31890 -2585
rect 31925 -2620 31935 -2585
rect 31970 -2620 31980 -2585
rect 32015 -2620 32025 -2585
rect 32060 -2620 32070 -2585
rect 32105 -2620 32115 -2585
rect 32150 -2620 32160 -2585
rect 32195 -2620 32205 -2585
rect 32240 -2620 32250 -2585
rect 32285 -2620 32295 -2585
rect 32330 -2620 32340 -2585
rect 32375 -2620 32385 -2585
rect 32420 -2620 32430 -2585
rect 32465 -2620 32475 -2585
rect 32510 -2620 32520 -2585
rect 32555 -2620 32565 -2585
rect 32600 -2620 32610 -2585
rect 32645 -2620 32655 -2585
rect 32690 -2620 32700 -2585
rect 32735 -2620 32745 -2585
rect 32780 -2620 32790 -2585
rect 32825 -2620 32835 -2585
rect 32870 -2620 32890 -2585
rect -120 -2630 32890 -2620
rect -120 -2650 31305 -2630
rect -120 -2690 -80 -2650
rect -40 -2690 270 -2650
rect 310 -2690 620 -2650
rect 660 -2690 970 -2650
rect 1010 -2690 1320 -2650
rect 1360 -2690 1670 -2650
rect 1710 -2690 2020 -2650
rect 2060 -2690 2370 -2650
rect 2410 -2690 2720 -2650
rect 2760 -2690 3070 -2650
rect 3110 -2690 5870 -2650
rect 5910 -2690 6220 -2650
rect 6260 -2690 6570 -2650
rect 6610 -2690 6920 -2650
rect 6960 -2690 7270 -2650
rect 7310 -2690 7620 -2650
rect 7660 -2690 7970 -2650
rect 8010 -2690 8320 -2650
rect 8360 -2690 8670 -2650
rect 8710 -2690 9020 -2650
rect 9060 -2665 31305 -2650
rect 31340 -2665 31350 -2630
rect 31385 -2665 31395 -2630
rect 31430 -2665 31440 -2630
rect 31475 -2665 31485 -2630
rect 31520 -2665 31530 -2630
rect 31565 -2665 31575 -2630
rect 31610 -2665 31620 -2630
rect 31655 -2665 31665 -2630
rect 31700 -2665 31710 -2630
rect 31745 -2665 31755 -2630
rect 31790 -2665 31800 -2630
rect 31835 -2665 31845 -2630
rect 31880 -2665 31890 -2630
rect 31925 -2665 31935 -2630
rect 31970 -2665 31980 -2630
rect 32015 -2665 32025 -2630
rect 32060 -2665 32070 -2630
rect 32105 -2665 32115 -2630
rect 32150 -2665 32160 -2630
rect 32195 -2665 32205 -2630
rect 32240 -2665 32250 -2630
rect 32285 -2665 32295 -2630
rect 32330 -2665 32340 -2630
rect 32375 -2665 32385 -2630
rect 32420 -2665 32430 -2630
rect 32465 -2665 32475 -2630
rect 32510 -2665 32520 -2630
rect 32555 -2665 32565 -2630
rect 32600 -2665 32610 -2630
rect 32645 -2665 32655 -2630
rect 32690 -2665 32700 -2630
rect 32735 -2665 32745 -2630
rect 32780 -2665 32790 -2630
rect 32825 -2665 32835 -2630
rect 32870 -2665 32890 -2630
rect 9060 -2675 32890 -2665
rect 9060 -2690 31305 -2675
rect -120 -2710 31305 -2690
rect 31340 -2710 31350 -2675
rect 31385 -2710 31395 -2675
rect 31430 -2710 31440 -2675
rect 31475 -2710 31485 -2675
rect 31520 -2710 31530 -2675
rect 31565 -2710 31575 -2675
rect 31610 -2710 31620 -2675
rect 31655 -2710 31665 -2675
rect 31700 -2710 31710 -2675
rect 31745 -2710 31755 -2675
rect 31790 -2710 31800 -2675
rect 31835 -2710 31845 -2675
rect 31880 -2710 31890 -2675
rect 31925 -2710 31935 -2675
rect 31970 -2710 31980 -2675
rect 32015 -2710 32025 -2675
rect 32060 -2710 32070 -2675
rect 32105 -2710 32115 -2675
rect 32150 -2710 32160 -2675
rect 32195 -2710 32205 -2675
rect 32240 -2710 32250 -2675
rect 32285 -2710 32295 -2675
rect 32330 -2710 32340 -2675
rect 32375 -2710 32385 -2675
rect 32420 -2710 32430 -2675
rect 32465 -2710 32475 -2675
rect 32510 -2710 32520 -2675
rect 32555 -2710 32565 -2675
rect 32600 -2710 32610 -2675
rect 32645 -2710 32655 -2675
rect 32690 -2710 32700 -2675
rect 32735 -2710 32745 -2675
rect 32780 -2710 32790 -2675
rect 32825 -2710 32835 -2675
rect 32870 -2710 32890 -2675
rect -120 -2720 32890 -2710
rect -120 -2760 -80 -2720
rect -40 -2760 270 -2720
rect 310 -2760 620 -2720
rect 660 -2760 970 -2720
rect 1010 -2760 1320 -2720
rect 1360 -2760 1670 -2720
rect 1710 -2760 2020 -2720
rect 2060 -2760 2370 -2720
rect 2410 -2760 2720 -2720
rect 2760 -2760 3070 -2720
rect 3110 -2760 5870 -2720
rect 5910 -2760 6220 -2720
rect 6260 -2760 6570 -2720
rect 6610 -2760 6920 -2720
rect 6960 -2760 7270 -2720
rect 7310 -2760 7620 -2720
rect 7660 -2760 7970 -2720
rect 8010 -2760 8320 -2720
rect 8360 -2760 8670 -2720
rect 8710 -2760 9020 -2720
rect 9060 -2755 31305 -2720
rect 31340 -2755 31350 -2720
rect 31385 -2755 31395 -2720
rect 31430 -2755 31440 -2720
rect 31475 -2755 31485 -2720
rect 31520 -2755 31530 -2720
rect 31565 -2755 31575 -2720
rect 31610 -2755 31620 -2720
rect 31655 -2755 31665 -2720
rect 31700 -2755 31710 -2720
rect 31745 -2755 31755 -2720
rect 31790 -2755 31800 -2720
rect 31835 -2755 31845 -2720
rect 31880 -2755 31890 -2720
rect 31925 -2755 31935 -2720
rect 31970 -2755 31980 -2720
rect 32015 -2755 32025 -2720
rect 32060 -2755 32070 -2720
rect 32105 -2755 32115 -2720
rect 32150 -2755 32160 -2720
rect 32195 -2755 32205 -2720
rect 32240 -2755 32250 -2720
rect 32285 -2755 32295 -2720
rect 32330 -2755 32340 -2720
rect 32375 -2755 32385 -2720
rect 32420 -2755 32430 -2720
rect 32465 -2755 32475 -2720
rect 32510 -2755 32520 -2720
rect 32555 -2755 32565 -2720
rect 32600 -2755 32610 -2720
rect 32645 -2755 32655 -2720
rect 32690 -2755 32700 -2720
rect 32735 -2755 32745 -2720
rect 32780 -2755 32790 -2720
rect 32825 -2755 32835 -2720
rect 32870 -2755 32890 -2720
rect 9060 -2760 32890 -2755
rect -120 -2765 32890 -2760
rect -120 -2790 31305 -2765
rect -120 -2830 -80 -2790
rect -40 -2830 270 -2790
rect 310 -2830 620 -2790
rect 660 -2830 970 -2790
rect 1010 -2830 1320 -2790
rect 1360 -2830 1670 -2790
rect 1710 -2830 2020 -2790
rect 2060 -2830 2370 -2790
rect 2410 -2830 2720 -2790
rect 2760 -2830 3070 -2790
rect 3110 -2830 5870 -2790
rect 5910 -2830 6220 -2790
rect 6260 -2830 6570 -2790
rect 6610 -2830 6920 -2790
rect 6960 -2830 7270 -2790
rect 7310 -2830 7620 -2790
rect 7660 -2830 7970 -2790
rect 8010 -2830 8320 -2790
rect 8360 -2830 8670 -2790
rect 8710 -2830 9020 -2790
rect 9060 -2800 31305 -2790
rect 31340 -2800 31350 -2765
rect 31385 -2800 31395 -2765
rect 31430 -2800 31440 -2765
rect 31475 -2800 31485 -2765
rect 31520 -2800 31530 -2765
rect 31565 -2800 31575 -2765
rect 31610 -2800 31620 -2765
rect 31655 -2800 31665 -2765
rect 31700 -2800 31710 -2765
rect 31745 -2800 31755 -2765
rect 31790 -2800 31800 -2765
rect 31835 -2800 31845 -2765
rect 31880 -2800 31890 -2765
rect 31925 -2800 31935 -2765
rect 31970 -2800 31980 -2765
rect 32015 -2800 32025 -2765
rect 32060 -2800 32070 -2765
rect 32105 -2800 32115 -2765
rect 32150 -2800 32160 -2765
rect 32195 -2800 32205 -2765
rect 32240 -2800 32250 -2765
rect 32285 -2800 32295 -2765
rect 32330 -2800 32340 -2765
rect 32375 -2800 32385 -2765
rect 32420 -2800 32430 -2765
rect 32465 -2800 32475 -2765
rect 32510 -2800 32520 -2765
rect 32555 -2800 32565 -2765
rect 32600 -2800 32610 -2765
rect 32645 -2800 32655 -2765
rect 32690 -2800 32700 -2765
rect 32735 -2800 32745 -2765
rect 32780 -2800 32790 -2765
rect 32825 -2800 32835 -2765
rect 32870 -2800 32890 -2765
rect 9060 -2810 32890 -2800
rect 9060 -2830 31305 -2810
rect -120 -2845 31305 -2830
rect 31340 -2845 31350 -2810
rect 31385 -2845 31395 -2810
rect 31430 -2845 31440 -2810
rect 31475 -2845 31485 -2810
rect 31520 -2845 31530 -2810
rect 31565 -2845 31575 -2810
rect 31610 -2845 31620 -2810
rect 31655 -2845 31665 -2810
rect 31700 -2845 31710 -2810
rect 31745 -2845 31755 -2810
rect 31790 -2845 31800 -2810
rect 31835 -2845 31845 -2810
rect 31880 -2845 31890 -2810
rect 31925 -2845 31935 -2810
rect 31970 -2845 31980 -2810
rect 32015 -2845 32025 -2810
rect 32060 -2845 32070 -2810
rect 32105 -2845 32115 -2810
rect 32150 -2845 32160 -2810
rect 32195 -2845 32205 -2810
rect 32240 -2845 32250 -2810
rect 32285 -2845 32295 -2810
rect 32330 -2845 32340 -2810
rect 32375 -2845 32385 -2810
rect 32420 -2845 32430 -2810
rect 32465 -2845 32475 -2810
rect 32510 -2845 32520 -2810
rect 32555 -2845 32565 -2810
rect 32600 -2845 32610 -2810
rect 32645 -2845 32655 -2810
rect 32690 -2845 32700 -2810
rect 32735 -2845 32745 -2810
rect 32780 -2845 32790 -2810
rect 32825 -2845 32835 -2810
rect 32870 -2845 32890 -2810
rect -120 -2855 32890 -2845
rect -120 -2895 -80 -2855
rect -40 -2895 270 -2855
rect 310 -2895 620 -2855
rect 660 -2895 970 -2855
rect 1010 -2895 1320 -2855
rect 1360 -2895 1670 -2855
rect 1710 -2895 2020 -2855
rect 2060 -2895 2370 -2855
rect 2410 -2895 2720 -2855
rect 2760 -2895 3070 -2855
rect 3110 -2895 5870 -2855
rect 5910 -2895 6220 -2855
rect 6260 -2895 6570 -2855
rect 6610 -2895 6920 -2855
rect 6960 -2895 7270 -2855
rect 7310 -2895 7620 -2855
rect 7660 -2895 7970 -2855
rect 8010 -2895 8320 -2855
rect 8360 -2895 8670 -2855
rect 8710 -2895 9020 -2855
rect 9060 -2890 31305 -2855
rect 31340 -2890 31350 -2855
rect 31385 -2890 31395 -2855
rect 31430 -2890 31440 -2855
rect 31475 -2890 31485 -2855
rect 31520 -2890 31530 -2855
rect 31565 -2890 31575 -2855
rect 31610 -2890 31620 -2855
rect 31655 -2890 31665 -2855
rect 31700 -2890 31710 -2855
rect 31745 -2890 31755 -2855
rect 31790 -2890 31800 -2855
rect 31835 -2890 31845 -2855
rect 31880 -2890 31890 -2855
rect 31925 -2890 31935 -2855
rect 31970 -2890 31980 -2855
rect 32015 -2890 32025 -2855
rect 32060 -2890 32070 -2855
rect 32105 -2890 32115 -2855
rect 32150 -2890 32160 -2855
rect 32195 -2890 32205 -2855
rect 32240 -2890 32250 -2855
rect 32285 -2890 32295 -2855
rect 32330 -2890 32340 -2855
rect 32375 -2890 32385 -2855
rect 32420 -2890 32430 -2855
rect 32465 -2890 32475 -2855
rect 32510 -2890 32520 -2855
rect 32555 -2890 32565 -2855
rect 32600 -2890 32610 -2855
rect 32645 -2890 32655 -2855
rect 32690 -2890 32700 -2855
rect 32735 -2890 32745 -2855
rect 32780 -2890 32790 -2855
rect 32825 -2890 32835 -2855
rect 32870 -2890 32890 -2855
rect 9060 -2895 32890 -2890
rect -120 -2905 32890 -2895
rect -38770 -3015 5600 -3005
rect -38770 -3055 3420 -3015
rect 3460 -3055 3770 -3015
rect 3810 -3055 4120 -3015
rect 4160 -3055 4470 -3015
rect 4510 -3055 4820 -3015
rect 4860 -3055 5170 -3015
rect 5210 -3055 5520 -3015
rect 5560 -3055 5600 -3015
rect -38770 -3080 5600 -3055
rect -38770 -3120 3420 -3080
rect 3460 -3120 3770 -3080
rect 3810 -3120 4120 -3080
rect 4160 -3120 4470 -3080
rect 4510 -3120 4820 -3080
rect 4860 -3120 5170 -3080
rect 5210 -3120 5520 -3080
rect 5560 -3120 5600 -3080
rect -38770 -3150 5600 -3120
rect -38770 -3190 3420 -3150
rect 3460 -3190 3770 -3150
rect 3810 -3190 4120 -3150
rect 4160 -3190 4470 -3150
rect 4510 -3190 4820 -3150
rect 4860 -3190 5170 -3150
rect 5210 -3190 5520 -3150
rect 5560 -3190 5600 -3150
rect -38770 -3220 5600 -3190
rect -38770 -3260 3420 -3220
rect 3460 -3260 3770 -3220
rect 3810 -3260 4120 -3220
rect 4160 -3260 4470 -3220
rect 4510 -3260 4820 -3220
rect 4860 -3260 5170 -3220
rect 5210 -3260 5520 -3220
rect 5560 -3260 5600 -3220
rect -38770 -3290 5600 -3260
rect -38770 -3330 3420 -3290
rect 3460 -3330 3770 -3290
rect 3810 -3330 4120 -3290
rect 4160 -3330 4470 -3290
rect 4510 -3330 4820 -3290
rect 4860 -3330 5170 -3290
rect 5210 -3330 5520 -3290
rect 5560 -3330 5600 -3290
rect -38770 -3355 5600 -3330
rect -38770 -3395 3420 -3355
rect 3460 -3395 3770 -3355
rect 3810 -3395 4120 -3355
rect 4160 -3395 4470 -3355
rect 4510 -3395 4820 -3355
rect 4860 -3395 5170 -3355
rect 5210 -3395 5520 -3355
rect 5560 -3395 5600 -3355
rect -38770 -3415 5600 -3395
rect -38770 -3455 3420 -3415
rect 3460 -3455 3770 -3415
rect 3810 -3455 4120 -3415
rect 4160 -3455 4470 -3415
rect 4510 -3455 4820 -3415
rect 4860 -3455 5170 -3415
rect 5210 -3455 5520 -3415
rect 5560 -3455 5600 -3415
rect -38770 -3480 5600 -3455
rect -38770 -3520 3420 -3480
rect 3460 -3520 3770 -3480
rect 3810 -3520 4120 -3480
rect 4160 -3520 4470 -3480
rect 4510 -3520 4820 -3480
rect 4860 -3520 5170 -3480
rect 5210 -3520 5520 -3480
rect 5560 -3520 5600 -3480
rect -38770 -3550 5600 -3520
rect -38770 -3590 3420 -3550
rect 3460 -3590 3770 -3550
rect 3810 -3590 4120 -3550
rect 4160 -3590 4470 -3550
rect 4510 -3590 4820 -3550
rect 4860 -3590 5170 -3550
rect 5210 -3590 5520 -3550
rect 5560 -3590 5600 -3550
rect -38770 -3620 5600 -3590
rect -38770 -3660 3420 -3620
rect 3460 -3660 3770 -3620
rect 3810 -3660 4120 -3620
rect 4160 -3660 4470 -3620
rect 4510 -3660 4820 -3620
rect 4860 -3660 5170 -3620
rect 5210 -3660 5520 -3620
rect 5560 -3660 5600 -3620
rect -38770 -3690 5600 -3660
rect -38770 -3730 3420 -3690
rect 3460 -3730 3770 -3690
rect 3810 -3730 4120 -3690
rect 4160 -3730 4470 -3690
rect 4510 -3730 4820 -3690
rect 4860 -3730 5170 -3690
rect 5210 -3730 5520 -3690
rect 5560 -3730 5600 -3690
rect -38770 -3755 5600 -3730
rect -38770 -3795 3420 -3755
rect 3460 -3795 3770 -3755
rect 3810 -3795 4120 -3755
rect 4160 -3795 4470 -3755
rect 4510 -3795 4820 -3755
rect 4860 -3795 5170 -3755
rect 5210 -3795 5520 -3755
rect 5560 -3795 5600 -3755
rect -38770 -3815 5600 -3795
rect -38770 -3855 3420 -3815
rect 3460 -3855 3770 -3815
rect 3810 -3855 4120 -3815
rect 4160 -3855 4470 -3815
rect 4510 -3855 4820 -3815
rect 4860 -3855 5170 -3815
rect 5210 -3855 5520 -3815
rect 5560 -3855 5600 -3815
rect -38770 -3880 5600 -3855
rect -38770 -3920 3420 -3880
rect 3460 -3920 3770 -3880
rect 3810 -3920 4120 -3880
rect 4160 -3920 4470 -3880
rect 4510 -3920 4820 -3880
rect 4860 -3920 5170 -3880
rect 5210 -3920 5520 -3880
rect 5560 -3920 5600 -3880
rect -38770 -3950 5600 -3920
rect -38770 -3990 3420 -3950
rect 3460 -3990 3770 -3950
rect 3810 -3990 4120 -3950
rect 4160 -3990 4470 -3950
rect 4510 -3990 4820 -3950
rect 4860 -3990 5170 -3950
rect 5210 -3990 5520 -3950
rect 5560 -3990 5600 -3950
rect -38770 -4020 5600 -3990
rect -38770 -4060 3420 -4020
rect 3460 -4060 3770 -4020
rect 3810 -4060 4120 -4020
rect 4160 -4060 4470 -4020
rect 4510 -4060 4820 -4020
rect 4860 -4060 5170 -4020
rect 5210 -4060 5520 -4020
rect 5560 -4060 5600 -4020
rect -38770 -4090 5600 -4060
rect -38770 -4130 3420 -4090
rect 3460 -4130 3770 -4090
rect 3810 -4130 4120 -4090
rect 4160 -4130 4470 -4090
rect 4510 -4130 4820 -4090
rect 4860 -4130 5170 -4090
rect 5210 -4130 5520 -4090
rect 5560 -4130 5600 -4090
rect -38770 -4155 5600 -4130
rect -38770 -4195 3420 -4155
rect 3460 -4195 3770 -4155
rect 3810 -4195 4120 -4155
rect 4160 -4195 4470 -4155
rect 4510 -4195 4820 -4155
rect 4860 -4195 5170 -4155
rect 5210 -4195 5520 -4155
rect 5560 -4195 5600 -4155
rect -38770 -4215 5600 -4195
rect -38770 -4255 3420 -4215
rect 3460 -4255 3770 -4215
rect 3810 -4255 4120 -4215
rect 4160 -4255 4470 -4215
rect 4510 -4255 4820 -4215
rect 4860 -4255 5170 -4215
rect 5210 -4255 5520 -4215
rect 5560 -4255 5600 -4215
rect -38770 -4280 5600 -4255
rect -38770 -4320 3420 -4280
rect 3460 -4320 3770 -4280
rect 3810 -4320 4120 -4280
rect 4160 -4320 4470 -4280
rect 4510 -4320 4820 -4280
rect 4860 -4320 5170 -4280
rect 5210 -4320 5520 -4280
rect 5560 -4320 5600 -4280
rect -38770 -4350 5600 -4320
rect -38770 -4390 3420 -4350
rect 3460 -4390 3770 -4350
rect 3810 -4390 4120 -4350
rect 4160 -4390 4470 -4350
rect 4510 -4390 4820 -4350
rect 4860 -4390 5170 -4350
rect 5210 -4390 5520 -4350
rect 5560 -4390 5600 -4350
rect -38770 -4420 5600 -4390
rect -38770 -4460 3420 -4420
rect 3460 -4460 3770 -4420
rect 3810 -4460 4120 -4420
rect 4160 -4460 4470 -4420
rect 4510 -4460 4820 -4420
rect 4860 -4460 5170 -4420
rect 5210 -4460 5520 -4420
rect 5560 -4460 5600 -4420
rect -38770 -4490 5600 -4460
rect -38770 -4530 3420 -4490
rect 3460 -4530 3770 -4490
rect 3810 -4530 4120 -4490
rect 4160 -4530 4470 -4490
rect 4510 -4530 4820 -4490
rect 4860 -4530 5170 -4490
rect 5210 -4530 5520 -4490
rect 5560 -4530 5600 -4490
rect -38770 -4555 5600 -4530
rect -38770 -4595 3420 -4555
rect 3460 -4595 3770 -4555
rect 3810 -4595 4120 -4555
rect 4160 -4595 4470 -4555
rect 4510 -4595 4820 -4555
rect 4860 -4595 5170 -4555
rect 5210 -4595 5520 -4555
rect 5560 -4595 5600 -4555
rect -38770 -4605 5600 -4595
use bgr_11  bgr_11_0
timestamp 1756070769
transform -1 0 22290 0 -1 11375
box 15640 -6260 19905 1640
use two_stage_opamp_dummy_magic_29  two_stage_opamp_dummy_magic_29_0
timestamp 1756064335
transform 1 0 -52410 0 1 85
box 51710 -1500 62090 6110
<< labels >>
flabel metal4 35620 6650 35620 6650 3 FreeSans 800 0 320 0 GNDA
port 2 e
flabel metal3 -37570 10155 -37570 10155 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal3 -38005 5940 -38005 5940 5 FreeSans 800 0 0 -400 VDDA_2
port 8 s
flabel metal4 -38770 -3785 -38770 -3785 7 FreeSans 800 0 -400 0 GNDA_2
port 7 w
flabel metal2 6795 850 6795 850 5 FreeSans 800 0 0 -400 VOUT-
port 4 s
flabel metal2 2185 850 2185 850 5 FreeSans 800 0 0 -400 VOUT+
port 3 s
flabel metal2 5375 1590 5375 1590 3 FreeSans 400 0 160 0 VIN-
port 6 e
flabel metal2 3605 1590 3605 1590 7 FreeSans 400 0 -160 0 VIN+
port 5 w
<< end >>
