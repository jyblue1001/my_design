* NGSPICE file created from bgr_opamp_dummy_magic_16.ext - technology: sky130A

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt bgr_11 ERR_AMP_REF V_CMFB_S3 VB1_CUR_BIAS TAIL_CUR_MIR_BIAS V_CMFB_S1 ERR_AMP_CUR_BIAS
+ VB3_CUR_BIAS V_CMFB_S4 V_CMFB_S2 VB2_CUR_BIAS a_34140_n1650# a_32560_n7778# a_37640_n2290#
+ w_32750_1090# a_33140_n1680# m1_35910_n8890# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ w_32720_n90# w_33500_2220# a_35550_n8610#
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23 Vin- sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
+ m=1
X0 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA V_CMFB_S2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X2 V_mir2 V_mir2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X3 VB2_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X4 a_38570_n6504# a_38690_n7778# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X5 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base V_CMFB_S2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA V_CMFB_S4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X8 V_p_1 Vin+ 1st_Vout_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X9 VB2_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X10 V_p_2 ERR_AMP_REF V_mir2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X11 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base START_UP_NFET1 START_UP_NFET1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X13 w_33500_2220# w_33500_2220# V_CMFB_S1 w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X14 V_TOP START_UP Vin- w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X15 V_CMFB_S3 w_33500_2220# w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA VB3_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X17 VB3_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X18 NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X19 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X21 1st_Vout_2 V_mir2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X22 V_p_1 Vin- V_mir1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X23 V_p_2 a_33140_n1680# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X24 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 V_CUR_REF_REG a_32320_n7778# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=4
X26 VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X27 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 w_32750_1090# V_TOP ERR_AMP_REF w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X30 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 w_33500_2220# PFET_GATE_10uA V_CMFB_S1 w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X32 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VB2_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X34 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 w_32750_1090# PFET_GATE_10uA VB1_CUR_BIAS w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X36 w_32750_1090# w_32750_1090# VB1_CUR_BIAS w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X37 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 w_32720_n90# V_mir1 V_mir1 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X41 Vin+ V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X42 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 V_mir1 Vin- V_p_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X45 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 TAIL_CUR_MIR_BIAS PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 w_32720_n90# V_mir2 V_mir2 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X49 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 ERR_AMP_REF w_32750_1090# w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X51 V_mir1 Vin- V_p_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X52 1st_Vout_1 V_mir1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 V_CMFB_S3 PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X56 w_32750_1090# V_TOP Vin+ w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X57 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Emitter Vin+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X59 w_33500_2220# PFET_GATE_10uA NFET_GATE_10uA w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X60 PFET_GATE_10uA 1st_Vout_2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X61 1st_Vout_1 Vin+ V_p_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X62 w_32720_n90# V_mir2 1st_Vout_2 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base VB3_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X64 TAIL_CUR_MIR_BIAS PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X65 w_32720_n90# 1st_Vout_2 PFET_GATE_10uA w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X66 V_p_1 Vin+ 1st_Vout_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X67 V_CMFB_S3 PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X68 w_32720_n90# w_32720_n90# V_TOP w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X69 V_CMFB_S2 NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X70 V_CMFB_S2 NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X71 V_CMFB_S1 PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X72 Vin+ a_38040_n7928# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=6
X73 1st_Vout_1 V_mir1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X74 TAIL_CUR_MIR_BIAS PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X75 V_mir1 V_mir1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X76 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base a_33140_n1680# PFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X78 w_32720_n90# 1st_Vout_1 V_TOP w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 PFET_GATE_10uA 1st_Vout_2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X80 V_p_2 ERR_AMP_REF V_mir2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X81 V_TOP a_33140_n1680# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X82 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VB3_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA ERR_AMP_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X85 w_32720_n90# V_mir1 1st_Vout_1 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X86 V_p_1 Vin+ 1st_Vout_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X87 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 V_CMFB_S1 w_33500_2220# w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X90 w_32720_n90# V_mir2 1st_Vout_2 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X91 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 w_32720_n90# 1st_Vout_2 PFET_GATE_10uA w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X93 V_p_2 V_CUR_REF_REG 1st_Vout_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X94 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 NFET_GATE_10uA w_33500_2220# w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X96 TAIL_CUR_MIR_BIAS PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X97 V_TOP w_32720_n90# w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X98 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 V_CUR_REF_REG PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X100 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 V_CMFB_S4 NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X103 V_mir2 V_mir2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X104 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA V_CMFB_S4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X106 1st_Vout_2 V_mir2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X107 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 Vin- a_32970_n7928# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=6
X111 w_32750_1090# w_32750_1090# V_TOP w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.2 ps=1.4 w=1 l=0.15
X112 w_32750_1090# V_TOP Vin- w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X113 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 a_32440_n6570# a_32320_n7778# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=4
X115 ERR_AMP_REF V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X116 w_32720_n90# V_mir1 1st_Vout_1 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X117 1st_Vout_2 V_CUR_REF_REG V_p_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X118 w_32720_n90# V_mir1 V_mir1 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X119 Vin+ V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X120 V_mir1 Vin- V_p_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X121 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 a_38570_n6504# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X123 a_33090_n6320# a_32560_n7778# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=6
X124 V_mir1 V_mir1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X125 w_32720_n90# w_32720_n90# PFET_GATE_10uA w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base a_33140_n1680# V_p_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X127 V_CMFB_S1 PFET_GATE_10uA w_33500_2220# w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X128 Vin- START_UP V_TOP w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X129 V_TOP 1st_Vout_1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 V_mir2 ERR_AMP_REF V_p_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X131 Vin- V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X132 a_37920_n6320# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=6
X133 V_mir2 V_mir2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X134 PFET_GATE_10uA cap_res2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_high_po_0p35 l=2.05
X135 w_32750_1090# V_TOP START_UP w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X136 1st_Vout_2 V_mir2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X137 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 w_32720_n90# 1st_Vout_2 PFET_GATE_10uA w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X139 V_TOP cap_res1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_high_po_0p35 l=2.05
X140 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 w_32750_1090# V_TOP ERR_AMP_REF w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X142 w_32720_n90# V_mir2 V_mir2 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X143 w_33500_2220# PFET_GATE_10uA TAIL_CUR_MIR_BIAS w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X144 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X147 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 w_32750_1090# V_TOP START_UP w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X149 VB1_CUR_BIAS w_32750_1090# w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X150 VB1_CUR_BIAS PFET_GATE_10uA w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X151 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X152 w_33500_2220# w_33500_2220# V_CMFB_S3 w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X153 START_UP_NFET1 START_UP START_UP sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X154 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 PFET_GATE_10uA w_32720_n90# w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X156 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 V_p_1 Vin- V_mir1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X158 V_p_2 V_CUR_REF_REG 1st_Vout_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X159 START_UP V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X160 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VB3_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X163 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA VB3_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X165 ERR_AMP_CUR_BIAS NFET_GATE_10uA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X166 w_33500_2220# PFET_GATE_10uA TAIL_CUR_MIR_BIAS w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X167 ERR_AMP_REF V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X168 V_TOP 1st_Vout_1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X169 V_p_2 ERR_AMP_REF V_mir2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X170 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 1st_Vout_1 V_mir1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X172 ERR_AMP_REF a_38690_n7778# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X173 START_UP V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X174 w_32720_n90# V_mir1 V_mir1 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X175 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X176 w_33500_2220# PFET_GATE_10uA V_CMFB_S3 w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X177 w_32720_n90# 1st_Vout_1 V_TOP w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X178 V_TOP w_32750_1090# w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X179 w_32720_n90# V_mir2 V_mir2 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X180 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base NFET_GATE_10uA VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X181 V_CMFB_S4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X182 w_32750_1090# V_TOP Vin- w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X183 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 w_32720_n90# V_mir2 1st_Vout_2 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X185 a_33090_n6320# a_32970_n7928# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=6
X186 w_33500_2220# PFET_GATE_10uA TAIL_CUR_MIR_BIAS w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X187 w_32750_1090# V_TOP Vin+ w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X188 PFET_GATE_10uA 1st_Vout_2 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X189 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 w_33500_2220# PFET_GATE_10uA V_CMFB_S3 w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X192 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 1st_Vout_1 Vin+ V_p_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X194 V_mir2 ERR_AMP_REF V_p_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X195 w_33500_2220# PFET_GATE_10uA V_CMFB_S1 w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X196 V_TOP 1st_Vout_1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X197 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 Vin- V_TOP w_32750_1090# w_32750_1090# sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X199 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 w_33500_2220# PFET_GATE_10uA TAIL_CUR_MIR_BIAS w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X201 w_33500_2220# w_33500_2220# V_CUR_REF_REG w_33500_2220# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X202 1st_Vout_2 V_CUR_REF_REG V_p_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X203 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 1st_Vout_1 cap_res1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 a_37920_n6320# a_38040_n7928# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=6
X206 w_32720_n90# 1st_Vout_1 V_TOP w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 1st_Vout_2 V_CUR_REF_REG V_p_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X209 w_32750_1090# w_32750_1090# ERR_AMP_REF w_32750_1090# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X210 w_32720_n90# V_mir1 1st_Vout_1 w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X211 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 1st_Vout_2 cap_res2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 a_32440_n6570# a_32560_n7778# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8/Base sky130_fd_pr__res_xhigh_po_0p35 l=4
X215 V_TOP m1_35910_n8890# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 V_mir1 V_mir1 w_32720_n90# w_32720_n90# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
.ends

.subckt two_stage_opamp_dummy_magic_23 V_CMFB_S1 V_CMFB_S3 Vb3 Vb2 Vb1 V_CMFB_S2 V_CMFB_S4
+ VOUT- VOUT+ V_err_amp_ref V_err_gate a_109830_3220# V_tail_gate w_109730_7340# VIN-
+ VIN+
X0 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1 VD2 VIN+ V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X2 w_109730_7340# Vb3 VD3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X3 V_err_p V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X4 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VD2 Vb1 Y a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X7 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 VD1 Vb1 X a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X11 VOUT- X w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X12 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 w_109730_7340# Y V_CMFB_S4 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X14 V_CMFB_S1 X a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X15 w_109730_7340# Y V_CMFB_S4 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X16 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 w_109730_7340# w_109730_7340# VD3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X18 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 w_109730_7340# V_err_gate a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X21 a_109830_3220# err_amp_mir err_amp_mir a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X22 a_109830_3220# a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=48.8 ps=279.2 w=2.5 l=0.15
X23 a_109830_3220# a_109830_3220# err_amp_mir a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X24 Y Vb1 VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X25 Vb1 Vb1 a_113080_1090# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X26 w_109730_7340# V_err_gate V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X27 V_source VIN- VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X28 Vb2_2 Vb2_2 Vb2_2 Vb2_2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=4.92 ps=27.8 w=3.5 l=0.2
X29 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 a_118270_3858# V_tot a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X31 a_109830_3220# V_b_2nd_stage VOUT- a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X32 VD4 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X33 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X34 VOUT+ Y w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X35 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 V_err_gate V_err_amp_ref a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X37 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 err_amp_out V_err_amp_ref V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X43 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X46 a_112280_5790# V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X47 V_CMFB_S3 Y a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X48 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X49 a_109830_3220# a_109830_3220# VOUT- a_109830_3220# sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X50 w_109730_7340# w_109730_7340# a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X51 VD1 Vb1 X a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X52 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VD4 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X54 VOUT- X w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X55 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 V_CMFB_S1 X a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X63 w_109730_7340# w_109730_7340# a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X64 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 w_109730_7340# V_err_gate V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 a_109830_3220# err_amp_mir err_amp_out a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X68 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X69 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 V_source VIN- VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X71 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 w_109730_7340# a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X75 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 w_109730_7340# a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X78 VOUT+ Y w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X79 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 w_109730_7340# Vb3 VD4 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X81 VOUT+ Y w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X82 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 V_err_gate V_tot a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X87 err_amp_out V_err_amp_ref V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X88 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 err_amp_mir V_tot V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X90 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X92 V_CMFB_S3 Y a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X93 a_109830_3220# a_109830_3220# V_tail_gate a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X94 VD2 VIN+ V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X95 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT- a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X98 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VD1 Vb1 X a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X100 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 V_CMFB_S2 X w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X102 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 a_112280_5790# V_tot V_err_gate w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X106 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VOUT- V_b_2nd_stage a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X109 V_CMFB_S1 X a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X110 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 Y Vb1 VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X115 w_109730_7340# Vb3 VD4 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X116 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 X VD3 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X123 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 V_CMFB_S4 Y w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X128 V_err_gate w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X129 a_109830_3220# a_109830_3220# w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X130 err_amp_mir V_tot V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X131 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 V_err_p V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X136 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X137 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X138 V_CMFB_S3 Y a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X139 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 V_p_mir VIN+ V_tail_gate a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X143 VD2 VIN+ V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 w_109730_7340# w_109730_7340# VD4 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X145 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VOUT+ w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X147 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT- w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X149 V_CMFB_S2 X w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X150 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 a_109830_3220# a_109830_3220# w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X152 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 a_109830_3220# a_109830_3220# V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X160 V_CMFB_S1 X a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X161 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 w_109730_7340# V_err_gate V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X163 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 Y Vb1 VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X165 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 w_109730_7340# X VOUT- w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X167 a_109830_3220# a_109830_3220# VOUT+ a_109830_3220# sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X168 VOUT- a_117950_946# a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X169 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 V_CMFB_S4 Y w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X171 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 err_amp_out V_err_amp_ref V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X177 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X180 a_112280_5790# V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X181 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X182 VD2 VIN+ V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X183 V_CMFB_S3 Y a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X184 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 VD1 VIN- V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X186 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 Vb2_Vb3 Vb2_Vb3 Vb2_Vb3 Vb2_Vb3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=5.6 ps=31.2 w=3.5 l=0.2
X188 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 w_109730_7340# Y VOUT+ w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X190 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 V_CMFB_S2 X w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X192 w_109730_7340# w_109730_7340# VOUT+ w_109730_7340# sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X193 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X200 w_109730_7340# w_109730_7340# V_err_gate w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X201 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 cap_res_X X a_109830_3220# sky130_fd_pr__res_high_po_1p41 l=1.41
X204 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X205 VD4 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X206 a_109830_3220# err_amp_mir err_amp_out a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X207 Y Vb1 VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X208 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X210 X Vb1 VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X211 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 w_109730_7340# X VOUT- w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X213 w_109730_7340# w_109730_7340# VOUT- w_109730_7340# sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X214 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 VOUT+ a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X216 Vb2_Vb3 w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X217 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 V_CMFB_S4 Y w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X221 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 err_amp_mir w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X223 err_amp_mir err_amp_mir a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X224 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X225 Vb2_Vb3 Vb2_Vb3 Vb3 Vb2_Vb3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X226 V_err_p V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X227 VD2 VIN+ V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X228 V_err_p V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X229 a_109830_3220# a_109830_3220# Vb1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X230 V_CMFB_S3 Y a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X231 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VOUT+ V_b_2nd_stage a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X234 VD1 VIN- V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X235 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VD1 VIN- V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X238 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 a_109020_3958# V_tot a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X242 w_109730_7340# Y VOUT+ w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X243 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 V_CMFB_S2 X w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X245 a_112280_5790# V_err_amp_ref V_err_gate w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X246 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 VD4 w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X248 VOUT+ V_b_2nd_stage a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X249 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X250 V_CMFB_S1 X a_109830_3220# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X251 Y VD4 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X252 VD3 w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X253 w_109730_7340# w_109730_7340# V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X254 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X255 V_source VIN+ VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X256 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 Y Vb1 VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X261 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 X Vb1 VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X263 X Vb1 VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X264 w_109730_7340# X VOUT- w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X265 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 V_CMFB_S4 Y w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X273 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X274 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 VD3 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X276 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 err_amp_out err_amp_mir a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X280 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 V_p_mir V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X282 VD2 Vb1 Y a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X283 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 a_112280_5790# V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X285 a_113080_1090# Vb1 Vb1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X286 VD2 a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X287 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 VD1 VIN- V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X289 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 Vb3 Vb2 Vb2_Vb3 Vb2_Vb3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X291 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X294 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 w_109730_7340# Y VOUT+ w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X296 a_112280_5790# V_err_amp_ref V_err_gate w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X297 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 w_109730_7340# Vb3 VD4 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X300 w_109730_7340# w_109730_7340# err_amp_out w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X301 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 w_109730_7340# V_err_gate a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X304 V_source Vb1 a_113080_1090# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X305 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X306 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 Y a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X309 X Vb1 VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X310 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 w_109730_7340# Vb3 Vb2_Vb3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X312 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X314 w_109730_7340# X VOUT- w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X315 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT- V_b_2nd_stage a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X321 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 V_CMFB_S4 Y w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X325 a_109830_3220# X V_CMFB_S1 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X326 V_b_2nd_stage a_109420_936# a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X327 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 a_112280_5790# V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X330 err_amp_mir err_amp_mir a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X331 err_amp_mir err_amp_mir a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X333 a_113080_1090# Vb1 Vb1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X334 VD1 VIN- V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X335 a_109020_3958# V_CMFB_S3 a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X336 Vb2_2 Vb2 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X337 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 V_CMFB_S2 X w_109730_7340# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X340 w_109730_7340# Y VOUT+ w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X341 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X347 a_112280_5790# V_tot V_err_gate w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X348 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 w_109730_7340# Vb3 VD3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X350 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 V_err_p V_err_amp_ref err_amp_out w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X353 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 V_err_p V_tot err_amp_mir w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X356 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X358 w_109730_7340# V_err_gate V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X359 a_109830_3220# Y V_CMFB_S3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X360 a_109830_3220# a_109830_3220# VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X361 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 X Vb1 VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X365 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X370 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 w_109730_7340# Vb3 VD3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X374 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 a_109830_3220# X V_CMFB_S1 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X376 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 a_109830_3220# X V_CMFB_S1 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X378 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 V_err_p w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X380 err_amp_out err_amp_mir a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X381 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X382 a_109830_3220# a_109830_3220# Y a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X383 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VD1 a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X386 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X387 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 a_109830_3220# V_b_2nd_stage VOUT- a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X393 w_109730_7340# w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=65.96 ps=373 w=1.8 l=0.2
X394 VD4 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X395 w_109730_7340# Y VOUT+ w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X396 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 a_112280_5790# V_err_amp_ref V_err_gate w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X398 V_err_p V_tot err_amp_mir w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X399 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X401 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 a_109830_3220# Y V_CMFB_S3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X404 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 V_tail_gate VIN- V_p_mir a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X406 V_source VIN+ VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X407 w_109730_7340# w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X408 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X410 w_109730_7340# Vb3 VD3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X411 X a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X412 w_109730_7340# X VOUT- w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X413 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 w_109730_7340# X V_CMFB_S2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X415 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 V_err_gate V_tot a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X417 VOUT+ a_109420_936# a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X418 Vb2 Vb2_2 Vb2_2 Vb2_2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X419 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 a_109830_3220# X V_CMFB_S1 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X425 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 a_108900_3958# V_CMFB_S4 a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X427 a_112280_5790# V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X428 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VD2 Vb1 Y a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X430 w_109730_7340# w_109730_7340# Vb2_2 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X431 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X433 VD3 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X434 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 w_109730_7340# Y V_CMFB_S4 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X436 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 V_err_p V_err_amp_ref err_amp_out w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X439 VD4 VD4 Y VD4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X440 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 w_109730_7340# V_err_gate a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X442 Vb1 a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X443 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X444 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X446 V_source VIN+ VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X447 a_109830_3220# Y V_CMFB_S3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X448 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 V_tail_gate a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X450 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 cap_res_Y Y a_109830_3220# sky130_fd_pr__res_high_po_1p41 l=1.41
X452 a_109830_3220# a_109830_3220# VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X453 VD3 VD3 X VD3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X454 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 w_109730_7340# X V_CMFB_S2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X456 VD3 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X457 V_b_2nd_stage a_117950_946# a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X458 w_109730_7340# X V_CMFB_S2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X459 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 a_109830_3220# X V_CMFB_S1 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X466 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 V_source err_amp_out a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X468 a_118270_3858# V_CMFB_S2 a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X469 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 w_109730_7340# Vb3 VD4 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X473 V_err_p V_err_gate w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X474 VD2 Vb1 Y a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X475 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X476 VD3 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X477 a_109830_3220# a_109830_3220# X a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X478 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VOUT- X w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X480 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 w_109730_7340# Y V_CMFB_S4 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X487 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 V_err_p V_tot err_amp_mir w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X492 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X493 a_109830_3220# err_amp_mir err_amp_mir a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X494 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 w_109730_7340# V_err_gate V_err_p w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X496 a_109830_3220# V_tail_gate V_source a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X497 V_source VIN+ VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X498 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X499 a_109830_3220# Y V_CMFB_S3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X500 VD3 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X501 a_109830_3220# Y V_CMFB_S3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X502 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 V_source VIN- VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X504 V_source VIN- VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X505 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 Vb2_2 Vb2 Vb2 Vb2_2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X509 VOUT+ Y w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X510 a_118390_3858# V_tot a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X511 w_109730_7340# X V_CMFB_S2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X512 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X517 V_err_gate V_tot a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X518 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 a_109830_3220# V_b_2nd_stage VOUT+ a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X521 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 V_source V_tail_gate a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X523 err_amp_out a_109830_3220# a_109830_3220# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X524 VD2 Vb1 Y a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X525 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X528 VD1 Vb1 X a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X529 VD1 Vb1 X a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X530 VOUT- X w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X531 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 w_109730_7340# Vb3 VD3 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X534 VOUT- X w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X535 a_108900_3958# V_tot a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X536 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 a_109830_3220# V_b_2nd_stage VOUT+ a_109830_3220# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X538 w_109730_7340# Vb3 VD4 w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X539 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 w_109730_7340# Y V_CMFB_S4 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X544 a_109830_3220# err_amp_mir err_amp_out a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X545 a_109830_3220# V_tail_gate V_p_mir a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X546 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 w_109730_7340# V_err_gate a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X548 w_109730_7340# V_err_gate a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X549 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 Vb1 Vb1 a_113080_1090# a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X552 V_source VIN+ VD2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X553 V_source VIN- VD1 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X554 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 VOUT+ Y w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X562 w_109730_7340# X V_CMFB_S2 a_109830_3220# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X563 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 V_err_gate V_err_amp_ref a_112280_5790# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X565 a_109830_3220# w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X566 a_118390_3858# V_CMFB_S1 a_109830_3220# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X567 VD4 Vb3 w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X568 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 a_109830_3220# w_109730_7340# w_109730_7340# w_109730_7340# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X571 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt bgr_opamp_dummy_magic_16 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
Xbgr_11_0 bgr_11_0/ERR_AMP_REF bgr_11_0/V_CMFB_S3 bgr_11_0/VB1_CUR_BIAS bgr_11_0/TAIL_CUR_MIR_BIAS
+ bgr_11_0/V_CMFB_S1 bgr_11_0/ERR_AMP_CUR_BIAS bgr_11_0/VB3_CUR_BIAS bgr_11_0/V_CMFB_S4
+ bgr_11_0/V_CMFB_S2 bgr_11_0/VB2_CUR_BIAS GNDA GNDA GNDA VDDA VDDA VDDA GNDA VDDA
+ VDDA GNDA bgr_11
Xtwo_stage_opamp_dummy_magic_23_0 bgr_11_0/V_CMFB_S1 bgr_11_0/V_CMFB_S3 bgr_11_0/VB3_CUR_BIAS
+ bgr_11_0/VB2_CUR_BIAS bgr_11_0/VB1_CUR_BIAS bgr_11_0/V_CMFB_S2 bgr_11_0/V_CMFB_S4
+ VOUT- VOUT+ bgr_11_0/ERR_AMP_REF bgr_11_0/ERR_AMP_CUR_BIAS GNDA bgr_11_0/TAIL_CUR_MIR_BIAS
+ VDDA VIN- VIN+ two_stage_opamp_dummy_magic_23
.ends

