* PEX produced on Sat Feb  1 12:18:36 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from div3_2.ext - technology: sky130A

.subckt div3_2
X0 C.t3 A.t2 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1 VDDA.t1 I.t2 VOUT.t2 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X2 VOUT.t0 I.t3 GNDA.t26 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X3 D.t1 CLK.t3 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X4 C.t0 CLK.t4 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X5 GNDA.t13 VIN CLK.t0 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X6 GNDA.t17 CLK.t5 H.t2 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X7 GNDA.t24 I.t4 G.t1 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 I.t0 CLK.t6 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 VDDA.t15 D.t2 E.t0 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X10 GNDA.t7 CLK.t7 C.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 GNDA.t15 CLK.t8 H.t1 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 A.t0 CLK.t9 B.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 F.t1 CLK.t10 E.t1 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 CLK.t2 VIN VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X15 VDDA.t11 VOUT.t3 A.t1 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 VOUT.t1 I.t5 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 I.t1 H.t4 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X18 GNDA.t9 CLK.t11 C.t2 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X19 VDDA.t5 VIN CLK.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X20 E.t2 I.t6 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X21 D.t0 C.t4 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X22 H.t0 CLK.t12 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X23 G.t0 D.t3 F.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X24 VDDA.t17 E.t3 H.t3 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X25 B.t0 VOUT.t4 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
R0 A.n0 A.t1 713.933
R1 A.n0 A.t2 314.233
R2 A.t0 A.n0 308.2
R3 VDDA.t12 VDDA.t14 2307.14
R4 VDDA.t8 VDDA.t2 2126.19
R5 VDDA.t18 VDDA.t16 1492.86
R6 VDDA.t10 VDDA.t6 1130.95
R7 VDDA.n4 VDDA.t20 927.381
R8 VDDA.n0 VDDA.t1 673.375
R9 VDDA.n0 VDDA.t3 673.101
R10 VDDA.n1 VDDA.t13 667.592
R11 VDDA.n4 VDDA.t12 610.715
R12 VDDA VDDA.n6 594.301
R13 VDDA.n0 VDDA.n5 594.301
R14 VDDA.n0 VDDA.n3 594.301
R15 VDDA.n0 VDDA.n2 594.301
R16 VDDA.t2 VDDA.t0 497.62
R17 VDDA.t16 VDDA.t8 497.62
R18 VDDA.t14 VDDA.t18 497.62
R19 VDDA.t20 VDDA.t10 497.62
R20 VDDA.t6 VDDA.t4 497.62
R21 VDDA.n1 VDDA.n4 373.793
R22 VDDA.n6 VDDA.t7 78.8005
R23 VDDA.n6 VDDA.t5 78.8005
R24 VDDA.n5 VDDA.t21 78.8005
R25 VDDA.n5 VDDA.t11 78.8005
R26 VDDA.n3 VDDA.t19 78.8005
R27 VDDA.n3 VDDA.t15 78.8005
R28 VDDA.n2 VDDA.t9 78.8005
R29 VDDA.n2 VDDA.t17 78.8005
R30 VDDA VDDA.n0 2.788
R31 VDDA.n1 VDDA.n0 2.75546
R32 C.n0 C.t3 721.4
R33 C.n1 C.t4 350.349
R34 C.n0 C.t2 276.733
R35 C.n2 C.n1 206.333
R36 C.n1 C.n0 48.0005
R37 C.n2 C.t1 48.0005
R38 C.t0 C.n2 48.0005
R39 I.n0 I.t0 663.801
R40 I.n0 I.t6 568.067
R41 I.t6 I.t4 514.134
R42 I.n3 I.n2 344.8
R43 I.n1 I.t2 289.2
R44 I.t1 I.n3 275.454
R45 I.n2 I.t3 241
R46 I.n1 I.t5 112.468
R47 I.n3 I.n0 97.9205
R48 I.n2 I.n1 64.2672
R49 VOUT.n0 VOUT.t4 4546.23
R50 VOUT.t4 VOUT.t3 819.4
R51 VOUT.n1 VOUT.n0 633
R52 VOUT.n0 VOUT.t0 261.8
R53 VOUT.t2 VOUT.n1 78.8005
R54 VOUT.n1 VOUT.t1 78.8005
R55 GNDA.t5 GNDA.t3 3723.08
R56 GNDA.t8 GNDA.t18 3723.08
R57 GNDA.t21 GNDA.t25 2820.51
R58 GNDA.n4 GNDA.t14 2200
R59 GNDA.n4 GNDA.t23 1523.08
R60 GNDA.t16 GNDA.t21 1241.03
R61 GNDA.t19 GNDA.t16 1241.03
R62 GNDA.t14 GNDA.t19 1241.03
R63 GNDA.t23 GNDA.t2 1241.03
R64 GNDA.t2 GNDA.t5 1241.03
R65 GNDA.t3 GNDA.t6 1241.03
R66 GNDA.t6 GNDA.t0 1241.03
R67 GNDA.t0 GNDA.t8 1241.03
R68 GNDA.t18 GNDA.t10 1241.03
R69 GNDA.t10 GNDA.t12 1241.03
R70 GNDA.n1 GNDA.n4 1173.79
R71 GNDA.n0 GNDA.t26 242.613
R72 GNDA GNDA.n7 194.3
R73 GNDA GNDA.n5 194.3
R74 GNDA.n0 GNDA.n3 194.3
R75 GNDA.n0 GNDA.n2 194.3
R76 GNDA GNDA.n6 194.3
R77 GNDA.n7 GNDA.t11 48.0005
R78 GNDA.n7 GNDA.t13 48.0005
R79 GNDA.n5 GNDA.t4 48.0005
R80 GNDA.n5 GNDA.t7 48.0005
R81 GNDA.n3 GNDA.t20 48.0005
R82 GNDA.n3 GNDA.t15 48.0005
R83 GNDA.n2 GNDA.t22 48.0005
R84 GNDA.n2 GNDA.t17 48.0005
R85 GNDA.n6 GNDA.t1 48.0005
R86 GNDA.n6 GNDA.t9 48.0005
R87 GNDA.t24 GNDA.n1 236.792
R88 GNDA.n0 GNDA.n1 2.75546
R89 GNDA GNDA.n0 2.4755
R90 CLK.n3 CLK.n2 742.51
R91 CLK.n8 CLK.t1 723.534
R92 CLK.t2 CLK.n9 723.534
R93 CLK.n2 CLK.n1 684.806
R94 CLK.n7 CLK.n6 366.856
R95 CLK.n0 CLK.t6 337.401
R96 CLK.n0 CLK.t5 305.267
R97 CLK.n8 CLK.t0 254.333
R98 CLK.n4 CLK.n3 224.934
R99 CLK.n7 CLK.t9 190.123
R100 CLK.n9 CLK.n7 187.201
R101 CLK.n1 CLK.n0 176.733
R102 CLK.n5 CLK.n4 176.733
R103 CLK.n6 CLK.n5 176.733
R104 CLK.n3 CLK.t3 144.601
R105 CLK.n2 CLK.t10 131.976
R106 CLK.n0 CLK.t12 128.534
R107 CLK.n1 CLK.t8 128.534
R108 CLK.n4 CLK.t7 112.468
R109 CLK.n6 CLK.t11 112.468
R110 CLK.n5 CLK.t4 112.468
R111 CLK.n9 CLK.n8 70.4005
R112 D.n1 D.n0 701.467
R113 D.n1 D.t1 694.201
R114 D.n0 D.t3 321.334
R115 D.t0 D.n1 314.921
R116 D.n0 D.t2 144.601
R117 H.n0 H.t3 723.534
R118 H.n1 H.t4 553.534
R119 H.n0 H.t1 254.333
R120 H.n2 H.n1 206.333
R121 H.n1 H.n0 70.4005
R122 H.t2 H.n2 48.0005
R123 H.n2 H.t0 48.0005
R124 G.t0 G.t1 96.0005
R125 E.n0 E.t2 685.134
R126 E.n1 E.t0 663.801
R127 E.n0 E.t3 534.268
R128 E.t1 E.n1 362.921
R129 E.n1 E.n0 91.7338
R130 B.t0 B.t1 96.0005
R131 F.t0 F.t1 96.0005
C0 VIN VDDA 0.126677f
C1 VIN GNDA 0.291288f
C2 VDDA GNDA 2.83767f
.ends

