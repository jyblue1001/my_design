* PEX produced on Fri Aug  1 04:21:51 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_17.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_17 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t421 GNDA.t727 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 GNDA.t883 two_stage_opamp_dummy_magic_24_0.Vb1.t217 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 VDDA.t422 GNDA.t726 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 GNDA.t884 two_stage_opamp_dummy_magic_24_0.Vb1.t216 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 VDDA.t133 two_stage_opamp_dummy_magic_24_0.Vb3.t8 two_stage_opamp_dummy_magic_24_0.VD4.t31 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X5 VDDA.t423 GNDA.t725 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VOUT+.t19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 two_stage_opamp_dummy_magic_24_0.Vb2.t10 bgr_11_0.NFET_GATE_10uA.t5 GNDA.t146 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X8 two_stage_opamp_dummy_magic_24_0.Y.t9 two_stage_opamp_dummy_magic_24_0.Vb2.t11 two_stage_opamp_dummy_magic_24_0.VD4.t3 two_stage_opamp_dummy_magic_24_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X9 two_stage_opamp_dummy_magic_24_0.VD2.t20 two_stage_opamp_dummy_magic_24_0.Vb1.t228 two_stage_opamp_dummy_magic_24_0.Y.t13 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X10 GNDA.t885 two_stage_opamp_dummy_magic_24_0.Vb1.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 GNDA.t886 two_stage_opamp_dummy_magic_24_0.Vb1.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDDA.t424 GNDA.t724 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 VDDA.t425 GNDA.t723 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 VDDA.t365 VDDA.t362 VDDA.t364 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X15 VDDA.t426 GNDA.t722 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 VDDA.t420 bgr_11_0.1st_Vout_1.t7 bgr_11_0.V_TOP.t5 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X17 GNDA.t887 two_stage_opamp_dummy_magic_24_0.Vb1.t213 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 VDDA.t427 GNDA.t721 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VDDA.t428 GNDA.t720 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VOUT-.t19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VOUT+.t20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t81 bgr_11_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t8 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X23 VDDA.t429 GNDA.t719 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 GNDA.t888 two_stage_opamp_dummy_magic_24_0.Vb1.t212 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 VDDA.t430 GNDA.t718 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 GNDA.t889 two_stage_opamp_dummy_magic_24_0.Vb1.t211 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 VDDA.t431 GNDA.t717 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VDDA.t432 GNDA.t716 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VDDA.t433 GNDA.t715 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 VDDA.t361 VDDA.t359 two_stage_opamp_dummy_magic_24_0.VD3.t27 VDDA.t360 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X31 GNDA.t890 two_stage_opamp_dummy_magic_24_0.Vb1.t210 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 GNDA.t891 two_stage_opamp_dummy_magic_24_0.Vb1.t209 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VDDA.t434 GNDA.t714 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VDDA.t435 GNDA.t713 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 a_13430_3858.t1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t11 GNDA.t867 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X36 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t14 bgr_11_0.NFET_GATE_10uA.t6 GNDA.t161 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X37 bgr_11_0.1st_Vout_1.t8 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VDDA.t436 GNDA.t712 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VDDA.t437 GNDA.t711 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VDDA.t438 GNDA.t710 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 GNDA.t892 two_stage_opamp_dummy_magic_24_0.Vb1.t208 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT-.t20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VDDA.t439 GNDA.t709 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT-.t21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 GNDA.t743 GNDA.t845 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X46 bgr_11_0.V_TOP.t14 VDDA.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VOUT-.t22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VDDA.t440 GNDA.t708 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VDDA.t441 GNDA.t707 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VDDA.t442 GNDA.t706 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT-.t23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VDDA.t443 GNDA.t705 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VDDA.t444 GNDA.t704 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 GNDA.t844 GNDA.t842 bgr_11_0.NFET_GATE_10uA.t2 GNDA.t843 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X55 GNDA.t893 two_stage_opamp_dummy_magic_24_0.Vb1.t207 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 two_stage_opamp_dummy_magic_24_0.V_err_gate.t5 bgr_11_0.NFET_GATE_10uA.t7 GNDA.t163 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X57 two_stage_opamp_dummy_magic_24_0.Vb2_2.t5 two_stage_opamp_dummy_magic_24_0.Vb2_2.t3 two_stage_opamp_dummy_magic_24_0.Vb2_2.t5 two_stage_opamp_dummy_magic_24_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X58 VDDA.t445 GNDA.t703 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VDDA.t148 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.t12 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X60 VDDA.t446 GNDA.t702 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 two_stage_opamp_dummy_magic_24_0.V_source.t25 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t12 GNDA.t857 GNDA.t856 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X62 VDDA.t447 GNDA.t701 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 GNDA.t743 GNDA.t841 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X64 GNDA.t894 two_stage_opamp_dummy_magic_24_0.Vb1.t206 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 VDDA.t448 GNDA.t700 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VDDA.t449 GNDA.t699 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 two_stage_opamp_dummy_magic_24_0.Y.t8 two_stage_opamp_dummy_magic_24_0.Vb2.t12 two_stage_opamp_dummy_magic_24_0.VD4.t7 two_stage_opamp_dummy_magic_24_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X68 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t1 VDDA.t356 VDDA.t358 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X69 GNDA.t895 two_stage_opamp_dummy_magic_24_0.Vb1.t205 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VDDA.t416 bgr_11_0.1st_Vout_1.t9 bgr_11_0.V_TOP.t4 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X71 VDDA.t166 bgr_11_0.V_TOP.t15 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t3 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X72 VDDA.t450 GNDA.t698 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VDDA.t451 GNDA.t697 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 VOUT-.t24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 bgr_11_0.V_TOP.t16 VDDA.t167 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VDDA.t452 GNDA.t696 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VDDA.t453 GNDA.t695 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_11_0.V_TOP.t11 VDDA.t353 VDDA.t355 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X79 VDDA.t454 GNDA.t694 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VOUT+.t2 a_4380_346.t1 GNDA.t28 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X81 VDDA.t455 GNDA.t693 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 GNDA.t896 two_stage_opamp_dummy_magic_24_0.Vb1.t204 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VDDA.t456 GNDA.t692 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VDDA.t457 GNDA.t691 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 GNDA.t897 two_stage_opamp_dummy_magic_24_0.Vb1.t203 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT+.t9 two_stage_opamp_dummy_magic_24_0.Y.t25 VDDA.t244 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X87 VDDA.t458 GNDA.t690 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 bgr_11_0.V_TOP.t17 VDDA.t228 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VDDA.t459 GNDA.t689 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 VOUT-.t25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 GNDA.t130 two_stage_opamp_dummy_magic_24_0.X.t25 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t9 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X92 GNDA.t898 two_stage_opamp_dummy_magic_24_0.Vb1.t202 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 VOUT-.t26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 VOUT-.t27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 two_stage_opamp_dummy_magic_24_0.VD3.t37 two_stage_opamp_dummy_magic_24_0.Vb3.t9 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X96 VDDA.t460 GNDA.t688 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT-.t28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 bgr_11_0.PFET_GATE_10uA.t7 bgr_11_0.1st_Vout_2.t7 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X99 GNDA.t899 two_stage_opamp_dummy_magic_24_0.Vb1.t201 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 VDDA.t461 GNDA.t687 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 VOUT-.t29 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 VOUT+.t18 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t2 GNDA.t876 GNDA.t875 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X103 VOUT+.t21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VDDA.t462 GNDA.t686 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 GNDA.t743 GNDA.t840 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X106 VDDA.t463 GNDA.t685 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VDDA.t464 GNDA.t684 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 GNDA.t900 two_stage_opamp_dummy_magic_24_0.Vb1.t200 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VDDA.t465 GNDA.t683 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 VOUT+.t22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VDDA.t352 VDDA.t350 bgr_11_0.NFET_GATE_10uA.t1 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X112 VDDA.t13 two_stage_opamp_dummy_magic_24_0.X.t26 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t1 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X113 GNDA.t901 two_stage_opamp_dummy_magic_24_0.Vb1.t199 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 VDDA.t466 GNDA.t682 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VDDA.t20 bgr_11_0.V_mir1.t9 bgr_11_0.V_mir1.t10 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X116 two_stage_opamp_dummy_magic_24_0.V_source.t0 VIN-.t0 two_stage_opamp_dummy_magic_24_0.VD1.t9 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X117 VDDA.t467 GNDA.t681 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+.t23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 two_stage_opamp_dummy_magic_24_0.V_err_gate.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t4 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t3 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X120 GNDA.t859 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_24_0.V_source.t24 GNDA.t858 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X121 bgr_11_0.V_TOP.t18 VDDA.t229 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 GNDA.t902 two_stage_opamp_dummy_magic_24_0.Vb1.t198 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 GNDA.t903 two_stage_opamp_dummy_magic_24_0.Vb1.t197 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t5 VDDA.t347 VDDA.t349 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X125 VDDA.t468 GNDA.t680 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VDDA.t469 GNDA.t679 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VDDA.t470 GNDA.t678 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VDDA.t471 GNDA.t677 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 GNDA.t904 two_stage_opamp_dummy_magic_24_0.Vb1.t196 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 GNDA.t905 two_stage_opamp_dummy_magic_24_0.Vb1.t195 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 VDDA.t472 GNDA.t676 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT+.t24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT-.t30 two_stage_opamp_dummy_magic_24_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VDDA.t405 bgr_11_0.1st_Vout_2.t8 bgr_11_0.PFET_GATE_10uA.t9 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X135 VOUT+.t25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 two_stage_opamp_dummy_magic_24_0.VD2.t19 two_stage_opamp_dummy_magic_24_0.Vb1.t229 two_stage_opamp_dummy_magic_24_0.Y.t15 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X137 VDDA.t111 GNDA.t837 GNDA.t839 GNDA.t838 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X138 VDDA.t370 two_stage_opamp_dummy_magic_24_0.Y.t26 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t11 GNDA.t847 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X139 VDDA.t473 GNDA.t675 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VDDA.t371 two_stage_opamp_dummy_magic_24_0.Y.t27 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t10 GNDA.t848 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X141 GNDA.t906 two_stage_opamp_dummy_magic_24_0.Vb1.t194 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 bgr_11_0.START_UP.t5 bgr_11_0.V_TOP.t19 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X143 VDDA.t474 GNDA.t674 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT-.t31 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VDDA.t475 GNDA.t673 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 two_stage_opamp_dummy_magic_24_0.VD1.t8 VIN-.t1 two_stage_opamp_dummy_magic_24_0.V_source.t29 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X147 VDDA.t476 GNDA.t672 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VDDA.t477 GNDA.t671 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 bgr_11_0.V_TOP.t20 VDDA.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 GNDA.t907 two_stage_opamp_dummy_magic_24_0.Vb1.t193 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 GNDA.t908 two_stage_opamp_dummy_magic_24_0.Vb1.t192 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VDDA.t478 GNDA.t670 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT-.t32 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 two_stage_opamp_dummy_magic_24_0.err_amp_out.t3 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t5 GNDA.t869 GNDA.t868 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X155 bgr_11_0.1st_Vout_2.t9 bgr_11_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VDDA.t479 GNDA.t669 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VDDA.t480 GNDA.t668 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT-.t33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VOUT-.t34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 GNDA.t909 two_stage_opamp_dummy_magic_24_0.Vb1.t191 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VDDA.t481 GNDA.t667 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VDDA.t482 GNDA.t666 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VDDA.t483 GNDA.t665 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VDDA.t484 GNDA.t664 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT+.t26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+.t27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 two_stage_opamp_dummy_magic_24_0.VD2.t4 VIN+.t0 two_stage_opamp_dummy_magic_24_0.V_source.t7 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X168 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_24_0.X.t27 VDDA.t176 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X169 GNDA.t910 two_stage_opamp_dummy_magic_24_0.Vb1.t190 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VDDA.t485 GNDA.t663 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VOUT+.t28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 bgr_11_0.Vin+.t5 bgr_11_0.V_TOP.t21 VDDA.t194 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X173 VDDA.t42 bgr_11_0.V_mir2.t13 bgr_11_0.1st_Vout_2.t1 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X174 GNDA.t911 two_stage_opamp_dummy_magic_24_0.Vb1.t189 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VDDA.t486 GNDA.t662 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 bgr_11_0.V_mir1.t0 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t1 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X177 GNDA.t912 two_stage_opamp_dummy_magic_24_0.Vb1.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VDDA.t487 GNDA.t661 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 GNDA.t913 two_stage_opamp_dummy_magic_24_0.Vb1.t187 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VDDA.t488 GNDA.t660 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT-.t35 two_stage_opamp_dummy_magic_24_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VDDA.t489 GNDA.t659 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 VOUT-.t36 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 VDDA.t490 GNDA.t658 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 two_stage_opamp_dummy_magic_24_0.V_source.t23 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t14 GNDA.t860 GNDA.t813 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X186 bgr_11_0.1st_Vout_2.t10 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 VDDA.t491 GNDA.t657 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VDDA.t492 GNDA.t656 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 GNDA.t914 two_stage_opamp_dummy_magic_24_0.Vb1.t186 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 VOUT-.t37 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 VDDA.t493 GNDA.t655 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 GNDA.t873 a_11300_28850.t1 GNDA.t872 sky130_fd_pr__res_xhigh_po_0p35 l=6
X193 VDDA.t346 VDDA.t343 VDDA.t345 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X194 a_4100_3858.t1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t0 GNDA.t147 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X195 VDDA.t494 GNDA.t654 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT-.t38 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VOUT-.t17 a_13390_346.t1 GNDA.t871 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X198 GNDA.t915 two_stage_opamp_dummy_magic_24_0.Vb1.t185 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VDDA.t495 GNDA.t653 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 bgr_11_0.1st_Vout_1.t10 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 GNDA.t916 two_stage_opamp_dummy_magic_24_0.Vb1.t184 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VOUT-.t39 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VOUT-.t40 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 two_stage_opamp_dummy_magic_24_0.VD4.t21 VDDA.t340 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X206 VDDA.t496 GNDA.t652 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VDDA.t497 GNDA.t651 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VDDA.t498 GNDA.t650 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 bgr_11_0.V_TOP.t22 VDDA.t195 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT-.t41 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 GNDA.t836 GNDA.t834 two_stage_opamp_dummy_magic_24_0.V_source.t37 GNDA.t835 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X212 VDDA.t499 GNDA.t649 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t6 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X214 VOUT+.t7 two_stage_opamp_dummy_magic_24_0.Y.t28 VDDA.t205 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X215 VOUT-.t5 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t3 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X216 VDDA.t500 GNDA.t648 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 GNDA.t917 two_stage_opamp_dummy_magic_24_0.Vb1.t183 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VDDA.t501 GNDA.t647 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VOUT+.t29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 VOUT+.t30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 VOUT+.t31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VDDA.t502 GNDA.t646 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 bgr_11_0.V_mir2.t12 bgr_11_0.V_mir2.t11 VDDA.t170 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X224 VDDA.t65 bgr_11_0.V_TOP.t23 bgr_11_0.Vin-.t6 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X225 VDDA.t503 GNDA.t645 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VOUT+.t32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VOUT-.t42 two_stage_opamp_dummy_magic_24_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 GNDA.t0 two_stage_opamp_dummy_magic_24_0.X.t28 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t8 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X230 GNDA.t918 two_stage_opamp_dummy_magic_24_0.Vb1.t182 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 GNDA.t919 two_stage_opamp_dummy_magic_24_0.Vb1.t181 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VDDA.t504 GNDA.t644 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 GNDA.t920 two_stage_opamp_dummy_magic_24_0.Vb1.t180 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VDDA.t505 GNDA.t643 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDDA.t506 GNDA.t642 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 GNDA.t921 two_stage_opamp_dummy_magic_24_0.Vb1.t179 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 two_stage_opamp_dummy_magic_24_0.VD1.t21 two_stage_opamp_dummy_magic_24_0.Vb1.t230 two_stage_opamp_dummy_magic_24_0.X.t16 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X238 VOUT-.t43 two_stage_opamp_dummy_magic_24_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDDA.t372 two_stage_opamp_dummy_magic_24_0.X.t29 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t8 GNDA.t852 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X240 VDDA.t507 GNDA.t641 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VDDA.t508 GNDA.t640 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 two_stage_opamp_dummy_magic_24_0.VD4.t9 two_stage_opamp_dummy_magic_24_0.Vb2.t13 two_stage_opamp_dummy_magic_24_0.Y.t7 two_stage_opamp_dummy_magic_24_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X243 GNDA.t738 VDDA.t337 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X244 GNDA.t922 two_stage_opamp_dummy_magic_24_0.Vb1.t178 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT-.t44 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VDDA.t158 two_stage_opamp_dummy_magic_24_0.V_err_gate.t6 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t2 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X247 GNDA.t142 two_stage_opamp_dummy_magic_24_0.Y.t29 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t16 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X248 GNDA.t833 GNDA.t831 two_stage_opamp_dummy_magic_24_0.Vb1.t219 GNDA.t832 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X249 VDDA.t509 GNDA.t639 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 GNDA.t923 two_stage_opamp_dummy_magic_24_0.Vb1.t177 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VOUT-.t45 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 VOUT+.t34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 GNDA.t138 two_stage_opamp_dummy_magic_24_0.Y.t30 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t15 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X254 VDDA.t510 GNDA.t638 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VDDA.t511 GNDA.t637 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VDDA.t75 two_stage_opamp_dummy_magic_24_0.X.t30 VOUT-.t2 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X257 VDDA.t512 GNDA.t636 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VOUT+.t35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 two_stage_opamp_dummy_magic_24_0.VD2.t18 two_stage_opamp_dummy_magic_24_0.Vb1.t231 two_stage_opamp_dummy_magic_24_0.Y.t14 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X260 GNDA.t924 two_stage_opamp_dummy_magic_24_0.Vb1.t176 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 VDDA.t513 GNDA.t635 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VDDA.t336 VDDA.t334 VOUT-.t13 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X263 VDDA.t201 two_stage_opamp_dummy_magic_24_0.Y.t31 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t9 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X264 GNDA.t925 two_stage_opamp_dummy_magic_24_0.Vb1.t175 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 GNDA.t926 two_stage_opamp_dummy_magic_24_0.Vb1.t174 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT-.t46 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 two_stage_opamp_dummy_magic_24_0.VD1.t20 two_stage_opamp_dummy_magic_24_0.Vb1.t232 two_stage_opamp_dummy_magic_24_0.X.t15 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X268 bgr_11_0.1st_Vout_2.t12 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDDA.t514 GNDA.t634 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VDDA.t515 GNDA.t633 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 a_5700_30308.t0 a_5820_29044.t1 GNDA.t34 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X272 VDDA.t516 GNDA.t632 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 VOUT-.t47 two_stage_opamp_dummy_magic_24_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 VDDA.t15 bgr_11_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t3 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X275 bgr_11_0.V_TOP.t24 VDDA.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 VDDA.t517 GNDA.t631 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VDDA.t518 GNDA.t630 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t6 VDDA.t331 VDDA.t333 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X279 a_13550_3858.t1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t16 GNDA.t846 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X280 VDDA.t519 GNDA.t629 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 VDDA.t109 bgr_11_0.V_TOP.t25 bgr_11_0.Vin+.t4 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X282 GNDA.t927 two_stage_opamp_dummy_magic_24_0.Vb1.t173 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VOUT+.t36 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VOUT+.t37 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VOUT-.t48 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VDDA.t520 GNDA.t628 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VOUT+.t38 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 VOUT-.t49 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 VDDA.t521 GNDA.t627 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 VDDA.t522 GNDA.t626 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VDDA.t523 GNDA.t625 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 GNDA.t830 GNDA.t828 two_stage_opamp_dummy_magic_24_0.Vb3.t6 GNDA.t829 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X293 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_24_0.X.t31 GNDA.t123 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X294 VDDA.t524 GNDA.t624 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 GNDA.t928 two_stage_opamp_dummy_magic_24_0.Vb1.t172 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 VDDA.t525 GNDA.t623 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 VDDA.t526 GNDA.t622 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 GNDA.t929 two_stage_opamp_dummy_magic_24_0.Vb1.t171 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 VDDA.t527 GNDA.t621 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VDDA.t150 bgr_11_0.V_mir1.t13 bgr_11_0.1st_Vout_1.t3 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X301 two_stage_opamp_dummy_magic_24_0.VD2.t5 VIN+.t1 two_stage_opamp_dummy_magic_24_0.V_source.t28 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X302 GNDA.t930 two_stage_opamp_dummy_magic_24_0.Vb1.t170 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 VDDA.t528 GNDA.t620 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VDDA.t529 GNDA.t619 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 VDDA.t530 GNDA.t618 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 VDDA.t531 GNDA.t617 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 two_stage_opamp_dummy_magic_24_0.VD2.t8 VIN+.t2 two_stage_opamp_dummy_magic_24_0.V_source.t36 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X308 two_stage_opamp_dummy_magic_24_0.V_p_mir.t3 VIN+.t3 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t0 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X309 GNDA.t931 two_stage_opamp_dummy_magic_24_0.Vb1.t169 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VDDA.t532 GNDA.t616 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT-.t50 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VDDA.t533 GNDA.t615 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 VOUT+.t39 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VOUT+.t40 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 bgr_11_0.V_p_2.t0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t7 bgr_11_0.V_mir2.t0 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X316 VDDA.t534 GNDA.t614 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VOUT-.t51 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 two_stage_opamp_dummy_magic_24_0.VD4.t37 two_stage_opamp_dummy_magic_24_0.VD4.t35 two_stage_opamp_dummy_magic_24_0.Y.t24 two_stage_opamp_dummy_magic_24_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X319 VOUT-.t52 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT-.t53 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 two_stage_opamp_dummy_magic_24_0.V_p_mir.t2 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t15 GNDA.t862 GNDA.t861 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X322 VDDA.t535 GNDA.t613 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VOUT-.t54 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 VOUT+.t41 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 two_stage_opamp_dummy_magic_24_0.V_source.t22 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t16 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X326 VDDA.t536 GNDA.t612 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VDDA.t537 GNDA.t611 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VDDA.t538 GNDA.t610 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VDDA.t539 GNDA.t609 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VDDA.t540 GNDA.t608 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 bgr_11_0.V_TOP.t26 VDDA.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 VDDA.t541 GNDA.t607 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VOUT+.t42 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VDDA.t542 GNDA.t606 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 VDDA.t543 GNDA.t605 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 VOUT-.t55 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 bgr_11_0.Vin+.t3 bgr_11_0.V_TOP.t27 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X338 VDDA.t544 GNDA.t604 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 GNDA.t932 two_stage_opamp_dummy_magic_24_0.Vb1.t168 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VDDA.t545 GNDA.t603 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VOUT+.t43 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VDDA.t546 GNDA.t602 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VOUT+.t44 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 VOUT+.t45 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 bgr_11_0.1st_Vout_2.t2 bgr_11_0.V_mir2.t14 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X346 VDDA.t547 GNDA.t601 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VDDA.t548 GNDA.t600 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT+.t46 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT+.t47 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VDDA.t418 bgr_11_0.1st_Vout_1.t11 bgr_11_0.V_TOP.t3 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X351 GNDA.t933 two_stage_opamp_dummy_magic_24_0.Vb1.t167 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 VDDA.t549 GNDA.t599 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 VDDA.t330 VDDA.t328 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X354 VDDA.t44 bgr_11_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t7 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X355 VDDA.t550 GNDA.t598 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 bgr_11_0.cap_res2.t0 bgr_11_0.PFET_GATE_10uA.t1 GNDA.t65 sky130_fd_pr__res_high_po_0p35 l=2.05
X357 VDDA.t223 bgr_11_0.V_mir1.t14 bgr_11_0.1st_Vout_1.t4 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X358 VDDA.t551 GNDA.t597 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 GNDA.t934 two_stage_opamp_dummy_magic_24_0.Vb1.t166 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 VDDA.t552 GNDA.t596 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 VDDA.t553 GNDA.t595 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 GNDA.t935 two_stage_opamp_dummy_magic_24_0.Vb1.t165 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 GNDA.t159 two_stage_opamp_dummy_magic_24_0.X.t32 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t6 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X364 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 VDDA.t554 GNDA.t594 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 VOUT-.t56 two_stage_opamp_dummy_magic_24_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 GNDA.t936 two_stage_opamp_dummy_magic_24_0.Vb1.t164 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 VOUT-.t57 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 VOUT-.t58 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 VOUT-.t59 two_stage_opamp_dummy_magic_24_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT-.t60 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 GNDA.t827 GNDA.t825 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t1 GNDA.t826 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X373 VDDA.t555 GNDA.t593 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 VDDA.t556 GNDA.t592 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VDDA.t557 GNDA.t591 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 GNDA.t743 GNDA.t742 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X377 two_stage_opamp_dummy_magic_24_0.VD1.t19 two_stage_opamp_dummy_magic_24_0.Vb1.t233 two_stage_opamp_dummy_magic_24_0.X.t18 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X378 two_stage_opamp_dummy_magic_24_0.X.t12 two_stage_opamp_dummy_magic_24_0.Vb2.t14 two_stage_opamp_dummy_magic_24_0.VD3.t25 two_stage_opamp_dummy_magic_24_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X379 VOUT+.t48 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VDDA.t558 GNDA.t590 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t13 bgr_11_0.PFET_GATE_10uA.t13 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X382 GNDA.t135 two_stage_opamp_dummy_magic_24_0.Y.t32 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t14 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X383 GNDA.t937 two_stage_opamp_dummy_magic_24_0.Vb1.t163 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 VOUT+.t49 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 GNDA.t880 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t14 GNDA.t879 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X386 VDDA.t559 GNDA.t589 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VOUT+.t50 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VDDA.t560 GNDA.t588 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 GNDA.t938 two_stage_opamp_dummy_magic_24_0.Vb1.t162 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VDDA.t561 GNDA.t587 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 VDDA.t562 GNDA.t586 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VDDA.t382 two_stage_opamp_dummy_magic_24_0.X.t33 VOUT-.t16 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X393 VDDA.t563 GNDA.t585 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 GNDA.t939 two_stage_opamp_dummy_magic_24_0.Vb1.t161 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 VOUT+.t51 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 a_6350_30458.t1 a_6470_28850.t1 GNDA.t51 sky130_fd_pr__res_xhigh_po_0p35 l=6
X397 two_stage_opamp_dummy_magic_24_0.VD2.t17 two_stage_opamp_dummy_magic_24_0.Vb1.t234 two_stage_opamp_dummy_magic_24_0.Y.t17 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X398 VDDA.t199 two_stage_opamp_dummy_magic_24_0.Y.t33 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t8 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X399 VDDA.t564 GNDA.t584 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT-.t61 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VDDA.t565 GNDA.t583 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VOUT+.t52 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 two_stage_opamp_dummy_magic_24_0.VD1.t18 two_stage_opamp_dummy_magic_24_0.Vb1.t235 two_stage_opamp_dummy_magic_24_0.X.t17 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X404 VDDA.t566 GNDA.t582 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 GNDA.t940 two_stage_opamp_dummy_magic_24_0.Vb1.t160 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VDDA.t567 GNDA.t581 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VOUT+.t53 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 GNDA.t941 two_stage_opamp_dummy_magic_24_0.Vb1.t159 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VDDA.t568 GNDA.t580 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VDDA.t569 GNDA.t579 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 GNDA.t942 two_stage_opamp_dummy_magic_24_0.Vb1.t158 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 GNDA.t943 two_stage_opamp_dummy_magic_24_0.Vb1.t157 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VDDA.t570 GNDA.t578 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VDDA.t571 GNDA.t577 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT-.t62 two_stage_opamp_dummy_magic_24_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 bgr_11_0.V_mir2.t10 bgr_11_0.V_mir2.t9 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X418 VOUT-.t63 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 two_stage_opamp_dummy_magic_24_0.Vb1_2.t4 two_stage_opamp_dummy_magic_24_0.Vb1.t224 two_stage_opamp_dummy_magic_24_0.Vb1.t225 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X420 GNDA.t944 two_stage_opamp_dummy_magic_24_0.Vb1.t156 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT-.t64 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VOUT-.t65 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 two_stage_opamp_dummy_magic_24_0.VD2.t7 VIN+.t4 two_stage_opamp_dummy_magic_24_0.V_source.t35 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X424 GNDA.t824 GNDA.t822 VOUT+.t15 GNDA.t823 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X425 VDDA.t572 GNDA.t576 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VDDA.t573 GNDA.t575 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VDDA.t574 GNDA.t574 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VDDA.t575 GNDA.t573 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VDDA.t576 GNDA.t572 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 GNDA.t945 two_stage_opamp_dummy_magic_24_0.Vb1.t155 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 GNDA.t946 two_stage_opamp_dummy_magic_24_0.Vb1.t154 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VDDA.t577 GNDA.t571 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 GNDA.t947 two_stage_opamp_dummy_magic_24_0.Vb1.t153 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VDDA.t578 GNDA.t570 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT+.t54 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 GNDA.t948 two_stage_opamp_dummy_magic_24_0.Vb1.t152 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 two_stage_opamp_dummy_magic_24_0.cap_res_X.t0 two_stage_opamp_dummy_magic_24_0.X.t0 GNDA.t29 sky130_fd_pr__res_high_po_1p41 l=1.41
X438 GNDA.t949 two_stage_opamp_dummy_magic_24_0.Vb1.t151 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 GNDA.t950 two_stage_opamp_dummy_magic_24_0.Vb1.t150 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VDDA.t579 GNDA.t569 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 GNDA.t743 GNDA.t821 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X442 a_12070_30308.t0 a_11950_29100.t0 GNDA.t5 sky130_fd_pr__res_xhigh_po_0p35 l=4
X443 two_stage_opamp_dummy_magic_24_0.V_source.t21 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t17 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X444 VDDA.t580 GNDA.t568 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VDDA.t581 GNDA.t567 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 VDDA.t582 GNDA.t566 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 GNDA.t951 two_stage_opamp_dummy_magic_24_0.Vb1.t149 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 bgr_11_0.1st_Vout_1.t13 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VDDA.t583 GNDA.t565 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 VOUT+.t55 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 VDDA.t584 GNDA.t564 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 VDDA.t585 GNDA.t563 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT-.t66 two_stage_opamp_dummy_magic_24_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VDDA.t144 two_stage_opamp_dummy_magic_24_0.Vb3.t10 two_stage_opamp_dummy_magic_24_0.VD4.t30 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X455 VDDA.t586 GNDA.t562 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 bgr_11_0.V_TOP.t28 VDDA.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 GNDA.t952 two_stage_opamp_dummy_magic_24_0.Vb1.t148 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 two_stage_opamp_dummy_magic_24_0.Vb3.t7 bgr_11_0.NFET_GATE_10uA.t9 GNDA.t882 GNDA.t881 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X459 bgr_11_0.PFET_GATE_10uA.t8 bgr_11_0.1st_Vout_2.t14 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X460 two_stage_opamp_dummy_magic_24_0.Vb3.t4 two_stage_opamp_dummy_magic_24_0.Vb2.t15 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X461 VDDA.t587 GNDA.t561 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 GNDA.t953 two_stage_opamp_dummy_magic_24_0.Vb1.t147 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 VDDA.t588 GNDA.t560 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 VDDA.t589 GNDA.t559 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 GNDA.t95 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t3 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t4 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X466 VDDA.t590 GNDA.t558 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 VDDA.t591 GNDA.t557 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VDDA.t592 GNDA.t556 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VDDA.t593 GNDA.t555 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 GNDA.t954 two_stage_opamp_dummy_magic_24_0.Vb1.t146 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT-.t67 two_stage_opamp_dummy_magic_24_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VDDA.t594 GNDA.t554 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VDDA.t595 GNDA.t553 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VOUT-.t68 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VDDA.t146 two_stage_opamp_dummy_magic_24_0.Vb3.t11 two_stage_opamp_dummy_magic_24_0.VD3.t36 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X477 VDDA.t596 GNDA.t552 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VOUT+.t56 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VDDA.t597 GNDA.t551 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VOUT-.t69 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VDDA.t598 GNDA.t550 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT+.t57 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 GNDA.t955 two_stage_opamp_dummy_magic_24_0.Vb1.t145 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT+.t58 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT+.t59 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 two_stage_opamp_dummy_magic_24_0.Y.t6 two_stage_opamp_dummy_magic_24_0.Vb2.t16 two_stage_opamp_dummy_magic_24_0.VD4.t1 two_stage_opamp_dummy_magic_24_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X487 VDDA.t599 GNDA.t549 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VOUT+.t60 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 VDDA.t600 GNDA.t548 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VDDA.t601 GNDA.t547 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 GNDA.t956 two_stage_opamp_dummy_magic_24_0.Vb1.t144 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VDDA.t602 GNDA.t546 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t13 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X494 VDDA.t603 GNDA.t545 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 GNDA.t133 two_stage_opamp_dummy_magic_24_0.Y.t34 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t13 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X496 VDDA.t604 GNDA.t544 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VDDA.t327 VDDA.t325 two_stage_opamp_dummy_magic_24_0.err_amp_out.t1 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X498 VDDA.t605 GNDA.t543 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VDDA.t606 GNDA.t542 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 VOUT+.t61 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VDDA.t607 GNDA.t541 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 GNDA.t180 bgr_11_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t12 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X503 bgr_11_0.V_TOP.t29 VDDA.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 VDDA.t608 GNDA.t540 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 VDDA.t48 bgr_11_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t6 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X506 GNDA.t957 two_stage_opamp_dummy_magic_24_0.Vb1.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 VDDA.t399 two_stage_opamp_dummy_magic_24_0.X.t34 VOUT-.t18 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X508 a_13550_3858.t0 two_stage_opamp_dummy_magic_24_0.V_tot.t1 GNDA.t52 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X509 VDDA.t609 GNDA.t539 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VDDA.t182 two_stage_opamp_dummy_magic_24_0.Y.t35 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t7 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X511 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t5 bgr_11_0.PFET_GATE_10uA.t15 VDDA.t83 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X512 VOUT-.t6 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t4 GNDA.t108 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X513 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 VDDA.t610 GNDA.t538 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VDDA.t611 GNDA.t537 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 two_stage_opamp_dummy_magic_24_0.VD1.t17 two_stage_opamp_dummy_magic_24_0.Vb1.t236 two_stage_opamp_dummy_magic_24_0.X.t23 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X517 GNDA.t958 two_stage_opamp_dummy_magic_24_0.Vb1.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VDDA.t612 GNDA.t536 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 GNDA.t959 two_stage_opamp_dummy_magic_24_0.Vb1.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VDDA.t613 GNDA.t535 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 bgr_11_0.V_TOP.t30 VDDA.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VDDA.t614 GNDA.t534 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VDDA.t615 GNDA.t533 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 bgr_11_0.START_UP.t4 bgr_11_0.V_TOP.t31 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X525 VDDA.t179 two_stage_opamp_dummy_magic_24_0.Y.t36 VOUT+.t6 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X526 GNDA.t960 two_stage_opamp_dummy_magic_24_0.Vb1.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 VOUT-.t70 two_stage_opamp_dummy_magic_24_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VDDA.t616 GNDA.t532 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 VDDA.t617 GNDA.t531 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT-.t71 two_stage_opamp_dummy_magic_24_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VDDA.t618 GNDA.t530 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 two_stage_opamp_dummy_magic_24_0.Vb2.t9 bgr_11_0.NFET_GATE_10uA.t12 GNDA.t169 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X533 bgr_11_0.1st_Vout_2.t3 bgr_11_0.V_mir2.t15 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X534 VDDA.t324 VDDA.t322 VOUT+.t13 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X535 VDDA.t619 GNDA.t529 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 GNDA.t961 two_stage_opamp_dummy_magic_24_0.Vb1.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 GNDA.t962 two_stage_opamp_dummy_magic_24_0.Vb1.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VDDA.t620 GNDA.t528 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 GNDA.t171 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_24_0.Vb2.t8 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X540 VOUT+.t62 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VOUT+.t63 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 two_stage_opamp_dummy_magic_24_0.VD2.t6 VIN+.t5 two_stage_opamp_dummy_magic_24_0.V_source.t32 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X543 GNDA.t963 two_stage_opamp_dummy_magic_24_0.Vb1.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VDDA.t621 GNDA.t527 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_24_0.X.t35 VDDA.t156 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X546 VDDA.t622 GNDA.t526 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 two_stage_opamp_dummy_magic_24_0.X.t22 two_stage_opamp_dummy_magic_24_0.Vb1.t237 two_stage_opamp_dummy_magic_24_0.VD1.t16 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X548 VDDA.t623 GNDA.t525 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 GNDA.t964 two_stage_opamp_dummy_magic_24_0.Vb1.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VDDA.t624 GNDA.t524 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VDDA.t625 GNDA.t523 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 bgr_11_0.NFET_GATE_10uA.t4 bgr_11_0.NFET_GATE_10uA.t3 GNDA.t182 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X553 GNDA.t820 GNDA.t818 VDDA.t378 GNDA.t819 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X554 VDDA.t626 GNDA.t522 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VDDA.t627 GNDA.t521 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VDDA.t628 GNDA.t520 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 bgr_11_0.V_TOP.t32 VDDA.t190 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 bgr_11_0.1st_Vout_2.t15 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VDDA.t629 GNDA.t519 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VOUT-.t72 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 two_stage_opamp_dummy_magic_24_0.V_source.t20 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t18 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X562 VOUT-.t4 two_stage_opamp_dummy_magic_24_0.X.t36 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X563 VDDA.t630 GNDA.t518 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 GNDA.t965 two_stage_opamp_dummy_magic_24_0.Vb1.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 bgr_11_0.V_mir1.t8 bgr_11_0.V_mir1.t7 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X566 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t9 VDDA.t319 VDDA.t321 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X567 two_stage_opamp_dummy_magic_24_0.Y.t16 two_stage_opamp_dummy_magic_24_0.Vb1.t238 two_stage_opamp_dummy_magic_24_0.VD2.t16 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X568 VDDA.t631 GNDA.t517 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT-.t73 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 GNDA.t966 two_stage_opamp_dummy_magic_24_0.Vb1.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 VDDA.t632 GNDA.t516 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 GNDA.t967 two_stage_opamp_dummy_magic_24_0.Vb1.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 bgr_11_0.V_TOP.t6 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t2 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X574 two_stage_opamp_dummy_magic_24_0.Vb1_2.t3 two_stage_opamp_dummy_magic_24_0.Vb1.t222 two_stage_opamp_dummy_magic_24_0.Vb1.t223 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X575 VDDA.t633 GNDA.t515 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 VDDA.t634 GNDA.t514 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VDDA.t318 VDDA.t316 bgr_11_0.V_TOP.t10 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X579 VDDA.t635 GNDA.t513 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 VOUT-.t74 two_stage_opamp_dummy_magic_24_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 GNDA.t968 two_stage_opamp_dummy_magic_24_0.Vb1.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 VDDA.t636 GNDA.t512 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 two_stage_opamp_dummy_magic_24_0.X.t2 two_stage_opamp_dummy_magic_24_0.VD3.t3 two_stage_opamp_dummy_magic_24_0.VD3.t5 two_stage_opamp_dummy_magic_24_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X584 VDDA.t637 GNDA.t511 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 VOUT+.t64 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 VOUT-.t75 two_stage_opamp_dummy_magic_24_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 VDDA.t638 GNDA.t510 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 bgr_11_0.1st_Vout_2.t16 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 VOUT+.t65 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 GNDA.t969 two_stage_opamp_dummy_magic_24_0.Vb1.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 VDDA.t639 GNDA.t509 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 VDDA.t640 GNDA.t508 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 VOUT+.t66 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VOUT+.t67 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 VDDA.t641 GNDA.t507 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 two_stage_opamp_dummy_magic_24_0.VD3.t23 two_stage_opamp_dummy_magic_24_0.Vb2.t17 two_stage_opamp_dummy_magic_24_0.X.t11 two_stage_opamp_dummy_magic_24_0.VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X597 GNDA.t970 two_stage_opamp_dummy_magic_24_0.Vb1.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 GNDA.t971 two_stage_opamp_dummy_magic_24_0.Vb1.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 VDDA.t642 GNDA.t506 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 VDDA.t643 GNDA.t505 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 GNDA.t972 two_stage_opamp_dummy_magic_24_0.Vb1.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VDDA.t644 GNDA.t504 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 GNDA.t973 two_stage_opamp_dummy_magic_24_0.Vb1.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VDDA.t645 GNDA.t503 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 bgr_11_0.1st_Vout_1.t17 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 VDDA.t646 GNDA.t502 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 bgr_11_0.NFET_GATE_10uA.t0 bgr_11_0.PFET_GATE_10uA.t16 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X608 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 GNDA.t46 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_24_0.V_source.t19 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X610 GNDA.t7 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_24_0.V_source.t18 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X611 GNDA.t974 two_stage_opamp_dummy_magic_24_0.Vb1.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VDDA.t647 GNDA.t501 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VDDA.t648 GNDA.t500 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 VOUT+.t68 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 two_stage_opamp_dummy_magic_24_0.V_err_p.t2 two_stage_opamp_dummy_magic_24_0.V_err_gate.t7 VDDA.t401 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X616 GNDA.t132 two_stage_opamp_dummy_magic_24_0.Y.t37 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t12 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X617 VDDA.t649 GNDA.t499 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 VDDA.t650 GNDA.t498 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 GNDA.t975 two_stage_opamp_dummy_magic_24_0.Vb1.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VOUT-.t76 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 VDDA.t60 bgr_11_0.V_TOP.t33 bgr_11_0.Vin+.t2 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X622 VDDA.t651 GNDA.t497 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 VDDA.t68 two_stage_opamp_dummy_magic_24_0.X.t37 VOUT-.t1 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X625 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 GNDA.t976 two_stage_opamp_dummy_magic_24_0.Vb1.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 VOUT-.t77 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 VDDA.t652 GNDA.t496 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 VDDA.t653 GNDA.t495 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 VDDA.t654 GNDA.t494 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 bgr_11_0.PFET_GATE_10uA.t2 bgr_11_0.1st_Vout_2.t19 VDDA.t140 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X632 GNDA.t977 two_stage_opamp_dummy_magic_24_0.Vb1.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 VDDA.t655 GNDA.t493 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 VOUT-.t78 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VOUT-.t79 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 two_stage_opamp_dummy_magic_24_0.VD1.t7 VIN-.t2 two_stage_opamp_dummy_magic_24_0.V_source.t5 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X637 VDDA.t656 GNDA.t492 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VDDA.t657 GNDA.t491 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 VOUT-.t80 two_stage_opamp_dummy_magic_24_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 VOUT+.t69 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 VOUT-.t81 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 two_stage_opamp_dummy_magic_24_0.VD3.t26 VDDA.t313 VDDA.t315 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X643 GNDA.t978 two_stage_opamp_dummy_magic_24_0.Vb1.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 VDDA.t658 GNDA.t490 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 VDDA.t246 two_stage_opamp_dummy_magic_24_0.Y.t38 VOUT+.t10 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X646 VDDA.t659 GNDA.t489 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 VOUT+.t70 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 GNDA.t979 two_stage_opamp_dummy_magic_24_0.Vb1.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 VDDA.t660 GNDA.t488 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_24_0.X.t38 GNDA.t53 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X651 VDDA.t661 GNDA.t487 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 VDDA.t662 GNDA.t486 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 GNDA.t980 two_stage_opamp_dummy_magic_24_0.Vb1.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 GNDA.t981 two_stage_opamp_dummy_magic_24_0.Vb1.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 VDDA.t663 GNDA.t485 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 GNDA.t982 two_stage_opamp_dummy_magic_24_0.Vb1.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VDDA.t312 VDDA.t310 GNDA.t737 VDDA.t311 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X658 bgr_11_0.1st_Vout_2.t20 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VDDA.t664 GNDA.t484 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 VDDA.t665 GNDA.t483 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 two_stage_opamp_dummy_magic_24_0.VD2.t10 GNDA.t815 GNDA.t817 GNDA.t816 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X662 GNDA.t983 two_stage_opamp_dummy_magic_24_0.Vb1.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t2 bgr_11_0.V_TOP.t34 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X664 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_24_0.X.t39 VDDA.t115 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X665 VDDA.t666 GNDA.t736 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 VOUT+.t71 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 VOUT+.t72 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 GNDA.t814 GNDA.t812 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t11 GNDA.t813 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X669 two_stage_opamp_dummy_magic_24_0.VD1.t6 VIN-.t3 two_stage_opamp_dummy_magic_24_0.V_source.t26 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X670 GNDA.t984 two_stage_opamp_dummy_magic_24_0.Vb1.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 VOUT-.t82 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 VOUT+.t73 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 VDDA.t667 GNDA.t735 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VOUT-.t83 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 VOUT-.t84 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 VDDA.t668 GNDA.t734 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 VOUT+.t74 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 two_stage_opamp_dummy_magic_24_0.VD4.t29 two_stage_opamp_dummy_magic_24_0.Vb3.t12 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X679 GNDA.t985 two_stage_opamp_dummy_magic_24_0.Vb1.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 VDDA.t669 GNDA.t733 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 bgr_11_0.1st_Vout_2.t5 bgr_11_0.V_mir2.t16 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X682 two_stage_opamp_dummy_magic_24_0.V_source.t17 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t21 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X683 bgr_11_0.1st_Vout_1.t19 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 GNDA.t986 two_stage_opamp_dummy_magic_24_0.Vb1.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VOUT-.t85 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 bgr_11_0.V_TOP.t2 bgr_11_0.1st_Vout_1.t20 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X687 two_stage_opamp_dummy_magic_24_0.Y.t19 two_stage_opamp_dummy_magic_24_0.Vb1.t239 two_stage_opamp_dummy_magic_24_0.VD2.t15 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X688 VDDA.t670 GNDA.t732 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VDDA.t671 GNDA.t731 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 VDDA.t672 GNDA.t730 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 GNDA.t729 VDDA.t673 bgr_11_0.V_TOP.t12 GNDA.t728 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X692 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_24_0.Vb3.t2 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X693 VOUT-.t3 two_stage_opamp_dummy_magic_24_0.X.t40 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X694 VDDA.t674 GNDA.t482 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 VDDA.t675 GNDA.t481 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 VDDA.t309 VDDA.t307 two_stage_opamp_dummy_magic_24_0.Vb1.t1 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X697 two_stage_opamp_dummy_magic_24_0.Y.t18 two_stage_opamp_dummy_magic_24_0.Vb1.t240 two_stage_opamp_dummy_magic_24_0.VD2.t14 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X698 bgr_11_0.V_TOP.t35 VDDA.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 VDDA.t676 GNDA.t480 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X700 VDDA.t677 GNDA.t479 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 VDDA.t678 GNDA.t478 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 VOUT-.t86 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 VOUT-.t87 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 two_stage_opamp_dummy_magic_24_0.VD3.t21 two_stage_opamp_dummy_magic_24_0.Vb2.t18 two_stage_opamp_dummy_magic_24_0.X.t10 two_stage_opamp_dummy_magic_24_0.VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X705 VDDA.t679 GNDA.t477 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 GNDA.t987 two_stage_opamp_dummy_magic_24_0.Vb1.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 GNDA.t988 two_stage_opamp_dummy_magic_24_0.Vb1.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT+.t75 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VOUT+.t76 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 VOUT-.t88 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 bgr_11_0.1st_Vout_1.t5 bgr_11_0.V_mir1.t15 VDDA.t225 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X712 VDDA.t680 GNDA.t476 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 VDDA.t681 GNDA.t475 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 VOUT+.t77 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VOUT+.t78 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 two_stage_opamp_dummy_magic_24_0.VD3.t35 two_stage_opamp_dummy_magic_24_0.Vb3.t13 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X717 GNDA.t854 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t5 VOUT+.t17 GNDA.t853 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X718 GNDA.t989 two_stage_opamp_dummy_magic_24_0.Vb1.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 GNDA.t990 two_stage_opamp_dummy_magic_24_0.Vb1.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 GNDA.t991 two_stage_opamp_dummy_magic_24_0.Vb1.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VOUT+.t79 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 VDDA.t682 GNDA.t474 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 VDDA.t683 GNDA.t473 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VDDA.t684 GNDA.t472 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VDDA.t685 GNDA.t471 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 bgr_11_0.V_p_1.t2 VDDA.t686 GNDA.t470 GNDA.t469 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X727 VDDA.t11 bgr_11_0.V_TOP.t36 bgr_11_0.START_UP.t3 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X728 VDDA.t687 GNDA.t444 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 GNDA.t811 GNDA.t808 GNDA.t810 GNDA.t809 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X730 VDDA.t688 GNDA.t443 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 GNDA.t992 two_stage_opamp_dummy_magic_24_0.Vb1.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 VOUT-.t89 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 GNDA.t743 GNDA.t744 bgr_11_0.Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X734 bgr_11_0.Vin-.t5 bgr_11_0.V_TOP.t37 VDDA.t212 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X735 VDDA.t689 GNDA.t442 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 VOUT-.t90 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VOUT-.t91 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 VDDA.t690 GNDA.t441 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 VDDA.t691 GNDA.t440 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 VOUT-.t92 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 VOUT+.t80 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 VDDA.t306 VDDA.t304 bgr_11_0.PFET_GATE_10uA.t5 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X743 VDDA.t692 GNDA.t439 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 VOUT+.t81 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 GNDA.t993 two_stage_opamp_dummy_magic_24_0.Vb1.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 VOUT-.t93 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VDDA.t693 GNDA.t438 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_24_0.VD4.t28 two_stage_opamp_dummy_magic_24_0.Vb3.t14 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X749 two_stage_opamp_dummy_magic_24_0.V_err_gate.t3 VDDA.t301 VDDA.t303 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X750 a_13430_3858.t0 two_stage_opamp_dummy_magic_24_0.V_tot.t2 GNDA.t102 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X751 VDDA.t694 GNDA.t437 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 GNDA.t155 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_24_0.V_source.t16 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X753 VDDA.t695 GNDA.t436 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VOUT+.t82 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 two_stage_opamp_dummy_magic_24_0.V_err_p.t3 two_stage_opamp_dummy_magic_24_0.V_tot.t5 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X756 VDDA.t696 GNDA.t435 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 GNDA.t994 two_stage_opamp_dummy_magic_24_0.Vb1.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VDDA.t697 GNDA.t434 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 VOUT+.t83 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VDDA.t698 GNDA.t433 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 VOUT-.t94 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 two_stage_opamp_dummy_magic_24_0.V_source.t38 two_stage_opamp_dummy_magic_24_0.Vb1.t241 two_stage_opamp_dummy_magic_24_0.Vb1_2.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X763 VDDA.t699 GNDA.t432 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 VDDA.t700 GNDA.t431 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VOUT+.t84 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 bgr_11_0.V_mir2.t8 bgr_11_0.V_mir2.t7 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X767 bgr_11_0.V_TOP.t38 VDDA.t213 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 GNDA.t995 two_stage_opamp_dummy_magic_24_0.Vb1.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 VDDA.t701 GNDA.t430 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 VDDA.t702 GNDA.t429 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 VDDA.t300 VDDA.t298 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t5 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X772 VDDA.t703 GNDA.t428 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X773 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t2 bgr_11_0.PFET_GATE_10uA.t17 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X774 GNDA.t996 two_stage_opamp_dummy_magic_24_0.Vb1.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 VDDA.t704 GNDA.t427 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_24_0.Y.t10 GNDA.t131 sky130_fd_pr__res_high_po_1p41 l=1.41
X777 VOUT+.t85 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 VDDA.t705 GNDA.t426 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 two_stage_opamp_dummy_magic_24_0.VD1.t5 VIN-.t4 two_stage_opamp_dummy_magic_24_0.V_source.t2 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X780 GNDA.t997 two_stage_opamp_dummy_magic_24_0.Vb1.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 VDDA.t706 GNDA.t425 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 VOUT+.t14 GNDA.t805 GNDA.t807 GNDA.t806 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X783 VDDA.t707 GNDA.t424 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 GNDA.t998 two_stage_opamp_dummy_magic_24_0.Vb1.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 VDDA.t248 two_stage_opamp_dummy_magic_24_0.Y.t39 VOUT+.t11 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X786 VDDA.t708 GNDA.t423 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 two_stage_opamp_dummy_magic_24_0.Vb3.t3 bgr_11_0.NFET_GATE_10uA.t14 GNDA.t173 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X788 VOUT-.t95 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X789 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_24_0.X.t41 GNDA.t87 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X790 VDDA.t709 GNDA.t422 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 VOUT-.t96 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X792 VDDA.t710 GNDA.t421 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 VOUT-.t97 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X794 GNDA.t999 two_stage_opamp_dummy_magic_24_0.Vb1.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X795 VDDA.t711 GNDA.t420 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 VOUT+.t86 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X797 GNDA.t1000 two_stage_opamp_dummy_magic_24_0.Vb1.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X798 VDDA.t712 GNDA.t419 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X799 VDDA.t713 GNDA.t418 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X800 bgr_11_0.1st_Vout_1.t1 bgr_11_0.V_mir1.t16 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X801 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_24_0.X.t42 VDDA.t119 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X802 GNDA.t1001 two_stage_opamp_dummy_magic_24_0.Vb1.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X803 VDDA.t714 GNDA.t417 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X804 VOUT+.t87 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X805 two_stage_opamp_dummy_magic_24_0.VD1.t4 VIN-.t5 two_stage_opamp_dummy_magic_24_0.V_source.t31 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X806 VOUT+.t88 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X807 VDDA.t297 VDDA.t295 two_stage_opamp_dummy_magic_24_0.V_err_gate.t2 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X808 VDDA.t715 GNDA.t416 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X809 VDDA.t29 two_stage_opamp_dummy_magic_24_0.Vb3.t15 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t10 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X810 VDDA.t716 GNDA.t415 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X811 VDDA.t717 GNDA.t414 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 VDDA.t718 GNDA.t413 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X813 GNDA.t1002 two_stage_opamp_dummy_magic_24_0.Vb1.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X814 VDDA.t719 GNDA.t412 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X815 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X816 VOUT-.t98 two_stage_opamp_dummy_magic_24_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X817 two_stage_opamp_dummy_magic_24_0.Y.t22 two_stage_opamp_dummy_magic_24_0.Vb1.t242 two_stage_opamp_dummy_magic_24_0.VD2.t13 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X818 VDDA.t720 GNDA.t411 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X819 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_24_0.Y.t40 VDDA.t171 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X820 GNDA.t1003 two_stage_opamp_dummy_magic_24_0.Vb1.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X821 VDDA.t721 GNDA.t410 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X822 VOUT+.t89 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X823 VOUT-.t99 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X824 GNDA.t804 GNDA.t802 VOUT-.t15 GNDA.t803 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X825 VDDA.t722 GNDA.t409 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X826 two_stage_opamp_dummy_magic_24_0.VD3.t19 two_stage_opamp_dummy_magic_24_0.Vb2.t19 two_stage_opamp_dummy_magic_24_0.X.t9 two_stage_opamp_dummy_magic_24_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X827 GNDA.t801 GNDA.t799 VDDA.t397 GNDA.t800 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X828 VOUT+.t90 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X829 VDDA.t723 GNDA.t408 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X830 VDDA.t724 GNDA.t407 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X831 VDDA.t725 GNDA.t406 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X832 GNDA.t798 GNDA.t796 two_stage_opamp_dummy_magic_24_0.VD1.t11 GNDA.t797 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X833 GNDA.t1004 two_stage_opamp_dummy_magic_24_0.Vb1.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X834 GNDA.t1005 two_stage_opamp_dummy_magic_24_0.Vb1.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X835 GNDA.t1006 two_stage_opamp_dummy_magic_24_0.Vb1.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X836 VDDA.t726 GNDA.t405 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X837 a_11420_30458.t0 a_11300_28850.t0 GNDA.t24 sky130_fd_pr__res_xhigh_po_0p35 l=6
X838 VDDA.t727 GNDA.t404 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X839 VDDA.t52 bgr_11_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t4 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X840 two_stage_opamp_dummy_magic_24_0.X.t8 two_stage_opamp_dummy_magic_24_0.Vb2.t20 two_stage_opamp_dummy_magic_24_0.VD3.t17 two_stage_opamp_dummy_magic_24_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X841 GNDA.t795 GNDA.t793 two_stage_opamp_dummy_magic_24_0.err_amp_out.t2 GNDA.t794 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X842 GNDA.t1007 two_stage_opamp_dummy_magic_24_0.Vb1.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X843 VOUT-.t100 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X844 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t3 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X845 two_stage_opamp_dummy_magic_24_0.VD4.t27 two_stage_opamp_dummy_magic_24_0.Vb3.t16 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X846 VDDA.t728 GNDA.t403 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X847 VDDA.t729 GNDA.t402 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X848 VOUT+.t91 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X849 bgr_11_0.V_TOP.t1 bgr_11_0.1st_Vout_1.t22 VDDA.t238 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X850 GNDA.t1008 two_stage_opamp_dummy_magic_24_0.Vb1.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X851 VDDA.t730 GNDA.t401 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X852 VOUT+.t92 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X853 VDDA.t731 GNDA.t400 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X854 VDDA.t732 GNDA.t399 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X855 two_stage_opamp_dummy_magic_24_0.VD4.t11 two_stage_opamp_dummy_magic_24_0.Vb2.t21 two_stage_opamp_dummy_magic_24_0.Y.t5 two_stage_opamp_dummy_magic_24_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X856 VOUT-.t101 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X857 VOUT+.t93 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X858 GNDA.t792 GNDA.t790 two_stage_opamp_dummy_magic_24_0.VD2.t9 GNDA.t791 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X859 VOUT+.t94 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X860 VDDA.t380 two_stage_opamp_dummy_magic_24_0.X.t43 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t10 GNDA.t864 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X861 VOUT+.t95 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X862 VOUT+.t96 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X863 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t13 bgr_11_0.NFET_GATE_10uA.t15 GNDA.t175 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X864 GNDA.t1009 two_stage_opamp_dummy_magic_24_0.Vb1.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X865 VDDA.t733 GNDA.t398 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X866 VDDA.t734 GNDA.t397 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X867 VDDA.t735 GNDA.t396 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X868 GNDA.t1010 two_stage_opamp_dummy_magic_24_0.Vb1.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X869 VDDA.t736 GNDA.t395 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X870 VDDA.t737 GNDA.t394 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X871 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X872 VOUT+.t97 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X873 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t12 bgr_11_0.PFET_GATE_10uA.t20 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X874 VDDA.t738 GNDA.t393 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X875 VDDA.t739 GNDA.t392 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X876 GNDA.t110 bgr_11_0.NFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_24_0.Vb2.t7 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X877 VDDA.t31 bgr_11_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t11 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X878 VDDA.t740 GNDA.t391 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X879 GNDA.t1011 two_stage_opamp_dummy_magic_24_0.Vb1.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X880 VDDA.t741 GNDA.t390 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X881 VOUT-.t102 two_stage_opamp_dummy_magic_24_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X882 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t7 GNDA.t787 GNDA.t789 GNDA.t788 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X883 bgr_11_0.V_TOP.t0 bgr_11_0.1st_Vout_1.t24 VDDA.t367 VDDA.t366 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X884 GNDA.t157 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_24_0.V_source.t15 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X885 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t1 a_13390_346.t0 GNDA.t166 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X886 VOUT+.t98 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X887 VDDA.t742 GNDA.t389 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X888 VDDA.t294 VDDA.t292 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t15 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X889 VDDA.t743 GNDA.t388 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X890 GNDA.t1012 two_stage_opamp_dummy_magic_24_0.Vb1.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X891 VOUT+.t99 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X892 GNDA.t1013 two_stage_opamp_dummy_magic_24_0.Vb1.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X893 VDDA.t744 GNDA.t387 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X894 GNDA.t1014 two_stage_opamp_dummy_magic_24_0.Vb1.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X895 VOUT+.t100 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X896 VDDA.t745 GNDA.t386 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X897 VDDA.t37 two_stage_opamp_dummy_magic_24_0.Vb3.t17 two_stage_opamp_dummy_magic_24_0.VD3.t34 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X898 GNDA.t1015 two_stage_opamp_dummy_magic_24_0.Vb1.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X899 bgr_11_0.1st_Vout_1.t25 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X900 VDDA.t746 GNDA.t468 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X901 VDDA.t747 GNDA.t467 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X902 bgr_11_0.PFET_GATE_10uA.t6 VDDA.t748 GNDA.t466 GNDA.t465 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X903 VOUT-.t103 two_stage_opamp_dummy_magic_24_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X904 VDDA.t749 GNDA.t385 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X905 VDDA.t750 GNDA.t384 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X906 GNDA.t35 a_5820_29044.t0 GNDA.t34 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X907 VDDA.t751 GNDA.t383 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X908 VOUT-.t104 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X909 VDDA.t752 GNDA.t382 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X910 VDDA.t753 GNDA.t381 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X911 VOUT-.t105 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X912 VOUT+.t101 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X913 VDDA.t173 two_stage_opamp_dummy_magic_24_0.Y.t41 VOUT+.t5 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X914 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t0 a_4380_346.t0 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X915 GNDA.t1016 two_stage_opamp_dummy_magic_24_0.Vb1.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X916 VOUT+.t102 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X917 VDDA.t754 GNDA.t380 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X918 VOUT+.t103 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X919 VOUT+.t104 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X920 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t3 two_stage_opamp_dummy_magic_24_0.X.t44 GNDA.t874 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X921 VDDA.t755 GNDA.t379 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X922 VDDA.t756 GNDA.t378 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X923 GNDA.t1017 two_stage_opamp_dummy_magic_24_0.Vb1.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X924 VDDA.t757 GNDA.t377 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X925 VOUT+.t105 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X926 GNDA.t743 GNDA.t786 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X927 bgr_11_0.V_mir1.t6 bgr_11_0.V_mir1.t5 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X928 VDDA.t160 two_stage_opamp_dummy_magic_24_0.Vb3.t18 two_stage_opamp_dummy_magic_24_0.VD4.t26 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X929 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X930 VDDA.t758 GNDA.t376 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X931 VDDA.t759 GNDA.t375 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X932 VDDA.t760 GNDA.t374 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X933 two_stage_opamp_dummy_magic_24_0.VD1.t10 GNDA.t783 GNDA.t785 GNDA.t784 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X934 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_24_0.X.t45 VDDA.t138 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X935 VDDA.t761 GNDA.t373 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X936 VDDA.t762 GNDA.t372 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X937 two_stage_opamp_dummy_magic_24_0.Y.t23 two_stage_opamp_dummy_magic_24_0.VD4.t32 two_stage_opamp_dummy_magic_24_0.VD4.t34 two_stage_opamp_dummy_magic_24_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X938 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_24_0.V_err_gate.t8 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X939 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t11 two_stage_opamp_dummy_magic_24_0.Y.t42 GNDA.t18 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X940 bgr_11_0.V_TOP.t39 VDDA.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X941 VDDA.t763 GNDA.t371 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X942 GNDA.t1018 two_stage_opamp_dummy_magic_24_0.Vb1.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X943 VOUT-.t106 two_stage_opamp_dummy_magic_24_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X944 bgr_11_0.V_TOP.t9 VDDA.t289 VDDA.t291 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X945 VDDA.t288 VDDA.t286 GNDA.t464 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X946 VDDA.t764 GNDA.t370 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X947 VDDA.t765 GNDA.t369 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X948 GNDA.t1019 two_stage_opamp_dummy_magic_24_0.Vb1.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X949 VOUT+.t106 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X950 VOUT-.t107 two_stage_opamp_dummy_magic_24_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X951 VDDA.t766 GNDA.t368 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X952 two_stage_opamp_dummy_magic_24_0.X.t7 two_stage_opamp_dummy_magic_24_0.Vb2.t22 two_stage_opamp_dummy_magic_24_0.VD3.t15 two_stage_opamp_dummy_magic_24_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X953 GNDA.t1020 two_stage_opamp_dummy_magic_24_0.Vb1.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X954 VDDA.t767 GNDA.t367 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X955 two_stage_opamp_dummy_magic_24_0.Y.t21 two_stage_opamp_dummy_magic_24_0.Vb1.t243 two_stage_opamp_dummy_magic_24_0.VD2.t12 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X956 VOUT+.t107 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X957 VDDA.t162 two_stage_opamp_dummy_magic_24_0.Vb3.t19 two_stage_opamp_dummy_magic_24_0.VD3.t33 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X958 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_24_0.Y.t43 VDDA.t8 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X959 GNDA.t1021 two_stage_opamp_dummy_magic_24_0.Vb1.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X960 VOUT-.t108 two_stage_opamp_dummy_magic_24_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X961 VDDA.t768 GNDA.t366 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X962 GNDA.t1022 two_stage_opamp_dummy_magic_24_0.Vb1.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X963 VDDA.t769 GNDA.t365 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X964 two_stage_opamp_dummy_magic_24_0.Vb3.t5 GNDA.t780 GNDA.t782 GNDA.t781 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X965 VDDA.t770 GNDA.t364 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X966 VDDA.t771 GNDA.t363 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X967 VDDA.t772 GNDA.t362 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X968 GNDA.t112 bgr_11_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_24_0.Vb3.t0 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X969 VDDA.t773 GNDA.t361 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 VDDA.t774 GNDA.t360 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X971 VDDA.t775 GNDA.t359 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X972 GNDA.t1023 two_stage_opamp_dummy_magic_24_0.Vb1.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X973 VDDA.t776 GNDA.t358 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X974 VOUT+.t108 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X975 VOUT-.t109 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X976 bgr_11_0.1st_Vout_2.t21 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X977 VOUT-.t110 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X978 VOUT+.t109 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X979 VOUT+.t110 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X980 VDDA.t413 bgr_11_0.V_mir2.t17 bgr_11_0.1st_Vout_2.t6 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X981 GNDA.t855 two_stage_opamp_dummy_magic_24_0.X.t46 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t2 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X982 GNDA.t1024 two_stage_opamp_dummy_magic_24_0.Vb1.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X983 VDDA.t777 GNDA.t357 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X984 VDDA.t778 GNDA.t356 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X985 VDDA.t779 GNDA.t355 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X986 VDDA.t780 GNDA.t354 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X987 VDDA.t781 GNDA.t353 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X988 VOUT+.t111 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X989 VDDA.t782 GNDA.t352 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X990 GNDA.t1025 two_stage_opamp_dummy_magic_24_0.Vb1.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X991 VDDA.t783 GNDA.t351 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X992 bgr_11_0.V_mir1.t4 bgr_11_0.V_mir1.t3 VDDA.t395 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X993 VDDA.t114 bgr_11_0.V_TOP.t40 bgr_11_0.START_UP.t2 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X994 two_stage_opamp_dummy_magic_24_0.V_source.t1 VIN+.t6 two_stage_opamp_dummy_magic_24_0.VD2.t0 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X995 VDDA.t784 GNDA.t350 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X996 VDDA.t785 GNDA.t349 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X997 VDDA.t407 two_stage_opamp_dummy_magic_24_0.Vb3.t20 two_stage_opamp_dummy_magic_24_0.VD4.t25 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X998 a_4100_3858.t0 two_stage_opamp_dummy_magic_24_0.V_tot.t3 GNDA.t119 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X999 VDDA.t12 two_stage_opamp_dummy_magic_24_0.X.t47 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t0 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1000 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1001 GNDA.t97 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_24_0.V_p_mir.t1 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1002 VDDA.t786 GNDA.t348 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1003 bgr_11_0.PFET_GATE_10uA.t4 VDDA.t283 VDDA.t285 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X1004 VDDA.t787 GNDA.t347 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1005 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1006 VDDA.t788 GNDA.t346 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1007 VDDA.t789 GNDA.t345 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1008 GNDA.t779 GNDA.t777 two_stage_opamp_dummy_magic_24_0.Vb2.t4 GNDA.t778 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X1009 GNDA.t99 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_24_0.V_source.t14 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1010 GNDA.t1026 two_stage_opamp_dummy_magic_24_0.Vb1.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1011 VDDA.t790 GNDA.t344 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1012 VDDA.t791 GNDA.t343 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1013 GNDA.t1027 two_stage_opamp_dummy_magic_24_0.Vb1.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1014 GNDA.t850 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t6 VOUT+.t16 GNDA.t849 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X1015 VDDA.t792 GNDA.t342 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1016 VDDA.t793 GNDA.t341 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1017 VDDA.t794 GNDA.t340 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1018 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t2 bgr_11_0.PFET_GATE_10uA.t22 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1019 VDDA.t795 GNDA.t339 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1020 VDDA.t282 VDDA.t279 VDDA.t281 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X1021 VDDA.t796 GNDA.t338 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1022 GNDA.t1028 two_stage_opamp_dummy_magic_24_0.Vb1.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1023 VDDA.t797 GNDA.t337 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1024 GNDA.t1029 two_stage_opamp_dummy_magic_24_0.Vb1.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1025 VOUT+.t112 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1026 GNDA.t59 a_6470_28850.t0 GNDA.t51 sky130_fd_pr__res_xhigh_po_0p35 l=6
X1027 VDDA.t798 GNDA.t336 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1028 VDDA.t409 two_stage_opamp_dummy_magic_24_0.Vb3.t21 two_stage_opamp_dummy_magic_24_0.VD4.t24 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1029 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1030 GNDA.t1030 two_stage_opamp_dummy_magic_24_0.Vb1.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1031 GNDA.t1031 two_stage_opamp_dummy_magic_24_0.Vb1.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 VOUT+.t113 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1033 GNDA.t1032 two_stage_opamp_dummy_magic_24_0.Vb1.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1034 VDDA.t799 GNDA.t335 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1035 VOUT+.t114 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1036 two_stage_opamp_dummy_magic_24_0.Y.t4 two_stage_opamp_dummy_magic_24_0.Vb2.t23 two_stage_opamp_dummy_magic_24_0.VD4.t5 two_stage_opamp_dummy_magic_24_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1037 two_stage_opamp_dummy_magic_24_0.V_source.t33 two_stage_opamp_dummy_magic_24_0.err_amp_out.t4 GNDA.t149 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1038 VDDA.t800 GNDA.t334 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1039 GNDA.t68 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t12 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1040 VDDA.t2 two_stage_opamp_dummy_magic_24_0.Y.t44 VOUT+.t0 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1041 VDDA.t801 GNDA.t333 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 VDDA.t802 GNDA.t332 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1043 GNDA.t1033 two_stage_opamp_dummy_magic_24_0.Vb1.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1044 VDDA.t803 GNDA.t331 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1045 two_stage_opamp_dummy_magic_24_0.Vb2.t3 GNDA.t774 GNDA.t776 GNDA.t775 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X1046 VDDA.t804 GNDA.t330 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1047 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t1 two_stage_opamp_dummy_magic_24_0.X.t48 GNDA.t64 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1048 bgr_11_0.1st_Vout_1.t28 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 VDDA.t805 GNDA.t329 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1050 bgr_11_0.V_p_1.t0 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t0 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X1051 bgr_11_0.1st_Vout_2.t24 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1052 VDDA.t92 bgr_11_0.V_mir2.t5 bgr_11_0.V_mir2.t6 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1053 VDDA.t278 VDDA.t276 VDDA.t278 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X1054 VDDA.t806 GNDA.t328 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1055 two_stage_opamp_dummy_magic_24_0.X.t24 two_stage_opamp_dummy_magic_24_0.Vb1.t244 two_stage_opamp_dummy_magic_24_0.VD1.t15 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1056 VDDA.t807 GNDA.t327 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1057 GNDA.t1034 two_stage_opamp_dummy_magic_24_0.Vb1.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1058 VOUT+.t115 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1059 VOUT+.t116 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1060 VDDA.t808 GNDA.t326 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1061 VDDA.t809 GNDA.t325 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1062 GNDA.t70 bgr_11_0.NFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_24_0.V_err_gate.t4 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1063 GNDA.t1035 two_stage_opamp_dummy_magic_24_0.Vb1.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1064 VOUT-.t111 two_stage_opamp_dummy_magic_24_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1065 VOUT-.t112 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1066 VOUT+.t117 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1067 GNDA.t1036 two_stage_opamp_dummy_magic_24_0.Vb1.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1068 VDDA.t810 GNDA.t324 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1069 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t10 two_stage_opamp_dummy_magic_24_0.Y.t45 GNDA.t12 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1070 bgr_11_0.1st_Vout_1.t29 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1071 VOUT-.t113 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1072 VOUT-.t114 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1073 two_stage_opamp_dummy_magic_24_0.X.t6 two_stage_opamp_dummy_magic_24_0.Vb2.t24 two_stage_opamp_dummy_magic_24_0.VD3.t13 two_stage_opamp_dummy_magic_24_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1074 VOUT-.t12 VDDA.t273 VDDA.t275 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X1075 VDDA.t811 GNDA.t323 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1076 VDDA.t812 GNDA.t322 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1077 a_12070_30308.t1 bgr_11_0.V_CUR_REF_REG.t1 GNDA.t143 sky130_fd_pr__res_xhigh_po_0p35 l=4
X1078 GNDA.t1037 two_stage_opamp_dummy_magic_24_0.Vb1.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1079 VDDA.t813 GNDA.t321 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1080 GNDA.t1038 two_stage_opamp_dummy_magic_24_0.Vb1.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1081 two_stage_opamp_dummy_magic_24_0.Y.t12 GNDA.t771 GNDA.t773 GNDA.t772 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X1082 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t4 two_stage_opamp_dummy_magic_24_0.Y.t46 VDDA.t21 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1083 bgr_11_0.1st_Vout_2.t25 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1084 VDDA.t814 GNDA.t320 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1085 VDDA.t815 GNDA.t319 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1086 VOUT-.t115 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1087 bgr_11_0.Vin-.t1 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t7 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1088 two_stage_opamp_dummy_magic_24_0.X.t19 two_stage_opamp_dummy_magic_24_0.Vb1.t245 two_stage_opamp_dummy_magic_24_0.VD1.t14 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1089 GNDA.t1039 two_stage_opamp_dummy_magic_24_0.Vb1.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1090 VDDA.t816 GNDA.t318 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1091 VDDA.t817 GNDA.t317 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1092 two_stage_opamp_dummy_magic_24_0.Vb2.t0 two_stage_opamp_dummy_magic_24_0.Vb2_2.t0 two_stage_opamp_dummy_magic_24_0.Vb2_2.t2 two_stage_opamp_dummy_magic_24_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X1093 two_stage_opamp_dummy_magic_24_0.Vb1.t221 two_stage_opamp_dummy_magic_24_0.Vb1.t220 two_stage_opamp_dummy_magic_24_0.Vb1_2.t2 GNDA.t878 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1094 VDDA.t818 GNDA.t316 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1095 VOUT+.t118 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1096 VOUT+.t119 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1097 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t1 bgr_11_0.V_TOP.t41 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1098 VDDA.t272 VDDA.t270 two_stage_opamp_dummy_magic_24_0.VD4.t20 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X1099 GNDA.t1040 two_stage_opamp_dummy_magic_24_0.Vb1.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1100 GNDA.t1041 two_stage_opamp_dummy_magic_24_0.Vb1.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1101 VDDA.t819 GNDA.t315 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1102 VDDA.t820 GNDA.t314 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1103 VOUT+.t120 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1104 two_stage_opamp_dummy_magic_24_0.Y.t3 two_stage_opamp_dummy_magic_24_0.Vb2.t25 two_stage_opamp_dummy_magic_24_0.VD4.t13 two_stage_opamp_dummy_magic_24_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1105 GNDA.t1042 two_stage_opamp_dummy_magic_24_0.Vb1.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1106 VDDA.t821 GNDA.t313 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1107 VDDA.t17 bgr_11_0.1st_Vout_2.t26 bgr_11_0.PFET_GATE_10uA.t0 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1108 bgr_11_0.1st_Vout_1.t30 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1109 VDDA.t822 GNDA.t312 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1110 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t63 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X1111 VDDA.t823 GNDA.t311 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1112 GNDA.t120 two_stage_opamp_dummy_magic_24_0.X.t49 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t0 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1113 VDDA.t824 GNDA.t310 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1114 two_stage_opamp_dummy_magic_24_0.V_source.t4 VIN+.t7 two_stage_opamp_dummy_magic_24_0.VD2.t2 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1115 GNDA.t1043 two_stage_opamp_dummy_magic_24_0.Vb1.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1116 GNDA.t1044 two_stage_opamp_dummy_magic_24_0.Vb1.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1117 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t10 GNDA.t769 GNDA.t770 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X1118 VDDA.t825 GNDA.t309 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1119 GNDA.t1045 two_stage_opamp_dummy_magic_24_0.Vb1.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1120 VDDA.t826 GNDA.t308 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1121 VOUT-.t116 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1122 VOUT-.t117 two_stage_opamp_dummy_magic_24_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1123 VOUT-.t118 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1124 VDDA.t827 GNDA.t307 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1125 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t267 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X1126 VDDA.t828 GNDA.t463 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1127 VDDA.t829 GNDA.t462 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1128 GNDA.t1046 two_stage_opamp_dummy_magic_24_0.Vb1.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1129 VDDA.t266 VDDA.t264 two_stage_opamp_dummy_magic_24_0.Vb2_2.t9 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X1130 GNDA.t1047 two_stage_opamp_dummy_magic_24_0.Vb1.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1131 VDDA.t77 bgr_11_0.PFET_GATE_10uA.t23 bgr_11_0.V_CUR_REF_REG.t0 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1132 GNDA.t1048 two_stage_opamp_dummy_magic_24_0.Vb1.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1133 VOUT-.t119 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1134 VOUT-.t120 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1135 GNDA.t31 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t7 VOUT-.t0 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X1136 VDDA.t830 GNDA.t461 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1137 VOUT-.t121 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1138 VDDA.t831 GNDA.t460 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1139 GNDA.t768 GNDA.t765 GNDA.t767 GNDA.t766 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X1140 GNDA.t151 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_24_0.V_source.t13 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1141 VDDA.t832 GNDA.t459 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1142 two_stage_opamp_dummy_magic_24_0.VD3.t32 two_stage_opamp_dummy_magic_24_0.Vb3.t22 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1143 VDDA.t833 GNDA.t458 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1144 VDDA.t263 VDDA.t261 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t4 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X1145 VDDA.t834 GNDA.t457 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1146 VDDA.t835 GNDA.t456 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1147 a_5700_30308.t1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t6 GNDA.t34 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X1148 VDDA.t836 GNDA.t455 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1149 bgr_11_0.V_TOP.t42 VDDA.t185 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1150 GNDA.t1049 two_stage_opamp_dummy_magic_24_0.Vb1.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1151 VDDA.t837 GNDA.t454 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1152 VDDA.t838 GNDA.t453 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1153 VDDA.t839 GNDA.t452 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1154 GNDA.t1050 two_stage_opamp_dummy_magic_24_0.Vb1.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1155 VDDA.t840 GNDA.t451 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1156 VOUT+.t121 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1157 VDDA.t841 GNDA.t450 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1158 VDDA.t842 GNDA.t449 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1159 VOUT+.t122 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1160 VDDA.t843 GNDA.t448 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1161 bgr_11_0.1st_Vout_1.t2 bgr_11_0.V_mir1.t17 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1162 GNDA.t447 VDDA.t844 bgr_11_0.V_p_2.t2 GNDA.t446 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X1163 VDDA.t845 GNDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1164 GNDA.t1051 two_stage_opamp_dummy_magic_24_0.Vb1.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1165 VDDA.t846 GNDA.t305 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1166 two_stage_opamp_dummy_magic_24_0.VD4.t23 two_stage_opamp_dummy_magic_24_0.Vb3.t23 VDDA.t392 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1167 two_stage_opamp_dummy_magic_24_0.X.t5 two_stage_opamp_dummy_magic_24_0.Vb2.t26 two_stage_opamp_dummy_magic_24_0.VD3.t11 two_stage_opamp_dummy_magic_24_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1168 VDDA.t847 GNDA.t304 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1169 VOUT-.t122 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1170 VDDA.t848 GNDA.t303 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1171 VOUT-.t123 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1172 two_stage_opamp_dummy_magic_24_0.VD4.t15 two_stage_opamp_dummy_magic_24_0.Vb2.t27 two_stage_opamp_dummy_magic_24_0.Y.t2 two_stage_opamp_dummy_magic_24_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1173 bgr_11_0.V_TOP.t43 VDDA.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1174 GNDA.t1052 two_stage_opamp_dummy_magic_24_0.Vb1.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1175 VDDA.t849 GNDA.t302 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1176 VOUT-.t124 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1177 GNDA.t743 GNDA.t764 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X1178 VDDA.t850 GNDA.t301 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1179 VDDA.t851 GNDA.t300 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1180 VDDA.t852 GNDA.t299 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1181 two_stage_opamp_dummy_magic_24_0.VD3.t2 two_stage_opamp_dummy_magic_24_0.VD3.t0 two_stage_opamp_dummy_magic_24_0.X.t1 two_stage_opamp_dummy_magic_24_0.VD3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X1182 two_stage_opamp_dummy_magic_24_0.X.t21 two_stage_opamp_dummy_magic_24_0.Vb1.t246 two_stage_opamp_dummy_magic_24_0.VD1.t13 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1183 VDDA.t853 GNDA.t298 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1184 VDDA.t854 GNDA.t297 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1185 VDDA.t855 GNDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1186 GNDA.t1053 two_stage_opamp_dummy_magic_24_0.Vb1.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1187 VDDA.t856 GNDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1188 VOUT+.t123 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1189 two_stage_opamp_dummy_magic_24_0.VD3.t31 two_stage_opamp_dummy_magic_24_0.Vb3.t24 VDDA.t208 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1190 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_24_0.Y.t47 GNDA.t48 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1191 VOUT-.t14 GNDA.t761 GNDA.t763 GNDA.t762 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X1192 VDDA.t857 GNDA.t294 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1193 VDDA.t858 GNDA.t293 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1194 VDDA.t216 bgr_11_0.V_TOP.t44 bgr_11_0.Vin-.t4 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1195 VOUT+.t124 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1196 bgr_11_0.V_TOP.t45 VDDA.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1197 GNDA.t1054 two_stage_opamp_dummy_magic_24_0.Vb1.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1198 GNDA.t1055 two_stage_opamp_dummy_magic_24_0.Vb1.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1199 VOUT-.t11 two_stage_opamp_dummy_magic_24_0.X.t50 VDDA.t220 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1200 VDDA.t859 GNDA.t292 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1201 VOUT+.t125 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1202 VDDA.t860 GNDA.t291 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1203 two_stage_opamp_dummy_magic_24_0.Vb1.t0 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1204 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t3 two_stage_opamp_dummy_magic_24_0.Y.t48 VDDA.t174 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1205 GNDA.t1056 two_stage_opamp_dummy_magic_24_0.Vb1.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1206 GNDA.t1057 two_stage_opamp_dummy_magic_24_0.Vb1.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1207 VDDA.t861 GNDA.t290 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1208 VOUT+.t126 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1209 VOUT-.t125 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1210 VDDA.t94 bgr_11_0.V_mir2.t3 bgr_11_0.V_mir2.t4 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1211 VOUT+.t127 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1212 VDDA.t862 GNDA.t289 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1213 VDDA.t152 bgr_11_0.V_mir1.t1 bgr_11_0.V_mir1.t2 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1214 two_stage_opamp_dummy_magic_24_0.X.t20 two_stage_opamp_dummy_magic_24_0.Vb1.t247 two_stage_opamp_dummy_magic_24_0.VD1.t12 GNDA.t865 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1215 VDDA.t863 GNDA.t288 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1216 GNDA.t1058 two_stage_opamp_dummy_magic_24_0.Vb1.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1217 VDDA.t864 GNDA.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1218 VDDA.t865 GNDA.t286 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1219 VDDA.t866 GNDA.t285 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1220 GNDA.t1059 two_stage_opamp_dummy_magic_24_0.Vb1.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1221 VDDA.t867 GNDA.t284 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1222 VOUT-.t126 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1223 VDDA.t868 GNDA.t283 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1224 VDDA.t869 GNDA.t282 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1225 VOUT+.t128 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1226 VOUT-.t127 two_stage_opamp_dummy_magic_24_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1227 a_4220_3858.t0 two_stage_opamp_dummy_magic_24_0.V_tot.t0 GNDA.t40 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X1228 GNDA.t1060 two_stage_opamp_dummy_magic_24_0.Vb1.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1229 VOUT-.t128 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1230 GNDA.t1061 two_stage_opamp_dummy_magic_24_0.Vb1.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1231 VDDA.t870 GNDA.t281 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1232 VOUT-.t129 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1233 VOUT-.t130 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1234 VDDA.t871 GNDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1235 VOUT-.t131 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1236 two_stage_opamp_dummy_magic_24_0.V_source.t39 VIN+.t8 two_stage_opamp_dummy_magic_24_0.VD2.t21 GNDA.t851 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1237 VDDA.t872 GNDA.t279 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1238 VOUT+.t129 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1239 GNDA.t760 GNDA.t758 two_stage_opamp_dummy_magic_24_0.X.t14 GNDA.t759 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X1240 VDDA.t873 GNDA.t278 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1241 GNDA.t1062 two_stage_opamp_dummy_magic_24_0.Vb1.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1242 VDDA.t874 GNDA.t277 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1243 VDDA.t875 GNDA.t276 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1244 VDDA.t876 GNDA.t275 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1245 GNDA.t1063 two_stage_opamp_dummy_magic_24_0.Vb1.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1246 VOUT+.t130 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1247 VDDA.t877 GNDA.t274 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1248 VDDA.t878 GNDA.t273 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1249 VOUT+.t131 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1250 two_stage_opamp_dummy_magic_24_0.Vb1.t227 two_stage_opamp_dummy_magic_24_0.Vb1.t226 two_stage_opamp_dummy_magic_24_0.Vb1_2.t1 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1251 bgr_11_0.V_TOP.t46 VDDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1252 VDDA.t879 GNDA.t272 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1253 GNDA.t1064 two_stage_opamp_dummy_magic_24_0.Vb1.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1254 GNDA.t1065 two_stage_opamp_dummy_magic_24_0.Vb1.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1255 GNDA.t1066 two_stage_opamp_dummy_magic_24_0.Vb1.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1256 VDDA.t880 GNDA.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1257 a_6350_30458.t0 bgr_11_0.Vin+.t1 GNDA.t51 sky130_fd_pr__res_xhigh_po_0p35 l=6
X1258 two_stage_opamp_dummy_magic_24_0.Vb2_2.t8 two_stage_opamp_dummy_magic_24_0.Vb2.t28 VDDA.t242 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X1259 GNDA.t153 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_24_0.V_source.t12 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1260 VDDA.t881 GNDA.t270 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1261 GNDA.t1067 two_stage_opamp_dummy_magic_24_0.Vb1.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1262 VDDA.t882 GNDA.t269 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1263 VOUT+.t132 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1264 GNDA.t1068 two_stage_opamp_dummy_magic_24_0.Vb1.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1265 VDDA.t883 GNDA.t268 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1266 VOUT+.t133 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1267 GNDA.t757 GNDA.t755 two_stage_opamp_dummy_magic_24_0.Y.t11 GNDA.t756 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X1268 VDDA.t884 GNDA.t267 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1269 VOUT+.t134 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1270 GNDA.t1069 two_stage_opamp_dummy_magic_24_0.Vb1.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1271 VDDA.t885 GNDA.t266 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1272 two_stage_opamp_dummy_magic_24_0.VD4.t22 two_stage_opamp_dummy_magic_24_0.Vb3.t25 VDDA.t210 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1273 bgr_11_0.Vin-.t3 bgr_11_0.V_TOP.t47 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1274 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t1 bgr_11_0.PFET_GATE_10uA.t25 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1275 two_stage_opamp_dummy_magic_24_0.VD4.t17 two_stage_opamp_dummy_magic_24_0.Vb2.t29 two_stage_opamp_dummy_magic_24_0.Y.t1 two_stage_opamp_dummy_magic_24_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1276 VOUT-.t132 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1277 VDDA.t886 GNDA.t265 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1278 VDDA.t125 bgr_11_0.PFET_GATE_10uA.t26 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t0 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1279 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t2 GNDA.t752 GNDA.t754 GNDA.t753 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X1280 VDDA.t887 GNDA.t264 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1281 VDDA.t888 GNDA.t263 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1282 GNDA.t1070 two_stage_opamp_dummy_magic_24_0.Vb1.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1283 VDDA.t889 GNDA.t262 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1284 bgr_11_0.cap_res1.t20 bgr_11_0.V_TOP.t13 GNDA.t877 sky130_fd_pr__res_high_po_0p35 l=2.05
X1285 VDDA.t203 bgr_11_0.1st_Vout_2.t27 bgr_11_0.PFET_GATE_10uA.t3 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1286 VDDA.t890 GNDA.t261 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1287 VOUT-.t133 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1288 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1289 GNDA.t1071 two_stage_opamp_dummy_magic_24_0.Vb1.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1290 VDDA.t891 GNDA.t260 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1291 VOUT-.t134 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1292 VOUT-.t135 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1293 VDDA.t892 GNDA.t259 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1294 VDDA.t893 GNDA.t258 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1295 VDDA.t894 GNDA.t257 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1296 GNDA.t114 bgr_11_0.NFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_24_0.Vb3.t1 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1297 two_stage_opamp_dummy_magic_24_0.VD3.t30 two_stage_opamp_dummy_magic_24_0.Vb3.t26 VDDA.t232 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1298 VOUT+.t135 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1299 GNDA.t1072 two_stage_opamp_dummy_magic_24_0.Vb1.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1300 GNDA.t1073 two_stage_opamp_dummy_magic_24_0.Vb1.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1301 VOUT+.t136 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1302 VDDA.t895 GNDA.t256 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1303 VOUT+.t137 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1304 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1305 VDDA.t896 GNDA.t255 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1306 VDDA.t897 GNDA.t254 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1307 GNDA.t1074 two_stage_opamp_dummy_magic_24_0.Vb1.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1308 two_stage_opamp_dummy_magic_24_0.VD3.t9 two_stage_opamp_dummy_magic_24_0.Vb2.t30 two_stage_opamp_dummy_magic_24_0.X.t4 two_stage_opamp_dummy_magic_24_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1309 VDDA.t898 GNDA.t253 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1310 two_stage_opamp_dummy_magic_24_0.V_source.t11 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t28 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1311 VDDA.t899 GNDA.t252 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1312 GNDA.t1075 two_stage_opamp_dummy_magic_24_0.Vb1.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1313 two_stage_opamp_dummy_magic_24_0.V_source.t10 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t29 GNDA.t39 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1314 VDDA.t900 GNDA.t251 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1315 VOUT-.t136 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1316 VOUT-.t137 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1317 two_stage_opamp_dummy_magic_24_0.err_amp_out.t0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_24_0.V_err_p.t0 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1318 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_24_0.Y.t49 GNDA.t128 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1319 VOUT+.t4 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t8 GNDA.t75 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X1320 VDDA.t901 GNDA.t250 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1321 VDDA.t902 GNDA.t249 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1322 GNDA.t1076 two_stage_opamp_dummy_magic_24_0.Vb1.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1323 VDDA.t903 GNDA.t248 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1324 VOUT-.t138 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1325 VOUT-.t139 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1326 VOUT+.t138 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1327 VDDA.t904 GNDA.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1328 GNDA.t743 GNDA.t751 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X1329 GNDA.t1077 two_stage_opamp_dummy_magic_24_0.Vb1.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1330 two_stage_opamp_dummy_magic_24_0.Vb2_2.t7 two_stage_opamp_dummy_magic_24_0.Vb2.t1 two_stage_opamp_dummy_magic_24_0.Vb2.t2 two_stage_opamp_dummy_magic_24_0.Vb2_2.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1331 VOUT+.t139 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1332 VOUT-.t9 two_stage_opamp_dummy_magic_24_0.X.t51 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1333 VOUT-.t140 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1334 VOUT-.t141 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1335 VDDA.t39 bgr_11_0.V_mir2.t18 bgr_11_0.1st_Vout_2.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1336 VDDA.t905 GNDA.t246 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1337 two_stage_opamp_dummy_magic_24_0.VD4.t19 two_stage_opamp_dummy_magic_24_0.Vb2.t31 two_stage_opamp_dummy_magic_24_0.Y.t0 two_stage_opamp_dummy_magic_24_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1338 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_24_0.Y.t50 VDDA.t4 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1339 VDDA.t906 GNDA.t245 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1340 two_stage_opamp_dummy_magic_24_0.X.t13 GNDA.t748 GNDA.t750 GNDA.t749 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X1341 GNDA.t1078 two_stage_opamp_dummy_magic_24_0.Vb1.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1342 VDDA.t907 GNDA.t244 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1343 VOUT-.t142 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1344 two_stage_opamp_dummy_magic_24_0.V_source.t27 VIN-.t6 two_stage_opamp_dummy_magic_24_0.VD1.t3 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1345 VOUT-.t143 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1346 VDDA.t908 GNDA.t243 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1347 VOUT+.t12 VDDA.t258 VDDA.t260 VDDA.t259 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X1348 VOUT+.t140 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1349 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t1 bgr_11_0.PFET_GATE_10uA.t27 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1350 VOUT+.t1 two_stage_opamp_dummy_magic_24_0.Y.t51 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1351 bgr_11_0.V_TOP.t48 VDDA.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1352 VDDA.t909 GNDA.t242 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1353 VDDA.t910 GNDA.t241 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1354 VDDA.t911 GNDA.t240 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1355 GNDA.t1079 two_stage_opamp_dummy_magic_24_0.Vb1.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1356 VDDA.t912 GNDA.t239 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1357 VDDA.t913 GNDA.t238 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1358 VOUT+.t3 two_stage_opamp_dummy_magic_24_0.Y.t52 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1359 GNDA.t1080 two_stage_opamp_dummy_magic_24_0.Vb1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1360 VDDA.t914 GNDA.t237 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1361 VOUT+.t141 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1362 VOUT+.t142 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1363 VOUT+.t143 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1364 VOUT-.t144 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1365 VDDA.t915 GNDA.t236 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1366 bgr_11_0.Vin+.t0 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t41 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X1367 VDDA.t916 GNDA.t235 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1368 two_stage_opamp_dummy_magic_24_0.V_source.t3 VIN+.t9 two_stage_opamp_dummy_magic_24_0.VD2.t1 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1369 VDDA.t917 GNDA.t234 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1370 GNDA.t1081 two_stage_opamp_dummy_magic_24_0.Vb1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1371 VDDA.t918 GNDA.t233 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1372 VDDA.t393 GNDA.t745 GNDA.t747 GNDA.t746 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X1373 VDDA.t919 GNDA.t232 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1374 GNDA.t116 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_24_0.Vb2.t6 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1375 two_stage_opamp_dummy_magic_24_0.V_source.t34 VIN-.t7 two_stage_opamp_dummy_magic_24_0.VD1.t2 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1376 GNDA.t1082 two_stage_opamp_dummy_magic_24_0.Vb1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1377 VDDA.t234 two_stage_opamp_dummy_magic_24_0.Vb3.t27 two_stage_opamp_dummy_magic_24_0.VD3.t29 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1378 VDDA.t920 GNDA.t231 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1379 VDDA.t921 GNDA.t230 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1380 GNDA.t1083 two_stage_opamp_dummy_magic_24_0.Vb1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1381 VDDA.t922 GNDA.t229 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1382 VOUT-.t145 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1383 VDDA.t99 bgr_11_0.V_TOP.t49 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t0 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1384 VDDA.t377 bgr_11_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t10 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1385 VDDA.t923 GNDA.t228 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1386 VOUT+.t144 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1387 two_stage_opamp_dummy_magic_24_0.Vb2.t5 bgr_11_0.NFET_GATE_10uA.t22 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1388 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t14 VDDA.t255 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X1389 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1390 VOUT-.t146 two_stage_opamp_dummy_magic_24_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1391 VDDA.t924 GNDA.t227 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1392 GNDA.t78 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_24_0.V_source.t9 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1393 VDDA.t925 GNDA.t226 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1394 VDDA.t218 two_stage_opamp_dummy_magic_24_0.X.t52 VOUT-.t10 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1395 VDDA.t926 GNDA.t225 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1396 VDDA.t927 GNDA.t224 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1397 GNDA.t1084 two_stage_opamp_dummy_magic_24_0.Vb1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1398 two_stage_opamp_dummy_magic_24_0.VD2.t11 two_stage_opamp_dummy_magic_24_0.Vb1.t248 two_stage_opamp_dummy_magic_24_0.Y.t20 GNDA.t866 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1399 VDDA.t928 GNDA.t223 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1400 VDDA.t929 GNDA.t222 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1401 VDDA.t930 GNDA.t221 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1402 VDDA.t931 GNDA.t220 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1403 GNDA.t1085 two_stage_opamp_dummy_magic_24_0.Vb1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1404 VDDA.t932 GNDA.t219 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1405 VOUT-.t147 two_stage_opamp_dummy_magic_24_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1406 VDDA.t933 GNDA.t218 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1407 VOUT+.t145 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1408 VDDA.t137 bgr_11_0.V_mir2.t1 bgr_11_0.V_mir2.t2 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1409 GNDA.t1086 two_stage_opamp_dummy_magic_24_0.Vb1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1410 VDDA.t934 GNDA.t217 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1411 VDDA.t935 GNDA.t216 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1412 VDDA.t936 GNDA.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1413 two_stage_opamp_dummy_magic_24_0.VD3.t7 two_stage_opamp_dummy_magic_24_0.Vb2.t32 two_stage_opamp_dummy_magic_24_0.X.t3 two_stage_opamp_dummy_magic_24_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1414 VOUT+.t146 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1415 VOUT+.t147 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1416 VDDA.t937 GNDA.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1417 VDDA.t938 GNDA.t213 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1418 VDDA.t939 GNDA.t212 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1419 two_stage_opamp_dummy_magic_24_0.Vb1.t218 GNDA.t739 GNDA.t741 GNDA.t740 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X1420 VDDA.t940 GNDA.t211 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1421 VDDA.t941 GNDA.t210 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1422 VDDA.t942 GNDA.t209 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1423 GNDA.t125 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t9 VOUT-.t7 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X1424 VDDA.t943 GNDA.t208 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1425 GNDA.t1087 two_stage_opamp_dummy_magic_24_0.Vb1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1426 VDDA.t944 GNDA.t207 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1427 VDDA.t945 GNDA.t206 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1428 VDDA.t236 two_stage_opamp_dummy_magic_24_0.Vb3.t28 two_stage_opamp_dummy_magic_24_0.VD3.t28 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1429 VDDA.t946 GNDA.t205 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1430 VDDA.t947 GNDA.t204 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1431 VOUT+.t148 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1432 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1433 VDDA.t948 GNDA.t203 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1434 VOUT+.t149 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1435 GNDA.t1088 two_stage_opamp_dummy_magic_24_0.Vb1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1436 GNDA.t1089 two_stage_opamp_dummy_magic_24_0.Vb1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1437 VOUT-.t148 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1438 VOUT-.t149 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1439 VOUT-.t150 two_stage_opamp_dummy_magic_24_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1440 VOUT+.t150 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1441 VDDA.t949 GNDA.t202 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1442 VDDA.t386 bgr_11_0.V_mir1.t18 bgr_11_0.1st_Vout_1.t6 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1443 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_24_0.V_err_gate.t0 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1444 two_stage_opamp_dummy_magic_24_0.V_source.t8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t31 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1445 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_24_0.Y.t53 GNDA.t49 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1446 VDDA.t950 GNDA.t201 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1447 VDDA.t951 GNDA.t200 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1448 VDDA.t197 two_stage_opamp_dummy_magic_24_0.V_err_gate.t9 two_stage_opamp_dummy_magic_24_0.V_err_p.t1 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1449 VDDA.t952 GNDA.t199 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1450 VDDA.t953 GNDA.t198 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1451 bgr_11_0.1st_Vout_2.t4 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t1 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X1452 GNDA.t1090 two_stage_opamp_dummy_magic_24_0.Vb1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1453 VOUT+.t151 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1454 VDDA.t954 GNDA.t197 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1455 VOUT-.t8 two_stage_opamp_dummy_magic_24_0.X.t53 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1456 bgr_11_0.1st_Vout_2.t31 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1457 VDDA.t955 GNDA.t196 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1458 bgr_11_0.START_UP.t1 bgr_11_0.START_UP.t0 bgr_11_0.START_UP_NFET1.t0 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X1459 GNDA.t1091 two_stage_opamp_dummy_magic_24_0.Vb1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1460 VDDA.t956 GNDA.t195 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1461 VDDA.t957 GNDA.t194 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1462 VDDA.t958 GNDA.t193 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1463 GNDA.t1092 two_stage_opamp_dummy_magic_24_0.Vb1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1464 VDDA.t959 GNDA.t192 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1465 VOUT+.t152 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1466 VOUT+.t153 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1467 VOUT+.t154 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1468 a_4220_3858.t1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t4 GNDA.t176 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X1469 two_stage_opamp_dummy_magic_24_0.V_source.t30 VIN-.t8 two_stage_opamp_dummy_magic_24_0.VD1.t1 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1470 VOUT+.t155 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1471 VDDA.t960 GNDA.t191 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1472 a_11420_30458.t1 bgr_11_0.Vin-.t0 GNDA.t33 sky130_fd_pr__res_xhigh_po_0p35 l=6
X1473 VOUT+.t8 two_stage_opamp_dummy_magic_24_0.Y.t54 VDDA.t240 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1474 bgr_11_0.1st_Vout_1.t32 bgr_11_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1475 VDDA.t961 GNDA.t190 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1476 GNDA.t61 a_11950_29100.t1 GNDA.t60 sky130_fd_pr__res_xhigh_po_0p35 l=4
X1477 GNDA.t445 VDDA.t252 VDDA.t254 VDDA.t253 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X1478 GNDA.t1093 two_stage_opamp_dummy_magic_24_0.Vb1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1479 VDDA.t962 GNDA.t189 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1480 VDDA.t963 GNDA.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1481 GNDA.t1094 two_stage_opamp_dummy_magic_24_0.Vb1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1482 GNDA.t1095 two_stage_opamp_dummy_magic_24_0.Vb1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1483 VDDA.t964 GNDA.t187 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1484 VDDA.t965 GNDA.t186 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1485 VDDA.t966 GNDA.t185 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1486 VOUT-.t151 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1487 VDDA.t251 VDDA.t249 bgr_11_0.V_TOP.t8 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X1488 bgr_11_0.1st_Vout_2.t32 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1489 GNDA.t1096 two_stage_opamp_dummy_magic_24_0.Vb1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1490 GNDA.t1097 two_stage_opamp_dummy_magic_24_0.Vb1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1491 VOUT-.t152 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1492 VOUT-.t153 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1493 VOUT+.t156 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1494 two_stage_opamp_dummy_magic_24_0.V_source.t6 VIN+.t10 two_stage_opamp_dummy_magic_24_0.VD2.t3 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1495 GNDA.t1098 two_stage_opamp_dummy_magic_24_0.Vb1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1496 VDDA.t967 GNDA.t184 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1497 VOUT-.t154 two_stage_opamp_dummy_magic_24_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1498 VDDA.t379 two_stage_opamp_dummy_magic_24_0.X.t54 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t9 GNDA.t863 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1499 VDDA.t968 GNDA.t183 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1500 VOUT-.t155 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1501 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t9 VIN-.t9 two_stage_opamp_dummy_magic_24_0.V_p_mir.t0 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1502 two_stage_opamp_dummy_magic_24_0.V_source.t40 VIN-.t10 two_stage_opamp_dummy_magic_24_0.VD1.t0 GNDA.t870 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1503 VOUT-.t156 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 VDDA.n2833 VDDA.t258 1231.74
R1 VDDA.n2836 VDDA.t322 1231.74
R2 VDDA.n2726 VDDA.t334 1231.74
R3 VDDA.n2729 VDDA.t273 1231.74
R4 VDDA.n2756 VDDA.t301 794.668
R5 VDDA.n2760 VDDA.t295 794.668
R6 VDDA.n2740 VDDA.t356 794.668
R7 VDDA.n2785 VDDA.t325 794.668
R8 VDDA.n2405 VDDA.t306 708.125
R9 VDDA.t306 VDDA.n2382 708.125
R10 VDDA.n2412 VDDA.t251 708.125
R11 VDDA.t251 VDDA.n2363 708.125
R12 VDDA.n1962 VDDA.t354 676.966
R13 VDDA.n2845 VDDA.t270 672.293
R14 VDDA.n2848 VDDA.t340 672.293
R15 VDDA.n2688 VDDA.t359 672.293
R16 VDDA.n2691 VDDA.t313 672.293
R17 VDDA.n2792 VDDA.t276 661.375
R18 VDDA.n2795 VDDA.t319 661.375
R19 VDDA.t290 VDDA.n2410 660.001
R20 VDDA.n2404 VDDA.t305 657.76
R21 VDDA.n2411 VDDA.t250 657.76
R22 VDDA.t317 VDDA.n1961 643.038
R23 VDDA.t299 VDDA.n2200 643.037
R24 VDDA.n2201 VDDA.t332 643.037
R25 VDDA.t293 VDDA.n2185 643.037
R26 VDDA.n2186 VDDA.t256 643.037
R27 VDDA.n2195 VDDA.t363 642.992
R28 VDDA.t329 VDDA.n2194 642.992
R29 VDDA.t268 VDDA.n2177 642.992
R30 VDDA.n2178 VDDA.t351 642.992
R31 VDDA.n2030 VDDA.t343 595.842
R32 VDDA.n2817 VDDA.t337 589.076
R33 VDDA.n2820 VDDA.t286 589.076
R34 VDDA.n2710 VDDA.t310 589.076
R35 VDDA.n2713 VDDA.t252 589.076
R36 VDDA.n1987 VDDA.n1955 587.407
R37 VDDA.n1983 VDDA.n1982 587.407
R38 VDDA.n2000 VDDA.n1999 587.407
R39 VDDA.n1994 VDDA.n1949 587.407
R40 VDDA.n1999 VDDA.n1998 585
R41 VDDA.n1997 VDDA.n1994 585
R42 VDDA.n1985 VDDA.n1955 585
R43 VDDA.n1984 VDDA.n1983 585
R44 VDDA.n2773 VDDA.n2772 585
R45 VDDA.n2770 VDDA.n2769 585
R46 VDDA.n2784 VDDA.n2733 585
R47 VDDA.n2755 VDDA.n2742 585
R48 VDDA.n2014 VDDA.t307 579.775
R49 VDDA.t284 VDDA.n2403 540.818
R50 VDDA.n2019 VDDA.t309 464.281
R51 VDDA.n2016 VDDA.t309 464.281
R52 VDDA.n2025 VDDA.t346 464.281
R53 VDDA.t346 VDDA.n2008 464.281
R54 VDDA.n2799 VDDA.t279 456.526
R55 VDDA.n2802 VDDA.t264 456.526
R56 VDDA.n2188 VDDA.t328 441.2
R57 VDDA.n2196 VDDA.t362 441.2
R58 VDDA.n2179 VDDA.t350 441.2
R59 VDDA.n2176 VDDA.t267 441.2
R60 VDDA.n1960 VDDA.t316 413.084
R61 VDDA.n1963 VDDA.t353 413.084
R62 VDDA.n2197 VDDA.t298 409.067
R63 VDDA.n2202 VDDA.t331 409.067
R64 VDDA.t305 VDDA.t387 407.144
R65 VDDA.t387 VDDA.t412 407.144
R66 VDDA.t412 VDDA.t126 407.144
R67 VDDA.t126 VDDA.t93 407.144
R68 VDDA.t93 VDDA.t169 407.144
R69 VDDA.t169 VDDA.t16 407.144
R70 VDDA.t16 VDDA.t402 407.144
R71 VDDA.t402 VDDA.t38 407.144
R72 VDDA.t38 VDDA.t410 407.144
R73 VDDA.t410 VDDA.t91 407.144
R74 VDDA.t91 VDDA.t141 407.144
R75 VDDA.t141 VDDA.t202 407.144
R76 VDDA.t202 VDDA.t139 407.144
R77 VDDA.t139 VDDA.t41 407.144
R78 VDDA.t41 VDDA.t128 407.144
R79 VDDA.t128 VDDA.t136 407.144
R80 VDDA.t136 VDDA.t153 407.144
R81 VDDA.t153 VDDA.t404 407.144
R82 VDDA.t404 VDDA.t284 407.144
R83 VDDA.t250 VDDA.t237 407.144
R84 VDDA.t237 VDDA.t151 407.144
R85 VDDA.t151 VDDA.t226 407.144
R86 VDDA.t226 VDDA.t385 407.144
R87 VDDA.t385 VDDA.t69 407.144
R88 VDDA.t69 VDDA.t417 407.144
R89 VDDA.t417 VDDA.t368 407.144
R90 VDDA.t368 VDDA.t147 407.144
R91 VDDA.t147 VDDA.t130 407.144
R92 VDDA.t130 VDDA.t149 407.144
R93 VDDA.t149 VDDA.t71 407.144
R94 VDDA.t71 VDDA.t419 407.144
R95 VDDA.t419 VDDA.t366 407.144
R96 VDDA.t366 VDDA.t19 407.144
R97 VDDA.t19 VDDA.t394 407.144
R98 VDDA.t394 VDDA.t222 407.144
R99 VDDA.t222 VDDA.t224 407.144
R100 VDDA.t224 VDDA.t415 407.144
R101 VDDA.t415 VDDA.t290 407.144
R102 VDDA.n2801 VDDA.t265 397.784
R103 VDDA.t280 VDDA.n2800 397.784
R104 VDDA.n2182 VDDA.t292 390.322
R105 VDDA.n2187 VDDA.t255 390.322
R106 VDDA.t304 VDDA.n2405 379.582
R107 VDDA.t249 VDDA.n2412 379.582
R108 VDDA.n2402 VDDA.t283 379.277
R109 VDDA.t122 VDDA.t299 373.214
R110 VDDA.t14 VDDA.t122 373.214
R111 VDDA.t49 VDDA.t14 373.214
R112 VDDA.t124 VDDA.t49 373.214
R113 VDDA.t332 VDDA.t124 373.214
R114 VDDA.t51 VDDA.t329 373.214
R115 VDDA.t374 VDDA.t51 373.214
R116 VDDA.t43 VDDA.t374 373.214
R117 VDDA.t86 VDDA.t43 373.214
R118 VDDA.t80 VDDA.t86 373.214
R119 VDDA.t82 VDDA.t80 373.214
R120 VDDA.t47 VDDA.t82 373.214
R121 VDDA.t32 VDDA.t47 373.214
R122 VDDA.t363 VDDA.t32 373.214
R123 VDDA.t88 VDDA.t293 373.214
R124 VDDA.t376 VDDA.t88 373.214
R125 VDDA.t45 VDDA.t376 373.214
R126 VDDA.t30 VDDA.t45 373.214
R127 VDDA.t256 VDDA.t30 373.214
R128 VDDA.t351 VDDA.t84 373.214
R129 VDDA.t84 VDDA.t76 373.214
R130 VDDA.t76 VDDA.t268 373.214
R131 VDDA.t163 VDDA.t317 373.214
R132 VDDA.t164 VDDA.t163 373.214
R133 VDDA.t354 VDDA.t164 373.214
R134 VDDA.n1980 VDDA.t261 360.868
R135 VDDA.n2005 VDDA.t347 360.868
R136 VDDA.t283 VDDA.n2400 358.858
R137 VDDA.n2406 VDDA.t304 358.858
R138 VDDA.n2409 VDDA.t289 358.858
R139 VDDA.n2413 VDDA.t249 358.858
R140 VDDA.n2195 VDDA.t365 354.154
R141 VDDA.n2194 VDDA.t330 354.154
R142 VDDA.n2177 VDDA.t269 354.154
R143 VDDA.n2178 VDDA.t352 354.154
R144 VDDA.n2410 VDDA.t291 354.065
R145 VDDA.n1961 VDDA.t318 354.063
R146 VDDA.n2401 VDDA.t285 351.793
R147 VDDA.n1962 VDDA.t355 347.224
R148 VDDA.n2819 VDDA.t287 343.882
R149 VDDA.t338 VDDA.n2818 343.882
R150 VDDA.t311 VDDA.n2711 343.882
R151 VDDA.n2712 VDDA.t253 343.882
R152 VDDA.n2214 VDDA.n2184 342.197
R153 VDDA.n2215 VDDA.n2183 342.197
R154 VDDA.n2203 VDDA.n2199 341.769
R155 VDDA.n2204 VDDA.n2198 341.769
R156 VDDA.n2399 VDDA.n2398 338.714
R157 VDDA.n2397 VDDA.n2396 338.714
R158 VDDA.n2395 VDDA.n2394 338.714
R159 VDDA.n2393 VDDA.n2392 338.714
R160 VDDA.n2391 VDDA.n2390 338.714
R161 VDDA.n2389 VDDA.n2388 338.714
R162 VDDA.n2387 VDDA.n2386 338.714
R163 VDDA.n2385 VDDA.n2384 338.714
R164 VDDA.n2381 VDDA.n2380 338.714
R165 VDDA.n2379 VDDA.n2378 338.714
R166 VDDA.n2377 VDDA.n2376 338.714
R167 VDDA.n2375 VDDA.n2374 338.714
R168 VDDA.n2373 VDDA.n2372 338.714
R169 VDDA.n2371 VDDA.n2370 338.714
R170 VDDA.n2369 VDDA.n2368 338.714
R171 VDDA.n2367 VDDA.n2366 338.714
R172 VDDA.n2365 VDDA.n2364 338.714
R173 VDDA.n2362 VDDA.n2361 338.714
R174 VDDA.n2207 VDDA.n2193 336.341
R175 VDDA.n2208 VDDA.n2192 336.341
R176 VDDA.n2209 VDDA.n2191 336.341
R177 VDDA.n2210 VDDA.n2190 336.341
R178 VDDA.n2211 VDDA.n2189 336.341
R179 VDDA.n2181 VDDA.n2180 336.341
R180 VDDA.n2185 VDDA.t294 332.267
R181 VDDA.n2186 VDDA.t257 332.267
R182 VDDA.n2200 VDDA.t300 332.084
R183 VDDA.n2201 VDDA.t333 332.084
R184 VDDA.n2772 VDDA.n2764 291.053
R185 VDDA.n2772 VDDA.n2771 291.053
R186 VDDA.n2769 VDDA.n2762 291.053
R187 VDDA.n2769 VDDA.n2768 291.053
R188 VDDA.n2777 VDDA.n2733 290.233
R189 VDDA.n2778 VDDA.n2733 290.233
R190 VDDA.n2747 VDDA.n2742 290.233
R191 VDDA.n2751 VDDA.n2742 290.233
R192 VDDA.t308 VDDA.n2021 267.188
R193 VDDA.n2027 VDDA.t344 267.188
R194 VDDA.t265 VDDA.t241 259.091
R195 VDDA.t241 VDDA.t280 259.091
R196 VDDA.t61 VDDA.t262 251.471
R197 VDDA.t10 VDDA.t61 251.471
R198 VDDA.t116 VDDA.t10 251.471
R199 VDDA.t215 VDDA.t116 251.471
R200 VDDA.t211 VDDA.t215 251.471
R201 VDDA.t108 VDDA.t211 251.471
R202 VDDA.t100 VDDA.t108 251.471
R203 VDDA.t98 VDDA.t100 251.471
R204 VDDA.t183 VDDA.t98 251.471
R205 VDDA.t59 VDDA.t183 251.471
R206 VDDA.t193 VDDA.t59 251.471
R207 VDDA.t64 VDDA.t193 251.471
R208 VDDA.t103 VDDA.t64 251.471
R209 VDDA.t113 VDDA.t103 251.471
R210 VDDA.t188 VDDA.t113 251.471
R211 VDDA.t165 VDDA.t188 251.471
R212 VDDA.t348 VDDA.t165 251.471
R213 VDDA.n2001 VDDA.n2000 243.698
R214 VDDA.n2026 VDDA.n2025 243.698
R215 VDDA.n2778 VDDA.n2736 242.903
R216 VDDA.n2752 VDDA.n2751 242.903
R217 VDDA.n2029 VDDA.n2028 238.367
R218 VDDA.n2403 VDDA.n2402 238.367
R219 VDDA.n2403 VDDA.n2383 238.367
R220 VDDA.n2774 VDDA.n2773 238.367
R221 VDDA.n2784 VDDA.n2783 238.367
R222 VDDA.n2770 VDDA.n2737 238.367
R223 VDDA.t262 VDDA.n1989 237.5
R224 VDDA.n2002 VDDA.t348 237.5
R225 VDDA.n2782 VDDA.t326 221.121
R226 VDDA.t357 VDDA.n2775 221.121
R227 VDDA.n2775 VDDA.t296 221.121
R228 VDDA.n2753 VDDA.t302 221.121
R229 VDDA.t78 VDDA.t308 217.708
R230 VDDA.t344 VDDA.t78 217.708
R231 VDDA.t287 VDDA.t200 217.708
R232 VDDA.t200 VDDA.t7 217.708
R233 VDDA.t7 VDDA.t206 217.708
R234 VDDA.t206 VDDA.t3 217.708
R235 VDDA.t3 VDDA.t198 217.708
R236 VDDA.t198 VDDA.t22 217.708
R237 VDDA.t22 VDDA.t181 217.708
R238 VDDA.t181 VDDA.t175 217.708
R239 VDDA.t175 VDDA.t180 217.708
R240 VDDA.t180 VDDA.t25 217.708
R241 VDDA.t25 VDDA.t338 217.708
R242 VDDA.t373 VDDA.t311 217.708
R243 VDDA.t168 VDDA.t373 217.708
R244 VDDA.t155 VDDA.t168 217.708
R245 VDDA.t90 VDDA.t155 217.708
R246 VDDA.t177 VDDA.t90 217.708
R247 VDDA.t396 VDDA.t177 217.708
R248 VDDA.t0 VDDA.t396 217.708
R249 VDDA.t63 VDDA.t0 217.708
R250 VDDA.t230 VDDA.t63 217.708
R251 VDDA.t40 VDDA.t230 217.708
R252 VDDA.t253 VDDA.t40 217.708
R253 VDDA.n2732 VDDA.n2731 213.186
R254 VDDA.n2758 VDDA.n2757 213.186
R255 VDDA.t277 VDDA.n2793 213.131
R256 VDDA.n2794 VDDA.t320 213.131
R257 VDDA.t271 VDDA.n2846 213.131
R258 VDDA.n2847 VDDA.t341 213.131
R259 VDDA.t360 VDDA.n2689 213.131
R260 VDDA.n2690 VDDA.t314 213.131
R261 VDDA.n2033 VDDA.n2032 201.169
R262 VDDA.n1988 VDDA.n1987 190.333
R263 VDDA.n2020 VDDA.n2019 190.333
R264 VDDA.n1993 VDDA.n1992 185
R265 VDDA.n1998 VDDA.n1991 185
R266 VDDA.n2002 VDDA.n1991 185
R267 VDDA.n1997 VDDA.n1996 185
R268 VDDA.n1995 VDDA.n1950 185
R269 VDDA.n2004 VDDA.n2003 185
R270 VDDA.n2003 VDDA.n2002 185
R271 VDDA.n1989 VDDA.n1988 185
R272 VDDA.n1986 VDDA.n1954 185
R273 VDDA.n1985 VDDA.n1956 185
R274 VDDA.n1984 VDDA.n1957 185
R275 VDDA.n1959 VDDA.n1958 185
R276 VDDA.n1981 VDDA.n1953 185
R277 VDDA.n1989 VDDA.n1953 185
R278 VDDA.n2024 VDDA.n2022 185
R279 VDDA.n2023 VDDA.n2009 185
R280 VDDA.n2021 VDDA.n2020 185
R281 VDDA.n2018 VDDA.n2012 185
R282 VDDA.n2017 VDDA.n2013 185
R283 VDDA.n2015 VDDA.n2011 185
R284 VDDA.n2021 VDDA.n2011 185
R285 VDDA.n2735 VDDA.n2734 185
R286 VDDA.n2781 VDDA.n2780 185
R287 VDDA.n2782 VDDA.n2781 185
R288 VDDA.n2779 VDDA.n2776 185
R289 VDDA.n2763 VDDA.n2739 185
R290 VDDA.n2767 VDDA.n2738 185
R291 VDDA.n2775 VDDA.n2738 185
R292 VDDA.n2766 VDDA.n2765 185
R293 VDDA.n2755 VDDA.n2754 185
R294 VDDA.n2754 VDDA.n2753 185
R295 VDDA.n2744 VDDA.n2743 185
R296 VDDA.n2749 VDDA.n2748 185
R297 VDDA.n2750 VDDA.n2746 185
R298 VDDA.t326 VDDA.t414 180.173
R299 VDDA.t414 VDDA.t400 180.173
R300 VDDA.t400 VDDA.t196 180.173
R301 VDDA.t196 VDDA.t18 180.173
R302 VDDA.t18 VDDA.t357 180.173
R303 VDDA.t221 VDDA.t296 180.173
R304 VDDA.t383 VDDA.t221 180.173
R305 VDDA.t157 VDDA.t383 180.173
R306 VDDA.t97 VDDA.t157 180.173
R307 VDDA.t302 VDDA.t97 180.173
R308 VDDA.n2801 VDDA.t266 168.139
R309 VDDA.n2800 VDDA.t282 168.139
R310 VDDA.n1948 VDDA.n1947 165.167
R311 VDDA.n1972 VDDA.n1971 165.167
R312 VDDA.n1973 VDDA.n1970 165.167
R313 VDDA.n1974 VDDA.n1969 165.167
R314 VDDA.n1975 VDDA.n1968 165.167
R315 VDDA.n1976 VDDA.n1967 165.167
R316 VDDA.n1977 VDDA.n1966 165.167
R317 VDDA.n1978 VDDA.n1965 165.167
R318 VDDA.n2798 VDDA.n2797 153.576
R319 VDDA.n1992 VDDA.n1991 150
R320 VDDA.n1996 VDDA.n1991 150
R321 VDDA.n2003 VDDA.n1950 150
R322 VDDA.n1988 VDDA.n1954 150
R323 VDDA.n1957 VDDA.n1956 150
R324 VDDA.n1958 VDDA.n1953 150
R325 VDDA.n2022 VDDA.n2009 150
R326 VDDA.n2020 VDDA.n2012 150
R327 VDDA.n2013 VDDA.n2011 150
R328 VDDA.n2739 VDDA.n2738 150
R329 VDDA.n2765 VDDA.n2738 150
R330 VDDA.n2781 VDDA.n2735 150
R331 VDDA.n2781 VDDA.n2776 150
R332 VDDA.n2754 VDDA.n2744 150
R333 VDDA.n2748 VDDA.n2746 150
R334 VDDA.t28 VDDA.t277 146.155
R335 VDDA.t320 VDDA.t28 146.155
R336 VDDA.t34 VDDA.t271 146.155
R337 VDDA.t406 VDDA.t34 146.155
R338 VDDA.t26 VDDA.t406 146.155
R339 VDDA.t132 VDDA.t26 146.155
R340 VDDA.t209 VDDA.t132 146.155
R341 VDDA.t408 VDDA.t209 146.155
R342 VDDA.t391 VDDA.t408 146.155
R343 VDDA.t159 VDDA.t391 146.155
R344 VDDA.t53 VDDA.t159 146.155
R345 VDDA.t143 VDDA.t53 146.155
R346 VDDA.t341 VDDA.t143 146.155
R347 VDDA.t231 VDDA.t360 146.155
R348 VDDA.t235 VDDA.t231 146.155
R349 VDDA.t207 VDDA.t235 146.155
R350 VDDA.t161 VDDA.t207 146.155
R351 VDDA.t55 VDDA.t161 146.155
R352 VDDA.t145 VDDA.t55 146.155
R353 VDDA.t134 VDDA.t145 146.155
R354 VDDA.t233 VDDA.t134 146.155
R355 VDDA.t389 VDDA.t233 146.155
R356 VDDA.t36 VDDA.t389 146.155
R357 VDDA.t314 VDDA.t36 146.155
R358 VDDA.n2819 VDDA.t288 136.701
R359 VDDA.n2818 VDDA.t339 136.701
R360 VDDA.n2711 VDDA.t312 136.701
R361 VDDA.n2712 VDDA.t254 136.701
R362 VDDA.t263 VDDA.n1955 123.126
R363 VDDA.n1983 VDDA.t263 123.126
R364 VDDA.n1999 VDDA.t349 123.126
R365 VDDA.n1994 VDDA.t349 123.126
R366 VDDA.n2835 VDDA.t323 122.829
R367 VDDA.t259 VDDA.n2834 122.829
R368 VDDA.t335 VDDA.n2727 122.829
R369 VDDA.n2728 VDDA.t274 122.829
R370 VDDA.t323 VDDA.t23 81.6411
R371 VDDA.t23 VDDA.t178 81.6411
R372 VDDA.t178 VDDA.t5 81.6411
R373 VDDA.t5 VDDA.t245 81.6411
R374 VDDA.t245 VDDA.t239 81.6411
R375 VDDA.t239 VDDA.t247 81.6411
R376 VDDA.t247 VDDA.t243 81.6411
R377 VDDA.t243 VDDA.t172 81.6411
R378 VDDA.t172 VDDA.t204 81.6411
R379 VDDA.t204 VDDA.t1 81.6411
R380 VDDA.t1 VDDA.t259 81.6411
R381 VDDA.t120 VDDA.t335 81.6411
R382 VDDA.t217 VDDA.t120 81.6411
R383 VDDA.t95 VDDA.t217 81.6411
R384 VDDA.t381 VDDA.t95 81.6411
R385 VDDA.t219 VDDA.t381 81.6411
R386 VDDA.t398 VDDA.t219 81.6411
R387 VDDA.t191 VDDA.t398 81.6411
R388 VDDA.t67 VDDA.t191 81.6411
R389 VDDA.t186 VDDA.t67 81.6411
R390 VDDA.t74 VDDA.t186 81.6411
R391 VDDA.t274 VDDA.t74 81.6411
R392 VDDA.n2793 VDDA.t278 76.2576
R393 VDDA.n2794 VDDA.t321 76.2576
R394 VDDA.n2846 VDDA.t272 76.2576
R395 VDDA.n2847 VDDA.t342 76.2576
R396 VDDA.n2689 VDDA.t361 76.2576
R397 VDDA.n2690 VDDA.t315 76.2576
R398 VDDA.n2791 VDDA.n2790 71.388
R399 VDDA.n2842 VDDA.n2841 71.3255
R400 VDDA.n2844 VDDA.n2843 71.3255
R401 VDDA.n2850 VDDA.n2849 71.3255
R402 VDDA.n2852 VDDA.n2851 71.3255
R403 VDDA.n2685 VDDA.n2684 71.3255
R404 VDDA.n2687 VDDA.n2686 71.3255
R405 VDDA.n2693 VDDA.n2692 71.3255
R406 VDDA.n2695 VDDA.n2694 71.3255
R407 VDDA.n2854 VDDA.n2840 66.8255
R408 VDDA.n2697 VDDA.n2683 66.8255
R409 VDDA.n2002 VDDA.n2001 65.8183
R410 VDDA.n2002 VDDA.n1990 65.8183
R411 VDDA.n1989 VDDA.n1951 65.8183
R412 VDDA.n1989 VDDA.n1952 65.8183
R413 VDDA.n2027 VDDA.n2026 65.8183
R414 VDDA.n2028 VDDA.n2027 65.8183
R415 VDDA.n2021 VDDA.n2010 65.8183
R416 VDDA.n2783 VDDA.n2782 65.8183
R417 VDDA.n2782 VDDA.n2736 65.8183
R418 VDDA.n2775 VDDA.n2774 65.8183
R419 VDDA.n2775 VDDA.n2737 65.8183
R420 VDDA.n2753 VDDA.n2745 65.8183
R421 VDDA.n2753 VDDA.n2752 65.8183
R422 VDDA.n2557 VDDA.t748 59.6762
R423 VDDA.n2558 VDDA.t673 59.6762
R424 VDDA.n1996 VDDA.n1990 53.3664
R425 VDDA.n2001 VDDA.n1992 53.3664
R426 VDDA.n1990 VDDA.n1950 53.3664
R427 VDDA.n1954 VDDA.n1951 53.3664
R428 VDDA.n1957 VDDA.n1952 53.3664
R429 VDDA.n1956 VDDA.n1951 53.3664
R430 VDDA.n1958 VDDA.n1952 53.3664
R431 VDDA.n2026 VDDA.n2022 53.3664
R432 VDDA.n2028 VDDA.n2009 53.3664
R433 VDDA.n2012 VDDA.n2010 53.3664
R434 VDDA.n2013 VDDA.n2010 53.3664
R435 VDDA.n2765 VDDA.n2737 53.3664
R436 VDDA.n2776 VDDA.n2736 53.3664
R437 VDDA.n2783 VDDA.n2735 53.3664
R438 VDDA.n2774 VDDA.n2739 53.3664
R439 VDDA.n2745 VDDA.n2744 53.3664
R440 VDDA.n2752 VDDA.n2746 53.3664
R441 VDDA.n2748 VDDA.n2745 53.3664
R442 VDDA.n2785 VDDA.n2784 51.6576
R443 VDDA.n2756 VDDA.n2755 51.6576
R444 VDDA.n2557 VDDA.t844 51.0443
R445 VDDA.n2559 VDDA.t686 49.1066
R446 VDDA.n2761 VDDA.n2760 48.0005
R447 VDDA.n2761 VDDA.n2740 48.0005
R448 VDDA.n2824 VDDA.n2823 41.1393
R449 VDDA.n2826 VDDA.n2825 41.1393
R450 VDDA.n2828 VDDA.n2827 41.1393
R451 VDDA.n2830 VDDA.n2829 41.1393
R452 VDDA.n2832 VDDA.n2831 41.1393
R453 VDDA.n2717 VDDA.n2716 41.1393
R454 VDDA.n2719 VDDA.n2718 41.1393
R455 VDDA.n2721 VDDA.n2720 41.1393
R456 VDDA.n2723 VDDA.n2722 41.1393
R457 VDDA.n2725 VDDA.n2724 41.1393
R458 VDDA.n2835 VDDA.t324 40.9789
R459 VDDA.n2834 VDDA.t260 40.9789
R460 VDDA.n2727 VDDA.t336 40.9789
R461 VDDA.n2728 VDDA.t275 40.9789
R462 VDDA.n237 VDDA.t73 39.4831
R463 VDDA.n2199 VDDA.t50 39.4005
R464 VDDA.n2199 VDDA.t125 39.4005
R465 VDDA.n2198 VDDA.t123 39.4005
R466 VDDA.n2198 VDDA.t15 39.4005
R467 VDDA.n2193 VDDA.t33 39.4005
R468 VDDA.n2193 VDDA.t364 39.4005
R469 VDDA.n2192 VDDA.t83 39.4005
R470 VDDA.n2192 VDDA.t48 39.4005
R471 VDDA.n2191 VDDA.t87 39.4005
R472 VDDA.n2191 VDDA.t81 39.4005
R473 VDDA.n2190 VDDA.t375 39.4005
R474 VDDA.n2190 VDDA.t44 39.4005
R475 VDDA.t330 VDDA.n2189 39.4005
R476 VDDA.n2189 VDDA.t52 39.4005
R477 VDDA.n2184 VDDA.t46 39.4005
R478 VDDA.n2184 VDDA.t31 39.4005
R479 VDDA.n2183 VDDA.t89 39.4005
R480 VDDA.n2183 VDDA.t377 39.4005
R481 VDDA.n2180 VDDA.t85 39.4005
R482 VDDA.n2180 VDDA.t77 39.4005
R483 VDDA.n2398 VDDA.t154 39.4005
R484 VDDA.n2398 VDDA.t405 39.4005
R485 VDDA.n2396 VDDA.t129 39.4005
R486 VDDA.n2396 VDDA.t137 39.4005
R487 VDDA.n2394 VDDA.t140 39.4005
R488 VDDA.n2394 VDDA.t42 39.4005
R489 VDDA.n2392 VDDA.t142 39.4005
R490 VDDA.n2392 VDDA.t203 39.4005
R491 VDDA.n2390 VDDA.t411 39.4005
R492 VDDA.n2390 VDDA.t92 39.4005
R493 VDDA.n2388 VDDA.t403 39.4005
R494 VDDA.n2388 VDDA.t39 39.4005
R495 VDDA.n2386 VDDA.t170 39.4005
R496 VDDA.n2386 VDDA.t17 39.4005
R497 VDDA.n2384 VDDA.t127 39.4005
R498 VDDA.n2384 VDDA.t94 39.4005
R499 VDDA.n2380 VDDA.t388 39.4005
R500 VDDA.n2380 VDDA.t413 39.4005
R501 VDDA.n2378 VDDA.t225 39.4005
R502 VDDA.n2378 VDDA.t416 39.4005
R503 VDDA.n2376 VDDA.t395 39.4005
R504 VDDA.n2376 VDDA.t223 39.4005
R505 VDDA.n2374 VDDA.t367 39.4005
R506 VDDA.n2374 VDDA.t20 39.4005
R507 VDDA.n2372 VDDA.t72 39.4005
R508 VDDA.n2372 VDDA.t420 39.4005
R509 VDDA.n2370 VDDA.t131 39.4005
R510 VDDA.n2370 VDDA.t150 39.4005
R511 VDDA.n2368 VDDA.t369 39.4005
R512 VDDA.n2368 VDDA.t148 39.4005
R513 VDDA.n2366 VDDA.t70 39.4005
R514 VDDA.n2366 VDDA.t418 39.4005
R515 VDDA.n2364 VDDA.t227 39.4005
R516 VDDA.n2364 VDDA.t386 39.4005
R517 VDDA.n2361 VDDA.t238 39.4005
R518 VDDA.n2361 VDDA.t152 39.4005
R519 VDDA.n2808 VDDA.n2806 30.2463
R520 VDDA.n2701 VDDA.n2699 30.2463
R521 VDDA.n2816 VDDA.n2815 29.6838
R522 VDDA.n2814 VDDA.n2813 29.6838
R523 VDDA.n2812 VDDA.n2811 29.6838
R524 VDDA.n2810 VDDA.n2809 29.6838
R525 VDDA.n2808 VDDA.n2807 29.6838
R526 VDDA.n2709 VDDA.n2708 29.6838
R527 VDDA.n2707 VDDA.n2706 29.6838
R528 VDDA.n2705 VDDA.n2704 29.6838
R529 VDDA.n2703 VDDA.n2702 29.6838
R530 VDDA.n2701 VDDA.n2700 29.6838
R531 VDDA.n2202 VDDA.n2201 27.2462
R532 VDDA.n2200 VDDA.n2197 27.2462
R533 VDDA.n2187 VDDA.n2186 27.2462
R534 VDDA.n2185 VDDA.n2182 27.2462
R535 VDDA.n2196 VDDA.n2195 24.9931
R536 VDDA.n2194 VDDA.n2188 24.9931
R537 VDDA.n2177 VDDA.n2176 24.9931
R538 VDDA.n2179 VDDA.n2178 24.9931
R539 VDDA.n1961 VDDA.n1960 22.9536
R540 VDDA.n2410 VDDA.n2409 22.9536
R541 VDDA.n2005 VDDA.n2004 22.8576
R542 VDDA.n1981 VDDA.n1980 22.8576
R543 VDDA.n2030 VDDA.n2029 22.8576
R544 VDDA.n2015 VDDA.n2014 22.8576
R545 VDDA.n2797 VDDA.t242 21.8894
R546 VDDA.n2797 VDDA.t281 21.8894
R547 VDDA.n2400 VDDA.n2383 20.7243
R548 VDDA.n2406 VDDA.n2382 20.7243
R549 VDDA.n2413 VDDA.n2363 20.7243
R550 VDDA.n1963 VDDA.n1962 20.4312
R551 VDDA.n2032 VDDA.t79 19.7005
R552 VDDA.n2032 VDDA.t345 19.7005
R553 VDDA.n2560 VDDA.n2559 19.1721
R554 VDDA.n2731 VDDA.t401 15.7605
R555 VDDA.n2731 VDDA.t197 15.7605
R556 VDDA.n2757 VDDA.t384 15.7605
R557 VDDA.n2757 VDDA.t158 15.7605
R558 VDDA.n2769 VDDA.t297 15.7605
R559 VDDA.n2772 VDDA.t358 15.7605
R560 VDDA.n2733 VDDA.t327 15.7605
R561 VDDA.n2742 VDDA.t303 15.7605
R562 VDDA.n2758 VDDA.n2756 14.7224
R563 VDDA.n2760 VDDA.n2759 13.8005
R564 VDDA.n2741 VDDA.n2740 13.8005
R565 VDDA.n2786 VDDA.n2785 13.8005
R566 VDDA.n1947 VDDA.t189 13.1338
R567 VDDA.n1947 VDDA.t166 13.1338
R568 VDDA.n1971 VDDA.t104 13.1338
R569 VDDA.n1971 VDDA.t114 13.1338
R570 VDDA.n1970 VDDA.t194 13.1338
R571 VDDA.n1970 VDDA.t65 13.1338
R572 VDDA.n1969 VDDA.t184 13.1338
R573 VDDA.n1969 VDDA.t60 13.1338
R574 VDDA.n1968 VDDA.t101 13.1338
R575 VDDA.n1968 VDDA.t99 13.1338
R576 VDDA.n1967 VDDA.t212 13.1338
R577 VDDA.n1967 VDDA.t109 13.1338
R578 VDDA.n1966 VDDA.t117 13.1338
R579 VDDA.n1966 VDDA.t216 13.1338
R580 VDDA.n1965 VDDA.t62 13.1338
R581 VDDA.n1965 VDDA.t11 13.1338
R582 VDDA.n2822 VDDA.n2816 11.9693
R583 VDDA.n2715 VDDA.n2709 11.9693
R584 VDDA.t278 VDDA.n2791 11.2576
R585 VDDA.n2791 VDDA.t29 11.2576
R586 VDDA.n2841 VDDA.t27 11.2576
R587 VDDA.n2841 VDDA.t133 11.2576
R588 VDDA.n2843 VDDA.t35 11.2576
R589 VDDA.n2843 VDDA.t407 11.2576
R590 VDDA.n2849 VDDA.t54 11.2576
R591 VDDA.n2849 VDDA.t144 11.2576
R592 VDDA.n2851 VDDA.t392 11.2576
R593 VDDA.n2851 VDDA.t160 11.2576
R594 VDDA.n2840 VDDA.t210 11.2576
R595 VDDA.n2840 VDDA.t409 11.2576
R596 VDDA.n2684 VDDA.t208 11.2576
R597 VDDA.n2684 VDDA.t162 11.2576
R598 VDDA.n2686 VDDA.t232 11.2576
R599 VDDA.n2686 VDDA.t236 11.2576
R600 VDDA.n2692 VDDA.t390 11.2576
R601 VDDA.n2692 VDDA.t37 11.2576
R602 VDDA.n2694 VDDA.t135 11.2576
R603 VDDA.n2694 VDDA.t234 11.2576
R604 VDDA.n2683 VDDA.t56 11.2576
R605 VDDA.n2683 VDDA.t146 11.2576
R606 VDDA.n2400 VDDA.n2399 11.2346
R607 VDDA.n1964 VDDA.n1960 11.205
R608 VDDA.n2407 VDDA.n2406 11.1096
R609 VDDA.n2414 VDDA.n2413 11.1096
R610 VDDA.n2409 VDDA.n2408 11.1096
R611 VDDA.n1964 VDDA.n1963 11.0331
R612 VDDA.n2181 VDDA.n2179 10.995
R613 VDDA.n2203 VDDA.n2202 10.9846
R614 VDDA.n2205 VDDA.n2197 10.87
R615 VDDA.n2212 VDDA.n2188 10.87
R616 VDDA.n2216 VDDA.n2182 10.87
R617 VDDA.n2213 VDDA.n2187 10.87
R618 VDDA.n2206 VDDA.n2196 10.87
R619 VDDA.n2031 VDDA.n2030 10.58
R620 VDDA.n1980 VDDA.n1979 10.5331
R621 VDDA.n2014 VDDA.n2007 10.5331
R622 VDDA.n2006 VDDA.n2005 10.5331
R623 VDDA.n2839 VDDA.n2838 10.1567
R624 VDDA.n2789 VDDA.n2788 10.1567
R625 VDDA.n2218 VDDA.n2176 9.42329
R626 VDDA.n1998 VDDA.n1993 9.14336
R627 VDDA.n1998 VDDA.n1997 9.14336
R628 VDDA.n1997 VDDA.n1995 9.14336
R629 VDDA.n1986 VDDA.n1985 9.14336
R630 VDDA.n1985 VDDA.n1984 9.14336
R631 VDDA.n1984 VDDA.n1959 9.14336
R632 VDDA.n2024 VDDA.n2023 9.14336
R633 VDDA.n2018 VDDA.n2017 9.14336
R634 VDDA.n2784 VDDA.n2734 9.14336
R635 VDDA.n2780 VDDA.n2779 9.14336
R636 VDDA.n2755 VDDA.n2743 9.14336
R637 VDDA.n2750 VDDA.n2749 9.14336
R638 VDDA.n2821 VDDA.n2817 8.79217
R639 VDDA.n2714 VDDA.n2710 8.79217
R640 VDDA.n2815 VDDA.t397 8.0005
R641 VDDA.n2815 VDDA.t371 8.0005
R642 VDDA.n2813 VDDA.t171 8.0005
R643 VDDA.n2813 VDDA.t370 8.0005
R644 VDDA.n2811 VDDA.t8 8.0005
R645 VDDA.n2811 VDDA.t201 8.0005
R646 VDDA.n2809 VDDA.t21 8.0005
R647 VDDA.n2809 VDDA.t199 8.0005
R648 VDDA.n2807 VDDA.t174 8.0005
R649 VDDA.n2807 VDDA.t182 8.0005
R650 VDDA.n2806 VDDA.t4 8.0005
R651 VDDA.n2806 VDDA.t111 8.0005
R652 VDDA.n2708 VDDA.t156 8.0005
R653 VDDA.n2708 VDDA.t393 8.0005
R654 VDDA.n2706 VDDA.t138 8.0005
R655 VDDA.n2706 VDDA.t372 8.0005
R656 VDDA.n2704 VDDA.t119 8.0005
R657 VDDA.n2704 VDDA.t13 8.0005
R658 VDDA.n2702 VDDA.t115 8.0005
R659 VDDA.n2702 VDDA.t379 8.0005
R660 VDDA.n2700 VDDA.t176 8.0005
R661 VDDA.n2700 VDDA.t12 8.0005
R662 VDDA.n2699 VDDA.t378 8.0005
R663 VDDA.n2699 VDDA.t380 8.0005
R664 VDDA.n2415 VDDA.n2414 7.55856
R665 VDDA.n2805 VDDA.n2804 7.1255
R666 VDDA.n2838 VDDA.n2822 6.688
R667 VDDA.n2788 VDDA.n2715 6.688
R668 VDDA.n2823 VDDA.t24 6.56717
R669 VDDA.n2823 VDDA.t179 6.56717
R670 VDDA.n2825 VDDA.t6 6.56717
R671 VDDA.n2825 VDDA.t246 6.56717
R672 VDDA.n2827 VDDA.t240 6.56717
R673 VDDA.n2827 VDDA.t248 6.56717
R674 VDDA.n2829 VDDA.t244 6.56717
R675 VDDA.n2829 VDDA.t173 6.56717
R676 VDDA.n2831 VDDA.t205 6.56717
R677 VDDA.n2831 VDDA.t2 6.56717
R678 VDDA.n2716 VDDA.t187 6.56717
R679 VDDA.n2716 VDDA.t75 6.56717
R680 VDDA.n2718 VDDA.t192 6.56717
R681 VDDA.n2718 VDDA.t68 6.56717
R682 VDDA.n2720 VDDA.t220 6.56717
R683 VDDA.n2720 VDDA.t399 6.56717
R684 VDDA.n2722 VDDA.t96 6.56717
R685 VDDA.n2722 VDDA.t382 6.56717
R686 VDDA.n2724 VDDA.t121 6.56717
R687 VDDA.n2724 VDDA.t218 6.56717
R688 VDDA.n2804 VDDA.n2796 6.21925
R689 VDDA.n2838 VDDA.n2837 6.0005
R690 VDDA.n2822 VDDA.n2821 6.0005
R691 VDDA.n2715 VDDA.n2714 6.0005
R692 VDDA.n2850 VDDA.n2848 5.91717
R693 VDDA.n2845 VDDA.n2844 5.91717
R694 VDDA.n2693 VDDA.n2691 5.91717
R695 VDDA.n2688 VDDA.n2687 5.91717
R696 VDDA.n2004 VDDA.n1949 5.33286
R697 VDDA.n1982 VDDA.n1981 5.33286
R698 VDDA.n2029 VDDA.n2008 5.33286
R699 VDDA.n2016 VDDA.n2015 5.33286
R700 VDDA.n2833 VDDA.n2832 5.313
R701 VDDA.n2726 VDDA.n2725 5.313
R702 VDDA.n2804 VDDA.n2803 5.28175
R703 VDDA.n2855 VDDA.n2854 5.21925
R704 VDDA.n2698 VDDA.n2697 5.21925
R705 VDDA.n687 VDDA.t463 4.8295
R706 VDDA.n694 VDDA.t578 4.8295
R707 VDDA.n702 VDDA.t855 4.8295
R708 VDDA.n709 VDDA.t423 4.8295
R709 VDDA.n717 VDDA.t446 4.8295
R710 VDDA.n724 VDDA.t559 4.8295
R711 VDDA.n732 VDDA.t835 4.8295
R712 VDDA.n739 VDDA.t954 4.8295
R713 VDDA.n747 VDDA.t679 4.8295
R714 VDDA.n754 VDDA.t798 4.8295
R715 VDDA.n762 VDDA.t814 4.8295
R716 VDDA.n769 VDDA.t932 4.8295
R717 VDDA.n777 VDDA.t656 4.8295
R718 VDDA.n784 VDDA.t776 4.8295
R719 VDDA.n792 VDDA.t522 4.8295
R720 VDDA.n799 VDDA.t639 4.8295
R721 VDDA.n807 VDDA.t659 4.8295
R722 VDDA.n814 VDDA.t777 4.8295
R723 VDDA.n822 VDDA.t503 4.8295
R724 VDDA.n829 VDDA.t621 4.8295
R725 VDDA.n837 VDDA.t896 4.8295
R726 VDDA.n844 VDDA.t466 4.8295
R727 VDDA.n852 VDDA.t738 4.8295
R728 VDDA.n859 VDDA.t858 4.8295
R729 VDDA.n867 VDDA.t879 4.8295
R730 VDDA.n874 VDDA.t447 4.8295
R731 VDDA.n882 VDDA.t720 4.8295
R732 VDDA.n889 VDDA.t836 4.8295
R733 VDDA.n897 VDDA.t565 4.8295
R734 VDDA.n904 VDDA.t681 4.8295
R735 VDDA.n912 VDDA.t699 4.8295
R736 VDDA.n919 VDDA.t816 4.8295
R737 VDDA.n927 VDDA.t547 4.8295
R738 VDDA.n934 VDDA.t658 4.8295
R739 VDDA.n942 VDDA.t938 4.8295
R740 VDDA.n949 VDDA.t502 4.8295
R741 VDDA.n957 VDDA.t523 4.8295
R742 VDDA.n964 VDDA.t640 4.8295
R743 VDDA.n972 VDDA.t916 4.8295
R744 VDDA.n979 VDDA.t485 4.8295
R745 VDDA.n987 VDDA.t760 4.8295
R746 VDDA.n994 VDDA.t878 4.8295
R747 VDDA.n1002 VDDA.t628 4.8295
R748 VDDA.n1009 VDDA.t741 4.8295
R749 VDDA.n1017 VDDA.t763 4.8295
R750 VDDA.n1024 VDDA.t880 4.8295
R751 VDDA.n1032 VDDA.t608 4.8295
R752 VDDA.n1039 VDDA.t721 4.8295
R753 VDDA.n1047 VDDA.t453 4.8295
R754 VDDA.n1054 VDDA.t567 4.8295
R755 VDDA.n1062 VDDA.t586 4.8295
R756 VDDA.n1069 VDDA.t701 4.8295
R757 VDDA.n1077 VDDA.t433 4.8295
R758 VDDA.n1084 VDDA.t549 4.8295
R759 VDDA.n1092 VDDA.t822 4.8295
R760 VDDA.n1099 VDDA.t942 4.8295
R761 VDDA.n1107 VDDA.t961 4.8295
R762 VDDA.n1114 VDDA.t525 4.8295
R763 VDDA.n1122 VDDA.t805 4.8295
R764 VDDA.n1129 VDDA.t918 4.8295
R765 VDDA.n1137 VDDA.t646 4.8295
R766 VDDA.n1144 VDDA.t762 4.8295
R767 VDDA.n1152 VDDA.t490 4.8295
R768 VDDA.n2821 VDDA.n2820 4.79217
R769 VDDA.n2714 VDDA.n2713 4.79217
R770 VDDA.n2799 VDDA.n2798 4.7505
R771 VDDA.n2792 VDDA.n2790 4.7505
R772 VDDA.n2837 VDDA.n2836 4.7505
R773 VDDA.n2730 VDDA.n2729 4.7505
R774 VDDA.n1496 VDDA.n1330 4.71259
R775 VDDA.n3357 VDDA.n3356 4.71245
R776 VDDA.n2787 VDDA.n2786 4.688
R777 VDDA.n2401 VDDA.n2383 4.54311
R778 VDDA.n2402 VDDA.n2401 4.54311
R779 VDDA.n2777 VDDA.n2734 4.53698
R780 VDDA.n2779 VDDA.n2778 4.53698
R781 VDDA.n2780 VDDA.n2777 4.53698
R782 VDDA.n2747 VDDA.n2743 4.53698
R783 VDDA.n2751 VDDA.n2750 4.53698
R784 VDDA.n2749 VDDA.n2747 4.53698
R785 VDDA.n2220 VDDA.n2219 4.5005
R786 VDDA.n2223 VDDA.n2222 4.5005
R787 VDDA.n2224 VDDA.n2175 4.5005
R788 VDDA.n2228 VDDA.n2225 4.5005
R789 VDDA.n2229 VDDA.n2174 4.5005
R790 VDDA.n2233 VDDA.n2232 4.5005
R791 VDDA.n2234 VDDA.n2173 4.5005
R792 VDDA.n2238 VDDA.n2235 4.5005
R793 VDDA.n2239 VDDA.n2172 4.5005
R794 VDDA.n2243 VDDA.n2242 4.5005
R795 VDDA.n2244 VDDA.n2171 4.5005
R796 VDDA.n2248 VDDA.n2245 4.5005
R797 VDDA.n2249 VDDA.n2170 4.5005
R798 VDDA.n2253 VDDA.n2252 4.5005
R799 VDDA.n2254 VDDA.n2169 4.5005
R800 VDDA.n2258 VDDA.n2255 4.5005
R801 VDDA.n2259 VDDA.n2168 4.5005
R802 VDDA.n2263 VDDA.n2262 4.5005
R803 VDDA.n2264 VDDA.n2167 4.5005
R804 VDDA.n2268 VDDA.n2265 4.5005
R805 VDDA.n2269 VDDA.n2166 4.5005
R806 VDDA.n2273 VDDA.n2272 4.5005
R807 VDDA.n2274 VDDA.n2165 4.5005
R808 VDDA.n2278 VDDA.n2275 4.5005
R809 VDDA.n2279 VDDA.n2164 4.5005
R810 VDDA.n2283 VDDA.n2282 4.5005
R811 VDDA.n2284 VDDA.n2163 4.5005
R812 VDDA.n2288 VDDA.n2285 4.5005
R813 VDDA.n2289 VDDA.n2162 4.5005
R814 VDDA.n2293 VDDA.n2292 4.5005
R815 VDDA.n2294 VDDA.n2161 4.5005
R816 VDDA.n2298 VDDA.n2295 4.5005
R817 VDDA.n2299 VDDA.n2160 4.5005
R818 VDDA.n2303 VDDA.n2302 4.5005
R819 VDDA.n2304 VDDA.n2159 4.5005
R820 VDDA.n2308 VDDA.n2305 4.5005
R821 VDDA.n2309 VDDA.n2158 4.5005
R822 VDDA.n2313 VDDA.n2312 4.5005
R823 VDDA.n2314 VDDA.n2157 4.5005
R824 VDDA.n2318 VDDA.n2315 4.5005
R825 VDDA.n2319 VDDA.n2156 4.5005
R826 VDDA.n2323 VDDA.n2322 4.5005
R827 VDDA.n2324 VDDA.n2155 4.5005
R828 VDDA.n2328 VDDA.n2325 4.5005
R829 VDDA.n2329 VDDA.n2154 4.5005
R830 VDDA.n2333 VDDA.n2332 4.5005
R831 VDDA.n2035 VDDA.n2034 4.5005
R832 VDDA.n2038 VDDA.n2037 4.5005
R833 VDDA.n2039 VDDA.n1946 4.5005
R834 VDDA.n2043 VDDA.n2040 4.5005
R835 VDDA.n2044 VDDA.n1945 4.5005
R836 VDDA.n2048 VDDA.n2047 4.5005
R837 VDDA.n2049 VDDA.n1944 4.5005
R838 VDDA.n2053 VDDA.n2050 4.5005
R839 VDDA.n2054 VDDA.n1943 4.5005
R840 VDDA.n2058 VDDA.n2057 4.5005
R841 VDDA.n2059 VDDA.n1942 4.5005
R842 VDDA.n2063 VDDA.n2060 4.5005
R843 VDDA.n2064 VDDA.n1941 4.5005
R844 VDDA.n2068 VDDA.n2067 4.5005
R845 VDDA.n2069 VDDA.n1940 4.5005
R846 VDDA.n2073 VDDA.n2070 4.5005
R847 VDDA.n2074 VDDA.n1939 4.5005
R848 VDDA.n2078 VDDA.n2077 4.5005
R849 VDDA.n2079 VDDA.n1938 4.5005
R850 VDDA.n2083 VDDA.n2080 4.5005
R851 VDDA.n2084 VDDA.n1937 4.5005
R852 VDDA.n2088 VDDA.n2087 4.5005
R853 VDDA.n2089 VDDA.n1936 4.5005
R854 VDDA.n2093 VDDA.n2090 4.5005
R855 VDDA.n2094 VDDA.n1935 4.5005
R856 VDDA.n2098 VDDA.n2097 4.5005
R857 VDDA.n2099 VDDA.n1934 4.5005
R858 VDDA.n2103 VDDA.n2100 4.5005
R859 VDDA.n2104 VDDA.n1933 4.5005
R860 VDDA.n2108 VDDA.n2107 4.5005
R861 VDDA.n2109 VDDA.n1932 4.5005
R862 VDDA.n2113 VDDA.n2110 4.5005
R863 VDDA.n2114 VDDA.n1931 4.5005
R864 VDDA.n2118 VDDA.n2117 4.5005
R865 VDDA.n2119 VDDA.n1930 4.5005
R866 VDDA.n2123 VDDA.n2120 4.5005
R867 VDDA.n2124 VDDA.n1929 4.5005
R868 VDDA.n2128 VDDA.n2127 4.5005
R869 VDDA.n2129 VDDA.n1928 4.5005
R870 VDDA.n2133 VDDA.n2130 4.5005
R871 VDDA.n2134 VDDA.n1927 4.5005
R872 VDDA.n2138 VDDA.n2137 4.5005
R873 VDDA.n2139 VDDA.n1926 4.5005
R874 VDDA.n2143 VDDA.n2140 4.5005
R875 VDDA.n2144 VDDA.n1925 4.5005
R876 VDDA.n2148 VDDA.n2147 4.5005
R877 VDDA.n238 VDDA.n237 4.5005
R878 VDDA.n241 VDDA.n240 4.5005
R879 VDDA.n242 VDDA.n231 4.5005
R880 VDDA.n246 VDDA.n243 4.5005
R881 VDDA.n247 VDDA.n230 4.5005
R882 VDDA.n251 VDDA.n250 4.5005
R883 VDDA.n252 VDDA.n229 4.5005
R884 VDDA.n256 VDDA.n253 4.5005
R885 VDDA.n257 VDDA.n228 4.5005
R886 VDDA.n261 VDDA.n260 4.5005
R887 VDDA.n262 VDDA.n227 4.5005
R888 VDDA.n266 VDDA.n263 4.5005
R889 VDDA.n267 VDDA.n226 4.5005
R890 VDDA.n271 VDDA.n270 4.5005
R891 VDDA.n272 VDDA.n225 4.5005
R892 VDDA.n276 VDDA.n273 4.5005
R893 VDDA.n277 VDDA.n224 4.5005
R894 VDDA.n281 VDDA.n280 4.5005
R895 VDDA.n282 VDDA.n223 4.5005
R896 VDDA.n286 VDDA.n283 4.5005
R897 VDDA.n287 VDDA.n222 4.5005
R898 VDDA.n291 VDDA.n290 4.5005
R899 VDDA.n292 VDDA.n221 4.5005
R900 VDDA.n296 VDDA.n293 4.5005
R901 VDDA.n297 VDDA.n220 4.5005
R902 VDDA.n301 VDDA.n300 4.5005
R903 VDDA.n302 VDDA.n219 4.5005
R904 VDDA.n306 VDDA.n303 4.5005
R905 VDDA.n307 VDDA.n218 4.5005
R906 VDDA.n311 VDDA.n310 4.5005
R907 VDDA.n312 VDDA.n217 4.5005
R908 VDDA.n316 VDDA.n313 4.5005
R909 VDDA.n317 VDDA.n216 4.5005
R910 VDDA.n321 VDDA.n320 4.5005
R911 VDDA.n322 VDDA.n215 4.5005
R912 VDDA.n326 VDDA.n323 4.5005
R913 VDDA.n327 VDDA.n214 4.5005
R914 VDDA.n331 VDDA.n330 4.5005
R915 VDDA.n332 VDDA.n213 4.5005
R916 VDDA.n336 VDDA.n333 4.5005
R917 VDDA.n337 VDDA.n212 4.5005
R918 VDDA.n341 VDDA.n340 4.5005
R919 VDDA.n342 VDDA.n211 4.5005
R920 VDDA.n346 VDDA.n343 4.5005
R921 VDDA.n347 VDDA.n210 4.5005
R922 VDDA.n351 VDDA.n350 4.5005
R923 VDDA.n2561 VDDA.n2560 4.5005
R924 VDDA.n2564 VDDA.n2563 4.5005
R925 VDDA.n2565 VDDA.n2556 4.5005
R926 VDDA.n2569 VDDA.n2566 4.5005
R927 VDDA.n2570 VDDA.n2555 4.5005
R928 VDDA.n2574 VDDA.n2573 4.5005
R929 VDDA.n2575 VDDA.n2554 4.5005
R930 VDDA.n2579 VDDA.n2576 4.5005
R931 VDDA.n2580 VDDA.n2553 4.5005
R932 VDDA.n2584 VDDA.n2583 4.5005
R933 VDDA.n2585 VDDA.n2552 4.5005
R934 VDDA.n2589 VDDA.n2586 4.5005
R935 VDDA.n2590 VDDA.n2551 4.5005
R936 VDDA.n2594 VDDA.n2593 4.5005
R937 VDDA.n2595 VDDA.n2550 4.5005
R938 VDDA.n2599 VDDA.n2596 4.5005
R939 VDDA.n2600 VDDA.n2549 4.5005
R940 VDDA.n2604 VDDA.n2603 4.5005
R941 VDDA.n2605 VDDA.n2548 4.5005
R942 VDDA.n2609 VDDA.n2606 4.5005
R943 VDDA.n2610 VDDA.n2547 4.5005
R944 VDDA.n2614 VDDA.n2613 4.5005
R945 VDDA.n2615 VDDA.n2546 4.5005
R946 VDDA.n2619 VDDA.n2616 4.5005
R947 VDDA.n2620 VDDA.n2545 4.5005
R948 VDDA.n2624 VDDA.n2623 4.5005
R949 VDDA.n2625 VDDA.n2544 4.5005
R950 VDDA.n2629 VDDA.n2626 4.5005
R951 VDDA.n2630 VDDA.n2543 4.5005
R952 VDDA.n2634 VDDA.n2633 4.5005
R953 VDDA.n2635 VDDA.n2542 4.5005
R954 VDDA.n2639 VDDA.n2636 4.5005
R955 VDDA.n2640 VDDA.n2541 4.5005
R956 VDDA.n2644 VDDA.n2643 4.5005
R957 VDDA.n2645 VDDA.n2540 4.5005
R958 VDDA.n2649 VDDA.n2646 4.5005
R959 VDDA.n2650 VDDA.n2539 4.5005
R960 VDDA.n2654 VDDA.n2653 4.5005
R961 VDDA.n2655 VDDA.n2538 4.5005
R962 VDDA.n2659 VDDA.n2656 4.5005
R963 VDDA.n2660 VDDA.n2537 4.5005
R964 VDDA.n2664 VDDA.n2663 4.5005
R965 VDDA.n2665 VDDA.n2536 4.5005
R966 VDDA.n2669 VDDA.n2666 4.5005
R967 VDDA.n2670 VDDA.n2535 4.5005
R968 VDDA.n2674 VDDA.n2673 4.5005
R969 VDDA.n2416 VDDA.n2415 4.5005
R970 VDDA.n2419 VDDA.n2418 4.5005
R971 VDDA.n2420 VDDA.n2360 4.5005
R972 VDDA.n2424 VDDA.n2421 4.5005
R973 VDDA.n2425 VDDA.n2359 4.5005
R974 VDDA.n2429 VDDA.n2428 4.5005
R975 VDDA.n2430 VDDA.n2358 4.5005
R976 VDDA.n2434 VDDA.n2431 4.5005
R977 VDDA.n2435 VDDA.n2357 4.5005
R978 VDDA.n2439 VDDA.n2438 4.5005
R979 VDDA.n2440 VDDA.n2356 4.5005
R980 VDDA.n2444 VDDA.n2441 4.5005
R981 VDDA.n2445 VDDA.n2355 4.5005
R982 VDDA.n2449 VDDA.n2448 4.5005
R983 VDDA.n2450 VDDA.n2354 4.5005
R984 VDDA.n2454 VDDA.n2451 4.5005
R985 VDDA.n2455 VDDA.n2353 4.5005
R986 VDDA.n2459 VDDA.n2458 4.5005
R987 VDDA.n2460 VDDA.n2352 4.5005
R988 VDDA.n2464 VDDA.n2461 4.5005
R989 VDDA.n2465 VDDA.n2351 4.5005
R990 VDDA.n2469 VDDA.n2468 4.5005
R991 VDDA.n2470 VDDA.n2350 4.5005
R992 VDDA.n2474 VDDA.n2471 4.5005
R993 VDDA.n2475 VDDA.n2349 4.5005
R994 VDDA.n2479 VDDA.n2478 4.5005
R995 VDDA.n2480 VDDA.n2348 4.5005
R996 VDDA.n2484 VDDA.n2481 4.5005
R997 VDDA.n2485 VDDA.n2347 4.5005
R998 VDDA.n2489 VDDA.n2488 4.5005
R999 VDDA.n2490 VDDA.n2346 4.5005
R1000 VDDA.n2494 VDDA.n2491 4.5005
R1001 VDDA.n2495 VDDA.n2345 4.5005
R1002 VDDA.n2499 VDDA.n2498 4.5005
R1003 VDDA.n2500 VDDA.n2344 4.5005
R1004 VDDA.n2504 VDDA.n2501 4.5005
R1005 VDDA.n2505 VDDA.n2343 4.5005
R1006 VDDA.n2509 VDDA.n2508 4.5005
R1007 VDDA.n2510 VDDA.n2342 4.5005
R1008 VDDA.n2514 VDDA.n2511 4.5005
R1009 VDDA.n2515 VDDA.n2341 4.5005
R1010 VDDA.n2519 VDDA.n2518 4.5005
R1011 VDDA.n2520 VDDA.n2340 4.5005
R1012 VDDA.n2524 VDDA.n2521 4.5005
R1013 VDDA.n2525 VDDA.n2339 4.5005
R1014 VDDA.n2529 VDDA.n2528 4.5005
R1015 VDDA.n91 VDDA.n85 4.5005
R1016 VDDA.n93 VDDA.n92 4.5005
R1017 VDDA.n94 VDDA.n84 4.5005
R1018 VDDA.n98 VDDA.n97 4.5005
R1019 VDDA.n99 VDDA.n81 4.5005
R1020 VDDA.n101 VDDA.n100 4.5005
R1021 VDDA.n102 VDDA.n80 4.5005
R1022 VDDA.n106 VDDA.n105 4.5005
R1023 VDDA.n107 VDDA.n77 4.5005
R1024 VDDA.n109 VDDA.n108 4.5005
R1025 VDDA.n110 VDDA.n76 4.5005
R1026 VDDA.n114 VDDA.n113 4.5005
R1027 VDDA.n115 VDDA.n73 4.5005
R1028 VDDA.n117 VDDA.n116 4.5005
R1029 VDDA.n118 VDDA.n72 4.5005
R1030 VDDA.n122 VDDA.n121 4.5005
R1031 VDDA.n123 VDDA.n69 4.5005
R1032 VDDA.n125 VDDA.n124 4.5005
R1033 VDDA.n126 VDDA.n68 4.5005
R1034 VDDA.n130 VDDA.n129 4.5005
R1035 VDDA.n131 VDDA.n65 4.5005
R1036 VDDA.n133 VDDA.n132 4.5005
R1037 VDDA.n134 VDDA.n64 4.5005
R1038 VDDA.n138 VDDA.n137 4.5005
R1039 VDDA.n139 VDDA.n61 4.5005
R1040 VDDA.n141 VDDA.n140 4.5005
R1041 VDDA.n142 VDDA.n60 4.5005
R1042 VDDA.n146 VDDA.n145 4.5005
R1043 VDDA.n147 VDDA.n57 4.5005
R1044 VDDA.n149 VDDA.n148 4.5005
R1045 VDDA.n150 VDDA.n56 4.5005
R1046 VDDA.n154 VDDA.n153 4.5005
R1047 VDDA.n155 VDDA.n53 4.5005
R1048 VDDA.n157 VDDA.n156 4.5005
R1049 VDDA.n158 VDDA.n52 4.5005
R1050 VDDA.n162 VDDA.n161 4.5005
R1051 VDDA.n163 VDDA.n49 4.5005
R1052 VDDA.n165 VDDA.n164 4.5005
R1053 VDDA.n166 VDDA.n48 4.5005
R1054 VDDA.n170 VDDA.n169 4.5005
R1055 VDDA.n171 VDDA.n45 4.5005
R1056 VDDA.n173 VDDA.n172 4.5005
R1057 VDDA.n174 VDDA.n44 4.5005
R1058 VDDA.n178 VDDA.n177 4.5005
R1059 VDDA.n179 VDDA.n43 4.5005
R1060 VDDA.n3358 VDDA.n3357 4.5005
R1061 VDDA.n3236 VDDA.n3235 4.5005
R1062 VDDA.n3246 VDDA.n3245 4.5005
R1063 VDDA.n3247 VDDA.n3234 4.5005
R1064 VDDA.n3249 VDDA.n3248 4.5005
R1065 VDDA.n3232 VDDA.n3231 4.5005
R1066 VDDA.n3256 VDDA.n3255 4.5005
R1067 VDDA.n3257 VDDA.n3230 4.5005
R1068 VDDA.n3259 VDDA.n3258 4.5005
R1069 VDDA.n3228 VDDA.n3227 4.5005
R1070 VDDA.n3266 VDDA.n3265 4.5005
R1071 VDDA.n3267 VDDA.n3226 4.5005
R1072 VDDA.n3269 VDDA.n3268 4.5005
R1073 VDDA.n3224 VDDA.n3223 4.5005
R1074 VDDA.n3276 VDDA.n3275 4.5005
R1075 VDDA.n3277 VDDA.n3222 4.5005
R1076 VDDA.n3279 VDDA.n3278 4.5005
R1077 VDDA.n3220 VDDA.n3219 4.5005
R1078 VDDA.n3286 VDDA.n3285 4.5005
R1079 VDDA.n3287 VDDA.n3218 4.5005
R1080 VDDA.n3289 VDDA.n3288 4.5005
R1081 VDDA.n3216 VDDA.n3215 4.5005
R1082 VDDA.n3296 VDDA.n3295 4.5005
R1083 VDDA.n3297 VDDA.n3214 4.5005
R1084 VDDA.n3299 VDDA.n3298 4.5005
R1085 VDDA.n3212 VDDA.n3211 4.5005
R1086 VDDA.n3306 VDDA.n3305 4.5005
R1087 VDDA.n3307 VDDA.n3210 4.5005
R1088 VDDA.n3309 VDDA.n3308 4.5005
R1089 VDDA.n3208 VDDA.n3207 4.5005
R1090 VDDA.n3316 VDDA.n3315 4.5005
R1091 VDDA.n3317 VDDA.n3206 4.5005
R1092 VDDA.n3319 VDDA.n3318 4.5005
R1093 VDDA.n3204 VDDA.n3203 4.5005
R1094 VDDA.n3326 VDDA.n3325 4.5005
R1095 VDDA.n3327 VDDA.n3202 4.5005
R1096 VDDA.n3329 VDDA.n3328 4.5005
R1097 VDDA.n3200 VDDA.n3199 4.5005
R1098 VDDA.n3336 VDDA.n3335 4.5005
R1099 VDDA.n3337 VDDA.n3198 4.5005
R1100 VDDA.n3339 VDDA.n3338 4.5005
R1101 VDDA.n3196 VDDA.n3195 4.5005
R1102 VDDA.n3346 VDDA.n3345 4.5005
R1103 VDDA.n3347 VDDA.n3194 4.5005
R1104 VDDA.n3349 VDDA.n3348 4.5005
R1105 VDDA.n3192 VDDA.n3191 4.5005
R1106 VDDA.n3355 VDDA.n3354 4.5005
R1107 VDDA.n3096 VDDA.n3092 4.5005
R1108 VDDA.n3100 VDDA.n3099 4.5005
R1109 VDDA.n3101 VDDA.n3089 4.5005
R1110 VDDA.n3103 VDDA.n3102 4.5005
R1111 VDDA.n3104 VDDA.n3088 4.5005
R1112 VDDA.n3108 VDDA.n3107 4.5005
R1113 VDDA.n3109 VDDA.n3085 4.5005
R1114 VDDA.n3111 VDDA.n3110 4.5005
R1115 VDDA.n3112 VDDA.n3084 4.5005
R1116 VDDA.n3116 VDDA.n3115 4.5005
R1117 VDDA.n3117 VDDA.n3081 4.5005
R1118 VDDA.n3119 VDDA.n3118 4.5005
R1119 VDDA.n3120 VDDA.n3080 4.5005
R1120 VDDA.n3124 VDDA.n3123 4.5005
R1121 VDDA.n3125 VDDA.n3077 4.5005
R1122 VDDA.n3127 VDDA.n3126 4.5005
R1123 VDDA.n3128 VDDA.n3076 4.5005
R1124 VDDA.n3132 VDDA.n3131 4.5005
R1125 VDDA.n3133 VDDA.n3073 4.5005
R1126 VDDA.n3135 VDDA.n3134 4.5005
R1127 VDDA.n3136 VDDA.n3072 4.5005
R1128 VDDA.n3140 VDDA.n3139 4.5005
R1129 VDDA.n3141 VDDA.n3069 4.5005
R1130 VDDA.n3143 VDDA.n3142 4.5005
R1131 VDDA.n3144 VDDA.n3068 4.5005
R1132 VDDA.n3148 VDDA.n3147 4.5005
R1133 VDDA.n3149 VDDA.n3065 4.5005
R1134 VDDA.n3151 VDDA.n3150 4.5005
R1135 VDDA.n3152 VDDA.n3064 4.5005
R1136 VDDA.n3156 VDDA.n3155 4.5005
R1137 VDDA.n3157 VDDA.n3061 4.5005
R1138 VDDA.n3159 VDDA.n3158 4.5005
R1139 VDDA.n3160 VDDA.n3060 4.5005
R1140 VDDA.n3164 VDDA.n3163 4.5005
R1141 VDDA.n3165 VDDA.n3057 4.5005
R1142 VDDA.n3167 VDDA.n3166 4.5005
R1143 VDDA.n3168 VDDA.n3056 4.5005
R1144 VDDA.n3172 VDDA.n3171 4.5005
R1145 VDDA.n3173 VDDA.n3053 4.5005
R1146 VDDA.n3175 VDDA.n3174 4.5005
R1147 VDDA.n3176 VDDA.n3052 4.5005
R1148 VDDA.n3180 VDDA.n3179 4.5005
R1149 VDDA.n3181 VDDA.n3051 4.5005
R1150 VDDA.n3183 VDDA.n3182 4.5005
R1151 VDDA.n182 VDDA.n181 4.5005
R1152 VDDA.n3189 VDDA.n3188 4.5005
R1153 VDDA.n2934 VDDA.n2928 4.5005
R1154 VDDA.n2936 VDDA.n2935 4.5005
R1155 VDDA.n2937 VDDA.n2927 4.5005
R1156 VDDA.n2941 VDDA.n2940 4.5005
R1157 VDDA.n2942 VDDA.n2924 4.5005
R1158 VDDA.n2944 VDDA.n2943 4.5005
R1159 VDDA.n2945 VDDA.n2923 4.5005
R1160 VDDA.n2949 VDDA.n2948 4.5005
R1161 VDDA.n2950 VDDA.n2920 4.5005
R1162 VDDA.n2952 VDDA.n2951 4.5005
R1163 VDDA.n2953 VDDA.n2919 4.5005
R1164 VDDA.n2957 VDDA.n2956 4.5005
R1165 VDDA.n2958 VDDA.n2916 4.5005
R1166 VDDA.n2960 VDDA.n2959 4.5005
R1167 VDDA.n2961 VDDA.n2915 4.5005
R1168 VDDA.n2965 VDDA.n2964 4.5005
R1169 VDDA.n2966 VDDA.n2912 4.5005
R1170 VDDA.n2968 VDDA.n2967 4.5005
R1171 VDDA.n2969 VDDA.n2911 4.5005
R1172 VDDA.n2973 VDDA.n2972 4.5005
R1173 VDDA.n2974 VDDA.n2908 4.5005
R1174 VDDA.n2976 VDDA.n2975 4.5005
R1175 VDDA.n2977 VDDA.n2907 4.5005
R1176 VDDA.n2981 VDDA.n2980 4.5005
R1177 VDDA.n2982 VDDA.n2904 4.5005
R1178 VDDA.n2984 VDDA.n2983 4.5005
R1179 VDDA.n2985 VDDA.n2903 4.5005
R1180 VDDA.n2989 VDDA.n2988 4.5005
R1181 VDDA.n2990 VDDA.n2900 4.5005
R1182 VDDA.n2992 VDDA.n2991 4.5005
R1183 VDDA.n2993 VDDA.n2899 4.5005
R1184 VDDA.n2997 VDDA.n2996 4.5005
R1185 VDDA.n2998 VDDA.n2896 4.5005
R1186 VDDA.n3000 VDDA.n2999 4.5005
R1187 VDDA.n3001 VDDA.n2895 4.5005
R1188 VDDA.n3005 VDDA.n3004 4.5005
R1189 VDDA.n3006 VDDA.n2892 4.5005
R1190 VDDA.n3008 VDDA.n3007 4.5005
R1191 VDDA.n3009 VDDA.n2891 4.5005
R1192 VDDA.n3013 VDDA.n3012 4.5005
R1193 VDDA.n3014 VDDA.n2888 4.5005
R1194 VDDA.n3016 VDDA.n3015 4.5005
R1195 VDDA.n3017 VDDA.n2887 4.5005
R1196 VDDA.n3021 VDDA.n3020 4.5005
R1197 VDDA.n3022 VDDA.n2886 4.5005
R1198 VDDA.n3024 VDDA.n3023 4.5005
R1199 VDDA.n428 VDDA.n422 4.5005
R1200 VDDA.n430 VDDA.n429 4.5005
R1201 VDDA.n431 VDDA.n421 4.5005
R1202 VDDA.n435 VDDA.n434 4.5005
R1203 VDDA.n436 VDDA.n418 4.5005
R1204 VDDA.n438 VDDA.n437 4.5005
R1205 VDDA.n439 VDDA.n417 4.5005
R1206 VDDA.n443 VDDA.n442 4.5005
R1207 VDDA.n444 VDDA.n414 4.5005
R1208 VDDA.n446 VDDA.n445 4.5005
R1209 VDDA.n447 VDDA.n413 4.5005
R1210 VDDA.n451 VDDA.n450 4.5005
R1211 VDDA.n452 VDDA.n410 4.5005
R1212 VDDA.n454 VDDA.n453 4.5005
R1213 VDDA.n455 VDDA.n409 4.5005
R1214 VDDA.n459 VDDA.n458 4.5005
R1215 VDDA.n460 VDDA.n406 4.5005
R1216 VDDA.n462 VDDA.n461 4.5005
R1217 VDDA.n463 VDDA.n405 4.5005
R1218 VDDA.n467 VDDA.n466 4.5005
R1219 VDDA.n468 VDDA.n402 4.5005
R1220 VDDA.n470 VDDA.n469 4.5005
R1221 VDDA.n471 VDDA.n401 4.5005
R1222 VDDA.n475 VDDA.n474 4.5005
R1223 VDDA.n476 VDDA.n398 4.5005
R1224 VDDA.n478 VDDA.n477 4.5005
R1225 VDDA.n479 VDDA.n397 4.5005
R1226 VDDA.n483 VDDA.n482 4.5005
R1227 VDDA.n484 VDDA.n394 4.5005
R1228 VDDA.n486 VDDA.n485 4.5005
R1229 VDDA.n487 VDDA.n393 4.5005
R1230 VDDA.n491 VDDA.n490 4.5005
R1231 VDDA.n492 VDDA.n390 4.5005
R1232 VDDA.n494 VDDA.n493 4.5005
R1233 VDDA.n495 VDDA.n389 4.5005
R1234 VDDA.n499 VDDA.n498 4.5005
R1235 VDDA.n500 VDDA.n386 4.5005
R1236 VDDA.n502 VDDA.n501 4.5005
R1237 VDDA.n503 VDDA.n385 4.5005
R1238 VDDA.n507 VDDA.n506 4.5005
R1239 VDDA.n508 VDDA.n382 4.5005
R1240 VDDA.n510 VDDA.n509 4.5005
R1241 VDDA.n511 VDDA.n381 4.5005
R1242 VDDA.n515 VDDA.n514 4.5005
R1243 VDDA.n516 VDDA.n380 4.5005
R1244 VDDA.n2858 VDDA.n2857 4.5005
R1245 VDDA.n1737 VDDA.n1733 4.5005
R1246 VDDA.n1741 VDDA.n1740 4.5005
R1247 VDDA.n1742 VDDA.n1730 4.5005
R1248 VDDA.n1744 VDDA.n1743 4.5005
R1249 VDDA.n1745 VDDA.n1729 4.5005
R1250 VDDA.n1749 VDDA.n1748 4.5005
R1251 VDDA.n1750 VDDA.n1726 4.5005
R1252 VDDA.n1752 VDDA.n1751 4.5005
R1253 VDDA.n1753 VDDA.n1725 4.5005
R1254 VDDA.n1757 VDDA.n1756 4.5005
R1255 VDDA.n1758 VDDA.n1722 4.5005
R1256 VDDA.n1760 VDDA.n1759 4.5005
R1257 VDDA.n1761 VDDA.n1721 4.5005
R1258 VDDA.n1765 VDDA.n1764 4.5005
R1259 VDDA.n1766 VDDA.n1718 4.5005
R1260 VDDA.n1768 VDDA.n1767 4.5005
R1261 VDDA.n1769 VDDA.n1717 4.5005
R1262 VDDA.n1773 VDDA.n1772 4.5005
R1263 VDDA.n1774 VDDA.n1714 4.5005
R1264 VDDA.n1776 VDDA.n1775 4.5005
R1265 VDDA.n1777 VDDA.n1713 4.5005
R1266 VDDA.n1781 VDDA.n1780 4.5005
R1267 VDDA.n1782 VDDA.n1710 4.5005
R1268 VDDA.n1784 VDDA.n1783 4.5005
R1269 VDDA.n1785 VDDA.n1709 4.5005
R1270 VDDA.n1789 VDDA.n1788 4.5005
R1271 VDDA.n1790 VDDA.n1706 4.5005
R1272 VDDA.n1792 VDDA.n1791 4.5005
R1273 VDDA.n1793 VDDA.n1705 4.5005
R1274 VDDA.n1797 VDDA.n1796 4.5005
R1275 VDDA.n1798 VDDA.n1702 4.5005
R1276 VDDA.n1800 VDDA.n1799 4.5005
R1277 VDDA.n1801 VDDA.n1701 4.5005
R1278 VDDA.n1805 VDDA.n1804 4.5005
R1279 VDDA.n1806 VDDA.n1698 4.5005
R1280 VDDA.n1808 VDDA.n1807 4.5005
R1281 VDDA.n1809 VDDA.n1697 4.5005
R1282 VDDA.n1813 VDDA.n1812 4.5005
R1283 VDDA.n1814 VDDA.n1694 4.5005
R1284 VDDA.n1816 VDDA.n1815 4.5005
R1285 VDDA.n1817 VDDA.n1693 4.5005
R1286 VDDA.n1821 VDDA.n1820 4.5005
R1287 VDDA.n1822 VDDA.n1692 4.5005
R1288 VDDA.n1824 VDDA.n1823 4.5005
R1289 VDDA.n519 VDDA.n518 4.5005
R1290 VDDA.n2681 VDDA.n2680 4.5005
R1291 VDDA.n2803 VDDA.n2802 4.5005
R1292 VDDA.n2796 VDDA.n2795 4.5005
R1293 VDDA.n2854 VDDA.n2853 4.5005
R1294 VDDA.n2788 VDDA.n2787 4.5005
R1295 VDDA.n2697 VDDA.n2696 4.5005
R1296 VDDA.n1575 VDDA.n1569 4.5005
R1297 VDDA.n1577 VDDA.n1576 4.5005
R1298 VDDA.n1578 VDDA.n1568 4.5005
R1299 VDDA.n1582 VDDA.n1581 4.5005
R1300 VDDA.n1583 VDDA.n1565 4.5005
R1301 VDDA.n1585 VDDA.n1584 4.5005
R1302 VDDA.n1586 VDDA.n1564 4.5005
R1303 VDDA.n1590 VDDA.n1589 4.5005
R1304 VDDA.n1591 VDDA.n1561 4.5005
R1305 VDDA.n1593 VDDA.n1592 4.5005
R1306 VDDA.n1594 VDDA.n1560 4.5005
R1307 VDDA.n1598 VDDA.n1597 4.5005
R1308 VDDA.n1599 VDDA.n1557 4.5005
R1309 VDDA.n1601 VDDA.n1600 4.5005
R1310 VDDA.n1602 VDDA.n1556 4.5005
R1311 VDDA.n1606 VDDA.n1605 4.5005
R1312 VDDA.n1607 VDDA.n1553 4.5005
R1313 VDDA.n1609 VDDA.n1608 4.5005
R1314 VDDA.n1610 VDDA.n1552 4.5005
R1315 VDDA.n1614 VDDA.n1613 4.5005
R1316 VDDA.n1615 VDDA.n1549 4.5005
R1317 VDDA.n1617 VDDA.n1616 4.5005
R1318 VDDA.n1618 VDDA.n1548 4.5005
R1319 VDDA.n1622 VDDA.n1621 4.5005
R1320 VDDA.n1623 VDDA.n1545 4.5005
R1321 VDDA.n1625 VDDA.n1624 4.5005
R1322 VDDA.n1626 VDDA.n1544 4.5005
R1323 VDDA.n1630 VDDA.n1629 4.5005
R1324 VDDA.n1631 VDDA.n1541 4.5005
R1325 VDDA.n1633 VDDA.n1632 4.5005
R1326 VDDA.n1634 VDDA.n1540 4.5005
R1327 VDDA.n1638 VDDA.n1637 4.5005
R1328 VDDA.n1639 VDDA.n1537 4.5005
R1329 VDDA.n1641 VDDA.n1640 4.5005
R1330 VDDA.n1642 VDDA.n1536 4.5005
R1331 VDDA.n1646 VDDA.n1645 4.5005
R1332 VDDA.n1647 VDDA.n1533 4.5005
R1333 VDDA.n1649 VDDA.n1648 4.5005
R1334 VDDA.n1650 VDDA.n1532 4.5005
R1335 VDDA.n1654 VDDA.n1653 4.5005
R1336 VDDA.n1655 VDDA.n1529 4.5005
R1337 VDDA.n1657 VDDA.n1656 4.5005
R1338 VDDA.n1658 VDDA.n1528 4.5005
R1339 VDDA.n1662 VDDA.n1661 4.5005
R1340 VDDA.n1663 VDDA.n1527 4.5005
R1341 VDDA.n1665 VDDA.n1664 4.5005
R1342 VDDA.n595 VDDA.n589 4.5005
R1343 VDDA.n597 VDDA.n596 4.5005
R1344 VDDA.n598 VDDA.n588 4.5005
R1345 VDDA.n602 VDDA.n601 4.5005
R1346 VDDA.n603 VDDA.n585 4.5005
R1347 VDDA.n605 VDDA.n604 4.5005
R1348 VDDA.n606 VDDA.n584 4.5005
R1349 VDDA.n610 VDDA.n609 4.5005
R1350 VDDA.n611 VDDA.n581 4.5005
R1351 VDDA.n613 VDDA.n612 4.5005
R1352 VDDA.n614 VDDA.n580 4.5005
R1353 VDDA.n618 VDDA.n617 4.5005
R1354 VDDA.n619 VDDA.n577 4.5005
R1355 VDDA.n621 VDDA.n620 4.5005
R1356 VDDA.n622 VDDA.n576 4.5005
R1357 VDDA.n626 VDDA.n625 4.5005
R1358 VDDA.n627 VDDA.n573 4.5005
R1359 VDDA.n629 VDDA.n628 4.5005
R1360 VDDA.n630 VDDA.n572 4.5005
R1361 VDDA.n634 VDDA.n633 4.5005
R1362 VDDA.n635 VDDA.n569 4.5005
R1363 VDDA.n637 VDDA.n636 4.5005
R1364 VDDA.n638 VDDA.n568 4.5005
R1365 VDDA.n642 VDDA.n641 4.5005
R1366 VDDA.n643 VDDA.n565 4.5005
R1367 VDDA.n645 VDDA.n644 4.5005
R1368 VDDA.n646 VDDA.n564 4.5005
R1369 VDDA.n650 VDDA.n649 4.5005
R1370 VDDA.n651 VDDA.n561 4.5005
R1371 VDDA.n653 VDDA.n652 4.5005
R1372 VDDA.n654 VDDA.n560 4.5005
R1373 VDDA.n658 VDDA.n657 4.5005
R1374 VDDA.n659 VDDA.n557 4.5005
R1375 VDDA.n661 VDDA.n660 4.5005
R1376 VDDA.n662 VDDA.n556 4.5005
R1377 VDDA.n666 VDDA.n665 4.5005
R1378 VDDA.n667 VDDA.n553 4.5005
R1379 VDDA.n669 VDDA.n668 4.5005
R1380 VDDA.n670 VDDA.n552 4.5005
R1381 VDDA.n674 VDDA.n673 4.5005
R1382 VDDA.n675 VDDA.n549 4.5005
R1383 VDDA.n677 VDDA.n676 4.5005
R1384 VDDA.n678 VDDA.n548 4.5005
R1385 VDDA.n682 VDDA.n681 4.5005
R1386 VDDA.n683 VDDA.n547 4.5005
R1387 VDDA.n1499 VDDA.n1498 4.5005
R1388 VDDA.n1376 VDDA.n1375 4.5005
R1389 VDDA.n1386 VDDA.n1385 4.5005
R1390 VDDA.n1387 VDDA.n1374 4.5005
R1391 VDDA.n1389 VDDA.n1388 4.5005
R1392 VDDA.n1372 VDDA.n1371 4.5005
R1393 VDDA.n1396 VDDA.n1395 4.5005
R1394 VDDA.n1397 VDDA.n1370 4.5005
R1395 VDDA.n1399 VDDA.n1398 4.5005
R1396 VDDA.n1368 VDDA.n1367 4.5005
R1397 VDDA.n1406 VDDA.n1405 4.5005
R1398 VDDA.n1407 VDDA.n1366 4.5005
R1399 VDDA.n1409 VDDA.n1408 4.5005
R1400 VDDA.n1364 VDDA.n1363 4.5005
R1401 VDDA.n1416 VDDA.n1415 4.5005
R1402 VDDA.n1417 VDDA.n1362 4.5005
R1403 VDDA.n1419 VDDA.n1418 4.5005
R1404 VDDA.n1360 VDDA.n1359 4.5005
R1405 VDDA.n1426 VDDA.n1425 4.5005
R1406 VDDA.n1427 VDDA.n1358 4.5005
R1407 VDDA.n1429 VDDA.n1428 4.5005
R1408 VDDA.n1356 VDDA.n1355 4.5005
R1409 VDDA.n1436 VDDA.n1435 4.5005
R1410 VDDA.n1437 VDDA.n1354 4.5005
R1411 VDDA.n1439 VDDA.n1438 4.5005
R1412 VDDA.n1352 VDDA.n1351 4.5005
R1413 VDDA.n1446 VDDA.n1445 4.5005
R1414 VDDA.n1447 VDDA.n1350 4.5005
R1415 VDDA.n1449 VDDA.n1448 4.5005
R1416 VDDA.n1348 VDDA.n1347 4.5005
R1417 VDDA.n1456 VDDA.n1455 4.5005
R1418 VDDA.n1457 VDDA.n1346 4.5005
R1419 VDDA.n1459 VDDA.n1458 4.5005
R1420 VDDA.n1344 VDDA.n1343 4.5005
R1421 VDDA.n1466 VDDA.n1465 4.5005
R1422 VDDA.n1467 VDDA.n1342 4.5005
R1423 VDDA.n1469 VDDA.n1468 4.5005
R1424 VDDA.n1340 VDDA.n1339 4.5005
R1425 VDDA.n1476 VDDA.n1475 4.5005
R1426 VDDA.n1477 VDDA.n1338 4.5005
R1427 VDDA.n1479 VDDA.n1478 4.5005
R1428 VDDA.n1336 VDDA.n1335 4.5005
R1429 VDDA.n1486 VDDA.n1485 4.5005
R1430 VDDA.n1487 VDDA.n1334 4.5005
R1431 VDDA.n1489 VDDA.n1488 4.5005
R1432 VDDA.n1332 VDDA.n1331 4.5005
R1433 VDDA.n1495 VDDA.n1494 4.5005
R1434 VDDA.n1217 VDDA.n1213 4.5005
R1435 VDDA.n1221 VDDA.n1220 4.5005
R1436 VDDA.n1222 VDDA.n1212 4.5005
R1437 VDDA.n1226 VDDA.n1223 4.5005
R1438 VDDA.n1227 VDDA.n1211 4.5005
R1439 VDDA.n1231 VDDA.n1230 4.5005
R1440 VDDA.n1232 VDDA.n1210 4.5005
R1441 VDDA.n1236 VDDA.n1233 4.5005
R1442 VDDA.n1237 VDDA.n1209 4.5005
R1443 VDDA.n1241 VDDA.n1240 4.5005
R1444 VDDA.n1242 VDDA.n1208 4.5005
R1445 VDDA.n1246 VDDA.n1243 4.5005
R1446 VDDA.n1247 VDDA.n1207 4.5005
R1447 VDDA.n1251 VDDA.n1250 4.5005
R1448 VDDA.n1252 VDDA.n1206 4.5005
R1449 VDDA.n1256 VDDA.n1253 4.5005
R1450 VDDA.n1257 VDDA.n1205 4.5005
R1451 VDDA.n1261 VDDA.n1260 4.5005
R1452 VDDA.n1262 VDDA.n1204 4.5005
R1453 VDDA.n1266 VDDA.n1263 4.5005
R1454 VDDA.n1267 VDDA.n1203 4.5005
R1455 VDDA.n1271 VDDA.n1270 4.5005
R1456 VDDA.n1272 VDDA.n1202 4.5005
R1457 VDDA.n1276 VDDA.n1273 4.5005
R1458 VDDA.n1277 VDDA.n1201 4.5005
R1459 VDDA.n1281 VDDA.n1280 4.5005
R1460 VDDA.n1282 VDDA.n1200 4.5005
R1461 VDDA.n1286 VDDA.n1283 4.5005
R1462 VDDA.n1287 VDDA.n1199 4.5005
R1463 VDDA.n1291 VDDA.n1290 4.5005
R1464 VDDA.n1292 VDDA.n1198 4.5005
R1465 VDDA.n1296 VDDA.n1293 4.5005
R1466 VDDA.n1297 VDDA.n1197 4.5005
R1467 VDDA.n1301 VDDA.n1300 4.5005
R1468 VDDA.n1302 VDDA.n1196 4.5005
R1469 VDDA.n1306 VDDA.n1303 4.5005
R1470 VDDA.n1307 VDDA.n1195 4.5005
R1471 VDDA.n1311 VDDA.n1310 4.5005
R1472 VDDA.n1312 VDDA.n1194 4.5005
R1473 VDDA.n1316 VDDA.n1313 4.5005
R1474 VDDA.n1317 VDDA.n1193 4.5005
R1475 VDDA.n1321 VDDA.n1320 4.5005
R1476 VDDA.n1322 VDDA.n1192 4.5005
R1477 VDDA.n1324 VDDA.n1323 4.5005
R1478 VDDA.n685 VDDA.n684 4.5005
R1479 VDDA.n1330 VDDA.n1329 4.5005
R1480 VDDA.n687 VDDA.t551 4.5005
R1481 VDDA.n688 VDDA.t952 4.5005
R1482 VDDA.n689 VDDA.t801 4.5005
R1483 VDDA.n690 VDDA.t887 4.5005
R1484 VDDA.n691 VDDA.t735 4.5005
R1485 VDDA.n692 VDDA.t590 4.5005
R1486 VDDA.n693 VDDA.t674 4.5005
R1487 VDDA.n701 VDDA.t526 4.5005
R1488 VDDA.n700 VDDA.t928 4.5005
R1489 VDDA.n699 VDDA.t782 4.5005
R1490 VDDA.n698 VDDA.t866 4.5005
R1491 VDDA.n697 VDDA.t715 4.5005
R1492 VDDA.n696 VDDA.t792 4.5005
R1493 VDDA.n695 VDDA.t877 4.5005
R1494 VDDA.n694 VDDA.t727 4.5005
R1495 VDDA.n702 VDDA.t943 4.5005
R1496 VDDA.n703 VDDA.t796 4.5005
R1497 VDDA.n704 VDDA.t643 4.5005
R1498 VDDA.n705 VDDA.t728 4.5005
R1499 VDDA.n706 VDDA.t580 4.5005
R1500 VDDA.n707 VDDA.t434 4.5005
R1501 VDDA.n708 VDDA.t516 4.5005
R1502 VDDA.n716 VDDA.t919 4.5005
R1503 VDDA.n715 VDDA.t772 4.5005
R1504 VDDA.n714 VDDA.t623 4.5005
R1505 VDDA.n713 VDDA.t708 4.5005
R1506 VDDA.n712 VDDA.t560 4.5005
R1507 VDDA.n711 VDDA.t633 4.5005
R1508 VDDA.n710 VDDA.t719 4.5005
R1509 VDDA.n709 VDDA.t571 4.5005
R1510 VDDA.n717 VDDA.t529 4.5005
R1511 VDDA.n718 VDDA.t931 4.5005
R1512 VDDA.n719 VDDA.t784 4.5005
R1513 VDDA.n720 VDDA.t867 4.5005
R1514 VDDA.n721 VDDA.t718 4.5005
R1515 VDDA.n722 VDDA.t569 4.5005
R1516 VDDA.n723 VDDA.t652 4.5005
R1517 VDDA.n731 VDDA.t505 4.5005
R1518 VDDA.n730 VDDA.t906 4.5005
R1519 VDDA.n729 VDDA.t758 4.5005
R1520 VDDA.n728 VDDA.t845 4.5005
R1521 VDDA.n727 VDDA.t695 4.5005
R1522 VDDA.n726 VDDA.t770 4.5005
R1523 VDDA.n725 VDDA.t857 4.5005
R1524 VDDA.n724 VDDA.t707 4.5005
R1525 VDDA.n732 VDDA.t920 4.5005
R1526 VDDA.n733 VDDA.t775 4.5005
R1527 VDDA.n734 VDDA.t626 4.5005
R1528 VDDA.n735 VDDA.t709 4.5005
R1529 VDDA.n736 VDDA.t563 4.5005
R1530 VDDA.n737 VDDA.t963 4.5005
R1531 VDDA.n738 VDDA.t496 4.5005
R1532 VDDA.n746 VDDA.t899 4.5005
R1533 VDDA.n745 VDDA.t750 4.5005
R1534 VDDA.n744 VDDA.t603 4.5005
R1535 VDDA.n743 VDDA.t688 4.5005
R1536 VDDA.n742 VDDA.t541 4.5005
R1537 VDDA.n741 VDDA.t614 4.5005
R1538 VDDA.n740 VDDA.t698 4.5005
R1539 VDDA.n739 VDDA.t553 4.5005
R1540 VDDA.n747 VDDA.t764 4.5005
R1541 VDDA.n748 VDDA.t619 4.5005
R1542 VDDA.n749 VDDA.t471 4.5005
R1543 VDDA.n750 VDDA.t555 4.5005
R1544 VDDA.n751 VDDA.t958 4.5005
R1545 VDDA.n752 VDDA.t807 4.5005
R1546 VDDA.n753 VDDA.t892 4.5005
R1547 VDDA.n761 VDDA.t743 4.5005
R1548 VDDA.n760 VDDA.t596 4.5005
R1549 VDDA.n759 VDDA.t448 4.5005
R1550 VDDA.n758 VDDA.t534 4.5005
R1551 VDDA.n757 VDDA.t933 4.5005
R1552 VDDA.n756 VDDA.t459 4.5005
R1553 VDDA.n755 VDDA.t546 4.5005
R1554 VDDA.n754 VDDA.t946 4.5005
R1555 VDDA.n762 VDDA.t901 4.5005
R1556 VDDA.n763 VDDA.t752 4.5005
R1557 VDDA.n764 VDDA.t605 4.5005
R1558 VDDA.n765 VDDA.t690 4.5005
R1559 VDDA.n766 VDDA.t544 4.5005
R1560 VDDA.n767 VDDA.t947 4.5005
R1561 VDDA.n768 VDDA.t481 4.5005
R1562 VDDA.n776 VDDA.t881 4.5005
R1563 VDDA.n775 VDDA.t730 4.5005
R1564 VDDA.n774 VDDA.t583 4.5005
R1565 VDDA.n773 VDDA.t666 4.5005
R1566 VDDA.n772 VDDA.t517 4.5005
R1567 VDDA.n771 VDDA.t594 4.5005
R1568 VDDA.n770 VDDA.t680 4.5005
R1569 VDDA.n769 VDDA.t533 4.5005
R1570 VDDA.n777 VDDA.t744 4.5005
R1571 VDDA.n778 VDDA.t598 4.5005
R1572 VDDA.n779 VDDA.t450 4.5005
R1573 VDDA.n780 VDDA.t535 4.5005
R1574 VDDA.n781 VDDA.t936 4.5005
R1575 VDDA.n782 VDDA.t787 4.5005
R1576 VDDA.n783 VDDA.t872 4.5005
R1577 VDDA.n791 VDDA.t722 4.5005
R1578 VDDA.n790 VDDA.t573 4.5005
R1579 VDDA.n789 VDDA.t427 4.5005
R1580 VDDA.n788 VDDA.t509 4.5005
R1581 VDDA.n787 VDDA.t909 4.5005
R1582 VDDA.n786 VDDA.t439 4.5005
R1583 VDDA.n785 VDDA.t520 4.5005
R1584 VDDA.n784 VDDA.t923 4.5005
R1585 VDDA.n792 VDDA.t610 4.5005
R1586 VDDA.n793 VDDA.t464 4.5005
R1587 VDDA.n794 VDDA.t863 4.5005
R1588 VDDA.n795 VDDA.t950 4.5005
R1589 VDDA.n796 VDDA.t802 4.5005
R1590 VDDA.n797 VDDA.t649 4.5005
R1591 VDDA.n798 VDDA.t733 4.5005
R1592 VDDA.n806 VDDA.t587 4.5005
R1593 VDDA.n805 VDDA.t443 4.5005
R1594 VDDA.n804 VDDA.t838 4.5005
R1595 VDDA.n803 VDDA.t926 4.5005
R1596 VDDA.n802 VDDA.t780 4.5005
R1597 VDDA.n801 VDDA.t850 4.5005
R1598 VDDA.n800 VDDA.t940 4.5005
R1599 VDDA.n799 VDDA.t790 4.5005
R1600 VDDA.n807 VDDA.t746 4.5005
R1601 VDDA.n808 VDDA.t599 4.5005
R1602 VDDA.n809 VDDA.t452 4.5005
R1603 VDDA.n810 VDDA.t537 4.5005
R1604 VDDA.n811 VDDA.t937 4.5005
R1605 VDDA.n812 VDDA.t791 4.5005
R1606 VDDA.n813 VDDA.t874 4.5005
R1607 VDDA.n821 VDDA.t723 4.5005
R1608 VDDA.n820 VDDA.t577 4.5005
R1609 VDDA.n819 VDDA.t431 4.5005
R1610 VDDA.n818 VDDA.t510 4.5005
R1611 VDDA.n817 VDDA.t914 4.5005
R1612 VDDA.n816 VDDA.t440 4.5005
R1613 VDDA.n815 VDDA.t524 4.5005
R1614 VDDA.n814 VDDA.t925 4.5005
R1615 VDDA.n822 VDDA.t591 4.5005
R1616 VDDA.n823 VDDA.t445 4.5005
R1617 VDDA.n824 VDDA.t842 4.5005
R1618 VDDA.n825 VDDA.t929 4.5005
R1619 VDDA.n826 VDDA.t783 4.5005
R1620 VDDA.n827 VDDA.t632 4.5005
R1621 VDDA.n828 VDDA.t716 4.5005
R1622 VDDA.n836 VDDA.t568 4.5005
R1623 VDDA.n835 VDDA.t422 4.5005
R1624 VDDA.n834 VDDA.t821 4.5005
R1625 VDDA.n833 VDDA.t905 4.5005
R1626 VDDA.n832 VDDA.t757 4.5005
R1627 VDDA.n831 VDDA.t830 4.5005
R1628 VDDA.n830 VDDA.t917 4.5005
R1629 VDDA.n829 VDDA.t769 4.5005
R1630 VDDA.n837 VDDA.t436 4.5005
R1631 VDDA.n838 VDDA.t834 4.5005
R1632 VDDA.n839 VDDA.t684 4.5005
R1633 VDDA.n840 VDDA.t773 4.5005
R1634 VDDA.n841 VDDA.t624 4.5005
R1635 VDDA.n842 VDDA.t476 4.5005
R1636 VDDA.n843 VDDA.t561 4.5005
R1637 VDDA.n851 VDDA.t962 4.5005
R1638 VDDA.n850 VDDA.t813 4.5005
R1639 VDDA.n849 VDDA.t663 4.5005
R1640 VDDA.n848 VDDA.t749 4.5005
R1641 VDDA.n847 VDDA.t602 4.5005
R1642 VDDA.n846 VDDA.t670 4.5005
R1643 VDDA.n845 VDDA.t761 4.5005
R1644 VDDA.n844 VDDA.t613 4.5005
R1645 VDDA.n852 VDDA.t825 4.5005
R1646 VDDA.n853 VDDA.t677 4.5005
R1647 VDDA.n854 VDDA.t530 4.5005
R1648 VDDA.n855 VDDA.t616 4.5005
R1649 VDDA.n856 VDDA.t468 4.5005
R1650 VDDA.n857 VDDA.t869 4.5005
R1651 VDDA.n858 VDDA.t956 4.5005
R1652 VDDA.n866 VDDA.t806 4.5005
R1653 VDDA.n865 VDDA.t655 4.5005
R1654 VDDA.n864 VDDA.t506 4.5005
R1655 VDDA.n863 VDDA.t595 4.5005
R1656 VDDA.n862 VDDA.t449 4.5005
R1657 VDDA.n861 VDDA.t514 4.5005
R1658 VDDA.n860 VDDA.t606 4.5005
R1659 VDDA.n859 VDDA.t458 4.5005
R1660 VDDA.n867 VDDA.t965 4.5005
R1661 VDDA.n868 VDDA.t815 4.5005
R1662 VDDA.n869 VDDA.t664 4.5005
R1663 VDDA.n870 VDDA.t751 4.5005
R1664 VDDA.n871 VDDA.t604 4.5005
R1665 VDDA.n872 VDDA.t457 4.5005
R1666 VDDA.n873 VDDA.t542 4.5005
R1667 VDDA.n881 VDDA.t944 4.5005
R1668 VDDA.n880 VDDA.t797 4.5005
R1669 VDDA.n879 VDDA.t645 4.5005
R1670 VDDA.n878 VDDA.t729 4.5005
R1671 VDDA.n877 VDDA.t581 4.5005
R1672 VDDA.n876 VDDA.t653 4.5005
R1673 VDDA.n875 VDDA.t740 4.5005
R1674 VDDA.n874 VDDA.t593 4.5005
R1675 VDDA.n882 VDDA.t809 4.5005
R1676 VDDA.n883 VDDA.t657 4.5005
R1677 VDDA.n884 VDDA.t507 4.5005
R1678 VDDA.n885 VDDA.t597 4.5005
R1679 VDDA.n886 VDDA.t451 4.5005
R1680 VDDA.n887 VDDA.t847 4.5005
R1681 VDDA.n888 VDDA.t934 4.5005
R1682 VDDA.n896 VDDA.t786 4.5005
R1683 VDDA.n895 VDDA.t636 4.5005
R1684 VDDA.n894 VDDA.t488 4.5005
R1685 VDDA.n893 VDDA.t572 4.5005
R1686 VDDA.n892 VDDA.t426 4.5005
R1687 VDDA.n891 VDDA.t497 4.5005
R1688 VDDA.n890 VDDA.t585 4.5005
R1689 VDDA.n889 VDDA.t438 4.5005
R1690 VDDA.n897 VDDA.t647 4.5005
R1691 VDDA.n898 VDDA.t500 4.5005
R1692 VDDA.n899 VDDA.t902 4.5005
R1693 VDDA.n900 VDDA.t441 4.5005
R1694 VDDA.n901 VDDA.t839 4.5005
R1695 VDDA.n902 VDDA.t691 4.5005
R1696 VDDA.n903 VDDA.t778 4.5005
R1697 VDDA.n911 VDDA.t630 4.5005
R1698 VDDA.n910 VDDA.t482 4.5005
R1699 VDDA.n909 VDDA.t883 4.5005
R1700 VDDA.n908 VDDA.t968 4.5005
R1701 VDDA.n907 VDDA.t818 4.5005
R1702 VDDA.n906 VDDA.t893 4.5005
R1703 VDDA.n905 VDDA.t432 4.5005
R1704 VDDA.n904 VDDA.t828 4.5005
R1705 VDDA.n912 VDDA.t788 4.5005
R1706 VDDA.n913 VDDA.t638 4.5005
R1707 VDDA.n914 VDDA.t491 4.5005
R1708 VDDA.n915 VDDA.t575 4.5005
R1709 VDDA.n916 VDDA.t429 4.5005
R1710 VDDA.n917 VDDA.t829 4.5005
R1711 VDDA.n918 VDDA.t912 4.5005
R1712 VDDA.n926 VDDA.t765 4.5005
R1713 VDDA.n925 VDDA.t620 4.5005
R1714 VDDA.n924 VDDA.t472 4.5005
R1715 VDDA.n923 VDDA.t556 4.5005
R1716 VDDA.n922 VDDA.t959 4.5005
R1717 VDDA.n921 VDDA.t479 4.5005
R1718 VDDA.n920 VDDA.t566 4.5005
R1719 VDDA.n919 VDDA.t967 4.5005
R1720 VDDA.n927 VDDA.t631 4.5005
R1721 VDDA.n928 VDDA.t484 4.5005
R1722 VDDA.n929 VDDA.t885 4.5005
R1723 VDDA.n930 VDDA.t421 4.5005
R1724 VDDA.n931 VDDA.t820 4.5005
R1725 VDDA.n932 VDDA.t668 4.5005
R1726 VDDA.n933 VDDA.t756 4.5005
R1727 VDDA.n941 VDDA.t609 4.5005
R1728 VDDA.n940 VDDA.t461 4.5005
R1729 VDDA.n939 VDDA.t861 4.5005
R1730 VDDA.n938 VDDA.t949 4.5005
R1731 VDDA.n937 VDDA.t799 4.5005
R1732 VDDA.n936 VDDA.t871 4.5005
R1733 VDDA.n935 VDDA.t960 4.5005
R1734 VDDA.n934 VDDA.t810 4.5005
R1735 VDDA.n942 VDDA.t474 4.5005
R1736 VDDA.n943 VDDA.t875 4.5005
R1737 VDDA.n944 VDDA.t724 4.5005
R1738 VDDA.n945 VDDA.t811 4.5005
R1739 VDDA.n946 VDDA.t661 4.5005
R1740 VDDA.n947 VDDA.t512 4.5005
R1741 VDDA.n948 VDDA.t601 4.5005
R1742 VDDA.n956 VDDA.t455 4.5005
R1743 VDDA.n955 VDDA.t853 4.5005
R1744 VDDA.n954 VDDA.t704 4.5005
R1745 VDDA.n953 VDDA.t793 4.5005
R1746 VDDA.n952 VDDA.t641 4.5005
R1747 VDDA.n951 VDDA.t714 4.5005
R1748 VDDA.n950 VDDA.t804 4.5005
R1749 VDDA.n949 VDDA.t651 4.5005
R1750 VDDA.n957 VDDA.t611 4.5005
R1751 VDDA.n958 VDDA.t465 4.5005
R1752 VDDA.n959 VDDA.t864 4.5005
R1753 VDDA.n960 VDDA.t951 4.5005
R1754 VDDA.n961 VDDA.t803 4.5005
R1755 VDDA.n962 VDDA.t650 4.5005
R1756 VDDA.n963 VDDA.t736 4.5005
R1757 VDDA.n971 VDDA.t588 4.5005
R1758 VDDA.n970 VDDA.t444 4.5005
R1759 VDDA.n969 VDDA.t841 4.5005
R1760 VDDA.n968 VDDA.t927 4.5005
R1761 VDDA.n967 VDDA.t781 4.5005
R1762 VDDA.n966 VDDA.t851 4.5005
R1763 VDDA.n965 VDDA.t941 4.5005
R1764 VDDA.n964 VDDA.t794 4.5005
R1765 VDDA.n972 VDDA.t456 4.5005
R1766 VDDA.n973 VDDA.t856 4.5005
R1767 VDDA.n974 VDDA.t706 4.5005
R1768 VDDA.n975 VDDA.t795 4.5005
R1769 VDDA.n976 VDDA.t644 4.5005
R1770 VDDA.n977 VDDA.t494 4.5005
R1771 VDDA.n978 VDDA.t582 4.5005
R1772 VDDA.n986 VDDA.t435 4.5005
R1773 VDDA.n985 VDDA.t832 4.5005
R1774 VDDA.n984 VDDA.t683 4.5005
R1775 VDDA.n983 VDDA.t771 4.5005
R1776 VDDA.n982 VDDA.t622 4.5005
R1777 VDDA.n981 VDDA.t694 4.5005
R1778 VDDA.n980 VDDA.t785 4.5005
R1779 VDDA.n979 VDDA.t634 4.5005
R1780 VDDA.n987 VDDA.t846 4.5005
R1781 VDDA.n988 VDDA.t697 4.5005
R1782 VDDA.n989 VDDA.t552 4.5005
R1783 VDDA.n990 VDDA.t635 4.5005
R1784 VDDA.n991 VDDA.t487 4.5005
R1785 VDDA.n992 VDDA.t888 4.5005
R1786 VDDA.n993 VDDA.t424 4.5005
R1787 VDDA.n1001 VDDA.t824 4.5005
R1788 VDDA.n1000 VDDA.t675 4.5005
R1789 VDDA.n999 VDDA.t528 4.5005
R1790 VDDA.n998 VDDA.t615 4.5005
R1791 VDDA.n997 VDDA.t467 4.5005
R1792 VDDA.n996 VDDA.t540 4.5005
R1793 VDDA.n995 VDDA.t627 4.5005
R1794 VDDA.n994 VDDA.t477 4.5005
R1795 VDDA.n1002 VDDA.t711 4.5005
R1796 VDDA.n1003 VDDA.t564 4.5005
R1797 VDDA.n1004 VDDA.t966 4.5005
R1798 VDDA.n1005 VDDA.t499 4.5005
R1799 VDDA.n1006 VDDA.t900 4.5005
R1800 VDDA.n1007 VDDA.t753 4.5005
R1801 VDDA.n1008 VDDA.t837 4.5005
R1802 VDDA.n1016 VDDA.t689 4.5005
R1803 VDDA.n1015 VDDA.t545 4.5005
R1804 VDDA.n1014 VDDA.t945 4.5005
R1805 VDDA.n1013 VDDA.t480 4.5005
R1806 VDDA.n1012 VDDA.t882 4.5005
R1807 VDDA.n1011 VDDA.t955 4.5005
R1808 VDDA.n1010 VDDA.t492 4.5005
R1809 VDDA.n1009 VDDA.t891 4.5005
R1810 VDDA.n1017 VDDA.t848 4.5005
R1811 VDDA.n1018 VDDA.t700 4.5005
R1812 VDDA.n1019 VDDA.t554 4.5005
R1813 VDDA.n1020 VDDA.t637 4.5005
R1814 VDDA.n1021 VDDA.t489 4.5005
R1815 VDDA.n1022 VDDA.t890 4.5005
R1816 VDDA.n1023 VDDA.t428 4.5005
R1817 VDDA.n1031 VDDA.t826 4.5005
R1818 VDDA.n1030 VDDA.t678 4.5005
R1819 VDDA.n1029 VDDA.t532 4.5005
R1820 VDDA.n1028 VDDA.t617 4.5005
R1821 VDDA.n1027 VDDA.t469 4.5005
R1822 VDDA.n1026 VDDA.t543 4.5005
R1823 VDDA.n1025 VDDA.t629 4.5005
R1824 VDDA.n1024 VDDA.t478 4.5005
R1825 VDDA.n1032 VDDA.t692 4.5005
R1826 VDDA.n1033 VDDA.t548 4.5005
R1827 VDDA.n1034 VDDA.t948 4.5005
R1828 VDDA.n1035 VDDA.t483 4.5005
R1829 VDDA.n1036 VDDA.t884 4.5005
R1830 VDDA.n1037 VDDA.t732 4.5005
R1831 VDDA.n1038 VDDA.t819 4.5005
R1832 VDDA.n1046 VDDA.t667 4.5005
R1833 VDDA.n1045 VDDA.t519 4.5005
R1834 VDDA.n1044 VDDA.t922 4.5005
R1835 VDDA.n1043 VDDA.t460 4.5005
R1836 VDDA.n1042 VDDA.t859 4.5005
R1837 VDDA.n1041 VDDA.t935 4.5005
R1838 VDDA.n1040 VDDA.t473 4.5005
R1839 VDDA.n1039 VDDA.t870 4.5005
R1840 VDDA.n1047 VDDA.t536 4.5005
R1841 VDDA.n1048 VDDA.t939 4.5005
R1842 VDDA.n1049 VDDA.t789 4.5005
R1843 VDDA.n1050 VDDA.t873 4.5005
R1844 VDDA.n1051 VDDA.t725 4.5005
R1845 VDDA.n1052 VDDA.t576 4.5005
R1846 VDDA.n1053 VDDA.t660 4.5005
R1847 VDDA.n1061 VDDA.t511 4.5005
R1848 VDDA.n1060 VDDA.t913 4.5005
R1849 VDDA.n1059 VDDA.t767 4.5005
R1850 VDDA.n1058 VDDA.t852 4.5005
R1851 VDDA.n1057 VDDA.t703 4.5005
R1852 VDDA.n1056 VDDA.t779 4.5005
R1853 VDDA.n1055 VDDA.t865 4.5005
R1854 VDDA.n1054 VDDA.t712 4.5005
R1855 VDDA.n1062 VDDA.t669 4.5005
R1856 VDDA.n1063 VDDA.t521 4.5005
R1857 VDDA.n1064 VDDA.t924 4.5005
R1858 VDDA.n1065 VDDA.t462 4.5005
R1859 VDDA.n1066 VDDA.t862 4.5005
R1860 VDDA.n1067 VDDA.t713 4.5005
R1861 VDDA.n1068 VDDA.t800 4.5005
R1862 VDDA.n1076 VDDA.t648 4.5005
R1863 VDDA.n1075 VDDA.t501 4.5005
R1864 VDDA.n1074 VDDA.t903 4.5005
R1865 VDDA.n1073 VDDA.t442 4.5005
R1866 VDDA.n1072 VDDA.t840 4.5005
R1867 VDDA.n1071 VDDA.t910 4.5005
R1868 VDDA.n1070 VDDA.t454 4.5005
R1869 VDDA.n1069 VDDA.t849 4.5005
R1870 VDDA.n1077 VDDA.t513 4.5005
R1871 VDDA.n1078 VDDA.t915 4.5005
R1872 VDDA.n1079 VDDA.t768 4.5005
R1873 VDDA.n1080 VDDA.t854 4.5005
R1874 VDDA.n1081 VDDA.t705 4.5005
R1875 VDDA.n1082 VDDA.t558 4.5005
R1876 VDDA.n1083 VDDA.t642 4.5005
R1877 VDDA.n1091 VDDA.t493 4.5005
R1878 VDDA.n1090 VDDA.t895 4.5005
R1879 VDDA.n1089 VDDA.t745 4.5005
R1880 VDDA.n1088 VDDA.t831 4.5005
R1881 VDDA.n1087 VDDA.t682 4.5005
R1882 VDDA.n1086 VDDA.t755 4.5005
R1883 VDDA.n1085 VDDA.t843 4.5005
R1884 VDDA.n1084 VDDA.t693 4.5005
R1885 VDDA.n1092 VDDA.t907 4.5005
R1886 VDDA.n1093 VDDA.t759 4.5005
R1887 VDDA.n1094 VDDA.t612 4.5005
R1888 VDDA.n1095 VDDA.t696 4.5005
R1889 VDDA.n1096 VDDA.t550 4.5005
R1890 VDDA.n1097 VDDA.t953 4.5005
R1891 VDDA.n1098 VDDA.t486 4.5005
R1892 VDDA.n1106 VDDA.t886 4.5005
R1893 VDDA.n1105 VDDA.t737 4.5005
R1894 VDDA.n1104 VDDA.t589 4.5005
R1895 VDDA.n1103 VDDA.t672 4.5005
R1896 VDDA.n1102 VDDA.t527 4.5005
R1897 VDDA.n1101 VDDA.t600 4.5005
R1898 VDDA.n1100 VDDA.t687 4.5005
R1899 VDDA.n1099 VDDA.t539 4.5005
R1900 VDDA.n1107 VDDA.t495 4.5005
R1901 VDDA.n1108 VDDA.t897 4.5005
R1902 VDDA.n1109 VDDA.t747 4.5005
R1903 VDDA.n1110 VDDA.t833 4.5005
R1904 VDDA.n1111 VDDA.t685 4.5005
R1905 VDDA.n1112 VDDA.t538 4.5005
R1906 VDDA.n1113 VDDA.t625 4.5005
R1907 VDDA.n1121 VDDA.t475 4.5005
R1908 VDDA.n1120 VDDA.t876 4.5005
R1909 VDDA.n1119 VDDA.t726 4.5005
R1910 VDDA.n1118 VDDA.t812 4.5005
R1911 VDDA.n1117 VDDA.t662 4.5005
R1912 VDDA.n1116 VDDA.t734 4.5005
R1913 VDDA.n1115 VDDA.t823 4.5005
R1914 VDDA.n1114 VDDA.t671 4.5005
R1915 VDDA.n1122 VDDA.t889 4.5005
R1916 VDDA.n1123 VDDA.t739 4.5005
R1917 VDDA.n1124 VDDA.t592 4.5005
R1918 VDDA.n1125 VDDA.t676 4.5005
R1919 VDDA.n1126 VDDA.t531 4.5005
R1920 VDDA.n1127 VDDA.t930 4.5005
R1921 VDDA.n1128 VDDA.t470 4.5005
R1922 VDDA.n1136 VDDA.t868 4.5005
R1923 VDDA.n1135 VDDA.t717 4.5005
R1924 VDDA.n1134 VDDA.t570 4.5005
R1925 VDDA.n1133 VDDA.t654 4.5005
R1926 VDDA.n1132 VDDA.t504 4.5005
R1927 VDDA.n1131 VDDA.t579 4.5005
R1928 VDDA.n1130 VDDA.t665 4.5005
R1929 VDDA.n1129 VDDA.t515 4.5005
R1930 VDDA.n1137 VDDA.t731 4.5005
R1931 VDDA.n1138 VDDA.t584 4.5005
R1932 VDDA.n1139 VDDA.t437 4.5005
R1933 VDDA.n1140 VDDA.t518 4.5005
R1934 VDDA.n1141 VDDA.t921 4.5005
R1935 VDDA.n1142 VDDA.t774 4.5005
R1936 VDDA.n1143 VDDA.t860 4.5005
R1937 VDDA.n1151 VDDA.t710 4.5005
R1938 VDDA.n1150 VDDA.t562 4.5005
R1939 VDDA.n1149 VDDA.t964 4.5005
R1940 VDDA.n1148 VDDA.t498 4.5005
R1941 VDDA.n1147 VDDA.t898 4.5005
R1942 VDDA.n1146 VDDA.t425 4.5005
R1943 VDDA.n1145 VDDA.t508 4.5005
R1944 VDDA.n1144 VDDA.t908 4.5005
R1945 VDDA.n1152 VDDA.t574 4.5005
R1946 VDDA.n1153 VDDA.t430 4.5005
R1947 VDDA.n1154 VDDA.t827 4.5005
R1948 VDDA.n1155 VDDA.t911 4.5005
R1949 VDDA.n1156 VDDA.t766 4.5005
R1950 VDDA.n1157 VDDA.t618 4.5005
R1951 VDDA.n1158 VDDA.t702 4.5005
R1952 VDDA.n1159 VDDA.t557 4.5005
R1953 VDDA.n1160 VDDA.t957 4.5005
R1954 VDDA.n1161 VDDA.t808 4.5005
R1955 VDDA.n1162 VDDA.t894 4.5005
R1956 VDDA.n1163 VDDA.t742 4.5005
R1957 VDDA.n1164 VDDA.t817 4.5005
R1958 VDDA.n1165 VDDA.t904 4.5005
R1959 VDDA.n1166 VDDA.t754 4.5005
R1960 VDDA.n1167 VDDA.t607 4.5005
R1961 VDDA.n2404 VDDA.n2382 4.48641
R1962 VDDA.n2405 VDDA.n2404 4.48641
R1963 VDDA.n2411 VDDA.n2363 4.48641
R1964 VDDA.n2412 VDDA.n2411 4.48641
R1965 VDDA.n2000 VDDA.n1993 3.75335
R1966 VDDA.n1995 VDDA.n1949 3.75335
R1967 VDDA.n1987 VDDA.n1986 3.75335
R1968 VDDA.n1982 VDDA.n1959 3.75335
R1969 VDDA.n2025 VDDA.n2024 3.75335
R1970 VDDA.n2023 VDDA.n2008 3.75335
R1971 VDDA.n2019 VDDA.n2018 3.75335
R1972 VDDA.n2017 VDDA.n2016 3.75335
R1973 VDDA.n3356 VDDA.n3355 3.62427
R1974 VDDA.n3190 VDDA.n3189 3.62427
R1975 VDDA.n3023 VDDA.n180 3.62427
R1976 VDDA.n2857 VDDA.n2856 3.62427
R1977 VDDA.n2682 VDDA.n2681 3.62427
R1978 VDDA.n1664 VDDA.n517 3.62427
R1979 VDDA.n1498 VDDA.n1497 3.62427
R1980 VDDA.n1496 VDDA.n1495 3.62427
R1981 VDDA.n2805 VDDA.n2789 3.563
R1982 VDDA.n2839 VDDA.n2805 3.563
R1983 VDDA.n2335 VDDA.n2334 3.47871
R1984 VDDA.n2150 VDDA.n2149 3.47871
R1985 VDDA.n353 VDDA.n352 3.47871
R1986 VDDA.n2676 VDDA.n2675 3.47871
R1987 VDDA.n2531 VDDA.n2530 3.47871
R1988 VDDA.n90 VDDA.n18 3.47821
R1989 VDDA.n3238 VDDA.n3237 3.47821
R1990 VDDA.n3093 VDDA.n3027 3.47821
R1991 VDDA.n2933 VDDA.n2861 3.47821
R1992 VDDA.n427 VDDA.n355 3.47821
R1993 VDDA.n1734 VDDA.n1668 3.47821
R1994 VDDA.n1574 VDDA.n1502 3.47821
R1995 VDDA.n594 VDDA.n522 3.47821
R1996 VDDA.n1378 VDDA.n1377 3.47821
R1997 VDDA.n1214 VDDA.n1168 3.47821
R1998 VDDA.n2153 VDDA.n2152 3.4105
R1999 VDDA.n2332 VDDA.n2331 3.4105
R2000 VDDA.n2330 VDDA.n2329 3.4105
R2001 VDDA.n2328 VDDA.n2327 3.4105
R2002 VDDA.n2326 VDDA.n2155 3.4105
R2003 VDDA.n2322 VDDA.n2321 3.4105
R2004 VDDA.n2320 VDDA.n2319 3.4105
R2005 VDDA.n2318 VDDA.n2317 3.4105
R2006 VDDA.n2316 VDDA.n2157 3.4105
R2007 VDDA.n2312 VDDA.n2311 3.4105
R2008 VDDA.n2310 VDDA.n2309 3.4105
R2009 VDDA.n2308 VDDA.n2307 3.4105
R2010 VDDA.n2306 VDDA.n2159 3.4105
R2011 VDDA.n2302 VDDA.n2301 3.4105
R2012 VDDA.n2300 VDDA.n2299 3.4105
R2013 VDDA.n2298 VDDA.n2297 3.4105
R2014 VDDA.n2296 VDDA.n2161 3.4105
R2015 VDDA.n2292 VDDA.n2291 3.4105
R2016 VDDA.n2290 VDDA.n2289 3.4105
R2017 VDDA.n2288 VDDA.n2287 3.4105
R2018 VDDA.n2286 VDDA.n2163 3.4105
R2019 VDDA.n2282 VDDA.n2281 3.4105
R2020 VDDA.n2280 VDDA.n2279 3.4105
R2021 VDDA.n2278 VDDA.n2277 3.4105
R2022 VDDA.n2276 VDDA.n2165 3.4105
R2023 VDDA.n2272 VDDA.n2271 3.4105
R2024 VDDA.n2270 VDDA.n2269 3.4105
R2025 VDDA.n2268 VDDA.n2267 3.4105
R2026 VDDA.n2266 VDDA.n2167 3.4105
R2027 VDDA.n2262 VDDA.n2261 3.4105
R2028 VDDA.n2260 VDDA.n2259 3.4105
R2029 VDDA.n2258 VDDA.n2257 3.4105
R2030 VDDA.n2256 VDDA.n2169 3.4105
R2031 VDDA.n2252 VDDA.n2251 3.4105
R2032 VDDA.n2250 VDDA.n2249 3.4105
R2033 VDDA.n2248 VDDA.n2247 3.4105
R2034 VDDA.n2246 VDDA.n2171 3.4105
R2035 VDDA.n2242 VDDA.n2241 3.4105
R2036 VDDA.n2240 VDDA.n2239 3.4105
R2037 VDDA.n2238 VDDA.n2237 3.4105
R2038 VDDA.n2236 VDDA.n2173 3.4105
R2039 VDDA.n2232 VDDA.n2231 3.4105
R2040 VDDA.n2230 VDDA.n2229 3.4105
R2041 VDDA.n2228 VDDA.n2227 3.4105
R2042 VDDA.n2226 VDDA.n2175 3.4105
R2043 VDDA.n2222 VDDA.n2221 3.4105
R2044 VDDA.n2220 VDDA.n1875 3.4105
R2045 VDDA.n1924 VDDA.n1923 3.4105
R2046 VDDA.n2147 VDDA.n2146 3.4105
R2047 VDDA.n2145 VDDA.n2144 3.4105
R2048 VDDA.n2143 VDDA.n2142 3.4105
R2049 VDDA.n2141 VDDA.n1926 3.4105
R2050 VDDA.n2137 VDDA.n2136 3.4105
R2051 VDDA.n2135 VDDA.n2134 3.4105
R2052 VDDA.n2133 VDDA.n2132 3.4105
R2053 VDDA.n2131 VDDA.n1928 3.4105
R2054 VDDA.n2127 VDDA.n2126 3.4105
R2055 VDDA.n2125 VDDA.n2124 3.4105
R2056 VDDA.n2123 VDDA.n2122 3.4105
R2057 VDDA.n2121 VDDA.n1930 3.4105
R2058 VDDA.n2117 VDDA.n2116 3.4105
R2059 VDDA.n2115 VDDA.n2114 3.4105
R2060 VDDA.n2113 VDDA.n2112 3.4105
R2061 VDDA.n2111 VDDA.n1932 3.4105
R2062 VDDA.n2107 VDDA.n2106 3.4105
R2063 VDDA.n2105 VDDA.n2104 3.4105
R2064 VDDA.n2103 VDDA.n2102 3.4105
R2065 VDDA.n2101 VDDA.n1934 3.4105
R2066 VDDA.n2097 VDDA.n2096 3.4105
R2067 VDDA.n2095 VDDA.n2094 3.4105
R2068 VDDA.n2093 VDDA.n2092 3.4105
R2069 VDDA.n2091 VDDA.n1936 3.4105
R2070 VDDA.n2087 VDDA.n2086 3.4105
R2071 VDDA.n2085 VDDA.n2084 3.4105
R2072 VDDA.n2083 VDDA.n2082 3.4105
R2073 VDDA.n2081 VDDA.n1938 3.4105
R2074 VDDA.n2077 VDDA.n2076 3.4105
R2075 VDDA.n2075 VDDA.n2074 3.4105
R2076 VDDA.n2073 VDDA.n2072 3.4105
R2077 VDDA.n2071 VDDA.n1940 3.4105
R2078 VDDA.n2067 VDDA.n2066 3.4105
R2079 VDDA.n2065 VDDA.n2064 3.4105
R2080 VDDA.n2063 VDDA.n2062 3.4105
R2081 VDDA.n2061 VDDA.n1942 3.4105
R2082 VDDA.n2057 VDDA.n2056 3.4105
R2083 VDDA.n2055 VDDA.n2054 3.4105
R2084 VDDA.n2053 VDDA.n2052 3.4105
R2085 VDDA.n2051 VDDA.n1944 3.4105
R2086 VDDA.n2047 VDDA.n2046 3.4105
R2087 VDDA.n2045 VDDA.n2044 3.4105
R2088 VDDA.n2043 VDDA.n2042 3.4105
R2089 VDDA.n2041 VDDA.n1946 3.4105
R2090 VDDA.n2037 VDDA.n2036 3.4105
R2091 VDDA.n2035 VDDA.n1899 3.4105
R2092 VDDA.n209 VDDA.n208 3.4105
R2093 VDDA.n350 VDDA.n349 3.4105
R2094 VDDA.n348 VDDA.n347 3.4105
R2095 VDDA.n346 VDDA.n345 3.4105
R2096 VDDA.n344 VDDA.n211 3.4105
R2097 VDDA.n340 VDDA.n339 3.4105
R2098 VDDA.n338 VDDA.n337 3.4105
R2099 VDDA.n336 VDDA.n335 3.4105
R2100 VDDA.n334 VDDA.n213 3.4105
R2101 VDDA.n330 VDDA.n329 3.4105
R2102 VDDA.n328 VDDA.n327 3.4105
R2103 VDDA.n326 VDDA.n325 3.4105
R2104 VDDA.n324 VDDA.n215 3.4105
R2105 VDDA.n320 VDDA.n319 3.4105
R2106 VDDA.n318 VDDA.n317 3.4105
R2107 VDDA.n316 VDDA.n315 3.4105
R2108 VDDA.n314 VDDA.n217 3.4105
R2109 VDDA.n310 VDDA.n309 3.4105
R2110 VDDA.n308 VDDA.n307 3.4105
R2111 VDDA.n306 VDDA.n305 3.4105
R2112 VDDA.n304 VDDA.n219 3.4105
R2113 VDDA.n300 VDDA.n299 3.4105
R2114 VDDA.n298 VDDA.n297 3.4105
R2115 VDDA.n296 VDDA.n295 3.4105
R2116 VDDA.n294 VDDA.n221 3.4105
R2117 VDDA.n290 VDDA.n289 3.4105
R2118 VDDA.n288 VDDA.n287 3.4105
R2119 VDDA.n286 VDDA.n285 3.4105
R2120 VDDA.n284 VDDA.n223 3.4105
R2121 VDDA.n280 VDDA.n279 3.4105
R2122 VDDA.n278 VDDA.n277 3.4105
R2123 VDDA.n276 VDDA.n275 3.4105
R2124 VDDA.n274 VDDA.n225 3.4105
R2125 VDDA.n270 VDDA.n269 3.4105
R2126 VDDA.n268 VDDA.n267 3.4105
R2127 VDDA.n266 VDDA.n265 3.4105
R2128 VDDA.n264 VDDA.n227 3.4105
R2129 VDDA.n260 VDDA.n259 3.4105
R2130 VDDA.n258 VDDA.n257 3.4105
R2131 VDDA.n256 VDDA.n255 3.4105
R2132 VDDA.n254 VDDA.n229 3.4105
R2133 VDDA.n250 VDDA.n249 3.4105
R2134 VDDA.n248 VDDA.n247 3.4105
R2135 VDDA.n246 VDDA.n245 3.4105
R2136 VDDA.n244 VDDA.n231 3.4105
R2137 VDDA.n240 VDDA.n239 3.4105
R2138 VDDA.n238 VDDA.n184 3.4105
R2139 VDDA.n2534 VDDA.n2533 3.4105
R2140 VDDA.n2673 VDDA.n2672 3.4105
R2141 VDDA.n2671 VDDA.n2670 3.4105
R2142 VDDA.n2669 VDDA.n2668 3.4105
R2143 VDDA.n2667 VDDA.n2536 3.4105
R2144 VDDA.n2663 VDDA.n2662 3.4105
R2145 VDDA.n2661 VDDA.n2660 3.4105
R2146 VDDA.n2659 VDDA.n2658 3.4105
R2147 VDDA.n2657 VDDA.n2538 3.4105
R2148 VDDA.n2653 VDDA.n2652 3.4105
R2149 VDDA.n2651 VDDA.n2650 3.4105
R2150 VDDA.n2649 VDDA.n2648 3.4105
R2151 VDDA.n2647 VDDA.n2540 3.4105
R2152 VDDA.n2643 VDDA.n2642 3.4105
R2153 VDDA.n2641 VDDA.n2640 3.4105
R2154 VDDA.n2639 VDDA.n2638 3.4105
R2155 VDDA.n2637 VDDA.n2542 3.4105
R2156 VDDA.n2633 VDDA.n2632 3.4105
R2157 VDDA.n2631 VDDA.n2630 3.4105
R2158 VDDA.n2629 VDDA.n2628 3.4105
R2159 VDDA.n2627 VDDA.n2544 3.4105
R2160 VDDA.n2623 VDDA.n2622 3.4105
R2161 VDDA.n2621 VDDA.n2620 3.4105
R2162 VDDA.n2619 VDDA.n2618 3.4105
R2163 VDDA.n2617 VDDA.n2546 3.4105
R2164 VDDA.n2613 VDDA.n2612 3.4105
R2165 VDDA.n2611 VDDA.n2610 3.4105
R2166 VDDA.n2609 VDDA.n2608 3.4105
R2167 VDDA.n2607 VDDA.n2548 3.4105
R2168 VDDA.n2603 VDDA.n2602 3.4105
R2169 VDDA.n2601 VDDA.n2600 3.4105
R2170 VDDA.n2599 VDDA.n2598 3.4105
R2171 VDDA.n2597 VDDA.n2550 3.4105
R2172 VDDA.n2593 VDDA.n2592 3.4105
R2173 VDDA.n2591 VDDA.n2590 3.4105
R2174 VDDA.n2589 VDDA.n2588 3.4105
R2175 VDDA.n2587 VDDA.n2552 3.4105
R2176 VDDA.n2583 VDDA.n2582 3.4105
R2177 VDDA.n2581 VDDA.n2580 3.4105
R2178 VDDA.n2579 VDDA.n2578 3.4105
R2179 VDDA.n2577 VDDA.n2554 3.4105
R2180 VDDA.n2573 VDDA.n2572 3.4105
R2181 VDDA.n2571 VDDA.n2570 3.4105
R2182 VDDA.n2569 VDDA.n2568 3.4105
R2183 VDDA.n2567 VDDA.n2556 3.4105
R2184 VDDA.n2563 VDDA.n2562 3.4105
R2185 VDDA.n2561 VDDA.n1827 3.4105
R2186 VDDA.n2338 VDDA.n2337 3.4105
R2187 VDDA.n2528 VDDA.n2527 3.4105
R2188 VDDA.n2526 VDDA.n2525 3.4105
R2189 VDDA.n2524 VDDA.n2523 3.4105
R2190 VDDA.n2522 VDDA.n2340 3.4105
R2191 VDDA.n2518 VDDA.n2517 3.4105
R2192 VDDA.n2516 VDDA.n2515 3.4105
R2193 VDDA.n2514 VDDA.n2513 3.4105
R2194 VDDA.n2512 VDDA.n2342 3.4105
R2195 VDDA.n2508 VDDA.n2507 3.4105
R2196 VDDA.n2506 VDDA.n2505 3.4105
R2197 VDDA.n2504 VDDA.n2503 3.4105
R2198 VDDA.n2502 VDDA.n2344 3.4105
R2199 VDDA.n2498 VDDA.n2497 3.4105
R2200 VDDA.n2496 VDDA.n2495 3.4105
R2201 VDDA.n2494 VDDA.n2493 3.4105
R2202 VDDA.n2492 VDDA.n2346 3.4105
R2203 VDDA.n2488 VDDA.n2487 3.4105
R2204 VDDA.n2486 VDDA.n2485 3.4105
R2205 VDDA.n2484 VDDA.n2483 3.4105
R2206 VDDA.n2482 VDDA.n2348 3.4105
R2207 VDDA.n2478 VDDA.n2477 3.4105
R2208 VDDA.n2476 VDDA.n2475 3.4105
R2209 VDDA.n2474 VDDA.n2473 3.4105
R2210 VDDA.n2472 VDDA.n2350 3.4105
R2211 VDDA.n2468 VDDA.n2467 3.4105
R2212 VDDA.n2466 VDDA.n2465 3.4105
R2213 VDDA.n2464 VDDA.n2463 3.4105
R2214 VDDA.n2462 VDDA.n2352 3.4105
R2215 VDDA.n2458 VDDA.n2457 3.4105
R2216 VDDA.n2456 VDDA.n2455 3.4105
R2217 VDDA.n2454 VDDA.n2453 3.4105
R2218 VDDA.n2452 VDDA.n2354 3.4105
R2219 VDDA.n2448 VDDA.n2447 3.4105
R2220 VDDA.n2446 VDDA.n2445 3.4105
R2221 VDDA.n2444 VDDA.n2443 3.4105
R2222 VDDA.n2442 VDDA.n2356 3.4105
R2223 VDDA.n2438 VDDA.n2437 3.4105
R2224 VDDA.n2436 VDDA.n2435 3.4105
R2225 VDDA.n2434 VDDA.n2433 3.4105
R2226 VDDA.n2432 VDDA.n2358 3.4105
R2227 VDDA.n2428 VDDA.n2427 3.4105
R2228 VDDA.n2426 VDDA.n2425 3.4105
R2229 VDDA.n2424 VDDA.n2423 3.4105
R2230 VDDA.n2422 VDDA.n2360 3.4105
R2231 VDDA.n2418 VDDA.n2417 3.4105
R2232 VDDA.n2416 VDDA.n1851 3.4105
R2233 VDDA.n43 VDDA.n42 3.4105
R2234 VDDA.n177 VDDA.n176 3.4105
R2235 VDDA.n175 VDDA.n174 3.4105
R2236 VDDA.n173 VDDA.n47 3.4105
R2237 VDDA.n46 VDDA.n45 3.4105
R2238 VDDA.n169 VDDA.n168 3.4105
R2239 VDDA.n167 VDDA.n166 3.4105
R2240 VDDA.n165 VDDA.n51 3.4105
R2241 VDDA.n50 VDDA.n49 3.4105
R2242 VDDA.n161 VDDA.n160 3.4105
R2243 VDDA.n159 VDDA.n158 3.4105
R2244 VDDA.n157 VDDA.n55 3.4105
R2245 VDDA.n54 VDDA.n53 3.4105
R2246 VDDA.n153 VDDA.n152 3.4105
R2247 VDDA.n151 VDDA.n150 3.4105
R2248 VDDA.n149 VDDA.n59 3.4105
R2249 VDDA.n58 VDDA.n57 3.4105
R2250 VDDA.n145 VDDA.n144 3.4105
R2251 VDDA.n143 VDDA.n142 3.4105
R2252 VDDA.n141 VDDA.n63 3.4105
R2253 VDDA.n62 VDDA.n61 3.4105
R2254 VDDA.n137 VDDA.n136 3.4105
R2255 VDDA.n135 VDDA.n134 3.4105
R2256 VDDA.n133 VDDA.n67 3.4105
R2257 VDDA.n66 VDDA.n65 3.4105
R2258 VDDA.n129 VDDA.n128 3.4105
R2259 VDDA.n127 VDDA.n126 3.4105
R2260 VDDA.n125 VDDA.n71 3.4105
R2261 VDDA.n70 VDDA.n69 3.4105
R2262 VDDA.n121 VDDA.n120 3.4105
R2263 VDDA.n119 VDDA.n118 3.4105
R2264 VDDA.n117 VDDA.n75 3.4105
R2265 VDDA.n74 VDDA.n73 3.4105
R2266 VDDA.n113 VDDA.n112 3.4105
R2267 VDDA.n111 VDDA.n110 3.4105
R2268 VDDA.n109 VDDA.n79 3.4105
R2269 VDDA.n78 VDDA.n77 3.4105
R2270 VDDA.n105 VDDA.n104 3.4105
R2271 VDDA.n103 VDDA.n102 3.4105
R2272 VDDA.n101 VDDA.n83 3.4105
R2273 VDDA.n82 VDDA.n81 3.4105
R2274 VDDA.n97 VDDA.n96 3.4105
R2275 VDDA.n95 VDDA.n94 3.4105
R2276 VDDA.n93 VDDA.n87 3.4105
R2277 VDDA.n86 VDDA.n85 3.4105
R2278 VDDA.n89 VDDA.n88 3.4105
R2279 VDDA.n3359 VDDA.n3358 3.4105
R2280 VDDA.n3352 VDDA.n3192 3.4105
R2281 VDDA.n3350 VDDA.n3349 3.4105
R2282 VDDA.n3194 VDDA.n3193 3.4105
R2283 VDDA.n3345 VDDA.n3344 3.4105
R2284 VDDA.n3342 VDDA.n3196 3.4105
R2285 VDDA.n3340 VDDA.n3339 3.4105
R2286 VDDA.n3198 VDDA.n3197 3.4105
R2287 VDDA.n3335 VDDA.n3334 3.4105
R2288 VDDA.n3332 VDDA.n3200 3.4105
R2289 VDDA.n3330 VDDA.n3329 3.4105
R2290 VDDA.n3202 VDDA.n3201 3.4105
R2291 VDDA.n3325 VDDA.n3324 3.4105
R2292 VDDA.n3322 VDDA.n3204 3.4105
R2293 VDDA.n3320 VDDA.n3319 3.4105
R2294 VDDA.n3206 VDDA.n3205 3.4105
R2295 VDDA.n3315 VDDA.n3314 3.4105
R2296 VDDA.n3312 VDDA.n3208 3.4105
R2297 VDDA.n3310 VDDA.n3309 3.4105
R2298 VDDA.n3210 VDDA.n3209 3.4105
R2299 VDDA.n3305 VDDA.n3304 3.4105
R2300 VDDA.n3302 VDDA.n3212 3.4105
R2301 VDDA.n3300 VDDA.n3299 3.4105
R2302 VDDA.n3214 VDDA.n3213 3.4105
R2303 VDDA.n3295 VDDA.n3294 3.4105
R2304 VDDA.n3292 VDDA.n3216 3.4105
R2305 VDDA.n3290 VDDA.n3289 3.4105
R2306 VDDA.n3218 VDDA.n3217 3.4105
R2307 VDDA.n3285 VDDA.n3284 3.4105
R2308 VDDA.n3282 VDDA.n3220 3.4105
R2309 VDDA.n3280 VDDA.n3279 3.4105
R2310 VDDA.n3222 VDDA.n3221 3.4105
R2311 VDDA.n3275 VDDA.n3274 3.4105
R2312 VDDA.n3272 VDDA.n3224 3.4105
R2313 VDDA.n3270 VDDA.n3269 3.4105
R2314 VDDA.n3226 VDDA.n3225 3.4105
R2315 VDDA.n3265 VDDA.n3264 3.4105
R2316 VDDA.n3262 VDDA.n3228 3.4105
R2317 VDDA.n3260 VDDA.n3259 3.4105
R2318 VDDA.n3230 VDDA.n3229 3.4105
R2319 VDDA.n3255 VDDA.n3254 3.4105
R2320 VDDA.n3252 VDDA.n3232 3.4105
R2321 VDDA.n3250 VDDA.n3249 3.4105
R2322 VDDA.n3234 VDDA.n3233 3.4105
R2323 VDDA.n3245 VDDA.n3244 3.4105
R2324 VDDA.n3242 VDDA.n3236 3.4105
R2325 VDDA.n3240 VDDA.n3239 3.4105
R2326 VDDA.n3354 VDDA.n3353 3.4105
R2327 VDDA.n183 VDDA.n182 3.4105
R2328 VDDA.n3184 VDDA.n3183 3.4105
R2329 VDDA.n3051 VDDA.n3050 3.4105
R2330 VDDA.n3179 VDDA.n3178 3.4105
R2331 VDDA.n3177 VDDA.n3176 3.4105
R2332 VDDA.n3175 VDDA.n3055 3.4105
R2333 VDDA.n3054 VDDA.n3053 3.4105
R2334 VDDA.n3171 VDDA.n3170 3.4105
R2335 VDDA.n3169 VDDA.n3168 3.4105
R2336 VDDA.n3167 VDDA.n3059 3.4105
R2337 VDDA.n3058 VDDA.n3057 3.4105
R2338 VDDA.n3163 VDDA.n3162 3.4105
R2339 VDDA.n3161 VDDA.n3160 3.4105
R2340 VDDA.n3159 VDDA.n3063 3.4105
R2341 VDDA.n3062 VDDA.n3061 3.4105
R2342 VDDA.n3155 VDDA.n3154 3.4105
R2343 VDDA.n3153 VDDA.n3152 3.4105
R2344 VDDA.n3151 VDDA.n3067 3.4105
R2345 VDDA.n3066 VDDA.n3065 3.4105
R2346 VDDA.n3147 VDDA.n3146 3.4105
R2347 VDDA.n3145 VDDA.n3144 3.4105
R2348 VDDA.n3143 VDDA.n3071 3.4105
R2349 VDDA.n3070 VDDA.n3069 3.4105
R2350 VDDA.n3139 VDDA.n3138 3.4105
R2351 VDDA.n3137 VDDA.n3136 3.4105
R2352 VDDA.n3135 VDDA.n3075 3.4105
R2353 VDDA.n3074 VDDA.n3073 3.4105
R2354 VDDA.n3131 VDDA.n3130 3.4105
R2355 VDDA.n3129 VDDA.n3128 3.4105
R2356 VDDA.n3127 VDDA.n3079 3.4105
R2357 VDDA.n3078 VDDA.n3077 3.4105
R2358 VDDA.n3123 VDDA.n3122 3.4105
R2359 VDDA.n3121 VDDA.n3120 3.4105
R2360 VDDA.n3119 VDDA.n3083 3.4105
R2361 VDDA.n3082 VDDA.n3081 3.4105
R2362 VDDA.n3115 VDDA.n3114 3.4105
R2363 VDDA.n3113 VDDA.n3112 3.4105
R2364 VDDA.n3111 VDDA.n3087 3.4105
R2365 VDDA.n3086 VDDA.n3085 3.4105
R2366 VDDA.n3107 VDDA.n3106 3.4105
R2367 VDDA.n3105 VDDA.n3104 3.4105
R2368 VDDA.n3103 VDDA.n3091 3.4105
R2369 VDDA.n3090 VDDA.n3089 3.4105
R2370 VDDA.n3099 VDDA.n3098 3.4105
R2371 VDDA.n3097 VDDA.n3096 3.4105
R2372 VDDA.n3095 VDDA.n3094 3.4105
R2373 VDDA.n3188 VDDA.n3187 3.4105
R2374 VDDA.n2886 VDDA.n2885 3.4105
R2375 VDDA.n3020 VDDA.n3019 3.4105
R2376 VDDA.n3018 VDDA.n3017 3.4105
R2377 VDDA.n3016 VDDA.n2890 3.4105
R2378 VDDA.n2889 VDDA.n2888 3.4105
R2379 VDDA.n3012 VDDA.n3011 3.4105
R2380 VDDA.n3010 VDDA.n3009 3.4105
R2381 VDDA.n3008 VDDA.n2894 3.4105
R2382 VDDA.n2893 VDDA.n2892 3.4105
R2383 VDDA.n3004 VDDA.n3003 3.4105
R2384 VDDA.n3002 VDDA.n3001 3.4105
R2385 VDDA.n3000 VDDA.n2898 3.4105
R2386 VDDA.n2897 VDDA.n2896 3.4105
R2387 VDDA.n2996 VDDA.n2995 3.4105
R2388 VDDA.n2994 VDDA.n2993 3.4105
R2389 VDDA.n2992 VDDA.n2902 3.4105
R2390 VDDA.n2901 VDDA.n2900 3.4105
R2391 VDDA.n2988 VDDA.n2987 3.4105
R2392 VDDA.n2986 VDDA.n2985 3.4105
R2393 VDDA.n2984 VDDA.n2906 3.4105
R2394 VDDA.n2905 VDDA.n2904 3.4105
R2395 VDDA.n2980 VDDA.n2979 3.4105
R2396 VDDA.n2978 VDDA.n2977 3.4105
R2397 VDDA.n2976 VDDA.n2910 3.4105
R2398 VDDA.n2909 VDDA.n2908 3.4105
R2399 VDDA.n2972 VDDA.n2971 3.4105
R2400 VDDA.n2970 VDDA.n2969 3.4105
R2401 VDDA.n2968 VDDA.n2914 3.4105
R2402 VDDA.n2913 VDDA.n2912 3.4105
R2403 VDDA.n2964 VDDA.n2963 3.4105
R2404 VDDA.n2962 VDDA.n2961 3.4105
R2405 VDDA.n2960 VDDA.n2918 3.4105
R2406 VDDA.n2917 VDDA.n2916 3.4105
R2407 VDDA.n2956 VDDA.n2955 3.4105
R2408 VDDA.n2954 VDDA.n2953 3.4105
R2409 VDDA.n2952 VDDA.n2922 3.4105
R2410 VDDA.n2921 VDDA.n2920 3.4105
R2411 VDDA.n2948 VDDA.n2947 3.4105
R2412 VDDA.n2946 VDDA.n2945 3.4105
R2413 VDDA.n2944 VDDA.n2926 3.4105
R2414 VDDA.n2925 VDDA.n2924 3.4105
R2415 VDDA.n2940 VDDA.n2939 3.4105
R2416 VDDA.n2938 VDDA.n2937 3.4105
R2417 VDDA.n2936 VDDA.n2930 3.4105
R2418 VDDA.n2929 VDDA.n2928 3.4105
R2419 VDDA.n2932 VDDA.n2931 3.4105
R2420 VDDA.n3025 VDDA.n3024 3.4105
R2421 VDDA.n380 VDDA.n379 3.4105
R2422 VDDA.n514 VDDA.n513 3.4105
R2423 VDDA.n512 VDDA.n511 3.4105
R2424 VDDA.n510 VDDA.n384 3.4105
R2425 VDDA.n383 VDDA.n382 3.4105
R2426 VDDA.n506 VDDA.n505 3.4105
R2427 VDDA.n504 VDDA.n503 3.4105
R2428 VDDA.n502 VDDA.n388 3.4105
R2429 VDDA.n387 VDDA.n386 3.4105
R2430 VDDA.n498 VDDA.n497 3.4105
R2431 VDDA.n496 VDDA.n495 3.4105
R2432 VDDA.n494 VDDA.n392 3.4105
R2433 VDDA.n391 VDDA.n390 3.4105
R2434 VDDA.n490 VDDA.n489 3.4105
R2435 VDDA.n488 VDDA.n487 3.4105
R2436 VDDA.n486 VDDA.n396 3.4105
R2437 VDDA.n395 VDDA.n394 3.4105
R2438 VDDA.n482 VDDA.n481 3.4105
R2439 VDDA.n480 VDDA.n479 3.4105
R2440 VDDA.n478 VDDA.n400 3.4105
R2441 VDDA.n399 VDDA.n398 3.4105
R2442 VDDA.n474 VDDA.n473 3.4105
R2443 VDDA.n472 VDDA.n471 3.4105
R2444 VDDA.n470 VDDA.n404 3.4105
R2445 VDDA.n403 VDDA.n402 3.4105
R2446 VDDA.n466 VDDA.n465 3.4105
R2447 VDDA.n464 VDDA.n463 3.4105
R2448 VDDA.n462 VDDA.n408 3.4105
R2449 VDDA.n407 VDDA.n406 3.4105
R2450 VDDA.n458 VDDA.n457 3.4105
R2451 VDDA.n456 VDDA.n455 3.4105
R2452 VDDA.n454 VDDA.n412 3.4105
R2453 VDDA.n411 VDDA.n410 3.4105
R2454 VDDA.n450 VDDA.n449 3.4105
R2455 VDDA.n448 VDDA.n447 3.4105
R2456 VDDA.n446 VDDA.n416 3.4105
R2457 VDDA.n415 VDDA.n414 3.4105
R2458 VDDA.n442 VDDA.n441 3.4105
R2459 VDDA.n440 VDDA.n439 3.4105
R2460 VDDA.n438 VDDA.n420 3.4105
R2461 VDDA.n419 VDDA.n418 3.4105
R2462 VDDA.n434 VDDA.n433 3.4105
R2463 VDDA.n432 VDDA.n431 3.4105
R2464 VDDA.n430 VDDA.n424 3.4105
R2465 VDDA.n423 VDDA.n422 3.4105
R2466 VDDA.n426 VDDA.n425 3.4105
R2467 VDDA.n2859 VDDA.n2858 3.4105
R2468 VDDA.n520 VDDA.n519 3.4105
R2469 VDDA.n1825 VDDA.n1824 3.4105
R2470 VDDA.n1692 VDDA.n1691 3.4105
R2471 VDDA.n1820 VDDA.n1819 3.4105
R2472 VDDA.n1818 VDDA.n1817 3.4105
R2473 VDDA.n1816 VDDA.n1696 3.4105
R2474 VDDA.n1695 VDDA.n1694 3.4105
R2475 VDDA.n1812 VDDA.n1811 3.4105
R2476 VDDA.n1810 VDDA.n1809 3.4105
R2477 VDDA.n1808 VDDA.n1700 3.4105
R2478 VDDA.n1699 VDDA.n1698 3.4105
R2479 VDDA.n1804 VDDA.n1803 3.4105
R2480 VDDA.n1802 VDDA.n1801 3.4105
R2481 VDDA.n1800 VDDA.n1704 3.4105
R2482 VDDA.n1703 VDDA.n1702 3.4105
R2483 VDDA.n1796 VDDA.n1795 3.4105
R2484 VDDA.n1794 VDDA.n1793 3.4105
R2485 VDDA.n1792 VDDA.n1708 3.4105
R2486 VDDA.n1707 VDDA.n1706 3.4105
R2487 VDDA.n1788 VDDA.n1787 3.4105
R2488 VDDA.n1786 VDDA.n1785 3.4105
R2489 VDDA.n1784 VDDA.n1712 3.4105
R2490 VDDA.n1711 VDDA.n1710 3.4105
R2491 VDDA.n1780 VDDA.n1779 3.4105
R2492 VDDA.n1778 VDDA.n1777 3.4105
R2493 VDDA.n1776 VDDA.n1716 3.4105
R2494 VDDA.n1715 VDDA.n1714 3.4105
R2495 VDDA.n1772 VDDA.n1771 3.4105
R2496 VDDA.n1770 VDDA.n1769 3.4105
R2497 VDDA.n1768 VDDA.n1720 3.4105
R2498 VDDA.n1719 VDDA.n1718 3.4105
R2499 VDDA.n1764 VDDA.n1763 3.4105
R2500 VDDA.n1762 VDDA.n1761 3.4105
R2501 VDDA.n1760 VDDA.n1724 3.4105
R2502 VDDA.n1723 VDDA.n1722 3.4105
R2503 VDDA.n1756 VDDA.n1755 3.4105
R2504 VDDA.n1754 VDDA.n1753 3.4105
R2505 VDDA.n1752 VDDA.n1728 3.4105
R2506 VDDA.n1727 VDDA.n1726 3.4105
R2507 VDDA.n1748 VDDA.n1747 3.4105
R2508 VDDA.n1746 VDDA.n1745 3.4105
R2509 VDDA.n1744 VDDA.n1732 3.4105
R2510 VDDA.n1731 VDDA.n1730 3.4105
R2511 VDDA.n1740 VDDA.n1739 3.4105
R2512 VDDA.n1738 VDDA.n1737 3.4105
R2513 VDDA.n1736 VDDA.n1735 3.4105
R2514 VDDA.n2680 VDDA.n2679 3.4105
R2515 VDDA.n1527 VDDA.n1526 3.4105
R2516 VDDA.n1661 VDDA.n1660 3.4105
R2517 VDDA.n1659 VDDA.n1658 3.4105
R2518 VDDA.n1657 VDDA.n1531 3.4105
R2519 VDDA.n1530 VDDA.n1529 3.4105
R2520 VDDA.n1653 VDDA.n1652 3.4105
R2521 VDDA.n1651 VDDA.n1650 3.4105
R2522 VDDA.n1649 VDDA.n1535 3.4105
R2523 VDDA.n1534 VDDA.n1533 3.4105
R2524 VDDA.n1645 VDDA.n1644 3.4105
R2525 VDDA.n1643 VDDA.n1642 3.4105
R2526 VDDA.n1641 VDDA.n1539 3.4105
R2527 VDDA.n1538 VDDA.n1537 3.4105
R2528 VDDA.n1637 VDDA.n1636 3.4105
R2529 VDDA.n1635 VDDA.n1634 3.4105
R2530 VDDA.n1633 VDDA.n1543 3.4105
R2531 VDDA.n1542 VDDA.n1541 3.4105
R2532 VDDA.n1629 VDDA.n1628 3.4105
R2533 VDDA.n1627 VDDA.n1626 3.4105
R2534 VDDA.n1625 VDDA.n1547 3.4105
R2535 VDDA.n1546 VDDA.n1545 3.4105
R2536 VDDA.n1621 VDDA.n1620 3.4105
R2537 VDDA.n1619 VDDA.n1618 3.4105
R2538 VDDA.n1617 VDDA.n1551 3.4105
R2539 VDDA.n1550 VDDA.n1549 3.4105
R2540 VDDA.n1613 VDDA.n1612 3.4105
R2541 VDDA.n1611 VDDA.n1610 3.4105
R2542 VDDA.n1609 VDDA.n1555 3.4105
R2543 VDDA.n1554 VDDA.n1553 3.4105
R2544 VDDA.n1605 VDDA.n1604 3.4105
R2545 VDDA.n1603 VDDA.n1602 3.4105
R2546 VDDA.n1601 VDDA.n1559 3.4105
R2547 VDDA.n1558 VDDA.n1557 3.4105
R2548 VDDA.n1597 VDDA.n1596 3.4105
R2549 VDDA.n1595 VDDA.n1594 3.4105
R2550 VDDA.n1593 VDDA.n1563 3.4105
R2551 VDDA.n1562 VDDA.n1561 3.4105
R2552 VDDA.n1589 VDDA.n1588 3.4105
R2553 VDDA.n1587 VDDA.n1586 3.4105
R2554 VDDA.n1585 VDDA.n1567 3.4105
R2555 VDDA.n1566 VDDA.n1565 3.4105
R2556 VDDA.n1581 VDDA.n1580 3.4105
R2557 VDDA.n1579 VDDA.n1578 3.4105
R2558 VDDA.n1577 VDDA.n1571 3.4105
R2559 VDDA.n1570 VDDA.n1569 3.4105
R2560 VDDA.n1573 VDDA.n1572 3.4105
R2561 VDDA.n1666 VDDA.n1665 3.4105
R2562 VDDA.n547 VDDA.n546 3.4105
R2563 VDDA.n681 VDDA.n680 3.4105
R2564 VDDA.n679 VDDA.n678 3.4105
R2565 VDDA.n677 VDDA.n551 3.4105
R2566 VDDA.n550 VDDA.n549 3.4105
R2567 VDDA.n673 VDDA.n672 3.4105
R2568 VDDA.n671 VDDA.n670 3.4105
R2569 VDDA.n669 VDDA.n555 3.4105
R2570 VDDA.n554 VDDA.n553 3.4105
R2571 VDDA.n665 VDDA.n664 3.4105
R2572 VDDA.n663 VDDA.n662 3.4105
R2573 VDDA.n661 VDDA.n559 3.4105
R2574 VDDA.n558 VDDA.n557 3.4105
R2575 VDDA.n657 VDDA.n656 3.4105
R2576 VDDA.n655 VDDA.n654 3.4105
R2577 VDDA.n653 VDDA.n563 3.4105
R2578 VDDA.n562 VDDA.n561 3.4105
R2579 VDDA.n649 VDDA.n648 3.4105
R2580 VDDA.n647 VDDA.n646 3.4105
R2581 VDDA.n645 VDDA.n567 3.4105
R2582 VDDA.n566 VDDA.n565 3.4105
R2583 VDDA.n641 VDDA.n640 3.4105
R2584 VDDA.n639 VDDA.n638 3.4105
R2585 VDDA.n637 VDDA.n571 3.4105
R2586 VDDA.n570 VDDA.n569 3.4105
R2587 VDDA.n633 VDDA.n632 3.4105
R2588 VDDA.n631 VDDA.n630 3.4105
R2589 VDDA.n629 VDDA.n575 3.4105
R2590 VDDA.n574 VDDA.n573 3.4105
R2591 VDDA.n625 VDDA.n624 3.4105
R2592 VDDA.n623 VDDA.n622 3.4105
R2593 VDDA.n621 VDDA.n579 3.4105
R2594 VDDA.n578 VDDA.n577 3.4105
R2595 VDDA.n617 VDDA.n616 3.4105
R2596 VDDA.n615 VDDA.n614 3.4105
R2597 VDDA.n613 VDDA.n583 3.4105
R2598 VDDA.n582 VDDA.n581 3.4105
R2599 VDDA.n609 VDDA.n608 3.4105
R2600 VDDA.n607 VDDA.n606 3.4105
R2601 VDDA.n605 VDDA.n587 3.4105
R2602 VDDA.n586 VDDA.n585 3.4105
R2603 VDDA.n601 VDDA.n600 3.4105
R2604 VDDA.n599 VDDA.n598 3.4105
R2605 VDDA.n597 VDDA.n591 3.4105
R2606 VDDA.n590 VDDA.n589 3.4105
R2607 VDDA.n593 VDDA.n592 3.4105
R2608 VDDA.n1500 VDDA.n1499 3.4105
R2609 VDDA.n1492 VDDA.n1332 3.4105
R2610 VDDA.n1490 VDDA.n1489 3.4105
R2611 VDDA.n1334 VDDA.n1333 3.4105
R2612 VDDA.n1485 VDDA.n1484 3.4105
R2613 VDDA.n1482 VDDA.n1336 3.4105
R2614 VDDA.n1480 VDDA.n1479 3.4105
R2615 VDDA.n1338 VDDA.n1337 3.4105
R2616 VDDA.n1475 VDDA.n1474 3.4105
R2617 VDDA.n1472 VDDA.n1340 3.4105
R2618 VDDA.n1470 VDDA.n1469 3.4105
R2619 VDDA.n1342 VDDA.n1341 3.4105
R2620 VDDA.n1465 VDDA.n1464 3.4105
R2621 VDDA.n1462 VDDA.n1344 3.4105
R2622 VDDA.n1460 VDDA.n1459 3.4105
R2623 VDDA.n1346 VDDA.n1345 3.4105
R2624 VDDA.n1455 VDDA.n1454 3.4105
R2625 VDDA.n1452 VDDA.n1348 3.4105
R2626 VDDA.n1450 VDDA.n1449 3.4105
R2627 VDDA.n1350 VDDA.n1349 3.4105
R2628 VDDA.n1445 VDDA.n1444 3.4105
R2629 VDDA.n1442 VDDA.n1352 3.4105
R2630 VDDA.n1440 VDDA.n1439 3.4105
R2631 VDDA.n1354 VDDA.n1353 3.4105
R2632 VDDA.n1435 VDDA.n1434 3.4105
R2633 VDDA.n1432 VDDA.n1356 3.4105
R2634 VDDA.n1430 VDDA.n1429 3.4105
R2635 VDDA.n1358 VDDA.n1357 3.4105
R2636 VDDA.n1425 VDDA.n1424 3.4105
R2637 VDDA.n1422 VDDA.n1360 3.4105
R2638 VDDA.n1420 VDDA.n1419 3.4105
R2639 VDDA.n1362 VDDA.n1361 3.4105
R2640 VDDA.n1415 VDDA.n1414 3.4105
R2641 VDDA.n1412 VDDA.n1364 3.4105
R2642 VDDA.n1410 VDDA.n1409 3.4105
R2643 VDDA.n1366 VDDA.n1365 3.4105
R2644 VDDA.n1405 VDDA.n1404 3.4105
R2645 VDDA.n1402 VDDA.n1368 3.4105
R2646 VDDA.n1400 VDDA.n1399 3.4105
R2647 VDDA.n1370 VDDA.n1369 3.4105
R2648 VDDA.n1395 VDDA.n1394 3.4105
R2649 VDDA.n1392 VDDA.n1372 3.4105
R2650 VDDA.n1390 VDDA.n1389 3.4105
R2651 VDDA.n1374 VDDA.n1373 3.4105
R2652 VDDA.n1385 VDDA.n1384 3.4105
R2653 VDDA.n1382 VDDA.n1376 3.4105
R2654 VDDA.n1380 VDDA.n1379 3.4105
R2655 VDDA.n1494 VDDA.n1493 3.4105
R2656 VDDA.n686 VDDA.n685 3.4105
R2657 VDDA.n1325 VDDA.n1324 3.4105
R2658 VDDA.n1192 VDDA.n1191 3.4105
R2659 VDDA.n1320 VDDA.n1319 3.4105
R2660 VDDA.n1318 VDDA.n1317 3.4105
R2661 VDDA.n1316 VDDA.n1315 3.4105
R2662 VDDA.n1314 VDDA.n1194 3.4105
R2663 VDDA.n1310 VDDA.n1309 3.4105
R2664 VDDA.n1308 VDDA.n1307 3.4105
R2665 VDDA.n1306 VDDA.n1305 3.4105
R2666 VDDA.n1304 VDDA.n1196 3.4105
R2667 VDDA.n1300 VDDA.n1299 3.4105
R2668 VDDA.n1298 VDDA.n1297 3.4105
R2669 VDDA.n1296 VDDA.n1295 3.4105
R2670 VDDA.n1294 VDDA.n1198 3.4105
R2671 VDDA.n1290 VDDA.n1289 3.4105
R2672 VDDA.n1288 VDDA.n1287 3.4105
R2673 VDDA.n1286 VDDA.n1285 3.4105
R2674 VDDA.n1284 VDDA.n1200 3.4105
R2675 VDDA.n1280 VDDA.n1279 3.4105
R2676 VDDA.n1278 VDDA.n1277 3.4105
R2677 VDDA.n1276 VDDA.n1275 3.4105
R2678 VDDA.n1274 VDDA.n1202 3.4105
R2679 VDDA.n1270 VDDA.n1269 3.4105
R2680 VDDA.n1268 VDDA.n1267 3.4105
R2681 VDDA.n1266 VDDA.n1265 3.4105
R2682 VDDA.n1264 VDDA.n1204 3.4105
R2683 VDDA.n1260 VDDA.n1259 3.4105
R2684 VDDA.n1258 VDDA.n1257 3.4105
R2685 VDDA.n1256 VDDA.n1255 3.4105
R2686 VDDA.n1254 VDDA.n1206 3.4105
R2687 VDDA.n1250 VDDA.n1249 3.4105
R2688 VDDA.n1248 VDDA.n1247 3.4105
R2689 VDDA.n1246 VDDA.n1245 3.4105
R2690 VDDA.n1244 VDDA.n1208 3.4105
R2691 VDDA.n1240 VDDA.n1239 3.4105
R2692 VDDA.n1238 VDDA.n1237 3.4105
R2693 VDDA.n1236 VDDA.n1235 3.4105
R2694 VDDA.n1234 VDDA.n1210 3.4105
R2695 VDDA.n1230 VDDA.n1229 3.4105
R2696 VDDA.n1228 VDDA.n1227 3.4105
R2697 VDDA.n1226 VDDA.n1225 3.4105
R2698 VDDA.n1224 VDDA.n1212 3.4105
R2699 VDDA.n1220 VDDA.n1219 3.4105
R2700 VDDA.n1218 VDDA.n1217 3.4105
R2701 VDDA.n1216 VDDA.n1215 3.4105
R2702 VDDA.n1329 VDDA.n1328 3.4105
R2703 VDDA.n1327 VDDA.n1168 3.4105
R2704 VDDA.n1328 VDDA.n1327 3.4105
R2705 VDDA.n1377 VDDA.n521 3.4105
R2706 VDDA.n1493 VDDA.n521 3.4105
R2707 VDDA.n1501 VDDA.n522 3.4105
R2708 VDDA.n1501 VDDA.n1500 3.4105
R2709 VDDA.n1667 VDDA.n1502 3.4105
R2710 VDDA.n1667 VDDA.n1666 3.4105
R2711 VDDA.n2678 VDDA.n1668 3.4105
R2712 VDDA.n2679 VDDA.n2678 3.4105
R2713 VDDA.n2860 VDDA.n355 3.4105
R2714 VDDA.n2860 VDDA.n2859 3.4105
R2715 VDDA.n3026 VDDA.n2861 3.4105
R2716 VDDA.n3026 VDDA.n3025 3.4105
R2717 VDDA.n3186 VDDA.n3027 3.4105
R2718 VDDA.n3187 VDDA.n3186 3.4105
R2719 VDDA.n3237 VDDA.n17 3.4105
R2720 VDDA.n3353 VDDA.n17 3.4105
R2721 VDDA.n3360 VDDA.n18 3.4105
R2722 VDDA.n3360 VDDA.n3359 3.4105
R2723 VDDA.n2532 VDDA.n1851 3.4105
R2724 VDDA.n2532 VDDA.n2531 3.4105
R2725 VDDA.n2677 VDDA.n1827 3.4105
R2726 VDDA.n2677 VDDA.n2676 3.4105
R2727 VDDA.n354 VDDA.n184 3.4105
R2728 VDDA.n354 VDDA.n353 3.4105
R2729 VDDA.n2151 VDDA.n1899 3.4105
R2730 VDDA.n2151 VDDA.n2150 3.4105
R2731 VDDA.n2336 VDDA.n1875 3.4105
R2732 VDDA.n2336 VDDA.n2335 3.4105
R2733 VDDA.n3467 VDDA.n15 3.4105
R2734 VDDA.n3467 VDDA.n16 3.4105
R2735 VDDA.n3467 VDDA.n3466 3.4105
R2736 VDDA.n3437 VDDA.n3378 3.4105
R2737 VDDA.n3466 VDDA.n3378 3.4105
R2738 VDDA.n3437 VDDA.n3375 3.4105
R2739 VDDA.n3436 VDDA.n3375 3.4105
R2740 VDDA.n3440 VDDA.n3375 3.4105
R2741 VDDA.n3435 VDDA.n3375 3.4105
R2742 VDDA.n3442 VDDA.n3375 3.4105
R2743 VDDA.n3434 VDDA.n3375 3.4105
R2744 VDDA.n3444 VDDA.n3375 3.4105
R2745 VDDA.n3433 VDDA.n3375 3.4105
R2746 VDDA.n3446 VDDA.n3375 3.4105
R2747 VDDA.n3432 VDDA.n3375 3.4105
R2748 VDDA.n3448 VDDA.n3375 3.4105
R2749 VDDA.n3431 VDDA.n3375 3.4105
R2750 VDDA.n3450 VDDA.n3375 3.4105
R2751 VDDA.n3430 VDDA.n3375 3.4105
R2752 VDDA.n3452 VDDA.n3375 3.4105
R2753 VDDA.n3429 VDDA.n3375 3.4105
R2754 VDDA.n3454 VDDA.n3375 3.4105
R2755 VDDA.n3428 VDDA.n3375 3.4105
R2756 VDDA.n3456 VDDA.n3375 3.4105
R2757 VDDA.n3427 VDDA.n3375 3.4105
R2758 VDDA.n3458 VDDA.n3375 3.4105
R2759 VDDA.n3426 VDDA.n3375 3.4105
R2760 VDDA.n3460 VDDA.n3375 3.4105
R2761 VDDA.n3425 VDDA.n3375 3.4105
R2762 VDDA.n3462 VDDA.n3375 3.4105
R2763 VDDA.n3424 VDDA.n3375 3.4105
R2764 VDDA.n3464 VDDA.n3375 3.4105
R2765 VDDA.n3423 VDDA.n3375 3.4105
R2766 VDDA.n3375 VDDA.n16 3.4105
R2767 VDDA.n3466 VDDA.n3375 3.4105
R2768 VDDA.n3437 VDDA.n3381 3.4105
R2769 VDDA.n3436 VDDA.n3381 3.4105
R2770 VDDA.n3440 VDDA.n3381 3.4105
R2771 VDDA.n3435 VDDA.n3381 3.4105
R2772 VDDA.n3442 VDDA.n3381 3.4105
R2773 VDDA.n3434 VDDA.n3381 3.4105
R2774 VDDA.n3444 VDDA.n3381 3.4105
R2775 VDDA.n3433 VDDA.n3381 3.4105
R2776 VDDA.n3446 VDDA.n3381 3.4105
R2777 VDDA.n3432 VDDA.n3381 3.4105
R2778 VDDA.n3448 VDDA.n3381 3.4105
R2779 VDDA.n3431 VDDA.n3381 3.4105
R2780 VDDA.n3450 VDDA.n3381 3.4105
R2781 VDDA.n3430 VDDA.n3381 3.4105
R2782 VDDA.n3452 VDDA.n3381 3.4105
R2783 VDDA.n3429 VDDA.n3381 3.4105
R2784 VDDA.n3454 VDDA.n3381 3.4105
R2785 VDDA.n3428 VDDA.n3381 3.4105
R2786 VDDA.n3456 VDDA.n3381 3.4105
R2787 VDDA.n3427 VDDA.n3381 3.4105
R2788 VDDA.n3458 VDDA.n3381 3.4105
R2789 VDDA.n3426 VDDA.n3381 3.4105
R2790 VDDA.n3460 VDDA.n3381 3.4105
R2791 VDDA.n3425 VDDA.n3381 3.4105
R2792 VDDA.n3462 VDDA.n3381 3.4105
R2793 VDDA.n3424 VDDA.n3381 3.4105
R2794 VDDA.n3464 VDDA.n3381 3.4105
R2795 VDDA.n3423 VDDA.n3381 3.4105
R2796 VDDA.n3381 VDDA.n16 3.4105
R2797 VDDA.n3466 VDDA.n3381 3.4105
R2798 VDDA.n3437 VDDA.n3374 3.4105
R2799 VDDA.n3436 VDDA.n3374 3.4105
R2800 VDDA.n3440 VDDA.n3374 3.4105
R2801 VDDA.n3435 VDDA.n3374 3.4105
R2802 VDDA.n3442 VDDA.n3374 3.4105
R2803 VDDA.n3434 VDDA.n3374 3.4105
R2804 VDDA.n3444 VDDA.n3374 3.4105
R2805 VDDA.n3433 VDDA.n3374 3.4105
R2806 VDDA.n3446 VDDA.n3374 3.4105
R2807 VDDA.n3432 VDDA.n3374 3.4105
R2808 VDDA.n3448 VDDA.n3374 3.4105
R2809 VDDA.n3431 VDDA.n3374 3.4105
R2810 VDDA.n3450 VDDA.n3374 3.4105
R2811 VDDA.n3430 VDDA.n3374 3.4105
R2812 VDDA.n3452 VDDA.n3374 3.4105
R2813 VDDA.n3429 VDDA.n3374 3.4105
R2814 VDDA.n3454 VDDA.n3374 3.4105
R2815 VDDA.n3428 VDDA.n3374 3.4105
R2816 VDDA.n3456 VDDA.n3374 3.4105
R2817 VDDA.n3427 VDDA.n3374 3.4105
R2818 VDDA.n3458 VDDA.n3374 3.4105
R2819 VDDA.n3426 VDDA.n3374 3.4105
R2820 VDDA.n3460 VDDA.n3374 3.4105
R2821 VDDA.n3425 VDDA.n3374 3.4105
R2822 VDDA.n3462 VDDA.n3374 3.4105
R2823 VDDA.n3424 VDDA.n3374 3.4105
R2824 VDDA.n3464 VDDA.n3374 3.4105
R2825 VDDA.n3423 VDDA.n3374 3.4105
R2826 VDDA.n3374 VDDA.n16 3.4105
R2827 VDDA.n3466 VDDA.n3374 3.4105
R2828 VDDA.n3437 VDDA.n3384 3.4105
R2829 VDDA.n3436 VDDA.n3384 3.4105
R2830 VDDA.n3440 VDDA.n3384 3.4105
R2831 VDDA.n3435 VDDA.n3384 3.4105
R2832 VDDA.n3442 VDDA.n3384 3.4105
R2833 VDDA.n3434 VDDA.n3384 3.4105
R2834 VDDA.n3444 VDDA.n3384 3.4105
R2835 VDDA.n3433 VDDA.n3384 3.4105
R2836 VDDA.n3446 VDDA.n3384 3.4105
R2837 VDDA.n3432 VDDA.n3384 3.4105
R2838 VDDA.n3448 VDDA.n3384 3.4105
R2839 VDDA.n3431 VDDA.n3384 3.4105
R2840 VDDA.n3450 VDDA.n3384 3.4105
R2841 VDDA.n3430 VDDA.n3384 3.4105
R2842 VDDA.n3452 VDDA.n3384 3.4105
R2843 VDDA.n3429 VDDA.n3384 3.4105
R2844 VDDA.n3454 VDDA.n3384 3.4105
R2845 VDDA.n3428 VDDA.n3384 3.4105
R2846 VDDA.n3456 VDDA.n3384 3.4105
R2847 VDDA.n3427 VDDA.n3384 3.4105
R2848 VDDA.n3458 VDDA.n3384 3.4105
R2849 VDDA.n3426 VDDA.n3384 3.4105
R2850 VDDA.n3460 VDDA.n3384 3.4105
R2851 VDDA.n3425 VDDA.n3384 3.4105
R2852 VDDA.n3462 VDDA.n3384 3.4105
R2853 VDDA.n3424 VDDA.n3384 3.4105
R2854 VDDA.n3464 VDDA.n3384 3.4105
R2855 VDDA.n3423 VDDA.n3384 3.4105
R2856 VDDA.n3384 VDDA.n16 3.4105
R2857 VDDA.n3466 VDDA.n3384 3.4105
R2858 VDDA.n3437 VDDA.n3373 3.4105
R2859 VDDA.n3436 VDDA.n3373 3.4105
R2860 VDDA.n3440 VDDA.n3373 3.4105
R2861 VDDA.n3435 VDDA.n3373 3.4105
R2862 VDDA.n3442 VDDA.n3373 3.4105
R2863 VDDA.n3434 VDDA.n3373 3.4105
R2864 VDDA.n3444 VDDA.n3373 3.4105
R2865 VDDA.n3433 VDDA.n3373 3.4105
R2866 VDDA.n3446 VDDA.n3373 3.4105
R2867 VDDA.n3432 VDDA.n3373 3.4105
R2868 VDDA.n3448 VDDA.n3373 3.4105
R2869 VDDA.n3431 VDDA.n3373 3.4105
R2870 VDDA.n3450 VDDA.n3373 3.4105
R2871 VDDA.n3430 VDDA.n3373 3.4105
R2872 VDDA.n3452 VDDA.n3373 3.4105
R2873 VDDA.n3429 VDDA.n3373 3.4105
R2874 VDDA.n3454 VDDA.n3373 3.4105
R2875 VDDA.n3428 VDDA.n3373 3.4105
R2876 VDDA.n3456 VDDA.n3373 3.4105
R2877 VDDA.n3427 VDDA.n3373 3.4105
R2878 VDDA.n3458 VDDA.n3373 3.4105
R2879 VDDA.n3426 VDDA.n3373 3.4105
R2880 VDDA.n3460 VDDA.n3373 3.4105
R2881 VDDA.n3425 VDDA.n3373 3.4105
R2882 VDDA.n3462 VDDA.n3373 3.4105
R2883 VDDA.n3424 VDDA.n3373 3.4105
R2884 VDDA.n3464 VDDA.n3373 3.4105
R2885 VDDA.n3423 VDDA.n3373 3.4105
R2886 VDDA.n3373 VDDA.n16 3.4105
R2887 VDDA.n3466 VDDA.n3373 3.4105
R2888 VDDA.n3437 VDDA.n3387 3.4105
R2889 VDDA.n3436 VDDA.n3387 3.4105
R2890 VDDA.n3440 VDDA.n3387 3.4105
R2891 VDDA.n3435 VDDA.n3387 3.4105
R2892 VDDA.n3442 VDDA.n3387 3.4105
R2893 VDDA.n3434 VDDA.n3387 3.4105
R2894 VDDA.n3444 VDDA.n3387 3.4105
R2895 VDDA.n3433 VDDA.n3387 3.4105
R2896 VDDA.n3446 VDDA.n3387 3.4105
R2897 VDDA.n3432 VDDA.n3387 3.4105
R2898 VDDA.n3448 VDDA.n3387 3.4105
R2899 VDDA.n3431 VDDA.n3387 3.4105
R2900 VDDA.n3450 VDDA.n3387 3.4105
R2901 VDDA.n3430 VDDA.n3387 3.4105
R2902 VDDA.n3452 VDDA.n3387 3.4105
R2903 VDDA.n3429 VDDA.n3387 3.4105
R2904 VDDA.n3454 VDDA.n3387 3.4105
R2905 VDDA.n3428 VDDA.n3387 3.4105
R2906 VDDA.n3456 VDDA.n3387 3.4105
R2907 VDDA.n3427 VDDA.n3387 3.4105
R2908 VDDA.n3458 VDDA.n3387 3.4105
R2909 VDDA.n3426 VDDA.n3387 3.4105
R2910 VDDA.n3460 VDDA.n3387 3.4105
R2911 VDDA.n3425 VDDA.n3387 3.4105
R2912 VDDA.n3462 VDDA.n3387 3.4105
R2913 VDDA.n3424 VDDA.n3387 3.4105
R2914 VDDA.n3464 VDDA.n3387 3.4105
R2915 VDDA.n3423 VDDA.n3387 3.4105
R2916 VDDA.n3387 VDDA.n16 3.4105
R2917 VDDA.n3466 VDDA.n3387 3.4105
R2918 VDDA.n3437 VDDA.n3372 3.4105
R2919 VDDA.n3436 VDDA.n3372 3.4105
R2920 VDDA.n3440 VDDA.n3372 3.4105
R2921 VDDA.n3435 VDDA.n3372 3.4105
R2922 VDDA.n3442 VDDA.n3372 3.4105
R2923 VDDA.n3434 VDDA.n3372 3.4105
R2924 VDDA.n3444 VDDA.n3372 3.4105
R2925 VDDA.n3433 VDDA.n3372 3.4105
R2926 VDDA.n3446 VDDA.n3372 3.4105
R2927 VDDA.n3432 VDDA.n3372 3.4105
R2928 VDDA.n3448 VDDA.n3372 3.4105
R2929 VDDA.n3431 VDDA.n3372 3.4105
R2930 VDDA.n3450 VDDA.n3372 3.4105
R2931 VDDA.n3430 VDDA.n3372 3.4105
R2932 VDDA.n3452 VDDA.n3372 3.4105
R2933 VDDA.n3429 VDDA.n3372 3.4105
R2934 VDDA.n3454 VDDA.n3372 3.4105
R2935 VDDA.n3428 VDDA.n3372 3.4105
R2936 VDDA.n3456 VDDA.n3372 3.4105
R2937 VDDA.n3427 VDDA.n3372 3.4105
R2938 VDDA.n3458 VDDA.n3372 3.4105
R2939 VDDA.n3426 VDDA.n3372 3.4105
R2940 VDDA.n3460 VDDA.n3372 3.4105
R2941 VDDA.n3425 VDDA.n3372 3.4105
R2942 VDDA.n3462 VDDA.n3372 3.4105
R2943 VDDA.n3424 VDDA.n3372 3.4105
R2944 VDDA.n3464 VDDA.n3372 3.4105
R2945 VDDA.n3423 VDDA.n3372 3.4105
R2946 VDDA.n3372 VDDA.n16 3.4105
R2947 VDDA.n3466 VDDA.n3372 3.4105
R2948 VDDA.n3437 VDDA.n3390 3.4105
R2949 VDDA.n3436 VDDA.n3390 3.4105
R2950 VDDA.n3440 VDDA.n3390 3.4105
R2951 VDDA.n3435 VDDA.n3390 3.4105
R2952 VDDA.n3442 VDDA.n3390 3.4105
R2953 VDDA.n3434 VDDA.n3390 3.4105
R2954 VDDA.n3444 VDDA.n3390 3.4105
R2955 VDDA.n3433 VDDA.n3390 3.4105
R2956 VDDA.n3446 VDDA.n3390 3.4105
R2957 VDDA.n3432 VDDA.n3390 3.4105
R2958 VDDA.n3448 VDDA.n3390 3.4105
R2959 VDDA.n3431 VDDA.n3390 3.4105
R2960 VDDA.n3450 VDDA.n3390 3.4105
R2961 VDDA.n3430 VDDA.n3390 3.4105
R2962 VDDA.n3452 VDDA.n3390 3.4105
R2963 VDDA.n3429 VDDA.n3390 3.4105
R2964 VDDA.n3454 VDDA.n3390 3.4105
R2965 VDDA.n3428 VDDA.n3390 3.4105
R2966 VDDA.n3456 VDDA.n3390 3.4105
R2967 VDDA.n3427 VDDA.n3390 3.4105
R2968 VDDA.n3458 VDDA.n3390 3.4105
R2969 VDDA.n3426 VDDA.n3390 3.4105
R2970 VDDA.n3460 VDDA.n3390 3.4105
R2971 VDDA.n3425 VDDA.n3390 3.4105
R2972 VDDA.n3462 VDDA.n3390 3.4105
R2973 VDDA.n3424 VDDA.n3390 3.4105
R2974 VDDA.n3464 VDDA.n3390 3.4105
R2975 VDDA.n3423 VDDA.n3390 3.4105
R2976 VDDA.n3390 VDDA.n16 3.4105
R2977 VDDA.n3466 VDDA.n3390 3.4105
R2978 VDDA.n3437 VDDA.n3371 3.4105
R2979 VDDA.n3436 VDDA.n3371 3.4105
R2980 VDDA.n3440 VDDA.n3371 3.4105
R2981 VDDA.n3435 VDDA.n3371 3.4105
R2982 VDDA.n3442 VDDA.n3371 3.4105
R2983 VDDA.n3434 VDDA.n3371 3.4105
R2984 VDDA.n3444 VDDA.n3371 3.4105
R2985 VDDA.n3433 VDDA.n3371 3.4105
R2986 VDDA.n3446 VDDA.n3371 3.4105
R2987 VDDA.n3432 VDDA.n3371 3.4105
R2988 VDDA.n3448 VDDA.n3371 3.4105
R2989 VDDA.n3431 VDDA.n3371 3.4105
R2990 VDDA.n3450 VDDA.n3371 3.4105
R2991 VDDA.n3430 VDDA.n3371 3.4105
R2992 VDDA.n3452 VDDA.n3371 3.4105
R2993 VDDA.n3429 VDDA.n3371 3.4105
R2994 VDDA.n3454 VDDA.n3371 3.4105
R2995 VDDA.n3428 VDDA.n3371 3.4105
R2996 VDDA.n3456 VDDA.n3371 3.4105
R2997 VDDA.n3427 VDDA.n3371 3.4105
R2998 VDDA.n3458 VDDA.n3371 3.4105
R2999 VDDA.n3426 VDDA.n3371 3.4105
R3000 VDDA.n3460 VDDA.n3371 3.4105
R3001 VDDA.n3425 VDDA.n3371 3.4105
R3002 VDDA.n3462 VDDA.n3371 3.4105
R3003 VDDA.n3424 VDDA.n3371 3.4105
R3004 VDDA.n3464 VDDA.n3371 3.4105
R3005 VDDA.n3423 VDDA.n3371 3.4105
R3006 VDDA.n3371 VDDA.n16 3.4105
R3007 VDDA.n3466 VDDA.n3371 3.4105
R3008 VDDA.n3437 VDDA.n3393 3.4105
R3009 VDDA.n3436 VDDA.n3393 3.4105
R3010 VDDA.n3440 VDDA.n3393 3.4105
R3011 VDDA.n3435 VDDA.n3393 3.4105
R3012 VDDA.n3442 VDDA.n3393 3.4105
R3013 VDDA.n3434 VDDA.n3393 3.4105
R3014 VDDA.n3444 VDDA.n3393 3.4105
R3015 VDDA.n3433 VDDA.n3393 3.4105
R3016 VDDA.n3446 VDDA.n3393 3.4105
R3017 VDDA.n3432 VDDA.n3393 3.4105
R3018 VDDA.n3448 VDDA.n3393 3.4105
R3019 VDDA.n3431 VDDA.n3393 3.4105
R3020 VDDA.n3450 VDDA.n3393 3.4105
R3021 VDDA.n3430 VDDA.n3393 3.4105
R3022 VDDA.n3452 VDDA.n3393 3.4105
R3023 VDDA.n3429 VDDA.n3393 3.4105
R3024 VDDA.n3454 VDDA.n3393 3.4105
R3025 VDDA.n3428 VDDA.n3393 3.4105
R3026 VDDA.n3456 VDDA.n3393 3.4105
R3027 VDDA.n3427 VDDA.n3393 3.4105
R3028 VDDA.n3458 VDDA.n3393 3.4105
R3029 VDDA.n3426 VDDA.n3393 3.4105
R3030 VDDA.n3460 VDDA.n3393 3.4105
R3031 VDDA.n3425 VDDA.n3393 3.4105
R3032 VDDA.n3462 VDDA.n3393 3.4105
R3033 VDDA.n3424 VDDA.n3393 3.4105
R3034 VDDA.n3464 VDDA.n3393 3.4105
R3035 VDDA.n3423 VDDA.n3393 3.4105
R3036 VDDA.n3393 VDDA.n16 3.4105
R3037 VDDA.n3466 VDDA.n3393 3.4105
R3038 VDDA.n3437 VDDA.n3370 3.4105
R3039 VDDA.n3436 VDDA.n3370 3.4105
R3040 VDDA.n3440 VDDA.n3370 3.4105
R3041 VDDA.n3435 VDDA.n3370 3.4105
R3042 VDDA.n3442 VDDA.n3370 3.4105
R3043 VDDA.n3434 VDDA.n3370 3.4105
R3044 VDDA.n3444 VDDA.n3370 3.4105
R3045 VDDA.n3433 VDDA.n3370 3.4105
R3046 VDDA.n3446 VDDA.n3370 3.4105
R3047 VDDA.n3432 VDDA.n3370 3.4105
R3048 VDDA.n3448 VDDA.n3370 3.4105
R3049 VDDA.n3431 VDDA.n3370 3.4105
R3050 VDDA.n3450 VDDA.n3370 3.4105
R3051 VDDA.n3430 VDDA.n3370 3.4105
R3052 VDDA.n3452 VDDA.n3370 3.4105
R3053 VDDA.n3429 VDDA.n3370 3.4105
R3054 VDDA.n3454 VDDA.n3370 3.4105
R3055 VDDA.n3428 VDDA.n3370 3.4105
R3056 VDDA.n3456 VDDA.n3370 3.4105
R3057 VDDA.n3427 VDDA.n3370 3.4105
R3058 VDDA.n3458 VDDA.n3370 3.4105
R3059 VDDA.n3426 VDDA.n3370 3.4105
R3060 VDDA.n3460 VDDA.n3370 3.4105
R3061 VDDA.n3425 VDDA.n3370 3.4105
R3062 VDDA.n3462 VDDA.n3370 3.4105
R3063 VDDA.n3424 VDDA.n3370 3.4105
R3064 VDDA.n3464 VDDA.n3370 3.4105
R3065 VDDA.n3423 VDDA.n3370 3.4105
R3066 VDDA.n3370 VDDA.n16 3.4105
R3067 VDDA.n3466 VDDA.n3370 3.4105
R3068 VDDA.n3437 VDDA.n3396 3.4105
R3069 VDDA.n3436 VDDA.n3396 3.4105
R3070 VDDA.n3440 VDDA.n3396 3.4105
R3071 VDDA.n3435 VDDA.n3396 3.4105
R3072 VDDA.n3442 VDDA.n3396 3.4105
R3073 VDDA.n3434 VDDA.n3396 3.4105
R3074 VDDA.n3444 VDDA.n3396 3.4105
R3075 VDDA.n3433 VDDA.n3396 3.4105
R3076 VDDA.n3446 VDDA.n3396 3.4105
R3077 VDDA.n3432 VDDA.n3396 3.4105
R3078 VDDA.n3448 VDDA.n3396 3.4105
R3079 VDDA.n3431 VDDA.n3396 3.4105
R3080 VDDA.n3450 VDDA.n3396 3.4105
R3081 VDDA.n3430 VDDA.n3396 3.4105
R3082 VDDA.n3452 VDDA.n3396 3.4105
R3083 VDDA.n3429 VDDA.n3396 3.4105
R3084 VDDA.n3454 VDDA.n3396 3.4105
R3085 VDDA.n3428 VDDA.n3396 3.4105
R3086 VDDA.n3456 VDDA.n3396 3.4105
R3087 VDDA.n3427 VDDA.n3396 3.4105
R3088 VDDA.n3458 VDDA.n3396 3.4105
R3089 VDDA.n3426 VDDA.n3396 3.4105
R3090 VDDA.n3460 VDDA.n3396 3.4105
R3091 VDDA.n3425 VDDA.n3396 3.4105
R3092 VDDA.n3462 VDDA.n3396 3.4105
R3093 VDDA.n3424 VDDA.n3396 3.4105
R3094 VDDA.n3464 VDDA.n3396 3.4105
R3095 VDDA.n3423 VDDA.n3396 3.4105
R3096 VDDA.n3396 VDDA.n16 3.4105
R3097 VDDA.n3466 VDDA.n3396 3.4105
R3098 VDDA.n3437 VDDA.n3369 3.4105
R3099 VDDA.n3436 VDDA.n3369 3.4105
R3100 VDDA.n3440 VDDA.n3369 3.4105
R3101 VDDA.n3435 VDDA.n3369 3.4105
R3102 VDDA.n3442 VDDA.n3369 3.4105
R3103 VDDA.n3434 VDDA.n3369 3.4105
R3104 VDDA.n3444 VDDA.n3369 3.4105
R3105 VDDA.n3433 VDDA.n3369 3.4105
R3106 VDDA.n3446 VDDA.n3369 3.4105
R3107 VDDA.n3432 VDDA.n3369 3.4105
R3108 VDDA.n3448 VDDA.n3369 3.4105
R3109 VDDA.n3431 VDDA.n3369 3.4105
R3110 VDDA.n3450 VDDA.n3369 3.4105
R3111 VDDA.n3430 VDDA.n3369 3.4105
R3112 VDDA.n3452 VDDA.n3369 3.4105
R3113 VDDA.n3429 VDDA.n3369 3.4105
R3114 VDDA.n3454 VDDA.n3369 3.4105
R3115 VDDA.n3428 VDDA.n3369 3.4105
R3116 VDDA.n3456 VDDA.n3369 3.4105
R3117 VDDA.n3427 VDDA.n3369 3.4105
R3118 VDDA.n3458 VDDA.n3369 3.4105
R3119 VDDA.n3426 VDDA.n3369 3.4105
R3120 VDDA.n3460 VDDA.n3369 3.4105
R3121 VDDA.n3425 VDDA.n3369 3.4105
R3122 VDDA.n3462 VDDA.n3369 3.4105
R3123 VDDA.n3424 VDDA.n3369 3.4105
R3124 VDDA.n3464 VDDA.n3369 3.4105
R3125 VDDA.n3423 VDDA.n3369 3.4105
R3126 VDDA.n3369 VDDA.n16 3.4105
R3127 VDDA.n3466 VDDA.n3369 3.4105
R3128 VDDA.n3437 VDDA.n3399 3.4105
R3129 VDDA.n3436 VDDA.n3399 3.4105
R3130 VDDA.n3440 VDDA.n3399 3.4105
R3131 VDDA.n3435 VDDA.n3399 3.4105
R3132 VDDA.n3442 VDDA.n3399 3.4105
R3133 VDDA.n3434 VDDA.n3399 3.4105
R3134 VDDA.n3444 VDDA.n3399 3.4105
R3135 VDDA.n3433 VDDA.n3399 3.4105
R3136 VDDA.n3446 VDDA.n3399 3.4105
R3137 VDDA.n3432 VDDA.n3399 3.4105
R3138 VDDA.n3448 VDDA.n3399 3.4105
R3139 VDDA.n3431 VDDA.n3399 3.4105
R3140 VDDA.n3450 VDDA.n3399 3.4105
R3141 VDDA.n3430 VDDA.n3399 3.4105
R3142 VDDA.n3452 VDDA.n3399 3.4105
R3143 VDDA.n3429 VDDA.n3399 3.4105
R3144 VDDA.n3454 VDDA.n3399 3.4105
R3145 VDDA.n3428 VDDA.n3399 3.4105
R3146 VDDA.n3456 VDDA.n3399 3.4105
R3147 VDDA.n3427 VDDA.n3399 3.4105
R3148 VDDA.n3458 VDDA.n3399 3.4105
R3149 VDDA.n3426 VDDA.n3399 3.4105
R3150 VDDA.n3460 VDDA.n3399 3.4105
R3151 VDDA.n3425 VDDA.n3399 3.4105
R3152 VDDA.n3462 VDDA.n3399 3.4105
R3153 VDDA.n3424 VDDA.n3399 3.4105
R3154 VDDA.n3464 VDDA.n3399 3.4105
R3155 VDDA.n3423 VDDA.n3399 3.4105
R3156 VDDA.n3399 VDDA.n16 3.4105
R3157 VDDA.n3466 VDDA.n3399 3.4105
R3158 VDDA.n3437 VDDA.n3368 3.4105
R3159 VDDA.n3436 VDDA.n3368 3.4105
R3160 VDDA.n3440 VDDA.n3368 3.4105
R3161 VDDA.n3435 VDDA.n3368 3.4105
R3162 VDDA.n3442 VDDA.n3368 3.4105
R3163 VDDA.n3434 VDDA.n3368 3.4105
R3164 VDDA.n3444 VDDA.n3368 3.4105
R3165 VDDA.n3433 VDDA.n3368 3.4105
R3166 VDDA.n3446 VDDA.n3368 3.4105
R3167 VDDA.n3432 VDDA.n3368 3.4105
R3168 VDDA.n3448 VDDA.n3368 3.4105
R3169 VDDA.n3431 VDDA.n3368 3.4105
R3170 VDDA.n3450 VDDA.n3368 3.4105
R3171 VDDA.n3430 VDDA.n3368 3.4105
R3172 VDDA.n3452 VDDA.n3368 3.4105
R3173 VDDA.n3429 VDDA.n3368 3.4105
R3174 VDDA.n3454 VDDA.n3368 3.4105
R3175 VDDA.n3428 VDDA.n3368 3.4105
R3176 VDDA.n3456 VDDA.n3368 3.4105
R3177 VDDA.n3427 VDDA.n3368 3.4105
R3178 VDDA.n3458 VDDA.n3368 3.4105
R3179 VDDA.n3426 VDDA.n3368 3.4105
R3180 VDDA.n3460 VDDA.n3368 3.4105
R3181 VDDA.n3425 VDDA.n3368 3.4105
R3182 VDDA.n3462 VDDA.n3368 3.4105
R3183 VDDA.n3424 VDDA.n3368 3.4105
R3184 VDDA.n3464 VDDA.n3368 3.4105
R3185 VDDA.n3423 VDDA.n3368 3.4105
R3186 VDDA.n3368 VDDA.n16 3.4105
R3187 VDDA.n3466 VDDA.n3368 3.4105
R3188 VDDA.n3437 VDDA.n3402 3.4105
R3189 VDDA.n3436 VDDA.n3402 3.4105
R3190 VDDA.n3440 VDDA.n3402 3.4105
R3191 VDDA.n3435 VDDA.n3402 3.4105
R3192 VDDA.n3442 VDDA.n3402 3.4105
R3193 VDDA.n3434 VDDA.n3402 3.4105
R3194 VDDA.n3444 VDDA.n3402 3.4105
R3195 VDDA.n3433 VDDA.n3402 3.4105
R3196 VDDA.n3446 VDDA.n3402 3.4105
R3197 VDDA.n3432 VDDA.n3402 3.4105
R3198 VDDA.n3448 VDDA.n3402 3.4105
R3199 VDDA.n3431 VDDA.n3402 3.4105
R3200 VDDA.n3450 VDDA.n3402 3.4105
R3201 VDDA.n3430 VDDA.n3402 3.4105
R3202 VDDA.n3452 VDDA.n3402 3.4105
R3203 VDDA.n3429 VDDA.n3402 3.4105
R3204 VDDA.n3454 VDDA.n3402 3.4105
R3205 VDDA.n3428 VDDA.n3402 3.4105
R3206 VDDA.n3456 VDDA.n3402 3.4105
R3207 VDDA.n3427 VDDA.n3402 3.4105
R3208 VDDA.n3458 VDDA.n3402 3.4105
R3209 VDDA.n3426 VDDA.n3402 3.4105
R3210 VDDA.n3460 VDDA.n3402 3.4105
R3211 VDDA.n3425 VDDA.n3402 3.4105
R3212 VDDA.n3462 VDDA.n3402 3.4105
R3213 VDDA.n3424 VDDA.n3402 3.4105
R3214 VDDA.n3464 VDDA.n3402 3.4105
R3215 VDDA.n3423 VDDA.n3402 3.4105
R3216 VDDA.n3402 VDDA.n16 3.4105
R3217 VDDA.n3466 VDDA.n3402 3.4105
R3218 VDDA.n3437 VDDA.n3367 3.4105
R3219 VDDA.n3436 VDDA.n3367 3.4105
R3220 VDDA.n3440 VDDA.n3367 3.4105
R3221 VDDA.n3435 VDDA.n3367 3.4105
R3222 VDDA.n3442 VDDA.n3367 3.4105
R3223 VDDA.n3434 VDDA.n3367 3.4105
R3224 VDDA.n3444 VDDA.n3367 3.4105
R3225 VDDA.n3433 VDDA.n3367 3.4105
R3226 VDDA.n3446 VDDA.n3367 3.4105
R3227 VDDA.n3432 VDDA.n3367 3.4105
R3228 VDDA.n3448 VDDA.n3367 3.4105
R3229 VDDA.n3431 VDDA.n3367 3.4105
R3230 VDDA.n3450 VDDA.n3367 3.4105
R3231 VDDA.n3430 VDDA.n3367 3.4105
R3232 VDDA.n3452 VDDA.n3367 3.4105
R3233 VDDA.n3429 VDDA.n3367 3.4105
R3234 VDDA.n3454 VDDA.n3367 3.4105
R3235 VDDA.n3428 VDDA.n3367 3.4105
R3236 VDDA.n3456 VDDA.n3367 3.4105
R3237 VDDA.n3427 VDDA.n3367 3.4105
R3238 VDDA.n3458 VDDA.n3367 3.4105
R3239 VDDA.n3426 VDDA.n3367 3.4105
R3240 VDDA.n3460 VDDA.n3367 3.4105
R3241 VDDA.n3425 VDDA.n3367 3.4105
R3242 VDDA.n3462 VDDA.n3367 3.4105
R3243 VDDA.n3424 VDDA.n3367 3.4105
R3244 VDDA.n3464 VDDA.n3367 3.4105
R3245 VDDA.n3423 VDDA.n3367 3.4105
R3246 VDDA.n3367 VDDA.n16 3.4105
R3247 VDDA.n3466 VDDA.n3367 3.4105
R3248 VDDA.n3437 VDDA.n3405 3.4105
R3249 VDDA.n3436 VDDA.n3405 3.4105
R3250 VDDA.n3440 VDDA.n3405 3.4105
R3251 VDDA.n3435 VDDA.n3405 3.4105
R3252 VDDA.n3442 VDDA.n3405 3.4105
R3253 VDDA.n3434 VDDA.n3405 3.4105
R3254 VDDA.n3444 VDDA.n3405 3.4105
R3255 VDDA.n3433 VDDA.n3405 3.4105
R3256 VDDA.n3446 VDDA.n3405 3.4105
R3257 VDDA.n3432 VDDA.n3405 3.4105
R3258 VDDA.n3448 VDDA.n3405 3.4105
R3259 VDDA.n3431 VDDA.n3405 3.4105
R3260 VDDA.n3450 VDDA.n3405 3.4105
R3261 VDDA.n3430 VDDA.n3405 3.4105
R3262 VDDA.n3452 VDDA.n3405 3.4105
R3263 VDDA.n3429 VDDA.n3405 3.4105
R3264 VDDA.n3454 VDDA.n3405 3.4105
R3265 VDDA.n3428 VDDA.n3405 3.4105
R3266 VDDA.n3456 VDDA.n3405 3.4105
R3267 VDDA.n3427 VDDA.n3405 3.4105
R3268 VDDA.n3458 VDDA.n3405 3.4105
R3269 VDDA.n3426 VDDA.n3405 3.4105
R3270 VDDA.n3460 VDDA.n3405 3.4105
R3271 VDDA.n3425 VDDA.n3405 3.4105
R3272 VDDA.n3462 VDDA.n3405 3.4105
R3273 VDDA.n3424 VDDA.n3405 3.4105
R3274 VDDA.n3464 VDDA.n3405 3.4105
R3275 VDDA.n3423 VDDA.n3405 3.4105
R3276 VDDA.n3405 VDDA.n16 3.4105
R3277 VDDA.n3466 VDDA.n3405 3.4105
R3278 VDDA.n3437 VDDA.n3366 3.4105
R3279 VDDA.n3436 VDDA.n3366 3.4105
R3280 VDDA.n3440 VDDA.n3366 3.4105
R3281 VDDA.n3435 VDDA.n3366 3.4105
R3282 VDDA.n3442 VDDA.n3366 3.4105
R3283 VDDA.n3434 VDDA.n3366 3.4105
R3284 VDDA.n3444 VDDA.n3366 3.4105
R3285 VDDA.n3433 VDDA.n3366 3.4105
R3286 VDDA.n3446 VDDA.n3366 3.4105
R3287 VDDA.n3432 VDDA.n3366 3.4105
R3288 VDDA.n3448 VDDA.n3366 3.4105
R3289 VDDA.n3431 VDDA.n3366 3.4105
R3290 VDDA.n3450 VDDA.n3366 3.4105
R3291 VDDA.n3430 VDDA.n3366 3.4105
R3292 VDDA.n3452 VDDA.n3366 3.4105
R3293 VDDA.n3429 VDDA.n3366 3.4105
R3294 VDDA.n3454 VDDA.n3366 3.4105
R3295 VDDA.n3428 VDDA.n3366 3.4105
R3296 VDDA.n3456 VDDA.n3366 3.4105
R3297 VDDA.n3427 VDDA.n3366 3.4105
R3298 VDDA.n3458 VDDA.n3366 3.4105
R3299 VDDA.n3426 VDDA.n3366 3.4105
R3300 VDDA.n3460 VDDA.n3366 3.4105
R3301 VDDA.n3425 VDDA.n3366 3.4105
R3302 VDDA.n3462 VDDA.n3366 3.4105
R3303 VDDA.n3424 VDDA.n3366 3.4105
R3304 VDDA.n3464 VDDA.n3366 3.4105
R3305 VDDA.n3423 VDDA.n3366 3.4105
R3306 VDDA.n3366 VDDA.n16 3.4105
R3307 VDDA.n3466 VDDA.n3366 3.4105
R3308 VDDA.n3437 VDDA.n3408 3.4105
R3309 VDDA.n3436 VDDA.n3408 3.4105
R3310 VDDA.n3440 VDDA.n3408 3.4105
R3311 VDDA.n3435 VDDA.n3408 3.4105
R3312 VDDA.n3442 VDDA.n3408 3.4105
R3313 VDDA.n3434 VDDA.n3408 3.4105
R3314 VDDA.n3444 VDDA.n3408 3.4105
R3315 VDDA.n3433 VDDA.n3408 3.4105
R3316 VDDA.n3446 VDDA.n3408 3.4105
R3317 VDDA.n3432 VDDA.n3408 3.4105
R3318 VDDA.n3448 VDDA.n3408 3.4105
R3319 VDDA.n3431 VDDA.n3408 3.4105
R3320 VDDA.n3450 VDDA.n3408 3.4105
R3321 VDDA.n3430 VDDA.n3408 3.4105
R3322 VDDA.n3452 VDDA.n3408 3.4105
R3323 VDDA.n3429 VDDA.n3408 3.4105
R3324 VDDA.n3454 VDDA.n3408 3.4105
R3325 VDDA.n3428 VDDA.n3408 3.4105
R3326 VDDA.n3456 VDDA.n3408 3.4105
R3327 VDDA.n3427 VDDA.n3408 3.4105
R3328 VDDA.n3458 VDDA.n3408 3.4105
R3329 VDDA.n3426 VDDA.n3408 3.4105
R3330 VDDA.n3460 VDDA.n3408 3.4105
R3331 VDDA.n3425 VDDA.n3408 3.4105
R3332 VDDA.n3462 VDDA.n3408 3.4105
R3333 VDDA.n3424 VDDA.n3408 3.4105
R3334 VDDA.n3464 VDDA.n3408 3.4105
R3335 VDDA.n3423 VDDA.n3408 3.4105
R3336 VDDA.n3408 VDDA.n16 3.4105
R3337 VDDA.n3466 VDDA.n3408 3.4105
R3338 VDDA.n3437 VDDA.n3365 3.4105
R3339 VDDA.n3436 VDDA.n3365 3.4105
R3340 VDDA.n3440 VDDA.n3365 3.4105
R3341 VDDA.n3435 VDDA.n3365 3.4105
R3342 VDDA.n3442 VDDA.n3365 3.4105
R3343 VDDA.n3434 VDDA.n3365 3.4105
R3344 VDDA.n3444 VDDA.n3365 3.4105
R3345 VDDA.n3433 VDDA.n3365 3.4105
R3346 VDDA.n3446 VDDA.n3365 3.4105
R3347 VDDA.n3432 VDDA.n3365 3.4105
R3348 VDDA.n3448 VDDA.n3365 3.4105
R3349 VDDA.n3431 VDDA.n3365 3.4105
R3350 VDDA.n3450 VDDA.n3365 3.4105
R3351 VDDA.n3430 VDDA.n3365 3.4105
R3352 VDDA.n3452 VDDA.n3365 3.4105
R3353 VDDA.n3429 VDDA.n3365 3.4105
R3354 VDDA.n3454 VDDA.n3365 3.4105
R3355 VDDA.n3428 VDDA.n3365 3.4105
R3356 VDDA.n3456 VDDA.n3365 3.4105
R3357 VDDA.n3427 VDDA.n3365 3.4105
R3358 VDDA.n3458 VDDA.n3365 3.4105
R3359 VDDA.n3426 VDDA.n3365 3.4105
R3360 VDDA.n3460 VDDA.n3365 3.4105
R3361 VDDA.n3425 VDDA.n3365 3.4105
R3362 VDDA.n3462 VDDA.n3365 3.4105
R3363 VDDA.n3424 VDDA.n3365 3.4105
R3364 VDDA.n3464 VDDA.n3365 3.4105
R3365 VDDA.n3423 VDDA.n3365 3.4105
R3366 VDDA.n3365 VDDA.n16 3.4105
R3367 VDDA.n3466 VDDA.n3365 3.4105
R3368 VDDA.n3437 VDDA.n3411 3.4105
R3369 VDDA.n3436 VDDA.n3411 3.4105
R3370 VDDA.n3440 VDDA.n3411 3.4105
R3371 VDDA.n3435 VDDA.n3411 3.4105
R3372 VDDA.n3442 VDDA.n3411 3.4105
R3373 VDDA.n3434 VDDA.n3411 3.4105
R3374 VDDA.n3444 VDDA.n3411 3.4105
R3375 VDDA.n3433 VDDA.n3411 3.4105
R3376 VDDA.n3446 VDDA.n3411 3.4105
R3377 VDDA.n3432 VDDA.n3411 3.4105
R3378 VDDA.n3448 VDDA.n3411 3.4105
R3379 VDDA.n3431 VDDA.n3411 3.4105
R3380 VDDA.n3450 VDDA.n3411 3.4105
R3381 VDDA.n3430 VDDA.n3411 3.4105
R3382 VDDA.n3452 VDDA.n3411 3.4105
R3383 VDDA.n3429 VDDA.n3411 3.4105
R3384 VDDA.n3454 VDDA.n3411 3.4105
R3385 VDDA.n3428 VDDA.n3411 3.4105
R3386 VDDA.n3456 VDDA.n3411 3.4105
R3387 VDDA.n3427 VDDA.n3411 3.4105
R3388 VDDA.n3458 VDDA.n3411 3.4105
R3389 VDDA.n3426 VDDA.n3411 3.4105
R3390 VDDA.n3460 VDDA.n3411 3.4105
R3391 VDDA.n3425 VDDA.n3411 3.4105
R3392 VDDA.n3462 VDDA.n3411 3.4105
R3393 VDDA.n3424 VDDA.n3411 3.4105
R3394 VDDA.n3464 VDDA.n3411 3.4105
R3395 VDDA.n3423 VDDA.n3411 3.4105
R3396 VDDA.n3411 VDDA.n16 3.4105
R3397 VDDA.n3466 VDDA.n3411 3.4105
R3398 VDDA.n3437 VDDA.n3364 3.4105
R3399 VDDA.n3436 VDDA.n3364 3.4105
R3400 VDDA.n3440 VDDA.n3364 3.4105
R3401 VDDA.n3435 VDDA.n3364 3.4105
R3402 VDDA.n3442 VDDA.n3364 3.4105
R3403 VDDA.n3434 VDDA.n3364 3.4105
R3404 VDDA.n3444 VDDA.n3364 3.4105
R3405 VDDA.n3433 VDDA.n3364 3.4105
R3406 VDDA.n3446 VDDA.n3364 3.4105
R3407 VDDA.n3432 VDDA.n3364 3.4105
R3408 VDDA.n3448 VDDA.n3364 3.4105
R3409 VDDA.n3431 VDDA.n3364 3.4105
R3410 VDDA.n3450 VDDA.n3364 3.4105
R3411 VDDA.n3430 VDDA.n3364 3.4105
R3412 VDDA.n3452 VDDA.n3364 3.4105
R3413 VDDA.n3429 VDDA.n3364 3.4105
R3414 VDDA.n3454 VDDA.n3364 3.4105
R3415 VDDA.n3428 VDDA.n3364 3.4105
R3416 VDDA.n3456 VDDA.n3364 3.4105
R3417 VDDA.n3427 VDDA.n3364 3.4105
R3418 VDDA.n3458 VDDA.n3364 3.4105
R3419 VDDA.n3426 VDDA.n3364 3.4105
R3420 VDDA.n3460 VDDA.n3364 3.4105
R3421 VDDA.n3425 VDDA.n3364 3.4105
R3422 VDDA.n3462 VDDA.n3364 3.4105
R3423 VDDA.n3424 VDDA.n3364 3.4105
R3424 VDDA.n3464 VDDA.n3364 3.4105
R3425 VDDA.n3423 VDDA.n3364 3.4105
R3426 VDDA.n3364 VDDA.n16 3.4105
R3427 VDDA.n3466 VDDA.n3364 3.4105
R3428 VDDA.n3437 VDDA.n3414 3.4105
R3429 VDDA.n3436 VDDA.n3414 3.4105
R3430 VDDA.n3440 VDDA.n3414 3.4105
R3431 VDDA.n3435 VDDA.n3414 3.4105
R3432 VDDA.n3442 VDDA.n3414 3.4105
R3433 VDDA.n3434 VDDA.n3414 3.4105
R3434 VDDA.n3444 VDDA.n3414 3.4105
R3435 VDDA.n3433 VDDA.n3414 3.4105
R3436 VDDA.n3446 VDDA.n3414 3.4105
R3437 VDDA.n3432 VDDA.n3414 3.4105
R3438 VDDA.n3448 VDDA.n3414 3.4105
R3439 VDDA.n3431 VDDA.n3414 3.4105
R3440 VDDA.n3450 VDDA.n3414 3.4105
R3441 VDDA.n3430 VDDA.n3414 3.4105
R3442 VDDA.n3452 VDDA.n3414 3.4105
R3443 VDDA.n3429 VDDA.n3414 3.4105
R3444 VDDA.n3454 VDDA.n3414 3.4105
R3445 VDDA.n3428 VDDA.n3414 3.4105
R3446 VDDA.n3456 VDDA.n3414 3.4105
R3447 VDDA.n3427 VDDA.n3414 3.4105
R3448 VDDA.n3458 VDDA.n3414 3.4105
R3449 VDDA.n3426 VDDA.n3414 3.4105
R3450 VDDA.n3460 VDDA.n3414 3.4105
R3451 VDDA.n3425 VDDA.n3414 3.4105
R3452 VDDA.n3462 VDDA.n3414 3.4105
R3453 VDDA.n3424 VDDA.n3414 3.4105
R3454 VDDA.n3464 VDDA.n3414 3.4105
R3455 VDDA.n3423 VDDA.n3414 3.4105
R3456 VDDA.n3414 VDDA.n16 3.4105
R3457 VDDA.n3466 VDDA.n3414 3.4105
R3458 VDDA.n3437 VDDA.n3363 3.4105
R3459 VDDA.n3436 VDDA.n3363 3.4105
R3460 VDDA.n3440 VDDA.n3363 3.4105
R3461 VDDA.n3435 VDDA.n3363 3.4105
R3462 VDDA.n3442 VDDA.n3363 3.4105
R3463 VDDA.n3434 VDDA.n3363 3.4105
R3464 VDDA.n3444 VDDA.n3363 3.4105
R3465 VDDA.n3433 VDDA.n3363 3.4105
R3466 VDDA.n3446 VDDA.n3363 3.4105
R3467 VDDA.n3432 VDDA.n3363 3.4105
R3468 VDDA.n3448 VDDA.n3363 3.4105
R3469 VDDA.n3431 VDDA.n3363 3.4105
R3470 VDDA.n3450 VDDA.n3363 3.4105
R3471 VDDA.n3430 VDDA.n3363 3.4105
R3472 VDDA.n3452 VDDA.n3363 3.4105
R3473 VDDA.n3429 VDDA.n3363 3.4105
R3474 VDDA.n3454 VDDA.n3363 3.4105
R3475 VDDA.n3428 VDDA.n3363 3.4105
R3476 VDDA.n3456 VDDA.n3363 3.4105
R3477 VDDA.n3427 VDDA.n3363 3.4105
R3478 VDDA.n3458 VDDA.n3363 3.4105
R3479 VDDA.n3426 VDDA.n3363 3.4105
R3480 VDDA.n3460 VDDA.n3363 3.4105
R3481 VDDA.n3425 VDDA.n3363 3.4105
R3482 VDDA.n3462 VDDA.n3363 3.4105
R3483 VDDA.n3424 VDDA.n3363 3.4105
R3484 VDDA.n3464 VDDA.n3363 3.4105
R3485 VDDA.n3423 VDDA.n3363 3.4105
R3486 VDDA.n3363 VDDA.n16 3.4105
R3487 VDDA.n3466 VDDA.n3363 3.4105
R3488 VDDA.n3437 VDDA.n3417 3.4105
R3489 VDDA.n3436 VDDA.n3417 3.4105
R3490 VDDA.n3440 VDDA.n3417 3.4105
R3491 VDDA.n3435 VDDA.n3417 3.4105
R3492 VDDA.n3442 VDDA.n3417 3.4105
R3493 VDDA.n3434 VDDA.n3417 3.4105
R3494 VDDA.n3444 VDDA.n3417 3.4105
R3495 VDDA.n3433 VDDA.n3417 3.4105
R3496 VDDA.n3446 VDDA.n3417 3.4105
R3497 VDDA.n3432 VDDA.n3417 3.4105
R3498 VDDA.n3448 VDDA.n3417 3.4105
R3499 VDDA.n3431 VDDA.n3417 3.4105
R3500 VDDA.n3450 VDDA.n3417 3.4105
R3501 VDDA.n3430 VDDA.n3417 3.4105
R3502 VDDA.n3452 VDDA.n3417 3.4105
R3503 VDDA.n3429 VDDA.n3417 3.4105
R3504 VDDA.n3454 VDDA.n3417 3.4105
R3505 VDDA.n3428 VDDA.n3417 3.4105
R3506 VDDA.n3456 VDDA.n3417 3.4105
R3507 VDDA.n3427 VDDA.n3417 3.4105
R3508 VDDA.n3458 VDDA.n3417 3.4105
R3509 VDDA.n3426 VDDA.n3417 3.4105
R3510 VDDA.n3460 VDDA.n3417 3.4105
R3511 VDDA.n3425 VDDA.n3417 3.4105
R3512 VDDA.n3462 VDDA.n3417 3.4105
R3513 VDDA.n3424 VDDA.n3417 3.4105
R3514 VDDA.n3464 VDDA.n3417 3.4105
R3515 VDDA.n3423 VDDA.n3417 3.4105
R3516 VDDA.n3417 VDDA.n16 3.4105
R3517 VDDA.n3466 VDDA.n3417 3.4105
R3518 VDDA.n3437 VDDA.n3362 3.4105
R3519 VDDA.n3436 VDDA.n3362 3.4105
R3520 VDDA.n3440 VDDA.n3362 3.4105
R3521 VDDA.n3435 VDDA.n3362 3.4105
R3522 VDDA.n3442 VDDA.n3362 3.4105
R3523 VDDA.n3434 VDDA.n3362 3.4105
R3524 VDDA.n3444 VDDA.n3362 3.4105
R3525 VDDA.n3433 VDDA.n3362 3.4105
R3526 VDDA.n3446 VDDA.n3362 3.4105
R3527 VDDA.n3432 VDDA.n3362 3.4105
R3528 VDDA.n3448 VDDA.n3362 3.4105
R3529 VDDA.n3431 VDDA.n3362 3.4105
R3530 VDDA.n3450 VDDA.n3362 3.4105
R3531 VDDA.n3430 VDDA.n3362 3.4105
R3532 VDDA.n3452 VDDA.n3362 3.4105
R3533 VDDA.n3429 VDDA.n3362 3.4105
R3534 VDDA.n3454 VDDA.n3362 3.4105
R3535 VDDA.n3428 VDDA.n3362 3.4105
R3536 VDDA.n3456 VDDA.n3362 3.4105
R3537 VDDA.n3427 VDDA.n3362 3.4105
R3538 VDDA.n3458 VDDA.n3362 3.4105
R3539 VDDA.n3426 VDDA.n3362 3.4105
R3540 VDDA.n3460 VDDA.n3362 3.4105
R3541 VDDA.n3425 VDDA.n3362 3.4105
R3542 VDDA.n3462 VDDA.n3362 3.4105
R3543 VDDA.n3424 VDDA.n3362 3.4105
R3544 VDDA.n3464 VDDA.n3362 3.4105
R3545 VDDA.n3423 VDDA.n3362 3.4105
R3546 VDDA.n3362 VDDA.n16 3.4105
R3547 VDDA.n3466 VDDA.n3362 3.4105
R3548 VDDA.n3437 VDDA.n3420 3.4105
R3549 VDDA.n3436 VDDA.n3420 3.4105
R3550 VDDA.n3440 VDDA.n3420 3.4105
R3551 VDDA.n3435 VDDA.n3420 3.4105
R3552 VDDA.n3442 VDDA.n3420 3.4105
R3553 VDDA.n3434 VDDA.n3420 3.4105
R3554 VDDA.n3444 VDDA.n3420 3.4105
R3555 VDDA.n3433 VDDA.n3420 3.4105
R3556 VDDA.n3446 VDDA.n3420 3.4105
R3557 VDDA.n3432 VDDA.n3420 3.4105
R3558 VDDA.n3448 VDDA.n3420 3.4105
R3559 VDDA.n3431 VDDA.n3420 3.4105
R3560 VDDA.n3450 VDDA.n3420 3.4105
R3561 VDDA.n3430 VDDA.n3420 3.4105
R3562 VDDA.n3452 VDDA.n3420 3.4105
R3563 VDDA.n3429 VDDA.n3420 3.4105
R3564 VDDA.n3454 VDDA.n3420 3.4105
R3565 VDDA.n3428 VDDA.n3420 3.4105
R3566 VDDA.n3456 VDDA.n3420 3.4105
R3567 VDDA.n3427 VDDA.n3420 3.4105
R3568 VDDA.n3458 VDDA.n3420 3.4105
R3569 VDDA.n3426 VDDA.n3420 3.4105
R3570 VDDA.n3460 VDDA.n3420 3.4105
R3571 VDDA.n3425 VDDA.n3420 3.4105
R3572 VDDA.n3462 VDDA.n3420 3.4105
R3573 VDDA.n3424 VDDA.n3420 3.4105
R3574 VDDA.n3464 VDDA.n3420 3.4105
R3575 VDDA.n3423 VDDA.n3420 3.4105
R3576 VDDA.n3420 VDDA.n16 3.4105
R3577 VDDA.n3466 VDDA.n3420 3.4105
R3578 VDDA.n3437 VDDA.n3361 3.4105
R3579 VDDA.n3436 VDDA.n3361 3.4105
R3580 VDDA.n3440 VDDA.n3361 3.4105
R3581 VDDA.n3435 VDDA.n3361 3.4105
R3582 VDDA.n3442 VDDA.n3361 3.4105
R3583 VDDA.n3434 VDDA.n3361 3.4105
R3584 VDDA.n3444 VDDA.n3361 3.4105
R3585 VDDA.n3433 VDDA.n3361 3.4105
R3586 VDDA.n3446 VDDA.n3361 3.4105
R3587 VDDA.n3432 VDDA.n3361 3.4105
R3588 VDDA.n3448 VDDA.n3361 3.4105
R3589 VDDA.n3431 VDDA.n3361 3.4105
R3590 VDDA.n3450 VDDA.n3361 3.4105
R3591 VDDA.n3430 VDDA.n3361 3.4105
R3592 VDDA.n3452 VDDA.n3361 3.4105
R3593 VDDA.n3429 VDDA.n3361 3.4105
R3594 VDDA.n3454 VDDA.n3361 3.4105
R3595 VDDA.n3428 VDDA.n3361 3.4105
R3596 VDDA.n3456 VDDA.n3361 3.4105
R3597 VDDA.n3427 VDDA.n3361 3.4105
R3598 VDDA.n3458 VDDA.n3361 3.4105
R3599 VDDA.n3426 VDDA.n3361 3.4105
R3600 VDDA.n3460 VDDA.n3361 3.4105
R3601 VDDA.n3425 VDDA.n3361 3.4105
R3602 VDDA.n3462 VDDA.n3361 3.4105
R3603 VDDA.n3424 VDDA.n3361 3.4105
R3604 VDDA.n3464 VDDA.n3361 3.4105
R3605 VDDA.n3423 VDDA.n3361 3.4105
R3606 VDDA.n3361 VDDA.n16 3.4105
R3607 VDDA.n3466 VDDA.n3361 3.4105
R3608 VDDA.n3465 VDDA.n3436 3.4105
R3609 VDDA.n3465 VDDA.n3440 3.4105
R3610 VDDA.n3465 VDDA.n3435 3.4105
R3611 VDDA.n3465 VDDA.n3442 3.4105
R3612 VDDA.n3465 VDDA.n3434 3.4105
R3613 VDDA.n3465 VDDA.n3444 3.4105
R3614 VDDA.n3465 VDDA.n3433 3.4105
R3615 VDDA.n3465 VDDA.n3446 3.4105
R3616 VDDA.n3465 VDDA.n3432 3.4105
R3617 VDDA.n3465 VDDA.n3448 3.4105
R3618 VDDA.n3465 VDDA.n3431 3.4105
R3619 VDDA.n3465 VDDA.n3450 3.4105
R3620 VDDA.n3465 VDDA.n3430 3.4105
R3621 VDDA.n3465 VDDA.n3452 3.4105
R3622 VDDA.n3465 VDDA.n3429 3.4105
R3623 VDDA.n3465 VDDA.n3454 3.4105
R3624 VDDA.n3465 VDDA.n3428 3.4105
R3625 VDDA.n3465 VDDA.n3456 3.4105
R3626 VDDA.n3465 VDDA.n3427 3.4105
R3627 VDDA.n3465 VDDA.n3458 3.4105
R3628 VDDA.n3465 VDDA.n3426 3.4105
R3629 VDDA.n3465 VDDA.n3460 3.4105
R3630 VDDA.n3465 VDDA.n3425 3.4105
R3631 VDDA.n3465 VDDA.n3462 3.4105
R3632 VDDA.n3465 VDDA.n3424 3.4105
R3633 VDDA.n3465 VDDA.n3464 3.4105
R3634 VDDA.n3465 VDDA.n3423 3.4105
R3635 VDDA.n3465 VDDA.n16 3.4105
R3636 VDDA.n3466 VDDA.n3465 3.4105
R3637 VDDA.n2034 VDDA.n2033 3.10304
R3638 VDDA.n2763 VDDA.n2762 2.8957
R3639 VDDA.n2764 VDDA.n2763 2.8957
R3640 VDDA.n2768 VDDA.n2766 2.8957
R3641 VDDA.n2771 VDDA.n2766 2.8957
R3642 VDDA.n2767 VDDA.n2764 2.8957
R3643 VDDA.n2771 VDDA.n2770 2.8957
R3644 VDDA.n2773 VDDA.n2762 2.8957
R3645 VDDA.n2768 VDDA.n2767 2.8957
R3646 VDDA.n2802 VDDA.n2801 2.8255
R3647 VDDA.n2800 VDDA.n2799 2.8255
R3648 VDDA.n2856 VDDA.n2855 2.65454
R3649 VDDA.n2698 VDDA.n2682 2.65418
R3650 VDDA.n2820 VDDA.n2819 2.423
R3651 VDDA.n2818 VDDA.n2817 2.423
R3652 VDDA.n2713 VDDA.n2712 2.423
R3653 VDDA.n2711 VDDA.n2710 2.423
R3654 VDDA.n2334 VDDA.n2333 2.39683
R3655 VDDA.n2149 VDDA.n2148 2.39683
R3656 VDDA.n352 VDDA.n351 2.39683
R3657 VDDA.n2675 VDDA.n2674 2.39683
R3658 VDDA.n2530 VDDA.n2529 2.39683
R3659 VDDA.n2773 VDDA.n2761 2.32777
R3660 VDDA.n91 VDDA.n90 2.30736
R3661 VDDA.n3238 VDDA.n3235 2.30736
R3662 VDDA.n3093 VDDA.n3092 2.30736
R3663 VDDA.n2934 VDDA.n2933 2.30736
R3664 VDDA.n428 VDDA.n427 2.30736
R3665 VDDA.n1734 VDDA.n1733 2.30736
R3666 VDDA.n1575 VDDA.n1574 2.30736
R3667 VDDA.n595 VDDA.n594 2.30736
R3668 VDDA.n1378 VDDA.n1375 2.30736
R3669 VDDA.n1214 VDDA.n1213 2.30736
R3670 VDDA.n2558 VDDA.n2557 2.251
R3671 VDDA.n1497 VDDA.n517 2.18322
R3672 VDDA.n3190 VDDA.n180 2.18322
R3673 VDDA.n2836 VDDA.n2835 1.97758
R3674 VDDA.n2834 VDDA.n2833 1.97758
R3675 VDDA.n2729 VDDA.n2728 1.97758
R3676 VDDA.n2727 VDDA.n2726 1.97758
R3677 VDDA.n2559 VDDA.n2558 1.93785
R3678 VDDA.n2795 VDDA.n2794 1.888
R3679 VDDA.n2793 VDDA.n2792 1.888
R3680 VDDA.n2219 VDDA.n2218 1.71668
R3681 VDDA.n3376 VDDA.n0 1.70567
R3682 VDDA.n3379 VDDA.n3376 1.70567
R3683 VDDA.n3382 VDDA.n3376 1.70567
R3684 VDDA.n3385 VDDA.n3376 1.70567
R3685 VDDA.n3388 VDDA.n3376 1.70567
R3686 VDDA.n3391 VDDA.n3376 1.70567
R3687 VDDA.n3394 VDDA.n3376 1.70567
R3688 VDDA.n3397 VDDA.n3376 1.70567
R3689 VDDA.n3400 VDDA.n3376 1.70567
R3690 VDDA.n3403 VDDA.n3376 1.70567
R3691 VDDA.n3406 VDDA.n3376 1.70567
R3692 VDDA.n3409 VDDA.n3376 1.70567
R3693 VDDA.n3412 VDDA.n3376 1.70567
R3694 VDDA.n3415 VDDA.n3376 1.70567
R3695 VDDA.n3418 VDDA.n3376 1.70567
R3696 VDDA.n3421 VDDA.n3376 1.70567
R3697 VDDA.n3467 VDDA.n14 1.70565
R3698 VDDA.n3467 VDDA.n12 1.70565
R3699 VDDA.n3467 VDDA.n10 1.70565
R3700 VDDA.n3467 VDDA.n8 1.70565
R3701 VDDA.n3467 VDDA.n6 1.70565
R3702 VDDA.n3467 VDDA.n4 1.70565
R3703 VDDA.n3467 VDDA.n2 1.70565
R3704 VDDA.n3443 VDDA.n3378 1.70565
R3705 VDDA.n3445 VDDA.n3378 1.70565
R3706 VDDA.n3451 VDDA.n3378 1.70565
R3707 VDDA.n3453 VDDA.n3378 1.70565
R3708 VDDA.n3459 VDDA.n3378 1.70565
R3709 VDDA.n3461 VDDA.n3378 1.70565
R3710 VDDA.n3465 VDDA.n3438 1.70565
R3711 VDDA.n3467 VDDA.n13 1.70563
R3712 VDDA.n3467 VDDA.n9 1.70563
R3713 VDDA.n3467 VDDA.n5 1.70563
R3714 VDDA.n3467 VDDA.n1 1.70563
R3715 VDDA.n3439 VDDA.n3378 1.70563
R3716 VDDA.n3441 VDDA.n3378 1.70563
R3717 VDDA.n3447 VDDA.n3378 1.70563
R3718 VDDA.n3449 VDDA.n3378 1.70563
R3719 VDDA.n3455 VDDA.n3378 1.70563
R3720 VDDA.n3457 VDDA.n3378 1.70563
R3721 VDDA.n3463 VDDA.n3378 1.70563
R3722 VDDA.n3422 VDDA.n3378 1.70563
R3723 VDDA.n3377 VDDA.n15 1.70563
R3724 VDDA.n3383 VDDA.n15 1.70563
R3725 VDDA.n3389 VDDA.n15 1.70563
R3726 VDDA.n3395 VDDA.n15 1.70563
R3727 VDDA.n3401 VDDA.n15 1.70563
R3728 VDDA.n3407 VDDA.n15 1.70563
R3729 VDDA.n3413 VDDA.n15 1.70563
R3730 VDDA.n3419 VDDA.n15 1.70563
R3731 VDDA.n3467 VDDA.n11 1.70556
R3732 VDDA.n3467 VDDA.n7 1.70556
R3733 VDDA.n3467 VDDA.n3 1.70556
R3734 VDDA.n3380 VDDA.n15 1.70556
R3735 VDDA.n3386 VDDA.n15 1.70556
R3736 VDDA.n3392 VDDA.n15 1.70556
R3737 VDDA.n3398 VDDA.n15 1.70556
R3738 VDDA.n3404 VDDA.n15 1.70556
R3739 VDDA.n3410 VDDA.n15 1.70556
R3740 VDDA.n3416 VDDA.n15 1.70556
R3741 VDDA.n1327 VDDA.n1189 1.69433
R3742 VDDA.n1327 VDDA.n1186 1.69433
R3743 VDDA.n1327 VDDA.n1183 1.69433
R3744 VDDA.n1327 VDDA.n1180 1.69433
R3745 VDDA.n1327 VDDA.n1177 1.69433
R3746 VDDA.n1327 VDDA.n1174 1.69433
R3747 VDDA.n1327 VDDA.n1171 1.69433
R3748 VDDA.n1481 VDDA.n521 1.69433
R3749 VDDA.n1463 VDDA.n521 1.69433
R3750 VDDA.n1451 VDDA.n521 1.69433
R3751 VDDA.n1433 VDDA.n521 1.69433
R3752 VDDA.n1421 VDDA.n521 1.69433
R3753 VDDA.n1403 VDDA.n521 1.69433
R3754 VDDA.n1391 VDDA.n521 1.69433
R3755 VDDA.n1501 VDDA.n543 1.69433
R3756 VDDA.n1501 VDDA.n540 1.69433
R3757 VDDA.n1501 VDDA.n537 1.69433
R3758 VDDA.n1501 VDDA.n534 1.69433
R3759 VDDA.n1501 VDDA.n531 1.69433
R3760 VDDA.n1501 VDDA.n528 1.69433
R3761 VDDA.n1501 VDDA.n525 1.69433
R3762 VDDA.n1667 VDDA.n1523 1.69433
R3763 VDDA.n1667 VDDA.n1520 1.69433
R3764 VDDA.n1667 VDDA.n1517 1.69433
R3765 VDDA.n1667 VDDA.n1514 1.69433
R3766 VDDA.n1667 VDDA.n1511 1.69433
R3767 VDDA.n1667 VDDA.n1508 1.69433
R3768 VDDA.n1667 VDDA.n1505 1.69433
R3769 VDDA.n2678 VDDA.n1689 1.69433
R3770 VDDA.n2678 VDDA.n1686 1.69433
R3771 VDDA.n2678 VDDA.n1683 1.69433
R3772 VDDA.n2678 VDDA.n1680 1.69433
R3773 VDDA.n2678 VDDA.n1677 1.69433
R3774 VDDA.n2678 VDDA.n1674 1.69433
R3775 VDDA.n2678 VDDA.n1671 1.69433
R3776 VDDA.n2860 VDDA.n376 1.69433
R3777 VDDA.n2860 VDDA.n373 1.69433
R3778 VDDA.n2860 VDDA.n370 1.69433
R3779 VDDA.n2860 VDDA.n367 1.69433
R3780 VDDA.n2860 VDDA.n364 1.69433
R3781 VDDA.n2860 VDDA.n361 1.69433
R3782 VDDA.n2860 VDDA.n358 1.69433
R3783 VDDA.n3026 VDDA.n2882 1.69433
R3784 VDDA.n3026 VDDA.n2879 1.69433
R3785 VDDA.n3026 VDDA.n2876 1.69433
R3786 VDDA.n3026 VDDA.n2873 1.69433
R3787 VDDA.n3026 VDDA.n2870 1.69433
R3788 VDDA.n3026 VDDA.n2867 1.69433
R3789 VDDA.n3026 VDDA.n2864 1.69433
R3790 VDDA.n3186 VDDA.n3048 1.69433
R3791 VDDA.n3186 VDDA.n3045 1.69433
R3792 VDDA.n3186 VDDA.n3042 1.69433
R3793 VDDA.n3186 VDDA.n3039 1.69433
R3794 VDDA.n3186 VDDA.n3036 1.69433
R3795 VDDA.n3186 VDDA.n3033 1.69433
R3796 VDDA.n3186 VDDA.n3030 1.69433
R3797 VDDA.n3341 VDDA.n17 1.69433
R3798 VDDA.n3323 VDDA.n17 1.69433
R3799 VDDA.n3311 VDDA.n17 1.69433
R3800 VDDA.n3293 VDDA.n17 1.69433
R3801 VDDA.n3281 VDDA.n17 1.69433
R3802 VDDA.n3263 VDDA.n17 1.69433
R3803 VDDA.n3251 VDDA.n17 1.69433
R3804 VDDA.n3360 VDDA.n39 1.69433
R3805 VDDA.n3360 VDDA.n36 1.69433
R3806 VDDA.n3360 VDDA.n33 1.69433
R3807 VDDA.n3360 VDDA.n30 1.69433
R3808 VDDA.n3360 VDDA.n27 1.69433
R3809 VDDA.n3360 VDDA.n24 1.69433
R3810 VDDA.n3360 VDDA.n21 1.69433
R3811 VDDA.n2532 VDDA.n1872 1.69433
R3812 VDDA.n2532 VDDA.n1869 1.69433
R3813 VDDA.n2532 VDDA.n1866 1.69433
R3814 VDDA.n2532 VDDA.n1863 1.69433
R3815 VDDA.n2532 VDDA.n1860 1.69433
R3816 VDDA.n2532 VDDA.n1857 1.69433
R3817 VDDA.n2532 VDDA.n1854 1.69433
R3818 VDDA.n2677 VDDA.n1848 1.69433
R3819 VDDA.n2677 VDDA.n1845 1.69433
R3820 VDDA.n2677 VDDA.n1842 1.69433
R3821 VDDA.n2677 VDDA.n1839 1.69433
R3822 VDDA.n2677 VDDA.n1836 1.69433
R3823 VDDA.n2677 VDDA.n1833 1.69433
R3824 VDDA.n2677 VDDA.n1830 1.69433
R3825 VDDA.n354 VDDA.n205 1.69433
R3826 VDDA.n354 VDDA.n202 1.69433
R3827 VDDA.n354 VDDA.n199 1.69433
R3828 VDDA.n354 VDDA.n196 1.69433
R3829 VDDA.n354 VDDA.n193 1.69433
R3830 VDDA.n354 VDDA.n190 1.69433
R3831 VDDA.n354 VDDA.n187 1.69433
R3832 VDDA.n2151 VDDA.n1920 1.69433
R3833 VDDA.n2151 VDDA.n1917 1.69433
R3834 VDDA.n2151 VDDA.n1914 1.69433
R3835 VDDA.n2151 VDDA.n1911 1.69433
R3836 VDDA.n2151 VDDA.n1908 1.69433
R3837 VDDA.n2151 VDDA.n1905 1.69433
R3838 VDDA.n2151 VDDA.n1902 1.69433
R3839 VDDA.n2336 VDDA.n1896 1.69433
R3840 VDDA.n2336 VDDA.n1893 1.69433
R3841 VDDA.n2336 VDDA.n1890 1.69433
R3842 VDDA.n2336 VDDA.n1887 1.69433
R3843 VDDA.n2336 VDDA.n1884 1.69433
R3844 VDDA.n2336 VDDA.n1881 1.69433
R3845 VDDA.n2336 VDDA.n1878 1.69433
R3846 VDDA.n1327 VDDA.n1326 1.6924
R3847 VDDA.n1327 VDDA.n1190 1.6924
R3848 VDDA.n1327 VDDA.n1188 1.6924
R3849 VDDA.n1327 VDDA.n1187 1.6924
R3850 VDDA.n1327 VDDA.n1185 1.6924
R3851 VDDA.n1327 VDDA.n1184 1.6924
R3852 VDDA.n1327 VDDA.n1182 1.6924
R3853 VDDA.n1327 VDDA.n1181 1.6924
R3854 VDDA.n1327 VDDA.n1179 1.6924
R3855 VDDA.n1327 VDDA.n1178 1.6924
R3856 VDDA.n1327 VDDA.n1176 1.6924
R3857 VDDA.n1327 VDDA.n1175 1.6924
R3858 VDDA.n1327 VDDA.n1173 1.6924
R3859 VDDA.n1327 VDDA.n1172 1.6924
R3860 VDDA.n1327 VDDA.n1170 1.6924
R3861 VDDA.n1327 VDDA.n1169 1.6924
R3862 VDDA.n1491 VDDA.n521 1.6924
R3863 VDDA.n1483 VDDA.n521 1.6924
R3864 VDDA.n1473 VDDA.n521 1.6924
R3865 VDDA.n1471 VDDA.n521 1.6924
R3866 VDDA.n1461 VDDA.n521 1.6924
R3867 VDDA.n1453 VDDA.n521 1.6924
R3868 VDDA.n1443 VDDA.n521 1.6924
R3869 VDDA.n1441 VDDA.n521 1.6924
R3870 VDDA.n1431 VDDA.n521 1.6924
R3871 VDDA.n1423 VDDA.n521 1.6924
R3872 VDDA.n1413 VDDA.n521 1.6924
R3873 VDDA.n1411 VDDA.n521 1.6924
R3874 VDDA.n1401 VDDA.n521 1.6924
R3875 VDDA.n1393 VDDA.n521 1.6924
R3876 VDDA.n1383 VDDA.n521 1.6924
R3877 VDDA.n1381 VDDA.n521 1.6924
R3878 VDDA.n1501 VDDA.n545 1.6924
R3879 VDDA.n1501 VDDA.n544 1.6924
R3880 VDDA.n1501 VDDA.n542 1.6924
R3881 VDDA.n1501 VDDA.n541 1.6924
R3882 VDDA.n1501 VDDA.n539 1.6924
R3883 VDDA.n1501 VDDA.n538 1.6924
R3884 VDDA.n1501 VDDA.n536 1.6924
R3885 VDDA.n1501 VDDA.n535 1.6924
R3886 VDDA.n1501 VDDA.n533 1.6924
R3887 VDDA.n1501 VDDA.n532 1.6924
R3888 VDDA.n1501 VDDA.n530 1.6924
R3889 VDDA.n1501 VDDA.n529 1.6924
R3890 VDDA.n1501 VDDA.n527 1.6924
R3891 VDDA.n1501 VDDA.n526 1.6924
R3892 VDDA.n1501 VDDA.n524 1.6924
R3893 VDDA.n1501 VDDA.n523 1.6924
R3894 VDDA.n1667 VDDA.n1525 1.6924
R3895 VDDA.n1667 VDDA.n1524 1.6924
R3896 VDDA.n1667 VDDA.n1522 1.6924
R3897 VDDA.n1667 VDDA.n1521 1.6924
R3898 VDDA.n1667 VDDA.n1519 1.6924
R3899 VDDA.n1667 VDDA.n1518 1.6924
R3900 VDDA.n1667 VDDA.n1516 1.6924
R3901 VDDA.n1667 VDDA.n1515 1.6924
R3902 VDDA.n1667 VDDA.n1513 1.6924
R3903 VDDA.n1667 VDDA.n1512 1.6924
R3904 VDDA.n1667 VDDA.n1510 1.6924
R3905 VDDA.n1667 VDDA.n1509 1.6924
R3906 VDDA.n1667 VDDA.n1507 1.6924
R3907 VDDA.n1667 VDDA.n1506 1.6924
R3908 VDDA.n1667 VDDA.n1504 1.6924
R3909 VDDA.n1667 VDDA.n1503 1.6924
R3910 VDDA.n2678 VDDA.n1826 1.6924
R3911 VDDA.n2678 VDDA.n1690 1.6924
R3912 VDDA.n2678 VDDA.n1688 1.6924
R3913 VDDA.n2678 VDDA.n1687 1.6924
R3914 VDDA.n2678 VDDA.n1685 1.6924
R3915 VDDA.n2678 VDDA.n1684 1.6924
R3916 VDDA.n2678 VDDA.n1682 1.6924
R3917 VDDA.n2678 VDDA.n1681 1.6924
R3918 VDDA.n2678 VDDA.n1679 1.6924
R3919 VDDA.n2678 VDDA.n1678 1.6924
R3920 VDDA.n2678 VDDA.n1676 1.6924
R3921 VDDA.n2678 VDDA.n1675 1.6924
R3922 VDDA.n2678 VDDA.n1673 1.6924
R3923 VDDA.n2678 VDDA.n1672 1.6924
R3924 VDDA.n2678 VDDA.n1670 1.6924
R3925 VDDA.n2678 VDDA.n1669 1.6924
R3926 VDDA.n2860 VDDA.n378 1.6924
R3927 VDDA.n2860 VDDA.n377 1.6924
R3928 VDDA.n2860 VDDA.n375 1.6924
R3929 VDDA.n2860 VDDA.n374 1.6924
R3930 VDDA.n2860 VDDA.n372 1.6924
R3931 VDDA.n2860 VDDA.n371 1.6924
R3932 VDDA.n2860 VDDA.n369 1.6924
R3933 VDDA.n2860 VDDA.n368 1.6924
R3934 VDDA.n2860 VDDA.n366 1.6924
R3935 VDDA.n2860 VDDA.n365 1.6924
R3936 VDDA.n2860 VDDA.n363 1.6924
R3937 VDDA.n2860 VDDA.n362 1.6924
R3938 VDDA.n2860 VDDA.n360 1.6924
R3939 VDDA.n2860 VDDA.n359 1.6924
R3940 VDDA.n2860 VDDA.n357 1.6924
R3941 VDDA.n2860 VDDA.n356 1.6924
R3942 VDDA.n3026 VDDA.n2884 1.6924
R3943 VDDA.n3026 VDDA.n2883 1.6924
R3944 VDDA.n3026 VDDA.n2881 1.6924
R3945 VDDA.n3026 VDDA.n2880 1.6924
R3946 VDDA.n3026 VDDA.n2878 1.6924
R3947 VDDA.n3026 VDDA.n2877 1.6924
R3948 VDDA.n3026 VDDA.n2875 1.6924
R3949 VDDA.n3026 VDDA.n2874 1.6924
R3950 VDDA.n3026 VDDA.n2872 1.6924
R3951 VDDA.n3026 VDDA.n2871 1.6924
R3952 VDDA.n3026 VDDA.n2869 1.6924
R3953 VDDA.n3026 VDDA.n2868 1.6924
R3954 VDDA.n3026 VDDA.n2866 1.6924
R3955 VDDA.n3026 VDDA.n2865 1.6924
R3956 VDDA.n3026 VDDA.n2863 1.6924
R3957 VDDA.n3026 VDDA.n2862 1.6924
R3958 VDDA.n3186 VDDA.n3185 1.6924
R3959 VDDA.n3186 VDDA.n3049 1.6924
R3960 VDDA.n3186 VDDA.n3047 1.6924
R3961 VDDA.n3186 VDDA.n3046 1.6924
R3962 VDDA.n3186 VDDA.n3044 1.6924
R3963 VDDA.n3186 VDDA.n3043 1.6924
R3964 VDDA.n3186 VDDA.n3041 1.6924
R3965 VDDA.n3186 VDDA.n3040 1.6924
R3966 VDDA.n3186 VDDA.n3038 1.6924
R3967 VDDA.n3186 VDDA.n3037 1.6924
R3968 VDDA.n3186 VDDA.n3035 1.6924
R3969 VDDA.n3186 VDDA.n3034 1.6924
R3970 VDDA.n3186 VDDA.n3032 1.6924
R3971 VDDA.n3186 VDDA.n3031 1.6924
R3972 VDDA.n3186 VDDA.n3029 1.6924
R3973 VDDA.n3186 VDDA.n3028 1.6924
R3974 VDDA.n3351 VDDA.n17 1.6924
R3975 VDDA.n3343 VDDA.n17 1.6924
R3976 VDDA.n3333 VDDA.n17 1.6924
R3977 VDDA.n3331 VDDA.n17 1.6924
R3978 VDDA.n3321 VDDA.n17 1.6924
R3979 VDDA.n3313 VDDA.n17 1.6924
R3980 VDDA.n3303 VDDA.n17 1.6924
R3981 VDDA.n3301 VDDA.n17 1.6924
R3982 VDDA.n3291 VDDA.n17 1.6924
R3983 VDDA.n3283 VDDA.n17 1.6924
R3984 VDDA.n3273 VDDA.n17 1.6924
R3985 VDDA.n3271 VDDA.n17 1.6924
R3986 VDDA.n3261 VDDA.n17 1.6924
R3987 VDDA.n3253 VDDA.n17 1.6924
R3988 VDDA.n3243 VDDA.n17 1.6924
R3989 VDDA.n3241 VDDA.n17 1.6924
R3990 VDDA.n3360 VDDA.n41 1.6924
R3991 VDDA.n3360 VDDA.n40 1.6924
R3992 VDDA.n3360 VDDA.n38 1.6924
R3993 VDDA.n3360 VDDA.n37 1.6924
R3994 VDDA.n3360 VDDA.n35 1.6924
R3995 VDDA.n3360 VDDA.n34 1.6924
R3996 VDDA.n3360 VDDA.n32 1.6924
R3997 VDDA.n3360 VDDA.n31 1.6924
R3998 VDDA.n3360 VDDA.n29 1.6924
R3999 VDDA.n3360 VDDA.n28 1.6924
R4000 VDDA.n3360 VDDA.n26 1.6924
R4001 VDDA.n3360 VDDA.n25 1.6924
R4002 VDDA.n3360 VDDA.n23 1.6924
R4003 VDDA.n3360 VDDA.n22 1.6924
R4004 VDDA.n3360 VDDA.n20 1.6924
R4005 VDDA.n3360 VDDA.n19 1.6924
R4006 VDDA.n2532 VDDA.n1874 1.6924
R4007 VDDA.n2532 VDDA.n1873 1.6924
R4008 VDDA.n2532 VDDA.n1871 1.6924
R4009 VDDA.n2532 VDDA.n1870 1.6924
R4010 VDDA.n2532 VDDA.n1868 1.6924
R4011 VDDA.n2532 VDDA.n1867 1.6924
R4012 VDDA.n2532 VDDA.n1865 1.6924
R4013 VDDA.n2532 VDDA.n1864 1.6924
R4014 VDDA.n2532 VDDA.n1862 1.6924
R4015 VDDA.n2532 VDDA.n1861 1.6924
R4016 VDDA.n2532 VDDA.n1859 1.6924
R4017 VDDA.n2532 VDDA.n1858 1.6924
R4018 VDDA.n2532 VDDA.n1856 1.6924
R4019 VDDA.n2532 VDDA.n1855 1.6924
R4020 VDDA.n2532 VDDA.n1853 1.6924
R4021 VDDA.n2532 VDDA.n1852 1.6924
R4022 VDDA.n2677 VDDA.n1850 1.6924
R4023 VDDA.n2677 VDDA.n1849 1.6924
R4024 VDDA.n2677 VDDA.n1847 1.6924
R4025 VDDA.n2677 VDDA.n1846 1.6924
R4026 VDDA.n2677 VDDA.n1844 1.6924
R4027 VDDA.n2677 VDDA.n1843 1.6924
R4028 VDDA.n2677 VDDA.n1841 1.6924
R4029 VDDA.n2677 VDDA.n1840 1.6924
R4030 VDDA.n2677 VDDA.n1838 1.6924
R4031 VDDA.n2677 VDDA.n1837 1.6924
R4032 VDDA.n2677 VDDA.n1835 1.6924
R4033 VDDA.n2677 VDDA.n1834 1.6924
R4034 VDDA.n2677 VDDA.n1832 1.6924
R4035 VDDA.n2677 VDDA.n1831 1.6924
R4036 VDDA.n2677 VDDA.n1829 1.6924
R4037 VDDA.n2677 VDDA.n1828 1.6924
R4038 VDDA.n354 VDDA.n207 1.6924
R4039 VDDA.n354 VDDA.n206 1.6924
R4040 VDDA.n354 VDDA.n204 1.6924
R4041 VDDA.n354 VDDA.n203 1.6924
R4042 VDDA.n354 VDDA.n201 1.6924
R4043 VDDA.n354 VDDA.n200 1.6924
R4044 VDDA.n354 VDDA.n198 1.6924
R4045 VDDA.n354 VDDA.n197 1.6924
R4046 VDDA.n354 VDDA.n195 1.6924
R4047 VDDA.n354 VDDA.n194 1.6924
R4048 VDDA.n354 VDDA.n192 1.6924
R4049 VDDA.n354 VDDA.n191 1.6924
R4050 VDDA.n354 VDDA.n189 1.6924
R4051 VDDA.n354 VDDA.n188 1.6924
R4052 VDDA.n354 VDDA.n186 1.6924
R4053 VDDA.n354 VDDA.n185 1.6924
R4054 VDDA.n2151 VDDA.n1922 1.6924
R4055 VDDA.n2151 VDDA.n1921 1.6924
R4056 VDDA.n2151 VDDA.n1919 1.6924
R4057 VDDA.n2151 VDDA.n1918 1.6924
R4058 VDDA.n2151 VDDA.n1916 1.6924
R4059 VDDA.n2151 VDDA.n1915 1.6924
R4060 VDDA.n2151 VDDA.n1913 1.6924
R4061 VDDA.n2151 VDDA.n1912 1.6924
R4062 VDDA.n2151 VDDA.n1910 1.6924
R4063 VDDA.n2151 VDDA.n1909 1.6924
R4064 VDDA.n2151 VDDA.n1907 1.6924
R4065 VDDA.n2151 VDDA.n1906 1.6924
R4066 VDDA.n2151 VDDA.n1904 1.6924
R4067 VDDA.n2151 VDDA.n1903 1.6924
R4068 VDDA.n2151 VDDA.n1901 1.6924
R4069 VDDA.n2151 VDDA.n1900 1.6924
R4070 VDDA.n2336 VDDA.n1898 1.6924
R4071 VDDA.n2336 VDDA.n1897 1.6924
R4072 VDDA.n2336 VDDA.n1895 1.6924
R4073 VDDA.n2336 VDDA.n1894 1.6924
R4074 VDDA.n2336 VDDA.n1892 1.6924
R4075 VDDA.n2336 VDDA.n1891 1.6924
R4076 VDDA.n2336 VDDA.n1889 1.6924
R4077 VDDA.n2336 VDDA.n1888 1.6924
R4078 VDDA.n2336 VDDA.n1886 1.6924
R4079 VDDA.n2336 VDDA.n1885 1.6924
R4080 VDDA.n2336 VDDA.n1883 1.6924
R4081 VDDA.n2336 VDDA.n1882 1.6924
R4082 VDDA.n2336 VDDA.n1880 1.6924
R4083 VDDA.n2336 VDDA.n1879 1.6924
R4084 VDDA.n2336 VDDA.n1877 1.6924
R4085 VDDA.n2336 VDDA.n1876 1.6924
R4086 VDDA.n2787 VDDA.n2730 1.5005
R4087 VDDA.n2218 VDDA.n2217 1.44719
R4088 VDDA.n2789 VDDA.n2698 1.438
R4089 VDDA.n2855 VDDA.n2839 1.438
R4090 VDDA.n1497 VDDA.n1496 1.08947
R4091 VDDA.n2682 VDDA.n517 1.08947
R4092 VDDA.n2856 VDDA.n180 1.08947
R4093 VDDA.n3356 VDDA.n3190 1.08947
R4094 VDDA.n2033 VDDA.n2031 1.05183
R4095 VDDA.n2848 VDDA.n2847 1.03383
R4096 VDDA.n2846 VDDA.n2845 1.03383
R4097 VDDA.n2691 VDDA.n2690 1.03383
R4098 VDDA.n2689 VDDA.n2688 1.03383
R4099 VDDA.n2759 VDDA.n2758 0.922375
R4100 VDDA.n2741 VDDA.n2732 0.922375
R4101 VDDA.n2786 VDDA.n2732 0.922375
R4102 VDDA.n2803 VDDA.n2798 0.6255
R4103 VDDA.n2796 VDDA.n2790 0.6255
R4104 VDDA.n2853 VDDA.n2852 0.6255
R4105 VDDA.n2852 VDDA.n2850 0.6255
R4106 VDDA.n2844 VDDA.n2842 0.6255
R4107 VDDA.n2853 VDDA.n2842 0.6255
R4108 VDDA.n2696 VDDA.n2695 0.6255
R4109 VDDA.n2695 VDDA.n2693 0.6255
R4110 VDDA.n2687 VDDA.n2685 0.6255
R4111 VDDA.n2696 VDDA.n2685 0.6255
R4112 VDDA.n2832 VDDA.n2830 0.563
R4113 VDDA.n2830 VDDA.n2828 0.563
R4114 VDDA.n2828 VDDA.n2826 0.563
R4115 VDDA.n2826 VDDA.n2824 0.563
R4116 VDDA.n2837 VDDA.n2824 0.563
R4117 VDDA.n2810 VDDA.n2808 0.563
R4118 VDDA.n2812 VDDA.n2810 0.563
R4119 VDDA.n2814 VDDA.n2812 0.563
R4120 VDDA.n2816 VDDA.n2814 0.563
R4121 VDDA.n2725 VDDA.n2723 0.563
R4122 VDDA.n2723 VDDA.n2721 0.563
R4123 VDDA.n2721 VDDA.n2719 0.563
R4124 VDDA.n2719 VDDA.n2717 0.563
R4125 VDDA.n2730 VDDA.n2717 0.563
R4126 VDDA.n2703 VDDA.n2701 0.563
R4127 VDDA.n2705 VDDA.n2703 0.563
R4128 VDDA.n2707 VDDA.n2705 0.563
R4129 VDDA.n2709 VDDA.n2707 0.563
R4130 VDDA.n2759 VDDA.n2741 0.3755
R4131 VDDA.n2408 VDDA.n2407 0.333833
R4132 VDDA.n688 VDDA.n687 0.3295
R4133 VDDA.n689 VDDA.n688 0.3295
R4134 VDDA.n690 VDDA.n689 0.3295
R4135 VDDA.n691 VDDA.n690 0.3295
R4136 VDDA.n692 VDDA.n691 0.3295
R4137 VDDA.n693 VDDA.n692 0.3295
R4138 VDDA.n701 VDDA.n693 0.3295
R4139 VDDA.n701 VDDA.n700 0.3295
R4140 VDDA.n700 VDDA.n699 0.3295
R4141 VDDA.n699 VDDA.n698 0.3295
R4142 VDDA.n698 VDDA.n697 0.3295
R4143 VDDA.n697 VDDA.n696 0.3295
R4144 VDDA.n696 VDDA.n695 0.3295
R4145 VDDA.n695 VDDA.n694 0.3295
R4146 VDDA.n703 VDDA.n702 0.3295
R4147 VDDA.n704 VDDA.n703 0.3295
R4148 VDDA.n705 VDDA.n704 0.3295
R4149 VDDA.n706 VDDA.n705 0.3295
R4150 VDDA.n707 VDDA.n706 0.3295
R4151 VDDA.n708 VDDA.n707 0.3295
R4152 VDDA.n716 VDDA.n708 0.3295
R4153 VDDA.n716 VDDA.n715 0.3295
R4154 VDDA.n715 VDDA.n714 0.3295
R4155 VDDA.n714 VDDA.n713 0.3295
R4156 VDDA.n713 VDDA.n712 0.3295
R4157 VDDA.n712 VDDA.n711 0.3295
R4158 VDDA.n711 VDDA.n710 0.3295
R4159 VDDA.n710 VDDA.n709 0.3295
R4160 VDDA.n718 VDDA.n717 0.3295
R4161 VDDA.n719 VDDA.n718 0.3295
R4162 VDDA.n720 VDDA.n719 0.3295
R4163 VDDA.n721 VDDA.n720 0.3295
R4164 VDDA.n722 VDDA.n721 0.3295
R4165 VDDA.n723 VDDA.n722 0.3295
R4166 VDDA.n731 VDDA.n723 0.3295
R4167 VDDA.n731 VDDA.n730 0.3295
R4168 VDDA.n730 VDDA.n729 0.3295
R4169 VDDA.n729 VDDA.n728 0.3295
R4170 VDDA.n728 VDDA.n727 0.3295
R4171 VDDA.n727 VDDA.n726 0.3295
R4172 VDDA.n726 VDDA.n725 0.3295
R4173 VDDA.n725 VDDA.n724 0.3295
R4174 VDDA.n733 VDDA.n732 0.3295
R4175 VDDA.n734 VDDA.n733 0.3295
R4176 VDDA.n735 VDDA.n734 0.3295
R4177 VDDA.n736 VDDA.n735 0.3295
R4178 VDDA.n737 VDDA.n736 0.3295
R4179 VDDA.n738 VDDA.n737 0.3295
R4180 VDDA.n746 VDDA.n738 0.3295
R4181 VDDA.n746 VDDA.n745 0.3295
R4182 VDDA.n745 VDDA.n744 0.3295
R4183 VDDA.n744 VDDA.n743 0.3295
R4184 VDDA.n743 VDDA.n742 0.3295
R4185 VDDA.n742 VDDA.n741 0.3295
R4186 VDDA.n741 VDDA.n740 0.3295
R4187 VDDA.n740 VDDA.n739 0.3295
R4188 VDDA.n748 VDDA.n747 0.3295
R4189 VDDA.n749 VDDA.n748 0.3295
R4190 VDDA.n750 VDDA.n749 0.3295
R4191 VDDA.n751 VDDA.n750 0.3295
R4192 VDDA.n752 VDDA.n751 0.3295
R4193 VDDA.n753 VDDA.n752 0.3295
R4194 VDDA.n761 VDDA.n753 0.3295
R4195 VDDA.n761 VDDA.n760 0.3295
R4196 VDDA.n760 VDDA.n759 0.3295
R4197 VDDA.n759 VDDA.n758 0.3295
R4198 VDDA.n758 VDDA.n757 0.3295
R4199 VDDA.n757 VDDA.n756 0.3295
R4200 VDDA.n756 VDDA.n755 0.3295
R4201 VDDA.n755 VDDA.n754 0.3295
R4202 VDDA.n763 VDDA.n762 0.3295
R4203 VDDA.n764 VDDA.n763 0.3295
R4204 VDDA.n765 VDDA.n764 0.3295
R4205 VDDA.n766 VDDA.n765 0.3295
R4206 VDDA.n767 VDDA.n766 0.3295
R4207 VDDA.n768 VDDA.n767 0.3295
R4208 VDDA.n776 VDDA.n768 0.3295
R4209 VDDA.n776 VDDA.n775 0.3295
R4210 VDDA.n775 VDDA.n774 0.3295
R4211 VDDA.n774 VDDA.n773 0.3295
R4212 VDDA.n773 VDDA.n772 0.3295
R4213 VDDA.n772 VDDA.n771 0.3295
R4214 VDDA.n771 VDDA.n770 0.3295
R4215 VDDA.n770 VDDA.n769 0.3295
R4216 VDDA.n778 VDDA.n777 0.3295
R4217 VDDA.n779 VDDA.n778 0.3295
R4218 VDDA.n780 VDDA.n779 0.3295
R4219 VDDA.n781 VDDA.n780 0.3295
R4220 VDDA.n782 VDDA.n781 0.3295
R4221 VDDA.n783 VDDA.n782 0.3295
R4222 VDDA.n791 VDDA.n783 0.3295
R4223 VDDA.n791 VDDA.n790 0.3295
R4224 VDDA.n790 VDDA.n789 0.3295
R4225 VDDA.n789 VDDA.n788 0.3295
R4226 VDDA.n788 VDDA.n787 0.3295
R4227 VDDA.n787 VDDA.n786 0.3295
R4228 VDDA.n786 VDDA.n785 0.3295
R4229 VDDA.n785 VDDA.n784 0.3295
R4230 VDDA.n793 VDDA.n792 0.3295
R4231 VDDA.n794 VDDA.n793 0.3295
R4232 VDDA.n795 VDDA.n794 0.3295
R4233 VDDA.n796 VDDA.n795 0.3295
R4234 VDDA.n797 VDDA.n796 0.3295
R4235 VDDA.n798 VDDA.n797 0.3295
R4236 VDDA.n806 VDDA.n798 0.3295
R4237 VDDA.n806 VDDA.n805 0.3295
R4238 VDDA.n805 VDDA.n804 0.3295
R4239 VDDA.n804 VDDA.n803 0.3295
R4240 VDDA.n803 VDDA.n802 0.3295
R4241 VDDA.n802 VDDA.n801 0.3295
R4242 VDDA.n801 VDDA.n800 0.3295
R4243 VDDA.n800 VDDA.n799 0.3295
R4244 VDDA.n808 VDDA.n807 0.3295
R4245 VDDA.n809 VDDA.n808 0.3295
R4246 VDDA.n810 VDDA.n809 0.3295
R4247 VDDA.n811 VDDA.n810 0.3295
R4248 VDDA.n812 VDDA.n811 0.3295
R4249 VDDA.n813 VDDA.n812 0.3295
R4250 VDDA.n821 VDDA.n813 0.3295
R4251 VDDA.n821 VDDA.n820 0.3295
R4252 VDDA.n820 VDDA.n819 0.3295
R4253 VDDA.n819 VDDA.n818 0.3295
R4254 VDDA.n818 VDDA.n817 0.3295
R4255 VDDA.n817 VDDA.n816 0.3295
R4256 VDDA.n816 VDDA.n815 0.3295
R4257 VDDA.n815 VDDA.n814 0.3295
R4258 VDDA.n823 VDDA.n822 0.3295
R4259 VDDA.n824 VDDA.n823 0.3295
R4260 VDDA.n825 VDDA.n824 0.3295
R4261 VDDA.n826 VDDA.n825 0.3295
R4262 VDDA.n827 VDDA.n826 0.3295
R4263 VDDA.n828 VDDA.n827 0.3295
R4264 VDDA.n836 VDDA.n828 0.3295
R4265 VDDA.n836 VDDA.n835 0.3295
R4266 VDDA.n835 VDDA.n834 0.3295
R4267 VDDA.n834 VDDA.n833 0.3295
R4268 VDDA.n833 VDDA.n832 0.3295
R4269 VDDA.n832 VDDA.n831 0.3295
R4270 VDDA.n831 VDDA.n830 0.3295
R4271 VDDA.n830 VDDA.n829 0.3295
R4272 VDDA.n838 VDDA.n837 0.3295
R4273 VDDA.n839 VDDA.n838 0.3295
R4274 VDDA.n840 VDDA.n839 0.3295
R4275 VDDA.n841 VDDA.n840 0.3295
R4276 VDDA.n842 VDDA.n841 0.3295
R4277 VDDA.n843 VDDA.n842 0.3295
R4278 VDDA.n851 VDDA.n843 0.3295
R4279 VDDA.n851 VDDA.n850 0.3295
R4280 VDDA.n850 VDDA.n849 0.3295
R4281 VDDA.n849 VDDA.n848 0.3295
R4282 VDDA.n848 VDDA.n847 0.3295
R4283 VDDA.n847 VDDA.n846 0.3295
R4284 VDDA.n846 VDDA.n845 0.3295
R4285 VDDA.n845 VDDA.n844 0.3295
R4286 VDDA.n853 VDDA.n852 0.3295
R4287 VDDA.n854 VDDA.n853 0.3295
R4288 VDDA.n855 VDDA.n854 0.3295
R4289 VDDA.n856 VDDA.n855 0.3295
R4290 VDDA.n857 VDDA.n856 0.3295
R4291 VDDA.n858 VDDA.n857 0.3295
R4292 VDDA.n866 VDDA.n858 0.3295
R4293 VDDA.n866 VDDA.n865 0.3295
R4294 VDDA.n865 VDDA.n864 0.3295
R4295 VDDA.n864 VDDA.n863 0.3295
R4296 VDDA.n863 VDDA.n862 0.3295
R4297 VDDA.n862 VDDA.n861 0.3295
R4298 VDDA.n861 VDDA.n860 0.3295
R4299 VDDA.n860 VDDA.n859 0.3295
R4300 VDDA.n868 VDDA.n867 0.3295
R4301 VDDA.n869 VDDA.n868 0.3295
R4302 VDDA.n870 VDDA.n869 0.3295
R4303 VDDA.n871 VDDA.n870 0.3295
R4304 VDDA.n872 VDDA.n871 0.3295
R4305 VDDA.n873 VDDA.n872 0.3295
R4306 VDDA.n881 VDDA.n873 0.3295
R4307 VDDA.n881 VDDA.n880 0.3295
R4308 VDDA.n880 VDDA.n879 0.3295
R4309 VDDA.n879 VDDA.n878 0.3295
R4310 VDDA.n878 VDDA.n877 0.3295
R4311 VDDA.n877 VDDA.n876 0.3295
R4312 VDDA.n876 VDDA.n875 0.3295
R4313 VDDA.n875 VDDA.n874 0.3295
R4314 VDDA.n883 VDDA.n882 0.3295
R4315 VDDA.n884 VDDA.n883 0.3295
R4316 VDDA.n885 VDDA.n884 0.3295
R4317 VDDA.n886 VDDA.n885 0.3295
R4318 VDDA.n887 VDDA.n886 0.3295
R4319 VDDA.n888 VDDA.n887 0.3295
R4320 VDDA.n896 VDDA.n888 0.3295
R4321 VDDA.n896 VDDA.n895 0.3295
R4322 VDDA.n895 VDDA.n894 0.3295
R4323 VDDA.n894 VDDA.n893 0.3295
R4324 VDDA.n893 VDDA.n892 0.3295
R4325 VDDA.n892 VDDA.n891 0.3295
R4326 VDDA.n891 VDDA.n890 0.3295
R4327 VDDA.n890 VDDA.n889 0.3295
R4328 VDDA.n898 VDDA.n897 0.3295
R4329 VDDA.n899 VDDA.n898 0.3295
R4330 VDDA.n900 VDDA.n899 0.3295
R4331 VDDA.n901 VDDA.n900 0.3295
R4332 VDDA.n902 VDDA.n901 0.3295
R4333 VDDA.n903 VDDA.n902 0.3295
R4334 VDDA.n911 VDDA.n903 0.3295
R4335 VDDA.n911 VDDA.n910 0.3295
R4336 VDDA.n910 VDDA.n909 0.3295
R4337 VDDA.n909 VDDA.n908 0.3295
R4338 VDDA.n908 VDDA.n907 0.3295
R4339 VDDA.n907 VDDA.n906 0.3295
R4340 VDDA.n906 VDDA.n905 0.3295
R4341 VDDA.n905 VDDA.n904 0.3295
R4342 VDDA.n913 VDDA.n912 0.3295
R4343 VDDA.n914 VDDA.n913 0.3295
R4344 VDDA.n915 VDDA.n914 0.3295
R4345 VDDA.n916 VDDA.n915 0.3295
R4346 VDDA.n917 VDDA.n916 0.3295
R4347 VDDA.n918 VDDA.n917 0.3295
R4348 VDDA.n926 VDDA.n918 0.3295
R4349 VDDA.n926 VDDA.n925 0.3295
R4350 VDDA.n925 VDDA.n924 0.3295
R4351 VDDA.n924 VDDA.n923 0.3295
R4352 VDDA.n923 VDDA.n922 0.3295
R4353 VDDA.n922 VDDA.n921 0.3295
R4354 VDDA.n921 VDDA.n920 0.3295
R4355 VDDA.n920 VDDA.n919 0.3295
R4356 VDDA.n928 VDDA.n927 0.3295
R4357 VDDA.n929 VDDA.n928 0.3295
R4358 VDDA.n930 VDDA.n929 0.3295
R4359 VDDA.n931 VDDA.n930 0.3295
R4360 VDDA.n932 VDDA.n931 0.3295
R4361 VDDA.n933 VDDA.n932 0.3295
R4362 VDDA.n941 VDDA.n933 0.3295
R4363 VDDA.n941 VDDA.n940 0.3295
R4364 VDDA.n940 VDDA.n939 0.3295
R4365 VDDA.n939 VDDA.n938 0.3295
R4366 VDDA.n938 VDDA.n937 0.3295
R4367 VDDA.n937 VDDA.n936 0.3295
R4368 VDDA.n936 VDDA.n935 0.3295
R4369 VDDA.n935 VDDA.n934 0.3295
R4370 VDDA.n943 VDDA.n942 0.3295
R4371 VDDA.n944 VDDA.n943 0.3295
R4372 VDDA.n945 VDDA.n944 0.3295
R4373 VDDA.n946 VDDA.n945 0.3295
R4374 VDDA.n947 VDDA.n946 0.3295
R4375 VDDA.n948 VDDA.n947 0.3295
R4376 VDDA.n956 VDDA.n948 0.3295
R4377 VDDA.n956 VDDA.n955 0.3295
R4378 VDDA.n955 VDDA.n954 0.3295
R4379 VDDA.n954 VDDA.n953 0.3295
R4380 VDDA.n953 VDDA.n952 0.3295
R4381 VDDA.n952 VDDA.n951 0.3295
R4382 VDDA.n951 VDDA.n950 0.3295
R4383 VDDA.n950 VDDA.n949 0.3295
R4384 VDDA.n958 VDDA.n957 0.3295
R4385 VDDA.n959 VDDA.n958 0.3295
R4386 VDDA.n960 VDDA.n959 0.3295
R4387 VDDA.n961 VDDA.n960 0.3295
R4388 VDDA.n962 VDDA.n961 0.3295
R4389 VDDA.n963 VDDA.n962 0.3295
R4390 VDDA.n971 VDDA.n963 0.3295
R4391 VDDA.n971 VDDA.n970 0.3295
R4392 VDDA.n970 VDDA.n969 0.3295
R4393 VDDA.n969 VDDA.n968 0.3295
R4394 VDDA.n968 VDDA.n967 0.3295
R4395 VDDA.n967 VDDA.n966 0.3295
R4396 VDDA.n966 VDDA.n965 0.3295
R4397 VDDA.n965 VDDA.n964 0.3295
R4398 VDDA.n973 VDDA.n972 0.3295
R4399 VDDA.n974 VDDA.n973 0.3295
R4400 VDDA.n975 VDDA.n974 0.3295
R4401 VDDA.n976 VDDA.n975 0.3295
R4402 VDDA.n977 VDDA.n976 0.3295
R4403 VDDA.n978 VDDA.n977 0.3295
R4404 VDDA.n986 VDDA.n978 0.3295
R4405 VDDA.n986 VDDA.n985 0.3295
R4406 VDDA.n985 VDDA.n984 0.3295
R4407 VDDA.n984 VDDA.n983 0.3295
R4408 VDDA.n983 VDDA.n982 0.3295
R4409 VDDA.n982 VDDA.n981 0.3295
R4410 VDDA.n981 VDDA.n980 0.3295
R4411 VDDA.n980 VDDA.n979 0.3295
R4412 VDDA.n988 VDDA.n987 0.3295
R4413 VDDA.n989 VDDA.n988 0.3295
R4414 VDDA.n990 VDDA.n989 0.3295
R4415 VDDA.n991 VDDA.n990 0.3295
R4416 VDDA.n992 VDDA.n991 0.3295
R4417 VDDA.n993 VDDA.n992 0.3295
R4418 VDDA.n1001 VDDA.n993 0.3295
R4419 VDDA.n1001 VDDA.n1000 0.3295
R4420 VDDA.n1000 VDDA.n999 0.3295
R4421 VDDA.n999 VDDA.n998 0.3295
R4422 VDDA.n998 VDDA.n997 0.3295
R4423 VDDA.n997 VDDA.n996 0.3295
R4424 VDDA.n996 VDDA.n995 0.3295
R4425 VDDA.n995 VDDA.n994 0.3295
R4426 VDDA.n1003 VDDA.n1002 0.3295
R4427 VDDA.n1004 VDDA.n1003 0.3295
R4428 VDDA.n1005 VDDA.n1004 0.3295
R4429 VDDA.n1006 VDDA.n1005 0.3295
R4430 VDDA.n1007 VDDA.n1006 0.3295
R4431 VDDA.n1008 VDDA.n1007 0.3295
R4432 VDDA.n1016 VDDA.n1008 0.3295
R4433 VDDA.n1016 VDDA.n1015 0.3295
R4434 VDDA.n1015 VDDA.n1014 0.3295
R4435 VDDA.n1014 VDDA.n1013 0.3295
R4436 VDDA.n1013 VDDA.n1012 0.3295
R4437 VDDA.n1012 VDDA.n1011 0.3295
R4438 VDDA.n1011 VDDA.n1010 0.3295
R4439 VDDA.n1010 VDDA.n1009 0.3295
R4440 VDDA.n1018 VDDA.n1017 0.3295
R4441 VDDA.n1019 VDDA.n1018 0.3295
R4442 VDDA.n1020 VDDA.n1019 0.3295
R4443 VDDA.n1021 VDDA.n1020 0.3295
R4444 VDDA.n1022 VDDA.n1021 0.3295
R4445 VDDA.n1023 VDDA.n1022 0.3295
R4446 VDDA.n1031 VDDA.n1023 0.3295
R4447 VDDA.n1031 VDDA.n1030 0.3295
R4448 VDDA.n1030 VDDA.n1029 0.3295
R4449 VDDA.n1029 VDDA.n1028 0.3295
R4450 VDDA.n1028 VDDA.n1027 0.3295
R4451 VDDA.n1027 VDDA.n1026 0.3295
R4452 VDDA.n1026 VDDA.n1025 0.3295
R4453 VDDA.n1025 VDDA.n1024 0.3295
R4454 VDDA.n1033 VDDA.n1032 0.3295
R4455 VDDA.n1034 VDDA.n1033 0.3295
R4456 VDDA.n1035 VDDA.n1034 0.3295
R4457 VDDA.n1036 VDDA.n1035 0.3295
R4458 VDDA.n1037 VDDA.n1036 0.3295
R4459 VDDA.n1038 VDDA.n1037 0.3295
R4460 VDDA.n1046 VDDA.n1038 0.3295
R4461 VDDA.n1046 VDDA.n1045 0.3295
R4462 VDDA.n1045 VDDA.n1044 0.3295
R4463 VDDA.n1044 VDDA.n1043 0.3295
R4464 VDDA.n1043 VDDA.n1042 0.3295
R4465 VDDA.n1042 VDDA.n1041 0.3295
R4466 VDDA.n1041 VDDA.n1040 0.3295
R4467 VDDA.n1040 VDDA.n1039 0.3295
R4468 VDDA.n1048 VDDA.n1047 0.3295
R4469 VDDA.n1049 VDDA.n1048 0.3295
R4470 VDDA.n1050 VDDA.n1049 0.3295
R4471 VDDA.n1051 VDDA.n1050 0.3295
R4472 VDDA.n1052 VDDA.n1051 0.3295
R4473 VDDA.n1053 VDDA.n1052 0.3295
R4474 VDDA.n1061 VDDA.n1053 0.3295
R4475 VDDA.n1061 VDDA.n1060 0.3295
R4476 VDDA.n1060 VDDA.n1059 0.3295
R4477 VDDA.n1059 VDDA.n1058 0.3295
R4478 VDDA.n1058 VDDA.n1057 0.3295
R4479 VDDA.n1057 VDDA.n1056 0.3295
R4480 VDDA.n1056 VDDA.n1055 0.3295
R4481 VDDA.n1055 VDDA.n1054 0.3295
R4482 VDDA.n1063 VDDA.n1062 0.3295
R4483 VDDA.n1064 VDDA.n1063 0.3295
R4484 VDDA.n1065 VDDA.n1064 0.3295
R4485 VDDA.n1066 VDDA.n1065 0.3295
R4486 VDDA.n1067 VDDA.n1066 0.3295
R4487 VDDA.n1068 VDDA.n1067 0.3295
R4488 VDDA.n1076 VDDA.n1068 0.3295
R4489 VDDA.n1076 VDDA.n1075 0.3295
R4490 VDDA.n1075 VDDA.n1074 0.3295
R4491 VDDA.n1074 VDDA.n1073 0.3295
R4492 VDDA.n1073 VDDA.n1072 0.3295
R4493 VDDA.n1072 VDDA.n1071 0.3295
R4494 VDDA.n1071 VDDA.n1070 0.3295
R4495 VDDA.n1070 VDDA.n1069 0.3295
R4496 VDDA.n1078 VDDA.n1077 0.3295
R4497 VDDA.n1079 VDDA.n1078 0.3295
R4498 VDDA.n1080 VDDA.n1079 0.3295
R4499 VDDA.n1081 VDDA.n1080 0.3295
R4500 VDDA.n1082 VDDA.n1081 0.3295
R4501 VDDA.n1083 VDDA.n1082 0.3295
R4502 VDDA.n1091 VDDA.n1083 0.3295
R4503 VDDA.n1091 VDDA.n1090 0.3295
R4504 VDDA.n1090 VDDA.n1089 0.3295
R4505 VDDA.n1089 VDDA.n1088 0.3295
R4506 VDDA.n1088 VDDA.n1087 0.3295
R4507 VDDA.n1087 VDDA.n1086 0.3295
R4508 VDDA.n1086 VDDA.n1085 0.3295
R4509 VDDA.n1085 VDDA.n1084 0.3295
R4510 VDDA.n1093 VDDA.n1092 0.3295
R4511 VDDA.n1094 VDDA.n1093 0.3295
R4512 VDDA.n1095 VDDA.n1094 0.3295
R4513 VDDA.n1096 VDDA.n1095 0.3295
R4514 VDDA.n1097 VDDA.n1096 0.3295
R4515 VDDA.n1098 VDDA.n1097 0.3295
R4516 VDDA.n1106 VDDA.n1098 0.3295
R4517 VDDA.n1106 VDDA.n1105 0.3295
R4518 VDDA.n1105 VDDA.n1104 0.3295
R4519 VDDA.n1104 VDDA.n1103 0.3295
R4520 VDDA.n1103 VDDA.n1102 0.3295
R4521 VDDA.n1102 VDDA.n1101 0.3295
R4522 VDDA.n1101 VDDA.n1100 0.3295
R4523 VDDA.n1100 VDDA.n1099 0.3295
R4524 VDDA.n1108 VDDA.n1107 0.3295
R4525 VDDA.n1109 VDDA.n1108 0.3295
R4526 VDDA.n1110 VDDA.n1109 0.3295
R4527 VDDA.n1111 VDDA.n1110 0.3295
R4528 VDDA.n1112 VDDA.n1111 0.3295
R4529 VDDA.n1113 VDDA.n1112 0.3295
R4530 VDDA.n1121 VDDA.n1113 0.3295
R4531 VDDA.n1121 VDDA.n1120 0.3295
R4532 VDDA.n1120 VDDA.n1119 0.3295
R4533 VDDA.n1119 VDDA.n1118 0.3295
R4534 VDDA.n1118 VDDA.n1117 0.3295
R4535 VDDA.n1117 VDDA.n1116 0.3295
R4536 VDDA.n1116 VDDA.n1115 0.3295
R4537 VDDA.n1115 VDDA.n1114 0.3295
R4538 VDDA.n1123 VDDA.n1122 0.3295
R4539 VDDA.n1124 VDDA.n1123 0.3295
R4540 VDDA.n1125 VDDA.n1124 0.3295
R4541 VDDA.n1126 VDDA.n1125 0.3295
R4542 VDDA.n1127 VDDA.n1126 0.3295
R4543 VDDA.n1128 VDDA.n1127 0.3295
R4544 VDDA.n1136 VDDA.n1128 0.3295
R4545 VDDA.n1136 VDDA.n1135 0.3295
R4546 VDDA.n1135 VDDA.n1134 0.3295
R4547 VDDA.n1134 VDDA.n1133 0.3295
R4548 VDDA.n1133 VDDA.n1132 0.3295
R4549 VDDA.n1132 VDDA.n1131 0.3295
R4550 VDDA.n1131 VDDA.n1130 0.3295
R4551 VDDA.n1130 VDDA.n1129 0.3295
R4552 VDDA.n1138 VDDA.n1137 0.3295
R4553 VDDA.n1139 VDDA.n1138 0.3295
R4554 VDDA.n1140 VDDA.n1139 0.3295
R4555 VDDA.n1141 VDDA.n1140 0.3295
R4556 VDDA.n1142 VDDA.n1141 0.3295
R4557 VDDA.n1143 VDDA.n1142 0.3295
R4558 VDDA.n1151 VDDA.n1143 0.3295
R4559 VDDA.n1151 VDDA.n1150 0.3295
R4560 VDDA.n1150 VDDA.n1149 0.3295
R4561 VDDA.n1149 VDDA.n1148 0.3295
R4562 VDDA.n1148 VDDA.n1147 0.3295
R4563 VDDA.n1147 VDDA.n1146 0.3295
R4564 VDDA.n1146 VDDA.n1145 0.3295
R4565 VDDA.n1145 VDDA.n1144 0.3295
R4566 VDDA.n1153 VDDA.n1152 0.3295
R4567 VDDA.n1154 VDDA.n1153 0.3295
R4568 VDDA.n1155 VDDA.n1154 0.3295
R4569 VDDA.n1156 VDDA.n1155 0.3295
R4570 VDDA.n1157 VDDA.n1156 0.3295
R4571 VDDA.n1158 VDDA.n1157 0.3295
R4572 VDDA.n1159 VDDA.n1158 0.3295
R4573 VDDA.n1160 VDDA.n1159 0.3295
R4574 VDDA.n1161 VDDA.n1160 0.3295
R4575 VDDA.n1162 VDDA.n1161 0.3295
R4576 VDDA.n1163 VDDA.n1162 0.3295
R4577 VDDA.n1164 VDDA.n1163 0.3295
R4578 VDDA.n1165 VDDA.n1164 0.3295
R4579 VDDA.n1166 VDDA.n1165 0.3295
R4580 VDDA.n1167 VDDA.n1166 0.3295
R4581 VDDA.n2217 VDDA.n2216 0.292167
R4582 VDDA.n2213 VDDA.n2212 0.292167
R4583 VDDA.n2206 VDDA.n2205 0.292167
R4584 VDDA.n716 VDDA.n701 0.2825
R4585 VDDA.n731 VDDA.n716 0.2825
R4586 VDDA.n746 VDDA.n731 0.2825
R4587 VDDA.n761 VDDA.n746 0.2825
R4588 VDDA.n776 VDDA.n761 0.2825
R4589 VDDA.n791 VDDA.n776 0.2825
R4590 VDDA.n806 VDDA.n791 0.2825
R4591 VDDA.n821 VDDA.n806 0.2825
R4592 VDDA.n836 VDDA.n821 0.2825
R4593 VDDA.n851 VDDA.n836 0.2825
R4594 VDDA.n866 VDDA.n851 0.2825
R4595 VDDA.n881 VDDA.n866 0.2825
R4596 VDDA.n896 VDDA.n881 0.2825
R4597 VDDA.n911 VDDA.n896 0.2825
R4598 VDDA.n926 VDDA.n911 0.2825
R4599 VDDA.n941 VDDA.n926 0.2825
R4600 VDDA.n956 VDDA.n941 0.2825
R4601 VDDA.n971 VDDA.n956 0.2825
R4602 VDDA.n986 VDDA.n971 0.2825
R4603 VDDA.n1001 VDDA.n986 0.2825
R4604 VDDA.n1016 VDDA.n1001 0.2825
R4605 VDDA.n1031 VDDA.n1016 0.2825
R4606 VDDA.n1046 VDDA.n1031 0.2825
R4607 VDDA.n1061 VDDA.n1046 0.2825
R4608 VDDA.n1076 VDDA.n1061 0.2825
R4609 VDDA.n1091 VDDA.n1076 0.2825
R4610 VDDA.n1106 VDDA.n1091 0.2825
R4611 VDDA.n1121 VDDA.n1106 0.2825
R4612 VDDA.n1136 VDDA.n1121 0.2825
R4613 VDDA.n1151 VDDA.n1136 0.2825
R4614 VDDA.n1159 VDDA.n1151 0.2825
R4615 VDDA.n1979 VDDA.n1964 0.246594
R4616 VDDA.n2007 VDDA.n2006 0.246594
R4617 VDDA.n1327 VDDA.n1167 0.194081
R4618 VDDA.t102 VDDA.t195 0.1603
R4619 VDDA.t167 VDDA.t105 0.1603
R4620 VDDA.t106 VDDA.t66 0.1603
R4621 VDDA.t112 VDDA.t9 0.1603
R4622 VDDA.t190 VDDA.t110 0.1603
R4623 VDDA.n233 VDDA.t118 0.159278
R4624 VDDA.n234 VDDA.t107 0.159278
R4625 VDDA.n235 VDDA.t228 0.159278
R4626 VDDA.n236 VDDA.t214 0.159278
R4627 VDDA.n2224 VDDA.n2223 0.146333
R4628 VDDA.n2225 VDDA.n2224 0.146333
R4629 VDDA.n2225 VDDA.n2174 0.146333
R4630 VDDA.n2235 VDDA.n2172 0.146333
R4631 VDDA.n2243 VDDA.n2172 0.146333
R4632 VDDA.n2244 VDDA.n2243 0.146333
R4633 VDDA.n2254 VDDA.n2253 0.146333
R4634 VDDA.n2255 VDDA.n2254 0.146333
R4635 VDDA.n2255 VDDA.n2168 0.146333
R4636 VDDA.n2265 VDDA.n2166 0.146333
R4637 VDDA.n2273 VDDA.n2166 0.146333
R4638 VDDA.n2274 VDDA.n2273 0.146333
R4639 VDDA.n2284 VDDA.n2283 0.146333
R4640 VDDA.n2285 VDDA.n2284 0.146333
R4641 VDDA.n2285 VDDA.n2162 0.146333
R4642 VDDA.n2295 VDDA.n2160 0.146333
R4643 VDDA.n2303 VDDA.n2160 0.146333
R4644 VDDA.n2304 VDDA.n2303 0.146333
R4645 VDDA.n2314 VDDA.n2313 0.146333
R4646 VDDA.n2315 VDDA.n2314 0.146333
R4647 VDDA.n2315 VDDA.n2156 0.146333
R4648 VDDA.n2325 VDDA.n2154 0.146333
R4649 VDDA.n2333 VDDA.n2154 0.146333
R4650 VDDA.n2222 VDDA.n2175 0.146333
R4651 VDDA.n2228 VDDA.n2175 0.146333
R4652 VDDA.n2229 VDDA.n2228 0.146333
R4653 VDDA.n2239 VDDA.n2238 0.146333
R4654 VDDA.n2242 VDDA.n2239 0.146333
R4655 VDDA.n2242 VDDA.n2171 0.146333
R4656 VDDA.n2252 VDDA.n2169 0.146333
R4657 VDDA.n2258 VDDA.n2169 0.146333
R4658 VDDA.n2259 VDDA.n2258 0.146333
R4659 VDDA.n2269 VDDA.n2268 0.146333
R4660 VDDA.n2272 VDDA.n2269 0.146333
R4661 VDDA.n2272 VDDA.n2165 0.146333
R4662 VDDA.n2282 VDDA.n2163 0.146333
R4663 VDDA.n2288 VDDA.n2163 0.146333
R4664 VDDA.n2289 VDDA.n2288 0.146333
R4665 VDDA.n2299 VDDA.n2298 0.146333
R4666 VDDA.n2302 VDDA.n2299 0.146333
R4667 VDDA.n2302 VDDA.n2159 0.146333
R4668 VDDA.n2312 VDDA.n2157 0.146333
R4669 VDDA.n2318 VDDA.n2157 0.146333
R4670 VDDA.n2319 VDDA.n2318 0.146333
R4671 VDDA.n2329 VDDA.n2328 0.146333
R4672 VDDA.n2332 VDDA.n2329 0.146333
R4673 VDDA.n2332 VDDA.n2153 0.146333
R4674 VDDA.n2039 VDDA.n2038 0.146333
R4675 VDDA.n2040 VDDA.n2039 0.146333
R4676 VDDA.n2040 VDDA.n1945 0.146333
R4677 VDDA.n2050 VDDA.n1943 0.146333
R4678 VDDA.n2058 VDDA.n1943 0.146333
R4679 VDDA.n2059 VDDA.n2058 0.146333
R4680 VDDA.n2069 VDDA.n2068 0.146333
R4681 VDDA.n2070 VDDA.n2069 0.146333
R4682 VDDA.n2070 VDDA.n1939 0.146333
R4683 VDDA.n2080 VDDA.n1937 0.146333
R4684 VDDA.n2088 VDDA.n1937 0.146333
R4685 VDDA.n2089 VDDA.n2088 0.146333
R4686 VDDA.n2099 VDDA.n2098 0.146333
R4687 VDDA.n2100 VDDA.n2099 0.146333
R4688 VDDA.n2100 VDDA.n1933 0.146333
R4689 VDDA.n2110 VDDA.n1931 0.146333
R4690 VDDA.n2118 VDDA.n1931 0.146333
R4691 VDDA.n2119 VDDA.n2118 0.146333
R4692 VDDA.n2129 VDDA.n2128 0.146333
R4693 VDDA.n2130 VDDA.n2129 0.146333
R4694 VDDA.n2130 VDDA.n1927 0.146333
R4695 VDDA.n2140 VDDA.n1925 0.146333
R4696 VDDA.n2148 VDDA.n1925 0.146333
R4697 VDDA.n2037 VDDA.n1946 0.146333
R4698 VDDA.n2043 VDDA.n1946 0.146333
R4699 VDDA.n2044 VDDA.n2043 0.146333
R4700 VDDA.n2054 VDDA.n2053 0.146333
R4701 VDDA.n2057 VDDA.n2054 0.146333
R4702 VDDA.n2057 VDDA.n1942 0.146333
R4703 VDDA.n2067 VDDA.n1940 0.146333
R4704 VDDA.n2073 VDDA.n1940 0.146333
R4705 VDDA.n2074 VDDA.n2073 0.146333
R4706 VDDA.n2084 VDDA.n2083 0.146333
R4707 VDDA.n2087 VDDA.n2084 0.146333
R4708 VDDA.n2087 VDDA.n1936 0.146333
R4709 VDDA.n2097 VDDA.n1934 0.146333
R4710 VDDA.n2103 VDDA.n1934 0.146333
R4711 VDDA.n2104 VDDA.n2103 0.146333
R4712 VDDA.n2114 VDDA.n2113 0.146333
R4713 VDDA.n2117 VDDA.n2114 0.146333
R4714 VDDA.n2117 VDDA.n1930 0.146333
R4715 VDDA.n2127 VDDA.n1928 0.146333
R4716 VDDA.n2133 VDDA.n1928 0.146333
R4717 VDDA.n2134 VDDA.n2133 0.146333
R4718 VDDA.n2144 VDDA.n2143 0.146333
R4719 VDDA.n2147 VDDA.n2144 0.146333
R4720 VDDA.n2147 VDDA.n1924 0.146333
R4721 VDDA.n242 VDDA.n241 0.146333
R4722 VDDA.n243 VDDA.n242 0.146333
R4723 VDDA.n243 VDDA.n230 0.146333
R4724 VDDA.n253 VDDA.n228 0.146333
R4725 VDDA.n261 VDDA.n228 0.146333
R4726 VDDA.n262 VDDA.n261 0.146333
R4727 VDDA.n272 VDDA.n271 0.146333
R4728 VDDA.n273 VDDA.n272 0.146333
R4729 VDDA.n273 VDDA.n224 0.146333
R4730 VDDA.n283 VDDA.n222 0.146333
R4731 VDDA.n291 VDDA.n222 0.146333
R4732 VDDA.n292 VDDA.n291 0.146333
R4733 VDDA.n302 VDDA.n301 0.146333
R4734 VDDA.n303 VDDA.n302 0.146333
R4735 VDDA.n303 VDDA.n218 0.146333
R4736 VDDA.n313 VDDA.n216 0.146333
R4737 VDDA.n321 VDDA.n216 0.146333
R4738 VDDA.n322 VDDA.n321 0.146333
R4739 VDDA.n332 VDDA.n331 0.146333
R4740 VDDA.n333 VDDA.n332 0.146333
R4741 VDDA.n333 VDDA.n212 0.146333
R4742 VDDA.n343 VDDA.n210 0.146333
R4743 VDDA.n351 VDDA.n210 0.146333
R4744 VDDA.n240 VDDA.n231 0.146333
R4745 VDDA.n246 VDDA.n231 0.146333
R4746 VDDA.n247 VDDA.n246 0.146333
R4747 VDDA.n257 VDDA.n256 0.146333
R4748 VDDA.n260 VDDA.n257 0.146333
R4749 VDDA.n260 VDDA.n227 0.146333
R4750 VDDA.n270 VDDA.n225 0.146333
R4751 VDDA.n276 VDDA.n225 0.146333
R4752 VDDA.n277 VDDA.n276 0.146333
R4753 VDDA.n287 VDDA.n286 0.146333
R4754 VDDA.n290 VDDA.n287 0.146333
R4755 VDDA.n290 VDDA.n221 0.146333
R4756 VDDA.n300 VDDA.n219 0.146333
R4757 VDDA.n306 VDDA.n219 0.146333
R4758 VDDA.n307 VDDA.n306 0.146333
R4759 VDDA.n317 VDDA.n316 0.146333
R4760 VDDA.n320 VDDA.n317 0.146333
R4761 VDDA.n320 VDDA.n215 0.146333
R4762 VDDA.n330 VDDA.n213 0.146333
R4763 VDDA.n336 VDDA.n213 0.146333
R4764 VDDA.n337 VDDA.n336 0.146333
R4765 VDDA.n347 VDDA.n346 0.146333
R4766 VDDA.n350 VDDA.n347 0.146333
R4767 VDDA.n350 VDDA.n209 0.146333
R4768 VDDA.n2565 VDDA.n2564 0.146333
R4769 VDDA.n2566 VDDA.n2565 0.146333
R4770 VDDA.n2566 VDDA.n2555 0.146333
R4771 VDDA.n2576 VDDA.n2553 0.146333
R4772 VDDA.n2584 VDDA.n2553 0.146333
R4773 VDDA.n2585 VDDA.n2584 0.146333
R4774 VDDA.n2595 VDDA.n2594 0.146333
R4775 VDDA.n2596 VDDA.n2595 0.146333
R4776 VDDA.n2596 VDDA.n2549 0.146333
R4777 VDDA.n2606 VDDA.n2547 0.146333
R4778 VDDA.n2614 VDDA.n2547 0.146333
R4779 VDDA.n2615 VDDA.n2614 0.146333
R4780 VDDA.n2625 VDDA.n2624 0.146333
R4781 VDDA.n2626 VDDA.n2625 0.146333
R4782 VDDA.n2626 VDDA.n2543 0.146333
R4783 VDDA.n2636 VDDA.n2541 0.146333
R4784 VDDA.n2644 VDDA.n2541 0.146333
R4785 VDDA.n2645 VDDA.n2644 0.146333
R4786 VDDA.n2655 VDDA.n2654 0.146333
R4787 VDDA.n2656 VDDA.n2655 0.146333
R4788 VDDA.n2656 VDDA.n2537 0.146333
R4789 VDDA.n2666 VDDA.n2535 0.146333
R4790 VDDA.n2674 VDDA.n2535 0.146333
R4791 VDDA.n2563 VDDA.n2556 0.146333
R4792 VDDA.n2569 VDDA.n2556 0.146333
R4793 VDDA.n2570 VDDA.n2569 0.146333
R4794 VDDA.n2580 VDDA.n2579 0.146333
R4795 VDDA.n2583 VDDA.n2580 0.146333
R4796 VDDA.n2583 VDDA.n2552 0.146333
R4797 VDDA.n2593 VDDA.n2550 0.146333
R4798 VDDA.n2599 VDDA.n2550 0.146333
R4799 VDDA.n2600 VDDA.n2599 0.146333
R4800 VDDA.n2610 VDDA.n2609 0.146333
R4801 VDDA.n2613 VDDA.n2610 0.146333
R4802 VDDA.n2613 VDDA.n2546 0.146333
R4803 VDDA.n2623 VDDA.n2544 0.146333
R4804 VDDA.n2629 VDDA.n2544 0.146333
R4805 VDDA.n2630 VDDA.n2629 0.146333
R4806 VDDA.n2640 VDDA.n2639 0.146333
R4807 VDDA.n2643 VDDA.n2640 0.146333
R4808 VDDA.n2643 VDDA.n2540 0.146333
R4809 VDDA.n2653 VDDA.n2538 0.146333
R4810 VDDA.n2659 VDDA.n2538 0.146333
R4811 VDDA.n2660 VDDA.n2659 0.146333
R4812 VDDA.n2670 VDDA.n2669 0.146333
R4813 VDDA.n2673 VDDA.n2670 0.146333
R4814 VDDA.n2673 VDDA.n2534 0.146333
R4815 VDDA.n2420 VDDA.n2419 0.146333
R4816 VDDA.n2421 VDDA.n2420 0.146333
R4817 VDDA.n2421 VDDA.n2359 0.146333
R4818 VDDA.n2431 VDDA.n2357 0.146333
R4819 VDDA.n2439 VDDA.n2357 0.146333
R4820 VDDA.n2440 VDDA.n2439 0.146333
R4821 VDDA.n2450 VDDA.n2449 0.146333
R4822 VDDA.n2451 VDDA.n2450 0.146333
R4823 VDDA.n2451 VDDA.n2353 0.146333
R4824 VDDA.n2461 VDDA.n2351 0.146333
R4825 VDDA.n2469 VDDA.n2351 0.146333
R4826 VDDA.n2470 VDDA.n2469 0.146333
R4827 VDDA.n2480 VDDA.n2479 0.146333
R4828 VDDA.n2481 VDDA.n2480 0.146333
R4829 VDDA.n2481 VDDA.n2347 0.146333
R4830 VDDA.n2491 VDDA.n2345 0.146333
R4831 VDDA.n2499 VDDA.n2345 0.146333
R4832 VDDA.n2500 VDDA.n2499 0.146333
R4833 VDDA.n2510 VDDA.n2509 0.146333
R4834 VDDA.n2511 VDDA.n2510 0.146333
R4835 VDDA.n2511 VDDA.n2341 0.146333
R4836 VDDA.n2521 VDDA.n2339 0.146333
R4837 VDDA.n2529 VDDA.n2339 0.146333
R4838 VDDA.n2418 VDDA.n2360 0.146333
R4839 VDDA.n2424 VDDA.n2360 0.146333
R4840 VDDA.n2425 VDDA.n2424 0.146333
R4841 VDDA.n2435 VDDA.n2434 0.146333
R4842 VDDA.n2438 VDDA.n2435 0.146333
R4843 VDDA.n2438 VDDA.n2356 0.146333
R4844 VDDA.n2448 VDDA.n2354 0.146333
R4845 VDDA.n2454 VDDA.n2354 0.146333
R4846 VDDA.n2455 VDDA.n2454 0.146333
R4847 VDDA.n2465 VDDA.n2464 0.146333
R4848 VDDA.n2468 VDDA.n2465 0.146333
R4849 VDDA.n2468 VDDA.n2350 0.146333
R4850 VDDA.n2478 VDDA.n2348 0.146333
R4851 VDDA.n2484 VDDA.n2348 0.146333
R4852 VDDA.n2485 VDDA.n2484 0.146333
R4853 VDDA.n2495 VDDA.n2494 0.146333
R4854 VDDA.n2498 VDDA.n2495 0.146333
R4855 VDDA.n2498 VDDA.n2344 0.146333
R4856 VDDA.n2508 VDDA.n2342 0.146333
R4857 VDDA.n2514 VDDA.n2342 0.146333
R4858 VDDA.n2515 VDDA.n2514 0.146333
R4859 VDDA.n2525 VDDA.n2524 0.146333
R4860 VDDA.n2528 VDDA.n2525 0.146333
R4861 VDDA.n2528 VDDA.n2338 0.146333
R4862 VDDA.n89 VDDA.n85 0.146333
R4863 VDDA.n93 VDDA.n85 0.146333
R4864 VDDA.n94 VDDA.n93 0.146333
R4865 VDDA.n102 VDDA.n101 0.146333
R4866 VDDA.n105 VDDA.n102 0.146333
R4867 VDDA.n105 VDDA.n77 0.146333
R4868 VDDA.n113 VDDA.n73 0.146333
R4869 VDDA.n117 VDDA.n73 0.146333
R4870 VDDA.n118 VDDA.n117 0.146333
R4871 VDDA.n126 VDDA.n125 0.146333
R4872 VDDA.n129 VDDA.n126 0.146333
R4873 VDDA.n129 VDDA.n65 0.146333
R4874 VDDA.n137 VDDA.n61 0.146333
R4875 VDDA.n141 VDDA.n61 0.146333
R4876 VDDA.n142 VDDA.n141 0.146333
R4877 VDDA.n150 VDDA.n149 0.146333
R4878 VDDA.n153 VDDA.n150 0.146333
R4879 VDDA.n153 VDDA.n53 0.146333
R4880 VDDA.n161 VDDA.n49 0.146333
R4881 VDDA.n165 VDDA.n49 0.146333
R4882 VDDA.n166 VDDA.n165 0.146333
R4883 VDDA.n174 VDDA.n173 0.146333
R4884 VDDA.n177 VDDA.n174 0.146333
R4885 VDDA.n177 VDDA.n43 0.146333
R4886 VDDA.n3239 VDDA.n3236 0.146333
R4887 VDDA.n3245 VDDA.n3236 0.146333
R4888 VDDA.n3245 VDDA.n3234 0.146333
R4889 VDDA.n3255 VDDA.n3230 0.146333
R4890 VDDA.n3259 VDDA.n3230 0.146333
R4891 VDDA.n3259 VDDA.n3228 0.146333
R4892 VDDA.n3269 VDDA.n3224 0.146333
R4893 VDDA.n3275 VDDA.n3224 0.146333
R4894 VDDA.n3275 VDDA.n3222 0.146333
R4895 VDDA.n3285 VDDA.n3218 0.146333
R4896 VDDA.n3289 VDDA.n3218 0.146333
R4897 VDDA.n3289 VDDA.n3216 0.146333
R4898 VDDA.n3299 VDDA.n3212 0.146333
R4899 VDDA.n3305 VDDA.n3212 0.146333
R4900 VDDA.n3305 VDDA.n3210 0.146333
R4901 VDDA.n3315 VDDA.n3206 0.146333
R4902 VDDA.n3319 VDDA.n3206 0.146333
R4903 VDDA.n3319 VDDA.n3204 0.146333
R4904 VDDA.n3329 VDDA.n3200 0.146333
R4905 VDDA.n3335 VDDA.n3200 0.146333
R4906 VDDA.n3335 VDDA.n3198 0.146333
R4907 VDDA.n3345 VDDA.n3194 0.146333
R4908 VDDA.n3349 VDDA.n3194 0.146333
R4909 VDDA.n3349 VDDA.n3192 0.146333
R4910 VDDA.n3096 VDDA.n3095 0.146333
R4911 VDDA.n3099 VDDA.n3096 0.146333
R4912 VDDA.n3099 VDDA.n3089 0.146333
R4913 VDDA.n3107 VDDA.n3085 0.146333
R4914 VDDA.n3111 VDDA.n3085 0.146333
R4915 VDDA.n3112 VDDA.n3111 0.146333
R4916 VDDA.n3120 VDDA.n3119 0.146333
R4917 VDDA.n3123 VDDA.n3120 0.146333
R4918 VDDA.n3123 VDDA.n3077 0.146333
R4919 VDDA.n3131 VDDA.n3073 0.146333
R4920 VDDA.n3135 VDDA.n3073 0.146333
R4921 VDDA.n3136 VDDA.n3135 0.146333
R4922 VDDA.n3144 VDDA.n3143 0.146333
R4923 VDDA.n3147 VDDA.n3144 0.146333
R4924 VDDA.n3147 VDDA.n3065 0.146333
R4925 VDDA.n3155 VDDA.n3061 0.146333
R4926 VDDA.n3159 VDDA.n3061 0.146333
R4927 VDDA.n3160 VDDA.n3159 0.146333
R4928 VDDA.n3168 VDDA.n3167 0.146333
R4929 VDDA.n3171 VDDA.n3168 0.146333
R4930 VDDA.n3171 VDDA.n3053 0.146333
R4931 VDDA.n3179 VDDA.n3051 0.146333
R4932 VDDA.n3183 VDDA.n3051 0.146333
R4933 VDDA.n3183 VDDA.n182 0.146333
R4934 VDDA.n2932 VDDA.n2928 0.146333
R4935 VDDA.n2936 VDDA.n2928 0.146333
R4936 VDDA.n2937 VDDA.n2936 0.146333
R4937 VDDA.n2945 VDDA.n2944 0.146333
R4938 VDDA.n2948 VDDA.n2945 0.146333
R4939 VDDA.n2948 VDDA.n2920 0.146333
R4940 VDDA.n2956 VDDA.n2916 0.146333
R4941 VDDA.n2960 VDDA.n2916 0.146333
R4942 VDDA.n2961 VDDA.n2960 0.146333
R4943 VDDA.n2969 VDDA.n2968 0.146333
R4944 VDDA.n2972 VDDA.n2969 0.146333
R4945 VDDA.n2972 VDDA.n2908 0.146333
R4946 VDDA.n2980 VDDA.n2904 0.146333
R4947 VDDA.n2984 VDDA.n2904 0.146333
R4948 VDDA.n2985 VDDA.n2984 0.146333
R4949 VDDA.n2993 VDDA.n2992 0.146333
R4950 VDDA.n2996 VDDA.n2993 0.146333
R4951 VDDA.n2996 VDDA.n2896 0.146333
R4952 VDDA.n3004 VDDA.n2892 0.146333
R4953 VDDA.n3008 VDDA.n2892 0.146333
R4954 VDDA.n3009 VDDA.n3008 0.146333
R4955 VDDA.n3017 VDDA.n3016 0.146333
R4956 VDDA.n3020 VDDA.n3017 0.146333
R4957 VDDA.n3020 VDDA.n2886 0.146333
R4958 VDDA.n426 VDDA.n422 0.146333
R4959 VDDA.n430 VDDA.n422 0.146333
R4960 VDDA.n431 VDDA.n430 0.146333
R4961 VDDA.n439 VDDA.n438 0.146333
R4962 VDDA.n442 VDDA.n439 0.146333
R4963 VDDA.n442 VDDA.n414 0.146333
R4964 VDDA.n450 VDDA.n410 0.146333
R4965 VDDA.n454 VDDA.n410 0.146333
R4966 VDDA.n455 VDDA.n454 0.146333
R4967 VDDA.n463 VDDA.n462 0.146333
R4968 VDDA.n466 VDDA.n463 0.146333
R4969 VDDA.n466 VDDA.n402 0.146333
R4970 VDDA.n474 VDDA.n398 0.146333
R4971 VDDA.n478 VDDA.n398 0.146333
R4972 VDDA.n479 VDDA.n478 0.146333
R4973 VDDA.n487 VDDA.n486 0.146333
R4974 VDDA.n490 VDDA.n487 0.146333
R4975 VDDA.n490 VDDA.n390 0.146333
R4976 VDDA.n498 VDDA.n386 0.146333
R4977 VDDA.n502 VDDA.n386 0.146333
R4978 VDDA.n503 VDDA.n502 0.146333
R4979 VDDA.n511 VDDA.n510 0.146333
R4980 VDDA.n514 VDDA.n511 0.146333
R4981 VDDA.n514 VDDA.n380 0.146333
R4982 VDDA.n1737 VDDA.n1736 0.146333
R4983 VDDA.n1740 VDDA.n1737 0.146333
R4984 VDDA.n1740 VDDA.n1730 0.146333
R4985 VDDA.n1748 VDDA.n1726 0.146333
R4986 VDDA.n1752 VDDA.n1726 0.146333
R4987 VDDA.n1753 VDDA.n1752 0.146333
R4988 VDDA.n1761 VDDA.n1760 0.146333
R4989 VDDA.n1764 VDDA.n1761 0.146333
R4990 VDDA.n1764 VDDA.n1718 0.146333
R4991 VDDA.n1772 VDDA.n1714 0.146333
R4992 VDDA.n1776 VDDA.n1714 0.146333
R4993 VDDA.n1777 VDDA.n1776 0.146333
R4994 VDDA.n1785 VDDA.n1784 0.146333
R4995 VDDA.n1788 VDDA.n1785 0.146333
R4996 VDDA.n1788 VDDA.n1706 0.146333
R4997 VDDA.n1796 VDDA.n1702 0.146333
R4998 VDDA.n1800 VDDA.n1702 0.146333
R4999 VDDA.n1801 VDDA.n1800 0.146333
R5000 VDDA.n1809 VDDA.n1808 0.146333
R5001 VDDA.n1812 VDDA.n1809 0.146333
R5002 VDDA.n1812 VDDA.n1694 0.146333
R5003 VDDA.n1820 VDDA.n1692 0.146333
R5004 VDDA.n1824 VDDA.n1692 0.146333
R5005 VDDA.n1824 VDDA.n519 0.146333
R5006 VDDA.n1573 VDDA.n1569 0.146333
R5007 VDDA.n1577 VDDA.n1569 0.146333
R5008 VDDA.n1578 VDDA.n1577 0.146333
R5009 VDDA.n1586 VDDA.n1585 0.146333
R5010 VDDA.n1589 VDDA.n1586 0.146333
R5011 VDDA.n1589 VDDA.n1561 0.146333
R5012 VDDA.n1597 VDDA.n1557 0.146333
R5013 VDDA.n1601 VDDA.n1557 0.146333
R5014 VDDA.n1602 VDDA.n1601 0.146333
R5015 VDDA.n1610 VDDA.n1609 0.146333
R5016 VDDA.n1613 VDDA.n1610 0.146333
R5017 VDDA.n1613 VDDA.n1549 0.146333
R5018 VDDA.n1621 VDDA.n1545 0.146333
R5019 VDDA.n1625 VDDA.n1545 0.146333
R5020 VDDA.n1626 VDDA.n1625 0.146333
R5021 VDDA.n1634 VDDA.n1633 0.146333
R5022 VDDA.n1637 VDDA.n1634 0.146333
R5023 VDDA.n1637 VDDA.n1537 0.146333
R5024 VDDA.n1645 VDDA.n1533 0.146333
R5025 VDDA.n1649 VDDA.n1533 0.146333
R5026 VDDA.n1650 VDDA.n1649 0.146333
R5027 VDDA.n1658 VDDA.n1657 0.146333
R5028 VDDA.n1661 VDDA.n1658 0.146333
R5029 VDDA.n1661 VDDA.n1527 0.146333
R5030 VDDA.n593 VDDA.n589 0.146333
R5031 VDDA.n597 VDDA.n589 0.146333
R5032 VDDA.n598 VDDA.n597 0.146333
R5033 VDDA.n606 VDDA.n605 0.146333
R5034 VDDA.n609 VDDA.n606 0.146333
R5035 VDDA.n609 VDDA.n581 0.146333
R5036 VDDA.n617 VDDA.n577 0.146333
R5037 VDDA.n621 VDDA.n577 0.146333
R5038 VDDA.n622 VDDA.n621 0.146333
R5039 VDDA.n630 VDDA.n629 0.146333
R5040 VDDA.n633 VDDA.n630 0.146333
R5041 VDDA.n633 VDDA.n569 0.146333
R5042 VDDA.n641 VDDA.n565 0.146333
R5043 VDDA.n645 VDDA.n565 0.146333
R5044 VDDA.n646 VDDA.n645 0.146333
R5045 VDDA.n654 VDDA.n653 0.146333
R5046 VDDA.n657 VDDA.n654 0.146333
R5047 VDDA.n657 VDDA.n557 0.146333
R5048 VDDA.n665 VDDA.n553 0.146333
R5049 VDDA.n669 VDDA.n553 0.146333
R5050 VDDA.n670 VDDA.n669 0.146333
R5051 VDDA.n678 VDDA.n677 0.146333
R5052 VDDA.n681 VDDA.n678 0.146333
R5053 VDDA.n681 VDDA.n547 0.146333
R5054 VDDA.n1379 VDDA.n1376 0.146333
R5055 VDDA.n1385 VDDA.n1376 0.146333
R5056 VDDA.n1385 VDDA.n1374 0.146333
R5057 VDDA.n1395 VDDA.n1370 0.146333
R5058 VDDA.n1399 VDDA.n1370 0.146333
R5059 VDDA.n1399 VDDA.n1368 0.146333
R5060 VDDA.n1409 VDDA.n1364 0.146333
R5061 VDDA.n1415 VDDA.n1364 0.146333
R5062 VDDA.n1415 VDDA.n1362 0.146333
R5063 VDDA.n1425 VDDA.n1358 0.146333
R5064 VDDA.n1429 VDDA.n1358 0.146333
R5065 VDDA.n1429 VDDA.n1356 0.146333
R5066 VDDA.n1439 VDDA.n1352 0.146333
R5067 VDDA.n1445 VDDA.n1352 0.146333
R5068 VDDA.n1445 VDDA.n1350 0.146333
R5069 VDDA.n1455 VDDA.n1346 0.146333
R5070 VDDA.n1459 VDDA.n1346 0.146333
R5071 VDDA.n1459 VDDA.n1344 0.146333
R5072 VDDA.n1469 VDDA.n1340 0.146333
R5073 VDDA.n1475 VDDA.n1340 0.146333
R5074 VDDA.n1475 VDDA.n1338 0.146333
R5075 VDDA.n1485 VDDA.n1334 0.146333
R5076 VDDA.n1489 VDDA.n1334 0.146333
R5077 VDDA.n1489 VDDA.n1332 0.146333
R5078 VDDA.n1217 VDDA.n1216 0.146333
R5079 VDDA.n1220 VDDA.n1217 0.146333
R5080 VDDA.n1220 VDDA.n1212 0.146333
R5081 VDDA.n1230 VDDA.n1210 0.146333
R5082 VDDA.n1236 VDDA.n1210 0.146333
R5083 VDDA.n1237 VDDA.n1236 0.146333
R5084 VDDA.n1247 VDDA.n1246 0.146333
R5085 VDDA.n1250 VDDA.n1247 0.146333
R5086 VDDA.n1250 VDDA.n1206 0.146333
R5087 VDDA.n1260 VDDA.n1204 0.146333
R5088 VDDA.n1266 VDDA.n1204 0.146333
R5089 VDDA.n1267 VDDA.n1266 0.146333
R5090 VDDA.n1277 VDDA.n1276 0.146333
R5091 VDDA.n1280 VDDA.n1277 0.146333
R5092 VDDA.n1280 VDDA.n1200 0.146333
R5093 VDDA.n1290 VDDA.n1198 0.146333
R5094 VDDA.n1296 VDDA.n1198 0.146333
R5095 VDDA.n1297 VDDA.n1296 0.146333
R5096 VDDA.n1307 VDDA.n1306 0.146333
R5097 VDDA.n1310 VDDA.n1307 0.146333
R5098 VDDA.n1310 VDDA.n1194 0.146333
R5099 VDDA.n1320 VDDA.n1192 0.146333
R5100 VDDA.n1324 VDDA.n1192 0.146333
R5101 VDDA.n1324 VDDA.n685 0.146333
R5102 VDDA.n1979 VDDA.n1978 0.141125
R5103 VDDA.n1978 VDDA.n1977 0.141125
R5104 VDDA.n1977 VDDA.n1976 0.141125
R5105 VDDA.n1976 VDDA.n1975 0.141125
R5106 VDDA.n1975 VDDA.n1974 0.141125
R5107 VDDA.n1974 VDDA.n1973 0.141125
R5108 VDDA.n1973 VDDA.n1972 0.141125
R5109 VDDA.n1972 VDDA.n1948 0.141125
R5110 VDDA.n2006 VDDA.n1948 0.141125
R5111 VDDA.n236 VDDA.t185 0.1368
R5112 VDDA.n236 VDDA.t102 0.1368
R5113 VDDA.n235 VDDA.t213 0.1368
R5114 VDDA.n235 VDDA.t167 0.1368
R5115 VDDA.n234 VDDA.t57 0.1368
R5116 VDDA.n234 VDDA.t106 0.1368
R5117 VDDA.n233 VDDA.t229 0.1368
R5118 VDDA.n233 VDDA.t112 0.1368
R5119 VDDA.n232 VDDA.t58 0.1368
R5120 VDDA.n232 VDDA.t190 0.1368
R5121 VDDA.n2223 VDDA.n2219 0.135917
R5122 VDDA.n2233 VDDA.n2174 0.135917
R5123 VDDA.n2235 VDDA.n2234 0.135917
R5124 VDDA.n2245 VDDA.n2244 0.135917
R5125 VDDA.n2253 VDDA.n2170 0.135917
R5126 VDDA.n2263 VDDA.n2168 0.135917
R5127 VDDA.n2265 VDDA.n2264 0.135917
R5128 VDDA.n2275 VDDA.n2274 0.135917
R5129 VDDA.n2283 VDDA.n2164 0.135917
R5130 VDDA.n2293 VDDA.n2162 0.135917
R5131 VDDA.n2295 VDDA.n2294 0.135917
R5132 VDDA.n2305 VDDA.n2304 0.135917
R5133 VDDA.n2313 VDDA.n2158 0.135917
R5134 VDDA.n2323 VDDA.n2156 0.135917
R5135 VDDA.n2325 VDDA.n2324 0.135917
R5136 VDDA.n2222 VDDA.n2220 0.135917
R5137 VDDA.n2232 VDDA.n2229 0.135917
R5138 VDDA.n2238 VDDA.n2173 0.135917
R5139 VDDA.n2248 VDDA.n2171 0.135917
R5140 VDDA.n2252 VDDA.n2249 0.135917
R5141 VDDA.n2262 VDDA.n2259 0.135917
R5142 VDDA.n2268 VDDA.n2167 0.135917
R5143 VDDA.n2278 VDDA.n2165 0.135917
R5144 VDDA.n2282 VDDA.n2279 0.135917
R5145 VDDA.n2292 VDDA.n2289 0.135917
R5146 VDDA.n2298 VDDA.n2161 0.135917
R5147 VDDA.n2308 VDDA.n2159 0.135917
R5148 VDDA.n2312 VDDA.n2309 0.135917
R5149 VDDA.n2322 VDDA.n2319 0.135917
R5150 VDDA.n2328 VDDA.n2155 0.135917
R5151 VDDA.n2038 VDDA.n2034 0.135917
R5152 VDDA.n2048 VDDA.n1945 0.135917
R5153 VDDA.n2050 VDDA.n2049 0.135917
R5154 VDDA.n2060 VDDA.n2059 0.135917
R5155 VDDA.n2068 VDDA.n1941 0.135917
R5156 VDDA.n2078 VDDA.n1939 0.135917
R5157 VDDA.n2080 VDDA.n2079 0.135917
R5158 VDDA.n2090 VDDA.n2089 0.135917
R5159 VDDA.n2098 VDDA.n1935 0.135917
R5160 VDDA.n2108 VDDA.n1933 0.135917
R5161 VDDA.n2110 VDDA.n2109 0.135917
R5162 VDDA.n2120 VDDA.n2119 0.135917
R5163 VDDA.n2128 VDDA.n1929 0.135917
R5164 VDDA.n2138 VDDA.n1927 0.135917
R5165 VDDA.n2140 VDDA.n2139 0.135917
R5166 VDDA.n2037 VDDA.n2035 0.135917
R5167 VDDA.n2047 VDDA.n2044 0.135917
R5168 VDDA.n2053 VDDA.n1944 0.135917
R5169 VDDA.n2063 VDDA.n1942 0.135917
R5170 VDDA.n2067 VDDA.n2064 0.135917
R5171 VDDA.n2077 VDDA.n2074 0.135917
R5172 VDDA.n2083 VDDA.n1938 0.135917
R5173 VDDA.n2093 VDDA.n1936 0.135917
R5174 VDDA.n2097 VDDA.n2094 0.135917
R5175 VDDA.n2107 VDDA.n2104 0.135917
R5176 VDDA.n2113 VDDA.n1932 0.135917
R5177 VDDA.n2123 VDDA.n1930 0.135917
R5178 VDDA.n2127 VDDA.n2124 0.135917
R5179 VDDA.n2137 VDDA.n2134 0.135917
R5180 VDDA.n2143 VDDA.n1926 0.135917
R5181 VDDA.n241 VDDA.n237 0.135917
R5182 VDDA.n251 VDDA.n230 0.135917
R5183 VDDA.n253 VDDA.n252 0.135917
R5184 VDDA.n263 VDDA.n262 0.135917
R5185 VDDA.n271 VDDA.n226 0.135917
R5186 VDDA.n281 VDDA.n224 0.135917
R5187 VDDA.n283 VDDA.n282 0.135917
R5188 VDDA.n293 VDDA.n292 0.135917
R5189 VDDA.n301 VDDA.n220 0.135917
R5190 VDDA.n311 VDDA.n218 0.135917
R5191 VDDA.n313 VDDA.n312 0.135917
R5192 VDDA.n323 VDDA.n322 0.135917
R5193 VDDA.n331 VDDA.n214 0.135917
R5194 VDDA.n341 VDDA.n212 0.135917
R5195 VDDA.n343 VDDA.n342 0.135917
R5196 VDDA.n240 VDDA.n238 0.135917
R5197 VDDA.n250 VDDA.n247 0.135917
R5198 VDDA.n256 VDDA.n229 0.135917
R5199 VDDA.n266 VDDA.n227 0.135917
R5200 VDDA.n270 VDDA.n267 0.135917
R5201 VDDA.n280 VDDA.n277 0.135917
R5202 VDDA.n286 VDDA.n223 0.135917
R5203 VDDA.n296 VDDA.n221 0.135917
R5204 VDDA.n300 VDDA.n297 0.135917
R5205 VDDA.n310 VDDA.n307 0.135917
R5206 VDDA.n316 VDDA.n217 0.135917
R5207 VDDA.n326 VDDA.n215 0.135917
R5208 VDDA.n330 VDDA.n327 0.135917
R5209 VDDA.n340 VDDA.n337 0.135917
R5210 VDDA.n346 VDDA.n211 0.135917
R5211 VDDA.n2564 VDDA.n2560 0.135917
R5212 VDDA.n2574 VDDA.n2555 0.135917
R5213 VDDA.n2576 VDDA.n2575 0.135917
R5214 VDDA.n2586 VDDA.n2585 0.135917
R5215 VDDA.n2594 VDDA.n2551 0.135917
R5216 VDDA.n2604 VDDA.n2549 0.135917
R5217 VDDA.n2606 VDDA.n2605 0.135917
R5218 VDDA.n2616 VDDA.n2615 0.135917
R5219 VDDA.n2624 VDDA.n2545 0.135917
R5220 VDDA.n2634 VDDA.n2543 0.135917
R5221 VDDA.n2636 VDDA.n2635 0.135917
R5222 VDDA.n2646 VDDA.n2645 0.135917
R5223 VDDA.n2654 VDDA.n2539 0.135917
R5224 VDDA.n2664 VDDA.n2537 0.135917
R5225 VDDA.n2666 VDDA.n2665 0.135917
R5226 VDDA.n2563 VDDA.n2561 0.135917
R5227 VDDA.n2573 VDDA.n2570 0.135917
R5228 VDDA.n2579 VDDA.n2554 0.135917
R5229 VDDA.n2589 VDDA.n2552 0.135917
R5230 VDDA.n2593 VDDA.n2590 0.135917
R5231 VDDA.n2603 VDDA.n2600 0.135917
R5232 VDDA.n2609 VDDA.n2548 0.135917
R5233 VDDA.n2619 VDDA.n2546 0.135917
R5234 VDDA.n2623 VDDA.n2620 0.135917
R5235 VDDA.n2633 VDDA.n2630 0.135917
R5236 VDDA.n2639 VDDA.n2542 0.135917
R5237 VDDA.n2649 VDDA.n2540 0.135917
R5238 VDDA.n2653 VDDA.n2650 0.135917
R5239 VDDA.n2663 VDDA.n2660 0.135917
R5240 VDDA.n2669 VDDA.n2536 0.135917
R5241 VDDA.n2419 VDDA.n2415 0.135917
R5242 VDDA.n2429 VDDA.n2359 0.135917
R5243 VDDA.n2431 VDDA.n2430 0.135917
R5244 VDDA.n2441 VDDA.n2440 0.135917
R5245 VDDA.n2449 VDDA.n2355 0.135917
R5246 VDDA.n2459 VDDA.n2353 0.135917
R5247 VDDA.n2461 VDDA.n2460 0.135917
R5248 VDDA.n2471 VDDA.n2470 0.135917
R5249 VDDA.n2479 VDDA.n2349 0.135917
R5250 VDDA.n2489 VDDA.n2347 0.135917
R5251 VDDA.n2491 VDDA.n2490 0.135917
R5252 VDDA.n2501 VDDA.n2500 0.135917
R5253 VDDA.n2509 VDDA.n2343 0.135917
R5254 VDDA.n2519 VDDA.n2341 0.135917
R5255 VDDA.n2521 VDDA.n2520 0.135917
R5256 VDDA.n2418 VDDA.n2416 0.135917
R5257 VDDA.n2428 VDDA.n2425 0.135917
R5258 VDDA.n2434 VDDA.n2358 0.135917
R5259 VDDA.n2444 VDDA.n2356 0.135917
R5260 VDDA.n2448 VDDA.n2445 0.135917
R5261 VDDA.n2458 VDDA.n2455 0.135917
R5262 VDDA.n2464 VDDA.n2352 0.135917
R5263 VDDA.n2474 VDDA.n2350 0.135917
R5264 VDDA.n2478 VDDA.n2475 0.135917
R5265 VDDA.n2488 VDDA.n2485 0.135917
R5266 VDDA.n2494 VDDA.n2346 0.135917
R5267 VDDA.n2504 VDDA.n2344 0.135917
R5268 VDDA.n2508 VDDA.n2505 0.135917
R5269 VDDA.n2518 VDDA.n2515 0.135917
R5270 VDDA.n2524 VDDA.n2340 0.135917
R5271 VDDA.n97 VDDA.n94 0.135917
R5272 VDDA.n101 VDDA.n81 0.135917
R5273 VDDA.n109 VDDA.n77 0.135917
R5274 VDDA.n113 VDDA.n110 0.135917
R5275 VDDA.n121 VDDA.n118 0.135917
R5276 VDDA.n125 VDDA.n69 0.135917
R5277 VDDA.n133 VDDA.n65 0.135917
R5278 VDDA.n137 VDDA.n134 0.135917
R5279 VDDA.n145 VDDA.n142 0.135917
R5280 VDDA.n149 VDDA.n57 0.135917
R5281 VDDA.n157 VDDA.n53 0.135917
R5282 VDDA.n161 VDDA.n158 0.135917
R5283 VDDA.n169 VDDA.n166 0.135917
R5284 VDDA.n173 VDDA.n45 0.135917
R5285 VDDA.n3358 VDDA.n43 0.135917
R5286 VDDA.n3249 VDDA.n3234 0.135917
R5287 VDDA.n3255 VDDA.n3232 0.135917
R5288 VDDA.n3265 VDDA.n3228 0.135917
R5289 VDDA.n3269 VDDA.n3226 0.135917
R5290 VDDA.n3279 VDDA.n3222 0.135917
R5291 VDDA.n3285 VDDA.n3220 0.135917
R5292 VDDA.n3295 VDDA.n3216 0.135917
R5293 VDDA.n3299 VDDA.n3214 0.135917
R5294 VDDA.n3309 VDDA.n3210 0.135917
R5295 VDDA.n3315 VDDA.n3208 0.135917
R5296 VDDA.n3325 VDDA.n3204 0.135917
R5297 VDDA.n3329 VDDA.n3202 0.135917
R5298 VDDA.n3339 VDDA.n3198 0.135917
R5299 VDDA.n3345 VDDA.n3196 0.135917
R5300 VDDA.n3354 VDDA.n3192 0.135917
R5301 VDDA.n3103 VDDA.n3089 0.135917
R5302 VDDA.n3107 VDDA.n3104 0.135917
R5303 VDDA.n3115 VDDA.n3112 0.135917
R5304 VDDA.n3119 VDDA.n3081 0.135917
R5305 VDDA.n3127 VDDA.n3077 0.135917
R5306 VDDA.n3131 VDDA.n3128 0.135917
R5307 VDDA.n3139 VDDA.n3136 0.135917
R5308 VDDA.n3143 VDDA.n3069 0.135917
R5309 VDDA.n3151 VDDA.n3065 0.135917
R5310 VDDA.n3155 VDDA.n3152 0.135917
R5311 VDDA.n3163 VDDA.n3160 0.135917
R5312 VDDA.n3167 VDDA.n3057 0.135917
R5313 VDDA.n3175 VDDA.n3053 0.135917
R5314 VDDA.n3179 VDDA.n3176 0.135917
R5315 VDDA.n3188 VDDA.n182 0.135917
R5316 VDDA.n2940 VDDA.n2937 0.135917
R5317 VDDA.n2944 VDDA.n2924 0.135917
R5318 VDDA.n2952 VDDA.n2920 0.135917
R5319 VDDA.n2956 VDDA.n2953 0.135917
R5320 VDDA.n2964 VDDA.n2961 0.135917
R5321 VDDA.n2968 VDDA.n2912 0.135917
R5322 VDDA.n2976 VDDA.n2908 0.135917
R5323 VDDA.n2980 VDDA.n2977 0.135917
R5324 VDDA.n2988 VDDA.n2985 0.135917
R5325 VDDA.n2992 VDDA.n2900 0.135917
R5326 VDDA.n3000 VDDA.n2896 0.135917
R5327 VDDA.n3004 VDDA.n3001 0.135917
R5328 VDDA.n3012 VDDA.n3009 0.135917
R5329 VDDA.n3016 VDDA.n2888 0.135917
R5330 VDDA.n3024 VDDA.n2886 0.135917
R5331 VDDA.n434 VDDA.n431 0.135917
R5332 VDDA.n438 VDDA.n418 0.135917
R5333 VDDA.n446 VDDA.n414 0.135917
R5334 VDDA.n450 VDDA.n447 0.135917
R5335 VDDA.n458 VDDA.n455 0.135917
R5336 VDDA.n462 VDDA.n406 0.135917
R5337 VDDA.n470 VDDA.n402 0.135917
R5338 VDDA.n474 VDDA.n471 0.135917
R5339 VDDA.n482 VDDA.n479 0.135917
R5340 VDDA.n486 VDDA.n394 0.135917
R5341 VDDA.n494 VDDA.n390 0.135917
R5342 VDDA.n498 VDDA.n495 0.135917
R5343 VDDA.n506 VDDA.n503 0.135917
R5344 VDDA.n510 VDDA.n382 0.135917
R5345 VDDA.n2858 VDDA.n380 0.135917
R5346 VDDA.n1744 VDDA.n1730 0.135917
R5347 VDDA.n1748 VDDA.n1745 0.135917
R5348 VDDA.n1756 VDDA.n1753 0.135917
R5349 VDDA.n1760 VDDA.n1722 0.135917
R5350 VDDA.n1768 VDDA.n1718 0.135917
R5351 VDDA.n1772 VDDA.n1769 0.135917
R5352 VDDA.n1780 VDDA.n1777 0.135917
R5353 VDDA.n1784 VDDA.n1710 0.135917
R5354 VDDA.n1792 VDDA.n1706 0.135917
R5355 VDDA.n1796 VDDA.n1793 0.135917
R5356 VDDA.n1804 VDDA.n1801 0.135917
R5357 VDDA.n1808 VDDA.n1698 0.135917
R5358 VDDA.n1816 VDDA.n1694 0.135917
R5359 VDDA.n1820 VDDA.n1817 0.135917
R5360 VDDA.n2680 VDDA.n519 0.135917
R5361 VDDA.n1581 VDDA.n1578 0.135917
R5362 VDDA.n1585 VDDA.n1565 0.135917
R5363 VDDA.n1593 VDDA.n1561 0.135917
R5364 VDDA.n1597 VDDA.n1594 0.135917
R5365 VDDA.n1605 VDDA.n1602 0.135917
R5366 VDDA.n1609 VDDA.n1553 0.135917
R5367 VDDA.n1617 VDDA.n1549 0.135917
R5368 VDDA.n1621 VDDA.n1618 0.135917
R5369 VDDA.n1629 VDDA.n1626 0.135917
R5370 VDDA.n1633 VDDA.n1541 0.135917
R5371 VDDA.n1641 VDDA.n1537 0.135917
R5372 VDDA.n1645 VDDA.n1642 0.135917
R5373 VDDA.n1653 VDDA.n1650 0.135917
R5374 VDDA.n1657 VDDA.n1529 0.135917
R5375 VDDA.n1665 VDDA.n1527 0.135917
R5376 VDDA.n601 VDDA.n598 0.135917
R5377 VDDA.n605 VDDA.n585 0.135917
R5378 VDDA.n613 VDDA.n581 0.135917
R5379 VDDA.n617 VDDA.n614 0.135917
R5380 VDDA.n625 VDDA.n622 0.135917
R5381 VDDA.n629 VDDA.n573 0.135917
R5382 VDDA.n637 VDDA.n569 0.135917
R5383 VDDA.n641 VDDA.n638 0.135917
R5384 VDDA.n649 VDDA.n646 0.135917
R5385 VDDA.n653 VDDA.n561 0.135917
R5386 VDDA.n661 VDDA.n557 0.135917
R5387 VDDA.n665 VDDA.n662 0.135917
R5388 VDDA.n673 VDDA.n670 0.135917
R5389 VDDA.n677 VDDA.n549 0.135917
R5390 VDDA.n1499 VDDA.n547 0.135917
R5391 VDDA.n1389 VDDA.n1374 0.135917
R5392 VDDA.n1395 VDDA.n1372 0.135917
R5393 VDDA.n1405 VDDA.n1368 0.135917
R5394 VDDA.n1409 VDDA.n1366 0.135917
R5395 VDDA.n1419 VDDA.n1362 0.135917
R5396 VDDA.n1425 VDDA.n1360 0.135917
R5397 VDDA.n1435 VDDA.n1356 0.135917
R5398 VDDA.n1439 VDDA.n1354 0.135917
R5399 VDDA.n1449 VDDA.n1350 0.135917
R5400 VDDA.n1455 VDDA.n1348 0.135917
R5401 VDDA.n1465 VDDA.n1344 0.135917
R5402 VDDA.n1469 VDDA.n1342 0.135917
R5403 VDDA.n1479 VDDA.n1338 0.135917
R5404 VDDA.n1485 VDDA.n1336 0.135917
R5405 VDDA.n1494 VDDA.n1332 0.135917
R5406 VDDA.n1226 VDDA.n1212 0.135917
R5407 VDDA.n1230 VDDA.n1227 0.135917
R5408 VDDA.n1240 VDDA.n1237 0.135917
R5409 VDDA.n1246 VDDA.n1208 0.135917
R5410 VDDA.n1256 VDDA.n1206 0.135917
R5411 VDDA.n1260 VDDA.n1257 0.135917
R5412 VDDA.n1270 VDDA.n1267 0.135917
R5413 VDDA.n1276 VDDA.n1202 0.135917
R5414 VDDA.n1286 VDDA.n1200 0.135917
R5415 VDDA.n1290 VDDA.n1287 0.135917
R5416 VDDA.n1300 VDDA.n1297 0.135917
R5417 VDDA.n1306 VDDA.n1196 0.135917
R5418 VDDA.n1316 VDDA.n1194 0.135917
R5419 VDDA.n1320 VDDA.n1317 0.135917
R5420 VDDA.n1329 VDDA.n685 0.135917
R5421 VDDA.n2217 VDDA.n2181 0.1255
R5422 VDDA.n2234 VDDA.n2233 0.1255
R5423 VDDA.n2245 VDDA.n2170 0.1255
R5424 VDDA.n2264 VDDA.n2263 0.1255
R5425 VDDA.n2275 VDDA.n2164 0.1255
R5426 VDDA.n2294 VDDA.n2293 0.1255
R5427 VDDA.n2305 VDDA.n2158 0.1255
R5428 VDDA.n2324 VDDA.n2323 0.1255
R5429 VDDA.n2232 VDDA.n2173 0.1255
R5430 VDDA.n2249 VDDA.n2248 0.1255
R5431 VDDA.n2262 VDDA.n2167 0.1255
R5432 VDDA.n2279 VDDA.n2278 0.1255
R5433 VDDA.n2292 VDDA.n2161 0.1255
R5434 VDDA.n2309 VDDA.n2308 0.1255
R5435 VDDA.n2322 VDDA.n2155 0.1255
R5436 VDDA.n2049 VDDA.n2048 0.1255
R5437 VDDA.n2060 VDDA.n1941 0.1255
R5438 VDDA.n2079 VDDA.n2078 0.1255
R5439 VDDA.n2090 VDDA.n1935 0.1255
R5440 VDDA.n2109 VDDA.n2108 0.1255
R5441 VDDA.n2120 VDDA.n1929 0.1255
R5442 VDDA.n2139 VDDA.n2138 0.1255
R5443 VDDA.n2047 VDDA.n1944 0.1255
R5444 VDDA.n2064 VDDA.n2063 0.1255
R5445 VDDA.n2077 VDDA.n1938 0.1255
R5446 VDDA.n2094 VDDA.n2093 0.1255
R5447 VDDA.n2107 VDDA.n1932 0.1255
R5448 VDDA.n2124 VDDA.n2123 0.1255
R5449 VDDA.n2137 VDDA.n1926 0.1255
R5450 VDDA.n252 VDDA.n251 0.1255
R5451 VDDA.n263 VDDA.n226 0.1255
R5452 VDDA.n282 VDDA.n281 0.1255
R5453 VDDA.n293 VDDA.n220 0.1255
R5454 VDDA.n312 VDDA.n311 0.1255
R5455 VDDA.n323 VDDA.n214 0.1255
R5456 VDDA.n342 VDDA.n341 0.1255
R5457 VDDA.n250 VDDA.n229 0.1255
R5458 VDDA.n267 VDDA.n266 0.1255
R5459 VDDA.n280 VDDA.n223 0.1255
R5460 VDDA.n297 VDDA.n296 0.1255
R5461 VDDA.n310 VDDA.n217 0.1255
R5462 VDDA.n327 VDDA.n326 0.1255
R5463 VDDA.n340 VDDA.n211 0.1255
R5464 VDDA.n2575 VDDA.n2574 0.1255
R5465 VDDA.n2586 VDDA.n2551 0.1255
R5466 VDDA.n2605 VDDA.n2604 0.1255
R5467 VDDA.n2616 VDDA.n2545 0.1255
R5468 VDDA.n2635 VDDA.n2634 0.1255
R5469 VDDA.n2646 VDDA.n2539 0.1255
R5470 VDDA.n2665 VDDA.n2664 0.1255
R5471 VDDA.n2573 VDDA.n2554 0.1255
R5472 VDDA.n2590 VDDA.n2589 0.1255
R5473 VDDA.n2603 VDDA.n2548 0.1255
R5474 VDDA.n2620 VDDA.n2619 0.1255
R5475 VDDA.n2633 VDDA.n2542 0.1255
R5476 VDDA.n2650 VDDA.n2649 0.1255
R5477 VDDA.n2663 VDDA.n2536 0.1255
R5478 VDDA.n2414 VDDA.n2362 0.1255
R5479 VDDA.n2365 VDDA.n2362 0.1255
R5480 VDDA.n2367 VDDA.n2365 0.1255
R5481 VDDA.n2369 VDDA.n2367 0.1255
R5482 VDDA.n2371 VDDA.n2369 0.1255
R5483 VDDA.n2373 VDDA.n2371 0.1255
R5484 VDDA.n2375 VDDA.n2373 0.1255
R5485 VDDA.n2377 VDDA.n2375 0.1255
R5486 VDDA.n2379 VDDA.n2377 0.1255
R5487 VDDA.n2408 VDDA.n2379 0.1255
R5488 VDDA.n2407 VDDA.n2381 0.1255
R5489 VDDA.n2385 VDDA.n2381 0.1255
R5490 VDDA.n2387 VDDA.n2385 0.1255
R5491 VDDA.n2389 VDDA.n2387 0.1255
R5492 VDDA.n2391 VDDA.n2389 0.1255
R5493 VDDA.n2393 VDDA.n2391 0.1255
R5494 VDDA.n2395 VDDA.n2393 0.1255
R5495 VDDA.n2397 VDDA.n2395 0.1255
R5496 VDDA.n2399 VDDA.n2397 0.1255
R5497 VDDA.n2430 VDDA.n2429 0.1255
R5498 VDDA.n2441 VDDA.n2355 0.1255
R5499 VDDA.n2460 VDDA.n2459 0.1255
R5500 VDDA.n2471 VDDA.n2349 0.1255
R5501 VDDA.n2490 VDDA.n2489 0.1255
R5502 VDDA.n2501 VDDA.n2343 0.1255
R5503 VDDA.n2520 VDDA.n2519 0.1255
R5504 VDDA.n2428 VDDA.n2358 0.1255
R5505 VDDA.n2445 VDDA.n2444 0.1255
R5506 VDDA.n2458 VDDA.n2352 0.1255
R5507 VDDA.n2475 VDDA.n2474 0.1255
R5508 VDDA.n2488 VDDA.n2346 0.1255
R5509 VDDA.n2505 VDDA.n2504 0.1255
R5510 VDDA.n2518 VDDA.n2340 0.1255
R5511 VDDA.n97 VDDA.n81 0.1255
R5512 VDDA.n110 VDDA.n109 0.1255
R5513 VDDA.n121 VDDA.n69 0.1255
R5514 VDDA.n134 VDDA.n133 0.1255
R5515 VDDA.n145 VDDA.n57 0.1255
R5516 VDDA.n158 VDDA.n157 0.1255
R5517 VDDA.n169 VDDA.n45 0.1255
R5518 VDDA.n3249 VDDA.n3232 0.1255
R5519 VDDA.n3265 VDDA.n3226 0.1255
R5520 VDDA.n3279 VDDA.n3220 0.1255
R5521 VDDA.n3295 VDDA.n3214 0.1255
R5522 VDDA.n3309 VDDA.n3208 0.1255
R5523 VDDA.n3325 VDDA.n3202 0.1255
R5524 VDDA.n3339 VDDA.n3196 0.1255
R5525 VDDA.n3104 VDDA.n3103 0.1255
R5526 VDDA.n3115 VDDA.n3081 0.1255
R5527 VDDA.n3128 VDDA.n3127 0.1255
R5528 VDDA.n3139 VDDA.n3069 0.1255
R5529 VDDA.n3152 VDDA.n3151 0.1255
R5530 VDDA.n3163 VDDA.n3057 0.1255
R5531 VDDA.n3176 VDDA.n3175 0.1255
R5532 VDDA.n2940 VDDA.n2924 0.1255
R5533 VDDA.n2953 VDDA.n2952 0.1255
R5534 VDDA.n2964 VDDA.n2912 0.1255
R5535 VDDA.n2977 VDDA.n2976 0.1255
R5536 VDDA.n2988 VDDA.n2900 0.1255
R5537 VDDA.n3001 VDDA.n3000 0.1255
R5538 VDDA.n3012 VDDA.n2888 0.1255
R5539 VDDA.n434 VDDA.n418 0.1255
R5540 VDDA.n447 VDDA.n446 0.1255
R5541 VDDA.n458 VDDA.n406 0.1255
R5542 VDDA.n471 VDDA.n470 0.1255
R5543 VDDA.n482 VDDA.n394 0.1255
R5544 VDDA.n495 VDDA.n494 0.1255
R5545 VDDA.n506 VDDA.n382 0.1255
R5546 VDDA.n1745 VDDA.n1744 0.1255
R5547 VDDA.n1756 VDDA.n1722 0.1255
R5548 VDDA.n1769 VDDA.n1768 0.1255
R5549 VDDA.n1780 VDDA.n1710 0.1255
R5550 VDDA.n1793 VDDA.n1792 0.1255
R5551 VDDA.n1804 VDDA.n1698 0.1255
R5552 VDDA.n1817 VDDA.n1816 0.1255
R5553 VDDA.n1581 VDDA.n1565 0.1255
R5554 VDDA.n1594 VDDA.n1593 0.1255
R5555 VDDA.n1605 VDDA.n1553 0.1255
R5556 VDDA.n1618 VDDA.n1617 0.1255
R5557 VDDA.n1629 VDDA.n1541 0.1255
R5558 VDDA.n1642 VDDA.n1641 0.1255
R5559 VDDA.n1653 VDDA.n1529 0.1255
R5560 VDDA.n601 VDDA.n585 0.1255
R5561 VDDA.n614 VDDA.n613 0.1255
R5562 VDDA.n625 VDDA.n573 0.1255
R5563 VDDA.n638 VDDA.n637 0.1255
R5564 VDDA.n649 VDDA.n561 0.1255
R5565 VDDA.n662 VDDA.n661 0.1255
R5566 VDDA.n673 VDDA.n549 0.1255
R5567 VDDA.n1389 VDDA.n1372 0.1255
R5568 VDDA.n1405 VDDA.n1366 0.1255
R5569 VDDA.n1419 VDDA.n1360 0.1255
R5570 VDDA.n1435 VDDA.n1354 0.1255
R5571 VDDA.n1449 VDDA.n1348 0.1255
R5572 VDDA.n1465 VDDA.n1342 0.1255
R5573 VDDA.n1479 VDDA.n1336 0.1255
R5574 VDDA.n1227 VDDA.n1226 0.1255
R5575 VDDA.n1240 VDDA.n1208 0.1255
R5576 VDDA.n1257 VDDA.n1256 0.1255
R5577 VDDA.n1270 VDDA.n1202 0.1255
R5578 VDDA.n1287 VDDA.n1286 0.1255
R5579 VDDA.n1300 VDDA.n1196 0.1255
R5580 VDDA.n1317 VDDA.n1316 0.1255
R5581 VDDA.n2216 VDDA.n2215 0.115083
R5582 VDDA.n2215 VDDA.n2214 0.115083
R5583 VDDA.n2214 VDDA.n2213 0.115083
R5584 VDDA.n2211 VDDA.n2210 0.115083
R5585 VDDA.n2210 VDDA.n2209 0.115083
R5586 VDDA.n2209 VDDA.n2208 0.115083
R5587 VDDA.n2208 VDDA.n2207 0.115083
R5588 VDDA.n2205 VDDA.n2204 0.115083
R5589 VDDA.n2204 VDDA.n2203 0.115083
R5590 VDDA.n2031 VDDA.n2007 0.0864375
R5591 VDDA.n92 VDDA.n91 0.0734167
R5592 VDDA.n92 VDDA.n84 0.0734167
R5593 VDDA.n100 VDDA.n80 0.0734167
R5594 VDDA.n106 VDDA.n80 0.0734167
R5595 VDDA.n107 VDDA.n106 0.0734167
R5596 VDDA.n115 VDDA.n114 0.0734167
R5597 VDDA.n116 VDDA.n115 0.0734167
R5598 VDDA.n116 VDDA.n72 0.0734167
R5599 VDDA.n124 VDDA.n68 0.0734167
R5600 VDDA.n130 VDDA.n68 0.0734167
R5601 VDDA.n131 VDDA.n130 0.0734167
R5602 VDDA.n139 VDDA.n138 0.0734167
R5603 VDDA.n140 VDDA.n139 0.0734167
R5604 VDDA.n140 VDDA.n60 0.0734167
R5605 VDDA.n148 VDDA.n56 0.0734167
R5606 VDDA.n154 VDDA.n56 0.0734167
R5607 VDDA.n155 VDDA.n154 0.0734167
R5608 VDDA.n163 VDDA.n162 0.0734167
R5609 VDDA.n164 VDDA.n163 0.0734167
R5610 VDDA.n164 VDDA.n48 0.0734167
R5611 VDDA.n172 VDDA.n44 0.0734167
R5612 VDDA.n178 VDDA.n44 0.0734167
R5613 VDDA.n179 VDDA.n178 0.0734167
R5614 VDDA.n3246 VDDA.n3235 0.0734167
R5615 VDDA.n3247 VDDA.n3246 0.0734167
R5616 VDDA.n3257 VDDA.n3256 0.0734167
R5617 VDDA.n3258 VDDA.n3257 0.0734167
R5618 VDDA.n3258 VDDA.n3227 0.0734167
R5619 VDDA.n3268 VDDA.n3223 0.0734167
R5620 VDDA.n3276 VDDA.n3223 0.0734167
R5621 VDDA.n3277 VDDA.n3276 0.0734167
R5622 VDDA.n3287 VDDA.n3286 0.0734167
R5623 VDDA.n3288 VDDA.n3287 0.0734167
R5624 VDDA.n3288 VDDA.n3215 0.0734167
R5625 VDDA.n3298 VDDA.n3211 0.0734167
R5626 VDDA.n3306 VDDA.n3211 0.0734167
R5627 VDDA.n3307 VDDA.n3306 0.0734167
R5628 VDDA.n3317 VDDA.n3316 0.0734167
R5629 VDDA.n3318 VDDA.n3317 0.0734167
R5630 VDDA.n3318 VDDA.n3203 0.0734167
R5631 VDDA.n3328 VDDA.n3199 0.0734167
R5632 VDDA.n3336 VDDA.n3199 0.0734167
R5633 VDDA.n3337 VDDA.n3336 0.0734167
R5634 VDDA.n3347 VDDA.n3346 0.0734167
R5635 VDDA.n3348 VDDA.n3347 0.0734167
R5636 VDDA.n3348 VDDA.n3191 0.0734167
R5637 VDDA.n3100 VDDA.n3092 0.0734167
R5638 VDDA.n3101 VDDA.n3100 0.0734167
R5639 VDDA.n3109 VDDA.n3108 0.0734167
R5640 VDDA.n3110 VDDA.n3109 0.0734167
R5641 VDDA.n3110 VDDA.n3084 0.0734167
R5642 VDDA.n3118 VDDA.n3080 0.0734167
R5643 VDDA.n3124 VDDA.n3080 0.0734167
R5644 VDDA.n3125 VDDA.n3124 0.0734167
R5645 VDDA.n3133 VDDA.n3132 0.0734167
R5646 VDDA.n3134 VDDA.n3133 0.0734167
R5647 VDDA.n3134 VDDA.n3072 0.0734167
R5648 VDDA.n3142 VDDA.n3068 0.0734167
R5649 VDDA.n3148 VDDA.n3068 0.0734167
R5650 VDDA.n3149 VDDA.n3148 0.0734167
R5651 VDDA.n3157 VDDA.n3156 0.0734167
R5652 VDDA.n3158 VDDA.n3157 0.0734167
R5653 VDDA.n3158 VDDA.n3060 0.0734167
R5654 VDDA.n3166 VDDA.n3056 0.0734167
R5655 VDDA.n3172 VDDA.n3056 0.0734167
R5656 VDDA.n3173 VDDA.n3172 0.0734167
R5657 VDDA.n3181 VDDA.n3180 0.0734167
R5658 VDDA.n3182 VDDA.n3181 0.0734167
R5659 VDDA.n3182 VDDA.n181 0.0734167
R5660 VDDA.n2935 VDDA.n2934 0.0734167
R5661 VDDA.n2935 VDDA.n2927 0.0734167
R5662 VDDA.n2943 VDDA.n2923 0.0734167
R5663 VDDA.n2949 VDDA.n2923 0.0734167
R5664 VDDA.n2950 VDDA.n2949 0.0734167
R5665 VDDA.n2958 VDDA.n2957 0.0734167
R5666 VDDA.n2959 VDDA.n2958 0.0734167
R5667 VDDA.n2959 VDDA.n2915 0.0734167
R5668 VDDA.n2967 VDDA.n2911 0.0734167
R5669 VDDA.n2973 VDDA.n2911 0.0734167
R5670 VDDA.n2974 VDDA.n2973 0.0734167
R5671 VDDA.n2982 VDDA.n2981 0.0734167
R5672 VDDA.n2983 VDDA.n2982 0.0734167
R5673 VDDA.n2983 VDDA.n2903 0.0734167
R5674 VDDA.n2991 VDDA.n2899 0.0734167
R5675 VDDA.n2997 VDDA.n2899 0.0734167
R5676 VDDA.n2998 VDDA.n2997 0.0734167
R5677 VDDA.n3006 VDDA.n3005 0.0734167
R5678 VDDA.n3007 VDDA.n3006 0.0734167
R5679 VDDA.n3007 VDDA.n2891 0.0734167
R5680 VDDA.n3015 VDDA.n2887 0.0734167
R5681 VDDA.n3021 VDDA.n2887 0.0734167
R5682 VDDA.n3022 VDDA.n3021 0.0734167
R5683 VDDA.n429 VDDA.n428 0.0734167
R5684 VDDA.n429 VDDA.n421 0.0734167
R5685 VDDA.n437 VDDA.n417 0.0734167
R5686 VDDA.n443 VDDA.n417 0.0734167
R5687 VDDA.n444 VDDA.n443 0.0734167
R5688 VDDA.n452 VDDA.n451 0.0734167
R5689 VDDA.n453 VDDA.n452 0.0734167
R5690 VDDA.n453 VDDA.n409 0.0734167
R5691 VDDA.n461 VDDA.n405 0.0734167
R5692 VDDA.n467 VDDA.n405 0.0734167
R5693 VDDA.n468 VDDA.n467 0.0734167
R5694 VDDA.n476 VDDA.n475 0.0734167
R5695 VDDA.n477 VDDA.n476 0.0734167
R5696 VDDA.n477 VDDA.n397 0.0734167
R5697 VDDA.n485 VDDA.n393 0.0734167
R5698 VDDA.n491 VDDA.n393 0.0734167
R5699 VDDA.n492 VDDA.n491 0.0734167
R5700 VDDA.n500 VDDA.n499 0.0734167
R5701 VDDA.n501 VDDA.n500 0.0734167
R5702 VDDA.n501 VDDA.n385 0.0734167
R5703 VDDA.n509 VDDA.n381 0.0734167
R5704 VDDA.n515 VDDA.n381 0.0734167
R5705 VDDA.n516 VDDA.n515 0.0734167
R5706 VDDA.n1741 VDDA.n1733 0.0734167
R5707 VDDA.n1742 VDDA.n1741 0.0734167
R5708 VDDA.n1750 VDDA.n1749 0.0734167
R5709 VDDA.n1751 VDDA.n1750 0.0734167
R5710 VDDA.n1751 VDDA.n1725 0.0734167
R5711 VDDA.n1759 VDDA.n1721 0.0734167
R5712 VDDA.n1765 VDDA.n1721 0.0734167
R5713 VDDA.n1766 VDDA.n1765 0.0734167
R5714 VDDA.n1774 VDDA.n1773 0.0734167
R5715 VDDA.n1775 VDDA.n1774 0.0734167
R5716 VDDA.n1775 VDDA.n1713 0.0734167
R5717 VDDA.n1783 VDDA.n1709 0.0734167
R5718 VDDA.n1789 VDDA.n1709 0.0734167
R5719 VDDA.n1790 VDDA.n1789 0.0734167
R5720 VDDA.n1798 VDDA.n1797 0.0734167
R5721 VDDA.n1799 VDDA.n1798 0.0734167
R5722 VDDA.n1799 VDDA.n1701 0.0734167
R5723 VDDA.n1807 VDDA.n1697 0.0734167
R5724 VDDA.n1813 VDDA.n1697 0.0734167
R5725 VDDA.n1814 VDDA.n1813 0.0734167
R5726 VDDA.n1822 VDDA.n1821 0.0734167
R5727 VDDA.n1823 VDDA.n1822 0.0734167
R5728 VDDA.n1823 VDDA.n518 0.0734167
R5729 VDDA.n1576 VDDA.n1575 0.0734167
R5730 VDDA.n1576 VDDA.n1568 0.0734167
R5731 VDDA.n1584 VDDA.n1564 0.0734167
R5732 VDDA.n1590 VDDA.n1564 0.0734167
R5733 VDDA.n1591 VDDA.n1590 0.0734167
R5734 VDDA.n1599 VDDA.n1598 0.0734167
R5735 VDDA.n1600 VDDA.n1599 0.0734167
R5736 VDDA.n1600 VDDA.n1556 0.0734167
R5737 VDDA.n1608 VDDA.n1552 0.0734167
R5738 VDDA.n1614 VDDA.n1552 0.0734167
R5739 VDDA.n1615 VDDA.n1614 0.0734167
R5740 VDDA.n1623 VDDA.n1622 0.0734167
R5741 VDDA.n1624 VDDA.n1623 0.0734167
R5742 VDDA.n1624 VDDA.n1544 0.0734167
R5743 VDDA.n1632 VDDA.n1540 0.0734167
R5744 VDDA.n1638 VDDA.n1540 0.0734167
R5745 VDDA.n1639 VDDA.n1638 0.0734167
R5746 VDDA.n1647 VDDA.n1646 0.0734167
R5747 VDDA.n1648 VDDA.n1647 0.0734167
R5748 VDDA.n1648 VDDA.n1532 0.0734167
R5749 VDDA.n1656 VDDA.n1528 0.0734167
R5750 VDDA.n1662 VDDA.n1528 0.0734167
R5751 VDDA.n1663 VDDA.n1662 0.0734167
R5752 VDDA.n596 VDDA.n595 0.0734167
R5753 VDDA.n596 VDDA.n588 0.0734167
R5754 VDDA.n604 VDDA.n584 0.0734167
R5755 VDDA.n610 VDDA.n584 0.0734167
R5756 VDDA.n611 VDDA.n610 0.0734167
R5757 VDDA.n619 VDDA.n618 0.0734167
R5758 VDDA.n620 VDDA.n619 0.0734167
R5759 VDDA.n620 VDDA.n576 0.0734167
R5760 VDDA.n628 VDDA.n572 0.0734167
R5761 VDDA.n634 VDDA.n572 0.0734167
R5762 VDDA.n635 VDDA.n634 0.0734167
R5763 VDDA.n643 VDDA.n642 0.0734167
R5764 VDDA.n644 VDDA.n643 0.0734167
R5765 VDDA.n644 VDDA.n564 0.0734167
R5766 VDDA.n652 VDDA.n560 0.0734167
R5767 VDDA.n658 VDDA.n560 0.0734167
R5768 VDDA.n659 VDDA.n658 0.0734167
R5769 VDDA.n667 VDDA.n666 0.0734167
R5770 VDDA.n668 VDDA.n667 0.0734167
R5771 VDDA.n668 VDDA.n552 0.0734167
R5772 VDDA.n676 VDDA.n548 0.0734167
R5773 VDDA.n682 VDDA.n548 0.0734167
R5774 VDDA.n683 VDDA.n682 0.0734167
R5775 VDDA.n1386 VDDA.n1375 0.0734167
R5776 VDDA.n1387 VDDA.n1386 0.0734167
R5777 VDDA.n1397 VDDA.n1396 0.0734167
R5778 VDDA.n1398 VDDA.n1397 0.0734167
R5779 VDDA.n1398 VDDA.n1367 0.0734167
R5780 VDDA.n1408 VDDA.n1363 0.0734167
R5781 VDDA.n1416 VDDA.n1363 0.0734167
R5782 VDDA.n1417 VDDA.n1416 0.0734167
R5783 VDDA.n1427 VDDA.n1426 0.0734167
R5784 VDDA.n1428 VDDA.n1427 0.0734167
R5785 VDDA.n1428 VDDA.n1355 0.0734167
R5786 VDDA.n1438 VDDA.n1351 0.0734167
R5787 VDDA.n1446 VDDA.n1351 0.0734167
R5788 VDDA.n1447 VDDA.n1446 0.0734167
R5789 VDDA.n1457 VDDA.n1456 0.0734167
R5790 VDDA.n1458 VDDA.n1457 0.0734167
R5791 VDDA.n1458 VDDA.n1343 0.0734167
R5792 VDDA.n1468 VDDA.n1339 0.0734167
R5793 VDDA.n1476 VDDA.n1339 0.0734167
R5794 VDDA.n1477 VDDA.n1476 0.0734167
R5795 VDDA.n1487 VDDA.n1486 0.0734167
R5796 VDDA.n1488 VDDA.n1487 0.0734167
R5797 VDDA.n1488 VDDA.n1331 0.0734167
R5798 VDDA.n1221 VDDA.n1213 0.0734167
R5799 VDDA.n1222 VDDA.n1221 0.0734167
R5800 VDDA.n1232 VDDA.n1231 0.0734167
R5801 VDDA.n1233 VDDA.n1232 0.0734167
R5802 VDDA.n1233 VDDA.n1209 0.0734167
R5803 VDDA.n1243 VDDA.n1207 0.0734167
R5804 VDDA.n1251 VDDA.n1207 0.0734167
R5805 VDDA.n1252 VDDA.n1251 0.0734167
R5806 VDDA.n1262 VDDA.n1261 0.0734167
R5807 VDDA.n1263 VDDA.n1262 0.0734167
R5808 VDDA.n1263 VDDA.n1203 0.0734167
R5809 VDDA.n1273 VDDA.n1201 0.0734167
R5810 VDDA.n1281 VDDA.n1201 0.0734167
R5811 VDDA.n1282 VDDA.n1281 0.0734167
R5812 VDDA.n1292 VDDA.n1291 0.0734167
R5813 VDDA.n1293 VDDA.n1292 0.0734167
R5814 VDDA.n1293 VDDA.n1197 0.0734167
R5815 VDDA.n1303 VDDA.n1195 0.0734167
R5816 VDDA.n1311 VDDA.n1195 0.0734167
R5817 VDDA.n1312 VDDA.n1311 0.0734167
R5818 VDDA.n1322 VDDA.n1321 0.0734167
R5819 VDDA.n1323 VDDA.n1322 0.0734167
R5820 VDDA.n1323 VDDA.n684 0.0734167
R5821 VDDA.n2212 VDDA.n2211 0.0682083
R5822 VDDA.n2207 VDDA.n2206 0.0682083
R5823 VDDA.n98 VDDA.n84 0.0682083
R5824 VDDA.n100 VDDA.n99 0.0682083
R5825 VDDA.n108 VDDA.n107 0.0682083
R5826 VDDA.n114 VDDA.n76 0.0682083
R5827 VDDA.n122 VDDA.n72 0.0682083
R5828 VDDA.n124 VDDA.n123 0.0682083
R5829 VDDA.n132 VDDA.n131 0.0682083
R5830 VDDA.n138 VDDA.n64 0.0682083
R5831 VDDA.n146 VDDA.n60 0.0682083
R5832 VDDA.n148 VDDA.n147 0.0682083
R5833 VDDA.n156 VDDA.n155 0.0682083
R5834 VDDA.n162 VDDA.n52 0.0682083
R5835 VDDA.n170 VDDA.n48 0.0682083
R5836 VDDA.n172 VDDA.n171 0.0682083
R5837 VDDA.n3357 VDDA.n179 0.0682083
R5838 VDDA.n3248 VDDA.n3247 0.0682083
R5839 VDDA.n3256 VDDA.n3231 0.0682083
R5840 VDDA.n3266 VDDA.n3227 0.0682083
R5841 VDDA.n3268 VDDA.n3267 0.0682083
R5842 VDDA.n3278 VDDA.n3277 0.0682083
R5843 VDDA.n3286 VDDA.n3219 0.0682083
R5844 VDDA.n3296 VDDA.n3215 0.0682083
R5845 VDDA.n3298 VDDA.n3297 0.0682083
R5846 VDDA.n3308 VDDA.n3307 0.0682083
R5847 VDDA.n3316 VDDA.n3207 0.0682083
R5848 VDDA.n3326 VDDA.n3203 0.0682083
R5849 VDDA.n3328 VDDA.n3327 0.0682083
R5850 VDDA.n3338 VDDA.n3337 0.0682083
R5851 VDDA.n3346 VDDA.n3195 0.0682083
R5852 VDDA.n3355 VDDA.n3191 0.0682083
R5853 VDDA.n3102 VDDA.n3101 0.0682083
R5854 VDDA.n3108 VDDA.n3088 0.0682083
R5855 VDDA.n3116 VDDA.n3084 0.0682083
R5856 VDDA.n3118 VDDA.n3117 0.0682083
R5857 VDDA.n3126 VDDA.n3125 0.0682083
R5858 VDDA.n3132 VDDA.n3076 0.0682083
R5859 VDDA.n3140 VDDA.n3072 0.0682083
R5860 VDDA.n3142 VDDA.n3141 0.0682083
R5861 VDDA.n3150 VDDA.n3149 0.0682083
R5862 VDDA.n3156 VDDA.n3064 0.0682083
R5863 VDDA.n3164 VDDA.n3060 0.0682083
R5864 VDDA.n3166 VDDA.n3165 0.0682083
R5865 VDDA.n3174 VDDA.n3173 0.0682083
R5866 VDDA.n3180 VDDA.n3052 0.0682083
R5867 VDDA.n3189 VDDA.n181 0.0682083
R5868 VDDA.n2941 VDDA.n2927 0.0682083
R5869 VDDA.n2943 VDDA.n2942 0.0682083
R5870 VDDA.n2951 VDDA.n2950 0.0682083
R5871 VDDA.n2957 VDDA.n2919 0.0682083
R5872 VDDA.n2965 VDDA.n2915 0.0682083
R5873 VDDA.n2967 VDDA.n2966 0.0682083
R5874 VDDA.n2975 VDDA.n2974 0.0682083
R5875 VDDA.n2981 VDDA.n2907 0.0682083
R5876 VDDA.n2989 VDDA.n2903 0.0682083
R5877 VDDA.n2991 VDDA.n2990 0.0682083
R5878 VDDA.n2999 VDDA.n2998 0.0682083
R5879 VDDA.n3005 VDDA.n2895 0.0682083
R5880 VDDA.n3013 VDDA.n2891 0.0682083
R5881 VDDA.n3015 VDDA.n3014 0.0682083
R5882 VDDA.n3023 VDDA.n3022 0.0682083
R5883 VDDA.n435 VDDA.n421 0.0682083
R5884 VDDA.n437 VDDA.n436 0.0682083
R5885 VDDA.n445 VDDA.n444 0.0682083
R5886 VDDA.n451 VDDA.n413 0.0682083
R5887 VDDA.n459 VDDA.n409 0.0682083
R5888 VDDA.n461 VDDA.n460 0.0682083
R5889 VDDA.n469 VDDA.n468 0.0682083
R5890 VDDA.n475 VDDA.n401 0.0682083
R5891 VDDA.n483 VDDA.n397 0.0682083
R5892 VDDA.n485 VDDA.n484 0.0682083
R5893 VDDA.n493 VDDA.n492 0.0682083
R5894 VDDA.n499 VDDA.n389 0.0682083
R5895 VDDA.n507 VDDA.n385 0.0682083
R5896 VDDA.n509 VDDA.n508 0.0682083
R5897 VDDA.n2857 VDDA.n516 0.0682083
R5898 VDDA.n1743 VDDA.n1742 0.0682083
R5899 VDDA.n1749 VDDA.n1729 0.0682083
R5900 VDDA.n1757 VDDA.n1725 0.0682083
R5901 VDDA.n1759 VDDA.n1758 0.0682083
R5902 VDDA.n1767 VDDA.n1766 0.0682083
R5903 VDDA.n1773 VDDA.n1717 0.0682083
R5904 VDDA.n1781 VDDA.n1713 0.0682083
R5905 VDDA.n1783 VDDA.n1782 0.0682083
R5906 VDDA.n1791 VDDA.n1790 0.0682083
R5907 VDDA.n1797 VDDA.n1705 0.0682083
R5908 VDDA.n1805 VDDA.n1701 0.0682083
R5909 VDDA.n1807 VDDA.n1806 0.0682083
R5910 VDDA.n1815 VDDA.n1814 0.0682083
R5911 VDDA.n1821 VDDA.n1693 0.0682083
R5912 VDDA.n2681 VDDA.n518 0.0682083
R5913 VDDA.n1582 VDDA.n1568 0.0682083
R5914 VDDA.n1584 VDDA.n1583 0.0682083
R5915 VDDA.n1592 VDDA.n1591 0.0682083
R5916 VDDA.n1598 VDDA.n1560 0.0682083
R5917 VDDA.n1606 VDDA.n1556 0.0682083
R5918 VDDA.n1608 VDDA.n1607 0.0682083
R5919 VDDA.n1616 VDDA.n1615 0.0682083
R5920 VDDA.n1622 VDDA.n1548 0.0682083
R5921 VDDA.n1630 VDDA.n1544 0.0682083
R5922 VDDA.n1632 VDDA.n1631 0.0682083
R5923 VDDA.n1640 VDDA.n1639 0.0682083
R5924 VDDA.n1646 VDDA.n1536 0.0682083
R5925 VDDA.n1654 VDDA.n1532 0.0682083
R5926 VDDA.n1656 VDDA.n1655 0.0682083
R5927 VDDA.n1664 VDDA.n1663 0.0682083
R5928 VDDA.n602 VDDA.n588 0.0682083
R5929 VDDA.n604 VDDA.n603 0.0682083
R5930 VDDA.n612 VDDA.n611 0.0682083
R5931 VDDA.n618 VDDA.n580 0.0682083
R5932 VDDA.n626 VDDA.n576 0.0682083
R5933 VDDA.n628 VDDA.n627 0.0682083
R5934 VDDA.n636 VDDA.n635 0.0682083
R5935 VDDA.n642 VDDA.n568 0.0682083
R5936 VDDA.n650 VDDA.n564 0.0682083
R5937 VDDA.n652 VDDA.n651 0.0682083
R5938 VDDA.n660 VDDA.n659 0.0682083
R5939 VDDA.n666 VDDA.n556 0.0682083
R5940 VDDA.n674 VDDA.n552 0.0682083
R5941 VDDA.n676 VDDA.n675 0.0682083
R5942 VDDA.n1498 VDDA.n683 0.0682083
R5943 VDDA.n1388 VDDA.n1387 0.0682083
R5944 VDDA.n1396 VDDA.n1371 0.0682083
R5945 VDDA.n1406 VDDA.n1367 0.0682083
R5946 VDDA.n1408 VDDA.n1407 0.0682083
R5947 VDDA.n1418 VDDA.n1417 0.0682083
R5948 VDDA.n1426 VDDA.n1359 0.0682083
R5949 VDDA.n1436 VDDA.n1355 0.0682083
R5950 VDDA.n1438 VDDA.n1437 0.0682083
R5951 VDDA.n1448 VDDA.n1447 0.0682083
R5952 VDDA.n1456 VDDA.n1347 0.0682083
R5953 VDDA.n1466 VDDA.n1343 0.0682083
R5954 VDDA.n1468 VDDA.n1467 0.0682083
R5955 VDDA.n1478 VDDA.n1477 0.0682083
R5956 VDDA.n1486 VDDA.n1335 0.0682083
R5957 VDDA.n1495 VDDA.n1331 0.0682083
R5958 VDDA.n1223 VDDA.n1222 0.0682083
R5959 VDDA.n1231 VDDA.n1211 0.0682083
R5960 VDDA.n1241 VDDA.n1209 0.0682083
R5961 VDDA.n1243 VDDA.n1242 0.0682083
R5962 VDDA.n1253 VDDA.n1252 0.0682083
R5963 VDDA.n1261 VDDA.n1205 0.0682083
R5964 VDDA.n1271 VDDA.n1203 0.0682083
R5965 VDDA.n1273 VDDA.n1272 0.0682083
R5966 VDDA.n1283 VDDA.n1282 0.0682083
R5967 VDDA.n1291 VDDA.n1199 0.0682083
R5968 VDDA.n1301 VDDA.n1197 0.0682083
R5969 VDDA.n1303 VDDA.n1302 0.0682083
R5970 VDDA.n1313 VDDA.n1312 0.0682083
R5971 VDDA.n1321 VDDA.n1193 0.0682083
R5972 VDDA.n1330 VDDA.n684 0.0682083
R5973 VDDA.n90 VDDA.n89 0.0672139
R5974 VDDA.n3239 VDDA.n3238 0.0672139
R5975 VDDA.n3095 VDDA.n3093 0.0672139
R5976 VDDA.n2933 VDDA.n2932 0.0672139
R5977 VDDA.n427 VDDA.n426 0.0672139
R5978 VDDA.n1736 VDDA.n1734 0.0672139
R5979 VDDA.n1574 VDDA.n1573 0.0672139
R5980 VDDA.n594 VDDA.n593 0.0672139
R5981 VDDA.n1379 VDDA.n1378 0.0672139
R5982 VDDA.n1216 VDDA.n1214 0.0672139
R5983 VDDA.n2334 VDDA.n2153 0.0667303
R5984 VDDA.n2149 VDDA.n1924 0.0667303
R5985 VDDA.n352 VDDA.n209 0.0667303
R5986 VDDA.n2675 VDDA.n2534 0.0667303
R5987 VDDA.n2530 VDDA.n2338 0.0667303
R5988 VDDA.n99 VDDA.n98 0.063
R5989 VDDA.n108 VDDA.n76 0.063
R5990 VDDA.n123 VDDA.n122 0.063
R5991 VDDA.n132 VDDA.n64 0.063
R5992 VDDA.n147 VDDA.n146 0.063
R5993 VDDA.n156 VDDA.n52 0.063
R5994 VDDA.n171 VDDA.n170 0.063
R5995 VDDA.n3248 VDDA.n3231 0.063
R5996 VDDA.n3267 VDDA.n3266 0.063
R5997 VDDA.n3278 VDDA.n3219 0.063
R5998 VDDA.n3297 VDDA.n3296 0.063
R5999 VDDA.n3308 VDDA.n3207 0.063
R6000 VDDA.n3327 VDDA.n3326 0.063
R6001 VDDA.n3338 VDDA.n3195 0.063
R6002 VDDA.n3102 VDDA.n3088 0.063
R6003 VDDA.n3117 VDDA.n3116 0.063
R6004 VDDA.n3126 VDDA.n3076 0.063
R6005 VDDA.n3141 VDDA.n3140 0.063
R6006 VDDA.n3150 VDDA.n3064 0.063
R6007 VDDA.n3165 VDDA.n3164 0.063
R6008 VDDA.n3174 VDDA.n3052 0.063
R6009 VDDA.n2942 VDDA.n2941 0.063
R6010 VDDA.n2951 VDDA.n2919 0.063
R6011 VDDA.n2966 VDDA.n2965 0.063
R6012 VDDA.n2975 VDDA.n2907 0.063
R6013 VDDA.n2990 VDDA.n2989 0.063
R6014 VDDA.n2999 VDDA.n2895 0.063
R6015 VDDA.n3014 VDDA.n3013 0.063
R6016 VDDA.n436 VDDA.n435 0.063
R6017 VDDA.n445 VDDA.n413 0.063
R6018 VDDA.n460 VDDA.n459 0.063
R6019 VDDA.n469 VDDA.n401 0.063
R6020 VDDA.n484 VDDA.n483 0.063
R6021 VDDA.n493 VDDA.n389 0.063
R6022 VDDA.n508 VDDA.n507 0.063
R6023 VDDA.n1743 VDDA.n1729 0.063
R6024 VDDA.n1758 VDDA.n1757 0.063
R6025 VDDA.n1767 VDDA.n1717 0.063
R6026 VDDA.n1782 VDDA.n1781 0.063
R6027 VDDA.n1791 VDDA.n1705 0.063
R6028 VDDA.n1806 VDDA.n1805 0.063
R6029 VDDA.n1815 VDDA.n1693 0.063
R6030 VDDA.n1583 VDDA.n1582 0.063
R6031 VDDA.n1592 VDDA.n1560 0.063
R6032 VDDA.n1607 VDDA.n1606 0.063
R6033 VDDA.n1616 VDDA.n1548 0.063
R6034 VDDA.n1631 VDDA.n1630 0.063
R6035 VDDA.n1640 VDDA.n1536 0.063
R6036 VDDA.n1655 VDDA.n1654 0.063
R6037 VDDA.n603 VDDA.n602 0.063
R6038 VDDA.n612 VDDA.n580 0.063
R6039 VDDA.n627 VDDA.n626 0.063
R6040 VDDA.n636 VDDA.n568 0.063
R6041 VDDA.n651 VDDA.n650 0.063
R6042 VDDA.n660 VDDA.n556 0.063
R6043 VDDA.n675 VDDA.n674 0.063
R6044 VDDA.n1388 VDDA.n1371 0.063
R6045 VDDA.n1407 VDDA.n1406 0.063
R6046 VDDA.n1418 VDDA.n1359 0.063
R6047 VDDA.n1437 VDDA.n1436 0.063
R6048 VDDA.n1448 VDDA.n1347 0.063
R6049 VDDA.n1467 VDDA.n1466 0.063
R6050 VDDA.n1478 VDDA.n1335 0.063
R6051 VDDA.n1223 VDDA.n1211 0.063
R6052 VDDA.n1242 VDDA.n1241 0.063
R6053 VDDA.n1253 VDDA.n1205 0.063
R6054 VDDA.n1272 VDDA.n1271 0.063
R6055 VDDA.n1283 VDDA.n1199 0.063
R6056 VDDA.n1302 VDDA.n1301 0.063
R6057 VDDA.n1313 VDDA.n1193 0.063
R6058 VDDA.n2227 VDDA.n2226 0.0553333
R6059 VDDA.n2241 VDDA.n2240 0.0553333
R6060 VDDA.n2257 VDDA.n2256 0.0553333
R6061 VDDA.n2271 VDDA.n2270 0.0553333
R6062 VDDA.n2287 VDDA.n2286 0.0553333
R6063 VDDA.n2301 VDDA.n2300 0.0553333
R6064 VDDA.n2317 VDDA.n2316 0.0553333
R6065 VDDA.n2331 VDDA.n2330 0.0553333
R6066 VDDA.n2042 VDDA.n2041 0.0553333
R6067 VDDA.n2056 VDDA.n2055 0.0553333
R6068 VDDA.n2072 VDDA.n2071 0.0553333
R6069 VDDA.n2086 VDDA.n2085 0.0553333
R6070 VDDA.n2102 VDDA.n2101 0.0553333
R6071 VDDA.n2116 VDDA.n2115 0.0553333
R6072 VDDA.n2132 VDDA.n2131 0.0553333
R6073 VDDA.n2146 VDDA.n2145 0.0553333
R6074 VDDA.n245 VDDA.n244 0.0553333
R6075 VDDA.n259 VDDA.n258 0.0553333
R6076 VDDA.n275 VDDA.n274 0.0553333
R6077 VDDA.n289 VDDA.n288 0.0553333
R6078 VDDA.n305 VDDA.n304 0.0553333
R6079 VDDA.n319 VDDA.n318 0.0553333
R6080 VDDA.n335 VDDA.n334 0.0553333
R6081 VDDA.n349 VDDA.n348 0.0553333
R6082 VDDA.n2568 VDDA.n2567 0.0553333
R6083 VDDA.n2582 VDDA.n2581 0.0553333
R6084 VDDA.n2598 VDDA.n2597 0.0553333
R6085 VDDA.n2612 VDDA.n2611 0.0553333
R6086 VDDA.n2628 VDDA.n2627 0.0553333
R6087 VDDA.n2642 VDDA.n2641 0.0553333
R6088 VDDA.n2658 VDDA.n2657 0.0553333
R6089 VDDA.n2672 VDDA.n2671 0.0553333
R6090 VDDA.n2423 VDDA.n2422 0.0553333
R6091 VDDA.n2437 VDDA.n2436 0.0553333
R6092 VDDA.n2453 VDDA.n2452 0.0553333
R6093 VDDA.n2467 VDDA.n2466 0.0553333
R6094 VDDA.n2483 VDDA.n2482 0.0553333
R6095 VDDA.n2497 VDDA.n2496 0.0553333
R6096 VDDA.n2513 VDDA.n2512 0.0553333
R6097 VDDA.n2527 VDDA.n2526 0.0553333
R6098 VDDA.n87 VDDA.n86 0.0553333
R6099 VDDA.n104 VDDA.n103 0.0553333
R6100 VDDA.n75 VDDA.n74 0.0553333
R6101 VDDA.n128 VDDA.n127 0.0553333
R6102 VDDA.n63 VDDA.n62 0.0553333
R6103 VDDA.n152 VDDA.n151 0.0553333
R6104 VDDA.n51 VDDA.n50 0.0553333
R6105 VDDA.n176 VDDA.n175 0.0553333
R6106 VDDA.n3244 VDDA.n3242 0.0553333
R6107 VDDA.n3260 VDDA.n3229 0.0553333
R6108 VDDA.n3274 VDDA.n3272 0.0553333
R6109 VDDA.n3290 VDDA.n3217 0.0553333
R6110 VDDA.n3304 VDDA.n3302 0.0553333
R6111 VDDA.n3320 VDDA.n3205 0.0553333
R6112 VDDA.n3334 VDDA.n3332 0.0553333
R6113 VDDA.n3350 VDDA.n3193 0.0553333
R6114 VDDA.n3098 VDDA.n3097 0.0553333
R6115 VDDA.n3087 VDDA.n3086 0.0553333
R6116 VDDA.n3122 VDDA.n3121 0.0553333
R6117 VDDA.n3075 VDDA.n3074 0.0553333
R6118 VDDA.n3146 VDDA.n3145 0.0553333
R6119 VDDA.n3063 VDDA.n3062 0.0553333
R6120 VDDA.n3170 VDDA.n3169 0.0553333
R6121 VDDA.n3184 VDDA.n3050 0.0553333
R6122 VDDA.n2930 VDDA.n2929 0.0553333
R6123 VDDA.n2947 VDDA.n2946 0.0553333
R6124 VDDA.n2918 VDDA.n2917 0.0553333
R6125 VDDA.n2971 VDDA.n2970 0.0553333
R6126 VDDA.n2906 VDDA.n2905 0.0553333
R6127 VDDA.n2995 VDDA.n2994 0.0553333
R6128 VDDA.n2894 VDDA.n2893 0.0553333
R6129 VDDA.n3019 VDDA.n3018 0.0553333
R6130 VDDA.n424 VDDA.n423 0.0553333
R6131 VDDA.n441 VDDA.n440 0.0553333
R6132 VDDA.n412 VDDA.n411 0.0553333
R6133 VDDA.n465 VDDA.n464 0.0553333
R6134 VDDA.n400 VDDA.n399 0.0553333
R6135 VDDA.n489 VDDA.n488 0.0553333
R6136 VDDA.n388 VDDA.n387 0.0553333
R6137 VDDA.n513 VDDA.n512 0.0553333
R6138 VDDA.n1739 VDDA.n1738 0.0553333
R6139 VDDA.n1728 VDDA.n1727 0.0553333
R6140 VDDA.n1763 VDDA.n1762 0.0553333
R6141 VDDA.n1716 VDDA.n1715 0.0553333
R6142 VDDA.n1787 VDDA.n1786 0.0553333
R6143 VDDA.n1704 VDDA.n1703 0.0553333
R6144 VDDA.n1811 VDDA.n1810 0.0553333
R6145 VDDA.n1825 VDDA.n1691 0.0553333
R6146 VDDA.n1571 VDDA.n1570 0.0553333
R6147 VDDA.n1588 VDDA.n1587 0.0553333
R6148 VDDA.n1559 VDDA.n1558 0.0553333
R6149 VDDA.n1612 VDDA.n1611 0.0553333
R6150 VDDA.n1547 VDDA.n1546 0.0553333
R6151 VDDA.n1636 VDDA.n1635 0.0553333
R6152 VDDA.n1535 VDDA.n1534 0.0553333
R6153 VDDA.n1660 VDDA.n1659 0.0553333
R6154 VDDA.n591 VDDA.n590 0.0553333
R6155 VDDA.n608 VDDA.n607 0.0553333
R6156 VDDA.n579 VDDA.n578 0.0553333
R6157 VDDA.n632 VDDA.n631 0.0553333
R6158 VDDA.n567 VDDA.n566 0.0553333
R6159 VDDA.n656 VDDA.n655 0.0553333
R6160 VDDA.n555 VDDA.n554 0.0553333
R6161 VDDA.n680 VDDA.n679 0.0553333
R6162 VDDA.n1384 VDDA.n1382 0.0553333
R6163 VDDA.n1400 VDDA.n1369 0.0553333
R6164 VDDA.n1414 VDDA.n1412 0.0553333
R6165 VDDA.n1430 VDDA.n1357 0.0553333
R6166 VDDA.n1444 VDDA.n1442 0.0553333
R6167 VDDA.n1460 VDDA.n1345 0.0553333
R6168 VDDA.n1474 VDDA.n1472 0.0553333
R6169 VDDA.n1490 VDDA.n1333 0.0553333
R6170 VDDA.n1219 VDDA.n1218 0.0553333
R6171 VDDA.n1235 VDDA.n1234 0.0553333
R6172 VDDA.n1249 VDDA.n1248 0.0553333
R6173 VDDA.n1265 VDDA.n1264 0.0553333
R6174 VDDA.n1279 VDDA.n1278 0.0553333
R6175 VDDA.n1295 VDDA.n1294 0.0553333
R6176 VDDA.n1309 VDDA.n1308 0.0553333
R6177 VDDA.n1325 VDDA.n1191 0.0553333
R6178 VDDA.n2221 VDDA.n1875 0.0514167
R6179 VDDA.n2231 VDDA.n2230 0.0514167
R6180 VDDA.n2237 VDDA.n2236 0.0514167
R6181 VDDA.n2247 VDDA.n2246 0.0514167
R6182 VDDA.n2251 VDDA.n2250 0.0514167
R6183 VDDA.n2261 VDDA.n2260 0.0514167
R6184 VDDA.n2267 VDDA.n2266 0.0514167
R6185 VDDA.n2277 VDDA.n2276 0.0514167
R6186 VDDA.n2281 VDDA.n2280 0.0514167
R6187 VDDA.n2291 VDDA.n2290 0.0514167
R6188 VDDA.n2297 VDDA.n2296 0.0514167
R6189 VDDA.n2307 VDDA.n2306 0.0514167
R6190 VDDA.n2311 VDDA.n2310 0.0514167
R6191 VDDA.n2321 VDDA.n2320 0.0514167
R6192 VDDA.n2327 VDDA.n2326 0.0514167
R6193 VDDA.n2335 VDDA.n2152 0.0514167
R6194 VDDA.n2036 VDDA.n1899 0.0514167
R6195 VDDA.n2046 VDDA.n2045 0.0514167
R6196 VDDA.n2052 VDDA.n2051 0.0514167
R6197 VDDA.n2062 VDDA.n2061 0.0514167
R6198 VDDA.n2066 VDDA.n2065 0.0514167
R6199 VDDA.n2076 VDDA.n2075 0.0514167
R6200 VDDA.n2082 VDDA.n2081 0.0514167
R6201 VDDA.n2092 VDDA.n2091 0.0514167
R6202 VDDA.n2096 VDDA.n2095 0.0514167
R6203 VDDA.n2106 VDDA.n2105 0.0514167
R6204 VDDA.n2112 VDDA.n2111 0.0514167
R6205 VDDA.n2122 VDDA.n2121 0.0514167
R6206 VDDA.n2126 VDDA.n2125 0.0514167
R6207 VDDA.n2136 VDDA.n2135 0.0514167
R6208 VDDA.n2142 VDDA.n2141 0.0514167
R6209 VDDA.n2150 VDDA.n1923 0.0514167
R6210 VDDA.n239 VDDA.n184 0.0514167
R6211 VDDA.n249 VDDA.n248 0.0514167
R6212 VDDA.n255 VDDA.n254 0.0514167
R6213 VDDA.n265 VDDA.n264 0.0514167
R6214 VDDA.n269 VDDA.n268 0.0514167
R6215 VDDA.n279 VDDA.n278 0.0514167
R6216 VDDA.n285 VDDA.n284 0.0514167
R6217 VDDA.n295 VDDA.n294 0.0514167
R6218 VDDA.n299 VDDA.n298 0.0514167
R6219 VDDA.n309 VDDA.n308 0.0514167
R6220 VDDA.n315 VDDA.n314 0.0514167
R6221 VDDA.n325 VDDA.n324 0.0514167
R6222 VDDA.n329 VDDA.n328 0.0514167
R6223 VDDA.n339 VDDA.n338 0.0514167
R6224 VDDA.n345 VDDA.n344 0.0514167
R6225 VDDA.n353 VDDA.n208 0.0514167
R6226 VDDA.n2562 VDDA.n1827 0.0514167
R6227 VDDA.n2572 VDDA.n2571 0.0514167
R6228 VDDA.n2578 VDDA.n2577 0.0514167
R6229 VDDA.n2588 VDDA.n2587 0.0514167
R6230 VDDA.n2592 VDDA.n2591 0.0514167
R6231 VDDA.n2602 VDDA.n2601 0.0514167
R6232 VDDA.n2608 VDDA.n2607 0.0514167
R6233 VDDA.n2618 VDDA.n2617 0.0514167
R6234 VDDA.n2622 VDDA.n2621 0.0514167
R6235 VDDA.n2632 VDDA.n2631 0.0514167
R6236 VDDA.n2638 VDDA.n2637 0.0514167
R6237 VDDA.n2648 VDDA.n2647 0.0514167
R6238 VDDA.n2652 VDDA.n2651 0.0514167
R6239 VDDA.n2662 VDDA.n2661 0.0514167
R6240 VDDA.n2668 VDDA.n2667 0.0514167
R6241 VDDA.n2676 VDDA.n2533 0.0514167
R6242 VDDA.n2417 VDDA.n1851 0.0514167
R6243 VDDA.n2427 VDDA.n2426 0.0514167
R6244 VDDA.n2433 VDDA.n2432 0.0514167
R6245 VDDA.n2443 VDDA.n2442 0.0514167
R6246 VDDA.n2447 VDDA.n2446 0.0514167
R6247 VDDA.n2457 VDDA.n2456 0.0514167
R6248 VDDA.n2463 VDDA.n2462 0.0514167
R6249 VDDA.n2473 VDDA.n2472 0.0514167
R6250 VDDA.n2477 VDDA.n2476 0.0514167
R6251 VDDA.n2487 VDDA.n2486 0.0514167
R6252 VDDA.n2493 VDDA.n2492 0.0514167
R6253 VDDA.n2503 VDDA.n2502 0.0514167
R6254 VDDA.n2507 VDDA.n2506 0.0514167
R6255 VDDA.n2517 VDDA.n2516 0.0514167
R6256 VDDA.n2523 VDDA.n2522 0.0514167
R6257 VDDA.n2531 VDDA.n2337 0.0514167
R6258 VDDA.n88 VDDA.n18 0.0514167
R6259 VDDA.n96 VDDA.n95 0.0514167
R6260 VDDA.n83 VDDA.n82 0.0514167
R6261 VDDA.n79 VDDA.n78 0.0514167
R6262 VDDA.n112 VDDA.n111 0.0514167
R6263 VDDA.n120 VDDA.n119 0.0514167
R6264 VDDA.n71 VDDA.n70 0.0514167
R6265 VDDA.n67 VDDA.n66 0.0514167
R6266 VDDA.n136 VDDA.n135 0.0514167
R6267 VDDA.n144 VDDA.n143 0.0514167
R6268 VDDA.n59 VDDA.n58 0.0514167
R6269 VDDA.n55 VDDA.n54 0.0514167
R6270 VDDA.n160 VDDA.n159 0.0514167
R6271 VDDA.n168 VDDA.n167 0.0514167
R6272 VDDA.n47 VDDA.n46 0.0514167
R6273 VDDA.n3359 VDDA.n42 0.0514167
R6274 VDDA.n3240 VDDA.n3237 0.0514167
R6275 VDDA.n3250 VDDA.n3233 0.0514167
R6276 VDDA.n3254 VDDA.n3252 0.0514167
R6277 VDDA.n3264 VDDA.n3262 0.0514167
R6278 VDDA.n3270 VDDA.n3225 0.0514167
R6279 VDDA.n3280 VDDA.n3221 0.0514167
R6280 VDDA.n3284 VDDA.n3282 0.0514167
R6281 VDDA.n3294 VDDA.n3292 0.0514167
R6282 VDDA.n3300 VDDA.n3213 0.0514167
R6283 VDDA.n3310 VDDA.n3209 0.0514167
R6284 VDDA.n3314 VDDA.n3312 0.0514167
R6285 VDDA.n3324 VDDA.n3322 0.0514167
R6286 VDDA.n3330 VDDA.n3201 0.0514167
R6287 VDDA.n3340 VDDA.n3197 0.0514167
R6288 VDDA.n3344 VDDA.n3342 0.0514167
R6289 VDDA.n3353 VDDA.n3352 0.0514167
R6290 VDDA.n3094 VDDA.n3027 0.0514167
R6291 VDDA.n3091 VDDA.n3090 0.0514167
R6292 VDDA.n3106 VDDA.n3105 0.0514167
R6293 VDDA.n3114 VDDA.n3113 0.0514167
R6294 VDDA.n3083 VDDA.n3082 0.0514167
R6295 VDDA.n3079 VDDA.n3078 0.0514167
R6296 VDDA.n3130 VDDA.n3129 0.0514167
R6297 VDDA.n3138 VDDA.n3137 0.0514167
R6298 VDDA.n3071 VDDA.n3070 0.0514167
R6299 VDDA.n3067 VDDA.n3066 0.0514167
R6300 VDDA.n3154 VDDA.n3153 0.0514167
R6301 VDDA.n3162 VDDA.n3161 0.0514167
R6302 VDDA.n3059 VDDA.n3058 0.0514167
R6303 VDDA.n3055 VDDA.n3054 0.0514167
R6304 VDDA.n3178 VDDA.n3177 0.0514167
R6305 VDDA.n3187 VDDA.n183 0.0514167
R6306 VDDA.n2931 VDDA.n2861 0.0514167
R6307 VDDA.n2939 VDDA.n2938 0.0514167
R6308 VDDA.n2926 VDDA.n2925 0.0514167
R6309 VDDA.n2922 VDDA.n2921 0.0514167
R6310 VDDA.n2955 VDDA.n2954 0.0514167
R6311 VDDA.n2963 VDDA.n2962 0.0514167
R6312 VDDA.n2914 VDDA.n2913 0.0514167
R6313 VDDA.n2910 VDDA.n2909 0.0514167
R6314 VDDA.n2979 VDDA.n2978 0.0514167
R6315 VDDA.n2987 VDDA.n2986 0.0514167
R6316 VDDA.n2902 VDDA.n2901 0.0514167
R6317 VDDA.n2898 VDDA.n2897 0.0514167
R6318 VDDA.n3003 VDDA.n3002 0.0514167
R6319 VDDA.n3011 VDDA.n3010 0.0514167
R6320 VDDA.n2890 VDDA.n2889 0.0514167
R6321 VDDA.n3025 VDDA.n2885 0.0514167
R6322 VDDA.n425 VDDA.n355 0.0514167
R6323 VDDA.n433 VDDA.n432 0.0514167
R6324 VDDA.n420 VDDA.n419 0.0514167
R6325 VDDA.n416 VDDA.n415 0.0514167
R6326 VDDA.n449 VDDA.n448 0.0514167
R6327 VDDA.n457 VDDA.n456 0.0514167
R6328 VDDA.n408 VDDA.n407 0.0514167
R6329 VDDA.n404 VDDA.n403 0.0514167
R6330 VDDA.n473 VDDA.n472 0.0514167
R6331 VDDA.n481 VDDA.n480 0.0514167
R6332 VDDA.n396 VDDA.n395 0.0514167
R6333 VDDA.n392 VDDA.n391 0.0514167
R6334 VDDA.n497 VDDA.n496 0.0514167
R6335 VDDA.n505 VDDA.n504 0.0514167
R6336 VDDA.n384 VDDA.n383 0.0514167
R6337 VDDA.n2859 VDDA.n379 0.0514167
R6338 VDDA.n1735 VDDA.n1668 0.0514167
R6339 VDDA.n1732 VDDA.n1731 0.0514167
R6340 VDDA.n1747 VDDA.n1746 0.0514167
R6341 VDDA.n1755 VDDA.n1754 0.0514167
R6342 VDDA.n1724 VDDA.n1723 0.0514167
R6343 VDDA.n1720 VDDA.n1719 0.0514167
R6344 VDDA.n1771 VDDA.n1770 0.0514167
R6345 VDDA.n1779 VDDA.n1778 0.0514167
R6346 VDDA.n1712 VDDA.n1711 0.0514167
R6347 VDDA.n1708 VDDA.n1707 0.0514167
R6348 VDDA.n1795 VDDA.n1794 0.0514167
R6349 VDDA.n1803 VDDA.n1802 0.0514167
R6350 VDDA.n1700 VDDA.n1699 0.0514167
R6351 VDDA.n1696 VDDA.n1695 0.0514167
R6352 VDDA.n1819 VDDA.n1818 0.0514167
R6353 VDDA.n2679 VDDA.n520 0.0514167
R6354 VDDA.n1572 VDDA.n1502 0.0514167
R6355 VDDA.n1580 VDDA.n1579 0.0514167
R6356 VDDA.n1567 VDDA.n1566 0.0514167
R6357 VDDA.n1563 VDDA.n1562 0.0514167
R6358 VDDA.n1596 VDDA.n1595 0.0514167
R6359 VDDA.n1604 VDDA.n1603 0.0514167
R6360 VDDA.n1555 VDDA.n1554 0.0514167
R6361 VDDA.n1551 VDDA.n1550 0.0514167
R6362 VDDA.n1620 VDDA.n1619 0.0514167
R6363 VDDA.n1628 VDDA.n1627 0.0514167
R6364 VDDA.n1543 VDDA.n1542 0.0514167
R6365 VDDA.n1539 VDDA.n1538 0.0514167
R6366 VDDA.n1644 VDDA.n1643 0.0514167
R6367 VDDA.n1652 VDDA.n1651 0.0514167
R6368 VDDA.n1531 VDDA.n1530 0.0514167
R6369 VDDA.n1666 VDDA.n1526 0.0514167
R6370 VDDA.n592 VDDA.n522 0.0514167
R6371 VDDA.n600 VDDA.n599 0.0514167
R6372 VDDA.n587 VDDA.n586 0.0514167
R6373 VDDA.n583 VDDA.n582 0.0514167
R6374 VDDA.n616 VDDA.n615 0.0514167
R6375 VDDA.n624 VDDA.n623 0.0514167
R6376 VDDA.n575 VDDA.n574 0.0514167
R6377 VDDA.n571 VDDA.n570 0.0514167
R6378 VDDA.n640 VDDA.n639 0.0514167
R6379 VDDA.n648 VDDA.n647 0.0514167
R6380 VDDA.n563 VDDA.n562 0.0514167
R6381 VDDA.n559 VDDA.n558 0.0514167
R6382 VDDA.n664 VDDA.n663 0.0514167
R6383 VDDA.n672 VDDA.n671 0.0514167
R6384 VDDA.n551 VDDA.n550 0.0514167
R6385 VDDA.n1500 VDDA.n546 0.0514167
R6386 VDDA.n1380 VDDA.n1377 0.0514167
R6387 VDDA.n1390 VDDA.n1373 0.0514167
R6388 VDDA.n1394 VDDA.n1392 0.0514167
R6389 VDDA.n1404 VDDA.n1402 0.0514167
R6390 VDDA.n1410 VDDA.n1365 0.0514167
R6391 VDDA.n1420 VDDA.n1361 0.0514167
R6392 VDDA.n1424 VDDA.n1422 0.0514167
R6393 VDDA.n1434 VDDA.n1432 0.0514167
R6394 VDDA.n1440 VDDA.n1353 0.0514167
R6395 VDDA.n1450 VDDA.n1349 0.0514167
R6396 VDDA.n1454 VDDA.n1452 0.0514167
R6397 VDDA.n1464 VDDA.n1462 0.0514167
R6398 VDDA.n1470 VDDA.n1341 0.0514167
R6399 VDDA.n1480 VDDA.n1337 0.0514167
R6400 VDDA.n1484 VDDA.n1482 0.0514167
R6401 VDDA.n1493 VDDA.n1492 0.0514167
R6402 VDDA.n1215 VDDA.n1168 0.0514167
R6403 VDDA.n1225 VDDA.n1224 0.0514167
R6404 VDDA.n1229 VDDA.n1228 0.0514167
R6405 VDDA.n1239 VDDA.n1238 0.0514167
R6406 VDDA.n1245 VDDA.n1244 0.0514167
R6407 VDDA.n1255 VDDA.n1254 0.0514167
R6408 VDDA.n1259 VDDA.n1258 0.0514167
R6409 VDDA.n1269 VDDA.n1268 0.0514167
R6410 VDDA.n1275 VDDA.n1274 0.0514167
R6411 VDDA.n1285 VDDA.n1284 0.0514167
R6412 VDDA.n1289 VDDA.n1288 0.0514167
R6413 VDDA.n1299 VDDA.n1298 0.0514167
R6414 VDDA.n1305 VDDA.n1304 0.0514167
R6415 VDDA.n1315 VDDA.n1314 0.0514167
R6416 VDDA.n1319 VDDA.n1318 0.0514167
R6417 VDDA.n1328 VDDA.n686 0.0514167
R6418 VDDA.n2336 VDDA.n2151 0.0358969
R6419 VDDA.n3466 VDDA.n3360 0.0297281
R6420 VDDA.n2226 VDDA.n1876 0.028198
R6421 VDDA.n2230 VDDA.n1877 0.028198
R6422 VDDA.n2240 VDDA.n1879 0.028198
R6423 VDDA.n2246 VDDA.n1880 0.028198
R6424 VDDA.n2256 VDDA.n1882 0.028198
R6425 VDDA.n2260 VDDA.n1883 0.028198
R6426 VDDA.n2270 VDDA.n1885 0.028198
R6427 VDDA.n2276 VDDA.n1886 0.028198
R6428 VDDA.n2286 VDDA.n1888 0.028198
R6429 VDDA.n2290 VDDA.n1889 0.028198
R6430 VDDA.n2300 VDDA.n1891 0.028198
R6431 VDDA.n2306 VDDA.n1892 0.028198
R6432 VDDA.n2316 VDDA.n1894 0.028198
R6433 VDDA.n2320 VDDA.n1895 0.028198
R6434 VDDA.n2330 VDDA.n1897 0.028198
R6435 VDDA.n2152 VDDA.n1898 0.028198
R6436 VDDA.n2041 VDDA.n1900 0.028198
R6437 VDDA.n2045 VDDA.n1901 0.028198
R6438 VDDA.n2055 VDDA.n1903 0.028198
R6439 VDDA.n2061 VDDA.n1904 0.028198
R6440 VDDA.n2071 VDDA.n1906 0.028198
R6441 VDDA.n2075 VDDA.n1907 0.028198
R6442 VDDA.n2085 VDDA.n1909 0.028198
R6443 VDDA.n2091 VDDA.n1910 0.028198
R6444 VDDA.n2101 VDDA.n1912 0.028198
R6445 VDDA.n2105 VDDA.n1913 0.028198
R6446 VDDA.n2115 VDDA.n1915 0.028198
R6447 VDDA.n2121 VDDA.n1916 0.028198
R6448 VDDA.n2131 VDDA.n1918 0.028198
R6449 VDDA.n2135 VDDA.n1919 0.028198
R6450 VDDA.n2145 VDDA.n1921 0.028198
R6451 VDDA.n1923 VDDA.n1922 0.028198
R6452 VDDA.n244 VDDA.n185 0.028198
R6453 VDDA.n248 VDDA.n186 0.028198
R6454 VDDA.n258 VDDA.n188 0.028198
R6455 VDDA.n264 VDDA.n189 0.028198
R6456 VDDA.n274 VDDA.n191 0.028198
R6457 VDDA.n278 VDDA.n192 0.028198
R6458 VDDA.n288 VDDA.n194 0.028198
R6459 VDDA.n294 VDDA.n195 0.028198
R6460 VDDA.n304 VDDA.n197 0.028198
R6461 VDDA.n308 VDDA.n198 0.028198
R6462 VDDA.n318 VDDA.n200 0.028198
R6463 VDDA.n324 VDDA.n201 0.028198
R6464 VDDA.n334 VDDA.n203 0.028198
R6465 VDDA.n338 VDDA.n204 0.028198
R6466 VDDA.n348 VDDA.n206 0.028198
R6467 VDDA.n208 VDDA.n207 0.028198
R6468 VDDA.n2567 VDDA.n1828 0.028198
R6469 VDDA.n2571 VDDA.n1829 0.028198
R6470 VDDA.n2581 VDDA.n1831 0.028198
R6471 VDDA.n2587 VDDA.n1832 0.028198
R6472 VDDA.n2597 VDDA.n1834 0.028198
R6473 VDDA.n2601 VDDA.n1835 0.028198
R6474 VDDA.n2611 VDDA.n1837 0.028198
R6475 VDDA.n2617 VDDA.n1838 0.028198
R6476 VDDA.n2627 VDDA.n1840 0.028198
R6477 VDDA.n2631 VDDA.n1841 0.028198
R6478 VDDA.n2641 VDDA.n1843 0.028198
R6479 VDDA.n2647 VDDA.n1844 0.028198
R6480 VDDA.n2657 VDDA.n1846 0.028198
R6481 VDDA.n2661 VDDA.n1847 0.028198
R6482 VDDA.n2671 VDDA.n1849 0.028198
R6483 VDDA.n2533 VDDA.n1850 0.028198
R6484 VDDA.n2422 VDDA.n1852 0.028198
R6485 VDDA.n2426 VDDA.n1853 0.028198
R6486 VDDA.n2436 VDDA.n1855 0.028198
R6487 VDDA.n2442 VDDA.n1856 0.028198
R6488 VDDA.n2452 VDDA.n1858 0.028198
R6489 VDDA.n2456 VDDA.n1859 0.028198
R6490 VDDA.n2466 VDDA.n1861 0.028198
R6491 VDDA.n2472 VDDA.n1862 0.028198
R6492 VDDA.n2482 VDDA.n1864 0.028198
R6493 VDDA.n2486 VDDA.n1865 0.028198
R6494 VDDA.n2496 VDDA.n1867 0.028198
R6495 VDDA.n2502 VDDA.n1868 0.028198
R6496 VDDA.n2512 VDDA.n1870 0.028198
R6497 VDDA.n2516 VDDA.n1871 0.028198
R6498 VDDA.n2526 VDDA.n1873 0.028198
R6499 VDDA.n2337 VDDA.n1874 0.028198
R6500 VDDA.n86 VDDA.n19 0.028198
R6501 VDDA.n95 VDDA.n20 0.028198
R6502 VDDA.n103 VDDA.n22 0.028198
R6503 VDDA.n78 VDDA.n23 0.028198
R6504 VDDA.n74 VDDA.n25 0.028198
R6505 VDDA.n119 VDDA.n26 0.028198
R6506 VDDA.n127 VDDA.n28 0.028198
R6507 VDDA.n66 VDDA.n29 0.028198
R6508 VDDA.n62 VDDA.n31 0.028198
R6509 VDDA.n143 VDDA.n32 0.028198
R6510 VDDA.n151 VDDA.n34 0.028198
R6511 VDDA.n54 VDDA.n35 0.028198
R6512 VDDA.n50 VDDA.n37 0.028198
R6513 VDDA.n167 VDDA.n38 0.028198
R6514 VDDA.n175 VDDA.n40 0.028198
R6515 VDDA.n42 VDDA.n41 0.028198
R6516 VDDA.n3242 VDDA.n3241 0.028198
R6517 VDDA.n3243 VDDA.n3233 0.028198
R6518 VDDA.n3253 VDDA.n3229 0.028198
R6519 VDDA.n3262 VDDA.n3261 0.028198
R6520 VDDA.n3272 VDDA.n3271 0.028198
R6521 VDDA.n3273 VDDA.n3221 0.028198
R6522 VDDA.n3283 VDDA.n3217 0.028198
R6523 VDDA.n3292 VDDA.n3291 0.028198
R6524 VDDA.n3302 VDDA.n3301 0.028198
R6525 VDDA.n3303 VDDA.n3209 0.028198
R6526 VDDA.n3313 VDDA.n3205 0.028198
R6527 VDDA.n3322 VDDA.n3321 0.028198
R6528 VDDA.n3332 VDDA.n3331 0.028198
R6529 VDDA.n3333 VDDA.n3197 0.028198
R6530 VDDA.n3343 VDDA.n3193 0.028198
R6531 VDDA.n3352 VDDA.n3351 0.028198
R6532 VDDA.n3097 VDDA.n3028 0.028198
R6533 VDDA.n3090 VDDA.n3029 0.028198
R6534 VDDA.n3086 VDDA.n3031 0.028198
R6535 VDDA.n3113 VDDA.n3032 0.028198
R6536 VDDA.n3121 VDDA.n3034 0.028198
R6537 VDDA.n3078 VDDA.n3035 0.028198
R6538 VDDA.n3074 VDDA.n3037 0.028198
R6539 VDDA.n3137 VDDA.n3038 0.028198
R6540 VDDA.n3145 VDDA.n3040 0.028198
R6541 VDDA.n3066 VDDA.n3041 0.028198
R6542 VDDA.n3062 VDDA.n3043 0.028198
R6543 VDDA.n3161 VDDA.n3044 0.028198
R6544 VDDA.n3169 VDDA.n3046 0.028198
R6545 VDDA.n3054 VDDA.n3047 0.028198
R6546 VDDA.n3050 VDDA.n3049 0.028198
R6547 VDDA.n3185 VDDA.n183 0.028198
R6548 VDDA.n2929 VDDA.n2862 0.028198
R6549 VDDA.n2938 VDDA.n2863 0.028198
R6550 VDDA.n2946 VDDA.n2865 0.028198
R6551 VDDA.n2921 VDDA.n2866 0.028198
R6552 VDDA.n2917 VDDA.n2868 0.028198
R6553 VDDA.n2962 VDDA.n2869 0.028198
R6554 VDDA.n2970 VDDA.n2871 0.028198
R6555 VDDA.n2909 VDDA.n2872 0.028198
R6556 VDDA.n2905 VDDA.n2874 0.028198
R6557 VDDA.n2986 VDDA.n2875 0.028198
R6558 VDDA.n2994 VDDA.n2877 0.028198
R6559 VDDA.n2897 VDDA.n2878 0.028198
R6560 VDDA.n2893 VDDA.n2880 0.028198
R6561 VDDA.n3010 VDDA.n2881 0.028198
R6562 VDDA.n3018 VDDA.n2883 0.028198
R6563 VDDA.n2885 VDDA.n2884 0.028198
R6564 VDDA.n423 VDDA.n356 0.028198
R6565 VDDA.n432 VDDA.n357 0.028198
R6566 VDDA.n440 VDDA.n359 0.028198
R6567 VDDA.n415 VDDA.n360 0.028198
R6568 VDDA.n411 VDDA.n362 0.028198
R6569 VDDA.n456 VDDA.n363 0.028198
R6570 VDDA.n464 VDDA.n365 0.028198
R6571 VDDA.n403 VDDA.n366 0.028198
R6572 VDDA.n399 VDDA.n368 0.028198
R6573 VDDA.n480 VDDA.n369 0.028198
R6574 VDDA.n488 VDDA.n371 0.028198
R6575 VDDA.n391 VDDA.n372 0.028198
R6576 VDDA.n387 VDDA.n374 0.028198
R6577 VDDA.n504 VDDA.n375 0.028198
R6578 VDDA.n512 VDDA.n377 0.028198
R6579 VDDA.n379 VDDA.n378 0.028198
R6580 VDDA.n1738 VDDA.n1669 0.028198
R6581 VDDA.n1731 VDDA.n1670 0.028198
R6582 VDDA.n1727 VDDA.n1672 0.028198
R6583 VDDA.n1754 VDDA.n1673 0.028198
R6584 VDDA.n1762 VDDA.n1675 0.028198
R6585 VDDA.n1719 VDDA.n1676 0.028198
R6586 VDDA.n1715 VDDA.n1678 0.028198
R6587 VDDA.n1778 VDDA.n1679 0.028198
R6588 VDDA.n1786 VDDA.n1681 0.028198
R6589 VDDA.n1707 VDDA.n1682 0.028198
R6590 VDDA.n1703 VDDA.n1684 0.028198
R6591 VDDA.n1802 VDDA.n1685 0.028198
R6592 VDDA.n1810 VDDA.n1687 0.028198
R6593 VDDA.n1695 VDDA.n1688 0.028198
R6594 VDDA.n1691 VDDA.n1690 0.028198
R6595 VDDA.n1826 VDDA.n520 0.028198
R6596 VDDA.n1570 VDDA.n1503 0.028198
R6597 VDDA.n1579 VDDA.n1504 0.028198
R6598 VDDA.n1587 VDDA.n1506 0.028198
R6599 VDDA.n1562 VDDA.n1507 0.028198
R6600 VDDA.n1558 VDDA.n1509 0.028198
R6601 VDDA.n1603 VDDA.n1510 0.028198
R6602 VDDA.n1611 VDDA.n1512 0.028198
R6603 VDDA.n1550 VDDA.n1513 0.028198
R6604 VDDA.n1546 VDDA.n1515 0.028198
R6605 VDDA.n1627 VDDA.n1516 0.028198
R6606 VDDA.n1635 VDDA.n1518 0.028198
R6607 VDDA.n1538 VDDA.n1519 0.028198
R6608 VDDA.n1534 VDDA.n1521 0.028198
R6609 VDDA.n1651 VDDA.n1522 0.028198
R6610 VDDA.n1659 VDDA.n1524 0.028198
R6611 VDDA.n1526 VDDA.n1525 0.028198
R6612 VDDA.n590 VDDA.n523 0.028198
R6613 VDDA.n599 VDDA.n524 0.028198
R6614 VDDA.n607 VDDA.n526 0.028198
R6615 VDDA.n582 VDDA.n527 0.028198
R6616 VDDA.n578 VDDA.n529 0.028198
R6617 VDDA.n623 VDDA.n530 0.028198
R6618 VDDA.n631 VDDA.n532 0.028198
R6619 VDDA.n570 VDDA.n533 0.028198
R6620 VDDA.n566 VDDA.n535 0.028198
R6621 VDDA.n647 VDDA.n536 0.028198
R6622 VDDA.n655 VDDA.n538 0.028198
R6623 VDDA.n558 VDDA.n539 0.028198
R6624 VDDA.n554 VDDA.n541 0.028198
R6625 VDDA.n671 VDDA.n542 0.028198
R6626 VDDA.n679 VDDA.n544 0.028198
R6627 VDDA.n546 VDDA.n545 0.028198
R6628 VDDA.n1382 VDDA.n1381 0.028198
R6629 VDDA.n1383 VDDA.n1373 0.028198
R6630 VDDA.n1393 VDDA.n1369 0.028198
R6631 VDDA.n1402 VDDA.n1401 0.028198
R6632 VDDA.n1412 VDDA.n1411 0.028198
R6633 VDDA.n1413 VDDA.n1361 0.028198
R6634 VDDA.n1423 VDDA.n1357 0.028198
R6635 VDDA.n1432 VDDA.n1431 0.028198
R6636 VDDA.n1442 VDDA.n1441 0.028198
R6637 VDDA.n1443 VDDA.n1349 0.028198
R6638 VDDA.n1453 VDDA.n1345 0.028198
R6639 VDDA.n1462 VDDA.n1461 0.028198
R6640 VDDA.n1472 VDDA.n1471 0.028198
R6641 VDDA.n1473 VDDA.n1337 0.028198
R6642 VDDA.n1483 VDDA.n1333 0.028198
R6643 VDDA.n1492 VDDA.n1491 0.028198
R6644 VDDA.n1218 VDDA.n1169 0.028198
R6645 VDDA.n1224 VDDA.n1170 0.028198
R6646 VDDA.n1234 VDDA.n1172 0.028198
R6647 VDDA.n1238 VDDA.n1173 0.028198
R6648 VDDA.n1248 VDDA.n1175 0.028198
R6649 VDDA.n1254 VDDA.n1176 0.028198
R6650 VDDA.n1264 VDDA.n1178 0.028198
R6651 VDDA.n1268 VDDA.n1179 0.028198
R6652 VDDA.n1278 VDDA.n1181 0.028198
R6653 VDDA.n1284 VDDA.n1182 0.028198
R6654 VDDA.n1294 VDDA.n1184 0.028198
R6655 VDDA.n1298 VDDA.n1185 0.028198
R6656 VDDA.n1308 VDDA.n1187 0.028198
R6657 VDDA.n1314 VDDA.n1188 0.028198
R6658 VDDA.n1191 VDDA.n1190 0.028198
R6659 VDDA.n1326 VDDA.n686 0.028198
R6660 VDDA.n1326 VDDA.n1325 0.028198
R6661 VDDA.n1319 VDDA.n1190 0.028198
R6662 VDDA.n1309 VDDA.n1188 0.028198
R6663 VDDA.n1305 VDDA.n1187 0.028198
R6664 VDDA.n1295 VDDA.n1185 0.028198
R6665 VDDA.n1289 VDDA.n1184 0.028198
R6666 VDDA.n1279 VDDA.n1182 0.028198
R6667 VDDA.n1275 VDDA.n1181 0.028198
R6668 VDDA.n1265 VDDA.n1179 0.028198
R6669 VDDA.n1259 VDDA.n1178 0.028198
R6670 VDDA.n1249 VDDA.n1176 0.028198
R6671 VDDA.n1245 VDDA.n1175 0.028198
R6672 VDDA.n1235 VDDA.n1173 0.028198
R6673 VDDA.n1229 VDDA.n1172 0.028198
R6674 VDDA.n1219 VDDA.n1170 0.028198
R6675 VDDA.n1215 VDDA.n1169 0.028198
R6676 VDDA.n1491 VDDA.n1490 0.028198
R6677 VDDA.n1484 VDDA.n1483 0.028198
R6678 VDDA.n1474 VDDA.n1473 0.028198
R6679 VDDA.n1471 VDDA.n1470 0.028198
R6680 VDDA.n1461 VDDA.n1460 0.028198
R6681 VDDA.n1454 VDDA.n1453 0.028198
R6682 VDDA.n1444 VDDA.n1443 0.028198
R6683 VDDA.n1441 VDDA.n1440 0.028198
R6684 VDDA.n1431 VDDA.n1430 0.028198
R6685 VDDA.n1424 VDDA.n1423 0.028198
R6686 VDDA.n1414 VDDA.n1413 0.028198
R6687 VDDA.n1411 VDDA.n1410 0.028198
R6688 VDDA.n1401 VDDA.n1400 0.028198
R6689 VDDA.n1394 VDDA.n1393 0.028198
R6690 VDDA.n1384 VDDA.n1383 0.028198
R6691 VDDA.n1381 VDDA.n1380 0.028198
R6692 VDDA.n680 VDDA.n545 0.028198
R6693 VDDA.n551 VDDA.n544 0.028198
R6694 VDDA.n555 VDDA.n542 0.028198
R6695 VDDA.n664 VDDA.n541 0.028198
R6696 VDDA.n656 VDDA.n539 0.028198
R6697 VDDA.n563 VDDA.n538 0.028198
R6698 VDDA.n567 VDDA.n536 0.028198
R6699 VDDA.n640 VDDA.n535 0.028198
R6700 VDDA.n632 VDDA.n533 0.028198
R6701 VDDA.n575 VDDA.n532 0.028198
R6702 VDDA.n579 VDDA.n530 0.028198
R6703 VDDA.n616 VDDA.n529 0.028198
R6704 VDDA.n608 VDDA.n527 0.028198
R6705 VDDA.n587 VDDA.n526 0.028198
R6706 VDDA.n591 VDDA.n524 0.028198
R6707 VDDA.n592 VDDA.n523 0.028198
R6708 VDDA.n1660 VDDA.n1525 0.028198
R6709 VDDA.n1531 VDDA.n1524 0.028198
R6710 VDDA.n1535 VDDA.n1522 0.028198
R6711 VDDA.n1644 VDDA.n1521 0.028198
R6712 VDDA.n1636 VDDA.n1519 0.028198
R6713 VDDA.n1543 VDDA.n1518 0.028198
R6714 VDDA.n1547 VDDA.n1516 0.028198
R6715 VDDA.n1620 VDDA.n1515 0.028198
R6716 VDDA.n1612 VDDA.n1513 0.028198
R6717 VDDA.n1555 VDDA.n1512 0.028198
R6718 VDDA.n1559 VDDA.n1510 0.028198
R6719 VDDA.n1596 VDDA.n1509 0.028198
R6720 VDDA.n1588 VDDA.n1507 0.028198
R6721 VDDA.n1567 VDDA.n1506 0.028198
R6722 VDDA.n1571 VDDA.n1504 0.028198
R6723 VDDA.n1572 VDDA.n1503 0.028198
R6724 VDDA.n1826 VDDA.n1825 0.028198
R6725 VDDA.n1819 VDDA.n1690 0.028198
R6726 VDDA.n1811 VDDA.n1688 0.028198
R6727 VDDA.n1700 VDDA.n1687 0.028198
R6728 VDDA.n1704 VDDA.n1685 0.028198
R6729 VDDA.n1795 VDDA.n1684 0.028198
R6730 VDDA.n1787 VDDA.n1682 0.028198
R6731 VDDA.n1712 VDDA.n1681 0.028198
R6732 VDDA.n1716 VDDA.n1679 0.028198
R6733 VDDA.n1771 VDDA.n1678 0.028198
R6734 VDDA.n1763 VDDA.n1676 0.028198
R6735 VDDA.n1724 VDDA.n1675 0.028198
R6736 VDDA.n1728 VDDA.n1673 0.028198
R6737 VDDA.n1747 VDDA.n1672 0.028198
R6738 VDDA.n1739 VDDA.n1670 0.028198
R6739 VDDA.n1735 VDDA.n1669 0.028198
R6740 VDDA.n513 VDDA.n378 0.028198
R6741 VDDA.n384 VDDA.n377 0.028198
R6742 VDDA.n388 VDDA.n375 0.028198
R6743 VDDA.n497 VDDA.n374 0.028198
R6744 VDDA.n489 VDDA.n372 0.028198
R6745 VDDA.n396 VDDA.n371 0.028198
R6746 VDDA.n400 VDDA.n369 0.028198
R6747 VDDA.n473 VDDA.n368 0.028198
R6748 VDDA.n465 VDDA.n366 0.028198
R6749 VDDA.n408 VDDA.n365 0.028198
R6750 VDDA.n412 VDDA.n363 0.028198
R6751 VDDA.n449 VDDA.n362 0.028198
R6752 VDDA.n441 VDDA.n360 0.028198
R6753 VDDA.n420 VDDA.n359 0.028198
R6754 VDDA.n424 VDDA.n357 0.028198
R6755 VDDA.n425 VDDA.n356 0.028198
R6756 VDDA.n3019 VDDA.n2884 0.028198
R6757 VDDA.n2890 VDDA.n2883 0.028198
R6758 VDDA.n2894 VDDA.n2881 0.028198
R6759 VDDA.n3003 VDDA.n2880 0.028198
R6760 VDDA.n2995 VDDA.n2878 0.028198
R6761 VDDA.n2902 VDDA.n2877 0.028198
R6762 VDDA.n2906 VDDA.n2875 0.028198
R6763 VDDA.n2979 VDDA.n2874 0.028198
R6764 VDDA.n2971 VDDA.n2872 0.028198
R6765 VDDA.n2914 VDDA.n2871 0.028198
R6766 VDDA.n2918 VDDA.n2869 0.028198
R6767 VDDA.n2955 VDDA.n2868 0.028198
R6768 VDDA.n2947 VDDA.n2866 0.028198
R6769 VDDA.n2926 VDDA.n2865 0.028198
R6770 VDDA.n2930 VDDA.n2863 0.028198
R6771 VDDA.n2931 VDDA.n2862 0.028198
R6772 VDDA.n3185 VDDA.n3184 0.028198
R6773 VDDA.n3178 VDDA.n3049 0.028198
R6774 VDDA.n3170 VDDA.n3047 0.028198
R6775 VDDA.n3059 VDDA.n3046 0.028198
R6776 VDDA.n3063 VDDA.n3044 0.028198
R6777 VDDA.n3154 VDDA.n3043 0.028198
R6778 VDDA.n3146 VDDA.n3041 0.028198
R6779 VDDA.n3071 VDDA.n3040 0.028198
R6780 VDDA.n3075 VDDA.n3038 0.028198
R6781 VDDA.n3130 VDDA.n3037 0.028198
R6782 VDDA.n3122 VDDA.n3035 0.028198
R6783 VDDA.n3083 VDDA.n3034 0.028198
R6784 VDDA.n3087 VDDA.n3032 0.028198
R6785 VDDA.n3106 VDDA.n3031 0.028198
R6786 VDDA.n3098 VDDA.n3029 0.028198
R6787 VDDA.n3094 VDDA.n3028 0.028198
R6788 VDDA.n3351 VDDA.n3350 0.028198
R6789 VDDA.n3344 VDDA.n3343 0.028198
R6790 VDDA.n3334 VDDA.n3333 0.028198
R6791 VDDA.n3331 VDDA.n3330 0.028198
R6792 VDDA.n3321 VDDA.n3320 0.028198
R6793 VDDA.n3314 VDDA.n3313 0.028198
R6794 VDDA.n3304 VDDA.n3303 0.028198
R6795 VDDA.n3301 VDDA.n3300 0.028198
R6796 VDDA.n3291 VDDA.n3290 0.028198
R6797 VDDA.n3284 VDDA.n3283 0.028198
R6798 VDDA.n3274 VDDA.n3273 0.028198
R6799 VDDA.n3271 VDDA.n3270 0.028198
R6800 VDDA.n3261 VDDA.n3260 0.028198
R6801 VDDA.n3254 VDDA.n3253 0.028198
R6802 VDDA.n3244 VDDA.n3243 0.028198
R6803 VDDA.n3241 VDDA.n3240 0.028198
R6804 VDDA.n176 VDDA.n41 0.028198
R6805 VDDA.n47 VDDA.n40 0.028198
R6806 VDDA.n51 VDDA.n38 0.028198
R6807 VDDA.n160 VDDA.n37 0.028198
R6808 VDDA.n152 VDDA.n35 0.028198
R6809 VDDA.n59 VDDA.n34 0.028198
R6810 VDDA.n63 VDDA.n32 0.028198
R6811 VDDA.n136 VDDA.n31 0.028198
R6812 VDDA.n128 VDDA.n29 0.028198
R6813 VDDA.n71 VDDA.n28 0.028198
R6814 VDDA.n75 VDDA.n26 0.028198
R6815 VDDA.n112 VDDA.n25 0.028198
R6816 VDDA.n104 VDDA.n23 0.028198
R6817 VDDA.n83 VDDA.n22 0.028198
R6818 VDDA.n87 VDDA.n20 0.028198
R6819 VDDA.n88 VDDA.n19 0.028198
R6820 VDDA.n2527 VDDA.n1874 0.028198
R6821 VDDA.n2523 VDDA.n1873 0.028198
R6822 VDDA.n2513 VDDA.n1871 0.028198
R6823 VDDA.n2507 VDDA.n1870 0.028198
R6824 VDDA.n2497 VDDA.n1868 0.028198
R6825 VDDA.n2493 VDDA.n1867 0.028198
R6826 VDDA.n2483 VDDA.n1865 0.028198
R6827 VDDA.n2477 VDDA.n1864 0.028198
R6828 VDDA.n2467 VDDA.n1862 0.028198
R6829 VDDA.n2463 VDDA.n1861 0.028198
R6830 VDDA.n2453 VDDA.n1859 0.028198
R6831 VDDA.n2447 VDDA.n1858 0.028198
R6832 VDDA.n2437 VDDA.n1856 0.028198
R6833 VDDA.n2433 VDDA.n1855 0.028198
R6834 VDDA.n2423 VDDA.n1853 0.028198
R6835 VDDA.n2417 VDDA.n1852 0.028198
R6836 VDDA.n2672 VDDA.n1850 0.028198
R6837 VDDA.n2668 VDDA.n1849 0.028198
R6838 VDDA.n2658 VDDA.n1847 0.028198
R6839 VDDA.n2652 VDDA.n1846 0.028198
R6840 VDDA.n2642 VDDA.n1844 0.028198
R6841 VDDA.n2638 VDDA.n1843 0.028198
R6842 VDDA.n2628 VDDA.n1841 0.028198
R6843 VDDA.n2622 VDDA.n1840 0.028198
R6844 VDDA.n2612 VDDA.n1838 0.028198
R6845 VDDA.n2608 VDDA.n1837 0.028198
R6846 VDDA.n2598 VDDA.n1835 0.028198
R6847 VDDA.n2592 VDDA.n1834 0.028198
R6848 VDDA.n2582 VDDA.n1832 0.028198
R6849 VDDA.n2578 VDDA.n1831 0.028198
R6850 VDDA.n2568 VDDA.n1829 0.028198
R6851 VDDA.n2562 VDDA.n1828 0.028198
R6852 VDDA.n349 VDDA.n207 0.028198
R6853 VDDA.n345 VDDA.n206 0.028198
R6854 VDDA.n335 VDDA.n204 0.028198
R6855 VDDA.n329 VDDA.n203 0.028198
R6856 VDDA.n319 VDDA.n201 0.028198
R6857 VDDA.n315 VDDA.n200 0.028198
R6858 VDDA.n305 VDDA.n198 0.028198
R6859 VDDA.n299 VDDA.n197 0.028198
R6860 VDDA.n289 VDDA.n195 0.028198
R6861 VDDA.n285 VDDA.n194 0.028198
R6862 VDDA.n275 VDDA.n192 0.028198
R6863 VDDA.n269 VDDA.n191 0.028198
R6864 VDDA.n259 VDDA.n189 0.028198
R6865 VDDA.n255 VDDA.n188 0.028198
R6866 VDDA.n245 VDDA.n186 0.028198
R6867 VDDA.n239 VDDA.n185 0.028198
R6868 VDDA.n2146 VDDA.n1922 0.028198
R6869 VDDA.n2142 VDDA.n1921 0.028198
R6870 VDDA.n2132 VDDA.n1919 0.028198
R6871 VDDA.n2126 VDDA.n1918 0.028198
R6872 VDDA.n2116 VDDA.n1916 0.028198
R6873 VDDA.n2112 VDDA.n1915 0.028198
R6874 VDDA.n2102 VDDA.n1913 0.028198
R6875 VDDA.n2096 VDDA.n1912 0.028198
R6876 VDDA.n2086 VDDA.n1910 0.028198
R6877 VDDA.n2082 VDDA.n1909 0.028198
R6878 VDDA.n2072 VDDA.n1907 0.028198
R6879 VDDA.n2066 VDDA.n1906 0.028198
R6880 VDDA.n2056 VDDA.n1904 0.028198
R6881 VDDA.n2052 VDDA.n1903 0.028198
R6882 VDDA.n2042 VDDA.n1901 0.028198
R6883 VDDA.n2036 VDDA.n1900 0.028198
R6884 VDDA.n2331 VDDA.n1898 0.028198
R6885 VDDA.n2327 VDDA.n1897 0.028198
R6886 VDDA.n2317 VDDA.n1895 0.028198
R6887 VDDA.n2311 VDDA.n1894 0.028198
R6888 VDDA.n2301 VDDA.n1892 0.028198
R6889 VDDA.n2297 VDDA.n1891 0.028198
R6890 VDDA.n2287 VDDA.n1889 0.028198
R6891 VDDA.n2281 VDDA.n1888 0.028198
R6892 VDDA.n2271 VDDA.n1886 0.028198
R6893 VDDA.n2267 VDDA.n1885 0.028198
R6894 VDDA.n2257 VDDA.n1883 0.028198
R6895 VDDA.n2251 VDDA.n1882 0.028198
R6896 VDDA.n2241 VDDA.n1880 0.028198
R6897 VDDA.n2237 VDDA.n1879 0.028198
R6898 VDDA.n2227 VDDA.n1877 0.028198
R6899 VDDA.n2221 VDDA.n1876 0.028198
R6900 VDDA.n2236 VDDA.n1878 0.0243392
R6901 VDDA.n2250 VDDA.n1881 0.0243392
R6902 VDDA.n2266 VDDA.n1884 0.0243392
R6903 VDDA.n2280 VDDA.n1887 0.0243392
R6904 VDDA.n2296 VDDA.n1890 0.0243392
R6905 VDDA.n2310 VDDA.n1893 0.0243392
R6906 VDDA.n2326 VDDA.n1896 0.0243392
R6907 VDDA.n2051 VDDA.n1902 0.0243392
R6908 VDDA.n2065 VDDA.n1905 0.0243392
R6909 VDDA.n2081 VDDA.n1908 0.0243392
R6910 VDDA.n2095 VDDA.n1911 0.0243392
R6911 VDDA.n2111 VDDA.n1914 0.0243392
R6912 VDDA.n2125 VDDA.n1917 0.0243392
R6913 VDDA.n2141 VDDA.n1920 0.0243392
R6914 VDDA.n254 VDDA.n187 0.0243392
R6915 VDDA.n268 VDDA.n190 0.0243392
R6916 VDDA.n284 VDDA.n193 0.0243392
R6917 VDDA.n298 VDDA.n196 0.0243392
R6918 VDDA.n314 VDDA.n199 0.0243392
R6919 VDDA.n328 VDDA.n202 0.0243392
R6920 VDDA.n344 VDDA.n205 0.0243392
R6921 VDDA.n2577 VDDA.n1830 0.0243392
R6922 VDDA.n2591 VDDA.n1833 0.0243392
R6923 VDDA.n2607 VDDA.n1836 0.0243392
R6924 VDDA.n2621 VDDA.n1839 0.0243392
R6925 VDDA.n2637 VDDA.n1842 0.0243392
R6926 VDDA.n2651 VDDA.n1845 0.0243392
R6927 VDDA.n2667 VDDA.n1848 0.0243392
R6928 VDDA.n2432 VDDA.n1854 0.0243392
R6929 VDDA.n2446 VDDA.n1857 0.0243392
R6930 VDDA.n2462 VDDA.n1860 0.0243392
R6931 VDDA.n2476 VDDA.n1863 0.0243392
R6932 VDDA.n2492 VDDA.n1866 0.0243392
R6933 VDDA.n2506 VDDA.n1869 0.0243392
R6934 VDDA.n2522 VDDA.n1872 0.0243392
R6935 VDDA.n82 VDDA.n21 0.0243392
R6936 VDDA.n111 VDDA.n24 0.0243392
R6937 VDDA.n70 VDDA.n27 0.0243392
R6938 VDDA.n135 VDDA.n30 0.0243392
R6939 VDDA.n58 VDDA.n33 0.0243392
R6940 VDDA.n159 VDDA.n36 0.0243392
R6941 VDDA.n46 VDDA.n39 0.0243392
R6942 VDDA.n3252 VDDA.n3251 0.0243392
R6943 VDDA.n3263 VDDA.n3225 0.0243392
R6944 VDDA.n3282 VDDA.n3281 0.0243392
R6945 VDDA.n3293 VDDA.n3213 0.0243392
R6946 VDDA.n3312 VDDA.n3311 0.0243392
R6947 VDDA.n3323 VDDA.n3201 0.0243392
R6948 VDDA.n3342 VDDA.n3341 0.0243392
R6949 VDDA.n3105 VDDA.n3030 0.0243392
R6950 VDDA.n3082 VDDA.n3033 0.0243392
R6951 VDDA.n3129 VDDA.n3036 0.0243392
R6952 VDDA.n3070 VDDA.n3039 0.0243392
R6953 VDDA.n3153 VDDA.n3042 0.0243392
R6954 VDDA.n3058 VDDA.n3045 0.0243392
R6955 VDDA.n3177 VDDA.n3048 0.0243392
R6956 VDDA.n2925 VDDA.n2864 0.0243392
R6957 VDDA.n2954 VDDA.n2867 0.0243392
R6958 VDDA.n2913 VDDA.n2870 0.0243392
R6959 VDDA.n2978 VDDA.n2873 0.0243392
R6960 VDDA.n2901 VDDA.n2876 0.0243392
R6961 VDDA.n3002 VDDA.n2879 0.0243392
R6962 VDDA.n2889 VDDA.n2882 0.0243392
R6963 VDDA.n419 VDDA.n358 0.0243392
R6964 VDDA.n448 VDDA.n361 0.0243392
R6965 VDDA.n407 VDDA.n364 0.0243392
R6966 VDDA.n472 VDDA.n367 0.0243392
R6967 VDDA.n395 VDDA.n370 0.0243392
R6968 VDDA.n496 VDDA.n373 0.0243392
R6969 VDDA.n383 VDDA.n376 0.0243392
R6970 VDDA.n1746 VDDA.n1671 0.0243392
R6971 VDDA.n1723 VDDA.n1674 0.0243392
R6972 VDDA.n1770 VDDA.n1677 0.0243392
R6973 VDDA.n1711 VDDA.n1680 0.0243392
R6974 VDDA.n1794 VDDA.n1683 0.0243392
R6975 VDDA.n1699 VDDA.n1686 0.0243392
R6976 VDDA.n1818 VDDA.n1689 0.0243392
R6977 VDDA.n1566 VDDA.n1505 0.0243392
R6978 VDDA.n1595 VDDA.n1508 0.0243392
R6979 VDDA.n1554 VDDA.n1511 0.0243392
R6980 VDDA.n1619 VDDA.n1514 0.0243392
R6981 VDDA.n1542 VDDA.n1517 0.0243392
R6982 VDDA.n1643 VDDA.n1520 0.0243392
R6983 VDDA.n1530 VDDA.n1523 0.0243392
R6984 VDDA.n586 VDDA.n525 0.0243392
R6985 VDDA.n615 VDDA.n528 0.0243392
R6986 VDDA.n574 VDDA.n531 0.0243392
R6987 VDDA.n639 VDDA.n534 0.0243392
R6988 VDDA.n562 VDDA.n537 0.0243392
R6989 VDDA.n663 VDDA.n540 0.0243392
R6990 VDDA.n550 VDDA.n543 0.0243392
R6991 VDDA.n1392 VDDA.n1391 0.0243392
R6992 VDDA.n1403 VDDA.n1365 0.0243392
R6993 VDDA.n1422 VDDA.n1421 0.0243392
R6994 VDDA.n1433 VDDA.n1353 0.0243392
R6995 VDDA.n1452 VDDA.n1451 0.0243392
R6996 VDDA.n1463 VDDA.n1341 0.0243392
R6997 VDDA.n1482 VDDA.n1481 0.0243392
R6998 VDDA.n1228 VDDA.n1171 0.0243392
R6999 VDDA.n1244 VDDA.n1174 0.0243392
R7000 VDDA.n1258 VDDA.n1177 0.0243392
R7001 VDDA.n1274 VDDA.n1180 0.0243392
R7002 VDDA.n1288 VDDA.n1183 0.0243392
R7003 VDDA.n1304 VDDA.n1186 0.0243392
R7004 VDDA.n1318 VDDA.n1189 0.0243392
R7005 VDDA.n1315 VDDA.n1189 0.0243392
R7006 VDDA.n1299 VDDA.n1186 0.0243392
R7007 VDDA.n1285 VDDA.n1183 0.0243392
R7008 VDDA.n1269 VDDA.n1180 0.0243392
R7009 VDDA.n1255 VDDA.n1177 0.0243392
R7010 VDDA.n1239 VDDA.n1174 0.0243392
R7011 VDDA.n1225 VDDA.n1171 0.0243392
R7012 VDDA.n1481 VDDA.n1480 0.0243392
R7013 VDDA.n1464 VDDA.n1463 0.0243392
R7014 VDDA.n1451 VDDA.n1450 0.0243392
R7015 VDDA.n1434 VDDA.n1433 0.0243392
R7016 VDDA.n1421 VDDA.n1420 0.0243392
R7017 VDDA.n1404 VDDA.n1403 0.0243392
R7018 VDDA.n1391 VDDA.n1390 0.0243392
R7019 VDDA.n672 VDDA.n543 0.0243392
R7020 VDDA.n559 VDDA.n540 0.0243392
R7021 VDDA.n648 VDDA.n537 0.0243392
R7022 VDDA.n571 VDDA.n534 0.0243392
R7023 VDDA.n624 VDDA.n531 0.0243392
R7024 VDDA.n583 VDDA.n528 0.0243392
R7025 VDDA.n600 VDDA.n525 0.0243392
R7026 VDDA.n1652 VDDA.n1523 0.0243392
R7027 VDDA.n1539 VDDA.n1520 0.0243392
R7028 VDDA.n1628 VDDA.n1517 0.0243392
R7029 VDDA.n1551 VDDA.n1514 0.0243392
R7030 VDDA.n1604 VDDA.n1511 0.0243392
R7031 VDDA.n1563 VDDA.n1508 0.0243392
R7032 VDDA.n1580 VDDA.n1505 0.0243392
R7033 VDDA.n1696 VDDA.n1689 0.0243392
R7034 VDDA.n1803 VDDA.n1686 0.0243392
R7035 VDDA.n1708 VDDA.n1683 0.0243392
R7036 VDDA.n1779 VDDA.n1680 0.0243392
R7037 VDDA.n1720 VDDA.n1677 0.0243392
R7038 VDDA.n1755 VDDA.n1674 0.0243392
R7039 VDDA.n1732 VDDA.n1671 0.0243392
R7040 VDDA.n505 VDDA.n376 0.0243392
R7041 VDDA.n392 VDDA.n373 0.0243392
R7042 VDDA.n481 VDDA.n370 0.0243392
R7043 VDDA.n404 VDDA.n367 0.0243392
R7044 VDDA.n457 VDDA.n364 0.0243392
R7045 VDDA.n416 VDDA.n361 0.0243392
R7046 VDDA.n433 VDDA.n358 0.0243392
R7047 VDDA.n3011 VDDA.n2882 0.0243392
R7048 VDDA.n2898 VDDA.n2879 0.0243392
R7049 VDDA.n2987 VDDA.n2876 0.0243392
R7050 VDDA.n2910 VDDA.n2873 0.0243392
R7051 VDDA.n2963 VDDA.n2870 0.0243392
R7052 VDDA.n2922 VDDA.n2867 0.0243392
R7053 VDDA.n2939 VDDA.n2864 0.0243392
R7054 VDDA.n3055 VDDA.n3048 0.0243392
R7055 VDDA.n3162 VDDA.n3045 0.0243392
R7056 VDDA.n3067 VDDA.n3042 0.0243392
R7057 VDDA.n3138 VDDA.n3039 0.0243392
R7058 VDDA.n3079 VDDA.n3036 0.0243392
R7059 VDDA.n3114 VDDA.n3033 0.0243392
R7060 VDDA.n3091 VDDA.n3030 0.0243392
R7061 VDDA.n3341 VDDA.n3340 0.0243392
R7062 VDDA.n3324 VDDA.n3323 0.0243392
R7063 VDDA.n3311 VDDA.n3310 0.0243392
R7064 VDDA.n3294 VDDA.n3293 0.0243392
R7065 VDDA.n3281 VDDA.n3280 0.0243392
R7066 VDDA.n3264 VDDA.n3263 0.0243392
R7067 VDDA.n3251 VDDA.n3250 0.0243392
R7068 VDDA.n168 VDDA.n39 0.0243392
R7069 VDDA.n55 VDDA.n36 0.0243392
R7070 VDDA.n144 VDDA.n33 0.0243392
R7071 VDDA.n67 VDDA.n30 0.0243392
R7072 VDDA.n120 VDDA.n27 0.0243392
R7073 VDDA.n79 VDDA.n24 0.0243392
R7074 VDDA.n96 VDDA.n21 0.0243392
R7075 VDDA.n2517 VDDA.n1872 0.0243392
R7076 VDDA.n2503 VDDA.n1869 0.0243392
R7077 VDDA.n2487 VDDA.n1866 0.0243392
R7078 VDDA.n2473 VDDA.n1863 0.0243392
R7079 VDDA.n2457 VDDA.n1860 0.0243392
R7080 VDDA.n2443 VDDA.n1857 0.0243392
R7081 VDDA.n2427 VDDA.n1854 0.0243392
R7082 VDDA.n2662 VDDA.n1848 0.0243392
R7083 VDDA.n2648 VDDA.n1845 0.0243392
R7084 VDDA.n2632 VDDA.n1842 0.0243392
R7085 VDDA.n2618 VDDA.n1839 0.0243392
R7086 VDDA.n2602 VDDA.n1836 0.0243392
R7087 VDDA.n2588 VDDA.n1833 0.0243392
R7088 VDDA.n2572 VDDA.n1830 0.0243392
R7089 VDDA.n339 VDDA.n205 0.0243392
R7090 VDDA.n325 VDDA.n202 0.0243392
R7091 VDDA.n309 VDDA.n199 0.0243392
R7092 VDDA.n295 VDDA.n196 0.0243392
R7093 VDDA.n279 VDDA.n193 0.0243392
R7094 VDDA.n265 VDDA.n190 0.0243392
R7095 VDDA.n249 VDDA.n187 0.0243392
R7096 VDDA.n2136 VDDA.n1920 0.0243392
R7097 VDDA.n2122 VDDA.n1917 0.0243392
R7098 VDDA.n2106 VDDA.n1914 0.0243392
R7099 VDDA.n2092 VDDA.n1911 0.0243392
R7100 VDDA.n2076 VDDA.n1908 0.0243392
R7101 VDDA.n2062 VDDA.n1905 0.0243392
R7102 VDDA.n2046 VDDA.n1902 0.0243392
R7103 VDDA.n2321 VDDA.n1896 0.0243392
R7104 VDDA.n2307 VDDA.n1893 0.0243392
R7105 VDDA.n2291 VDDA.n1890 0.0243392
R7106 VDDA.n2277 VDDA.n1887 0.0243392
R7107 VDDA.n2261 VDDA.n1884 0.0243392
R7108 VDDA.n2247 VDDA.n1881 0.0243392
R7109 VDDA.n2231 VDDA.n1878 0.0243392
R7110 VDDA.n2151 VDDA.n354 0.0129844
R7111 VDDA.n1667 VDDA.n1501 0.0107812
R7112 VDDA.n3186 VDDA.n3026 0.0107812
R7113 VDDA.n2532 VDDA.n2336 0.0101203
R7114 VDDA VDDA.n3467 0.00879844
R7115 VDDA.n2860 VDDA.n354 0.00586094
R7116 VDDA.n1327 VDDA.n521 0.00564062
R7117 VDDA.n1501 VDDA.n521 0.00564062
R7118 VDDA.n2678 VDDA.n1667 0.00564062
R7119 VDDA.n3026 VDDA.n2860 0.00564062
R7120 VDDA.n3186 VDDA.n17 0.00564062
R7121 VDDA.n3360 VDDA.n17 0.00564062
R7122 VDDA.n2678 VDDA.n2677 0.00534688
R7123 VDDA.n2677 VDDA.n2532 0.00475937
R7124 VDDA.n3466 VDDA.n3376 0.00189531
R7125 VDDA.n3376 VDDA.n16 0.00189531
R7126 VDDA.n3425 VDDA.n3 0.00188102
R7127 VDDA.n3429 VDDA.n7 0.00188102
R7128 VDDA.n3433 VDDA.n11 0.00188102
R7129 VDDA.n3380 VDDA.n3374 0.00188102
R7130 VDDA.n3386 VDDA.n3372 0.00188102
R7131 VDDA.n3392 VDDA.n3370 0.00188102
R7132 VDDA.n3398 VDDA.n3368 0.00188102
R7133 VDDA.n3404 VDDA.n3366 0.00188102
R7134 VDDA.n3410 VDDA.n3364 0.00188102
R7135 VDDA.n3416 VDDA.n3362 0.00188102
R7136 VDDA.n3444 VDDA.n11 0.00188102
R7137 VDDA.n3452 VDDA.n7 0.00188102
R7138 VDDA.n3460 VDDA.n3 0.00188102
R7139 VDDA.n3381 VDDA.n3380 0.00188102
R7140 VDDA.n3387 VDDA.n3386 0.00188102
R7141 VDDA.n3393 VDDA.n3392 0.00188102
R7142 VDDA.n3399 VDDA.n3398 0.00188102
R7143 VDDA.n3405 VDDA.n3404 0.00188102
R7144 VDDA.n3411 VDDA.n3410 0.00188102
R7145 VDDA.n3417 VDDA.n3416 0.00188102
R7146 VDDA.n3423 VDDA.n3422 0.00173422
R7147 VDDA.n3423 VDDA.n1 0.00173422
R7148 VDDA.n3463 VDDA.n3424 0.00173422
R7149 VDDA.n3457 VDDA.n3427 0.00173422
R7150 VDDA.n3427 VDDA.n5 0.00173422
R7151 VDDA.n3455 VDDA.n3428 0.00173422
R7152 VDDA.n3449 VDDA.n3431 0.00173422
R7153 VDDA.n3431 VDDA.n9 0.00173422
R7154 VDDA.n3447 VDDA.n3432 0.00173422
R7155 VDDA.n3441 VDDA.n3435 0.00173422
R7156 VDDA.n3435 VDDA.n13 0.00173422
R7157 VDDA.n3439 VDDA.n3436 0.00173422
R7158 VDDA.n3377 VDDA.n3375 0.00173422
R7159 VDDA.n3383 VDDA.n3373 0.00173422
R7160 VDDA.n3389 VDDA.n3371 0.00173422
R7161 VDDA.n3395 VDDA.n3369 0.00173422
R7162 VDDA.n3401 VDDA.n3367 0.00173422
R7163 VDDA.n3407 VDDA.n3365 0.00173422
R7164 VDDA.n3413 VDDA.n3363 0.00173422
R7165 VDDA.n3419 VDDA.n3361 0.00173422
R7166 VDDA.n3440 VDDA.n13 0.00173422
R7167 VDDA.n3448 VDDA.n9 0.00173422
R7168 VDDA.n3456 VDDA.n5 0.00173422
R7169 VDDA.n3464 VDDA.n1 0.00173422
R7170 VDDA.n3378 VDDA.n3377 0.00173422
R7171 VDDA.n3440 VDDA.n3439 0.00173422
R7172 VDDA.n3442 VDDA.n3441 0.00173422
R7173 VDDA.n3448 VDDA.n3447 0.00173422
R7174 VDDA.n3450 VDDA.n3449 0.00173422
R7175 VDDA.n3456 VDDA.n3455 0.00173422
R7176 VDDA.n3458 VDDA.n3457 0.00173422
R7177 VDDA.n3464 VDDA.n3463 0.00173422
R7178 VDDA.n3422 VDDA.n16 0.00173422
R7179 VDDA.n3384 VDDA.n3383 0.00173422
R7180 VDDA.n3390 VDDA.n3389 0.00173422
R7181 VDDA.n3396 VDDA.n3395 0.00173422
R7182 VDDA.n3402 VDDA.n3401 0.00173422
R7183 VDDA.n3408 VDDA.n3407 0.00173422
R7184 VDDA.n3414 VDDA.n3413 0.00173422
R7185 VDDA.n3420 VDDA.n3419 0.00173422
R7186 VDDA.n3424 VDDA.n2 0.00169751
R7187 VDDA.n3461 VDDA.n3425 0.00169751
R7188 VDDA.n3459 VDDA.n3426 0.00169751
R7189 VDDA.n3426 VDDA.n4 0.00169751
R7190 VDDA.n3428 VDDA.n6 0.00169751
R7191 VDDA.n3453 VDDA.n3429 0.00169751
R7192 VDDA.n3451 VDDA.n3430 0.00169751
R7193 VDDA.n3430 VDDA.n8 0.00169751
R7194 VDDA.n3432 VDDA.n10 0.00169751
R7195 VDDA.n3445 VDDA.n3433 0.00169751
R7196 VDDA.n3443 VDDA.n3434 0.00169751
R7197 VDDA.n3434 VDDA.n12 0.00169751
R7198 VDDA.n3436 VDDA.n14 0.00169751
R7199 VDDA.n3438 VDDA.n15 0.00169751
R7200 VDDA.n3437 VDDA.n14 0.00169751
R7201 VDDA.n3442 VDDA.n12 0.00169751
R7202 VDDA.n3446 VDDA.n10 0.00169751
R7203 VDDA.n3450 VDDA.n8 0.00169751
R7204 VDDA.n3454 VDDA.n6 0.00169751
R7205 VDDA.n3458 VDDA.n4 0.00169751
R7206 VDDA.n3462 VDDA.n2 0.00169751
R7207 VDDA.n3444 VDDA.n3443 0.00169751
R7208 VDDA.n3446 VDDA.n3445 0.00169751
R7209 VDDA.n3452 VDDA.n3451 0.00169751
R7210 VDDA.n3454 VDDA.n3453 0.00169751
R7211 VDDA.n3460 VDDA.n3459 0.00169751
R7212 VDDA.n3462 VDDA.n3461 0.00169751
R7213 VDDA.n3438 VDDA.n3437 0.00169751
R7214 VDDA.n3378 VDDA.n0 0.00166081
R7215 VDDA.n3381 VDDA.n3379 0.00166081
R7216 VDDA.n3384 VDDA.n3382 0.00166081
R7217 VDDA.n3387 VDDA.n3385 0.00166081
R7218 VDDA.n3390 VDDA.n3388 0.00166081
R7219 VDDA.n3393 VDDA.n3391 0.00166081
R7220 VDDA.n3396 VDDA.n3394 0.00166081
R7221 VDDA.n3399 VDDA.n3397 0.00166081
R7222 VDDA.n3402 VDDA.n3400 0.00166081
R7223 VDDA.n3405 VDDA.n3403 0.00166081
R7224 VDDA.n3408 VDDA.n3406 0.00166081
R7225 VDDA.n3411 VDDA.n3409 0.00166081
R7226 VDDA.n3414 VDDA.n3412 0.00166081
R7227 VDDA.n3417 VDDA.n3415 0.00166081
R7228 VDDA.n3420 VDDA.n3418 0.00166081
R7229 VDDA.n3465 VDDA.n3421 0.00166081
R7230 VDDA.n3467 VDDA.n0 0.00166081
R7231 VDDA.n3379 VDDA.n3375 0.00166081
R7232 VDDA.n3382 VDDA.n3374 0.00166081
R7233 VDDA.n3385 VDDA.n3373 0.00166081
R7234 VDDA.n3388 VDDA.n3372 0.00166081
R7235 VDDA.n3391 VDDA.n3371 0.00166081
R7236 VDDA.n3394 VDDA.n3370 0.00166081
R7237 VDDA.n3397 VDDA.n3369 0.00166081
R7238 VDDA.n3400 VDDA.n3368 0.00166081
R7239 VDDA.n3403 VDDA.n3367 0.00166081
R7240 VDDA.n3406 VDDA.n3366 0.00166081
R7241 VDDA.n3409 VDDA.n3365 0.00166081
R7242 VDDA.n3412 VDDA.n3364 0.00166081
R7243 VDDA.n3415 VDDA.n3363 0.00166081
R7244 VDDA.n3418 VDDA.n3362 0.00166081
R7245 VDDA.n3421 VDDA.n3361 0.00166081
R7246 VDDA.t118 VDDA.n232 0.00152174
R7247 VDDA.t107 VDDA.n233 0.00152174
R7248 VDDA.t228 VDDA.n234 0.00152174
R7249 VDDA.t214 VDDA.n235 0.00152174
R7250 VDDA.t73 VDDA.n236 0.00152174
R7251 GNDA.n632 GNDA.n631 458822
R7252 GNDA.n1344 GNDA.n626 164529
R7253 GNDA.n631 GNDA.n628 112519
R7254 GNDA.n631 GNDA.n625 86240
R7255 GNDA.n632 GNDA.t33 63867.8
R7256 GNDA.n4101 GNDA.n4100 50290
R7257 GNDA.n6098 GNDA.n1344 41014.3
R7258 GNDA.n6096 GNDA.n6095 30702.9
R7259 GNDA.n6099 GNDA.n626 25923.2
R7260 GNDA.n6098 GNDA.n6097 25066.7
R7261 GNDA.n6099 GNDA.n628 23672.9
R7262 GNDA.n4102 GNDA.n632 20341
R7263 GNDA.n6102 GNDA.n6101 18211.5
R7264 GNDA.n1345 GNDA.n633 13528.5
R7265 GNDA.n4105 GNDA.n4104 11440
R7266 GNDA.n6097 GNDA.n6096 10513.3
R7267 GNDA.n4102 GNDA.n4101 10148.9
R7268 GNDA.n6101 GNDA.n6100 9910.09
R7269 GNDA.n6100 GNDA.n627 9724.16
R7270 GNDA.n4107 GNDA.n4099 9626.42
R7271 GNDA.n6094 GNDA.n1347 9611.7
R7272 GNDA.n6102 GNDA.n625 8404
R7273 GNDA.n4106 GNDA.n4105 8346.79
R7274 GNDA.n4105 GNDA.n1346 8346.79
R7275 GNDA.n6100 GNDA.n6099 7676.92
R7276 GNDA.n6099 GNDA.n633 6600
R7277 GNDA.n4103 GNDA.n4102 6089.82
R7278 GNDA.n4103 GNDA.n633 5672.23
R7279 GNDA.n4104 GNDA.n1345 4754.02
R7280 GNDA.n4100 GNDA.t29 4218.68
R7281 GNDA.n627 GNDA.n625 4106.67
R7282 GNDA.n6097 GNDA.n1345 4096.55
R7283 GNDA.n6103 GNDA.n6102 3974.19
R7284 GNDA.n6099 GNDA.n6098 3666.67
R7285 GNDA.n6099 GNDA.n632 2975.41
R7286 GNDA.n1344 GNDA.t446 2523.88
R7287 GNDA.n6095 GNDA.t131 2149.15
R7288 GNDA.n6095 GNDA.n1344 2057.79
R7289 GNDA.n4104 GNDA.n4103 2042.87
R7290 GNDA.n4100 GNDA.t877 1916.55
R7291 GNDA.n6703 GNDA.n6702 1422.12
R7292 GNDA.n6230 GNDA.n560 1185.07
R7293 GNDA.n6230 GNDA.n6229 1185.07
R7294 GNDA.n4106 GNDA.n4101 1141.98
R7295 GNDA.n6096 GNDA.n1346 1141.98
R7296 GNDA.n6101 GNDA.n626 927.471
R7297 GNDA.n628 GNDA.n627 776.471
R7298 GNDA.n6091 GNDA.t837 747.734
R7299 GNDA.n4796 GNDA.t799 747.734
R7300 GNDA.n4093 GNDA.t745 747.734
R7301 GNDA.n4096 GNDA.t818 747.734
R7302 GNDA.n6244 GNDA.n6243 686.717
R7303 GNDA.n961 GNDA.n559 686.717
R7304 GNDA.n1333 GNDA.n1332 686.717
R7305 GNDA.n1332 GNDA.n634 686.717
R7306 GNDA.n955 GNDA.n948 686.717
R7307 GNDA.n6240 GNDA.n556 686.717
R7308 GNDA.n6744 GNDA.n6621 669.307
R7309 GNDA.n1595 GNDA.t765 659.367
R7310 GNDA.n4162 GNDA.t834 659.367
R7311 GNDA.n4120 GNDA.t793 659.367
R7312 GNDA.n4124 GNDA.t752 659.367
R7313 GNDA.n630 GNDA.n629 585.003
R7314 GNDA.n926 GNDA.n925 585.001
R7315 GNDA.n1051 GNDA.n1050 585.001
R7316 GNDA.n583 GNDA.n582 585.001
R7317 GNDA.n599 GNDA.n598 585.001
R7318 GNDA.n562 GNDA.n561 585.001
R7319 GNDA.n564 GNDA.n563 585.001
R7320 GNDA.n6262 GNDA.n6261 585.001
R7321 GNDA.n6759 GNDA.n6758 585
R7322 GNDA.n6760 GNDA.n6759 585
R7323 GNDA.n300 GNDA.n299 585
R7324 GNDA.n6761 GNDA.n300 585
R7325 GNDA.n6764 GNDA.n6763 585
R7326 GNDA.n6763 GNDA.n6762 585
R7327 GNDA.n6765 GNDA.n298 585
R7328 GNDA.n298 GNDA.n297 585
R7329 GNDA.n6767 GNDA.n6766 585
R7330 GNDA.n6768 GNDA.n6767 585
R7331 GNDA.n296 GNDA.n295 585
R7332 GNDA.n6769 GNDA.n296 585
R7333 GNDA.n6772 GNDA.n6771 585
R7334 GNDA.n6771 GNDA.n6770 585
R7335 GNDA.n6773 GNDA.n294 585
R7336 GNDA.n294 GNDA.n293 585
R7337 GNDA.n6775 GNDA.n6774 585
R7338 GNDA.n6776 GNDA.n6775 585
R7339 GNDA.n292 GNDA.n291 585
R7340 GNDA.n6777 GNDA.n292 585
R7341 GNDA.n6780 GNDA.n6779 585
R7342 GNDA.n6779 GNDA.n6778 585
R7343 GNDA.n6781 GNDA.n290 585
R7344 GNDA.n290 GNDA.n99 585
R7345 GNDA.n6743 GNDA.n6742 585
R7346 GNDA.n6741 GNDA.n356 585
R7347 GNDA.t743 GNDA.n356 585
R7348 GNDA.n7140 GNDA.n7139 585
R7349 GNDA.n132 GNDA.n130 585
R7350 GNDA.n243 GNDA.n242 585
R7351 GNDA.n245 GNDA.n244 585
R7352 GNDA.n247 GNDA.n246 585
R7353 GNDA.n249 GNDA.n248 585
R7354 GNDA.n251 GNDA.n250 585
R7355 GNDA.n253 GNDA.n252 585
R7356 GNDA.n255 GNDA.n254 585
R7357 GNDA.n257 GNDA.n256 585
R7358 GNDA.n259 GNDA.n258 585
R7359 GNDA.n261 GNDA.n260 585
R7360 GNDA.n692 GNDA.n691 585
R7361 GNDA.n689 GNDA.n688 585
R7362 GNDA.n687 GNDA.n686 585
R7363 GNDA.n685 GNDA.n684 585
R7364 GNDA.n683 GNDA.n682 585
R7365 GNDA.n681 GNDA.n680 585
R7366 GNDA.n679 GNDA.n678 585
R7367 GNDA.n677 GNDA.n676 585
R7368 GNDA.n675 GNDA.n674 585
R7369 GNDA.n673 GNDA.n672 585
R7370 GNDA.n671 GNDA.n670 585
R7371 GNDA.n136 GNDA.n133 585
R7372 GNDA.n846 GNDA.n845 585
R7373 GNDA.n848 GNDA.n847 585
R7374 GNDA.n850 GNDA.n849 585
R7375 GNDA.n852 GNDA.n851 585
R7376 GNDA.n854 GNDA.n853 585
R7377 GNDA.n856 GNDA.n855 585
R7378 GNDA.n858 GNDA.n857 585
R7379 GNDA.n860 GNDA.n859 585
R7380 GNDA.n862 GNDA.n861 585
R7381 GNDA.n864 GNDA.n863 585
R7382 GNDA.n866 GNDA.n865 585
R7383 GNDA.n868 GNDA.n867 585
R7384 GNDA.n7320 GNDA.n7319 585
R7385 GNDA.n7317 GNDA.n54 585
R7386 GNDA.n59 GNDA.n58 585
R7387 GNDA.n7312 GNDA.n7311 585
R7388 GNDA.n7310 GNDA.n7309 585
R7389 GNDA.n7236 GNDA.n63 585
R7390 GNDA.n7238 GNDA.n7237 585
R7391 GNDA.n7243 GNDA.n7242 585
R7392 GNDA.n7241 GNDA.n7234 585
R7393 GNDA.n7249 GNDA.n7248 585
R7394 GNDA.n7251 GNDA.n7250 585
R7395 GNDA.n7232 GNDA.n7231 585
R7396 GNDA.n6897 GNDA.n6896 585
R7397 GNDA.n6894 GNDA.n6893 585
R7398 GNDA.n6892 GNDA.n6891 585
R7399 GNDA.n6808 GNDA.n6784 585
R7400 GNDA.n6810 GNDA.n6809 585
R7401 GNDA.n6814 GNDA.n6813 585
R7402 GNDA.n6816 GNDA.n6815 585
R7403 GNDA.n6823 GNDA.n6822 585
R7404 GNDA.n6821 GNDA.n6806 585
R7405 GNDA.n6829 GNDA.n6828 585
R7406 GNDA.n6831 GNDA.n6830 585
R7407 GNDA.n6804 GNDA.n6803 585
R7408 GNDA.n329 GNDA.n326 585
R7409 GNDA.n330 GNDA.n324 585
R7410 GNDA.n331 GNDA.n323 585
R7411 GNDA.n321 GNDA.n319 585
R7412 GNDA.n337 GNDA.n318 585
R7413 GNDA.n338 GNDA.n316 585
R7414 GNDA.n339 GNDA.n315 585
R7415 GNDA.n313 GNDA.n311 585
R7416 GNDA.n345 GNDA.n310 585
R7417 GNDA.n346 GNDA.n308 585
R7418 GNDA.n347 GNDA.n307 585
R7419 GNDA.n303 GNDA.n302 585
R7420 GNDA.n134 GNDA.n85 585
R7421 GNDA.n7229 GNDA.n85 585
R7422 GNDA.n350 GNDA.n303 585
R7423 GNDA.n348 GNDA.n347 585
R7424 GNDA.n346 GNDA.n305 585
R7425 GNDA.n345 GNDA.n344 585
R7426 GNDA.n342 GNDA.n311 585
R7427 GNDA.n340 GNDA.n339 585
R7428 GNDA.n338 GNDA.n312 585
R7429 GNDA.n337 GNDA.n336 585
R7430 GNDA.n334 GNDA.n319 585
R7431 GNDA.n332 GNDA.n331 585
R7432 GNDA.n330 GNDA.n320 585
R7433 GNDA.n329 GNDA.n328 585
R7434 GNDA.n134 GNDA.n55 585
R7435 GNDA.n7229 GNDA.n55 585
R7436 GNDA.n7115 GNDA.n160 585
R7437 GNDA.n7116 GNDA.n151 585
R7438 GNDA.n7119 GNDA.n150 585
R7439 GNDA.n7120 GNDA.n149 585
R7440 GNDA.n7123 GNDA.n148 585
R7441 GNDA.n7124 GNDA.n147 585
R7442 GNDA.n7127 GNDA.n146 585
R7443 GNDA.n7129 GNDA.n145 585
R7444 GNDA.n7130 GNDA.n144 585
R7445 GNDA.n7131 GNDA.n143 585
R7446 GNDA.n152 GNDA.n135 585
R7447 GNDA.n7137 GNDA.n131 585
R7448 GNDA.n7137 GNDA.n7136 585
R7449 GNDA.n137 GNDA.n135 585
R7450 GNDA.n7132 GNDA.n7131 585
R7451 GNDA.n7130 GNDA.n142 585
R7452 GNDA.n7129 GNDA.n7128 585
R7453 GNDA.n7127 GNDA.n7126 585
R7454 GNDA.n7125 GNDA.n7124 585
R7455 GNDA.n7123 GNDA.n7122 585
R7456 GNDA.n7121 GNDA.n7120 585
R7457 GNDA.n7119 GNDA.n7118 585
R7458 GNDA.n7117 GNDA.n7116 585
R7459 GNDA.n7115 GNDA.n7114 585
R7460 GNDA.n6206 GNDA.n587 585
R7461 GNDA.n6209 GNDA.n6208 585
R7462 GNDA.n590 GNDA.n589 585
R7463 GNDA.n1118 GNDA.n1117 585
R7464 GNDA.n1119 GNDA.n1115 585
R7465 GNDA.n1113 GNDA.n1110 585
R7466 GNDA.n1125 GNDA.n1109 585
R7467 GNDA.n1126 GNDA.n1107 585
R7468 GNDA.n1127 GNDA.n1106 585
R7469 GNDA.n1103 GNDA.n1102 585
R7470 GNDA.n1134 GNDA.n1133 585
R7471 GNDA.n1136 GNDA.n914 585
R7472 GNDA.n914 GNDA.n913 585
R7473 GNDA.n1133 GNDA.n1132 585
R7474 GNDA.n1130 GNDA.n1103 585
R7475 GNDA.n1128 GNDA.n1127 585
R7476 GNDA.n1126 GNDA.n1104 585
R7477 GNDA.n1125 GNDA.n1124 585
R7478 GNDA.n1122 GNDA.n1110 585
R7479 GNDA.n1120 GNDA.n1119 585
R7480 GNDA.n1118 GNDA.n1112 585
R7481 GNDA.n589 GNDA.n588 585
R7482 GNDA.n6210 GNDA.n6209 585
R7483 GNDA.n6212 GNDA.n587 585
R7484 GNDA.n1138 GNDA.n1137 585
R7485 GNDA.n1100 GNDA.n915 585
R7486 GNDA.n1099 GNDA.n1098 585
R7487 GNDA.n1097 GNDA.n1096 585
R7488 GNDA.n1095 GNDA.n917 585
R7489 GNDA.n1093 GNDA.n1092 585
R7490 GNDA.n1091 GNDA.n918 585
R7491 GNDA.n1090 GNDA.n1089 585
R7492 GNDA.n1087 GNDA.n919 585
R7493 GNDA.n1085 GNDA.n1084 585
R7494 GNDA.n1083 GNDA.n920 585
R7495 GNDA.n1082 GNDA.n1081 585
R7496 GNDA.n1163 GNDA.n1162 585
R7497 GNDA.n1161 GNDA.n1160 585
R7498 GNDA.n1159 GNDA.n908 585
R7499 GNDA.n1157 GNDA.n1156 585
R7500 GNDA.n1155 GNDA.n909 585
R7501 GNDA.n1154 GNDA.n1153 585
R7502 GNDA.n1151 GNDA.n910 585
R7503 GNDA.n1149 GNDA.n1148 585
R7504 GNDA.n1147 GNDA.n911 585
R7505 GNDA.n1146 GNDA.n1145 585
R7506 GNDA.n1143 GNDA.n912 585
R7507 GNDA.n1141 GNDA.n1140 585
R7508 GNDA.n1218 GNDA.n648 585
R7509 GNDA.n1216 GNDA.n1215 585
R7510 GNDA.n1214 GNDA.n649 585
R7511 GNDA.n1213 GNDA.n1212 585
R7512 GNDA.n1210 GNDA.n650 585
R7513 GNDA.n1208 GNDA.n1207 585
R7514 GNDA.n1206 GNDA.n651 585
R7515 GNDA.n1205 GNDA.n1204 585
R7516 GNDA.n1202 GNDA.n652 585
R7517 GNDA.n1200 GNDA.n1199 585
R7518 GNDA.n1198 GNDA.n653 585
R7519 GNDA.n1197 GNDA.n1196 585
R7520 GNDA.n6951 GNDA.n163 585
R7521 GNDA.n6951 GNDA.n162 585
R7522 GNDA.n7041 GNDA.n7040 585
R7523 GNDA.n7038 GNDA.n227 585
R7524 GNDA.n6928 GNDA.n6927 585
R7525 GNDA.n7033 GNDA.n7032 585
R7526 GNDA.n7031 GNDA.n7030 585
R7527 GNDA.n6957 GNDA.n6932 585
R7528 GNDA.n6959 GNDA.n6958 585
R7529 GNDA.n6964 GNDA.n6963 585
R7530 GNDA.n6962 GNDA.n6955 585
R7531 GNDA.n6970 GNDA.n6969 585
R7532 GNDA.n6972 GNDA.n6971 585
R7533 GNDA.n6953 GNDA.n6952 585
R7534 GNDA.n7113 GNDA.n163 585
R7535 GNDA.n7113 GNDA.n162 585
R7536 GNDA.n7112 GNDA.n7111 585
R7537 GNDA.n7109 GNDA.n7108 585
R7538 GNDA.n7107 GNDA.n7106 585
R7539 GNDA.n200 GNDA.n168 585
R7540 GNDA.n220 GNDA.n219 585
R7541 GNDA.n216 GNDA.n199 585
R7542 GNDA.n203 GNDA.n202 585
R7543 GNDA.n211 GNDA.n210 585
R7544 GNDA.n209 GNDA.n208 585
R7545 GNDA.n189 GNDA.n188 585
R7546 GNDA.n7046 GNDA.n7045 585
R7547 GNDA.n654 GNDA.n190 585
R7548 GNDA.n781 GNDA.n657 585
R7549 GNDA.n805 GNDA.n783 585
R7550 GNDA.n807 GNDA.n806 585
R7551 GNDA.n803 GNDA.n802 585
R7552 GNDA.n801 GNDA.n800 585
R7553 GNDA.n796 GNDA.n795 585
R7554 GNDA.n794 GNDA.n793 585
R7555 GNDA.n789 GNDA.n788 585
R7556 GNDA.n787 GNDA.n708 585
R7557 GNDA.n815 GNDA.n814 585
R7558 GNDA.n817 GNDA.n816 585
R7559 GNDA.n820 GNDA.n819 585
R7560 GNDA.n1335 GNDA.n640 585
R7561 GNDA.n1338 GNDA.n1337 585
R7562 GNDA.n1337 GNDA.n1336 585
R7563 GNDA.n639 GNDA.n638 585
R7564 GNDA.n1236 GNDA.n639 585
R7565 GNDA.n1234 GNDA.n1233 585
R7566 GNDA.n1235 GNDA.n1234 585
R7567 GNDA.n1232 GNDA.n642 585
R7568 GNDA.n642 GNDA.n641 585
R7569 GNDA.n1231 GNDA.n1230 585
R7570 GNDA.n1230 GNDA.n553 585
R7571 GNDA.n1229 GNDA.n643 585
R7572 GNDA.n1229 GNDA.n552 585
R7573 GNDA.n1228 GNDA.n645 585
R7574 GNDA.n1228 GNDA.n1227 585
R7575 GNDA.n1222 GNDA.n644 585
R7576 GNDA.n1226 GNDA.n644 585
R7577 GNDA.n1224 GNDA.n1223 585
R7578 GNDA.n1225 GNDA.n1224 585
R7579 GNDA.n1221 GNDA.n647 585
R7580 GNDA.n647 GNDA.n646 585
R7581 GNDA.n1220 GNDA.n1219 585
R7582 GNDA.n1219 GNDA.n102 585
R7583 GNDA.n1334 GNDA.n635 585
R7584 GNDA.n705 GNDA.n704 585
R7585 GNDA.n825 GNDA.n824 585
R7586 GNDA.n826 GNDA.n825 585
R7587 GNDA.n702 GNDA.n701 585
R7588 GNDA.n827 GNDA.n702 585
R7589 GNDA.n830 GNDA.n829 585
R7590 GNDA.n829 GNDA.n828 585
R7591 GNDA.n831 GNDA.n700 585
R7592 GNDA.n703 GNDA.n700 585
R7593 GNDA.n833 GNDA.n832 585
R7594 GNDA.n833 GNDA.n109 585
R7595 GNDA.n834 GNDA.n699 585
R7596 GNDA.n834 GNDA.n110 585
R7597 GNDA.n837 GNDA.n836 585
R7598 GNDA.n836 GNDA.n835 585
R7599 GNDA.n838 GNDA.n697 585
R7600 GNDA.n697 GNDA.n696 585
R7601 GNDA.n840 GNDA.n839 585
R7602 GNDA.n841 GNDA.n840 585
R7603 GNDA.n698 GNDA.n695 585
R7604 GNDA.n842 GNDA.n695 585
R7605 GNDA.n844 GNDA.n694 585
R7606 GNDA.n844 GNDA.n843 585
R7607 GNDA.n821 GNDA.n103 585
R7608 GNDA.n7154 GNDA.n7153 585
R7609 GNDA.n7156 GNDA.n88 585
R7610 GNDA.n7227 GNDA.n7226 585
R7611 GNDA.n24 GNDA.n22 585
R7612 GNDA.n7325 GNDA.n7324 585
R7613 GNDA.n32 GNDA.n25 585
R7614 GNDA.n40 GNDA.n39 585
R7615 GNDA.n35 GNDA.n31 585
R7616 GNDA.n30 GNDA.n0 585
R7617 GNDA.n7161 GNDA.n1 585
R7618 GNDA.n7163 GNDA.n7162 585
R7619 GNDA.n7167 GNDA.n7166 585
R7620 GNDA.n7169 GNDA.n7168 585
R7621 GNDA.n7158 GNDA.n7157 585
R7622 GNDA.n7148 GNDA.n89 585
R7623 GNDA.n7152 GNDA.n89 585
R7624 GNDA.n7150 GNDA.n7149 585
R7625 GNDA.n7151 GNDA.n7150 585
R7626 GNDA.n7147 GNDA.n91 585
R7627 GNDA.n91 GNDA.n90 585
R7628 GNDA.n7146 GNDA.n7145 585
R7629 GNDA.n7145 GNDA.n7144 585
R7630 GNDA.n93 GNDA.n92 585
R7631 GNDA.n7143 GNDA.n93 585
R7632 GNDA.n6691 GNDA.n6690 585
R7633 GNDA.n6690 GNDA.n111 585
R7634 GNDA.n6693 GNDA.n6692 585
R7635 GNDA.n6694 GNDA.n6693 585
R7636 GNDA.n6689 GNDA.n6688 585
R7637 GNDA.n6695 GNDA.n6689 585
R7638 GNDA.n6698 GNDA.n6697 585
R7639 GNDA.n6697 GNDA.n6696 585
R7640 GNDA.n6699 GNDA.n6687 585
R7641 GNDA.n6687 GNDA.n6686 585
R7642 GNDA.n6701 GNDA.n6700 585
R7643 GNDA.n6702 GNDA.n6701 585
R7644 GNDA.n6685 GNDA.n6684 585
R7645 GNDA.n6703 GNDA.n6685 585
R7646 GNDA.n6706 GNDA.n6705 585
R7647 GNDA.n6705 GNDA.n6704 585
R7648 GNDA.n6707 GNDA.n6683 585
R7649 GNDA.n6683 GNDA.n6682 585
R7650 GNDA.n6709 GNDA.n6708 585
R7651 GNDA.n6710 GNDA.n6709 585
R7652 GNDA.n6681 GNDA.n6680 585
R7653 GNDA.n6711 GNDA.n6681 585
R7654 GNDA.n6714 GNDA.n6713 585
R7655 GNDA.n6713 GNDA.n6712 585
R7656 GNDA.n6715 GNDA.n6679 585
R7657 GNDA.n6679 GNDA.n6678 585
R7658 GNDA.n6717 GNDA.n6716 585
R7659 GNDA.n6718 GNDA.n6717 585
R7660 GNDA.n6677 GNDA.n6676 585
R7661 GNDA.n6719 GNDA.n6677 585
R7662 GNDA.n6722 GNDA.n6721 585
R7663 GNDA.n6721 GNDA.n6720 585
R7664 GNDA.n6723 GNDA.n6675 585
R7665 GNDA.n6675 GNDA.n6629 585
R7666 GNDA.n6725 GNDA.n6724 585
R7667 GNDA.n6726 GNDA.n6725 585
R7668 GNDA.n6730 GNDA.n6729 585
R7669 GNDA.n6729 GNDA.n6728 585
R7670 GNDA.n6731 GNDA.n6625 585
R7671 GNDA.n6625 GNDA.n6624 585
R7672 GNDA.n6733 GNDA.n6732 585
R7673 GNDA.n6734 GNDA.n6733 585
R7674 GNDA.n6626 GNDA.n6623 585
R7675 GNDA.n6735 GNDA.n6623 585
R7676 GNDA.n6737 GNDA.n6622 585
R7677 GNDA.n6737 GNDA.n6736 585
R7678 GNDA.n6739 GNDA.n6738 585
R7679 GNDA.n6738 GNDA.n357 585
R7680 GNDA.n355 GNDA.n354 585
R7681 GNDA.n6745 GNDA.n355 585
R7682 GNDA.n6748 GNDA.n6747 585
R7683 GNDA.n6747 GNDA.n6746 585
R7684 GNDA.n6749 GNDA.n353 585
R7685 GNDA.n353 GNDA.n352 585
R7686 GNDA.n6751 GNDA.n6750 585
R7687 GNDA.n6752 GNDA.n6751 585
R7688 GNDA.n351 GNDA.n304 585
R7689 GNDA.n6753 GNDA.n351 585
R7690 GNDA.n6756 GNDA.n6755 585
R7691 GNDA.n6755 GNDA.n6754 585
R7692 GNDA.n6651 GNDA.n83 585
R7693 GNDA.n6652 GNDA.n6650 585
R7694 GNDA.n6657 GNDA.n6648 585
R7695 GNDA.n6658 GNDA.n6646 585
R7696 GNDA.n6659 GNDA.n6645 585
R7697 GNDA.n6643 GNDA.n6641 585
R7698 GNDA.n6665 GNDA.n6640 585
R7699 GNDA.n6666 GNDA.n6638 585
R7700 GNDA.n6667 GNDA.n6637 585
R7701 GNDA.n6635 GNDA.n6633 585
R7702 GNDA.n6672 GNDA.n6632 585
R7703 GNDA.n6673 GNDA.n6628 585
R7704 GNDA.n7230 GNDA.n84 585
R7705 GNDA.n7230 GNDA.n7229 585
R7706 GNDA.n6674 GNDA.n6673 585
R7707 GNDA.n6672 GNDA.n6671 585
R7708 GNDA.n6670 GNDA.n6633 585
R7709 GNDA.n6668 GNDA.n6667 585
R7710 GNDA.n6666 GNDA.n6634 585
R7711 GNDA.n6665 GNDA.n6664 585
R7712 GNDA.n6662 GNDA.n6641 585
R7713 GNDA.n6660 GNDA.n6659 585
R7714 GNDA.n6658 GNDA.n6642 585
R7715 GNDA.n6657 GNDA.n6656 585
R7716 GNDA.n6654 GNDA.n6652 585
R7717 GNDA.n6651 GNDA.n86 585
R7718 GNDA.n7228 GNDA.n84 585
R7719 GNDA.n7229 GNDA.n7228 585
R7720 GNDA.n901 GNDA.n900 585
R7721 GNDA.n898 GNDA.n659 585
R7722 GNDA.n897 GNDA.n896 585
R7723 GNDA.n888 GNDA.n661 585
R7724 GNDA.n890 GNDA.n889 585
R7725 GNDA.n886 GNDA.n663 585
R7726 GNDA.n885 GNDA.n884 585
R7727 GNDA.n876 GNDA.n665 585
R7728 GNDA.n878 GNDA.n877 585
R7729 GNDA.n874 GNDA.n667 585
R7730 GNDA.n873 GNDA.n872 585
R7731 GNDA.n690 GNDA.n669 585
R7732 GNDA.n904 GNDA.n656 585
R7733 GNDA.n656 GNDA.n162 585
R7734 GNDA.n869 GNDA.n669 585
R7735 GNDA.n872 GNDA.n871 585
R7736 GNDA.n667 GNDA.n666 585
R7737 GNDA.n666 GNDA.n112 585
R7738 GNDA.n879 GNDA.n878 585
R7739 GNDA.n881 GNDA.n665 585
R7740 GNDA.n884 GNDA.n883 585
R7741 GNDA.n663 GNDA.n662 585
R7742 GNDA.n891 GNDA.n890 585
R7743 GNDA.n893 GNDA.n661 585
R7744 GNDA.n896 GNDA.n895 585
R7745 GNDA.n659 GNDA.n658 585
R7746 GNDA.n902 GNDA.n901 585
R7747 GNDA.n902 GNDA.n112 585
R7748 GNDA.n904 GNDA.n903 585
R7749 GNDA.n903 GNDA.n162 585
R7750 GNDA.n6216 GNDA.n569 585
R7751 GNDA.n6219 GNDA.n6218 585
R7752 GNDA.n574 GNDA.n573 585
R7753 GNDA.n1178 GNDA.n1177 585
R7754 GNDA.n1179 GNDA.n1176 585
R7755 GNDA.n1173 GNDA.n1172 585
R7756 GNDA.n1185 GNDA.n1171 585
R7757 GNDA.n1186 GNDA.n1170 585
R7758 GNDA.n1187 GNDA.n1169 585
R7759 GNDA.n1167 GNDA.n1166 585
R7760 GNDA.n1192 GNDA.n1165 585
R7761 GNDA.n1193 GNDA.n1164 585
R7762 GNDA.n1194 GNDA.n1193 585
R7763 GNDA.n1192 GNDA.n1191 585
R7764 GNDA.n1190 GNDA.n1167 585
R7765 GNDA.n1188 GNDA.n1187 585
R7766 GNDA.n1186 GNDA.n1168 585
R7767 GNDA.n1185 GNDA.n1184 585
R7768 GNDA.n1182 GNDA.n1173 585
R7769 GNDA.n1180 GNDA.n1179 585
R7770 GNDA.n1178 GNDA.n1175 585
R7771 GNDA.n573 GNDA.n572 585
R7772 GNDA.n6220 GNDA.n6219 585
R7773 GNDA.n6222 GNDA.n569 585
R7774 GNDA.n960 GNDA.n959 585
R7775 GNDA.n950 GNDA.n949 585
R7776 GNDA.n962 GNDA.n949 585
R7777 GNDA.n954 GNDA.n953 585
R7778 GNDA.n6233 GNDA.n558 585
R7779 GNDA.n6237 GNDA.n557 585
R7780 GNDA.n6245 GNDA.n557 585
R7781 GNDA.n6236 GNDA.n6235 585
R7782 GNDA.n6205 GNDA.n584 585
R7783 GNDA.n6205 GNDA.n6204 585
R7784 GNDA.n1056 GNDA.n1055 585
R7785 GNDA.n1055 GNDA.n106 585
R7786 GNDA.n1054 GNDA.n924 585
R7787 GNDA.n1054 GNDA.n1053 585
R7788 GNDA.n1040 GNDA.n923 585
R7789 GNDA.n1052 GNDA.n923 585
R7790 GNDA.n1048 GNDA.n1047 585
R7791 GNDA.n1049 GNDA.n1048 585
R7792 GNDA.n930 GNDA.n928 585
R7793 GNDA.n928 GNDA.n927 585
R7794 GNDA.n966 GNDA.n963 585
R7795 GNDA.n963 GNDA.n107 585
R7796 GNDA.n974 GNDA.n973 585
R7797 GNDA.n975 GNDA.n974 585
R7798 GNDA.n964 GNDA.n947 585
R7799 GNDA.n976 GNDA.n947 585
R7800 GNDA.n980 GNDA.n979 585
R7801 GNDA.n979 GNDA.n978 585
R7802 GNDA.n981 GNDA.n592 585
R7803 GNDA.n977 GNDA.n592 585
R7804 GNDA.n6201 GNDA.n6200 585
R7805 GNDA.n6202 GNDA.n6201 585
R7806 GNDA.n6198 GNDA.n591 585
R7807 GNDA.n6203 GNDA.n591 585
R7808 GNDA.n6224 GNDA.n566 585
R7809 GNDA.n580 GNDA.n566 585
R7810 GNDA.n6213 GNDA.n584 585
R7811 GNDA.n6214 GNDA.n6213 585
R7812 GNDA.n6196 GNDA.n586 585
R7813 GNDA.n586 GNDA.n585 585
R7814 GNDA.n6194 GNDA.n6193 585
R7815 GNDA.n6193 GNDA.n6192 585
R7816 GNDA.n601 GNDA.n597 585
R7817 GNDA.n6191 GNDA.n597 585
R7818 GNDA.n6189 GNDA.n6188 585
R7819 GNDA.n6190 GNDA.n6189 585
R7820 GNDA.n603 GNDA.n600 585
R7821 GNDA.n6107 GNDA.n600 585
R7822 GNDA.n6110 GNDA.n6109 585
R7823 GNDA.n6109 GNDA.n6108 585
R7824 GNDA.n6111 GNDA.n6105 585
R7825 GNDA.n6105 GNDA.n6104 585
R7826 GNDA.n6120 GNDA.n6119 585
R7827 GNDA.n6121 GNDA.n6120 585
R7828 GNDA.n624 GNDA.n623 585
R7829 GNDA.n6122 GNDA.n624 585
R7830 GNDA.n6126 GNDA.n6125 585
R7831 GNDA.n6125 GNDA.n6124 585
R7832 GNDA.n620 GNDA.n565 585
R7833 GNDA.n6123 GNDA.n565 585
R7834 GNDA.n6227 GNDA.n6226 585
R7835 GNDA.n6228 GNDA.n6227 585
R7836 GNDA.n6224 GNDA.n6223 585
R7837 GNDA.n6223 GNDA.n570 585
R7838 GNDA.n571 GNDA.n568 585
R7839 GNDA.n1237 GNDA.n571 585
R7840 GNDA.n1307 GNDA.n1239 585
R7841 GNDA.n1239 GNDA.n1238 585
R7842 GNDA.n1330 GNDA.n1329 585
R7843 GNDA.n1331 GNDA.n1330 585
R7844 GNDA.n1242 GNDA.n1240 585
R7845 GNDA.n1320 GNDA.n1240 585
R7846 GNDA.n1323 GNDA.n1322 585
R7847 GNDA.n1322 GNDA.n1321 585
R7848 GNDA.n1319 GNDA.n1318 585
R7849 GNDA.n1319 GNDA.n555 585
R7850 GNDA.n1316 GNDA.n551 585
R7851 GNDA.n6246 GNDA.n551 585
R7852 GNDA.n6249 GNDA.n6248 585
R7853 GNDA.n6248 GNDA.n6247 585
R7854 GNDA.n548 GNDA.n543 585
R7855 GNDA.n543 GNDA.n541 585
R7856 GNDA.n6259 GNDA.n6258 585
R7857 GNDA.n6260 GNDA.n6259 585
R7858 GNDA.n546 GNDA.n544 585
R7859 GNDA.n544 GNDA.n542 585
R7860 GNDA.n1341 GNDA.n1340 585
R7861 GNDA.n1342 GNDA.n1341 585
R7862 GNDA.n1079 GNDA.n1078 585
R7863 GNDA.n1077 GNDA.n1076 585
R7864 GNDA.n1075 GNDA.n1074 585
R7865 GNDA.n1073 GNDA.n1072 585
R7866 GNDA.n1071 GNDA.n1070 585
R7867 GNDA.n1069 GNDA.n1068 585
R7868 GNDA.n1067 GNDA.n1066 585
R7869 GNDA.n1065 GNDA.n1064 585
R7870 GNDA.n1063 GNDA.n1062 585
R7871 GNDA.n1061 GNDA.n1060 585
R7872 GNDA.n1059 GNDA.n1058 585
R7873 GNDA.n6922 GNDA.n281 585
R7874 GNDA.n263 GNDA.n262 585
R7875 GNDA.n265 GNDA.n264 585
R7876 GNDA.n267 GNDA.n266 585
R7877 GNDA.n269 GNDA.n268 585
R7878 GNDA.n271 GNDA.n270 585
R7879 GNDA.n273 GNDA.n272 585
R7880 GNDA.n275 GNDA.n274 585
R7881 GNDA.n276 GNDA.n241 585
R7882 GNDA.n279 GNDA.n278 585
R7883 GNDA.n277 GNDA.n240 585
R7884 GNDA.n230 GNDA.n229 585
R7885 GNDA.n6922 GNDA.n230 585
R7886 GNDA.n6925 GNDA.n6924 585
R7887 GNDA.n6925 GNDA.n228 585
R7888 GNDA.n6920 GNDA.n6919 585
R7889 GNDA.n6918 GNDA.n289 585
R7890 GNDA.n6917 GNDA.n288 585
R7891 GNDA.n6922 GNDA.n288 585
R7892 GNDA.n6916 GNDA.n6915 585
R7893 GNDA.n6914 GNDA.n6913 585
R7894 GNDA.n6912 GNDA.n6911 585
R7895 GNDA.n6910 GNDA.n6909 585
R7896 GNDA.n6908 GNDA.n6907 585
R7897 GNDA.n6906 GNDA.n6905 585
R7898 GNDA.n6904 GNDA.n6903 585
R7899 GNDA.n6902 GNDA.n6901 585
R7900 GNDA.n6900 GNDA.n6899 585
R7901 GNDA.n6899 GNDA.n6898 585
R7902 GNDA.n1366 GNDA.t805 524.808
R7903 GNDA.n4801 GNDA.t822 524.808
R7904 GNDA.n4085 GNDA.t761 524.808
R7905 GNDA.n3462 GNDA.t802 524.808
R7906 GNDA.n4116 GNDA.t748 508.743
R7907 GNDA.n4113 GNDA.t755 508.743
R7908 GNDA.n4782 GNDA.t739 508.743
R7909 GNDA.n4127 GNDA.t831 508.743
R7910 GNDA.n4109 GNDA.t758 499.442
R7911 GNDA.n4112 GNDA.t771 499.442
R7912 GNDA.n4793 GNDA.t815 499.442
R7913 GNDA.n4088 GNDA.t796 499.442
R7914 GNDA.n4789 GNDA.t790 475.976
R7915 GNDA.n4789 GNDA.t769 475.976
R7916 GNDA.n4132 GNDA.t812 475.976
R7917 GNDA.n4132 GNDA.t783 475.976
R7918 GNDA.n1334 GNDA.n1333 466.925
R7919 GNDA.n527 GNDA.t808 425.134
R7920 GNDA.n524 GNDA.t842 409.067
R7921 GNDA.n6263 GNDA.t774 409.067
R7922 GNDA.n537 GNDA.t825 409.067
R7923 GNDA.n536 GNDA.t780 409.067
R7924 GNDA.n533 GNDA.t828 409.067
R7925 GNDA.n532 GNDA.t787 409.067
R7926 GNDA.n528 GNDA.t777 409.067
R7927 GNDA.n1332 GNDA.t63 377.332
R7928 GNDA.n301 GNDA.n96 370.214
R7929 GNDA.n6727 GNDA.n98 370.214
R7930 GNDA.n301 GNDA.n95 365.957
R7931 GNDA.n6727 GNDA.n97 365.957
R7932 GNDA.n4091 GNDA.n4090 344.954
R7933 GNDA.n4798 GNDA.n4795 344.954
R7934 GNDA.t743 GNDA.n94 172.876
R7935 GNDA.t743 GNDA.n95 327.661
R7936 GNDA.t743 GNDA.n97 327.661
R7937 GNDA.n6215 GNDA.t743 172.876
R7938 GNDA.n581 GNDA.t743 172.615
R7939 GNDA.t743 GNDA.n96 323.404
R7940 GNDA.t743 GNDA.n98 323.404
R7941 GNDA.t743 GNDA.n554 172.615
R7942 GNDA.n4118 GNDA.n4117 296.158
R7943 GNDA.n4126 GNDA.n1815 296.158
R7944 GNDA.n4784 GNDA.n4783 296.158
R7945 GNDA.n4129 GNDA.n4128 296.158
R7946 GNDA.n4108 GNDA.n4107 292.5
R7947 GNDA.n4111 GNDA.n1347 292.5
R7948 GNDA.n4090 GNDA.n4089 292.5
R7949 GNDA.n4137 GNDA.n4136 292.5
R7950 GNDA.n4786 GNDA.n4785 292.5
R7951 GNDA.n4795 GNDA.n4794 292.5
R7952 GNDA.n4118 GNDA.t749 277.57
R7953 GNDA.n4118 GNDA.t794 277.57
R7954 GNDA.t753 GNDA.n4126 277.57
R7955 GNDA.n4126 GNDA.t756 277.57
R7956 GNDA.n1339 GNDA.n637 264.301
R7957 GNDA.n823 GNDA.n822 264.301
R7958 GNDA.n7155 GNDA.n87 264.301
R7959 GNDA.n1057 GNDA.n921 264.301
R7960 GNDA.n6923 GNDA.n6922 264.301
R7961 GNDA.n6922 GNDA.n235 264.301
R7962 GNDA.n1219 GNDA.n1218 259.416
R7963 GNDA.n1164 GNDA.n1163 259.416
R7964 GNDA.n1137 GNDA.n1136 259.416
R7965 GNDA.n6729 GNDA.n6628 259.416
R7966 GNDA.n845 GNDA.n844 259.416
R7967 GNDA.n691 GNDA.n690 259.416
R7968 GNDA.n7140 GNDA.n131 259.416
R7969 GNDA.n6759 GNDA.n302 259.416
R7970 GNDA.n6701 GNDA.n6685 259.416
R7971 GNDA.n1292 GNDA.n1247 258.334
R7972 GNDA.n6166 GNDA.n6164 258.334
R7973 GNDA.n7085 GNDA.n7084 258.334
R7974 GNDA.n6870 GNDA.n6869 258.334
R7975 GNDA.n764 GNDA.n763 258.334
R7976 GNDA.n7009 GNDA.n6949 258.334
R7977 GNDA.n7288 GNDA.n80 258.334
R7978 GNDA.n1022 GNDA.n936 258.334
R7979 GNDA.n7208 GNDA.n7207 258.334
R7980 GNDA.n4106 GNDA.t759 257.01
R7981 GNDA.t772 GNDA.n1346 257.01
R7982 GNDA.n7142 GNDA.n7141 254.34
R7983 GNDA.n7142 GNDA.n129 254.34
R7984 GNDA.n7142 GNDA.n128 254.34
R7985 GNDA.n7142 GNDA.n127 254.34
R7986 GNDA.n7142 GNDA.n126 254.34
R7987 GNDA.n7142 GNDA.n125 254.34
R7988 GNDA.n7142 GNDA.n124 254.34
R7989 GNDA.n7142 GNDA.n123 254.34
R7990 GNDA.n7142 GNDA.n122 254.34
R7991 GNDA.n7142 GNDA.n121 254.34
R7992 GNDA.n7142 GNDA.n120 254.34
R7993 GNDA.n7142 GNDA.n119 254.34
R7994 GNDA.n7142 GNDA.n118 254.34
R7995 GNDA.n7142 GNDA.n117 254.34
R7996 GNDA.n7142 GNDA.n116 254.34
R7997 GNDA.n7142 GNDA.n115 254.34
R7998 GNDA.n7142 GNDA.n114 254.34
R7999 GNDA.n7142 GNDA.n113 254.34
R8000 GNDA.n7322 GNDA.n7321 254.34
R8001 GNDA.n7322 GNDA.n53 254.34
R8002 GNDA.n7322 GNDA.n52 254.34
R8003 GNDA.n7322 GNDA.n51 254.34
R8004 GNDA.n7322 GNDA.n50 254.34
R8005 GNDA.n7322 GNDA.n49 254.34
R8006 GNDA.n7322 GNDA.n48 254.34
R8007 GNDA.n7322 GNDA.n47 254.34
R8008 GNDA.n7322 GNDA.n46 254.34
R8009 GNDA.n7322 GNDA.n45 254.34
R8010 GNDA.n7322 GNDA.n44 254.34
R8011 GNDA.n7322 GNDA.n43 254.34
R8012 GNDA.n325 GNDA.n95 254.34
R8013 GNDA.n322 GNDA.n95 254.34
R8014 GNDA.n317 GNDA.n95 254.34
R8015 GNDA.n314 GNDA.n95 254.34
R8016 GNDA.n309 GNDA.n95 254.34
R8017 GNDA.n306 GNDA.n95 254.34
R8018 GNDA.n349 GNDA.n96 254.34
R8019 GNDA.n343 GNDA.n96 254.34
R8020 GNDA.n341 GNDA.n96 254.34
R8021 GNDA.n335 GNDA.n96 254.34
R8022 GNDA.n333 GNDA.n96 254.34
R8023 GNDA.n327 GNDA.n96 254.34
R8024 GNDA.n159 GNDA.n158 254.34
R8025 GNDA.n158 GNDA.n157 254.34
R8026 GNDA.n158 GNDA.n156 254.34
R8027 GNDA.n158 GNDA.n155 254.34
R8028 GNDA.n158 GNDA.n154 254.34
R8029 GNDA.n158 GNDA.n153 254.34
R8030 GNDA.n7135 GNDA.n7134 254.34
R8031 GNDA.n7134 GNDA.n7133 254.34
R8032 GNDA.n7134 GNDA.n141 254.34
R8033 GNDA.n7134 GNDA.n140 254.34
R8034 GNDA.n7134 GNDA.n139 254.34
R8035 GNDA.n7134 GNDA.n138 254.34
R8036 GNDA.n6207 GNDA.n94 254.34
R8037 GNDA.n1116 GNDA.n94 254.34
R8038 GNDA.n1114 GNDA.n94 254.34
R8039 GNDA.n1108 GNDA.n94 254.34
R8040 GNDA.n1105 GNDA.n94 254.34
R8041 GNDA.n1135 GNDA.n94 254.34
R8042 GNDA.n1131 GNDA.n581 254.34
R8043 GNDA.n1129 GNDA.n581 254.34
R8044 GNDA.n1123 GNDA.n581 254.34
R8045 GNDA.n1121 GNDA.n581 254.34
R8046 GNDA.n1111 GNDA.n581 254.34
R8047 GNDA.n6211 GNDA.n581 254.34
R8048 GNDA.n1101 GNDA.n104 254.34
R8049 GNDA.n916 GNDA.n104 254.34
R8050 GNDA.n1094 GNDA.n104 254.34
R8051 GNDA.n1088 GNDA.n104 254.34
R8052 GNDA.n1086 GNDA.n104 254.34
R8053 GNDA.n1080 GNDA.n104 254.34
R8054 GNDA.n907 GNDA.n104 254.34
R8055 GNDA.n1158 GNDA.n104 254.34
R8056 GNDA.n1152 GNDA.n104 254.34
R8057 GNDA.n1150 GNDA.n104 254.34
R8058 GNDA.n1144 GNDA.n104 254.34
R8059 GNDA.n1142 GNDA.n104 254.34
R8060 GNDA.n1217 GNDA.n104 254.34
R8061 GNDA.n1211 GNDA.n104 254.34
R8062 GNDA.n1209 GNDA.n104 254.34
R8063 GNDA.n1203 GNDA.n104 254.34
R8064 GNDA.n1201 GNDA.n104 254.34
R8065 GNDA.n1195 GNDA.n104 254.34
R8066 GNDA.n7043 GNDA.n7042 254.34
R8067 GNDA.n7043 GNDA.n226 254.34
R8068 GNDA.n7043 GNDA.n225 254.34
R8069 GNDA.n7043 GNDA.n224 254.34
R8070 GNDA.n7043 GNDA.n223 254.34
R8071 GNDA.n7043 GNDA.n222 254.34
R8072 GNDA.n7043 GNDA.n164 254.34
R8073 GNDA.n7043 GNDA.n167 254.34
R8074 GNDA.n7043 GNDA.n221 254.34
R8075 GNDA.n7043 GNDA.n198 254.34
R8076 GNDA.n7043 GNDA.n197 254.34
R8077 GNDA.n7044 GNDA.n7043 254.34
R8078 GNDA.n7043 GNDA.n196 254.34
R8079 GNDA.n7043 GNDA.n195 254.34
R8080 GNDA.n7043 GNDA.n194 254.34
R8081 GNDA.n7043 GNDA.n193 254.34
R8082 GNDA.n7043 GNDA.n192 254.34
R8083 GNDA.n7043 GNDA.n191 254.34
R8084 GNDA.n7322 GNDA.n42 254.34
R8085 GNDA.n7323 GNDA.n7322 254.34
R8086 GNDA.n7322 GNDA.n41 254.34
R8087 GNDA.n7322 GNDA.n29 254.34
R8088 GNDA.n7322 GNDA.n28 254.34
R8089 GNDA.n7322 GNDA.n27 254.34
R8090 GNDA.n6649 GNDA.n97 254.34
R8091 GNDA.n6647 GNDA.n97 254.34
R8092 GNDA.n6644 GNDA.n97 254.34
R8093 GNDA.n6639 GNDA.n97 254.34
R8094 GNDA.n6636 GNDA.n97 254.34
R8095 GNDA.n6631 GNDA.n97 254.34
R8096 GNDA.n6630 GNDA.n98 254.34
R8097 GNDA.n6669 GNDA.n98 254.34
R8098 GNDA.n6663 GNDA.n98 254.34
R8099 GNDA.n6661 GNDA.n98 254.34
R8100 GNDA.n6655 GNDA.n98 254.34
R8101 GNDA.n6653 GNDA.n98 254.34
R8102 GNDA.n899 GNDA.n101 254.34
R8103 GNDA.n660 GNDA.n101 254.34
R8104 GNDA.n887 GNDA.n101 254.34
R8105 GNDA.n664 GNDA.n101 254.34
R8106 GNDA.n875 GNDA.n101 254.34
R8107 GNDA.n668 GNDA.n101 254.34
R8108 GNDA.n870 GNDA.n112 254.34
R8109 GNDA.n880 GNDA.n112 254.34
R8110 GNDA.n882 GNDA.n112 254.34
R8111 GNDA.n892 GNDA.n112 254.34
R8112 GNDA.n894 GNDA.n112 254.34
R8113 GNDA.n6217 GNDA.n6215 254.34
R8114 GNDA.n6215 GNDA.n579 254.34
R8115 GNDA.n6215 GNDA.n578 254.34
R8116 GNDA.n6215 GNDA.n577 254.34
R8117 GNDA.n6215 GNDA.n576 254.34
R8118 GNDA.n6215 GNDA.n575 254.34
R8119 GNDA.n906 GNDA.n554 254.34
R8120 GNDA.n1189 GNDA.n554 254.34
R8121 GNDA.n1183 GNDA.n554 254.34
R8122 GNDA.n1181 GNDA.n554 254.34
R8123 GNDA.n1174 GNDA.n554 254.34
R8124 GNDA.n6221 GNDA.n554 254.34
R8125 GNDA.n6922 GNDA.n287 254.34
R8126 GNDA.n6922 GNDA.n286 254.34
R8127 GNDA.n6922 GNDA.n285 254.34
R8128 GNDA.n6922 GNDA.n284 254.34
R8129 GNDA.n6922 GNDA.n283 254.34
R8130 GNDA.n6922 GNDA.n282 254.34
R8131 GNDA.n6922 GNDA.n236 254.34
R8132 GNDA.n6922 GNDA.n237 254.34
R8133 GNDA.n6922 GNDA.n238 254.34
R8134 GNDA.n6922 GNDA.n239 254.34
R8135 GNDA.n6922 GNDA.n280 254.34
R8136 GNDA.n6922 GNDA.n6921 254.34
R8137 GNDA.n6922 GNDA.n231 254.34
R8138 GNDA.n6922 GNDA.n232 254.34
R8139 GNDA.n6922 GNDA.n233 254.34
R8140 GNDA.n6922 GNDA.n234 254.34
R8141 GNDA.t743 GNDA.n6744 250.349
R8142 GNDA.n1196 GNDA.n1194 249.663
R8143 GNDA.n1141 GNDA.n913 249.663
R8144 GNDA.n1081 GNDA.n1079 249.663
R8145 GNDA.n6755 GNDA.n350 249.663
R8146 GNDA.n869 GNDA.n868 249.663
R8147 GNDA.n7136 GNDA.n136 249.663
R8148 GNDA.n262 GNDA.n261 249.663
R8149 GNDA.n6920 GNDA.n290 249.663
R8150 GNDA.n6725 GNDA.n6674 249.663
R8151 GNDA.n558 GNDA.n557 246.25
R8152 GNDA.n6235 GNDA.n557 246.25
R8153 GNDA.n960 GNDA.n949 246.25
R8154 GNDA.n953 GNDA.n949 246.25
R8155 GNDA.n962 GNDA.n961 241.643
R8156 GNDA.n962 GNDA.n948 241.643
R8157 GNDA.n6245 GNDA.n6244 241.643
R8158 GNDA.n6245 GNDA.n556 241.643
R8159 GNDA.t759 GNDA.t3 226.168
R8160 GNDA.t3 GNDA.t141 226.168
R8161 GNDA.t141 GNDA.t2 226.168
R8162 GNDA.t2 GNDA.t82 226.168
R8163 GNDA.t82 GNDA.t86 226.168
R8164 GNDA.t86 GNDA.t15 226.168
R8165 GNDA.t15 GNDA.t85 226.168
R8166 GNDA.t85 GNDA.t22 226.168
R8167 GNDA.t22 GNDA.t865 226.168
R8168 GNDA.t865 GNDA.t23 226.168
R8169 GNDA.t23 GNDA.t749 226.168
R8170 GNDA.t794 GNDA.t868 226.168
R8171 GNDA.t94 GNDA.t753 226.168
R8172 GNDA.t756 GNDA.t4 226.168
R8173 GNDA.t4 GNDA.t866 226.168
R8174 GNDA.t866 GNDA.t73 226.168
R8175 GNDA.t73 GNDA.t83 226.168
R8176 GNDA.t83 GNDA.t72 226.168
R8177 GNDA.t72 GNDA.t42 226.168
R8178 GNDA.t42 GNDA.t21 226.168
R8179 GNDA.t21 GNDA.t140 226.168
R8180 GNDA.t140 GNDA.t1 226.168
R8181 GNDA.t1 GNDA.t14 226.168
R8182 GNDA.t14 GNDA.t772 226.168
R8183 GNDA.t743 GNDA.t25 199.179
R8184 GNDA.n4139 GNDA.n4138 197.133
R8185 GNDA.n1594 GNDA.n1593 197.133
R8186 GNDA.n4119 GNDA.n4118 197.133
R8187 GNDA.n4126 GNDA.n4125 197.133
R8188 GNDA.n1341 GNDA.n635 197
R8189 GNDA.n6227 GNDA.n566 197
R8190 GNDA.n6205 GNDA.n591 197
R8191 GNDA.n821 GNDA.n820 197
R8192 GNDA.n656 GNDA.n190 197
R8193 GNDA.n6952 GNDA.n6951 197
R8194 GNDA.n6743 GNDA.n356 197
R8195 GNDA.n6803 GNDA.n85 197
R8196 GNDA.n7231 GNDA.n7230 197
R8197 GNDA.n7157 GNDA.n7156 197
R8198 GNDA.n6223 GNDA.n571 187.249
R8199 GNDA.n6213 GNDA.n586 187.249
R8200 GNDA.n1055 GNDA.n281 187.249
R8201 GNDA.n903 GNDA.n657 187.249
R8202 GNDA.n7113 GNDA.n7112 187.249
R8203 GNDA.n7041 GNDA.n228 187.249
R8204 GNDA.n6898 GNDA.n6897 187.249
R8205 GNDA.n7320 GNDA.n55 187.249
R8206 GNDA.n7228 GNDA.n7227 187.249
R8207 GNDA.n6243 GNDA.n6242 185
R8208 GNDA.n6240 GNDA.n6239 185
R8209 GNDA.n957 GNDA.n559 185
R8210 GNDA.n957 GNDA.n950 185
R8211 GNDA.n951 GNDA.n559 185
R8212 GNDA.n955 GNDA.n951 185
R8213 GNDA.n1292 GNDA.n1291 185
R8214 GNDA.n1294 GNDA.n1246 185
R8215 GNDA.n1297 GNDA.n1296 185
R8216 GNDA.n1298 GNDA.n1245 185
R8217 GNDA.n1300 GNDA.n1299 185
R8218 GNDA.n1302 GNDA.n1244 185
R8219 GNDA.n1305 GNDA.n1304 185
R8220 GNDA.n1306 GNDA.n1243 185
R8221 GNDA.n1310 GNDA.n1309 185
R8222 GNDA.n1274 GNDA.n1251 185
R8223 GNDA.n1276 GNDA.n1275 185
R8224 GNDA.n1278 GNDA.n1250 185
R8225 GNDA.n1281 GNDA.n1280 185
R8226 GNDA.n1282 GNDA.n1249 185
R8227 GNDA.n1284 GNDA.n1283 185
R8228 GNDA.n1286 GNDA.n1248 185
R8229 GNDA.n1289 GNDA.n1288 185
R8230 GNDA.n1290 GNDA.n1247 185
R8231 GNDA.n1258 GNDA.n547 185
R8232 GNDA.n1259 GNDA.n1257 185
R8233 GNDA.n1261 GNDA.n1260 185
R8234 GNDA.n1263 GNDA.n1254 185
R8235 GNDA.n1265 GNDA.n1264 185
R8236 GNDA.n1266 GNDA.n1253 185
R8237 GNDA.n1268 GNDA.n1267 185
R8238 GNDA.n1270 GNDA.n1252 185
R8239 GNDA.n1273 GNDA.n1272 185
R8240 GNDA.n6257 GNDA.n6256 185
R8241 GNDA.n6254 GNDA.n545 185
R8242 GNDA.n6253 GNDA.n549 185
R8243 GNDA.n6251 GNDA.n6250 185
R8244 GNDA.n1317 GNDA.n550 185
R8245 GNDA.n1315 GNDA.n1314 185
R8246 GNDA.n1325 GNDA.n1324 185
R8247 GNDA.n1328 GNDA.n1327 185
R8248 GNDA.n1312 GNDA.n1241 185
R8249 GNDA.n6167 GNDA.n6166 185
R8250 GNDA.n6168 GNDA.n608 185
R8251 GNDA.n6170 GNDA.n6169 185
R8252 GNDA.n6172 GNDA.n607 185
R8253 GNDA.n6175 GNDA.n6174 185
R8254 GNDA.n6176 GNDA.n606 185
R8255 GNDA.n6178 GNDA.n6177 185
R8256 GNDA.n6180 GNDA.n605 185
R8257 GNDA.n6181 GNDA.n595 185
R8258 GNDA.n6148 GNDA.n613 185
R8259 GNDA.n6151 GNDA.n6150 185
R8260 GNDA.n6152 GNDA.n612 185
R8261 GNDA.n6154 GNDA.n6153 185
R8262 GNDA.n6156 GNDA.n611 185
R8263 GNDA.n6159 GNDA.n6158 185
R8264 GNDA.n6160 GNDA.n610 185
R8265 GNDA.n6162 GNDA.n6161 185
R8266 GNDA.n6164 GNDA.n609 185
R8267 GNDA.n6132 GNDA.n6131 185
R8268 GNDA.n6134 GNDA.n618 185
R8269 GNDA.n6136 GNDA.n6135 185
R8270 GNDA.n6137 GNDA.n617 185
R8271 GNDA.n6139 GNDA.n6138 185
R8272 GNDA.n6141 GNDA.n615 185
R8273 GNDA.n6143 GNDA.n6142 185
R8274 GNDA.n6144 GNDA.n614 185
R8275 GNDA.n6146 GNDA.n6145 185
R8276 GNDA.n6130 GNDA.n621 185
R8277 GNDA.n6128 GNDA.n6127 185
R8278 GNDA.n6118 GNDA.n622 185
R8279 GNDA.n6117 GNDA.n6116 185
R8280 GNDA.n6114 GNDA.n6112 185
R8281 GNDA.n6106 GNDA.n604 185
R8282 GNDA.n6187 GNDA.n6186 185
R8283 GNDA.n6184 GNDA.n602 185
R8284 GNDA.n6183 GNDA.n596 185
R8285 GNDA.n7086 GNDA.n7085 185
R8286 GNDA.n7088 GNDA.n7087 185
R8287 GNDA.n7090 GNDA.n7089 185
R8288 GNDA.n7092 GNDA.n7091 185
R8289 GNDA.n7094 GNDA.n7093 185
R8290 GNDA.n7096 GNDA.n7095 185
R8291 GNDA.n7098 GNDA.n7097 185
R8292 GNDA.n7100 GNDA.n7099 185
R8293 GNDA.n7101 GNDA.n165 185
R8294 GNDA.n7068 GNDA.n7067 185
R8295 GNDA.n7070 GNDA.n7069 185
R8296 GNDA.n7072 GNDA.n7071 185
R8297 GNDA.n7074 GNDA.n7073 185
R8298 GNDA.n7076 GNDA.n7075 185
R8299 GNDA.n7078 GNDA.n7077 185
R8300 GNDA.n7080 GNDA.n7079 185
R8301 GNDA.n7082 GNDA.n7081 185
R8302 GNDA.n7084 GNDA.n7083 185
R8303 GNDA.n7050 GNDA.n7049 185
R8304 GNDA.n7052 GNDA.n7051 185
R8305 GNDA.n7054 GNDA.n7053 185
R8306 GNDA.n7056 GNDA.n7055 185
R8307 GNDA.n7058 GNDA.n7057 185
R8308 GNDA.n7060 GNDA.n7059 185
R8309 GNDA.n7062 GNDA.n7061 185
R8310 GNDA.n7064 GNDA.n7063 185
R8311 GNDA.n7066 GNDA.n7065 185
R8312 GNDA.n7048 GNDA.n7047 185
R8313 GNDA.n207 GNDA.n206 185
R8314 GNDA.n205 GNDA.n204 185
R8315 GNDA.n213 GNDA.n212 185
R8316 GNDA.n215 GNDA.n214 185
R8317 GNDA.n218 GNDA.n217 185
R8318 GNDA.n201 GNDA.n170 185
R8319 GNDA.n7105 GNDA.n7104 185
R8320 GNDA.n169 GNDA.n166 185
R8321 GNDA.n6871 GNDA.n6870 185
R8322 GNDA.n6873 GNDA.n6872 185
R8323 GNDA.n6875 GNDA.n6874 185
R8324 GNDA.n6877 GNDA.n6876 185
R8325 GNDA.n6879 GNDA.n6878 185
R8326 GNDA.n6881 GNDA.n6880 185
R8327 GNDA.n6883 GNDA.n6882 185
R8328 GNDA.n6885 GNDA.n6884 185
R8329 GNDA.n6886 GNDA.n6782 185
R8330 GNDA.n6853 GNDA.n6852 185
R8331 GNDA.n6855 GNDA.n6854 185
R8332 GNDA.n6857 GNDA.n6856 185
R8333 GNDA.n6859 GNDA.n6858 185
R8334 GNDA.n6861 GNDA.n6860 185
R8335 GNDA.n6863 GNDA.n6862 185
R8336 GNDA.n6865 GNDA.n6864 185
R8337 GNDA.n6867 GNDA.n6866 185
R8338 GNDA.n6869 GNDA.n6868 185
R8339 GNDA.n6835 GNDA.n6834 185
R8340 GNDA.n6837 GNDA.n6836 185
R8341 GNDA.n6839 GNDA.n6838 185
R8342 GNDA.n6841 GNDA.n6840 185
R8343 GNDA.n6843 GNDA.n6842 185
R8344 GNDA.n6845 GNDA.n6844 185
R8345 GNDA.n6847 GNDA.n6846 185
R8346 GNDA.n6849 GNDA.n6848 185
R8347 GNDA.n6851 GNDA.n6850 185
R8348 GNDA.n765 GNDA.n764 185
R8349 GNDA.n767 GNDA.n766 185
R8350 GNDA.n769 GNDA.n768 185
R8351 GNDA.n771 GNDA.n770 185
R8352 GNDA.n773 GNDA.n772 185
R8353 GNDA.n775 GNDA.n774 185
R8354 GNDA.n777 GNDA.n776 185
R8355 GNDA.n779 GNDA.n778 185
R8356 GNDA.n780 GNDA.n728 185
R8357 GNDA.n747 GNDA.n746 185
R8358 GNDA.n749 GNDA.n748 185
R8359 GNDA.n751 GNDA.n750 185
R8360 GNDA.n753 GNDA.n752 185
R8361 GNDA.n755 GNDA.n754 185
R8362 GNDA.n757 GNDA.n756 185
R8363 GNDA.n759 GNDA.n758 185
R8364 GNDA.n761 GNDA.n760 185
R8365 GNDA.n763 GNDA.n762 185
R8366 GNDA.n720 GNDA.n706 185
R8367 GNDA.n731 GNDA.n730 185
R8368 GNDA.n733 GNDA.n732 185
R8369 GNDA.n735 GNDA.n734 185
R8370 GNDA.n737 GNDA.n736 185
R8371 GNDA.n739 GNDA.n738 185
R8372 GNDA.n741 GNDA.n740 185
R8373 GNDA.n743 GNDA.n742 185
R8374 GNDA.n745 GNDA.n744 185
R8375 GNDA.n710 GNDA.n707 185
R8376 GNDA.n813 GNDA.n812 185
R8377 GNDA.n786 GNDA.n709 185
R8378 GNDA.n792 GNDA.n791 185
R8379 GNDA.n790 GNDA.n785 185
R8380 GNDA.n799 GNDA.n798 185
R8381 GNDA.n797 GNDA.n784 185
R8382 GNDA.n804 GNDA.n729 185
R8383 GNDA.n809 GNDA.n808 185
R8384 GNDA.n7011 GNDA.n6949 185
R8385 GNDA.n7025 GNDA.n7024 185
R8386 GNDA.n7023 GNDA.n6950 185
R8387 GNDA.n7022 GNDA.n7021 185
R8388 GNDA.n7020 GNDA.n7019 185
R8389 GNDA.n7018 GNDA.n7017 185
R8390 GNDA.n7016 GNDA.n7015 185
R8391 GNDA.n7014 GNDA.n7013 185
R8392 GNDA.n7012 GNDA.n6926 185
R8393 GNDA.n6994 GNDA.n6993 185
R8394 GNDA.n6996 GNDA.n6995 185
R8395 GNDA.n6998 GNDA.n6997 185
R8396 GNDA.n7000 GNDA.n6999 185
R8397 GNDA.n7002 GNDA.n7001 185
R8398 GNDA.n7004 GNDA.n7003 185
R8399 GNDA.n7006 GNDA.n7005 185
R8400 GNDA.n7008 GNDA.n7007 185
R8401 GNDA.n7010 GNDA.n7009 185
R8402 GNDA.n6976 GNDA.n6975 185
R8403 GNDA.n6978 GNDA.n6977 185
R8404 GNDA.n6980 GNDA.n6979 185
R8405 GNDA.n6982 GNDA.n6981 185
R8406 GNDA.n6984 GNDA.n6983 185
R8407 GNDA.n6986 GNDA.n6985 185
R8408 GNDA.n6988 GNDA.n6987 185
R8409 GNDA.n6990 GNDA.n6989 185
R8410 GNDA.n6992 GNDA.n6991 185
R8411 GNDA.n6974 GNDA.n6973 185
R8412 GNDA.n6968 GNDA.n6967 185
R8413 GNDA.n6966 GNDA.n6965 185
R8414 GNDA.n6961 GNDA.n6960 185
R8415 GNDA.n6956 GNDA.n6934 185
R8416 GNDA.n7029 GNDA.n7028 185
R8417 GNDA.n6933 GNDA.n6931 185
R8418 GNDA.n7035 GNDA.n7034 185
R8419 GNDA.n7037 GNDA.n7036 185
R8420 GNDA.n7290 GNDA.n80 185
R8421 GNDA.n7304 GNDA.n7303 185
R8422 GNDA.n7302 GNDA.n81 185
R8423 GNDA.n7301 GNDA.n7300 185
R8424 GNDA.n7299 GNDA.n7298 185
R8425 GNDA.n7297 GNDA.n7296 185
R8426 GNDA.n7295 GNDA.n7294 185
R8427 GNDA.n7293 GNDA.n7292 185
R8428 GNDA.n7291 GNDA.n57 185
R8429 GNDA.n7273 GNDA.n7272 185
R8430 GNDA.n7275 GNDA.n7274 185
R8431 GNDA.n7277 GNDA.n7276 185
R8432 GNDA.n7279 GNDA.n7278 185
R8433 GNDA.n7281 GNDA.n7280 185
R8434 GNDA.n7283 GNDA.n7282 185
R8435 GNDA.n7285 GNDA.n7284 185
R8436 GNDA.n7287 GNDA.n7286 185
R8437 GNDA.n7289 GNDA.n7288 185
R8438 GNDA.n7255 GNDA.n7254 185
R8439 GNDA.n7257 GNDA.n7256 185
R8440 GNDA.n7259 GNDA.n7258 185
R8441 GNDA.n7261 GNDA.n7260 185
R8442 GNDA.n7263 GNDA.n7262 185
R8443 GNDA.n7265 GNDA.n7264 185
R8444 GNDA.n7267 GNDA.n7266 185
R8445 GNDA.n7269 GNDA.n7268 185
R8446 GNDA.n7271 GNDA.n7270 185
R8447 GNDA.n7253 GNDA.n7252 185
R8448 GNDA.n7247 GNDA.n7246 185
R8449 GNDA.n7245 GNDA.n7244 185
R8450 GNDA.n7240 GNDA.n7239 185
R8451 GNDA.n7235 GNDA.n65 185
R8452 GNDA.n7308 GNDA.n7307 185
R8453 GNDA.n64 GNDA.n62 185
R8454 GNDA.n7314 GNDA.n7313 185
R8455 GNDA.n7316 GNDA.n7315 185
R8456 GNDA.n6833 GNDA.n6832 185
R8457 GNDA.n6827 GNDA.n6826 185
R8458 GNDA.n6825 GNDA.n6824 185
R8459 GNDA.n6820 GNDA.n6819 185
R8460 GNDA.n6818 GNDA.n6817 185
R8461 GNDA.n6812 GNDA.n6811 185
R8462 GNDA.n6807 GNDA.n6786 185
R8463 GNDA.n6890 GNDA.n6889 185
R8464 GNDA.n6785 GNDA.n6783 185
R8465 GNDA.n1022 GNDA.n1021 185
R8466 GNDA.n1024 GNDA.n935 185
R8467 GNDA.n1027 GNDA.n1026 185
R8468 GNDA.n1028 GNDA.n934 185
R8469 GNDA.n1030 GNDA.n1029 185
R8470 GNDA.n1032 GNDA.n933 185
R8471 GNDA.n1035 GNDA.n1034 185
R8472 GNDA.n1036 GNDA.n932 185
R8473 GNDA.n1038 GNDA.n1037 185
R8474 GNDA.n1004 GNDA.n940 185
R8475 GNDA.n1006 GNDA.n1005 185
R8476 GNDA.n1008 GNDA.n939 185
R8477 GNDA.n1011 GNDA.n1010 185
R8478 GNDA.n1012 GNDA.n938 185
R8479 GNDA.n1014 GNDA.n1013 185
R8480 GNDA.n1016 GNDA.n937 185
R8481 GNDA.n1019 GNDA.n1018 185
R8482 GNDA.n1020 GNDA.n936 185
R8483 GNDA.n986 GNDA.n594 185
R8484 GNDA.n989 GNDA.n988 185
R8485 GNDA.n991 GNDA.n990 185
R8486 GNDA.n993 GNDA.n943 185
R8487 GNDA.n995 GNDA.n994 185
R8488 GNDA.n996 GNDA.n942 185
R8489 GNDA.n998 GNDA.n997 185
R8490 GNDA.n1000 GNDA.n941 185
R8491 GNDA.n1003 GNDA.n1002 185
R8492 GNDA.n985 GNDA.n593 185
R8493 GNDA.n983 GNDA.n982 185
R8494 GNDA.n946 GNDA.n945 185
R8495 GNDA.n972 GNDA.n971 185
R8496 GNDA.n969 GNDA.n967 185
R8497 GNDA.n965 GNDA.n931 185
R8498 GNDA.n1046 GNDA.n1045 185
R8499 GNDA.n1043 GNDA.n929 185
R8500 GNDA.n1042 GNDA.n1041 185
R8501 GNDA.n7209 GNDA.n7208 185
R8502 GNDA.n7211 GNDA.n7210 185
R8503 GNDA.n7213 GNDA.n7212 185
R8504 GNDA.n7215 GNDA.n7214 185
R8505 GNDA.n7217 GNDA.n7216 185
R8506 GNDA.n7219 GNDA.n7218 185
R8507 GNDA.n7221 GNDA.n7220 185
R8508 GNDA.n7223 GNDA.n7222 185
R8509 GNDA.n7224 GNDA.n20 185
R8510 GNDA.n7191 GNDA.n7190 185
R8511 GNDA.n7193 GNDA.n7192 185
R8512 GNDA.n7195 GNDA.n7194 185
R8513 GNDA.n7197 GNDA.n7196 185
R8514 GNDA.n7199 GNDA.n7198 185
R8515 GNDA.n7201 GNDA.n7200 185
R8516 GNDA.n7203 GNDA.n7202 185
R8517 GNDA.n7205 GNDA.n7204 185
R8518 GNDA.n7207 GNDA.n7206 185
R8519 GNDA.n7173 GNDA.n7172 185
R8520 GNDA.n7175 GNDA.n7174 185
R8521 GNDA.n7177 GNDA.n7176 185
R8522 GNDA.n7179 GNDA.n7178 185
R8523 GNDA.n7181 GNDA.n7180 185
R8524 GNDA.n7183 GNDA.n7182 185
R8525 GNDA.n7185 GNDA.n7184 185
R8526 GNDA.n7187 GNDA.n7186 185
R8527 GNDA.n7189 GNDA.n7188 185
R8528 GNDA.n7171 GNDA.n7170 185
R8529 GNDA.n7165 GNDA.n7164 185
R8530 GNDA.n7160 GNDA.n3 185
R8531 GNDA.n7331 GNDA.n7330 185
R8532 GNDA.n34 GNDA.n2 185
R8533 GNDA.n38 GNDA.n37 185
R8534 GNDA.n36 GNDA.n33 185
R8535 GNDA.n23 GNDA.n21 185
R8536 GNDA.n7327 GNDA.n7326 185
R8537 GNDA.n1219 GNDA.n647 175.546
R8538 GNDA.n1224 GNDA.n647 175.546
R8539 GNDA.n1224 GNDA.n644 175.546
R8540 GNDA.n1228 GNDA.n644 175.546
R8541 GNDA.n1229 GNDA.n1228 175.546
R8542 GNDA.n1230 GNDA.n1229 175.546
R8543 GNDA.n1230 GNDA.n642 175.546
R8544 GNDA.n1234 GNDA.n642 175.546
R8545 GNDA.n1234 GNDA.n639 175.546
R8546 GNDA.n1337 GNDA.n639 175.546
R8547 GNDA.n1337 GNDA.n640 175.546
R8548 GNDA.n1239 GNDA.n571 175.546
R8549 GNDA.n1330 GNDA.n1239 175.546
R8550 GNDA.n1330 GNDA.n1240 175.546
R8551 GNDA.n1322 GNDA.n1240 175.546
R8552 GNDA.n1322 GNDA.n1319 175.546
R8553 GNDA.n1319 GNDA.n551 175.546
R8554 GNDA.n6248 GNDA.n551 175.546
R8555 GNDA.n6248 GNDA.n543 175.546
R8556 GNDA.n6259 GNDA.n543 175.546
R8557 GNDA.n6259 GNDA.n544 175.546
R8558 GNDA.n1341 GNDA.n544 175.546
R8559 GNDA.n1191 GNDA.n1190 175.546
R8560 GNDA.n1188 GNDA.n1168 175.546
R8561 GNDA.n1184 GNDA.n1182 175.546
R8562 GNDA.n1180 GNDA.n1175 175.546
R8563 GNDA.n6220 GNDA.n572 175.546
R8564 GNDA.n1200 GNDA.n653 175.546
R8565 GNDA.n1204 GNDA.n1202 175.546
R8566 GNDA.n1208 GNDA.n651 175.546
R8567 GNDA.n1212 GNDA.n1210 175.546
R8568 GNDA.n1216 GNDA.n649 175.546
R8569 GNDA.n1166 GNDA.n1165 175.546
R8570 GNDA.n1170 GNDA.n1169 175.546
R8571 GNDA.n1172 GNDA.n1171 175.546
R8572 GNDA.n1177 GNDA.n1176 175.546
R8573 GNDA.n6218 GNDA.n574 175.546
R8574 GNDA.n1145 GNDA.n1143 175.546
R8575 GNDA.n1149 GNDA.n911 175.546
R8576 GNDA.n1153 GNDA.n1151 175.546
R8577 GNDA.n1157 GNDA.n909 175.546
R8578 GNDA.n1160 GNDA.n1159 175.546
R8579 GNDA.n6193 GNDA.n586 175.546
R8580 GNDA.n6193 GNDA.n597 175.546
R8581 GNDA.n6189 GNDA.n597 175.546
R8582 GNDA.n6189 GNDA.n600 175.546
R8583 GNDA.n6109 GNDA.n600 175.546
R8584 GNDA.n6109 GNDA.n6105 175.546
R8585 GNDA.n6120 GNDA.n6105 175.546
R8586 GNDA.n6120 GNDA.n624 175.546
R8587 GNDA.n6125 GNDA.n624 175.546
R8588 GNDA.n6125 GNDA.n565 175.546
R8589 GNDA.n6227 GNDA.n565 175.546
R8590 GNDA.n1132 GNDA.n1130 175.546
R8591 GNDA.n1128 GNDA.n1104 175.546
R8592 GNDA.n1124 GNDA.n1122 175.546
R8593 GNDA.n1120 GNDA.n1112 175.546
R8594 GNDA.n6210 GNDA.n588 175.546
R8595 GNDA.n1076 GNDA.n1075 175.546
R8596 GNDA.n1072 GNDA.n1071 175.546
R8597 GNDA.n1068 GNDA.n1067 175.546
R8598 GNDA.n1064 GNDA.n1063 175.546
R8599 GNDA.n1060 GNDA.n1059 175.546
R8600 GNDA.n1085 GNDA.n920 175.546
R8601 GNDA.n1089 GNDA.n1087 175.546
R8602 GNDA.n1093 GNDA.n918 175.546
R8603 GNDA.n1096 GNDA.n1095 175.546
R8604 GNDA.n1100 GNDA.n1099 175.546
R8605 GNDA.n1055 GNDA.n1054 175.546
R8606 GNDA.n1054 GNDA.n923 175.546
R8607 GNDA.n1048 GNDA.n923 175.546
R8608 GNDA.n1048 GNDA.n928 175.546
R8609 GNDA.n963 GNDA.n928 175.546
R8610 GNDA.n974 GNDA.n963 175.546
R8611 GNDA.n974 GNDA.n947 175.546
R8612 GNDA.n979 GNDA.n947 175.546
R8613 GNDA.n979 GNDA.n592 175.546
R8614 GNDA.n6201 GNDA.n592 175.546
R8615 GNDA.n6201 GNDA.n591 175.546
R8616 GNDA.n1134 GNDA.n1102 175.546
R8617 GNDA.n1107 GNDA.n1106 175.546
R8618 GNDA.n1113 GNDA.n1109 175.546
R8619 GNDA.n1117 GNDA.n1115 175.546
R8620 GNDA.n6208 GNDA.n590 175.546
R8621 GNDA.n6635 GNDA.n6632 175.546
R8622 GNDA.n6638 GNDA.n6637 175.546
R8623 GNDA.n6643 GNDA.n6640 175.546
R8624 GNDA.n6646 GNDA.n6645 175.546
R8625 GNDA.n6650 GNDA.n6648 175.546
R8626 GNDA.n6755 GNDA.n351 175.546
R8627 GNDA.n6751 GNDA.n351 175.546
R8628 GNDA.n6751 GNDA.n353 175.546
R8629 GNDA.n6747 GNDA.n353 175.546
R8630 GNDA.n6747 GNDA.n355 175.546
R8631 GNDA.n6738 GNDA.n355 175.546
R8632 GNDA.n6738 GNDA.n6737 175.546
R8633 GNDA.n6737 GNDA.n6623 175.546
R8634 GNDA.n6733 GNDA.n6623 175.546
R8635 GNDA.n6733 GNDA.n6625 175.546
R8636 GNDA.n6729 GNDA.n6625 175.546
R8637 GNDA.n348 GNDA.n305 175.546
R8638 GNDA.n344 GNDA.n342 175.546
R8639 GNDA.n340 GNDA.n312 175.546
R8640 GNDA.n336 GNDA.n334 175.546
R8641 GNDA.n332 GNDA.n320 175.546
R8642 GNDA.n844 GNDA.n695 175.546
R8643 GNDA.n840 GNDA.n695 175.546
R8644 GNDA.n840 GNDA.n697 175.546
R8645 GNDA.n836 GNDA.n697 175.546
R8646 GNDA.n836 GNDA.n834 175.546
R8647 GNDA.n834 GNDA.n833 175.546
R8648 GNDA.n833 GNDA.n700 175.546
R8649 GNDA.n829 GNDA.n700 175.546
R8650 GNDA.n829 GNDA.n702 175.546
R8651 GNDA.n825 GNDA.n702 175.546
R8652 GNDA.n825 GNDA.n705 175.546
R8653 GNDA.n806 GNDA.n805 175.546
R8654 GNDA.n802 GNDA.n801 175.546
R8655 GNDA.n795 GNDA.n794 175.546
R8656 GNDA.n788 GNDA.n787 175.546
R8657 GNDA.n816 GNDA.n815 175.546
R8658 GNDA.n871 GNDA.n666 175.546
R8659 GNDA.n879 GNDA.n666 175.546
R8660 GNDA.n883 GNDA.n881 175.546
R8661 GNDA.n891 GNDA.n662 175.546
R8662 GNDA.n895 GNDA.n893 175.546
R8663 GNDA.n902 GNDA.n658 175.546
R8664 GNDA.n865 GNDA.n864 175.546
R8665 GNDA.n861 GNDA.n860 175.546
R8666 GNDA.n857 GNDA.n856 175.546
R8667 GNDA.n853 GNDA.n852 175.546
R8668 GNDA.n849 GNDA.n848 175.546
R8669 GNDA.n874 GNDA.n873 175.546
R8670 GNDA.n877 GNDA.n876 175.546
R8671 GNDA.n886 GNDA.n885 175.546
R8672 GNDA.n889 GNDA.n888 175.546
R8673 GNDA.n898 GNDA.n897 175.546
R8674 GNDA.n7108 GNDA.n7107 175.546
R8675 GNDA.n220 GNDA.n200 175.546
R8676 GNDA.n202 GNDA.n199 175.546
R8677 GNDA.n210 GNDA.n209 175.546
R8678 GNDA.n7045 GNDA.n189 175.546
R8679 GNDA.n7132 GNDA.n137 175.546
R8680 GNDA.n7128 GNDA.n142 175.546
R8681 GNDA.n7126 GNDA.n7125 175.546
R8682 GNDA.n7122 GNDA.n7121 175.546
R8683 GNDA.n7118 GNDA.n7117 175.546
R8684 GNDA.n672 GNDA.n671 175.546
R8685 GNDA.n676 GNDA.n675 175.546
R8686 GNDA.n680 GNDA.n679 175.546
R8687 GNDA.n684 GNDA.n683 175.546
R8688 GNDA.n688 GNDA.n687 175.546
R8689 GNDA.n152 GNDA.n143 175.546
R8690 GNDA.n145 GNDA.n144 175.546
R8691 GNDA.n147 GNDA.n146 175.546
R8692 GNDA.n149 GNDA.n148 175.546
R8693 GNDA.n151 GNDA.n150 175.546
R8694 GNDA.n6927 GNDA.n227 175.546
R8695 GNDA.n7032 GNDA.n7031 175.546
R8696 GNDA.n6958 GNDA.n6957 175.546
R8697 GNDA.n6963 GNDA.n6962 175.546
R8698 GNDA.n6971 GNDA.n6970 175.546
R8699 GNDA.n266 GNDA.n265 175.546
R8700 GNDA.n270 GNDA.n269 175.546
R8701 GNDA.n274 GNDA.n273 175.546
R8702 GNDA.n279 GNDA.n241 175.546
R8703 GNDA.n240 GNDA.n230 175.546
R8704 GNDA.n6924 GNDA.n230 175.546
R8705 GNDA.n258 GNDA.n257 175.546
R8706 GNDA.n254 GNDA.n253 175.546
R8707 GNDA.n250 GNDA.n249 175.546
R8708 GNDA.n246 GNDA.n245 175.546
R8709 GNDA.n242 GNDA.n130 175.546
R8710 GNDA.n308 GNDA.n307 175.546
R8711 GNDA.n313 GNDA.n310 175.546
R8712 GNDA.n316 GNDA.n315 175.546
R8713 GNDA.n321 GNDA.n318 175.546
R8714 GNDA.n324 GNDA.n323 175.546
R8715 GNDA.n6893 GNDA.n6892 175.546
R8716 GNDA.n6809 GNDA.n6808 175.546
R8717 GNDA.n6815 GNDA.n6814 175.546
R8718 GNDA.n6822 GNDA.n6821 175.546
R8719 GNDA.n6830 GNDA.n6829 175.546
R8720 GNDA.n289 GNDA.n288 175.546
R8721 GNDA.n6915 GNDA.n288 175.546
R8722 GNDA.n6913 GNDA.n6912 175.546
R8723 GNDA.n6909 GNDA.n6908 175.546
R8724 GNDA.n6905 GNDA.n6904 175.546
R8725 GNDA.n6901 GNDA.n6900 175.546
R8726 GNDA.n6779 GNDA.n290 175.546
R8727 GNDA.n6779 GNDA.n292 175.546
R8728 GNDA.n6775 GNDA.n292 175.546
R8729 GNDA.n6775 GNDA.n294 175.546
R8730 GNDA.n6771 GNDA.n294 175.546
R8731 GNDA.n6771 GNDA.n296 175.546
R8732 GNDA.n6767 GNDA.n296 175.546
R8733 GNDA.n6767 GNDA.n298 175.546
R8734 GNDA.n6763 GNDA.n298 175.546
R8735 GNDA.n6763 GNDA.n300 175.546
R8736 GNDA.n6759 GNDA.n300 175.546
R8737 GNDA.n58 GNDA.n54 175.546
R8738 GNDA.n7311 GNDA.n7310 175.546
R8739 GNDA.n7237 GNDA.n7236 175.546
R8740 GNDA.n7242 GNDA.n7241 175.546
R8741 GNDA.n7250 GNDA.n7249 175.546
R8742 GNDA.n6671 GNDA.n6670 175.546
R8743 GNDA.n6668 GNDA.n6634 175.546
R8744 GNDA.n6664 GNDA.n6662 175.546
R8745 GNDA.n6660 GNDA.n6642 175.546
R8746 GNDA.n6656 GNDA.n6654 175.546
R8747 GNDA.n6725 GNDA.n6675 175.546
R8748 GNDA.n6721 GNDA.n6675 175.546
R8749 GNDA.n6721 GNDA.n6677 175.546
R8750 GNDA.n6717 GNDA.n6677 175.546
R8751 GNDA.n6717 GNDA.n6679 175.546
R8752 GNDA.n6713 GNDA.n6679 175.546
R8753 GNDA.n6713 GNDA.n6681 175.546
R8754 GNDA.n6709 GNDA.n6681 175.546
R8755 GNDA.n6709 GNDA.n6683 175.546
R8756 GNDA.n6705 GNDA.n6683 175.546
R8757 GNDA.n6705 GNDA.n6685 175.546
R8758 GNDA.n7324 GNDA.n24 175.546
R8759 GNDA.n40 GNDA.n25 175.546
R8760 GNDA.n31 GNDA.n30 175.546
R8761 GNDA.n7162 GNDA.n7161 175.546
R8762 GNDA.n7168 GNDA.n7167 175.546
R8763 GNDA.n6701 GNDA.n6687 175.546
R8764 GNDA.n6697 GNDA.n6687 175.546
R8765 GNDA.n6697 GNDA.n6689 175.546
R8766 GNDA.n6693 GNDA.n6689 175.546
R8767 GNDA.n6693 GNDA.n6690 175.546
R8768 GNDA.n6690 GNDA.n93 175.546
R8769 GNDA.n7145 GNDA.n93 175.546
R8770 GNDA.n7145 GNDA.n91 175.546
R8771 GNDA.n7150 GNDA.n91 175.546
R8772 GNDA.n7150 GNDA.n89 175.546
R8773 GNDA.n7154 GNDA.n89 175.546
R8774 GNDA.n158 GNDA.n100 173.881
R8775 GNDA.t743 GNDA.n101 172.876
R8776 GNDA.t743 GNDA.n112 172.615
R8777 GNDA.n7134 GNDA.n100 171.624
R8778 GNDA.n6256 GNDA.n547 163.333
R8779 GNDA.n6132 GNDA.n6130 163.333
R8780 GNDA.n7049 GNDA.n7048 163.333
R8781 GNDA.n6834 GNDA.n6833 163.333
R8782 GNDA.n720 GNDA.n710 163.333
R8783 GNDA.n6975 GNDA.n6974 163.333
R8784 GNDA.n7254 GNDA.n7253 163.333
R8785 GNDA.n986 GNDA.n985 163.333
R8786 GNDA.n7172 GNDA.n7171 163.333
R8787 GNDA.n4790 GNDA.n4789 161.3
R8788 GNDA.n4133 GNDA.n4132 161.3
R8789 GNDA.n1288 GNDA.n1286 150
R8790 GNDA.n1284 GNDA.n1249 150
R8791 GNDA.n1280 GNDA.n1278 150
R8792 GNDA.n1276 GNDA.n1251 150
R8793 GNDA.n1272 GNDA.n1270 150
R8794 GNDA.n1268 GNDA.n1253 150
R8795 GNDA.n1264 GNDA.n1263 150
R8796 GNDA.n1261 GNDA.n1257 150
R8797 GNDA.n1327 GNDA.n1312 150
R8798 GNDA.n1325 GNDA.n1314 150
R8799 GNDA.n6251 GNDA.n550 150
R8800 GNDA.n6254 GNDA.n6253 150
R8801 GNDA.n1296 GNDA.n1294 150
R8802 GNDA.n1300 GNDA.n1245 150
R8803 GNDA.n1304 GNDA.n1302 150
R8804 GNDA.n1310 GNDA.n1243 150
R8805 GNDA.n6162 GNDA.n610 150
R8806 GNDA.n6158 GNDA.n6156 150
R8807 GNDA.n6154 GNDA.n612 150
R8808 GNDA.n6150 GNDA.n6148 150
R8809 GNDA.n6146 GNDA.n614 150
R8810 GNDA.n6142 GNDA.n6141 150
R8811 GNDA.n6139 GNDA.n617 150
R8812 GNDA.n6135 GNDA.n6134 150
R8813 GNDA.n6184 GNDA.n6183 150
R8814 GNDA.n6186 GNDA.n604 150
R8815 GNDA.n6116 GNDA.n6114 150
R8816 GNDA.n6128 GNDA.n622 150
R8817 GNDA.n6170 GNDA.n608 150
R8818 GNDA.n6174 GNDA.n6172 150
R8819 GNDA.n6178 GNDA.n606 150
R8820 GNDA.n6181 GNDA.n6180 150
R8821 GNDA.n7081 GNDA.n7080 150
R8822 GNDA.n7077 GNDA.n7076 150
R8823 GNDA.n7073 GNDA.n7072 150
R8824 GNDA.n7069 GNDA.n7068 150
R8825 GNDA.n7065 GNDA.n7064 150
R8826 GNDA.n7061 GNDA.n7060 150
R8827 GNDA.n7057 GNDA.n7056 150
R8828 GNDA.n7053 GNDA.n7052 150
R8829 GNDA.n7104 GNDA.n169 150
R8830 GNDA.n217 GNDA.n170 150
R8831 GNDA.n214 GNDA.n213 150
R8832 GNDA.n206 GNDA.n205 150
R8833 GNDA.n7089 GNDA.n7088 150
R8834 GNDA.n7093 GNDA.n7092 150
R8835 GNDA.n7097 GNDA.n7096 150
R8836 GNDA.n7101 GNDA.n7100 150
R8837 GNDA.n6866 GNDA.n6865 150
R8838 GNDA.n6862 GNDA.n6861 150
R8839 GNDA.n6858 GNDA.n6857 150
R8840 GNDA.n6854 GNDA.n6853 150
R8841 GNDA.n6850 GNDA.n6849 150
R8842 GNDA.n6846 GNDA.n6845 150
R8843 GNDA.n6842 GNDA.n6841 150
R8844 GNDA.n6838 GNDA.n6837 150
R8845 GNDA.n6889 GNDA.n6785 150
R8846 GNDA.n6811 GNDA.n6786 150
R8847 GNDA.n6819 GNDA.n6818 150
R8848 GNDA.n6826 GNDA.n6825 150
R8849 GNDA.n6874 GNDA.n6873 150
R8850 GNDA.n6878 GNDA.n6877 150
R8851 GNDA.n6882 GNDA.n6881 150
R8852 GNDA.n6886 GNDA.n6885 150
R8853 GNDA.n760 GNDA.n759 150
R8854 GNDA.n756 GNDA.n755 150
R8855 GNDA.n752 GNDA.n751 150
R8856 GNDA.n748 GNDA.n747 150
R8857 GNDA.n744 GNDA.n743 150
R8858 GNDA.n740 GNDA.n739 150
R8859 GNDA.n736 GNDA.n735 150
R8860 GNDA.n732 GNDA.n731 150
R8861 GNDA.n809 GNDA.n729 150
R8862 GNDA.n798 GNDA.n797 150
R8863 GNDA.n791 GNDA.n790 150
R8864 GNDA.n812 GNDA.n709 150
R8865 GNDA.n768 GNDA.n767 150
R8866 GNDA.n772 GNDA.n771 150
R8867 GNDA.n776 GNDA.n775 150
R8868 GNDA.n778 GNDA.n728 150
R8869 GNDA.n7007 GNDA.n7006 150
R8870 GNDA.n7003 GNDA.n7002 150
R8871 GNDA.n6999 GNDA.n6998 150
R8872 GNDA.n6995 GNDA.n6994 150
R8873 GNDA.n6991 GNDA.n6990 150
R8874 GNDA.n6987 GNDA.n6986 150
R8875 GNDA.n6983 GNDA.n6982 150
R8876 GNDA.n6979 GNDA.n6978 150
R8877 GNDA.n7036 GNDA.n7035 150
R8878 GNDA.n7028 GNDA.n6933 150
R8879 GNDA.n6960 GNDA.n6934 150
R8880 GNDA.n6967 GNDA.n6966 150
R8881 GNDA.n7025 GNDA.n6950 150
R8882 GNDA.n7021 GNDA.n7020 150
R8883 GNDA.n7017 GNDA.n7016 150
R8884 GNDA.n7013 GNDA.n7012 150
R8885 GNDA.n7286 GNDA.n7285 150
R8886 GNDA.n7282 GNDA.n7281 150
R8887 GNDA.n7278 GNDA.n7277 150
R8888 GNDA.n7274 GNDA.n7273 150
R8889 GNDA.n7270 GNDA.n7269 150
R8890 GNDA.n7266 GNDA.n7265 150
R8891 GNDA.n7262 GNDA.n7261 150
R8892 GNDA.n7258 GNDA.n7257 150
R8893 GNDA.n7315 GNDA.n7314 150
R8894 GNDA.n7307 GNDA.n64 150
R8895 GNDA.n7239 GNDA.n65 150
R8896 GNDA.n7246 GNDA.n7245 150
R8897 GNDA.n7304 GNDA.n81 150
R8898 GNDA.n7300 GNDA.n7299 150
R8899 GNDA.n7296 GNDA.n7295 150
R8900 GNDA.n7292 GNDA.n7291 150
R8901 GNDA.n1018 GNDA.n1016 150
R8902 GNDA.n1014 GNDA.n938 150
R8903 GNDA.n1010 GNDA.n1008 150
R8904 GNDA.n1006 GNDA.n940 150
R8905 GNDA.n1002 GNDA.n1000 150
R8906 GNDA.n998 GNDA.n942 150
R8907 GNDA.n994 GNDA.n993 150
R8908 GNDA.n991 GNDA.n988 150
R8909 GNDA.n1043 GNDA.n1042 150
R8910 GNDA.n1045 GNDA.n931 150
R8911 GNDA.n971 GNDA.n969 150
R8912 GNDA.n983 GNDA.n945 150
R8913 GNDA.n1026 GNDA.n1024 150
R8914 GNDA.n1030 GNDA.n934 150
R8915 GNDA.n1034 GNDA.n1032 150
R8916 GNDA.n1038 GNDA.n932 150
R8917 GNDA.n7204 GNDA.n7203 150
R8918 GNDA.n7200 GNDA.n7199 150
R8919 GNDA.n7196 GNDA.n7195 150
R8920 GNDA.n7192 GNDA.n7191 150
R8921 GNDA.n7188 GNDA.n7187 150
R8922 GNDA.n7184 GNDA.n7183 150
R8923 GNDA.n7180 GNDA.n7179 150
R8924 GNDA.n7176 GNDA.n7175 150
R8925 GNDA.n7327 GNDA.n21 150
R8926 GNDA.n37 GNDA.n36 150
R8927 GNDA.n7330 GNDA.n2 150
R8928 GNDA.n7164 GNDA.n3 150
R8929 GNDA.n7212 GNDA.n7211 150
R8930 GNDA.n7216 GNDA.n7215 150
R8931 GNDA.n7220 GNDA.n7219 150
R8932 GNDA.n7222 GNDA.n20 150
R8933 GNDA.n6093 GNDA.n6092 148.017
R8934 GNDA.n4798 GNDA.n4797 148.017
R8935 GNDA.n4092 GNDA.n4091 148.017
R8936 GNDA.n4098 GNDA.n4097 148.017
R8937 GNDA.n6264 GNDA.n540 136.145
R8938 GNDA.n6265 GNDA.n539 136.145
R8939 GNDA.n6266 GNDA.n538 136.145
R8940 GNDA.n6269 GNDA.n535 136.145
R8941 GNDA.n6270 GNDA.n534 136.145
R8942 GNDA.n6273 GNDA.n531 136.145
R8943 GNDA.n6274 GNDA.n530 136.145
R8944 GNDA.n6275 GNDA.n529 136.145
R8945 GNDA.n6278 GNDA.n526 136.145
R8946 GNDA.n6279 GNDA.n525 136.145
R8947 GNDA.n958 GNDA.n957 134.268
R8948 GNDA.n958 GNDA.n951 134.268
R8949 GNDA.n921 GNDA.n282 132.721
R8950 GNDA.n6262 GNDA.t776 130.001
R8951 GNDA.n563 GNDA.t827 130.001
R8952 GNDA.n561 GNDA.t782 130.001
R8953 GNDA.n598 GNDA.t830 130.001
R8954 GNDA.n582 GNDA.t789 130.001
R8955 GNDA.n1050 GNDA.t779 130.001
R8956 GNDA.n925 GNDA.t811 130.001
R8957 GNDA.n629 GNDA.t844 130
R8958 GNDA.n6223 GNDA.n6222 124.832
R8959 GNDA.n6216 GNDA.n566 124.832
R8960 GNDA.n6213 GNDA.n6212 124.832
R8961 GNDA.n6206 GNDA.n6205 124.832
R8962 GNDA.n7230 GNDA.n83 124.832
R8963 GNDA.n328 GNDA.n55 124.832
R8964 GNDA.n903 GNDA.n902 124.832
R8965 GNDA.n900 GNDA.n656 124.832
R8966 GNDA.n7114 GNDA.n7113 124.832
R8967 GNDA.n6951 GNDA.n160 124.832
R8968 GNDA.n326 GNDA.n85 124.832
R8969 GNDA.n7228 GNDA.n86 124.832
R8970 GNDA.n1352 GNDA.n1350 124.59
R8971 GNDA.n1819 GNDA.n1818 124.028
R8972 GNDA.n1821 GNDA.n1820 124.028
R8973 GNDA.n1823 GNDA.n1822 124.028
R8974 GNDA.n1825 GNDA.n1824 124.028
R8975 GNDA.n1827 GNDA.n1826 124.028
R8976 GNDA.n1829 GNDA.n1828 124.028
R8977 GNDA.n1360 GNDA.n1359 124.028
R8978 GNDA.n1358 GNDA.n1357 124.028
R8979 GNDA.n1356 GNDA.n1355 124.028
R8980 GNDA.n1354 GNDA.n1353 124.028
R8981 GNDA.n1352 GNDA.n1351 124.028
R8982 GNDA.t131 GNDA.t119 121.772
R8983 GNDA.t29 GNDA.t102 121.772
R8984 GNDA.n6281 GNDA.t873 116.073
R8985 GNDA.n6619 GNDA.t35 115.105
R8986 GNDA.n6620 GNDA.t59 114.635
R8987 GNDA.n6281 GNDA.t61 114.635
R8988 GNDA.n4130 GNDA.t868 113.085
R8989 GNDA.n4130 GNDA.t94 113.085
R8990 GNDA.n6235 GNDA.n556 101.718
R8991 GNDA.n953 GNDA.n948 101.718
R8992 GNDA.n961 GNDA.n960 101.718
R8993 GNDA.n6244 GNDA.n558 101.718
R8994 GNDA.n1053 GNDA.n1052 99.6733
R8995 GNDA.n978 GNDA.n976 99.6733
R8996 GNDA.n6192 GNDA.n6191 99.6733
R8997 GNDA.n6124 GNDA.n6123 99.6733
R8998 GNDA.n1321 GNDA.n1320 99.6733
R8999 GNDA.n6260 GNDA.n542 99.6733
R9000 GNDA.n1342 GNDA.n542 99.6733
R9001 GNDA.t743 GNDA.n104 47.6748
R9002 GNDA.n1052 GNDA.n1051 96.3509
R9003 GNDA.t743 GNDA.n6214 96.3509
R9004 GNDA.n6247 GNDA.t88 96.3509
R9005 GNDA.t743 GNDA.n580 95.2434
R9006 GNDA.n1053 GNDA.n926 91.921
R9007 GNDA.n927 GNDA.t17 91.921
R9008 GNDA.n6261 GNDA.n6260 91.921
R9009 GNDA.n6242 GNDA.n6234 91.069
R9010 GNDA.n6242 GNDA.n6241 91.069
R9011 GNDA.n6239 GNDA.n6232 91.069
R9012 GNDA.n6239 GNDA.n6238 91.069
R9013 GNDA.n957 GNDA.n956 91.069
R9014 GNDA.n952 GNDA.n951 91.069
R9015 GNDA.t179 GNDA.n975 90.8135
R9016 GNDA.t113 GNDA.n6107 90.8135
R9017 GNDA.n1331 GNDA.t67 90.8135
R9018 GNDA.t177 GNDA.n977 86.3836
R9019 GNDA.n6121 GNDA.t881 86.3836
R9020 GNDA.t160 GNDA.n555 86.3836
R9021 GNDA.n6744 GNDA.n6743 84.306
R9022 GNDA.t879 GNDA.n6203 79.7387
R9023 GNDA.n6760 GNDA.n301 76.4476
R9024 GNDA.n6728 GNDA.n6727 76.4476
R9025 GNDA.t743 GNDA.n100 76.3879
R9026 GNDA.n1194 GNDA.n906 76.3222
R9027 GNDA.n1190 GNDA.n1189 76.3222
R9028 GNDA.n1183 GNDA.n1168 76.3222
R9029 GNDA.n1182 GNDA.n1181 76.3222
R9030 GNDA.n1175 GNDA.n1174 76.3222
R9031 GNDA.n6221 GNDA.n6220 76.3222
R9032 GNDA.n1195 GNDA.n653 76.3222
R9033 GNDA.n1202 GNDA.n1201 76.3222
R9034 GNDA.n1203 GNDA.n651 76.3222
R9035 GNDA.n1210 GNDA.n1209 76.3222
R9036 GNDA.n1211 GNDA.n649 76.3222
R9037 GNDA.n1218 GNDA.n1217 76.3222
R9038 GNDA.n1165 GNDA.n575 76.3222
R9039 GNDA.n1169 GNDA.n576 76.3222
R9040 GNDA.n1171 GNDA.n577 76.3222
R9041 GNDA.n1176 GNDA.n578 76.3222
R9042 GNDA.n579 GNDA.n574 76.3222
R9043 GNDA.n6217 GNDA.n6216 76.3222
R9044 GNDA.n1143 GNDA.n1142 76.3222
R9045 GNDA.n1144 GNDA.n911 76.3222
R9046 GNDA.n1151 GNDA.n1150 76.3222
R9047 GNDA.n1152 GNDA.n909 76.3222
R9048 GNDA.n1159 GNDA.n1158 76.3222
R9049 GNDA.n1163 GNDA.n907 76.3222
R9050 GNDA.n1131 GNDA.n913 76.3222
R9051 GNDA.n1130 GNDA.n1129 76.3222
R9052 GNDA.n1123 GNDA.n1104 76.3222
R9053 GNDA.n1122 GNDA.n1121 76.3222
R9054 GNDA.n1112 GNDA.n1111 76.3222
R9055 GNDA.n6211 GNDA.n6210 76.3222
R9056 GNDA.n1079 GNDA.n287 76.3222
R9057 GNDA.n1075 GNDA.n286 76.3222
R9058 GNDA.n1071 GNDA.n285 76.3222
R9059 GNDA.n1067 GNDA.n284 76.3222
R9060 GNDA.n1063 GNDA.n283 76.3222
R9061 GNDA.n1059 GNDA.n282 76.3222
R9062 GNDA.n1080 GNDA.n920 76.3222
R9063 GNDA.n1087 GNDA.n1086 76.3222
R9064 GNDA.n1088 GNDA.n918 76.3222
R9065 GNDA.n1095 GNDA.n1094 76.3222
R9066 GNDA.n1099 GNDA.n916 76.3222
R9067 GNDA.n1137 GNDA.n1101 76.3222
R9068 GNDA.n1136 GNDA.n1135 76.3222
R9069 GNDA.n1105 GNDA.n1102 76.3222
R9070 GNDA.n1108 GNDA.n1107 76.3222
R9071 GNDA.n1114 GNDA.n1113 76.3222
R9072 GNDA.n1117 GNDA.n1116 76.3222
R9073 GNDA.n6208 GNDA.n6207 76.3222
R9074 GNDA.n6632 GNDA.n6631 76.3222
R9075 GNDA.n6637 GNDA.n6636 76.3222
R9076 GNDA.n6640 GNDA.n6639 76.3222
R9077 GNDA.n6645 GNDA.n6644 76.3222
R9078 GNDA.n6648 GNDA.n6647 76.3222
R9079 GNDA.n6649 GNDA.n83 76.3222
R9080 GNDA.n350 GNDA.n349 76.3222
R9081 GNDA.n343 GNDA.n305 76.3222
R9082 GNDA.n342 GNDA.n341 76.3222
R9083 GNDA.n335 GNDA.n312 76.3222
R9084 GNDA.n334 GNDA.n333 76.3222
R9085 GNDA.n327 GNDA.n320 76.3222
R9086 GNDA.n657 GNDA.n196 76.3222
R9087 GNDA.n806 GNDA.n195 76.3222
R9088 GNDA.n801 GNDA.n194 76.3222
R9089 GNDA.n794 GNDA.n193 76.3222
R9090 GNDA.n787 GNDA.n192 76.3222
R9091 GNDA.n816 GNDA.n191 76.3222
R9092 GNDA.n870 GNDA.n869 76.3222
R9093 GNDA.n880 GNDA.n879 76.3222
R9094 GNDA.n883 GNDA.n882 76.3222
R9095 GNDA.n892 GNDA.n891 76.3222
R9096 GNDA.n895 GNDA.n894 76.3222
R9097 GNDA.n865 GNDA.n113 76.3222
R9098 GNDA.n861 GNDA.n114 76.3222
R9099 GNDA.n857 GNDA.n115 76.3222
R9100 GNDA.n853 GNDA.n116 76.3222
R9101 GNDA.n849 GNDA.n117 76.3222
R9102 GNDA.n845 GNDA.n118 76.3222
R9103 GNDA.n873 GNDA.n668 76.3222
R9104 GNDA.n877 GNDA.n875 76.3222
R9105 GNDA.n885 GNDA.n664 76.3222
R9106 GNDA.n889 GNDA.n887 76.3222
R9107 GNDA.n897 GNDA.n660 76.3222
R9108 GNDA.n900 GNDA.n899 76.3222
R9109 GNDA.n7112 GNDA.n164 76.3222
R9110 GNDA.n7107 GNDA.n167 76.3222
R9111 GNDA.n221 GNDA.n220 76.3222
R9112 GNDA.n202 GNDA.n198 76.3222
R9113 GNDA.n209 GNDA.n197 76.3222
R9114 GNDA.n7045 GNDA.n7044 76.3222
R9115 GNDA.n7136 GNDA.n7135 76.3222
R9116 GNDA.n7133 GNDA.n7132 76.3222
R9117 GNDA.n7128 GNDA.n141 76.3222
R9118 GNDA.n7125 GNDA.n140 76.3222
R9119 GNDA.n7121 GNDA.n139 76.3222
R9120 GNDA.n7117 GNDA.n138 76.3222
R9121 GNDA.n671 GNDA.n119 76.3222
R9122 GNDA.n675 GNDA.n120 76.3222
R9123 GNDA.n679 GNDA.n121 76.3222
R9124 GNDA.n683 GNDA.n122 76.3222
R9125 GNDA.n687 GNDA.n123 76.3222
R9126 GNDA.n691 GNDA.n124 76.3222
R9127 GNDA.n153 GNDA.n152 76.3222
R9128 GNDA.n154 GNDA.n144 76.3222
R9129 GNDA.n155 GNDA.n146 76.3222
R9130 GNDA.n156 GNDA.n148 76.3222
R9131 GNDA.n157 GNDA.n150 76.3222
R9132 GNDA.n160 GNDA.n159 76.3222
R9133 GNDA.n7042 GNDA.n7041 76.3222
R9134 GNDA.n6927 GNDA.n226 76.3222
R9135 GNDA.n7031 GNDA.n225 76.3222
R9136 GNDA.n6958 GNDA.n224 76.3222
R9137 GNDA.n6962 GNDA.n223 76.3222
R9138 GNDA.n6971 GNDA.n222 76.3222
R9139 GNDA.n262 GNDA.n236 76.3222
R9140 GNDA.n266 GNDA.n237 76.3222
R9141 GNDA.n270 GNDA.n238 76.3222
R9142 GNDA.n274 GNDA.n239 76.3222
R9143 GNDA.n280 GNDA.n279 76.3222
R9144 GNDA.n258 GNDA.n125 76.3222
R9145 GNDA.n254 GNDA.n126 76.3222
R9146 GNDA.n250 GNDA.n127 76.3222
R9147 GNDA.n246 GNDA.n128 76.3222
R9148 GNDA.n242 GNDA.n129 76.3222
R9149 GNDA.n7141 GNDA.n7140 76.3222
R9150 GNDA.n307 GNDA.n306 76.3222
R9151 GNDA.n310 GNDA.n309 76.3222
R9152 GNDA.n315 GNDA.n314 76.3222
R9153 GNDA.n318 GNDA.n317 76.3222
R9154 GNDA.n323 GNDA.n322 76.3222
R9155 GNDA.n326 GNDA.n325 76.3222
R9156 GNDA.n6893 GNDA.n48 76.3222
R9157 GNDA.n6808 GNDA.n47 76.3222
R9158 GNDA.n6814 GNDA.n46 76.3222
R9159 GNDA.n6822 GNDA.n45 76.3222
R9160 GNDA.n6829 GNDA.n44 76.3222
R9161 GNDA.n6803 GNDA.n43 76.3222
R9162 GNDA.n6921 GNDA.n6920 76.3222
R9163 GNDA.n6915 GNDA.n231 76.3222
R9164 GNDA.n6912 GNDA.n232 76.3222
R9165 GNDA.n6908 GNDA.n233 76.3222
R9166 GNDA.n6904 GNDA.n234 76.3222
R9167 GNDA.n7141 GNDA.n130 76.3222
R9168 GNDA.n245 GNDA.n129 76.3222
R9169 GNDA.n249 GNDA.n128 76.3222
R9170 GNDA.n253 GNDA.n127 76.3222
R9171 GNDA.n257 GNDA.n126 76.3222
R9172 GNDA.n261 GNDA.n125 76.3222
R9173 GNDA.n688 GNDA.n124 76.3222
R9174 GNDA.n684 GNDA.n123 76.3222
R9175 GNDA.n680 GNDA.n122 76.3222
R9176 GNDA.n676 GNDA.n121 76.3222
R9177 GNDA.n672 GNDA.n120 76.3222
R9178 GNDA.n136 GNDA.n119 76.3222
R9179 GNDA.n848 GNDA.n118 76.3222
R9180 GNDA.n852 GNDA.n117 76.3222
R9181 GNDA.n856 GNDA.n116 76.3222
R9182 GNDA.n860 GNDA.n115 76.3222
R9183 GNDA.n864 GNDA.n114 76.3222
R9184 GNDA.n868 GNDA.n113 76.3222
R9185 GNDA.n7321 GNDA.n54 76.3222
R9186 GNDA.n7311 GNDA.n53 76.3222
R9187 GNDA.n7236 GNDA.n52 76.3222
R9188 GNDA.n7242 GNDA.n51 76.3222
R9189 GNDA.n7249 GNDA.n50 76.3222
R9190 GNDA.n7231 GNDA.n49 76.3222
R9191 GNDA.n7321 GNDA.n7320 76.3222
R9192 GNDA.n58 GNDA.n53 76.3222
R9193 GNDA.n7310 GNDA.n52 76.3222
R9194 GNDA.n7237 GNDA.n51 76.3222
R9195 GNDA.n7241 GNDA.n50 76.3222
R9196 GNDA.n7250 GNDA.n49 76.3222
R9197 GNDA.n6897 GNDA.n48 76.3222
R9198 GNDA.n6892 GNDA.n47 76.3222
R9199 GNDA.n6809 GNDA.n46 76.3222
R9200 GNDA.n6815 GNDA.n45 76.3222
R9201 GNDA.n6821 GNDA.n44 76.3222
R9202 GNDA.n6830 GNDA.n43 76.3222
R9203 GNDA.n325 GNDA.n324 76.3222
R9204 GNDA.n322 GNDA.n321 76.3222
R9205 GNDA.n317 GNDA.n316 76.3222
R9206 GNDA.n314 GNDA.n313 76.3222
R9207 GNDA.n309 GNDA.n308 76.3222
R9208 GNDA.n306 GNDA.n302 76.3222
R9209 GNDA.n349 GNDA.n348 76.3222
R9210 GNDA.n344 GNDA.n343 76.3222
R9211 GNDA.n341 GNDA.n340 76.3222
R9212 GNDA.n336 GNDA.n335 76.3222
R9213 GNDA.n333 GNDA.n332 76.3222
R9214 GNDA.n328 GNDA.n327 76.3222
R9215 GNDA.n159 GNDA.n151 76.3222
R9216 GNDA.n157 GNDA.n149 76.3222
R9217 GNDA.n156 GNDA.n147 76.3222
R9218 GNDA.n155 GNDA.n145 76.3222
R9219 GNDA.n154 GNDA.n143 76.3222
R9220 GNDA.n153 GNDA.n131 76.3222
R9221 GNDA.n7135 GNDA.n137 76.3222
R9222 GNDA.n7133 GNDA.n142 76.3222
R9223 GNDA.n7126 GNDA.n141 76.3222
R9224 GNDA.n7122 GNDA.n140 76.3222
R9225 GNDA.n7118 GNDA.n139 76.3222
R9226 GNDA.n7114 GNDA.n138 76.3222
R9227 GNDA.n6207 GNDA.n6206 76.3222
R9228 GNDA.n1116 GNDA.n590 76.3222
R9229 GNDA.n1115 GNDA.n1114 76.3222
R9230 GNDA.n1109 GNDA.n1108 76.3222
R9231 GNDA.n1106 GNDA.n1105 76.3222
R9232 GNDA.n1135 GNDA.n1134 76.3222
R9233 GNDA.n1132 GNDA.n1131 76.3222
R9234 GNDA.n1129 GNDA.n1128 76.3222
R9235 GNDA.n1124 GNDA.n1123 76.3222
R9236 GNDA.n1121 GNDA.n1120 76.3222
R9237 GNDA.n1111 GNDA.n588 76.3222
R9238 GNDA.n6212 GNDA.n6211 76.3222
R9239 GNDA.n1101 GNDA.n1100 76.3222
R9240 GNDA.n1096 GNDA.n916 76.3222
R9241 GNDA.n1094 GNDA.n1093 76.3222
R9242 GNDA.n1089 GNDA.n1088 76.3222
R9243 GNDA.n1086 GNDA.n1085 76.3222
R9244 GNDA.n1081 GNDA.n1080 76.3222
R9245 GNDA.n1160 GNDA.n907 76.3222
R9246 GNDA.n1158 GNDA.n1157 76.3222
R9247 GNDA.n1153 GNDA.n1152 76.3222
R9248 GNDA.n1150 GNDA.n1149 76.3222
R9249 GNDA.n1145 GNDA.n1144 76.3222
R9250 GNDA.n1142 GNDA.n1141 76.3222
R9251 GNDA.n1217 GNDA.n1216 76.3222
R9252 GNDA.n1212 GNDA.n1211 76.3222
R9253 GNDA.n1209 GNDA.n1208 76.3222
R9254 GNDA.n1204 GNDA.n1203 76.3222
R9255 GNDA.n1201 GNDA.n1200 76.3222
R9256 GNDA.n1196 GNDA.n1195 76.3222
R9257 GNDA.n7042 GNDA.n227 76.3222
R9258 GNDA.n7032 GNDA.n226 76.3222
R9259 GNDA.n6957 GNDA.n225 76.3222
R9260 GNDA.n6963 GNDA.n224 76.3222
R9261 GNDA.n6970 GNDA.n223 76.3222
R9262 GNDA.n6952 GNDA.n222 76.3222
R9263 GNDA.n7108 GNDA.n164 76.3222
R9264 GNDA.n200 GNDA.n167 76.3222
R9265 GNDA.n221 GNDA.n199 76.3222
R9266 GNDA.n210 GNDA.n198 76.3222
R9267 GNDA.n197 GNDA.n189 76.3222
R9268 GNDA.n7044 GNDA.n190 76.3222
R9269 GNDA.n805 GNDA.n196 76.3222
R9270 GNDA.n802 GNDA.n195 76.3222
R9271 GNDA.n795 GNDA.n194 76.3222
R9272 GNDA.n788 GNDA.n193 76.3222
R9273 GNDA.n815 GNDA.n192 76.3222
R9274 GNDA.n820 GNDA.n191 76.3222
R9275 GNDA.n6674 GNDA.n6630 76.3222
R9276 GNDA.n6670 GNDA.n6669 76.3222
R9277 GNDA.n6663 GNDA.n6634 76.3222
R9278 GNDA.n6662 GNDA.n6661 76.3222
R9279 GNDA.n6655 GNDA.n6642 76.3222
R9280 GNDA.n6654 GNDA.n6653 76.3222
R9281 GNDA.n42 GNDA.n24 76.3222
R9282 GNDA.n7323 GNDA.n25 76.3222
R9283 GNDA.n41 GNDA.n31 76.3222
R9284 GNDA.n7161 GNDA.n29 76.3222
R9285 GNDA.n7167 GNDA.n28 76.3222
R9286 GNDA.n7157 GNDA.n27 76.3222
R9287 GNDA.n7227 GNDA.n42 76.3222
R9288 GNDA.n7324 GNDA.n7323 76.3222
R9289 GNDA.n41 GNDA.n40 76.3222
R9290 GNDA.n30 GNDA.n29 76.3222
R9291 GNDA.n7162 GNDA.n28 76.3222
R9292 GNDA.n7168 GNDA.n27 76.3222
R9293 GNDA.n6650 GNDA.n6649 76.3222
R9294 GNDA.n6647 GNDA.n6646 76.3222
R9295 GNDA.n6644 GNDA.n6643 76.3222
R9296 GNDA.n6639 GNDA.n6638 76.3222
R9297 GNDA.n6636 GNDA.n6635 76.3222
R9298 GNDA.n6631 GNDA.n6628 76.3222
R9299 GNDA.n6671 GNDA.n6630 76.3222
R9300 GNDA.n6669 GNDA.n6668 76.3222
R9301 GNDA.n6664 GNDA.n6663 76.3222
R9302 GNDA.n6661 GNDA.n6660 76.3222
R9303 GNDA.n6656 GNDA.n6655 76.3222
R9304 GNDA.n6653 GNDA.n86 76.3222
R9305 GNDA.n899 GNDA.n898 76.3222
R9306 GNDA.n888 GNDA.n660 76.3222
R9307 GNDA.n887 GNDA.n886 76.3222
R9308 GNDA.n876 GNDA.n664 76.3222
R9309 GNDA.n875 GNDA.n874 76.3222
R9310 GNDA.n690 GNDA.n668 76.3222
R9311 GNDA.n871 GNDA.n870 76.3222
R9312 GNDA.n881 GNDA.n880 76.3222
R9313 GNDA.n882 GNDA.n662 76.3222
R9314 GNDA.n893 GNDA.n892 76.3222
R9315 GNDA.n894 GNDA.n658 76.3222
R9316 GNDA.n6218 GNDA.n6217 76.3222
R9317 GNDA.n1177 GNDA.n579 76.3222
R9318 GNDA.n1172 GNDA.n578 76.3222
R9319 GNDA.n1170 GNDA.n577 76.3222
R9320 GNDA.n1166 GNDA.n576 76.3222
R9321 GNDA.n1164 GNDA.n575 76.3222
R9322 GNDA.n1191 GNDA.n906 76.3222
R9323 GNDA.n1189 GNDA.n1188 76.3222
R9324 GNDA.n1184 GNDA.n1183 76.3222
R9325 GNDA.n1181 GNDA.n1180 76.3222
R9326 GNDA.n1174 GNDA.n572 76.3222
R9327 GNDA.n6222 GNDA.n6221 76.3222
R9328 GNDA.n1076 GNDA.n287 76.3222
R9329 GNDA.n1072 GNDA.n286 76.3222
R9330 GNDA.n1068 GNDA.n285 76.3222
R9331 GNDA.n1064 GNDA.n284 76.3222
R9332 GNDA.n1060 GNDA.n283 76.3222
R9333 GNDA.n265 GNDA.n236 76.3222
R9334 GNDA.n269 GNDA.n237 76.3222
R9335 GNDA.n273 GNDA.n238 76.3222
R9336 GNDA.n241 GNDA.n239 76.3222
R9337 GNDA.n280 GNDA.n240 76.3222
R9338 GNDA.n6921 GNDA.n289 76.3222
R9339 GNDA.n6913 GNDA.n231 76.3222
R9340 GNDA.n6909 GNDA.n232 76.3222
R9341 GNDA.n6905 GNDA.n233 76.3222
R9342 GNDA.n6901 GNDA.n234 76.3222
R9343 GNDA.n1237 GNDA.t174 75.3088
R9344 GNDA.n6754 GNDA.n301 74.8124
R9345 GNDA.n6727 GNDA.n6726 74.8124
R9346 GNDA.n1271 GNDA.n1251 74.5978
R9347 GNDA.n1272 GNDA.n1271 74.5978
R9348 GNDA.n6148 GNDA.n6147 74.5978
R9349 GNDA.n6147 GNDA.n6146 74.5978
R9350 GNDA.n7068 GNDA.n176 74.5978
R9351 GNDA.n7065 GNDA.n176 74.5978
R9352 GNDA.n6853 GNDA.n6792 74.5978
R9353 GNDA.n6850 GNDA.n6792 74.5978
R9354 GNDA.n747 GNDA.n716 74.5978
R9355 GNDA.n744 GNDA.n716 74.5978
R9356 GNDA.n6994 GNDA.n6939 74.5978
R9357 GNDA.n6991 GNDA.n6939 74.5978
R9358 GNDA.n7273 GNDA.n70 74.5978
R9359 GNDA.n7270 GNDA.n70 74.5978
R9360 GNDA.n1001 GNDA.n940 74.5978
R9361 GNDA.n1002 GNDA.n1001 74.5978
R9362 GNDA.n7191 GNDA.n9 74.5978
R9363 GNDA.n7188 GNDA.n9 74.5978
R9364 GNDA.n1312 GNDA.n1311 69.3109
R9365 GNDA.n1311 GNDA.n1310 69.3109
R9366 GNDA.n6183 GNDA.n6182 69.3109
R9367 GNDA.n6182 GNDA.n6181 69.3109
R9368 GNDA.n7102 GNDA.n169 69.3109
R9369 GNDA.n7102 GNDA.n7101 69.3109
R9370 GNDA.n6887 GNDA.n6785 69.3109
R9371 GNDA.n6887 GNDA.n6886 69.3109
R9372 GNDA.n810 GNDA.n809 69.3109
R9373 GNDA.n810 GNDA.n728 69.3109
R9374 GNDA.n7036 GNDA.n6929 69.3109
R9375 GNDA.n7012 GNDA.n6929 69.3109
R9376 GNDA.n7315 GNDA.n60 69.3109
R9377 GNDA.n7291 GNDA.n60 69.3109
R9378 GNDA.n1042 GNDA.n1039 69.3109
R9379 GNDA.n1039 GNDA.n1038 69.3109
R9380 GNDA.n7328 GNDA.n7327 69.3109
R9381 GNDA.n7328 GNDA.n20 69.3109
R9382 GNDA.n6190 GNDA.t172 68.664
R9383 GNDA.n1238 GNDA.t168 68.664
R9384 GNDA.n1293 GNDA.t841 65.8183
R9385 GNDA.n1295 GNDA.t841 65.8183
R9386 GNDA.n1301 GNDA.t841 65.8183
R9387 GNDA.n1303 GNDA.t841 65.8183
R9388 GNDA.n1277 GNDA.t841 65.8183
R9389 GNDA.n1279 GNDA.t841 65.8183
R9390 GNDA.n1285 GNDA.t841 65.8183
R9391 GNDA.n1287 GNDA.t841 65.8183
R9392 GNDA.n1256 GNDA.t841 65.8183
R9393 GNDA.n1262 GNDA.t841 65.8183
R9394 GNDA.n1255 GNDA.t841 65.8183
R9395 GNDA.n1269 GNDA.t841 65.8183
R9396 GNDA.n6255 GNDA.t841 65.8183
R9397 GNDA.n6252 GNDA.t841 65.8183
R9398 GNDA.n1313 GNDA.t841 65.8183
R9399 GNDA.n1326 GNDA.t841 65.8183
R9400 GNDA.n6165 GNDA.t821 65.8183
R9401 GNDA.n6171 GNDA.t821 65.8183
R9402 GNDA.n6173 GNDA.t821 65.8183
R9403 GNDA.n6179 GNDA.t821 65.8183
R9404 GNDA.n6149 GNDA.t821 65.8183
R9405 GNDA.n6155 GNDA.t821 65.8183
R9406 GNDA.n6157 GNDA.t821 65.8183
R9407 GNDA.n6163 GNDA.t821 65.8183
R9408 GNDA.n6133 GNDA.t821 65.8183
R9409 GNDA.n619 GNDA.t821 65.8183
R9410 GNDA.n6140 GNDA.t821 65.8183
R9411 GNDA.n616 GNDA.t821 65.8183
R9412 GNDA.n6129 GNDA.t821 65.8183
R9413 GNDA.n6115 GNDA.t821 65.8183
R9414 GNDA.n6113 GNDA.t821 65.8183
R9415 GNDA.n6185 GNDA.t821 65.8183
R9416 GNDA.t744 GNDA.n186 65.8183
R9417 GNDA.t744 GNDA.n185 65.8183
R9418 GNDA.t744 GNDA.n184 65.8183
R9419 GNDA.t744 GNDA.n183 65.8183
R9420 GNDA.t744 GNDA.n174 65.8183
R9421 GNDA.t744 GNDA.n181 65.8183
R9422 GNDA.t744 GNDA.n171 65.8183
R9423 GNDA.t744 GNDA.n182 65.8183
R9424 GNDA.t744 GNDA.n180 65.8183
R9425 GNDA.t744 GNDA.n179 65.8183
R9426 GNDA.t744 GNDA.n178 65.8183
R9427 GNDA.t744 GNDA.n177 65.8183
R9428 GNDA.t744 GNDA.n175 65.8183
R9429 GNDA.t744 GNDA.n173 65.8183
R9430 GNDA.t744 GNDA.n172 65.8183
R9431 GNDA.n7103 GNDA.t744 65.8183
R9432 GNDA.t786 GNDA.n6802 65.8183
R9433 GNDA.t786 GNDA.n6801 65.8183
R9434 GNDA.t786 GNDA.n6800 65.8183
R9435 GNDA.t786 GNDA.n6799 65.8183
R9436 GNDA.t786 GNDA.n6790 65.8183
R9437 GNDA.t786 GNDA.n6797 65.8183
R9438 GNDA.t786 GNDA.n6787 65.8183
R9439 GNDA.t786 GNDA.n6798 65.8183
R9440 GNDA.t786 GNDA.n6796 65.8183
R9441 GNDA.t786 GNDA.n6795 65.8183
R9442 GNDA.t786 GNDA.n6794 65.8183
R9443 GNDA.t786 GNDA.n6793 65.8183
R9444 GNDA.t742 GNDA.n727 65.8183
R9445 GNDA.t742 GNDA.n726 65.8183
R9446 GNDA.t742 GNDA.n725 65.8183
R9447 GNDA.t742 GNDA.n724 65.8183
R9448 GNDA.t742 GNDA.n715 65.8183
R9449 GNDA.t742 GNDA.n722 65.8183
R9450 GNDA.t742 GNDA.n712 65.8183
R9451 GNDA.t742 GNDA.n723 65.8183
R9452 GNDA.t742 GNDA.n721 65.8183
R9453 GNDA.t742 GNDA.n719 65.8183
R9454 GNDA.t742 GNDA.n718 65.8183
R9455 GNDA.t742 GNDA.n717 65.8183
R9456 GNDA.n811 GNDA.t742 65.8183
R9457 GNDA.t742 GNDA.n714 65.8183
R9458 GNDA.t742 GNDA.n713 65.8183
R9459 GNDA.t742 GNDA.n711 65.8183
R9460 GNDA.t840 GNDA.n7026 65.8183
R9461 GNDA.t840 GNDA.n6948 65.8183
R9462 GNDA.t840 GNDA.n6947 65.8183
R9463 GNDA.t840 GNDA.n6946 65.8183
R9464 GNDA.t840 GNDA.n6937 65.8183
R9465 GNDA.t840 GNDA.n6944 65.8183
R9466 GNDA.t840 GNDA.n6935 65.8183
R9467 GNDA.t840 GNDA.n6945 65.8183
R9468 GNDA.t840 GNDA.n6943 65.8183
R9469 GNDA.t840 GNDA.n6942 65.8183
R9470 GNDA.t840 GNDA.n6941 65.8183
R9471 GNDA.t840 GNDA.n6940 65.8183
R9472 GNDA.t840 GNDA.n6938 65.8183
R9473 GNDA.t840 GNDA.n6936 65.8183
R9474 GNDA.n7027 GNDA.t840 65.8183
R9475 GNDA.t840 GNDA.n6930 65.8183
R9476 GNDA.t845 GNDA.n7305 65.8183
R9477 GNDA.t845 GNDA.n79 65.8183
R9478 GNDA.t845 GNDA.n78 65.8183
R9479 GNDA.t845 GNDA.n77 65.8183
R9480 GNDA.t845 GNDA.n68 65.8183
R9481 GNDA.t845 GNDA.n75 65.8183
R9482 GNDA.t845 GNDA.n66 65.8183
R9483 GNDA.t845 GNDA.n76 65.8183
R9484 GNDA.t845 GNDA.n74 65.8183
R9485 GNDA.t845 GNDA.n73 65.8183
R9486 GNDA.t845 GNDA.n72 65.8183
R9487 GNDA.t845 GNDA.n71 65.8183
R9488 GNDA.t845 GNDA.n69 65.8183
R9489 GNDA.t845 GNDA.n67 65.8183
R9490 GNDA.n7306 GNDA.t845 65.8183
R9491 GNDA.t845 GNDA.n61 65.8183
R9492 GNDA.t786 GNDA.n6791 65.8183
R9493 GNDA.t786 GNDA.n6789 65.8183
R9494 GNDA.t786 GNDA.n6788 65.8183
R9495 GNDA.n6888 GNDA.t786 65.8183
R9496 GNDA.n1023 GNDA.t751 65.8183
R9497 GNDA.n1025 GNDA.t751 65.8183
R9498 GNDA.n1031 GNDA.t751 65.8183
R9499 GNDA.n1033 GNDA.t751 65.8183
R9500 GNDA.n1007 GNDA.t751 65.8183
R9501 GNDA.n1009 GNDA.t751 65.8183
R9502 GNDA.n1015 GNDA.t751 65.8183
R9503 GNDA.n1017 GNDA.t751 65.8183
R9504 GNDA.n987 GNDA.t751 65.8183
R9505 GNDA.n992 GNDA.t751 65.8183
R9506 GNDA.n944 GNDA.t751 65.8183
R9507 GNDA.n999 GNDA.t751 65.8183
R9508 GNDA.n984 GNDA.t751 65.8183
R9509 GNDA.n970 GNDA.t751 65.8183
R9510 GNDA.n968 GNDA.t751 65.8183
R9511 GNDA.n1044 GNDA.t751 65.8183
R9512 GNDA.t764 GNDA.n19 65.8183
R9513 GNDA.t764 GNDA.n18 65.8183
R9514 GNDA.t764 GNDA.n17 65.8183
R9515 GNDA.t764 GNDA.n16 65.8183
R9516 GNDA.t764 GNDA.n7 65.8183
R9517 GNDA.t764 GNDA.n14 65.8183
R9518 GNDA.t764 GNDA.n5 65.8183
R9519 GNDA.t764 GNDA.n15 65.8183
R9520 GNDA.t764 GNDA.n13 65.8183
R9521 GNDA.t764 GNDA.n12 65.8183
R9522 GNDA.t764 GNDA.n11 65.8183
R9523 GNDA.t764 GNDA.n10 65.8183
R9524 GNDA.t764 GNDA.n8 65.8183
R9525 GNDA.n7329 GNDA.t764 65.8183
R9526 GNDA.t764 GNDA.n6 65.8183
R9527 GNDA.t764 GNDA.n4 65.8183
R9528 GNDA.n6202 GNDA.t109 64.2341
R9529 GNDA.n6122 GNDA.t111 64.2341
R9530 GNDA.n585 GNDA.n560 63.1266
R9531 GNDA.n6228 GNDA.n564 63.1266
R9532 GNDA.n4108 GNDA.t760 62.2505
R9533 GNDA.n4117 GNDA.t750 62.2505
R9534 GNDA.n1815 GNDA.t757 62.2505
R9535 GNDA.n4111 GNDA.t773 62.2505
R9536 GNDA.n4783 GNDA.t741 62.2505
R9537 GNDA.n4128 GNDA.t833 62.2505
R9538 GNDA.n4794 GNDA.t817 62.2505
R9539 GNDA.n4787 GNDA.t792 62.2505
R9540 GNDA.n1590 GNDA.t770 62.2505
R9541 GNDA.n4135 GNDA.t814 62.2505
R9542 GNDA.n4131 GNDA.t785 62.2505
R9543 GNDA.n4089 GNDA.t798 62.2505
R9544 GNDA.n1365 GNDA.n1348 59.2425
R9545 GNDA.n4800 GNDA.n4799 59.2425
R9546 GNDA.n4087 GNDA.n4086 59.2425
R9547 GNDA.n3461 GNDA.n1817 59.2425
R9548 GNDA.n585 GNDA.n583 58.6967
R9549 GNDA.n6229 GNDA.n6228 58.6967
R9550 GNDA.n1311 GNDA.t841 57.8461
R9551 GNDA.n6182 GNDA.t821 57.8461
R9552 GNDA.t744 GNDA.n7102 57.8461
R9553 GNDA.t742 GNDA.n810 57.8461
R9554 GNDA.t840 GNDA.n6929 57.8461
R9555 GNDA.t845 GNDA.n60 57.8461
R9556 GNDA.t786 GNDA.n6887 57.8461
R9557 GNDA.n1039 GNDA.t751 57.8461
R9558 GNDA.t764 GNDA.n7328 57.8461
R9559 GNDA.t117 GNDA.n6202 57.5892
R9560 GNDA.t781 GNDA.n6122 57.5892
R9561 GNDA.t775 GNDA.n6246 57.5892
R9562 GNDA.n640 GNDA.n637 56.3995
R9563 GNDA.n822 GNDA.n705 56.3995
R9564 GNDA.n6924 GNDA.n6923 56.3995
R9565 GNDA.n6900 GNDA.n235 56.3995
R9566 GNDA.n637 GNDA.n635 56.3995
R9567 GNDA.n822 GNDA.n821 56.3995
R9568 GNDA.n7155 GNDA.n7154 56.3995
R9569 GNDA.n7156 GNDA.n7155 56.3995
R9570 GNDA.n921 GNDA.n281 56.3995
R9571 GNDA.n6923 GNDA.n228 56.3995
R9572 GNDA.n6898 GNDA.n235 56.3995
R9573 GNDA.n1271 GNDA.t841 55.2026
R9574 GNDA.n6147 GNDA.t821 55.2026
R9575 GNDA.t744 GNDA.n176 55.2026
R9576 GNDA.t786 GNDA.n6792 55.2026
R9577 GNDA.t742 GNDA.n716 55.2026
R9578 GNDA.t840 GNDA.n6939 55.2026
R9579 GNDA.t845 GNDA.n70 55.2026
R9580 GNDA.n1001 GNDA.t751 55.2026
R9581 GNDA.t764 GNDA.n9 55.2026
R9582 GNDA.t877 GNDA.t143 55.1153
R9583 GNDA.t446 GNDA.n1343 54.2977
R9584 GNDA.n1287 GNDA.n1247 53.3664
R9585 GNDA.n1286 GNDA.n1285 53.3664
R9586 GNDA.n1279 GNDA.n1249 53.3664
R9587 GNDA.n1278 GNDA.n1277 53.3664
R9588 GNDA.n1269 GNDA.n1268 53.3664
R9589 GNDA.n1264 GNDA.n1255 53.3664
R9590 GNDA.n1262 GNDA.n1261 53.3664
R9591 GNDA.n1256 GNDA.n547 53.3664
R9592 GNDA.n1327 GNDA.n1326 53.3664
R9593 GNDA.n1314 GNDA.n1313 53.3664
R9594 GNDA.n6252 GNDA.n6251 53.3664
R9595 GNDA.n6255 GNDA.n6254 53.3664
R9596 GNDA.n1294 GNDA.n1293 53.3664
R9597 GNDA.n1296 GNDA.n1295 53.3664
R9598 GNDA.n1301 GNDA.n1300 53.3664
R9599 GNDA.n1304 GNDA.n1303 53.3664
R9600 GNDA.n1293 GNDA.n1292 53.3664
R9601 GNDA.n1295 GNDA.n1245 53.3664
R9602 GNDA.n1302 GNDA.n1301 53.3664
R9603 GNDA.n1303 GNDA.n1243 53.3664
R9604 GNDA.n1277 GNDA.n1276 53.3664
R9605 GNDA.n1280 GNDA.n1279 53.3664
R9606 GNDA.n1285 GNDA.n1284 53.3664
R9607 GNDA.n1288 GNDA.n1287 53.3664
R9608 GNDA.n1257 GNDA.n1256 53.3664
R9609 GNDA.n1263 GNDA.n1262 53.3664
R9610 GNDA.n1255 GNDA.n1253 53.3664
R9611 GNDA.n1270 GNDA.n1269 53.3664
R9612 GNDA.n6256 GNDA.n6255 53.3664
R9613 GNDA.n6253 GNDA.n6252 53.3664
R9614 GNDA.n1313 GNDA.n550 53.3664
R9615 GNDA.n1326 GNDA.n1325 53.3664
R9616 GNDA.n6164 GNDA.n6163 53.3664
R9617 GNDA.n6157 GNDA.n610 53.3664
R9618 GNDA.n6156 GNDA.n6155 53.3664
R9619 GNDA.n6149 GNDA.n612 53.3664
R9620 GNDA.n6142 GNDA.n616 53.3664
R9621 GNDA.n6140 GNDA.n6139 53.3664
R9622 GNDA.n6135 GNDA.n619 53.3664
R9623 GNDA.n6133 GNDA.n6132 53.3664
R9624 GNDA.n6185 GNDA.n6184 53.3664
R9625 GNDA.n6113 GNDA.n604 53.3664
R9626 GNDA.n6116 GNDA.n6115 53.3664
R9627 GNDA.n6129 GNDA.n6128 53.3664
R9628 GNDA.n6165 GNDA.n608 53.3664
R9629 GNDA.n6171 GNDA.n6170 53.3664
R9630 GNDA.n6174 GNDA.n6173 53.3664
R9631 GNDA.n6179 GNDA.n6178 53.3664
R9632 GNDA.n6166 GNDA.n6165 53.3664
R9633 GNDA.n6172 GNDA.n6171 53.3664
R9634 GNDA.n6173 GNDA.n606 53.3664
R9635 GNDA.n6180 GNDA.n6179 53.3664
R9636 GNDA.n6150 GNDA.n6149 53.3664
R9637 GNDA.n6155 GNDA.n6154 53.3664
R9638 GNDA.n6158 GNDA.n6157 53.3664
R9639 GNDA.n6163 GNDA.n6162 53.3664
R9640 GNDA.n6134 GNDA.n6133 53.3664
R9641 GNDA.n619 GNDA.n617 53.3664
R9642 GNDA.n6141 GNDA.n6140 53.3664
R9643 GNDA.n616 GNDA.n614 53.3664
R9644 GNDA.n6130 GNDA.n6129 53.3664
R9645 GNDA.n6115 GNDA.n622 53.3664
R9646 GNDA.n6114 GNDA.n6113 53.3664
R9647 GNDA.n6186 GNDA.n6185 53.3664
R9648 GNDA.n7084 GNDA.n182 53.3664
R9649 GNDA.n7080 GNDA.n171 53.3664
R9650 GNDA.n7076 GNDA.n181 53.3664
R9651 GNDA.n7072 GNDA.n174 53.3664
R9652 GNDA.n7061 GNDA.n177 53.3664
R9653 GNDA.n7057 GNDA.n178 53.3664
R9654 GNDA.n7053 GNDA.n179 53.3664
R9655 GNDA.n7049 GNDA.n180 53.3664
R9656 GNDA.n7104 GNDA.n7103 53.3664
R9657 GNDA.n217 GNDA.n172 53.3664
R9658 GNDA.n213 GNDA.n173 53.3664
R9659 GNDA.n206 GNDA.n175 53.3664
R9660 GNDA.n7088 GNDA.n186 53.3664
R9661 GNDA.n7089 GNDA.n185 53.3664
R9662 GNDA.n7093 GNDA.n184 53.3664
R9663 GNDA.n7097 GNDA.n183 53.3664
R9664 GNDA.n7085 GNDA.n186 53.3664
R9665 GNDA.n7092 GNDA.n185 53.3664
R9666 GNDA.n7096 GNDA.n184 53.3664
R9667 GNDA.n7100 GNDA.n183 53.3664
R9668 GNDA.n7069 GNDA.n174 53.3664
R9669 GNDA.n7073 GNDA.n181 53.3664
R9670 GNDA.n7077 GNDA.n171 53.3664
R9671 GNDA.n7081 GNDA.n182 53.3664
R9672 GNDA.n7052 GNDA.n180 53.3664
R9673 GNDA.n7056 GNDA.n179 53.3664
R9674 GNDA.n7060 GNDA.n178 53.3664
R9675 GNDA.n7064 GNDA.n177 53.3664
R9676 GNDA.n7048 GNDA.n175 53.3664
R9677 GNDA.n205 GNDA.n173 53.3664
R9678 GNDA.n214 GNDA.n172 53.3664
R9679 GNDA.n7103 GNDA.n170 53.3664
R9680 GNDA.n6869 GNDA.n6798 53.3664
R9681 GNDA.n6865 GNDA.n6787 53.3664
R9682 GNDA.n6861 GNDA.n6797 53.3664
R9683 GNDA.n6857 GNDA.n6790 53.3664
R9684 GNDA.n6846 GNDA.n6793 53.3664
R9685 GNDA.n6842 GNDA.n6794 53.3664
R9686 GNDA.n6838 GNDA.n6795 53.3664
R9687 GNDA.n6834 GNDA.n6796 53.3664
R9688 GNDA.n6889 GNDA.n6888 53.3664
R9689 GNDA.n6811 GNDA.n6788 53.3664
R9690 GNDA.n6819 GNDA.n6789 53.3664
R9691 GNDA.n6826 GNDA.n6791 53.3664
R9692 GNDA.n6873 GNDA.n6802 53.3664
R9693 GNDA.n6874 GNDA.n6801 53.3664
R9694 GNDA.n6878 GNDA.n6800 53.3664
R9695 GNDA.n6882 GNDA.n6799 53.3664
R9696 GNDA.n6870 GNDA.n6802 53.3664
R9697 GNDA.n6877 GNDA.n6801 53.3664
R9698 GNDA.n6881 GNDA.n6800 53.3664
R9699 GNDA.n6885 GNDA.n6799 53.3664
R9700 GNDA.n6854 GNDA.n6790 53.3664
R9701 GNDA.n6858 GNDA.n6797 53.3664
R9702 GNDA.n6862 GNDA.n6787 53.3664
R9703 GNDA.n6866 GNDA.n6798 53.3664
R9704 GNDA.n6837 GNDA.n6796 53.3664
R9705 GNDA.n6841 GNDA.n6795 53.3664
R9706 GNDA.n6845 GNDA.n6794 53.3664
R9707 GNDA.n6849 GNDA.n6793 53.3664
R9708 GNDA.n763 GNDA.n723 53.3664
R9709 GNDA.n759 GNDA.n712 53.3664
R9710 GNDA.n755 GNDA.n722 53.3664
R9711 GNDA.n751 GNDA.n715 53.3664
R9712 GNDA.n740 GNDA.n717 53.3664
R9713 GNDA.n736 GNDA.n718 53.3664
R9714 GNDA.n732 GNDA.n719 53.3664
R9715 GNDA.n721 GNDA.n720 53.3664
R9716 GNDA.n729 GNDA.n711 53.3664
R9717 GNDA.n798 GNDA.n713 53.3664
R9718 GNDA.n791 GNDA.n714 53.3664
R9719 GNDA.n812 GNDA.n811 53.3664
R9720 GNDA.n767 GNDA.n727 53.3664
R9721 GNDA.n768 GNDA.n726 53.3664
R9722 GNDA.n772 GNDA.n725 53.3664
R9723 GNDA.n776 GNDA.n724 53.3664
R9724 GNDA.n764 GNDA.n727 53.3664
R9725 GNDA.n771 GNDA.n726 53.3664
R9726 GNDA.n775 GNDA.n725 53.3664
R9727 GNDA.n778 GNDA.n724 53.3664
R9728 GNDA.n748 GNDA.n715 53.3664
R9729 GNDA.n752 GNDA.n722 53.3664
R9730 GNDA.n756 GNDA.n712 53.3664
R9731 GNDA.n760 GNDA.n723 53.3664
R9732 GNDA.n731 GNDA.n721 53.3664
R9733 GNDA.n735 GNDA.n719 53.3664
R9734 GNDA.n739 GNDA.n718 53.3664
R9735 GNDA.n743 GNDA.n717 53.3664
R9736 GNDA.n811 GNDA.n710 53.3664
R9737 GNDA.n714 GNDA.n709 53.3664
R9738 GNDA.n790 GNDA.n713 53.3664
R9739 GNDA.n797 GNDA.n711 53.3664
R9740 GNDA.n7009 GNDA.n6945 53.3664
R9741 GNDA.n7006 GNDA.n6935 53.3664
R9742 GNDA.n7002 GNDA.n6944 53.3664
R9743 GNDA.n6998 GNDA.n6937 53.3664
R9744 GNDA.n6987 GNDA.n6940 53.3664
R9745 GNDA.n6983 GNDA.n6941 53.3664
R9746 GNDA.n6979 GNDA.n6942 53.3664
R9747 GNDA.n6975 GNDA.n6943 53.3664
R9748 GNDA.n7035 GNDA.n6930 53.3664
R9749 GNDA.n7028 GNDA.n7027 53.3664
R9750 GNDA.n6960 GNDA.n6936 53.3664
R9751 GNDA.n6967 GNDA.n6938 53.3664
R9752 GNDA.n7026 GNDA.n7025 53.3664
R9753 GNDA.n6950 GNDA.n6948 53.3664
R9754 GNDA.n7020 GNDA.n6947 53.3664
R9755 GNDA.n7016 GNDA.n6946 53.3664
R9756 GNDA.n7026 GNDA.n6949 53.3664
R9757 GNDA.n7021 GNDA.n6948 53.3664
R9758 GNDA.n7017 GNDA.n6947 53.3664
R9759 GNDA.n7013 GNDA.n6946 53.3664
R9760 GNDA.n6995 GNDA.n6937 53.3664
R9761 GNDA.n6999 GNDA.n6944 53.3664
R9762 GNDA.n7003 GNDA.n6935 53.3664
R9763 GNDA.n7007 GNDA.n6945 53.3664
R9764 GNDA.n6978 GNDA.n6943 53.3664
R9765 GNDA.n6982 GNDA.n6942 53.3664
R9766 GNDA.n6986 GNDA.n6941 53.3664
R9767 GNDA.n6990 GNDA.n6940 53.3664
R9768 GNDA.n6974 GNDA.n6938 53.3664
R9769 GNDA.n6966 GNDA.n6936 53.3664
R9770 GNDA.n7027 GNDA.n6934 53.3664
R9771 GNDA.n6933 GNDA.n6930 53.3664
R9772 GNDA.n7288 GNDA.n76 53.3664
R9773 GNDA.n7285 GNDA.n66 53.3664
R9774 GNDA.n7281 GNDA.n75 53.3664
R9775 GNDA.n7277 GNDA.n68 53.3664
R9776 GNDA.n7266 GNDA.n71 53.3664
R9777 GNDA.n7262 GNDA.n72 53.3664
R9778 GNDA.n7258 GNDA.n73 53.3664
R9779 GNDA.n7254 GNDA.n74 53.3664
R9780 GNDA.n7314 GNDA.n61 53.3664
R9781 GNDA.n7307 GNDA.n7306 53.3664
R9782 GNDA.n7239 GNDA.n67 53.3664
R9783 GNDA.n7246 GNDA.n69 53.3664
R9784 GNDA.n7305 GNDA.n7304 53.3664
R9785 GNDA.n81 GNDA.n79 53.3664
R9786 GNDA.n7299 GNDA.n78 53.3664
R9787 GNDA.n7295 GNDA.n77 53.3664
R9788 GNDA.n7305 GNDA.n80 53.3664
R9789 GNDA.n7300 GNDA.n79 53.3664
R9790 GNDA.n7296 GNDA.n78 53.3664
R9791 GNDA.n7292 GNDA.n77 53.3664
R9792 GNDA.n7274 GNDA.n68 53.3664
R9793 GNDA.n7278 GNDA.n75 53.3664
R9794 GNDA.n7282 GNDA.n66 53.3664
R9795 GNDA.n7286 GNDA.n76 53.3664
R9796 GNDA.n7257 GNDA.n74 53.3664
R9797 GNDA.n7261 GNDA.n73 53.3664
R9798 GNDA.n7265 GNDA.n72 53.3664
R9799 GNDA.n7269 GNDA.n71 53.3664
R9800 GNDA.n7253 GNDA.n69 53.3664
R9801 GNDA.n7245 GNDA.n67 53.3664
R9802 GNDA.n7306 GNDA.n65 53.3664
R9803 GNDA.n64 GNDA.n61 53.3664
R9804 GNDA.n6833 GNDA.n6791 53.3664
R9805 GNDA.n6825 GNDA.n6789 53.3664
R9806 GNDA.n6818 GNDA.n6788 53.3664
R9807 GNDA.n6888 GNDA.n6786 53.3664
R9808 GNDA.n1017 GNDA.n936 53.3664
R9809 GNDA.n1016 GNDA.n1015 53.3664
R9810 GNDA.n1009 GNDA.n938 53.3664
R9811 GNDA.n1008 GNDA.n1007 53.3664
R9812 GNDA.n999 GNDA.n998 53.3664
R9813 GNDA.n994 GNDA.n944 53.3664
R9814 GNDA.n992 GNDA.n991 53.3664
R9815 GNDA.n987 GNDA.n986 53.3664
R9816 GNDA.n1044 GNDA.n1043 53.3664
R9817 GNDA.n968 GNDA.n931 53.3664
R9818 GNDA.n971 GNDA.n970 53.3664
R9819 GNDA.n984 GNDA.n983 53.3664
R9820 GNDA.n1024 GNDA.n1023 53.3664
R9821 GNDA.n1026 GNDA.n1025 53.3664
R9822 GNDA.n1031 GNDA.n1030 53.3664
R9823 GNDA.n1034 GNDA.n1033 53.3664
R9824 GNDA.n1023 GNDA.n1022 53.3664
R9825 GNDA.n1025 GNDA.n934 53.3664
R9826 GNDA.n1032 GNDA.n1031 53.3664
R9827 GNDA.n1033 GNDA.n932 53.3664
R9828 GNDA.n1007 GNDA.n1006 53.3664
R9829 GNDA.n1010 GNDA.n1009 53.3664
R9830 GNDA.n1015 GNDA.n1014 53.3664
R9831 GNDA.n1018 GNDA.n1017 53.3664
R9832 GNDA.n988 GNDA.n987 53.3664
R9833 GNDA.n993 GNDA.n992 53.3664
R9834 GNDA.n944 GNDA.n942 53.3664
R9835 GNDA.n1000 GNDA.n999 53.3664
R9836 GNDA.n985 GNDA.n984 53.3664
R9837 GNDA.n970 GNDA.n945 53.3664
R9838 GNDA.n969 GNDA.n968 53.3664
R9839 GNDA.n1045 GNDA.n1044 53.3664
R9840 GNDA.n7207 GNDA.n15 53.3664
R9841 GNDA.n7203 GNDA.n5 53.3664
R9842 GNDA.n7199 GNDA.n14 53.3664
R9843 GNDA.n7195 GNDA.n7 53.3664
R9844 GNDA.n7184 GNDA.n10 53.3664
R9845 GNDA.n7180 GNDA.n11 53.3664
R9846 GNDA.n7176 GNDA.n12 53.3664
R9847 GNDA.n7172 GNDA.n13 53.3664
R9848 GNDA.n21 GNDA.n4 53.3664
R9849 GNDA.n37 GNDA.n6 53.3664
R9850 GNDA.n7330 GNDA.n7329 53.3664
R9851 GNDA.n7164 GNDA.n8 53.3664
R9852 GNDA.n7211 GNDA.n19 53.3664
R9853 GNDA.n7212 GNDA.n18 53.3664
R9854 GNDA.n7216 GNDA.n17 53.3664
R9855 GNDA.n7220 GNDA.n16 53.3664
R9856 GNDA.n7208 GNDA.n19 53.3664
R9857 GNDA.n7215 GNDA.n18 53.3664
R9858 GNDA.n7219 GNDA.n17 53.3664
R9859 GNDA.n7222 GNDA.n16 53.3664
R9860 GNDA.n7192 GNDA.n7 53.3664
R9861 GNDA.n7196 GNDA.n14 53.3664
R9862 GNDA.n7200 GNDA.n5 53.3664
R9863 GNDA.n7204 GNDA.n15 53.3664
R9864 GNDA.n7175 GNDA.n13 53.3664
R9865 GNDA.n7179 GNDA.n12 53.3664
R9866 GNDA.n7183 GNDA.n11 53.3664
R9867 GNDA.n7187 GNDA.n10 53.3664
R9868 GNDA.n7171 GNDA.n8 53.3664
R9869 GNDA.n7329 GNDA.n3 53.3664
R9870 GNDA.n6 GNDA.n2 53.3664
R9871 GNDA.n36 GNDA.n4 53.3664
R9872 GNDA.t778 GNDA.n107 53.1593
R9873 GNDA.t829 GNDA.n6190 53.1593
R9874 GNDA.n1238 GNDA.t115 53.1593
R9875 GNDA.t743 GNDA.n107 52.0518
R9876 GNDA.t465 GNDA.n570 52.0518
R9877 GNDA.n6204 GNDA.t728 50.9444
R9878 GNDA.n4090 GNDA.t797 49.5418
R9879 GNDA.n4795 GNDA.t816 49.5418
R9880 GNDA.t28 GNDA.n6094 49.4893
R9881 GNDA.t871 GNDA.n4099 49.4893
R9882 GNDA.n580 GNDA.n564 48.7294
R9883 GNDA.t743 GNDA.n7142 47.6748
R9884 GNDA.n6214 GNDA.n583 47.6219
R9885 GNDA.n6246 GNDA.t743 47.6219
R9886 GNDA.n6191 GNDA.t829 46.5145
R9887 GNDA.t115 GNDA.n1237 46.5145
R9888 GNDA.n6108 GNDA.t41 45.407
R9889 GNDA.t743 GNDA.n102 44.3072
R9890 GNDA.t819 GNDA.n1817 42.2023
R9891 GNDA.t838 GNDA.n1348 42.2023
R9892 GNDA.n6203 GNDA.t117 42.0846
R9893 GNDA.n6104 GNDA.n6103 42.0846
R9894 GNDA.n6124 GNDA.t781 42.0846
R9895 GNDA.n927 GNDA.t58 40.9771
R9896 GNDA.n4139 GNDA.t836 40.4338
R9897 GNDA.n1594 GNDA.t768 40.4338
R9898 GNDA.n4119 GNDA.t795 40.4338
R9899 GNDA.n4125 GNDA.t754 40.4338
R9900 GNDA.t129 GNDA.t864 40.3675
R9901 GNDA.t90 GNDA.t26 40.3675
R9902 GNDA.t93 GNDA.t863 40.3675
R9903 GNDA.t852 GNDA.t106 40.3675
R9904 GNDA.t746 GNDA.t121 40.3675
R9905 GNDA.t797 GNDA.t105 40.3675
R9906 GNDA.t105 GNDA.t100 40.3675
R9907 GNDA.t100 GNDA.t76 40.3675
R9908 GNDA.t156 GNDA.t813 40.3675
R9909 GNDA.t813 GNDA.t98 40.3675
R9910 GNDA.t45 GNDA.t54 40.3675
R9911 GNDA.t144 GNDA.t50 40.3675
R9912 GNDA.t50 GNDA.t816 40.3675
R9913 GNDA.t800 GNDA.t848 40.3675
R9914 GNDA.t126 GNDA.t847 40.3675
R9915 GNDA.t139 GNDA.t47 40.3675
R9916 GNDA.t136 GNDA.t127 40.3675
R9917 GNDA.t134 GNDA.t13 40.3675
R9918 GNDA.n843 GNDA.t51 40.1125
R9919 GNDA.n6243 GNDA.n6231 39.3903
R9920 GNDA.n6231 GNDA.n559 39.3903
R9921 GNDA.t728 GNDA.t788 38.7621
R9922 GNDA.t826 GNDA.t465 38.7621
R9923 GNDA.t27 GNDA.t107 38.5326
R9924 GNDA.t36 GNDA.n4129 38.5326
R9925 GNDA.t19 GNDA.t853 38.5326
R9926 GNDA.n4141 GNDA.n4140 37.5297
R9927 GNDA.n4143 GNDA.n4142 37.5297
R9928 GNDA.n4145 GNDA.n4144 37.5297
R9929 GNDA.n4147 GNDA.n4146 37.5297
R9930 GNDA.n4149 GNDA.n4148 37.5297
R9931 GNDA.n4151 GNDA.n4150 37.5297
R9932 GNDA.n4153 GNDA.n4152 37.5297
R9933 GNDA.n4155 GNDA.n4154 37.5297
R9934 GNDA.n4157 GNDA.n4156 37.5297
R9935 GNDA.n4159 GNDA.n4158 37.5297
R9936 GNDA.n4161 GNDA.n4160 37.5297
R9937 GNDA.n4123 GNDA.n4122 37.5297
R9938 GNDA.n6778 GNDA.n99 36.7932
R9939 GNDA.n6778 GNDA.n6777 36.7932
R9940 GNDA.n6777 GNDA.n6776 36.7932
R9941 GNDA.n6776 GNDA.n293 36.7932
R9942 GNDA.n6770 GNDA.n293 36.7932
R9943 GNDA.n6769 GNDA.n6768 36.7932
R9944 GNDA.n6768 GNDA.n297 36.7932
R9945 GNDA.n6762 GNDA.n297 36.7932
R9946 GNDA.n6762 GNDA.n6761 36.7932
R9947 GNDA.n6761 GNDA.n6760 36.7932
R9948 GNDA.n6754 GNDA.n6753 36.7932
R9949 GNDA.n6753 GNDA.n6752 36.7932
R9950 GNDA.n6752 GNDA.n352 36.7932
R9951 GNDA.n6746 GNDA.n352 36.7932
R9952 GNDA.n6746 GNDA.n6745 36.7932
R9953 GNDA.n6736 GNDA.n357 36.7932
R9954 GNDA.n6736 GNDA.n6735 36.7932
R9955 GNDA.n6735 GNDA.n6734 36.7932
R9956 GNDA.n6734 GNDA.n6624 36.7932
R9957 GNDA.n6728 GNDA.n6624 36.7932
R9958 GNDA.n6726 GNDA.n6629 36.7932
R9959 GNDA.n6720 GNDA.n6629 36.7932
R9960 GNDA.n6720 GNDA.n6719 36.7932
R9961 GNDA.n6719 GNDA.n6718 36.7932
R9962 GNDA.n6718 GNDA.n6678 36.7932
R9963 GNDA.n6712 GNDA.n6711 36.7932
R9964 GNDA.n6711 GNDA.n6710 36.7932
R9965 GNDA.n6710 GNDA.n6682 36.7932
R9966 GNDA.n6704 GNDA.n6682 36.7932
R9967 GNDA.n6704 GNDA.n6703 36.7932
R9968 GNDA.n4091 GNDA.n4087 36.6977
R9969 GNDA.n4799 GNDA.n4798 36.6977
R9970 GNDA.n6247 GNDA.t165 36.5472
R9971 GNDA.t40 GNDA.t176 35.9923
R9972 GNDA.t119 GNDA.t40 35.9923
R9973 GNDA.t102 GNDA.t52 35.9923
R9974 GNDA.t52 GNDA.t846 35.9923
R9975 GNDA.t111 GNDA.n6121 35.4397
R9976 GNDA.t124 GNDA.t27 34.8629
R9977 GNDA.t74 GNDA.t19 34.8629
R9978 GNDA.n599 GNDA.n560 33.2248
R9979 GNDA.n6229 GNDA.n562 33.2248
R9980 GNDA.t743 GNDA.n26 32.9056
R9981 GNDA.t743 GNDA.n108 32.9056
R9982 GNDA.n6204 GNDA.t879 32.1173
R9983 GNDA.n4794 GNDA.n4793 31.5738
R9984 GNDA.t863 GNDA.t30 31.1932
R9985 GNDA.n4138 GNDA.t122 31.1932
R9986 GNDA.n4785 GNDA.t150 31.1932
R9987 GNDA.n1593 GNDA.t851 31.1932
R9988 GNDA.t47 GNDA.t875 31.1932
R9989 GNDA.n6092 GNDA.t839 31.1255
R9990 GNDA.n4797 GNDA.t801 31.1255
R9991 GNDA.n4092 GNDA.t747 31.1255
R9992 GNDA.n4097 GNDA.t820 31.1255
R9993 GNDA.n6107 GNDA.t172 31.0098
R9994 GNDA.t174 GNDA.n570 31.0098
R9995 GNDA.n6245 GNDA.n555 29.9023
R9996 GNDA.n4112 GNDA.n4111 29.8672
R9997 GNDA.n4089 GNDA.n4088 29.8672
R9998 GNDA.n4109 GNDA.n4108 29.8672
R9999 GNDA.n4099 GNDA.n4098 29.3583
R10000 GNDA.n6094 GNDA.n6093 29.3583
R10001 GNDA.t743 GNDA.n103 29.1014
R10002 GNDA.t109 GNDA.t25 27.6874
R10003 GNDA.t62 GNDA.t168 27.6874
R10004 GNDA.n1291 GNDA.n1290 27.5561
R10005 GNDA.n6167 GNDA.n609 27.5561
R10006 GNDA.n7086 GNDA.n7083 27.5561
R10007 GNDA.n6871 GNDA.n6868 27.5561
R10008 GNDA.n765 GNDA.n762 27.5561
R10009 GNDA.n7011 GNDA.n7010 27.5561
R10010 GNDA.n7290 GNDA.n7289 27.5561
R10011 GNDA.n1021 GNDA.n1020 27.5561
R10012 GNDA.n7209 GNDA.n7206 27.5561
R10013 GNDA.t762 GNDA.t852 27.5234
R10014 GNDA.t823 GNDA.t126 27.5234
R10015 GNDA.n1274 GNDA.n1273 26.6672
R10016 GNDA.n6145 GNDA.n613 26.6672
R10017 GNDA.n7067 GNDA.n7066 26.6672
R10018 GNDA.n6852 GNDA.n6851 26.6672
R10019 GNDA.n746 GNDA.n745 26.6672
R10020 GNDA.n6993 GNDA.n6992 26.6672
R10021 GNDA.n7272 GNDA.n7271 26.6672
R10022 GNDA.n1004 GNDA.n1003 26.6672
R10023 GNDA.n7190 GNDA.n7189 26.6672
R10024 GNDA.n1343 GNDA.n1342 26.5799
R10025 GNDA.t181 GNDA.t69 26.1768
R10026 GNDA.t69 GNDA.t162 26.1768
R10027 GNDA.t162 GNDA.t809 26.1768
R10028 GNDA.n975 GNDA.n962 25.4724
R10029 GNDA.n959 GNDA.n958 25.3679
R10030 GNDA.n540 GNDA.t161 24.0005
R10031 GNDA.n540 GNDA.t171 24.0005
R10032 GNDA.n539 GNDA.t169 24.0005
R10033 GNDA.n539 GNDA.t68 24.0005
R10034 GNDA.n538 GNDA.t175 24.0005
R10035 GNDA.n538 GNDA.t116 24.0005
R10036 GNDA.n535 GNDA.t882 24.0005
R10037 GNDA.n535 GNDA.t112 24.0005
R10038 GNDA.n534 GNDA.t173 24.0005
R10039 GNDA.n534 GNDA.t114 24.0005
R10040 GNDA.n531 GNDA.t118 24.0005
R10041 GNDA.n531 GNDA.t880 24.0005
R10042 GNDA.n530 GNDA.t178 24.0005
R10043 GNDA.n530 GNDA.t110 24.0005
R10044 GNDA.n529 GNDA.t146 24.0005
R10045 GNDA.n529 GNDA.t180 24.0005
R10046 GNDA.n526 GNDA.t163 24.0005
R10047 GNDA.n526 GNDA.t810 24.0005
R10048 GNDA.n525 GNDA.t182 24.0005
R10049 GNDA.n525 GNDA.t70 24.0005
R10050 GNDA.t11 GNDA.t147 23.995
R10051 GNDA.t166 GNDA.t867 23.995
R10052 GNDA.t803 GNDA.t819 23.8537
R10053 GNDA.t26 GNDA.t103 23.8537
R10054 GNDA.t856 GNDA.t20 23.8537
R10055 GNDA.t127 GNDA.t849 23.8537
R10056 GNDA.t806 GNDA.t838 23.8537
R10057 GNDA.n6702 GNDA.n6686 23.5958
R10058 GNDA.n6696 GNDA.n6686 23.5958
R10059 GNDA.n6696 GNDA.n6695 23.5958
R10060 GNDA.n6695 GNDA.n6694 23.5958
R10061 GNDA.n6694 GNDA.n111 23.5958
R10062 GNDA.n7144 GNDA.n7143 23.5958
R10063 GNDA.n7144 GNDA.n90 23.5958
R10064 GNDA.n7151 GNDA.n90 23.5958
R10065 GNDA.n7152 GNDA.n7151 23.5958
R10066 GNDA.n7153 GNDA.n7152 23.5958
R10067 GNDA.n7153 GNDA.n88 23.5958
R10068 GNDA.t65 GNDA.n88 23.5958
R10069 GNDA.n843 GNDA.n842 23.5958
R10070 GNDA.n842 GNDA.n841 23.5958
R10071 GNDA.n841 GNDA.n696 23.5958
R10072 GNDA.n835 GNDA.n696 23.5958
R10073 GNDA.n835 GNDA.n110 23.5958
R10074 GNDA.n703 GNDA.n109 23.5958
R10075 GNDA.n828 GNDA.n703 23.5958
R10076 GNDA.n828 GNDA.n827 23.5958
R10077 GNDA.n827 GNDA.n826 23.5958
R10078 GNDA.n826 GNDA.n704 23.5958
R10079 GNDA.n704 GNDA.n103 23.5958
R10080 GNDA.n646 GNDA.n102 23.5958
R10081 GNDA.n1225 GNDA.n646 23.5958
R10082 GNDA.n1226 GNDA.n1225 23.5958
R10083 GNDA.n1227 GNDA.n1226 23.5958
R10084 GNDA.n1227 GNDA.n552 23.5958
R10085 GNDA.n641 GNDA.n553 23.5958
R10086 GNDA.n1235 GNDA.n641 23.5958
R10087 GNDA.n1236 GNDA.n1235 23.5958
R10088 GNDA.n1336 GNDA.n1236 23.5958
R10089 GNDA.n1336 GNDA.n1335 23.5958
R10090 GNDA.n1335 GNDA.n1334 23.5958
R10091 GNDA.t743 GNDA.n106 22.15
R10092 GNDA.t835 GNDA.t32 22.0188
R10093 GNDA.t148 GNDA.t158 22.0188
R10094 GNDA.t858 GNDA.t92 22.0188
R10095 GNDA.t38 GNDA.t870 22.0188
R10096 GNDA.t6 GNDA.t137 22.0188
R10097 GNDA.t79 GNDA.t10 22.0188
R10098 GNDA.t154 GNDA.t784 22.0188
R10099 GNDA.t791 GNDA.t56 22.0188
R10100 GNDA.t89 GNDA.t152 22.0188
R10101 GNDA.t16 GNDA.t43 22.0188
R10102 GNDA.t167 GNDA.t77 22.0188
R10103 GNDA.t81 GNDA.t8 22.0188
R10104 GNDA.t96 GNDA.t101 22.0188
R10105 GNDA.t861 GNDA.t66 22.0188
R10106 GNDA.t766 GNDA.t164 22.0188
R10107 GNDA.n6621 GNDA.n6620 21.0192
R10108 GNDA.n6263 GNDA.n6262 20.8233
R10109 GNDA.n563 GNDA.n537 20.8233
R10110 GNDA.n561 GNDA.n536 20.8233
R10111 GNDA.n598 GNDA.n533 20.8233
R10112 GNDA.n582 GNDA.n532 20.8233
R10113 GNDA.n1050 GNDA.n528 20.8233
R10114 GNDA.n925 GNDA.n527 20.8233
R10115 GNDA.n629 GNDA.n524 20.8233
R10116 GNDA.n4107 GNDA.n4106 20.5612
R10117 GNDA.n1347 GNDA.n1346 20.5612
R10118 GNDA.n630 GNDA.t24 20.2276
R10119 GNDA.t98 GNDA.n4130 20.184
R10120 GNDA.n4130 GNDA.t36 20.184
R10121 GNDA.n1818 GNDA.t53 19.7005
R10122 GNDA.n1818 GNDA.t445 19.7005
R10123 GNDA.n1820 GNDA.t64 19.7005
R10124 GNDA.n1820 GNDA.t159 19.7005
R10125 GNDA.n1822 GNDA.t874 19.7005
R10126 GNDA.n1822 GNDA.t0 19.7005
R10127 GNDA.n1824 GNDA.t87 19.7005
R10128 GNDA.n1824 GNDA.t130 19.7005
R10129 GNDA.n1826 GNDA.t123 19.7005
R10130 GNDA.n1826 GNDA.t120 19.7005
R10131 GNDA.n1828 GNDA.t737 19.7005
R10132 GNDA.n1828 GNDA.t855 19.7005
R10133 GNDA.n1359 GNDA.t49 19.7005
R10134 GNDA.n1359 GNDA.t738 19.7005
R10135 GNDA.n1357 GNDA.t128 19.7005
R10136 GNDA.n1357 GNDA.t132 19.7005
R10137 GNDA.n1355 GNDA.t48 19.7005
R10138 GNDA.n1355 GNDA.t133 19.7005
R10139 GNDA.n1353 GNDA.t12 19.7005
R10140 GNDA.n1353 GNDA.t135 19.7005
R10141 GNDA.n1351 GNDA.t18 19.7005
R10142 GNDA.n1351 GNDA.t142 19.7005
R10143 GNDA.n1350 GNDA.t464 19.7005
R10144 GNDA.n1350 GNDA.t138 19.7005
R10145 GNDA.n6770 GNDA.t743 19.2145
R10146 GNDA.n6745 GNDA.t743 19.2145
R10147 GNDA.t743 GNDA.n6678 19.2145
R10148 GNDA.n6741 GNDA.n6740 18.5605
R10149 GNDA.t122 GNDA.t835 18.3491
R10150 GNDA.t32 GNDA.t148 18.3491
R10151 GNDA.t158 GNDA.t858 18.3491
R10152 GNDA.t92 GNDA.t38 18.3491
R10153 GNDA.t870 GNDA.t6 18.3491
R10154 GNDA.t137 GNDA.t79 18.3491
R10155 GNDA.t10 GNDA.t154 18.3491
R10156 GNDA.t784 GNDA.t856 18.3491
R10157 GNDA.t66 GNDA.t96 18.3491
R10158 GNDA.t164 GNDA.t861 18.3491
R10159 GNDA.t851 GNDA.t766 18.3491
R10160 GNDA.n4114 GNDA.n4112 18.0922
R10161 GNDA.n1220 GNDA.n648 17.5843
R10162 GNDA.n846 GNDA.n694 17.5843
R10163 GNDA.n6700 GNDA.n6684 17.5843
R10164 GNDA.t743 GNDA.n6769 17.5792
R10165 GNDA.t743 GNDA.n357 17.5792
R10166 GNDA.n6712 GNDA.t743 17.5792
R10167 GNDA.n263 GNDA.n260 16.9379
R10168 GNDA.n6919 GNDA.n6781 16.9379
R10169 GNDA.n1082 GNDA.n1078 16.9379
R10170 GNDA.n7138 GNDA.n134 16.7709
R10171 GNDA.n1139 GNDA.n163 16.7709
R10172 GNDA.n693 GNDA.n84 16.7709
R10173 GNDA.n905 GNDA.n904 16.7709
R10174 GNDA.t843 GNDA.t872 16.6582
R10175 GNDA.t743 GNDA.t145 16.6126
R10176 GNDA.t743 GNDA.t170 16.6126
R10177 GNDA.t864 GNDA.t803 16.5143
R10178 GNDA.t103 GNDA.t129 16.5143
R10179 GNDA.t8 GNDA.n4784 16.5143
R10180 GNDA.t849 GNDA.t134 16.5143
R10181 GNDA.t13 GNDA.t806 16.5143
R10182 GNDA.n1291 GNDA.n1246 16.0005
R10183 GNDA.n1297 GNDA.n1246 16.0005
R10184 GNDA.n1298 GNDA.n1297 16.0005
R10185 GNDA.n1299 GNDA.n1298 16.0005
R10186 GNDA.n1299 GNDA.n1244 16.0005
R10187 GNDA.n1305 GNDA.n1244 16.0005
R10188 GNDA.n1306 GNDA.n1305 16.0005
R10189 GNDA.n1309 GNDA.n1306 16.0005
R10190 GNDA.n1290 GNDA.n1289 16.0005
R10191 GNDA.n1289 GNDA.n1248 16.0005
R10192 GNDA.n1283 GNDA.n1248 16.0005
R10193 GNDA.n1283 GNDA.n1282 16.0005
R10194 GNDA.n1282 GNDA.n1281 16.0005
R10195 GNDA.n1281 GNDA.n1250 16.0005
R10196 GNDA.n1275 GNDA.n1250 16.0005
R10197 GNDA.n1275 GNDA.n1274 16.0005
R10198 GNDA.n1273 GNDA.n1252 16.0005
R10199 GNDA.n1267 GNDA.n1252 16.0005
R10200 GNDA.n1267 GNDA.n1266 16.0005
R10201 GNDA.n1266 GNDA.n1265 16.0005
R10202 GNDA.n1265 GNDA.n1254 16.0005
R10203 GNDA.n1260 GNDA.n1254 16.0005
R10204 GNDA.n1260 GNDA.n1259 16.0005
R10205 GNDA.n1259 GNDA.n1258 16.0005
R10206 GNDA.n6168 GNDA.n6167 16.0005
R10207 GNDA.n6169 GNDA.n6168 16.0005
R10208 GNDA.n6169 GNDA.n607 16.0005
R10209 GNDA.n6175 GNDA.n607 16.0005
R10210 GNDA.n6176 GNDA.n6175 16.0005
R10211 GNDA.n6177 GNDA.n6176 16.0005
R10212 GNDA.n6177 GNDA.n605 16.0005
R10213 GNDA.n605 GNDA.n595 16.0005
R10214 GNDA.n6161 GNDA.n609 16.0005
R10215 GNDA.n6161 GNDA.n6160 16.0005
R10216 GNDA.n6160 GNDA.n6159 16.0005
R10217 GNDA.n6159 GNDA.n611 16.0005
R10218 GNDA.n6153 GNDA.n611 16.0005
R10219 GNDA.n6153 GNDA.n6152 16.0005
R10220 GNDA.n6152 GNDA.n6151 16.0005
R10221 GNDA.n6151 GNDA.n613 16.0005
R10222 GNDA.n6145 GNDA.n6144 16.0005
R10223 GNDA.n6144 GNDA.n6143 16.0005
R10224 GNDA.n6143 GNDA.n615 16.0005
R10225 GNDA.n6138 GNDA.n615 16.0005
R10226 GNDA.n6138 GNDA.n6137 16.0005
R10227 GNDA.n6137 GNDA.n6136 16.0005
R10228 GNDA.n6136 GNDA.n618 16.0005
R10229 GNDA.n6131 GNDA.n618 16.0005
R10230 GNDA.n7087 GNDA.n7086 16.0005
R10231 GNDA.n7090 GNDA.n7087 16.0005
R10232 GNDA.n7091 GNDA.n7090 16.0005
R10233 GNDA.n7094 GNDA.n7091 16.0005
R10234 GNDA.n7095 GNDA.n7094 16.0005
R10235 GNDA.n7098 GNDA.n7095 16.0005
R10236 GNDA.n7099 GNDA.n7098 16.0005
R10237 GNDA.n7099 GNDA.n165 16.0005
R10238 GNDA.n7083 GNDA.n7082 16.0005
R10239 GNDA.n7082 GNDA.n7079 16.0005
R10240 GNDA.n7079 GNDA.n7078 16.0005
R10241 GNDA.n7078 GNDA.n7075 16.0005
R10242 GNDA.n7075 GNDA.n7074 16.0005
R10243 GNDA.n7074 GNDA.n7071 16.0005
R10244 GNDA.n7071 GNDA.n7070 16.0005
R10245 GNDA.n7070 GNDA.n7067 16.0005
R10246 GNDA.n7066 GNDA.n7063 16.0005
R10247 GNDA.n7063 GNDA.n7062 16.0005
R10248 GNDA.n7062 GNDA.n7059 16.0005
R10249 GNDA.n7059 GNDA.n7058 16.0005
R10250 GNDA.n7058 GNDA.n7055 16.0005
R10251 GNDA.n7055 GNDA.n7054 16.0005
R10252 GNDA.n7054 GNDA.n7051 16.0005
R10253 GNDA.n7051 GNDA.n7050 16.0005
R10254 GNDA.n6872 GNDA.n6871 16.0005
R10255 GNDA.n6875 GNDA.n6872 16.0005
R10256 GNDA.n6876 GNDA.n6875 16.0005
R10257 GNDA.n6879 GNDA.n6876 16.0005
R10258 GNDA.n6880 GNDA.n6879 16.0005
R10259 GNDA.n6883 GNDA.n6880 16.0005
R10260 GNDA.n6884 GNDA.n6883 16.0005
R10261 GNDA.n6884 GNDA.n6782 16.0005
R10262 GNDA.n6868 GNDA.n6867 16.0005
R10263 GNDA.n6867 GNDA.n6864 16.0005
R10264 GNDA.n6864 GNDA.n6863 16.0005
R10265 GNDA.n6863 GNDA.n6860 16.0005
R10266 GNDA.n6860 GNDA.n6859 16.0005
R10267 GNDA.n6859 GNDA.n6856 16.0005
R10268 GNDA.n6856 GNDA.n6855 16.0005
R10269 GNDA.n6855 GNDA.n6852 16.0005
R10270 GNDA.n6851 GNDA.n6848 16.0005
R10271 GNDA.n6848 GNDA.n6847 16.0005
R10272 GNDA.n6847 GNDA.n6844 16.0005
R10273 GNDA.n6844 GNDA.n6843 16.0005
R10274 GNDA.n6843 GNDA.n6840 16.0005
R10275 GNDA.n6840 GNDA.n6839 16.0005
R10276 GNDA.n6839 GNDA.n6836 16.0005
R10277 GNDA.n6836 GNDA.n6835 16.0005
R10278 GNDA.n766 GNDA.n765 16.0005
R10279 GNDA.n769 GNDA.n766 16.0005
R10280 GNDA.n770 GNDA.n769 16.0005
R10281 GNDA.n773 GNDA.n770 16.0005
R10282 GNDA.n774 GNDA.n773 16.0005
R10283 GNDA.n777 GNDA.n774 16.0005
R10284 GNDA.n779 GNDA.n777 16.0005
R10285 GNDA.n780 GNDA.n779 16.0005
R10286 GNDA.n762 GNDA.n761 16.0005
R10287 GNDA.n761 GNDA.n758 16.0005
R10288 GNDA.n758 GNDA.n757 16.0005
R10289 GNDA.n757 GNDA.n754 16.0005
R10290 GNDA.n754 GNDA.n753 16.0005
R10291 GNDA.n753 GNDA.n750 16.0005
R10292 GNDA.n750 GNDA.n749 16.0005
R10293 GNDA.n749 GNDA.n746 16.0005
R10294 GNDA.n745 GNDA.n742 16.0005
R10295 GNDA.n742 GNDA.n741 16.0005
R10296 GNDA.n741 GNDA.n738 16.0005
R10297 GNDA.n738 GNDA.n737 16.0005
R10298 GNDA.n737 GNDA.n734 16.0005
R10299 GNDA.n734 GNDA.n733 16.0005
R10300 GNDA.n733 GNDA.n730 16.0005
R10301 GNDA.n730 GNDA.n706 16.0005
R10302 GNDA.n7024 GNDA.n7011 16.0005
R10303 GNDA.n7024 GNDA.n7023 16.0005
R10304 GNDA.n7023 GNDA.n7022 16.0005
R10305 GNDA.n7022 GNDA.n7019 16.0005
R10306 GNDA.n7019 GNDA.n7018 16.0005
R10307 GNDA.n7018 GNDA.n7015 16.0005
R10308 GNDA.n7015 GNDA.n7014 16.0005
R10309 GNDA.n7014 GNDA.n6926 16.0005
R10310 GNDA.n7010 GNDA.n7008 16.0005
R10311 GNDA.n7008 GNDA.n7005 16.0005
R10312 GNDA.n7005 GNDA.n7004 16.0005
R10313 GNDA.n7004 GNDA.n7001 16.0005
R10314 GNDA.n7001 GNDA.n7000 16.0005
R10315 GNDA.n7000 GNDA.n6997 16.0005
R10316 GNDA.n6997 GNDA.n6996 16.0005
R10317 GNDA.n6996 GNDA.n6993 16.0005
R10318 GNDA.n6992 GNDA.n6989 16.0005
R10319 GNDA.n6989 GNDA.n6988 16.0005
R10320 GNDA.n6988 GNDA.n6985 16.0005
R10321 GNDA.n6985 GNDA.n6984 16.0005
R10322 GNDA.n6984 GNDA.n6981 16.0005
R10323 GNDA.n6981 GNDA.n6980 16.0005
R10324 GNDA.n6980 GNDA.n6977 16.0005
R10325 GNDA.n6977 GNDA.n6976 16.0005
R10326 GNDA.n6742 GNDA.n6621 16.0005
R10327 GNDA.n6742 GNDA.n6741 16.0005
R10328 GNDA.n7303 GNDA.n7290 16.0005
R10329 GNDA.n7303 GNDA.n7302 16.0005
R10330 GNDA.n7302 GNDA.n7301 16.0005
R10331 GNDA.n7301 GNDA.n7298 16.0005
R10332 GNDA.n7298 GNDA.n7297 16.0005
R10333 GNDA.n7297 GNDA.n7294 16.0005
R10334 GNDA.n7294 GNDA.n7293 16.0005
R10335 GNDA.n7293 GNDA.n57 16.0005
R10336 GNDA.n7289 GNDA.n7287 16.0005
R10337 GNDA.n7287 GNDA.n7284 16.0005
R10338 GNDA.n7284 GNDA.n7283 16.0005
R10339 GNDA.n7283 GNDA.n7280 16.0005
R10340 GNDA.n7280 GNDA.n7279 16.0005
R10341 GNDA.n7279 GNDA.n7276 16.0005
R10342 GNDA.n7276 GNDA.n7275 16.0005
R10343 GNDA.n7275 GNDA.n7272 16.0005
R10344 GNDA.n7271 GNDA.n7268 16.0005
R10345 GNDA.n7268 GNDA.n7267 16.0005
R10346 GNDA.n7267 GNDA.n7264 16.0005
R10347 GNDA.n7264 GNDA.n7263 16.0005
R10348 GNDA.n7263 GNDA.n7260 16.0005
R10349 GNDA.n7260 GNDA.n7259 16.0005
R10350 GNDA.n7259 GNDA.n7256 16.0005
R10351 GNDA.n7256 GNDA.n7255 16.0005
R10352 GNDA.n1021 GNDA.n935 16.0005
R10353 GNDA.n1027 GNDA.n935 16.0005
R10354 GNDA.n1028 GNDA.n1027 16.0005
R10355 GNDA.n1029 GNDA.n1028 16.0005
R10356 GNDA.n1029 GNDA.n933 16.0005
R10357 GNDA.n1035 GNDA.n933 16.0005
R10358 GNDA.n1036 GNDA.n1035 16.0005
R10359 GNDA.n1037 GNDA.n1036 16.0005
R10360 GNDA.n1020 GNDA.n1019 16.0005
R10361 GNDA.n1019 GNDA.n937 16.0005
R10362 GNDA.n1013 GNDA.n937 16.0005
R10363 GNDA.n1013 GNDA.n1012 16.0005
R10364 GNDA.n1012 GNDA.n1011 16.0005
R10365 GNDA.n1011 GNDA.n939 16.0005
R10366 GNDA.n1005 GNDA.n939 16.0005
R10367 GNDA.n1005 GNDA.n1004 16.0005
R10368 GNDA.n1003 GNDA.n941 16.0005
R10369 GNDA.n997 GNDA.n941 16.0005
R10370 GNDA.n997 GNDA.n996 16.0005
R10371 GNDA.n996 GNDA.n995 16.0005
R10372 GNDA.n995 GNDA.n943 16.0005
R10373 GNDA.n990 GNDA.n943 16.0005
R10374 GNDA.n990 GNDA.n989 16.0005
R10375 GNDA.n989 GNDA.n594 16.0005
R10376 GNDA.n7210 GNDA.n7209 16.0005
R10377 GNDA.n7213 GNDA.n7210 16.0005
R10378 GNDA.n7214 GNDA.n7213 16.0005
R10379 GNDA.n7217 GNDA.n7214 16.0005
R10380 GNDA.n7218 GNDA.n7217 16.0005
R10381 GNDA.n7221 GNDA.n7218 16.0005
R10382 GNDA.n7223 GNDA.n7221 16.0005
R10383 GNDA.n7224 GNDA.n7223 16.0005
R10384 GNDA.n7206 GNDA.n7205 16.0005
R10385 GNDA.n7205 GNDA.n7202 16.0005
R10386 GNDA.n7202 GNDA.n7201 16.0005
R10387 GNDA.n7201 GNDA.n7198 16.0005
R10388 GNDA.n7198 GNDA.n7197 16.0005
R10389 GNDA.n7197 GNDA.n7194 16.0005
R10390 GNDA.n7194 GNDA.n7193 16.0005
R10391 GNDA.n7193 GNDA.n7190 16.0005
R10392 GNDA.n7189 GNDA.n7186 16.0005
R10393 GNDA.n7186 GNDA.n7185 16.0005
R10394 GNDA.n7185 GNDA.n7182 16.0005
R10395 GNDA.n7182 GNDA.n7181 16.0005
R10396 GNDA.n7181 GNDA.n7178 16.0005
R10397 GNDA.n7178 GNDA.n7177 16.0005
R10398 GNDA.n7177 GNDA.n7174 16.0005
R10399 GNDA.n7174 GNDA.n7173 16.0005
R10400 GNDA.t743 GNDA.n111 15.9929
R10401 GNDA.t743 GNDA.n110 15.9929
R10402 GNDA.t743 GNDA.n552 15.9929
R10403 GNDA.n1421 GNDA.n1420 15.99
R10404 GNDA.n4805 GNDA.n4804 15.99
R10405 GNDA.n1834 GNDA.n1833 15.99
R10406 GNDA.n3466 GNDA.n3465 15.99
R10407 GNDA.t143 GNDA.t5 15.7476
R10408 GNDA.t5 GNDA.t60 15.7476
R10409 GNDA.t743 GNDA.n105 14.8877
R10410 GNDA.n6089 GNDA.n1360 14.813
R10411 GNDA.n1830 GNDA.n1829 14.813
R10412 GNDA.n6619 GNDA.n6618 14.563
R10413 GNDA.n7322 GNDA.n26 14.555
R10414 GNDA.n7043 GNDA.n108 14.555
R10415 GNDA.n4793 GNDA.n4792 14.3838
R10416 GNDA.n4088 GNDA.n1831 14.3838
R10417 GNDA.n1343 GNDA.n634 14.1577
R10418 GNDA.n4110 GNDA.n4109 14.0922
R10419 GNDA.n6231 GNDA.n6230 13.313
R10420 GNDA.n978 GNDA.t177 13.2902
R10421 GNDA.n6104 GNDA.t881 13.2902
R10422 GNDA.n1321 GNDA.t160 13.2902
R10423 GNDA.n1333 GNDA.t62 13.109
R10424 GNDA.t62 GNDA.n634 13.109
R10425 GNDA.t121 GNDA.t762 12.8445
R10426 GNDA.n4087 GNDA.t746 12.8445
R10427 GNDA.n4799 GNDA.t800 12.8445
R10428 GNDA.t848 GNDA.t823 12.8445
R10429 GNDA.n1365 GNDA.t807 12.6791
R10430 GNDA.n4800 GNDA.t824 12.6791
R10431 GNDA.n4086 GNDA.t763 12.6791
R10432 GNDA.n3461 GNDA.t804 12.6791
R10433 GNDA.t147 GNDA.t28 11.9978
R10434 GNDA.t176 GNDA.t11 11.9978
R10435 GNDA.t846 GNDA.t166 11.9978
R10436 GNDA.t867 GNDA.t871 11.9978
R10437 GNDA.t24 GNDA.t843 11.8988
R10438 GNDA.n1221 GNDA.n1220 11.6369
R10439 GNDA.n1223 GNDA.n1221 11.6369
R10440 GNDA.n1223 GNDA.n1222 11.6369
R10441 GNDA.n1222 GNDA.n645 11.6369
R10442 GNDA.n645 GNDA.n643 11.6369
R10443 GNDA.n1231 GNDA.n643 11.6369
R10444 GNDA.n1232 GNDA.n1231 11.6369
R10445 GNDA.n1233 GNDA.n1232 11.6369
R10446 GNDA.n1233 GNDA.n638 11.6369
R10447 GNDA.n1338 GNDA.n638 11.6369
R10448 GNDA.n1198 GNDA.n1197 11.6369
R10449 GNDA.n1199 GNDA.n1198 11.6369
R10450 GNDA.n1199 GNDA.n652 11.6369
R10451 GNDA.n1205 GNDA.n652 11.6369
R10452 GNDA.n1206 GNDA.n1205 11.6369
R10453 GNDA.n1207 GNDA.n1206 11.6369
R10454 GNDA.n1207 GNDA.n650 11.6369
R10455 GNDA.n1213 GNDA.n650 11.6369
R10456 GNDA.n1214 GNDA.n1213 11.6369
R10457 GNDA.n1215 GNDA.n1214 11.6369
R10458 GNDA.n1215 GNDA.n648 11.6369
R10459 GNDA.n1140 GNDA.n912 11.6369
R10460 GNDA.n1146 GNDA.n912 11.6369
R10461 GNDA.n1147 GNDA.n1146 11.6369
R10462 GNDA.n1148 GNDA.n1147 11.6369
R10463 GNDA.n1148 GNDA.n910 11.6369
R10464 GNDA.n1154 GNDA.n910 11.6369
R10465 GNDA.n1155 GNDA.n1154 11.6369
R10466 GNDA.n1156 GNDA.n1155 11.6369
R10467 GNDA.n1156 GNDA.n908 11.6369
R10468 GNDA.n1161 GNDA.n908 11.6369
R10469 GNDA.n1162 GNDA.n1161 11.6369
R10470 GNDA.n698 GNDA.n694 11.6369
R10471 GNDA.n839 GNDA.n698 11.6369
R10472 GNDA.n839 GNDA.n838 11.6369
R10473 GNDA.n838 GNDA.n837 11.6369
R10474 GNDA.n837 GNDA.n699 11.6369
R10475 GNDA.n832 GNDA.n699 11.6369
R10476 GNDA.n832 GNDA.n831 11.6369
R10477 GNDA.n831 GNDA.n830 11.6369
R10478 GNDA.n830 GNDA.n701 11.6369
R10479 GNDA.n824 GNDA.n701 11.6369
R10480 GNDA.n867 GNDA.n866 11.6369
R10481 GNDA.n866 GNDA.n863 11.6369
R10482 GNDA.n863 GNDA.n862 11.6369
R10483 GNDA.n862 GNDA.n859 11.6369
R10484 GNDA.n859 GNDA.n858 11.6369
R10485 GNDA.n858 GNDA.n855 11.6369
R10486 GNDA.n855 GNDA.n854 11.6369
R10487 GNDA.n854 GNDA.n851 11.6369
R10488 GNDA.n851 GNDA.n850 11.6369
R10489 GNDA.n850 GNDA.n847 11.6369
R10490 GNDA.n847 GNDA.n846 11.6369
R10491 GNDA.n670 GNDA.n133 11.6369
R10492 GNDA.n673 GNDA.n670 11.6369
R10493 GNDA.n674 GNDA.n673 11.6369
R10494 GNDA.n677 GNDA.n674 11.6369
R10495 GNDA.n678 GNDA.n677 11.6369
R10496 GNDA.n681 GNDA.n678 11.6369
R10497 GNDA.n682 GNDA.n681 11.6369
R10498 GNDA.n685 GNDA.n682 11.6369
R10499 GNDA.n686 GNDA.n685 11.6369
R10500 GNDA.n689 GNDA.n686 11.6369
R10501 GNDA.n692 GNDA.n689 11.6369
R10502 GNDA.n264 GNDA.n263 11.6369
R10503 GNDA.n267 GNDA.n264 11.6369
R10504 GNDA.n268 GNDA.n267 11.6369
R10505 GNDA.n271 GNDA.n268 11.6369
R10506 GNDA.n272 GNDA.n271 11.6369
R10507 GNDA.n275 GNDA.n272 11.6369
R10508 GNDA.n276 GNDA.n275 11.6369
R10509 GNDA.n278 GNDA.n276 11.6369
R10510 GNDA.n278 GNDA.n277 11.6369
R10511 GNDA.n277 GNDA.n229 11.6369
R10512 GNDA.n260 GNDA.n259 11.6369
R10513 GNDA.n259 GNDA.n256 11.6369
R10514 GNDA.n256 GNDA.n255 11.6369
R10515 GNDA.n255 GNDA.n252 11.6369
R10516 GNDA.n252 GNDA.n251 11.6369
R10517 GNDA.n251 GNDA.n248 11.6369
R10518 GNDA.n248 GNDA.n247 11.6369
R10519 GNDA.n247 GNDA.n244 11.6369
R10520 GNDA.n244 GNDA.n243 11.6369
R10521 GNDA.n243 GNDA.n132 11.6369
R10522 GNDA.n7139 GNDA.n132 11.6369
R10523 GNDA.n6919 GNDA.n6918 11.6369
R10524 GNDA.n6918 GNDA.n6917 11.6369
R10525 GNDA.n6917 GNDA.n6916 11.6369
R10526 GNDA.n6916 GNDA.n6914 11.6369
R10527 GNDA.n6914 GNDA.n6911 11.6369
R10528 GNDA.n6911 GNDA.n6910 11.6369
R10529 GNDA.n6910 GNDA.n6907 11.6369
R10530 GNDA.n6907 GNDA.n6906 11.6369
R10531 GNDA.n6906 GNDA.n6903 11.6369
R10532 GNDA.n6903 GNDA.n6902 11.6369
R10533 GNDA.n6781 GNDA.n6780 11.6369
R10534 GNDA.n6780 GNDA.n291 11.6369
R10535 GNDA.n6774 GNDA.n291 11.6369
R10536 GNDA.n6774 GNDA.n6773 11.6369
R10537 GNDA.n6773 GNDA.n6772 11.6369
R10538 GNDA.n6772 GNDA.n295 11.6369
R10539 GNDA.n6766 GNDA.n295 11.6369
R10540 GNDA.n6766 GNDA.n6765 11.6369
R10541 GNDA.n6765 GNDA.n6764 11.6369
R10542 GNDA.n6764 GNDA.n299 11.6369
R10543 GNDA.n6758 GNDA.n299 11.6369
R10544 GNDA.n1078 GNDA.n1077 11.6369
R10545 GNDA.n1077 GNDA.n1074 11.6369
R10546 GNDA.n1074 GNDA.n1073 11.6369
R10547 GNDA.n1073 GNDA.n1070 11.6369
R10548 GNDA.n1070 GNDA.n1069 11.6369
R10549 GNDA.n1069 GNDA.n1066 11.6369
R10550 GNDA.n1066 GNDA.n1065 11.6369
R10551 GNDA.n1065 GNDA.n1062 11.6369
R10552 GNDA.n1062 GNDA.n1061 11.6369
R10553 GNDA.n1061 GNDA.n1058 11.6369
R10554 GNDA.n1083 GNDA.n1082 11.6369
R10555 GNDA.n1084 GNDA.n1083 11.6369
R10556 GNDA.n1084 GNDA.n919 11.6369
R10557 GNDA.n1090 GNDA.n919 11.6369
R10558 GNDA.n1091 GNDA.n1090 11.6369
R10559 GNDA.n1092 GNDA.n1091 11.6369
R10560 GNDA.n1092 GNDA.n917 11.6369
R10561 GNDA.n1097 GNDA.n917 11.6369
R10562 GNDA.n1098 GNDA.n1097 11.6369
R10563 GNDA.n1098 GNDA.n915 11.6369
R10564 GNDA.n1138 GNDA.n915 11.6369
R10565 GNDA.n6700 GNDA.n6699 11.6369
R10566 GNDA.n6699 GNDA.n6698 11.6369
R10567 GNDA.n6698 GNDA.n6688 11.6369
R10568 GNDA.n6692 GNDA.n6688 11.6369
R10569 GNDA.n6692 GNDA.n6691 11.6369
R10570 GNDA.n6691 GNDA.n92 11.6369
R10571 GNDA.n7146 GNDA.n92 11.6369
R10572 GNDA.n7147 GNDA.n7146 11.6369
R10573 GNDA.n7149 GNDA.n7147 11.6369
R10574 GNDA.n7149 GNDA.n7148 11.6369
R10575 GNDA.n6724 GNDA.n6723 11.6369
R10576 GNDA.n6723 GNDA.n6722 11.6369
R10577 GNDA.n6722 GNDA.n6676 11.6369
R10578 GNDA.n6716 GNDA.n6676 11.6369
R10579 GNDA.n6716 GNDA.n6715 11.6369
R10580 GNDA.n6715 GNDA.n6714 11.6369
R10581 GNDA.n6714 GNDA.n6680 11.6369
R10582 GNDA.n6708 GNDA.n6680 11.6369
R10583 GNDA.n6708 GNDA.n6707 11.6369
R10584 GNDA.n6707 GNDA.n6706 11.6369
R10585 GNDA.n6706 GNDA.n6684 11.6369
R10586 GNDA.n6756 GNDA.n304 11.6369
R10587 GNDA.n6750 GNDA.n304 11.6369
R10588 GNDA.n6750 GNDA.n6749 11.6369
R10589 GNDA.n6749 GNDA.n6748 11.6369
R10590 GNDA.n6748 GNDA.n354 11.6369
R10591 GNDA.n6739 GNDA.n6622 11.6369
R10592 GNDA.n6626 GNDA.n6622 11.6369
R10593 GNDA.n6732 GNDA.n6626 11.6369
R10594 GNDA.n6732 GNDA.n6731 11.6369
R10595 GNDA.n6731 GNDA.n6730 11.6369
R10596 GNDA.n6282 GNDA.n6280 11.0384
R10597 GNDA.t878 GNDA.t791 11.0097
R10598 GNDA.t71 GNDA.t89 11.0097
R10599 GNDA.t84 GNDA.t16 11.0097
R10600 GNDA.t91 GNDA.t167 11.0097
R10601 GNDA.t740 GNDA.t81 11.0097
R10602 GNDA.n6264 GNDA.n6263 10.9846
R10603 GNDA.n6280 GNDA.n524 10.87
R10604 GNDA.n6277 GNDA.n527 10.87
R10605 GNDA.n6276 GNDA.n528 10.87
R10606 GNDA.n6272 GNDA.n532 10.87
R10607 GNDA.n6271 GNDA.n533 10.87
R10608 GNDA.n6268 GNDA.n536 10.87
R10609 GNDA.n6267 GNDA.n537 10.87
R10610 GNDA.n4121 GNDA.n1816 10.563
R10611 GNDA.n4140 GNDA.t862 9.6005
R10612 GNDA.n4140 GNDA.t767 9.6005
R10613 GNDA.n4142 GNDA.t9 9.6005
R10614 GNDA.n4142 GNDA.t97 9.6005
R10615 GNDA.n4144 GNDA.t44 9.6005
R10616 GNDA.n4144 GNDA.t78 9.6005
R10617 GNDA.n4146 GNDA.t57 9.6005
R10618 GNDA.n4146 GNDA.t153 9.6005
R10619 GNDA.n4148 GNDA.t55 9.6005
R10620 GNDA.n4148 GNDA.t151 9.6005
R10621 GNDA.n4150 GNDA.t37 9.6005
R10622 GNDA.n4150 GNDA.t46 9.6005
R10623 GNDA.n4152 GNDA.t860 9.6005
R10624 GNDA.n4152 GNDA.t99 9.6005
R10625 GNDA.n4154 GNDA.t857 9.6005
R10626 GNDA.n4154 GNDA.t157 9.6005
R10627 GNDA.n4156 GNDA.t80 9.6005
R10628 GNDA.n4156 GNDA.t155 9.6005
R10629 GNDA.n4158 GNDA.t39 9.6005
R10630 GNDA.n4158 GNDA.t7 9.6005
R10631 GNDA.n4160 GNDA.t149 9.6005
R10632 GNDA.n4160 GNDA.t859 9.6005
R10633 GNDA.n4122 GNDA.t869 9.6005
R10634 GNDA.n4122 GNDA.t95 9.6005
R10635 GNDA.n6239 GNDA.t447 9.6005
R10636 GNDA.n6242 GNDA.t466 9.6005
R10637 GNDA.n951 GNDA.t470 9.6005
R10638 GNDA.n957 GNDA.t729 9.6005
R10639 GNDA.t872 GNDA.t181 9.51916
R10640 GNDA.t30 GNDA.t90 9.17481
R10641 GNDA.n4138 GNDA.t76 9.17481
R10642 GNDA.n4137 GNDA.t156 9.17481
R10643 GNDA.n1593 GNDA.t144 9.17481
R10644 GNDA.t875 GNDA.t136 9.17481
R10645 GNDA.n6282 GNDA.n6281 8.938
R10646 GNDA.n976 GNDA.t179 8.8603
R10647 GNDA.n6108 GNDA.t113 8.8603
R10648 GNDA.n1320 GNDA.t67 8.8603
R10649 GNDA.n4095 GNDA.n1830 8.78175
R10650 GNDA.n6090 GNDA.n6089 8.78175
R10651 GNDA.n7229 GNDA.n26 8.60107
R10652 GNDA.n162 GNDA.n108 8.60107
R10653 GNDA.n4163 GNDA.n4162 8.3755
R10654 GNDA.t33 GNDA.n630 8.32933
R10655 GNDA.t743 GNDA.n99 8.17666
R10656 GNDA.n6089 GNDA.n6088 7.77133
R10657 GNDA.n1888 GNDA.n1830 7.77133
R10658 GNDA.n926 GNDA.n106 7.75283
R10659 GNDA.n1049 GNDA.t17 7.75283
R10660 GNDA.n977 GNDA.t25 7.75283
R10661 GNDA.n6123 GNDA.n562 7.75283
R10662 GNDA.n6261 GNDA.n541 7.75283
R10663 GNDA.n7143 GNDA.t743 7.60343
R10664 GNDA.t743 GNDA.n109 7.60343
R10665 GNDA.t743 GNDA.n553 7.60343
R10666 GNDA.n4110 GNDA.n1816 7.438
R10667 GNDA.n4098 GNDA.n1817 7.33995
R10668 GNDA.t20 GNDA.n4137 7.33995
R10669 GNDA.t54 GNDA.t832 7.33995
R10670 GNDA.t150 GNDA.t878 7.33995
R10671 GNDA.t56 GNDA.t71 7.33995
R10672 GNDA.t152 GNDA.t84 7.33995
R10673 GNDA.t43 GNDA.t91 7.33995
R10674 GNDA.t77 GNDA.t740 7.33995
R10675 GNDA.n6093 GNDA.n1348 7.33995
R10676 GNDA.n1819 GNDA.n1816 6.90675
R10677 GNDA.n1162 GNDA.n905 6.72373
R10678 GNDA.n693 GNDA.n692 6.72373
R10679 GNDA.n7139 GNDA.n7138 6.72373
R10680 GNDA.n6758 GNDA.n6757 6.72373
R10681 GNDA.n1139 GNDA.n1138 6.72373
R10682 GNDA.n6730 GNDA.n6627 6.72373
R10683 GNDA.t41 GNDA.t743 6.64535
R10684 GNDA.n6283 GNDA.n6282 6.42238
R10685 GNDA.n1197 GNDA.n905 6.20656
R10686 GNDA.n1140 GNDA.n1139 6.20656
R10687 GNDA.n867 GNDA.n693 6.20656
R10688 GNDA.n7138 GNDA.n133 6.20656
R10689 GNDA.n6724 GNDA.n6627 6.20656
R10690 GNDA.n6757 GNDA.n6756 6.20656
R10691 GNDA.n6740 GNDA.n354 6.07727
R10692 GNDA.t809 GNDA.t469 5.94966
R10693 GNDA.n959 GNDA.n559 5.81868
R10694 GNDA.n959 GNDA.n950 5.81868
R10695 GNDA.n6740 GNDA.n6739 5.5601
R10696 GNDA.t58 GNDA.t778 5.53788
R10697 GNDA.n962 GNDA.t145 5.53788
R10698 GNDA.t743 GNDA.t788 5.53788
R10699 GNDA.n6103 GNDA.t743 5.53788
R10700 GNDA.t743 GNDA.t826 5.53788
R10701 GNDA.t170 GNDA.n6245 5.53788
R10702 GNDA.t165 GNDA.t775 5.53788
R10703 GNDA.n1258 GNDA.n636 5.51161
R10704 GNDA.n6131 GNDA.n567 5.51161
R10705 GNDA.n7050 GNDA.n187 5.51161
R10706 GNDA.n6835 GNDA.n6805 5.51161
R10707 GNDA.n818 GNDA.n706 5.51161
R10708 GNDA.n6976 GNDA.n6954 5.51161
R10709 GNDA.n7255 GNDA.n7233 5.51161
R10710 GNDA.n6199 GNDA.n594 5.51161
R10711 GNDA.n7173 GNDA.n7159 5.51161
R10712 GNDA.t106 GNDA.t124 5.50509
R10713 GNDA.t847 GNDA.t74 5.50509
R10714 GNDA.n1340 GNDA.n1339 5.1717
R10715 GNDA.n823 GNDA.n819 5.1717
R10716 GNDA.n7158 GNDA.n87 5.1717
R10717 GNDA.n4791 GNDA.n4790 5.08383
R10718 GNDA.n4133 GNDA.n1589 5.08383
R10719 GNDA.n4162 GNDA.n4161 5.063
R10720 GNDA.n4124 GNDA.n4123 5.063
R10721 GNDA.n7040 GNDA.n6925 4.9157
R10722 GNDA.n6899 GNDA.n6896 4.9157
R10723 GNDA.n1057 GNDA.n1056 4.9157
R10724 GNDA.n6091 GNDA.n6090 4.85467
R10725 GNDA.n4796 GNDA.n1349 4.85467
R10726 GNDA.n4094 GNDA.n4093 4.85467
R10727 GNDA.n4096 GNDA.n4095 4.85467
R10728 GNDA.n4782 GNDA.n4781 4.83383
R10729 GNDA.n4127 GNDA.n1648 4.83383
R10730 GNDA.n6446 GNDA.t888 4.8295
R10731 GNDA.n6449 GNDA.t948 4.8295
R10732 GNDA.n6453 GNDA.t939 4.8295
R10733 GNDA.n6456 GNDA.t1000 4.8295
R10734 GNDA.n6460 GNDA.t1002 4.8295
R10735 GNDA.n6463 GNDA.t1061 4.8295
R10736 GNDA.n6467 GNDA.t1063 4.8295
R10737 GNDA.n6470 GNDA.t908 4.8295
R10738 GNDA.n6474 GNDA.t1010 4.8295
R10739 GNDA.n6477 GNDA.t1071 4.8295
R10740 GNDA.n6481 GNDA.t1073 4.8295
R10741 GNDA.n6484 GNDA.t916 4.8295
R10742 GNDA.n6488 GNDA.t917 4.8295
R10743 GNDA.n6491 GNDA.t976 4.8295
R10744 GNDA.n6495 GNDA.t1079 4.8295
R10745 GNDA.n6498 GNDA.t925 4.8295
R10746 GNDA.n6502 GNDA.t927 4.8295
R10747 GNDA.n6505 GNDA.t986 4.8295
R10748 GNDA.n6509 GNDA.t987 4.8295
R10749 GNDA.n6512 GNDA.t1048 4.8295
R10750 GNDA.n6516 GNDA.t932 4.8295
R10751 GNDA.n6519 GNDA.t993 4.8295
R10752 GNDA.n6523 GNDA.t994 4.8295
R10753 GNDA.n6526 GNDA.t1052 4.8295
R10754 GNDA.n6530 GNDA.t1053 4.8295
R10755 GNDA.n6533 GNDA.t898 4.8295
R10756 GNDA.n6537 GNDA.t900 4.8295
R10757 GNDA.n6540 GNDA.t960 4.8295
R10758 GNDA.n6544 GNDA.t1062 4.8295
R10759 GNDA.n6547 GNDA.t907 4.8295
R10760 GNDA.n6551 GNDA.t899 4.8295
R10761 GNDA.n6554 GNDA.t959 4.8295
R10762 GNDA.n6558 GNDA.t961 4.8295
R10763 GNDA.n6561 GNDA.t1022 4.8295
R10764 GNDA.n6565 GNDA.t909 4.8295
R10765 GNDA.n6568 GNDA.t966 4.8295
R10766 GNDA.n6572 GNDA.t968 4.8295
R10767 GNDA.n6575 GNDA.t1026 4.8295
R10768 GNDA.n6579 GNDA.t1028 4.8295
R10769 GNDA.n6582 GNDA.t1088 4.8295
R10770 GNDA.n6586 GNDA.t977 4.8295
R10771 GNDA.n6589 GNDA.t1036 4.8295
R10772 GNDA.n6593 GNDA.t1037 4.8295
R10773 GNDA.n6596 GNDA.t1098 4.8295
R10774 GNDA.n6600 GNDA.t883 4.8295
R10775 GNDA.n6603 GNDA.t944 4.8295
R10776 GNDA.n6607 GNDA.t1007 4.8295
R10777 GNDA.n4116 GNDA.n4115 4.79217
R10778 GNDA.n4114 GNDA.n4113 4.79217
R10779 GNDA.n4141 GNDA.n1595 4.71925
R10780 GNDA.t60 GNDA.n632 4.5934
R10781 GNDA.n4778 GNDA.n4777 4.5005
R10782 GNDA.n1597 GNDA.n1596 4.5005
R10783 GNDA.n4663 GNDA.n4662 4.5005
R10784 GNDA.n4667 GNDA.n4664 4.5005
R10785 GNDA.n4668 GNDA.n4661 4.5005
R10786 GNDA.n4672 GNDA.n4671 4.5005
R10787 GNDA.n4673 GNDA.n4660 4.5005
R10788 GNDA.n4677 GNDA.n4674 4.5005
R10789 GNDA.n4678 GNDA.n4659 4.5005
R10790 GNDA.n4682 GNDA.n4681 4.5005
R10791 GNDA.n4683 GNDA.n4658 4.5005
R10792 GNDA.n4687 GNDA.n4684 4.5005
R10793 GNDA.n4688 GNDA.n4657 4.5005
R10794 GNDA.n4692 GNDA.n4691 4.5005
R10795 GNDA.n4693 GNDA.n4656 4.5005
R10796 GNDA.n4697 GNDA.n4694 4.5005
R10797 GNDA.n4698 GNDA.n4655 4.5005
R10798 GNDA.n4702 GNDA.n4701 4.5005
R10799 GNDA.n4703 GNDA.n4654 4.5005
R10800 GNDA.n4707 GNDA.n4704 4.5005
R10801 GNDA.n4708 GNDA.n4653 4.5005
R10802 GNDA.n4712 GNDA.n4711 4.5005
R10803 GNDA.n4713 GNDA.n4652 4.5005
R10804 GNDA.n4717 GNDA.n4714 4.5005
R10805 GNDA.n4718 GNDA.n4651 4.5005
R10806 GNDA.n4722 GNDA.n4721 4.5005
R10807 GNDA.n4723 GNDA.n4650 4.5005
R10808 GNDA.n4727 GNDA.n4724 4.5005
R10809 GNDA.n4728 GNDA.n4649 4.5005
R10810 GNDA.n4732 GNDA.n4731 4.5005
R10811 GNDA.n4733 GNDA.n4648 4.5005
R10812 GNDA.n4737 GNDA.n4734 4.5005
R10813 GNDA.n4738 GNDA.n4647 4.5005
R10814 GNDA.n4742 GNDA.n4741 4.5005
R10815 GNDA.n4743 GNDA.n4646 4.5005
R10816 GNDA.n4747 GNDA.n4744 4.5005
R10817 GNDA.n4748 GNDA.n4645 4.5005
R10818 GNDA.n4752 GNDA.n4751 4.5005
R10819 GNDA.n4753 GNDA.n4644 4.5005
R10820 GNDA.n4757 GNDA.n4754 4.5005
R10821 GNDA.n4758 GNDA.n4643 4.5005
R10822 GNDA.n4762 GNDA.n4761 4.5005
R10823 GNDA.n4763 GNDA.n4642 4.5005
R10824 GNDA.n4767 GNDA.n4764 4.5005
R10825 GNDA.n4768 GNDA.n4641 4.5005
R10826 GNDA.n4772 GNDA.n4771 4.5005
R10827 GNDA.n5686 GNDA.n1361 4.5005
R10828 GNDA.n5689 GNDA.n5688 4.5005
R10829 GNDA.n5690 GNDA.n5685 4.5005
R10830 GNDA.n5694 GNDA.n5691 4.5005
R10831 GNDA.n5695 GNDA.n5684 4.5005
R10832 GNDA.n5699 GNDA.n5698 4.5005
R10833 GNDA.n5700 GNDA.n5683 4.5005
R10834 GNDA.n5704 GNDA.n5701 4.5005
R10835 GNDA.n5705 GNDA.n5682 4.5005
R10836 GNDA.n5709 GNDA.n5708 4.5005
R10837 GNDA.n5710 GNDA.n5681 4.5005
R10838 GNDA.n5714 GNDA.n5711 4.5005
R10839 GNDA.n5715 GNDA.n5680 4.5005
R10840 GNDA.n5719 GNDA.n5718 4.5005
R10841 GNDA.n5720 GNDA.n5679 4.5005
R10842 GNDA.n5724 GNDA.n5721 4.5005
R10843 GNDA.n5725 GNDA.n5678 4.5005
R10844 GNDA.n5729 GNDA.n5728 4.5005
R10845 GNDA.n5730 GNDA.n5677 4.5005
R10846 GNDA.n5734 GNDA.n5731 4.5005
R10847 GNDA.n5735 GNDA.n5676 4.5005
R10848 GNDA.n5739 GNDA.n5738 4.5005
R10849 GNDA.n5740 GNDA.n5675 4.5005
R10850 GNDA.n5744 GNDA.n5741 4.5005
R10851 GNDA.n5745 GNDA.n5674 4.5005
R10852 GNDA.n5749 GNDA.n5748 4.5005
R10853 GNDA.n5750 GNDA.n5673 4.5005
R10854 GNDA.n5754 GNDA.n5751 4.5005
R10855 GNDA.n5755 GNDA.n5672 4.5005
R10856 GNDA.n5759 GNDA.n5758 4.5005
R10857 GNDA.n5760 GNDA.n5671 4.5005
R10858 GNDA.n5764 GNDA.n5761 4.5005
R10859 GNDA.n5765 GNDA.n5670 4.5005
R10860 GNDA.n5769 GNDA.n5768 4.5005
R10861 GNDA.n5770 GNDA.n5669 4.5005
R10862 GNDA.n5774 GNDA.n5771 4.5005
R10863 GNDA.n5775 GNDA.n5668 4.5005
R10864 GNDA.n5779 GNDA.n5778 4.5005
R10865 GNDA.n5780 GNDA.n5667 4.5005
R10866 GNDA.n5784 GNDA.n5781 4.5005
R10867 GNDA.n5785 GNDA.n5666 4.5005
R10868 GNDA.n5789 GNDA.n5788 4.5005
R10869 GNDA.n5790 GNDA.n5665 4.5005
R10870 GNDA.n5794 GNDA.n5791 4.5005
R10871 GNDA.n5795 GNDA.n5664 4.5005
R10872 GNDA.n5799 GNDA.n5798 4.5005
R10873 GNDA.n6083 GNDA.n6082 4.5005
R10874 GNDA.n1369 GNDA.n1368 4.5005
R10875 GNDA.n5968 GNDA.n5967 4.5005
R10876 GNDA.n5972 GNDA.n5969 4.5005
R10877 GNDA.n5973 GNDA.n5966 4.5005
R10878 GNDA.n5977 GNDA.n5976 4.5005
R10879 GNDA.n5978 GNDA.n5965 4.5005
R10880 GNDA.n5982 GNDA.n5979 4.5005
R10881 GNDA.n5983 GNDA.n5964 4.5005
R10882 GNDA.n5987 GNDA.n5986 4.5005
R10883 GNDA.n5988 GNDA.n5963 4.5005
R10884 GNDA.n5992 GNDA.n5989 4.5005
R10885 GNDA.n5993 GNDA.n5962 4.5005
R10886 GNDA.n5997 GNDA.n5996 4.5005
R10887 GNDA.n5998 GNDA.n5961 4.5005
R10888 GNDA.n6002 GNDA.n5999 4.5005
R10889 GNDA.n6003 GNDA.n5960 4.5005
R10890 GNDA.n6007 GNDA.n6006 4.5005
R10891 GNDA.n6008 GNDA.n5959 4.5005
R10892 GNDA.n6012 GNDA.n6009 4.5005
R10893 GNDA.n6013 GNDA.n5958 4.5005
R10894 GNDA.n6017 GNDA.n6016 4.5005
R10895 GNDA.n6018 GNDA.n5957 4.5005
R10896 GNDA.n6022 GNDA.n6019 4.5005
R10897 GNDA.n6023 GNDA.n5956 4.5005
R10898 GNDA.n6027 GNDA.n6026 4.5005
R10899 GNDA.n6028 GNDA.n5955 4.5005
R10900 GNDA.n6032 GNDA.n6029 4.5005
R10901 GNDA.n6033 GNDA.n5954 4.5005
R10902 GNDA.n6037 GNDA.n6036 4.5005
R10903 GNDA.n6038 GNDA.n5953 4.5005
R10904 GNDA.n6042 GNDA.n6039 4.5005
R10905 GNDA.n6043 GNDA.n5952 4.5005
R10906 GNDA.n6047 GNDA.n6046 4.5005
R10907 GNDA.n6048 GNDA.n5951 4.5005
R10908 GNDA.n6052 GNDA.n6049 4.5005
R10909 GNDA.n6053 GNDA.n5950 4.5005
R10910 GNDA.n6057 GNDA.n6056 4.5005
R10911 GNDA.n6058 GNDA.n5949 4.5005
R10912 GNDA.n6062 GNDA.n6059 4.5005
R10913 GNDA.n6063 GNDA.n5948 4.5005
R10914 GNDA.n6067 GNDA.n6066 4.5005
R10915 GNDA.n6068 GNDA.n5947 4.5005
R10916 GNDA.n6072 GNDA.n6069 4.5005
R10917 GNDA.n6073 GNDA.n5946 4.5005
R10918 GNDA.n6077 GNDA.n6076 4.5005
R10919 GNDA.n1587 GNDA.n1586 4.5005
R10920 GNDA.n1424 GNDA.n1423 4.5005
R10921 GNDA.n1470 GNDA.n1425 4.5005
R10922 GNDA.n1471 GNDA.n1426 4.5005
R10923 GNDA.n1472 GNDA.n1427 4.5005
R10924 GNDA.n1473 GNDA.n1428 4.5005
R10925 GNDA.n1474 GNDA.n1429 4.5005
R10926 GNDA.n1475 GNDA.n1430 4.5005
R10927 GNDA.n1476 GNDA.n1431 4.5005
R10928 GNDA.n1477 GNDA.n1432 4.5005
R10929 GNDA.n1478 GNDA.n1433 4.5005
R10930 GNDA.n1479 GNDA.n1434 4.5005
R10931 GNDA.n1480 GNDA.n1435 4.5005
R10932 GNDA.n1481 GNDA.n1436 4.5005
R10933 GNDA.n1482 GNDA.n1437 4.5005
R10934 GNDA.n1483 GNDA.n1438 4.5005
R10935 GNDA.n1484 GNDA.n1439 4.5005
R10936 GNDA.n1485 GNDA.n1440 4.5005
R10937 GNDA.n1486 GNDA.n1441 4.5005
R10938 GNDA.n1487 GNDA.n1442 4.5005
R10939 GNDA.n1488 GNDA.n1443 4.5005
R10940 GNDA.n1489 GNDA.n1444 4.5005
R10941 GNDA.n1490 GNDA.n1445 4.5005
R10942 GNDA.n1491 GNDA.n1446 4.5005
R10943 GNDA.n1492 GNDA.n1447 4.5005
R10944 GNDA.n1493 GNDA.n1448 4.5005
R10945 GNDA.n1494 GNDA.n1449 4.5005
R10946 GNDA.n1495 GNDA.n1450 4.5005
R10947 GNDA.n1496 GNDA.n1451 4.5005
R10948 GNDA.n1497 GNDA.n1452 4.5005
R10949 GNDA.n1498 GNDA.n1453 4.5005
R10950 GNDA.n1499 GNDA.n1454 4.5005
R10951 GNDA.n1500 GNDA.n1455 4.5005
R10952 GNDA.n1501 GNDA.n1456 4.5005
R10953 GNDA.n1502 GNDA.n1457 4.5005
R10954 GNDA.n1503 GNDA.n1458 4.5005
R10955 GNDA.n1504 GNDA.n1459 4.5005
R10956 GNDA.n1505 GNDA.n1460 4.5005
R10957 GNDA.n1506 GNDA.n1461 4.5005
R10958 GNDA.n1507 GNDA.n1462 4.5005
R10959 GNDA.n1508 GNDA.n1463 4.5005
R10960 GNDA.n1509 GNDA.n1464 4.5005
R10961 GNDA.n1510 GNDA.n1465 4.5005
R10962 GNDA.n1511 GNDA.n1466 4.5005
R10963 GNDA.n1512 GNDA.n1467 4.5005
R10964 GNDA.n1513 GNDA.n1468 4.5005
R10965 GNDA.n3635 GNDA.n3634 4.5005
R10966 GNDA.n3638 GNDA.n3637 4.5005
R10967 GNDA.n3639 GNDA.n3633 4.5005
R10968 GNDA.n3643 GNDA.n3640 4.5005
R10969 GNDA.n3644 GNDA.n3632 4.5005
R10970 GNDA.n3648 GNDA.n3647 4.5005
R10971 GNDA.n3649 GNDA.n3631 4.5005
R10972 GNDA.n3653 GNDA.n3650 4.5005
R10973 GNDA.n3654 GNDA.n3630 4.5005
R10974 GNDA.n3658 GNDA.n3657 4.5005
R10975 GNDA.n3659 GNDA.n3629 4.5005
R10976 GNDA.n3663 GNDA.n3660 4.5005
R10977 GNDA.n3664 GNDA.n3628 4.5005
R10978 GNDA.n3668 GNDA.n3667 4.5005
R10979 GNDA.n3669 GNDA.n3627 4.5005
R10980 GNDA.n3673 GNDA.n3670 4.5005
R10981 GNDA.n3674 GNDA.n3626 4.5005
R10982 GNDA.n3678 GNDA.n3677 4.5005
R10983 GNDA.n3679 GNDA.n3625 4.5005
R10984 GNDA.n3683 GNDA.n3680 4.5005
R10985 GNDA.n3684 GNDA.n3624 4.5005
R10986 GNDA.n3688 GNDA.n3687 4.5005
R10987 GNDA.n3689 GNDA.n3623 4.5005
R10988 GNDA.n3693 GNDA.n3690 4.5005
R10989 GNDA.n3694 GNDA.n3622 4.5005
R10990 GNDA.n3698 GNDA.n3697 4.5005
R10991 GNDA.n3699 GNDA.n3621 4.5005
R10992 GNDA.n3703 GNDA.n3700 4.5005
R10993 GNDA.n3704 GNDA.n3620 4.5005
R10994 GNDA.n3708 GNDA.n3707 4.5005
R10995 GNDA.n3709 GNDA.n3619 4.5005
R10996 GNDA.n3713 GNDA.n3710 4.5005
R10997 GNDA.n3714 GNDA.n3618 4.5005
R10998 GNDA.n3718 GNDA.n3717 4.5005
R10999 GNDA.n3719 GNDA.n3617 4.5005
R11000 GNDA.n3723 GNDA.n3720 4.5005
R11001 GNDA.n3724 GNDA.n3616 4.5005
R11002 GNDA.n3728 GNDA.n3727 4.5005
R11003 GNDA.n3729 GNDA.n3615 4.5005
R11004 GNDA.n3733 GNDA.n3730 4.5005
R11005 GNDA.n3734 GNDA.n3614 4.5005
R11006 GNDA.n3738 GNDA.n3737 4.5005
R11007 GNDA.n3739 GNDA.n3613 4.5005
R11008 GNDA.n3743 GNDA.n3740 4.5005
R11009 GNDA.n3744 GNDA.n3612 4.5005
R11010 GNDA.n3748 GNDA.n3747 4.5005
R11011 GNDA.n3459 GNDA.n3458 4.5005
R11012 GNDA.n3296 GNDA.n3295 4.5005
R11013 GNDA.n3342 GNDA.n3297 4.5005
R11014 GNDA.n3343 GNDA.n3298 4.5005
R11015 GNDA.n3344 GNDA.n3299 4.5005
R11016 GNDA.n3345 GNDA.n3300 4.5005
R11017 GNDA.n3346 GNDA.n3301 4.5005
R11018 GNDA.n3347 GNDA.n3302 4.5005
R11019 GNDA.n3348 GNDA.n3303 4.5005
R11020 GNDA.n3349 GNDA.n3304 4.5005
R11021 GNDA.n3350 GNDA.n3305 4.5005
R11022 GNDA.n3351 GNDA.n3306 4.5005
R11023 GNDA.n3352 GNDA.n3307 4.5005
R11024 GNDA.n3353 GNDA.n3308 4.5005
R11025 GNDA.n3354 GNDA.n3309 4.5005
R11026 GNDA.n3355 GNDA.n3310 4.5005
R11027 GNDA.n3356 GNDA.n3311 4.5005
R11028 GNDA.n3357 GNDA.n3312 4.5005
R11029 GNDA.n3358 GNDA.n3313 4.5005
R11030 GNDA.n3359 GNDA.n3314 4.5005
R11031 GNDA.n3360 GNDA.n3315 4.5005
R11032 GNDA.n3361 GNDA.n3316 4.5005
R11033 GNDA.n3362 GNDA.n3317 4.5005
R11034 GNDA.n3363 GNDA.n3318 4.5005
R11035 GNDA.n3364 GNDA.n3319 4.5005
R11036 GNDA.n3365 GNDA.n3320 4.5005
R11037 GNDA.n3366 GNDA.n3321 4.5005
R11038 GNDA.n3367 GNDA.n3322 4.5005
R11039 GNDA.n3368 GNDA.n3323 4.5005
R11040 GNDA.n3369 GNDA.n3324 4.5005
R11041 GNDA.n3370 GNDA.n3325 4.5005
R11042 GNDA.n3371 GNDA.n3326 4.5005
R11043 GNDA.n3372 GNDA.n3327 4.5005
R11044 GNDA.n3373 GNDA.n3328 4.5005
R11045 GNDA.n3374 GNDA.n3329 4.5005
R11046 GNDA.n3375 GNDA.n3330 4.5005
R11047 GNDA.n3376 GNDA.n3331 4.5005
R11048 GNDA.n3377 GNDA.n3332 4.5005
R11049 GNDA.n3378 GNDA.n3333 4.5005
R11050 GNDA.n3379 GNDA.n3334 4.5005
R11051 GNDA.n3380 GNDA.n3335 4.5005
R11052 GNDA.n3381 GNDA.n3336 4.5005
R11053 GNDA.n3382 GNDA.n3337 4.5005
R11054 GNDA.n3383 GNDA.n3338 4.5005
R11055 GNDA.n3384 GNDA.n3339 4.5005
R11056 GNDA.n3385 GNDA.n3340 4.5005
R11057 GNDA.n5234 GNDA.n5233 4.5005
R11058 GNDA.n5070 GNDA.n5069 4.5005
R11059 GNDA.n5119 GNDA.n5118 4.5005
R11060 GNDA.n5123 GNDA.n5120 4.5005
R11061 GNDA.n5124 GNDA.n5117 4.5005
R11062 GNDA.n5128 GNDA.n5127 4.5005
R11063 GNDA.n5129 GNDA.n5116 4.5005
R11064 GNDA.n5133 GNDA.n5130 4.5005
R11065 GNDA.n5134 GNDA.n5115 4.5005
R11066 GNDA.n5138 GNDA.n5137 4.5005
R11067 GNDA.n5139 GNDA.n5114 4.5005
R11068 GNDA.n5143 GNDA.n5140 4.5005
R11069 GNDA.n5144 GNDA.n5113 4.5005
R11070 GNDA.n5148 GNDA.n5147 4.5005
R11071 GNDA.n5149 GNDA.n5112 4.5005
R11072 GNDA.n5153 GNDA.n5150 4.5005
R11073 GNDA.n5154 GNDA.n5111 4.5005
R11074 GNDA.n5158 GNDA.n5157 4.5005
R11075 GNDA.n5159 GNDA.n5110 4.5005
R11076 GNDA.n5163 GNDA.n5160 4.5005
R11077 GNDA.n5164 GNDA.n5109 4.5005
R11078 GNDA.n5168 GNDA.n5167 4.5005
R11079 GNDA.n5169 GNDA.n5108 4.5005
R11080 GNDA.n5173 GNDA.n5170 4.5005
R11081 GNDA.n5174 GNDA.n5107 4.5005
R11082 GNDA.n5178 GNDA.n5177 4.5005
R11083 GNDA.n5179 GNDA.n5106 4.5005
R11084 GNDA.n5183 GNDA.n5180 4.5005
R11085 GNDA.n5184 GNDA.n5105 4.5005
R11086 GNDA.n5188 GNDA.n5187 4.5005
R11087 GNDA.n5189 GNDA.n5104 4.5005
R11088 GNDA.n5193 GNDA.n5190 4.5005
R11089 GNDA.n5194 GNDA.n5103 4.5005
R11090 GNDA.n5198 GNDA.n5197 4.5005
R11091 GNDA.n5199 GNDA.n5102 4.5005
R11092 GNDA.n5203 GNDA.n5200 4.5005
R11093 GNDA.n5204 GNDA.n5101 4.5005
R11094 GNDA.n5208 GNDA.n5207 4.5005
R11095 GNDA.n5209 GNDA.n5100 4.5005
R11096 GNDA.n5213 GNDA.n5210 4.5005
R11097 GNDA.n5214 GNDA.n5099 4.5005
R11098 GNDA.n5218 GNDA.n5217 4.5005
R11099 GNDA.n5219 GNDA.n5098 4.5005
R11100 GNDA.n5223 GNDA.n5220 4.5005
R11101 GNDA.n5224 GNDA.n5097 4.5005
R11102 GNDA.n5228 GNDA.n5227 4.5005
R11103 GNDA.n5399 GNDA.n5398 4.5005
R11104 GNDA.n5236 GNDA.n5235 4.5005
R11105 GNDA.n5282 GNDA.n5237 4.5005
R11106 GNDA.n5283 GNDA.n5238 4.5005
R11107 GNDA.n5284 GNDA.n5239 4.5005
R11108 GNDA.n5285 GNDA.n5240 4.5005
R11109 GNDA.n5286 GNDA.n5241 4.5005
R11110 GNDA.n5287 GNDA.n5242 4.5005
R11111 GNDA.n5288 GNDA.n5243 4.5005
R11112 GNDA.n5289 GNDA.n5244 4.5005
R11113 GNDA.n5290 GNDA.n5245 4.5005
R11114 GNDA.n5291 GNDA.n5246 4.5005
R11115 GNDA.n5292 GNDA.n5247 4.5005
R11116 GNDA.n5293 GNDA.n5248 4.5005
R11117 GNDA.n5294 GNDA.n5249 4.5005
R11118 GNDA.n5295 GNDA.n5250 4.5005
R11119 GNDA.n5296 GNDA.n5251 4.5005
R11120 GNDA.n5297 GNDA.n5252 4.5005
R11121 GNDA.n5298 GNDA.n5253 4.5005
R11122 GNDA.n5299 GNDA.n5254 4.5005
R11123 GNDA.n5300 GNDA.n5255 4.5005
R11124 GNDA.n5301 GNDA.n5256 4.5005
R11125 GNDA.n5302 GNDA.n5257 4.5005
R11126 GNDA.n5303 GNDA.n5258 4.5005
R11127 GNDA.n5304 GNDA.n5259 4.5005
R11128 GNDA.n5305 GNDA.n5260 4.5005
R11129 GNDA.n5306 GNDA.n5261 4.5005
R11130 GNDA.n5307 GNDA.n5262 4.5005
R11131 GNDA.n5308 GNDA.n5263 4.5005
R11132 GNDA.n5309 GNDA.n5264 4.5005
R11133 GNDA.n5310 GNDA.n5265 4.5005
R11134 GNDA.n5311 GNDA.n5266 4.5005
R11135 GNDA.n5312 GNDA.n5267 4.5005
R11136 GNDA.n5313 GNDA.n5268 4.5005
R11137 GNDA.n5314 GNDA.n5269 4.5005
R11138 GNDA.n5315 GNDA.n5270 4.5005
R11139 GNDA.n5316 GNDA.n5271 4.5005
R11140 GNDA.n5317 GNDA.n5272 4.5005
R11141 GNDA.n5318 GNDA.n5273 4.5005
R11142 GNDA.n5319 GNDA.n5274 4.5005
R11143 GNDA.n5320 GNDA.n5275 4.5005
R11144 GNDA.n5321 GNDA.n5276 4.5005
R11145 GNDA.n5322 GNDA.n5277 4.5005
R11146 GNDA.n5323 GNDA.n5278 4.5005
R11147 GNDA.n5324 GNDA.n5279 4.5005
R11148 GNDA.n5325 GNDA.n5280 4.5005
R11149 GNDA.n5403 GNDA.n5402 4.5005
R11150 GNDA.n5406 GNDA.n5405 4.5005
R11151 GNDA.n5407 GNDA.n5068 4.5005
R11152 GNDA.n5411 GNDA.n5408 4.5005
R11153 GNDA.n5412 GNDA.n5067 4.5005
R11154 GNDA.n5416 GNDA.n5415 4.5005
R11155 GNDA.n5417 GNDA.n5066 4.5005
R11156 GNDA.n5421 GNDA.n5418 4.5005
R11157 GNDA.n5422 GNDA.n5065 4.5005
R11158 GNDA.n5426 GNDA.n5425 4.5005
R11159 GNDA.n5427 GNDA.n5064 4.5005
R11160 GNDA.n5431 GNDA.n5428 4.5005
R11161 GNDA.n5432 GNDA.n5063 4.5005
R11162 GNDA.n5436 GNDA.n5435 4.5005
R11163 GNDA.n5437 GNDA.n5062 4.5005
R11164 GNDA.n5441 GNDA.n5438 4.5005
R11165 GNDA.n5442 GNDA.n5061 4.5005
R11166 GNDA.n5446 GNDA.n5445 4.5005
R11167 GNDA.n5447 GNDA.n5060 4.5005
R11168 GNDA.n5451 GNDA.n5448 4.5005
R11169 GNDA.n5452 GNDA.n5059 4.5005
R11170 GNDA.n5456 GNDA.n5455 4.5005
R11171 GNDA.n5457 GNDA.n5058 4.5005
R11172 GNDA.n5461 GNDA.n5458 4.5005
R11173 GNDA.n5462 GNDA.n5057 4.5005
R11174 GNDA.n5466 GNDA.n5465 4.5005
R11175 GNDA.n5467 GNDA.n5056 4.5005
R11176 GNDA.n5471 GNDA.n5468 4.5005
R11177 GNDA.n5472 GNDA.n5055 4.5005
R11178 GNDA.n5476 GNDA.n5475 4.5005
R11179 GNDA.n5477 GNDA.n5054 4.5005
R11180 GNDA.n5481 GNDA.n5478 4.5005
R11181 GNDA.n5482 GNDA.n5053 4.5005
R11182 GNDA.n5486 GNDA.n5485 4.5005
R11183 GNDA.n5487 GNDA.n5052 4.5005
R11184 GNDA.n5491 GNDA.n5488 4.5005
R11185 GNDA.n5492 GNDA.n5051 4.5005
R11186 GNDA.n5496 GNDA.n5495 4.5005
R11187 GNDA.n5497 GNDA.n5050 4.5005
R11188 GNDA.n5501 GNDA.n5498 4.5005
R11189 GNDA.n5502 GNDA.n5049 4.5005
R11190 GNDA.n5506 GNDA.n5505 4.5005
R11191 GNDA.n5507 GNDA.n5048 4.5005
R11192 GNDA.n5511 GNDA.n5508 4.5005
R11193 GNDA.n5512 GNDA.n5047 4.5005
R11194 GNDA.n5516 GNDA.n5515 4.5005
R11195 GNDA.n5545 GNDA.n5544 4.5005
R11196 GNDA.n5548 GNDA.n5547 4.5005
R11197 GNDA.n5549 GNDA.n5543 4.5005
R11198 GNDA.n5553 GNDA.n5550 4.5005
R11199 GNDA.n5554 GNDA.n5542 4.5005
R11200 GNDA.n5558 GNDA.n5557 4.5005
R11201 GNDA.n5559 GNDA.n5541 4.5005
R11202 GNDA.n5563 GNDA.n5560 4.5005
R11203 GNDA.n5564 GNDA.n5540 4.5005
R11204 GNDA.n5568 GNDA.n5567 4.5005
R11205 GNDA.n5569 GNDA.n5539 4.5005
R11206 GNDA.n5573 GNDA.n5570 4.5005
R11207 GNDA.n5574 GNDA.n5538 4.5005
R11208 GNDA.n5578 GNDA.n5577 4.5005
R11209 GNDA.n5579 GNDA.n5537 4.5005
R11210 GNDA.n5583 GNDA.n5580 4.5005
R11211 GNDA.n5584 GNDA.n5536 4.5005
R11212 GNDA.n5588 GNDA.n5587 4.5005
R11213 GNDA.n5589 GNDA.n5535 4.5005
R11214 GNDA.n5593 GNDA.n5590 4.5005
R11215 GNDA.n5594 GNDA.n5534 4.5005
R11216 GNDA.n5598 GNDA.n5597 4.5005
R11217 GNDA.n5599 GNDA.n5533 4.5005
R11218 GNDA.n5603 GNDA.n5600 4.5005
R11219 GNDA.n5604 GNDA.n5532 4.5005
R11220 GNDA.n5608 GNDA.n5607 4.5005
R11221 GNDA.n5609 GNDA.n5531 4.5005
R11222 GNDA.n5613 GNDA.n5610 4.5005
R11223 GNDA.n5614 GNDA.n5530 4.5005
R11224 GNDA.n5618 GNDA.n5617 4.5005
R11225 GNDA.n5619 GNDA.n5529 4.5005
R11226 GNDA.n5623 GNDA.n5620 4.5005
R11227 GNDA.n5624 GNDA.n5528 4.5005
R11228 GNDA.n5628 GNDA.n5627 4.5005
R11229 GNDA.n5629 GNDA.n5527 4.5005
R11230 GNDA.n5633 GNDA.n5630 4.5005
R11231 GNDA.n5634 GNDA.n5526 4.5005
R11232 GNDA.n5638 GNDA.n5637 4.5005
R11233 GNDA.n5639 GNDA.n5525 4.5005
R11234 GNDA.n5643 GNDA.n5640 4.5005
R11235 GNDA.n5644 GNDA.n5524 4.5005
R11236 GNDA.n5648 GNDA.n5647 4.5005
R11237 GNDA.n5649 GNDA.n5523 4.5005
R11238 GNDA.n5653 GNDA.n5650 4.5005
R11239 GNDA.n5654 GNDA.n5522 4.5005
R11240 GNDA.n5658 GNDA.n5657 4.5005
R11241 GNDA.n5827 GNDA.n1363 4.5005
R11242 GNDA.n5830 GNDA.n5829 4.5005
R11243 GNDA.n5831 GNDA.n5826 4.5005
R11244 GNDA.n5835 GNDA.n5832 4.5005
R11245 GNDA.n5836 GNDA.n5825 4.5005
R11246 GNDA.n5840 GNDA.n5839 4.5005
R11247 GNDA.n5841 GNDA.n5824 4.5005
R11248 GNDA.n5845 GNDA.n5842 4.5005
R11249 GNDA.n5846 GNDA.n5823 4.5005
R11250 GNDA.n5850 GNDA.n5849 4.5005
R11251 GNDA.n5851 GNDA.n5822 4.5005
R11252 GNDA.n5855 GNDA.n5852 4.5005
R11253 GNDA.n5856 GNDA.n5821 4.5005
R11254 GNDA.n5860 GNDA.n5859 4.5005
R11255 GNDA.n5861 GNDA.n5820 4.5005
R11256 GNDA.n5865 GNDA.n5862 4.5005
R11257 GNDA.n5866 GNDA.n5819 4.5005
R11258 GNDA.n5870 GNDA.n5869 4.5005
R11259 GNDA.n5871 GNDA.n5818 4.5005
R11260 GNDA.n5875 GNDA.n5872 4.5005
R11261 GNDA.n5876 GNDA.n5817 4.5005
R11262 GNDA.n5880 GNDA.n5879 4.5005
R11263 GNDA.n5881 GNDA.n5816 4.5005
R11264 GNDA.n5885 GNDA.n5882 4.5005
R11265 GNDA.n5886 GNDA.n5815 4.5005
R11266 GNDA.n5890 GNDA.n5889 4.5005
R11267 GNDA.n5891 GNDA.n5814 4.5005
R11268 GNDA.n5895 GNDA.n5892 4.5005
R11269 GNDA.n5896 GNDA.n5813 4.5005
R11270 GNDA.n5900 GNDA.n5899 4.5005
R11271 GNDA.n5901 GNDA.n5812 4.5005
R11272 GNDA.n5905 GNDA.n5902 4.5005
R11273 GNDA.n5906 GNDA.n5811 4.5005
R11274 GNDA.n5910 GNDA.n5909 4.5005
R11275 GNDA.n5911 GNDA.n5810 4.5005
R11276 GNDA.n5915 GNDA.n5912 4.5005
R11277 GNDA.n5916 GNDA.n5809 4.5005
R11278 GNDA.n5920 GNDA.n5919 4.5005
R11279 GNDA.n5921 GNDA.n5808 4.5005
R11280 GNDA.n5925 GNDA.n5922 4.5005
R11281 GNDA.n5926 GNDA.n5807 4.5005
R11282 GNDA.n5930 GNDA.n5929 4.5005
R11283 GNDA.n5931 GNDA.n5806 4.5005
R11284 GNDA.n5935 GNDA.n5932 4.5005
R11285 GNDA.n5936 GNDA.n5805 4.5005
R11286 GNDA.n5940 GNDA.n5939 4.5005
R11287 GNDA.n4808 GNDA.n4807 4.5005
R11288 GNDA.n4811 GNDA.n4810 4.5005
R11289 GNDA.n4812 GNDA.n1419 4.5005
R11290 GNDA.n4816 GNDA.n4813 4.5005
R11291 GNDA.n4817 GNDA.n1418 4.5005
R11292 GNDA.n4821 GNDA.n4820 4.5005
R11293 GNDA.n4822 GNDA.n1417 4.5005
R11294 GNDA.n4826 GNDA.n4823 4.5005
R11295 GNDA.n4827 GNDA.n1416 4.5005
R11296 GNDA.n4831 GNDA.n4830 4.5005
R11297 GNDA.n4832 GNDA.n1415 4.5005
R11298 GNDA.n4836 GNDA.n4833 4.5005
R11299 GNDA.n4837 GNDA.n1414 4.5005
R11300 GNDA.n4841 GNDA.n4840 4.5005
R11301 GNDA.n4842 GNDA.n1413 4.5005
R11302 GNDA.n4846 GNDA.n4843 4.5005
R11303 GNDA.n4847 GNDA.n1412 4.5005
R11304 GNDA.n4851 GNDA.n4850 4.5005
R11305 GNDA.n4852 GNDA.n1411 4.5005
R11306 GNDA.n4856 GNDA.n4853 4.5005
R11307 GNDA.n4857 GNDA.n1410 4.5005
R11308 GNDA.n4861 GNDA.n4860 4.5005
R11309 GNDA.n4862 GNDA.n1409 4.5005
R11310 GNDA.n4866 GNDA.n4863 4.5005
R11311 GNDA.n4867 GNDA.n1408 4.5005
R11312 GNDA.n4871 GNDA.n4870 4.5005
R11313 GNDA.n4872 GNDA.n1407 4.5005
R11314 GNDA.n4876 GNDA.n4873 4.5005
R11315 GNDA.n4877 GNDA.n1406 4.5005
R11316 GNDA.n4881 GNDA.n4880 4.5005
R11317 GNDA.n4882 GNDA.n1405 4.5005
R11318 GNDA.n4886 GNDA.n4883 4.5005
R11319 GNDA.n4887 GNDA.n1404 4.5005
R11320 GNDA.n4891 GNDA.n4890 4.5005
R11321 GNDA.n4892 GNDA.n1403 4.5005
R11322 GNDA.n4896 GNDA.n4893 4.5005
R11323 GNDA.n4897 GNDA.n1402 4.5005
R11324 GNDA.n4901 GNDA.n4900 4.5005
R11325 GNDA.n4902 GNDA.n1401 4.5005
R11326 GNDA.n4906 GNDA.n4903 4.5005
R11327 GNDA.n4907 GNDA.n1400 4.5005
R11328 GNDA.n4911 GNDA.n4910 4.5005
R11329 GNDA.n4912 GNDA.n1399 4.5005
R11330 GNDA.n4916 GNDA.n4913 4.5005
R11331 GNDA.n4917 GNDA.n1398 4.5005
R11332 GNDA.n4921 GNDA.n4920 4.5005
R11333 GNDA.n4522 GNDA.n4521 4.5005
R11334 GNDA.n4525 GNDA.n4524 4.5005
R11335 GNDA.n4526 GNDA.n4520 4.5005
R11336 GNDA.n4530 GNDA.n4527 4.5005
R11337 GNDA.n4531 GNDA.n4519 4.5005
R11338 GNDA.n4535 GNDA.n4534 4.5005
R11339 GNDA.n4536 GNDA.n4518 4.5005
R11340 GNDA.n4540 GNDA.n4537 4.5005
R11341 GNDA.n4541 GNDA.n4517 4.5005
R11342 GNDA.n4545 GNDA.n4544 4.5005
R11343 GNDA.n4546 GNDA.n4516 4.5005
R11344 GNDA.n4550 GNDA.n4547 4.5005
R11345 GNDA.n4551 GNDA.n4515 4.5005
R11346 GNDA.n4555 GNDA.n4554 4.5005
R11347 GNDA.n4556 GNDA.n4514 4.5005
R11348 GNDA.n4560 GNDA.n4557 4.5005
R11349 GNDA.n4561 GNDA.n4513 4.5005
R11350 GNDA.n4565 GNDA.n4564 4.5005
R11351 GNDA.n4566 GNDA.n4512 4.5005
R11352 GNDA.n4570 GNDA.n4567 4.5005
R11353 GNDA.n4571 GNDA.n4511 4.5005
R11354 GNDA.n4575 GNDA.n4574 4.5005
R11355 GNDA.n4576 GNDA.n4510 4.5005
R11356 GNDA.n4580 GNDA.n4577 4.5005
R11357 GNDA.n4581 GNDA.n4509 4.5005
R11358 GNDA.n4585 GNDA.n4584 4.5005
R11359 GNDA.n4586 GNDA.n4508 4.5005
R11360 GNDA.n4590 GNDA.n4587 4.5005
R11361 GNDA.n4591 GNDA.n4507 4.5005
R11362 GNDA.n4595 GNDA.n4594 4.5005
R11363 GNDA.n4596 GNDA.n4506 4.5005
R11364 GNDA.n4600 GNDA.n4597 4.5005
R11365 GNDA.n4601 GNDA.n4505 4.5005
R11366 GNDA.n4605 GNDA.n4604 4.5005
R11367 GNDA.n4606 GNDA.n4504 4.5005
R11368 GNDA.n4610 GNDA.n4607 4.5005
R11369 GNDA.n4611 GNDA.n4503 4.5005
R11370 GNDA.n4615 GNDA.n4614 4.5005
R11371 GNDA.n4616 GNDA.n4502 4.5005
R11372 GNDA.n4620 GNDA.n4617 4.5005
R11373 GNDA.n4621 GNDA.n4501 4.5005
R11374 GNDA.n4625 GNDA.n4624 4.5005
R11375 GNDA.n4626 GNDA.n4500 4.5005
R11376 GNDA.n4630 GNDA.n4627 4.5005
R11377 GNDA.n4631 GNDA.n4499 4.5005
R11378 GNDA.n4635 GNDA.n4634 4.5005
R11379 GNDA.n4333 GNDA.n4332 4.5005
R11380 GNDA.n4336 GNDA.n4335 4.5005
R11381 GNDA.n4337 GNDA.n4331 4.5005
R11382 GNDA.n4341 GNDA.n4338 4.5005
R11383 GNDA.n4342 GNDA.n4330 4.5005
R11384 GNDA.n4346 GNDA.n4345 4.5005
R11385 GNDA.n4347 GNDA.n4329 4.5005
R11386 GNDA.n4351 GNDA.n4348 4.5005
R11387 GNDA.n4352 GNDA.n4328 4.5005
R11388 GNDA.n4356 GNDA.n4355 4.5005
R11389 GNDA.n4357 GNDA.n4327 4.5005
R11390 GNDA.n4361 GNDA.n4358 4.5005
R11391 GNDA.n4362 GNDA.n4326 4.5005
R11392 GNDA.n4366 GNDA.n4365 4.5005
R11393 GNDA.n4367 GNDA.n4325 4.5005
R11394 GNDA.n4371 GNDA.n4368 4.5005
R11395 GNDA.n4372 GNDA.n4324 4.5005
R11396 GNDA.n4376 GNDA.n4375 4.5005
R11397 GNDA.n4377 GNDA.n4323 4.5005
R11398 GNDA.n4381 GNDA.n4378 4.5005
R11399 GNDA.n4382 GNDA.n4322 4.5005
R11400 GNDA.n4386 GNDA.n4385 4.5005
R11401 GNDA.n4387 GNDA.n4321 4.5005
R11402 GNDA.n4391 GNDA.n4388 4.5005
R11403 GNDA.n4392 GNDA.n4320 4.5005
R11404 GNDA.n4396 GNDA.n4395 4.5005
R11405 GNDA.n4397 GNDA.n4319 4.5005
R11406 GNDA.n4401 GNDA.n4398 4.5005
R11407 GNDA.n4402 GNDA.n4318 4.5005
R11408 GNDA.n4406 GNDA.n4405 4.5005
R11409 GNDA.n4407 GNDA.n4317 4.5005
R11410 GNDA.n4411 GNDA.n4408 4.5005
R11411 GNDA.n4412 GNDA.n4316 4.5005
R11412 GNDA.n4416 GNDA.n4415 4.5005
R11413 GNDA.n4417 GNDA.n4315 4.5005
R11414 GNDA.n4421 GNDA.n4418 4.5005
R11415 GNDA.n4422 GNDA.n4314 4.5005
R11416 GNDA.n4426 GNDA.n4425 4.5005
R11417 GNDA.n4427 GNDA.n4313 4.5005
R11418 GNDA.n4431 GNDA.n4428 4.5005
R11419 GNDA.n4432 GNDA.n4312 4.5005
R11420 GNDA.n4436 GNDA.n4435 4.5005
R11421 GNDA.n4437 GNDA.n4311 4.5005
R11422 GNDA.n4441 GNDA.n4438 4.5005
R11423 GNDA.n4442 GNDA.n4310 4.5005
R11424 GNDA.n4446 GNDA.n4445 4.5005
R11425 GNDA.n4167 GNDA.n4166 4.5005
R11426 GNDA.n4170 GNDA.n4169 4.5005
R11427 GNDA.n4171 GNDA.n1647 4.5005
R11428 GNDA.n4175 GNDA.n4172 4.5005
R11429 GNDA.n4176 GNDA.n1646 4.5005
R11430 GNDA.n4180 GNDA.n4179 4.5005
R11431 GNDA.n4181 GNDA.n1645 4.5005
R11432 GNDA.n4185 GNDA.n4182 4.5005
R11433 GNDA.n4186 GNDA.n1644 4.5005
R11434 GNDA.n4190 GNDA.n4189 4.5005
R11435 GNDA.n4191 GNDA.n1643 4.5005
R11436 GNDA.n4195 GNDA.n4192 4.5005
R11437 GNDA.n4196 GNDA.n1642 4.5005
R11438 GNDA.n4200 GNDA.n4199 4.5005
R11439 GNDA.n4201 GNDA.n1641 4.5005
R11440 GNDA.n4205 GNDA.n4202 4.5005
R11441 GNDA.n4206 GNDA.n1640 4.5005
R11442 GNDA.n4210 GNDA.n4209 4.5005
R11443 GNDA.n4211 GNDA.n1639 4.5005
R11444 GNDA.n4215 GNDA.n4212 4.5005
R11445 GNDA.n4216 GNDA.n1638 4.5005
R11446 GNDA.n4220 GNDA.n4219 4.5005
R11447 GNDA.n4221 GNDA.n1637 4.5005
R11448 GNDA.n4225 GNDA.n4222 4.5005
R11449 GNDA.n4226 GNDA.n1636 4.5005
R11450 GNDA.n4230 GNDA.n4229 4.5005
R11451 GNDA.n4231 GNDA.n1635 4.5005
R11452 GNDA.n4235 GNDA.n4232 4.5005
R11453 GNDA.n4236 GNDA.n1634 4.5005
R11454 GNDA.n4240 GNDA.n4239 4.5005
R11455 GNDA.n4241 GNDA.n1633 4.5005
R11456 GNDA.n4245 GNDA.n4242 4.5005
R11457 GNDA.n4246 GNDA.n1632 4.5005
R11458 GNDA.n4250 GNDA.n4249 4.5005
R11459 GNDA.n4251 GNDA.n1631 4.5005
R11460 GNDA.n4255 GNDA.n4252 4.5005
R11461 GNDA.n4256 GNDA.n1630 4.5005
R11462 GNDA.n4260 GNDA.n4259 4.5005
R11463 GNDA.n4261 GNDA.n1629 4.5005
R11464 GNDA.n4265 GNDA.n4262 4.5005
R11465 GNDA.n4266 GNDA.n1628 4.5005
R11466 GNDA.n4270 GNDA.n4269 4.5005
R11467 GNDA.n4271 GNDA.n1627 4.5005
R11468 GNDA.n4275 GNDA.n4272 4.5005
R11469 GNDA.n4276 GNDA.n1626 4.5005
R11470 GNDA.n4280 GNDA.n4279 4.5005
R11471 GNDA.n1813 GNDA.n1812 4.5005
R11472 GNDA.n1650 GNDA.n1649 4.5005
R11473 GNDA.n1696 GNDA.n1651 4.5005
R11474 GNDA.n1697 GNDA.n1652 4.5005
R11475 GNDA.n1698 GNDA.n1653 4.5005
R11476 GNDA.n1699 GNDA.n1654 4.5005
R11477 GNDA.n1700 GNDA.n1655 4.5005
R11478 GNDA.n1701 GNDA.n1656 4.5005
R11479 GNDA.n1702 GNDA.n1657 4.5005
R11480 GNDA.n1703 GNDA.n1658 4.5005
R11481 GNDA.n1704 GNDA.n1659 4.5005
R11482 GNDA.n1705 GNDA.n1660 4.5005
R11483 GNDA.n1706 GNDA.n1661 4.5005
R11484 GNDA.n1707 GNDA.n1662 4.5005
R11485 GNDA.n1708 GNDA.n1663 4.5005
R11486 GNDA.n1709 GNDA.n1664 4.5005
R11487 GNDA.n1710 GNDA.n1665 4.5005
R11488 GNDA.n1711 GNDA.n1666 4.5005
R11489 GNDA.n1712 GNDA.n1667 4.5005
R11490 GNDA.n1713 GNDA.n1668 4.5005
R11491 GNDA.n1714 GNDA.n1669 4.5005
R11492 GNDA.n1715 GNDA.n1670 4.5005
R11493 GNDA.n1716 GNDA.n1671 4.5005
R11494 GNDA.n1717 GNDA.n1672 4.5005
R11495 GNDA.n1718 GNDA.n1673 4.5005
R11496 GNDA.n1719 GNDA.n1674 4.5005
R11497 GNDA.n1720 GNDA.n1675 4.5005
R11498 GNDA.n1721 GNDA.n1676 4.5005
R11499 GNDA.n1722 GNDA.n1677 4.5005
R11500 GNDA.n1723 GNDA.n1678 4.5005
R11501 GNDA.n1724 GNDA.n1679 4.5005
R11502 GNDA.n1725 GNDA.n1680 4.5005
R11503 GNDA.n1726 GNDA.n1681 4.5005
R11504 GNDA.n1727 GNDA.n1682 4.5005
R11505 GNDA.n1728 GNDA.n1683 4.5005
R11506 GNDA.n1729 GNDA.n1684 4.5005
R11507 GNDA.n1730 GNDA.n1685 4.5005
R11508 GNDA.n1731 GNDA.n1686 4.5005
R11509 GNDA.n1732 GNDA.n1687 4.5005
R11510 GNDA.n1733 GNDA.n1688 4.5005
R11511 GNDA.n1734 GNDA.n1689 4.5005
R11512 GNDA.n1735 GNDA.n1690 4.5005
R11513 GNDA.n1736 GNDA.n1691 4.5005
R11514 GNDA.n1737 GNDA.n1692 4.5005
R11515 GNDA.n1738 GNDA.n1693 4.5005
R11516 GNDA.n1739 GNDA.n1694 4.5005
R11517 GNDA.n3824 GNDA.n3823 4.5005
R11518 GNDA.n3827 GNDA.n3826 4.5005
R11519 GNDA.n3828 GNDA.n3822 4.5005
R11520 GNDA.n3832 GNDA.n3829 4.5005
R11521 GNDA.n3833 GNDA.n3821 4.5005
R11522 GNDA.n3837 GNDA.n3836 4.5005
R11523 GNDA.n3838 GNDA.n3820 4.5005
R11524 GNDA.n3842 GNDA.n3839 4.5005
R11525 GNDA.n3843 GNDA.n3819 4.5005
R11526 GNDA.n3847 GNDA.n3846 4.5005
R11527 GNDA.n3848 GNDA.n3818 4.5005
R11528 GNDA.n3852 GNDA.n3849 4.5005
R11529 GNDA.n3853 GNDA.n3817 4.5005
R11530 GNDA.n3857 GNDA.n3856 4.5005
R11531 GNDA.n3858 GNDA.n3816 4.5005
R11532 GNDA.n3862 GNDA.n3859 4.5005
R11533 GNDA.n3863 GNDA.n3815 4.5005
R11534 GNDA.n3867 GNDA.n3866 4.5005
R11535 GNDA.n3868 GNDA.n3814 4.5005
R11536 GNDA.n3872 GNDA.n3869 4.5005
R11537 GNDA.n3873 GNDA.n3813 4.5005
R11538 GNDA.n3877 GNDA.n3876 4.5005
R11539 GNDA.n3878 GNDA.n3812 4.5005
R11540 GNDA.n3882 GNDA.n3879 4.5005
R11541 GNDA.n3883 GNDA.n3811 4.5005
R11542 GNDA.n3887 GNDA.n3886 4.5005
R11543 GNDA.n3888 GNDA.n3810 4.5005
R11544 GNDA.n3892 GNDA.n3889 4.5005
R11545 GNDA.n3893 GNDA.n3809 4.5005
R11546 GNDA.n3897 GNDA.n3896 4.5005
R11547 GNDA.n3898 GNDA.n3808 4.5005
R11548 GNDA.n3902 GNDA.n3899 4.5005
R11549 GNDA.n3903 GNDA.n3807 4.5005
R11550 GNDA.n3907 GNDA.n3906 4.5005
R11551 GNDA.n3908 GNDA.n3806 4.5005
R11552 GNDA.n3912 GNDA.n3909 4.5005
R11553 GNDA.n3913 GNDA.n3805 4.5005
R11554 GNDA.n3917 GNDA.n3916 4.5005
R11555 GNDA.n3918 GNDA.n3804 4.5005
R11556 GNDA.n3922 GNDA.n3919 4.5005
R11557 GNDA.n3923 GNDA.n3803 4.5005
R11558 GNDA.n3927 GNDA.n3926 4.5005
R11559 GNDA.n3928 GNDA.n3802 4.5005
R11560 GNDA.n3932 GNDA.n3929 4.5005
R11561 GNDA.n3933 GNDA.n3801 4.5005
R11562 GNDA.n3937 GNDA.n3936 4.5005
R11563 GNDA.n4080 GNDA.n4079 4.5005
R11564 GNDA.n1836 GNDA.n1835 4.5005
R11565 GNDA.n3965 GNDA.n3964 4.5005
R11566 GNDA.n3969 GNDA.n3966 4.5005
R11567 GNDA.n3970 GNDA.n3963 4.5005
R11568 GNDA.n3974 GNDA.n3973 4.5005
R11569 GNDA.n3975 GNDA.n3962 4.5005
R11570 GNDA.n3979 GNDA.n3976 4.5005
R11571 GNDA.n3980 GNDA.n3961 4.5005
R11572 GNDA.n3984 GNDA.n3983 4.5005
R11573 GNDA.n3985 GNDA.n3960 4.5005
R11574 GNDA.n3989 GNDA.n3986 4.5005
R11575 GNDA.n3990 GNDA.n3959 4.5005
R11576 GNDA.n3994 GNDA.n3993 4.5005
R11577 GNDA.n3995 GNDA.n3958 4.5005
R11578 GNDA.n3999 GNDA.n3996 4.5005
R11579 GNDA.n4000 GNDA.n3957 4.5005
R11580 GNDA.n4004 GNDA.n4003 4.5005
R11581 GNDA.n4005 GNDA.n3956 4.5005
R11582 GNDA.n4009 GNDA.n4006 4.5005
R11583 GNDA.n4010 GNDA.n3955 4.5005
R11584 GNDA.n4014 GNDA.n4013 4.5005
R11585 GNDA.n4015 GNDA.n3954 4.5005
R11586 GNDA.n4019 GNDA.n4016 4.5005
R11587 GNDA.n4020 GNDA.n3953 4.5005
R11588 GNDA.n4024 GNDA.n4023 4.5005
R11589 GNDA.n4025 GNDA.n3952 4.5005
R11590 GNDA.n4029 GNDA.n4026 4.5005
R11591 GNDA.n4030 GNDA.n3951 4.5005
R11592 GNDA.n4034 GNDA.n4033 4.5005
R11593 GNDA.n4035 GNDA.n3950 4.5005
R11594 GNDA.n4039 GNDA.n4036 4.5005
R11595 GNDA.n4040 GNDA.n3949 4.5005
R11596 GNDA.n4044 GNDA.n4043 4.5005
R11597 GNDA.n4045 GNDA.n3948 4.5005
R11598 GNDA.n4049 GNDA.n4046 4.5005
R11599 GNDA.n4050 GNDA.n3947 4.5005
R11600 GNDA.n4054 GNDA.n4053 4.5005
R11601 GNDA.n4055 GNDA.n3946 4.5005
R11602 GNDA.n4059 GNDA.n4056 4.5005
R11603 GNDA.n4060 GNDA.n3945 4.5005
R11604 GNDA.n4064 GNDA.n4063 4.5005
R11605 GNDA.n4065 GNDA.n3944 4.5005
R11606 GNDA.n4069 GNDA.n4066 4.5005
R11607 GNDA.n4070 GNDA.n3943 4.5005
R11608 GNDA.n4074 GNDA.n4073 4.5005
R11609 GNDA.n3469 GNDA.n3468 4.5005
R11610 GNDA.n3472 GNDA.n3471 4.5005
R11611 GNDA.n3473 GNDA.n1886 4.5005
R11612 GNDA.n3477 GNDA.n3474 4.5005
R11613 GNDA.n3478 GNDA.n1885 4.5005
R11614 GNDA.n3482 GNDA.n3481 4.5005
R11615 GNDA.n3483 GNDA.n1884 4.5005
R11616 GNDA.n3487 GNDA.n3484 4.5005
R11617 GNDA.n3488 GNDA.n1883 4.5005
R11618 GNDA.n3492 GNDA.n3491 4.5005
R11619 GNDA.n3493 GNDA.n1882 4.5005
R11620 GNDA.n3497 GNDA.n3494 4.5005
R11621 GNDA.n3498 GNDA.n1881 4.5005
R11622 GNDA.n3502 GNDA.n3501 4.5005
R11623 GNDA.n3503 GNDA.n1880 4.5005
R11624 GNDA.n3507 GNDA.n3504 4.5005
R11625 GNDA.n3508 GNDA.n1879 4.5005
R11626 GNDA.n3512 GNDA.n3511 4.5005
R11627 GNDA.n3513 GNDA.n1878 4.5005
R11628 GNDA.n3517 GNDA.n3514 4.5005
R11629 GNDA.n3518 GNDA.n1877 4.5005
R11630 GNDA.n3522 GNDA.n3521 4.5005
R11631 GNDA.n3523 GNDA.n1876 4.5005
R11632 GNDA.n3527 GNDA.n3524 4.5005
R11633 GNDA.n3528 GNDA.n1875 4.5005
R11634 GNDA.n3532 GNDA.n3531 4.5005
R11635 GNDA.n3533 GNDA.n1874 4.5005
R11636 GNDA.n3537 GNDA.n3534 4.5005
R11637 GNDA.n3538 GNDA.n1873 4.5005
R11638 GNDA.n3542 GNDA.n3541 4.5005
R11639 GNDA.n3543 GNDA.n1872 4.5005
R11640 GNDA.n3547 GNDA.n3544 4.5005
R11641 GNDA.n3548 GNDA.n1871 4.5005
R11642 GNDA.n3552 GNDA.n3551 4.5005
R11643 GNDA.n3553 GNDA.n1870 4.5005
R11644 GNDA.n3557 GNDA.n3554 4.5005
R11645 GNDA.n3558 GNDA.n1869 4.5005
R11646 GNDA.n3562 GNDA.n3561 4.5005
R11647 GNDA.n3563 GNDA.n1868 4.5005
R11648 GNDA.n3567 GNDA.n3564 4.5005
R11649 GNDA.n3568 GNDA.n1867 4.5005
R11650 GNDA.n3572 GNDA.n3571 4.5005
R11651 GNDA.n3573 GNDA.n1866 4.5005
R11652 GNDA.n3577 GNDA.n3574 4.5005
R11653 GNDA.n3578 GNDA.n1865 4.5005
R11654 GNDA.n3582 GNDA.n3581 4.5005
R11655 GNDA.n2534 GNDA.n1887 4.5005
R11656 GNDA.n2537 GNDA.n2536 4.5005
R11657 GNDA.n2538 GNDA.n2533 4.5005
R11658 GNDA.n2542 GNDA.n2539 4.5005
R11659 GNDA.n2543 GNDA.n2532 4.5005
R11660 GNDA.n2547 GNDA.n2546 4.5005
R11661 GNDA.n2548 GNDA.n2531 4.5005
R11662 GNDA.n2552 GNDA.n2549 4.5005
R11663 GNDA.n2553 GNDA.n2530 4.5005
R11664 GNDA.n2557 GNDA.n2556 4.5005
R11665 GNDA.n2558 GNDA.n2529 4.5005
R11666 GNDA.n2562 GNDA.n2559 4.5005
R11667 GNDA.n2563 GNDA.n2528 4.5005
R11668 GNDA.n2567 GNDA.n2566 4.5005
R11669 GNDA.n2568 GNDA.n2527 4.5005
R11670 GNDA.n2572 GNDA.n2569 4.5005
R11671 GNDA.n2573 GNDA.n2526 4.5005
R11672 GNDA.n2577 GNDA.n2576 4.5005
R11673 GNDA.n2578 GNDA.n2525 4.5005
R11674 GNDA.n2582 GNDA.n2579 4.5005
R11675 GNDA.n2583 GNDA.n2524 4.5005
R11676 GNDA.n2587 GNDA.n2586 4.5005
R11677 GNDA.n2588 GNDA.n2523 4.5005
R11678 GNDA.n2592 GNDA.n2589 4.5005
R11679 GNDA.n2593 GNDA.n2522 4.5005
R11680 GNDA.n2597 GNDA.n2596 4.5005
R11681 GNDA.n2598 GNDA.n2521 4.5005
R11682 GNDA.n2602 GNDA.n2599 4.5005
R11683 GNDA.n2603 GNDA.n2520 4.5005
R11684 GNDA.n2607 GNDA.n2606 4.5005
R11685 GNDA.n2608 GNDA.n2519 4.5005
R11686 GNDA.n2612 GNDA.n2609 4.5005
R11687 GNDA.n2613 GNDA.n2518 4.5005
R11688 GNDA.n2617 GNDA.n2616 4.5005
R11689 GNDA.n2618 GNDA.n2517 4.5005
R11690 GNDA.n2622 GNDA.n2619 4.5005
R11691 GNDA.n2623 GNDA.n2516 4.5005
R11692 GNDA.n2627 GNDA.n2626 4.5005
R11693 GNDA.n2628 GNDA.n2515 4.5005
R11694 GNDA.n2632 GNDA.n2629 4.5005
R11695 GNDA.n2633 GNDA.n2514 4.5005
R11696 GNDA.n2637 GNDA.n2636 4.5005
R11697 GNDA.n2638 GNDA.n2513 4.5005
R11698 GNDA.n2642 GNDA.n2639 4.5005
R11699 GNDA.n2643 GNDA.n2512 4.5005
R11700 GNDA.n2647 GNDA.n2646 4.5005
R11701 GNDA.n2817 GNDA.n1889 4.5005
R11702 GNDA.n2820 GNDA.n2819 4.5005
R11703 GNDA.n2821 GNDA.n2816 4.5005
R11704 GNDA.n2825 GNDA.n2822 4.5005
R11705 GNDA.n2826 GNDA.n2815 4.5005
R11706 GNDA.n2830 GNDA.n2829 4.5005
R11707 GNDA.n2831 GNDA.n2814 4.5005
R11708 GNDA.n2835 GNDA.n2832 4.5005
R11709 GNDA.n2836 GNDA.n2813 4.5005
R11710 GNDA.n2840 GNDA.n2839 4.5005
R11711 GNDA.n2841 GNDA.n2812 4.5005
R11712 GNDA.n2845 GNDA.n2842 4.5005
R11713 GNDA.n2846 GNDA.n2811 4.5005
R11714 GNDA.n2850 GNDA.n2849 4.5005
R11715 GNDA.n2851 GNDA.n2810 4.5005
R11716 GNDA.n2855 GNDA.n2852 4.5005
R11717 GNDA.n2856 GNDA.n2809 4.5005
R11718 GNDA.n2860 GNDA.n2859 4.5005
R11719 GNDA.n2861 GNDA.n2808 4.5005
R11720 GNDA.n2865 GNDA.n2862 4.5005
R11721 GNDA.n2866 GNDA.n2807 4.5005
R11722 GNDA.n2870 GNDA.n2869 4.5005
R11723 GNDA.n2871 GNDA.n2806 4.5005
R11724 GNDA.n2875 GNDA.n2872 4.5005
R11725 GNDA.n2876 GNDA.n2805 4.5005
R11726 GNDA.n2880 GNDA.n2879 4.5005
R11727 GNDA.n2881 GNDA.n2804 4.5005
R11728 GNDA.n2885 GNDA.n2882 4.5005
R11729 GNDA.n2886 GNDA.n2803 4.5005
R11730 GNDA.n2890 GNDA.n2889 4.5005
R11731 GNDA.n2891 GNDA.n2802 4.5005
R11732 GNDA.n2895 GNDA.n2892 4.5005
R11733 GNDA.n2896 GNDA.n2801 4.5005
R11734 GNDA.n2900 GNDA.n2899 4.5005
R11735 GNDA.n2901 GNDA.n2800 4.5005
R11736 GNDA.n2905 GNDA.n2902 4.5005
R11737 GNDA.n2906 GNDA.n2799 4.5005
R11738 GNDA.n2910 GNDA.n2909 4.5005
R11739 GNDA.n2911 GNDA.n2798 4.5005
R11740 GNDA.n2915 GNDA.n2912 4.5005
R11741 GNDA.n2916 GNDA.n2797 4.5005
R11742 GNDA.n2920 GNDA.n2919 4.5005
R11743 GNDA.n2921 GNDA.n2796 4.5005
R11744 GNDA.n2925 GNDA.n2922 4.5005
R11745 GNDA.n2926 GNDA.n2795 4.5005
R11746 GNDA.n2930 GNDA.n2929 4.5005
R11747 GNDA.n2958 GNDA.n1890 4.5005
R11748 GNDA.n2961 GNDA.n2960 4.5005
R11749 GNDA.n2962 GNDA.n2957 4.5005
R11750 GNDA.n2966 GNDA.n2963 4.5005
R11751 GNDA.n2967 GNDA.n2956 4.5005
R11752 GNDA.n2971 GNDA.n2970 4.5005
R11753 GNDA.n2972 GNDA.n2955 4.5005
R11754 GNDA.n2976 GNDA.n2973 4.5005
R11755 GNDA.n2977 GNDA.n2954 4.5005
R11756 GNDA.n2981 GNDA.n2980 4.5005
R11757 GNDA.n2982 GNDA.n2953 4.5005
R11758 GNDA.n2986 GNDA.n2983 4.5005
R11759 GNDA.n2987 GNDA.n2952 4.5005
R11760 GNDA.n2991 GNDA.n2990 4.5005
R11761 GNDA.n2992 GNDA.n2951 4.5005
R11762 GNDA.n2996 GNDA.n2993 4.5005
R11763 GNDA.n2997 GNDA.n2950 4.5005
R11764 GNDA.n3001 GNDA.n3000 4.5005
R11765 GNDA.n3002 GNDA.n2949 4.5005
R11766 GNDA.n3006 GNDA.n3003 4.5005
R11767 GNDA.n3007 GNDA.n2948 4.5005
R11768 GNDA.n3011 GNDA.n3010 4.5005
R11769 GNDA.n3012 GNDA.n2947 4.5005
R11770 GNDA.n3016 GNDA.n3013 4.5005
R11771 GNDA.n3017 GNDA.n2946 4.5005
R11772 GNDA.n3021 GNDA.n3020 4.5005
R11773 GNDA.n3022 GNDA.n2945 4.5005
R11774 GNDA.n3026 GNDA.n3023 4.5005
R11775 GNDA.n3027 GNDA.n2944 4.5005
R11776 GNDA.n3031 GNDA.n3030 4.5005
R11777 GNDA.n3032 GNDA.n2943 4.5005
R11778 GNDA.n3036 GNDA.n3033 4.5005
R11779 GNDA.n3037 GNDA.n2942 4.5005
R11780 GNDA.n3041 GNDA.n3040 4.5005
R11781 GNDA.n3042 GNDA.n2941 4.5005
R11782 GNDA.n3046 GNDA.n3043 4.5005
R11783 GNDA.n3047 GNDA.n2940 4.5005
R11784 GNDA.n3051 GNDA.n3050 4.5005
R11785 GNDA.n3052 GNDA.n2939 4.5005
R11786 GNDA.n3056 GNDA.n3053 4.5005
R11787 GNDA.n3057 GNDA.n2938 4.5005
R11788 GNDA.n3061 GNDA.n3060 4.5005
R11789 GNDA.n3062 GNDA.n2937 4.5005
R11790 GNDA.n3066 GNDA.n3063 4.5005
R11791 GNDA.n3067 GNDA.n2936 4.5005
R11792 GNDA.n3071 GNDA.n3070 4.5005
R11793 GNDA.n3099 GNDA.n1891 4.5005
R11794 GNDA.n3102 GNDA.n3101 4.5005
R11795 GNDA.n3103 GNDA.n3098 4.5005
R11796 GNDA.n3107 GNDA.n3104 4.5005
R11797 GNDA.n3108 GNDA.n3097 4.5005
R11798 GNDA.n3112 GNDA.n3111 4.5005
R11799 GNDA.n3113 GNDA.n3096 4.5005
R11800 GNDA.n3117 GNDA.n3114 4.5005
R11801 GNDA.n3118 GNDA.n3095 4.5005
R11802 GNDA.n3122 GNDA.n3121 4.5005
R11803 GNDA.n3123 GNDA.n3094 4.5005
R11804 GNDA.n3127 GNDA.n3124 4.5005
R11805 GNDA.n3128 GNDA.n3093 4.5005
R11806 GNDA.n3132 GNDA.n3131 4.5005
R11807 GNDA.n3133 GNDA.n3092 4.5005
R11808 GNDA.n3137 GNDA.n3134 4.5005
R11809 GNDA.n3138 GNDA.n3091 4.5005
R11810 GNDA.n3142 GNDA.n3141 4.5005
R11811 GNDA.n3143 GNDA.n3090 4.5005
R11812 GNDA.n3147 GNDA.n3144 4.5005
R11813 GNDA.n3148 GNDA.n3089 4.5005
R11814 GNDA.n3152 GNDA.n3151 4.5005
R11815 GNDA.n3153 GNDA.n3088 4.5005
R11816 GNDA.n3157 GNDA.n3154 4.5005
R11817 GNDA.n3158 GNDA.n3087 4.5005
R11818 GNDA.n3162 GNDA.n3161 4.5005
R11819 GNDA.n3163 GNDA.n3086 4.5005
R11820 GNDA.n3167 GNDA.n3164 4.5005
R11821 GNDA.n3168 GNDA.n3085 4.5005
R11822 GNDA.n3172 GNDA.n3171 4.5005
R11823 GNDA.n3173 GNDA.n3084 4.5005
R11824 GNDA.n3177 GNDA.n3174 4.5005
R11825 GNDA.n3178 GNDA.n3083 4.5005
R11826 GNDA.n3182 GNDA.n3181 4.5005
R11827 GNDA.n3183 GNDA.n3082 4.5005
R11828 GNDA.n3187 GNDA.n3184 4.5005
R11829 GNDA.n3188 GNDA.n3081 4.5005
R11830 GNDA.n3192 GNDA.n3191 4.5005
R11831 GNDA.n3193 GNDA.n3080 4.5005
R11832 GNDA.n3197 GNDA.n3194 4.5005
R11833 GNDA.n3198 GNDA.n3079 4.5005
R11834 GNDA.n3202 GNDA.n3201 4.5005
R11835 GNDA.n3203 GNDA.n3078 4.5005
R11836 GNDA.n3207 GNDA.n3204 4.5005
R11837 GNDA.n3208 GNDA.n3077 4.5005
R11838 GNDA.n3212 GNDA.n3211 4.5005
R11839 GNDA.n3288 GNDA.n3287 4.5005
R11840 GNDA.n3286 GNDA.n1892 4.5005
R11841 GNDA.n3285 GNDA.n3284 4.5005
R11842 GNDA.n3283 GNDA.n1896 4.5005
R11843 GNDA.n3282 GNDA.n3281 4.5005
R11844 GNDA.n3280 GNDA.n1897 4.5005
R11845 GNDA.n3279 GNDA.n3278 4.5005
R11846 GNDA.n3277 GNDA.n1901 4.5005
R11847 GNDA.n3276 GNDA.n3275 4.5005
R11848 GNDA.n3274 GNDA.n1902 4.5005
R11849 GNDA.n3273 GNDA.n3272 4.5005
R11850 GNDA.n3271 GNDA.n1906 4.5005
R11851 GNDA.n3270 GNDA.n3269 4.5005
R11852 GNDA.n3268 GNDA.n1907 4.5005
R11853 GNDA.n3267 GNDA.n3266 4.5005
R11854 GNDA.n3265 GNDA.n1911 4.5005
R11855 GNDA.n3264 GNDA.n3263 4.5005
R11856 GNDA.n3262 GNDA.n1912 4.5005
R11857 GNDA.n3261 GNDA.n3260 4.5005
R11858 GNDA.n3259 GNDA.n1916 4.5005
R11859 GNDA.n3258 GNDA.n3257 4.5005
R11860 GNDA.n3256 GNDA.n1917 4.5005
R11861 GNDA.n3255 GNDA.n3254 4.5005
R11862 GNDA.n3253 GNDA.n1921 4.5005
R11863 GNDA.n3252 GNDA.n3251 4.5005
R11864 GNDA.n3250 GNDA.n1922 4.5005
R11865 GNDA.n3249 GNDA.n3248 4.5005
R11866 GNDA.n3247 GNDA.n1926 4.5005
R11867 GNDA.n3246 GNDA.n3245 4.5005
R11868 GNDA.n3244 GNDA.n1927 4.5005
R11869 GNDA.n3243 GNDA.n3242 4.5005
R11870 GNDA.n3241 GNDA.n1931 4.5005
R11871 GNDA.n3240 GNDA.n3239 4.5005
R11872 GNDA.n3238 GNDA.n1932 4.5005
R11873 GNDA.n3237 GNDA.n3236 4.5005
R11874 GNDA.n3235 GNDA.n1936 4.5005
R11875 GNDA.n3234 GNDA.n3233 4.5005
R11876 GNDA.n3232 GNDA.n1937 4.5005
R11877 GNDA.n3231 GNDA.n3230 4.5005
R11878 GNDA.n3229 GNDA.n1941 4.5005
R11879 GNDA.n3228 GNDA.n3227 4.5005
R11880 GNDA.n3226 GNDA.n1942 4.5005
R11881 GNDA.n3225 GNDA.n3224 4.5005
R11882 GNDA.n3223 GNDA.n1946 4.5005
R11883 GNDA.n3222 GNDA.n3221 4.5005
R11884 GNDA.n3220 GNDA.n1947 4.5005
R11885 GNDA.n3464 GNDA.n3463 4.5005
R11886 GNDA.n4084 GNDA.n4083 4.5005
R11887 GNDA.n4803 GNDA.n4802 4.5005
R11888 GNDA.n1367 GNDA.n1364 4.5005
R11889 GNDA.n2698 GNDA.n2697 4.5005
R11890 GNDA.n2701 GNDA.n2700 4.5005
R11891 GNDA.n2702 GNDA.n2694 4.5005
R11892 GNDA.n2704 GNDA.n2703 4.5005
R11893 GNDA.n2705 GNDA.n2693 4.5005
R11894 GNDA.n2709 GNDA.n2708 4.5005
R11895 GNDA.n2710 GNDA.n2690 4.5005
R11896 GNDA.n2712 GNDA.n2711 4.5005
R11897 GNDA.n2713 GNDA.n2689 4.5005
R11898 GNDA.n2717 GNDA.n2716 4.5005
R11899 GNDA.n2718 GNDA.n2686 4.5005
R11900 GNDA.n2720 GNDA.n2719 4.5005
R11901 GNDA.n2721 GNDA.n2685 4.5005
R11902 GNDA.n2725 GNDA.n2724 4.5005
R11903 GNDA.n2726 GNDA.n2682 4.5005
R11904 GNDA.n2728 GNDA.n2727 4.5005
R11905 GNDA.n2729 GNDA.n2681 4.5005
R11906 GNDA.n2733 GNDA.n2732 4.5005
R11907 GNDA.n2734 GNDA.n2678 4.5005
R11908 GNDA.n2736 GNDA.n2735 4.5005
R11909 GNDA.n2737 GNDA.n2677 4.5005
R11910 GNDA.n2741 GNDA.n2740 4.5005
R11911 GNDA.n2742 GNDA.n2674 4.5005
R11912 GNDA.n2744 GNDA.n2743 4.5005
R11913 GNDA.n2745 GNDA.n2673 4.5005
R11914 GNDA.n2749 GNDA.n2748 4.5005
R11915 GNDA.n2750 GNDA.n2670 4.5005
R11916 GNDA.n2752 GNDA.n2751 4.5005
R11917 GNDA.n2753 GNDA.n2669 4.5005
R11918 GNDA.n2757 GNDA.n2756 4.5005
R11919 GNDA.n2758 GNDA.n2666 4.5005
R11920 GNDA.n2760 GNDA.n2759 4.5005
R11921 GNDA.n2761 GNDA.n2665 4.5005
R11922 GNDA.n2765 GNDA.n2764 4.5005
R11923 GNDA.n2766 GNDA.n2662 4.5005
R11924 GNDA.n2768 GNDA.n2767 4.5005
R11925 GNDA.n2769 GNDA.n2661 4.5005
R11926 GNDA.n2773 GNDA.n2772 4.5005
R11927 GNDA.n2774 GNDA.n2658 4.5005
R11928 GNDA.n2776 GNDA.n2775 4.5005
R11929 GNDA.n2777 GNDA.n2657 4.5005
R11930 GNDA.n2781 GNDA.n2780 4.5005
R11931 GNDA.n2782 GNDA.n2654 4.5005
R11932 GNDA.n2784 GNDA.n2783 4.5005
R11933 GNDA.n2785 GNDA.n2653 4.5005
R11934 GNDA.n2789 GNDA.n2788 4.5005
R11935 GNDA.n4121 GNDA.n4120 4.5005
R11936 GNDA.n6356 GNDA.n6352 4.5005
R11937 GNDA.n6360 GNDA.n6359 4.5005
R11938 GNDA.n6361 GNDA.n6349 4.5005
R11939 GNDA.n6363 GNDA.n6362 4.5005
R11940 GNDA.n6364 GNDA.n6348 4.5005
R11941 GNDA.n6368 GNDA.n6367 4.5005
R11942 GNDA.n6369 GNDA.n6345 4.5005
R11943 GNDA.n6371 GNDA.n6370 4.5005
R11944 GNDA.n6372 GNDA.n6344 4.5005
R11945 GNDA.n6376 GNDA.n6375 4.5005
R11946 GNDA.n6377 GNDA.n6341 4.5005
R11947 GNDA.n6379 GNDA.n6378 4.5005
R11948 GNDA.n6380 GNDA.n6340 4.5005
R11949 GNDA.n6384 GNDA.n6383 4.5005
R11950 GNDA.n6385 GNDA.n6337 4.5005
R11951 GNDA.n6387 GNDA.n6386 4.5005
R11952 GNDA.n6388 GNDA.n6336 4.5005
R11953 GNDA.n6392 GNDA.n6391 4.5005
R11954 GNDA.n6393 GNDA.n6333 4.5005
R11955 GNDA.n6395 GNDA.n6394 4.5005
R11956 GNDA.n6396 GNDA.n6332 4.5005
R11957 GNDA.n6400 GNDA.n6399 4.5005
R11958 GNDA.n6401 GNDA.n6329 4.5005
R11959 GNDA.n6403 GNDA.n6402 4.5005
R11960 GNDA.n6404 GNDA.n6328 4.5005
R11961 GNDA.n6408 GNDA.n6407 4.5005
R11962 GNDA.n6409 GNDA.n6325 4.5005
R11963 GNDA.n6411 GNDA.n6410 4.5005
R11964 GNDA.n6412 GNDA.n6324 4.5005
R11965 GNDA.n6416 GNDA.n6415 4.5005
R11966 GNDA.n6417 GNDA.n6321 4.5005
R11967 GNDA.n6419 GNDA.n6418 4.5005
R11968 GNDA.n6420 GNDA.n6320 4.5005
R11969 GNDA.n6424 GNDA.n6423 4.5005
R11970 GNDA.n6425 GNDA.n6317 4.5005
R11971 GNDA.n6427 GNDA.n6426 4.5005
R11972 GNDA.n6428 GNDA.n6316 4.5005
R11973 GNDA.n6432 GNDA.n6431 4.5005
R11974 GNDA.n6433 GNDA.n6313 4.5005
R11975 GNDA.n6435 GNDA.n6434 4.5005
R11976 GNDA.n6436 GNDA.n6312 4.5005
R11977 GNDA.n6440 GNDA.n6439 4.5005
R11978 GNDA.n6441 GNDA.n6311 4.5005
R11979 GNDA.n6443 GNDA.n6442 4.5005
R11980 GNDA.n359 GNDA.n358 4.5005
R11981 GNDA.n6618 GNDA.n6617 4.5005
R11982 GNDA.n413 GNDA.n409 4.5005
R11983 GNDA.n417 GNDA.n414 4.5005
R11984 GNDA.n418 GNDA.n408 4.5005
R11985 GNDA.n422 GNDA.n421 4.5005
R11986 GNDA.n423 GNDA.n407 4.5005
R11987 GNDA.n427 GNDA.n424 4.5005
R11988 GNDA.n428 GNDA.n406 4.5005
R11989 GNDA.n432 GNDA.n431 4.5005
R11990 GNDA.n433 GNDA.n405 4.5005
R11991 GNDA.n437 GNDA.n434 4.5005
R11992 GNDA.n438 GNDA.n404 4.5005
R11993 GNDA.n442 GNDA.n441 4.5005
R11994 GNDA.n443 GNDA.n403 4.5005
R11995 GNDA.n447 GNDA.n444 4.5005
R11996 GNDA.n448 GNDA.n402 4.5005
R11997 GNDA.n452 GNDA.n451 4.5005
R11998 GNDA.n453 GNDA.n401 4.5005
R11999 GNDA.n457 GNDA.n454 4.5005
R12000 GNDA.n458 GNDA.n400 4.5005
R12001 GNDA.n462 GNDA.n461 4.5005
R12002 GNDA.n463 GNDA.n399 4.5005
R12003 GNDA.n467 GNDA.n464 4.5005
R12004 GNDA.n468 GNDA.n398 4.5005
R12005 GNDA.n472 GNDA.n471 4.5005
R12006 GNDA.n473 GNDA.n397 4.5005
R12007 GNDA.n477 GNDA.n474 4.5005
R12008 GNDA.n478 GNDA.n396 4.5005
R12009 GNDA.n482 GNDA.n481 4.5005
R12010 GNDA.n483 GNDA.n395 4.5005
R12011 GNDA.n487 GNDA.n484 4.5005
R12012 GNDA.n488 GNDA.n394 4.5005
R12013 GNDA.n492 GNDA.n491 4.5005
R12014 GNDA.n493 GNDA.n393 4.5005
R12015 GNDA.n497 GNDA.n494 4.5005
R12016 GNDA.n498 GNDA.n392 4.5005
R12017 GNDA.n502 GNDA.n501 4.5005
R12018 GNDA.n503 GNDA.n391 4.5005
R12019 GNDA.n507 GNDA.n504 4.5005
R12020 GNDA.n508 GNDA.n390 4.5005
R12021 GNDA.n512 GNDA.n511 4.5005
R12022 GNDA.n513 GNDA.n389 4.5005
R12023 GNDA.n517 GNDA.n514 4.5005
R12024 GNDA.n518 GNDA.n388 4.5005
R12025 GNDA.n522 GNDA.n521 4.5005
R12026 GNDA.n523 GNDA.n387 4.5005
R12027 GNDA.n6284 GNDA.n6283 4.5005
R12028 GNDA.n6446 GNDA.t1045 4.5005
R12029 GNDA.n6447 GNDA.t988 4.5005
R12030 GNDA.n6448 GNDA.t1019 4.5005
R12031 GNDA.n6452 GNDA.t1012 4.5005
R12032 GNDA.n6451 GNDA.t1084 4.5005
R12033 GNDA.n6450 GNDA.t926 4.5005
R12034 GNDA.n6449 GNDA.t890 4.5005
R12035 GNDA.n6453 GNDA.t1095 4.5005
R12036 GNDA.n6454 GNDA.t1038 4.5005
R12037 GNDA.n6455 GNDA.t1075 4.5005
R12038 GNDA.n6459 GNDA.t1066 4.5005
R12039 GNDA.n6458 GNDA.t923 4.5005
R12040 GNDA.n6457 GNDA.t975 4.5005
R12041 GNDA.n6456 GNDA.t940 4.5005
R12042 GNDA.n6460 GNDA.t943 4.5005
R12043 GNDA.n6461 GNDA.t884 4.5005
R12044 GNDA.n6462 GNDA.t921 4.5005
R12045 GNDA.n6466 GNDA.t911 4.5005
R12046 GNDA.n6465 GNDA.t984 4.5005
R12047 GNDA.n6464 GNDA.t1035 4.5005
R12048 GNDA.n6463 GNDA.t1003 4.5005
R12049 GNDA.n6467 GNDA.t1006 4.5005
R12050 GNDA.n6468 GNDA.t947 4.5005
R12051 GNDA.n6469 GNDA.t982 4.5005
R12052 GNDA.n6473 GNDA.t971 4.5005
R12053 GNDA.n6472 GNDA.t1044 4.5005
R12054 GNDA.n6471 GNDA.t1097 4.5005
R12055 GNDA.n6470 GNDA.t1065 4.5005
R12056 GNDA.n6474 GNDA.t953 4.5005
R12057 GNDA.n6475 GNDA.t893 4.5005
R12058 GNDA.n6476 GNDA.t929 4.5005
R12059 GNDA.n6480 GNDA.t919 4.5005
R12060 GNDA.n6479 GNDA.t992 4.5005
R12061 GNDA.n6478 GNDA.t1046 4.5005
R12062 GNDA.n6477 GNDA.t1011 4.5005
R12063 GNDA.n6481 GNDA.t1014 4.5005
R12064 GNDA.n6482 GNDA.t955 4.5005
R12065 GNDA.n6483 GNDA.t991 4.5005
R12066 GNDA.n6487 GNDA.t979 4.5005
R12067 GNDA.n6486 GNDA.t1051 4.5005
R12068 GNDA.n6485 GNDA.t892 4.5005
R12069 GNDA.n6484 GNDA.t1074 4.5005
R12070 GNDA.n6488 GNDA.t1076 4.5005
R12071 GNDA.n6489 GNDA.t1016 4.5005
R12072 GNDA.n6490 GNDA.t1050 4.5005
R12073 GNDA.n6494 GNDA.t1041 4.5005
R12074 GNDA.n6493 GNDA.t896 4.5005
R12075 GNDA.n6492 GNDA.t954 4.5005
R12076 GNDA.n6491 GNDA.t918 4.5005
R12077 GNDA.n6495 GNDA.t1020 4.5005
R12078 GNDA.n6496 GNDA.t962 4.5005
R12079 GNDA.n6497 GNDA.t996 4.5005
R12080 GNDA.n6501 GNDA.t990 4.5005
R12081 GNDA.n6500 GNDA.t1059 4.5005
R12082 GNDA.n6499 GNDA.t897 4.5005
R12083 GNDA.n6498 GNDA.t1081 4.5005
R12084 GNDA.n6502 GNDA.t1083 4.5005
R12085 GNDA.n6503 GNDA.t1023 4.5005
R12086 GNDA.n6504 GNDA.t1057 4.5005
R12087 GNDA.n6508 GNDA.t1049 4.5005
R12088 GNDA.n6507 GNDA.t906 4.5005
R12089 GNDA.n6506 GNDA.t958 4.5005
R12090 GNDA.n6505 GNDA.t928 4.5005
R12091 GNDA.n6509 GNDA.t931 4.5005
R12092 GNDA.n6510 GNDA.t1085 4.5005
R12093 GNDA.n6511 GNDA.t905 4.5005
R12094 GNDA.n6515 GNDA.t895 4.5005
R12095 GNDA.n6514 GNDA.t965 4.5005
R12096 GNDA.n6513 GNDA.t1021 4.5005
R12097 GNDA.n6512 GNDA.t989 4.5005
R12098 GNDA.n6516 GNDA.t1087 4.5005
R12099 GNDA.n6517 GNDA.t1029 4.5005
R12100 GNDA.n6518 GNDA.t1067 4.5005
R12101 GNDA.n6522 GNDA.t1055 4.5005
R12102 GNDA.n6521 GNDA.t914 4.5005
R12103 GNDA.n6520 GNDA.t967 4.5005
R12104 GNDA.n6519 GNDA.t933 4.5005
R12105 GNDA.n6523 GNDA.t934 4.5005
R12106 GNDA.n6524 GNDA.t1090 4.5005
R12107 GNDA.n6525 GNDA.t912 4.5005
R12108 GNDA.n6529 GNDA.t903 4.5005
R12109 GNDA.n6528 GNDA.t974 4.5005
R12110 GNDA.n6527 GNDA.t1027 4.5005
R12111 GNDA.n6526 GNDA.t995 4.5005
R12112 GNDA.n6530 GNDA.t997 4.5005
R12113 GNDA.n6531 GNDA.t937 4.5005
R12114 GNDA.n6532 GNDA.t972 4.5005
R12115 GNDA.n6536 GNDA.t964 4.5005
R12116 GNDA.n6535 GNDA.t1034 4.5005
R12117 GNDA.n6534 GNDA.t1089 4.5005
R12118 GNDA.n6533 GNDA.t1054 4.5005
R12119 GNDA.n6537 GNDA.t1058 4.5005
R12120 GNDA.n6538 GNDA.t1001 4.5005
R12121 GNDA.n6539 GNDA.t1033 4.5005
R12122 GNDA.n6543 GNDA.t1025 4.5005
R12123 GNDA.n6542 GNDA.t1094 4.5005
R12124 GNDA.n6541 GNDA.t936 4.5005
R12125 GNDA.n6540 GNDA.t902 4.5005
R12126 GNDA.n6544 GNDA.t1005 4.5005
R12127 GNDA.n6545 GNDA.t946 4.5005
R12128 GNDA.n6546 GNDA.t981 4.5005
R12129 GNDA.n6550 GNDA.t970 4.5005
R12130 GNDA.n6549 GNDA.t1043 4.5005
R12131 GNDA.n6548 GNDA.t1096 4.5005
R12132 GNDA.n6547 GNDA.t1064 4.5005
R12133 GNDA.n6551 GNDA.t1056 4.5005
R12134 GNDA.n6552 GNDA.t999 4.5005
R12135 GNDA.n6553 GNDA.t1032 4.5005
R12136 GNDA.n6557 GNDA.t1024 4.5005
R12137 GNDA.n6556 GNDA.t1093 4.5005
R12138 GNDA.n6555 GNDA.t935 4.5005
R12139 GNDA.n6554 GNDA.t901 4.5005
R12140 GNDA.n6558 GNDA.t904 4.5005
R12141 GNDA.n6559 GNDA.t1060 4.5005
R12142 GNDA.n6560 GNDA.t1092 4.5005
R12143 GNDA.n6564 GNDA.t1086 4.5005
R12144 GNDA.n6563 GNDA.t941 4.5005
R12145 GNDA.n6562 GNDA.t998 4.5005
R12146 GNDA.n6561 GNDA.t963 4.5005
R12147 GNDA.n6565 GNDA.t1068 4.5005
R12148 GNDA.n6566 GNDA.t1008 4.5005
R12149 GNDA.n6567 GNDA.t1040 4.5005
R12150 GNDA.n6571 GNDA.t1031 4.5005
R12151 GNDA.n6570 GNDA.t891 4.5005
R12152 GNDA.n6569 GNDA.t942 4.5005
R12153 GNDA.n6568 GNDA.t910 4.5005
R12154 GNDA.n6572 GNDA.t913 4.5005
R12155 GNDA.n6573 GNDA.t1070 4.5005
R12156 GNDA.n6574 GNDA.t887 4.5005
R12157 GNDA.n6578 GNDA.t1091 4.5005
R12158 GNDA.n6577 GNDA.t952 4.5005
R12159 GNDA.n6576 GNDA.t1004 4.5005
R12160 GNDA.n6575 GNDA.t969 4.5005
R12161 GNDA.n6579 GNDA.t973 4.5005
R12162 GNDA.n6580 GNDA.t915 4.5005
R12163 GNDA.n6581 GNDA.t951 4.5005
R12164 GNDA.n6585 GNDA.t938 4.5005
R12165 GNDA.n6584 GNDA.t1013 4.5005
R12166 GNDA.n6583 GNDA.t1069 4.5005
R12167 GNDA.n6582 GNDA.t1030 4.5005
R12168 GNDA.n6586 GNDA.t920 4.5005
R12169 GNDA.n6587 GNDA.t1078 4.5005
R12170 GNDA.n6588 GNDA.t894 4.5005
R12171 GNDA.n6592 GNDA.t886 4.5005
R12172 GNDA.n6591 GNDA.t957 4.5005
R12173 GNDA.n6590 GNDA.t1015 4.5005
R12174 GNDA.n6589 GNDA.t978 4.5005
R12175 GNDA.n6593 GNDA.t980 4.5005
R12176 GNDA.n6594 GNDA.t924 4.5005
R12177 GNDA.n6595 GNDA.t956 4.5005
R12178 GNDA.n6599 GNDA.t950 4.5005
R12179 GNDA.n6598 GNDA.t1018 4.5005
R12180 GNDA.n6597 GNDA.t1077 4.5005
R12181 GNDA.n6596 GNDA.t1039 4.5005
R12182 GNDA.n6600 GNDA.t1042 4.5005
R12183 GNDA.n6601 GNDA.t985 4.5005
R12184 GNDA.n6602 GNDA.t1017 4.5005
R12185 GNDA.n6606 GNDA.t1009 4.5005
R12186 GNDA.n6605 GNDA.t1082 4.5005
R12187 GNDA.n6604 GNDA.t922 4.5005
R12188 GNDA.n6603 GNDA.t885 4.5005
R12189 GNDA.n6614 GNDA.t945 4.5005
R12190 GNDA.n6613 GNDA.t889 4.5005
R12191 GNDA.n6612 GNDA.t1047 4.5005
R12192 GNDA.n6611 GNDA.t1080 4.5005
R12193 GNDA.n6610 GNDA.t1072 4.5005
R12194 GNDA.n6609 GNDA.t930 4.5005
R12195 GNDA.n6608 GNDA.t983 4.5005
R12196 GNDA.n6607 GNDA.t949 4.5005
R12197 GNDA.n347 GNDA.n303 4.26717
R12198 GNDA.n347 GNDA.n346 4.26717
R12199 GNDA.n346 GNDA.n345 4.26717
R12200 GNDA.n345 GNDA.n311 4.26717
R12201 GNDA.n339 GNDA.n311 4.26717
R12202 GNDA.n339 GNDA.n338 4.26717
R12203 GNDA.n338 GNDA.n337 4.26717
R12204 GNDA.n337 GNDA.n319 4.26717
R12205 GNDA.n331 GNDA.n319 4.26717
R12206 GNDA.n331 GNDA.n330 4.26717
R12207 GNDA.n330 GNDA.n329 4.26717
R12208 GNDA.n7137 GNDA.n135 4.26717
R12209 GNDA.n7131 GNDA.n135 4.26717
R12210 GNDA.n7131 GNDA.n7130 4.26717
R12211 GNDA.n7130 GNDA.n7129 4.26717
R12212 GNDA.n7129 GNDA.n7127 4.26717
R12213 GNDA.n7127 GNDA.n7124 4.26717
R12214 GNDA.n7124 GNDA.n7123 4.26717
R12215 GNDA.n7123 GNDA.n7120 4.26717
R12216 GNDA.n7120 GNDA.n7119 4.26717
R12217 GNDA.n7119 GNDA.n7116 4.26717
R12218 GNDA.n7116 GNDA.n7115 4.26717
R12219 GNDA.n1133 GNDA.n914 4.26717
R12220 GNDA.n1133 GNDA.n1103 4.26717
R12221 GNDA.n1127 GNDA.n1103 4.26717
R12222 GNDA.n1127 GNDA.n1126 4.26717
R12223 GNDA.n1126 GNDA.n1125 4.26717
R12224 GNDA.n1125 GNDA.n1110 4.26717
R12225 GNDA.n1119 GNDA.n1110 4.26717
R12226 GNDA.n1119 GNDA.n1118 4.26717
R12227 GNDA.n1118 GNDA.n589 4.26717
R12228 GNDA.n6209 GNDA.n589 4.26717
R12229 GNDA.n6209 GNDA.n587 4.26717
R12230 GNDA.n6673 GNDA.n6672 4.26717
R12231 GNDA.n6672 GNDA.n6633 4.26717
R12232 GNDA.n6667 GNDA.n6633 4.26717
R12233 GNDA.n6667 GNDA.n6666 4.26717
R12234 GNDA.n6666 GNDA.n6665 4.26717
R12235 GNDA.n6665 GNDA.n6641 4.26717
R12236 GNDA.n6659 GNDA.n6641 4.26717
R12237 GNDA.n6659 GNDA.n6658 4.26717
R12238 GNDA.n6658 GNDA.n6657 4.26717
R12239 GNDA.n6657 GNDA.n6652 4.26717
R12240 GNDA.n6652 GNDA.n6651 4.26717
R12241 GNDA.n872 GNDA.n669 4.26717
R12242 GNDA.n872 GNDA.n667 4.26717
R12243 GNDA.n878 GNDA.n667 4.26717
R12244 GNDA.n878 GNDA.n665 4.26717
R12245 GNDA.n884 GNDA.n665 4.26717
R12246 GNDA.n884 GNDA.n663 4.26717
R12247 GNDA.n890 GNDA.n663 4.26717
R12248 GNDA.n890 GNDA.n661 4.26717
R12249 GNDA.n896 GNDA.n661 4.26717
R12250 GNDA.n896 GNDA.n659 4.26717
R12251 GNDA.n901 GNDA.n659 4.26717
R12252 GNDA.n1193 GNDA.n1192 4.26717
R12253 GNDA.n1192 GNDA.n1167 4.26717
R12254 GNDA.n1187 GNDA.n1167 4.26717
R12255 GNDA.n1187 GNDA.n1186 4.26717
R12256 GNDA.n1186 GNDA.n1185 4.26717
R12257 GNDA.n1185 GNDA.n1173 4.26717
R12258 GNDA.n1179 GNDA.n1173 4.26717
R12259 GNDA.n1179 GNDA.n1178 4.26717
R12260 GNDA.n1178 GNDA.n573 4.26717
R12261 GNDA.n6219 GNDA.n573 4.26717
R12262 GNDA.n6219 GNDA.n569 4.26717
R12263 GNDA.n1831 GNDA.n1589 4.2505
R12264 GNDA.n4792 GNDA.n4791 4.2505
R12265 GNDA.t743 GNDA.t51 4.19522
R12266 GNDA.n4115 GNDA.n4110 4.0005
R12267 GNDA.n4095 GNDA.n4094 4.0005
R12268 GNDA.n6090 GNDA.n1349 4.0005
R12269 GNDA.n6757 GNDA.n303 3.93531
R12270 GNDA.n7138 GNDA.n7137 3.93531
R12271 GNDA.n1139 GNDA.n914 3.93531
R12272 GNDA.n6673 GNDA.n6627 3.93531
R12273 GNDA.n693 GNDA.n669 3.93531
R12274 GNDA.n1193 GNDA.n905 3.93531
R12275 GNDA.t34 GNDA.t65 3.93305
R12276 GNDA.n4779 GNDA.n1595 3.83383
R12277 GNDA.n1307 GNDA.n1241 3.7893
R12278 GNDA.n1329 GNDA.n1328 3.7893
R12279 GNDA.n1324 GNDA.n1242 3.7893
R12280 GNDA.n1323 GNDA.n1315 3.7893
R12281 GNDA.n1318 GNDA.n1317 3.7893
R12282 GNDA.n6249 GNDA.n549 3.7893
R12283 GNDA.n548 GNDA.n545 3.7893
R12284 GNDA.n6258 GNDA.n6257 3.7893
R12285 GNDA.n6194 GNDA.n596 3.7893
R12286 GNDA.n602 GNDA.n601 3.7893
R12287 GNDA.n6188 GNDA.n6187 3.7893
R12288 GNDA.n6106 GNDA.n603 3.7893
R12289 GNDA.n6112 GNDA.n6110 3.7893
R12290 GNDA.n6119 GNDA.n6118 3.7893
R12291 GNDA.n6127 GNDA.n623 3.7893
R12292 GNDA.n6126 GNDA.n621 3.7893
R12293 GNDA.n7109 GNDA.n166 3.7893
R12294 GNDA.n7106 GNDA.n7105 3.7893
R12295 GNDA.n201 GNDA.n168 3.7893
R12296 GNDA.n219 GNDA.n218 3.7893
R12297 GNDA.n216 GNDA.n215 3.7893
R12298 GNDA.n211 GNDA.n204 3.7893
R12299 GNDA.n208 GNDA.n207 3.7893
R12300 GNDA.n7047 GNDA.n188 3.7893
R12301 GNDA.n808 GNDA.n783 3.7893
R12302 GNDA.n807 GNDA.n804 3.7893
R12303 GNDA.n803 GNDA.n784 3.7893
R12304 GNDA.n800 GNDA.n799 3.7893
R12305 GNDA.n796 GNDA.n785 3.7893
R12306 GNDA.n789 GNDA.n786 3.7893
R12307 GNDA.n813 GNDA.n708 3.7893
R12308 GNDA.n814 GNDA.n707 3.7893
R12309 GNDA.n7038 GNDA.n7037 3.7893
R12310 GNDA.n7034 GNDA.n6928 3.7893
R12311 GNDA.n7033 GNDA.n6931 3.7893
R12312 GNDA.n7030 GNDA.n7029 3.7893
R12313 GNDA.n6956 GNDA.n6932 3.7893
R12314 GNDA.n6965 GNDA.n6964 3.7893
R12315 GNDA.n6968 GNDA.n6955 3.7893
R12316 GNDA.n6973 GNDA.n6969 3.7893
R12317 GNDA.n7317 GNDA.n7316 3.7893
R12318 GNDA.n7313 GNDA.n59 3.7893
R12319 GNDA.n7312 GNDA.n62 3.7893
R12320 GNDA.n7309 GNDA.n7308 3.7893
R12321 GNDA.n7235 GNDA.n63 3.7893
R12322 GNDA.n7244 GNDA.n7243 3.7893
R12323 GNDA.n7247 GNDA.n7234 3.7893
R12324 GNDA.n7252 GNDA.n7248 3.7893
R12325 GNDA.n6894 GNDA.n6783 3.7893
R12326 GNDA.n6891 GNDA.n6890 3.7893
R12327 GNDA.n6807 GNDA.n6784 3.7893
R12328 GNDA.n6812 GNDA.n6810 3.7893
R12329 GNDA.n6817 GNDA.n6813 3.7893
R12330 GNDA.n6824 GNDA.n6823 3.7893
R12331 GNDA.n6827 GNDA.n6806 3.7893
R12332 GNDA.n6832 GNDA.n6828 3.7893
R12333 GNDA.n1041 GNDA.n924 3.7893
R12334 GNDA.n1040 GNDA.n929 3.7893
R12335 GNDA.n1047 GNDA.n1046 3.7893
R12336 GNDA.n965 GNDA.n930 3.7893
R12337 GNDA.n967 GNDA.n966 3.7893
R12338 GNDA.n964 GNDA.n946 3.7893
R12339 GNDA.n982 GNDA.n980 3.7893
R12340 GNDA.n981 GNDA.n593 3.7893
R12341 GNDA.n7326 GNDA.n22 3.7893
R12342 GNDA.n7325 GNDA.n23 3.7893
R12343 GNDA.n33 GNDA.n32 3.7893
R12344 GNDA.n39 GNDA.n38 3.7893
R12345 GNDA.n35 GNDA.n34 3.7893
R12346 GNDA.n7160 GNDA.n1 3.7893
R12347 GNDA.n7165 GNDA.n7163 3.7893
R12348 GNDA.n7170 GNDA.n7166 3.7893
R12349 GNDA.n6250 GNDA 3.7381
R12350 GNDA.n6117 GNDA 3.7381
R12351 GNDA.n212 GNDA 3.7381
R12352 GNDA GNDA.n792 3.7381
R12353 GNDA.n6961 GNDA 3.7381
R12354 GNDA.n7240 GNDA 3.7381
R12355 GNDA.n6820 GNDA 3.7381
R12356 GNDA GNDA.n972 3.7381
R12357 GNDA GNDA.n7331 3.7381
R12358 GNDA.n4786 GNDA.n1590 3.65764
R12359 GNDA.n4787 GNDA.n4786 3.65764
R12360 GNDA.n4136 GNDA.n4131 3.65764
R12361 GNDA.n4136 GNDA.n4135 3.65764
R12362 GNDA.n3218 GNDA.n3217 3.50398
R12363 GNDA.n3289 GNDA.n3288 3.48371
R12364 GNDA.n5400 GNDA.n5234 3.48265
R12365 GNDA.n6353 GNDA.n6287 3.47871
R12366 GNDA.n412 GNDA.n362 3.47871
R12367 GNDA.n4774 GNDA.n4773 3.47821
R12368 GNDA.n5801 GNDA.n5800 3.47821
R12369 GNDA.n2791 GNDA.n2790 3.47821
R12370 GNDA.n6079 GNDA.n6078 3.47821
R12371 GNDA.n1515 GNDA.n1514 3.47821
R12372 GNDA.n3750 GNDA.n3749 3.47821
R12373 GNDA.n3387 GNDA.n3386 3.47821
R12374 GNDA.n5230 GNDA.n5229 3.47821
R12375 GNDA.n5327 GNDA.n5326 3.47821
R12376 GNDA.n5518 GNDA.n5517 3.47821
R12377 GNDA.n5660 GNDA.n5659 3.47821
R12378 GNDA.n5942 GNDA.n5941 3.47821
R12379 GNDA.n4923 GNDA.n4922 3.47821
R12380 GNDA.n4637 GNDA.n4636 3.47821
R12381 GNDA.n4448 GNDA.n4447 3.47821
R12382 GNDA.n4282 GNDA.n4281 3.47821
R12383 GNDA.n1741 GNDA.n1740 3.47821
R12384 GNDA.n3939 GNDA.n3938 3.47821
R12385 GNDA.n4076 GNDA.n4075 3.47821
R12386 GNDA.n3584 GNDA.n3583 3.47821
R12387 GNDA.n2649 GNDA.n2648 3.47821
R12388 GNDA.n2932 GNDA.n2931 3.47821
R12389 GNDA.n3073 GNDA.n3072 3.47821
R12390 GNDA.n3214 GNDA.n3213 3.47821
R12391 GNDA.n3287 GNDA.n1893 3.43627
R12392 GNDA.n1420 GNDA.t876 3.42907
R12393 GNDA.n1420 GNDA.t850 3.42907
R12394 GNDA.n4804 GNDA.t75 3.42907
R12395 GNDA.n4804 GNDA.t854 3.42907
R12396 GNDA.n1833 GNDA.t108 3.42907
R12397 GNDA.n1833 GNDA.t125 3.42907
R12398 GNDA.n3465 GNDA.t104 3.42907
R12399 GNDA.n3465 GNDA.t31 3.42907
R12400 GNDA.n4640 GNDA.n4639 3.4105
R12401 GNDA.n4771 GNDA.n4770 3.4105
R12402 GNDA.n4769 GNDA.n4768 3.4105
R12403 GNDA.n4767 GNDA.n4766 3.4105
R12404 GNDA.n4765 GNDA.n4642 3.4105
R12405 GNDA.n4761 GNDA.n4760 3.4105
R12406 GNDA.n4759 GNDA.n4758 3.4105
R12407 GNDA.n4757 GNDA.n4756 3.4105
R12408 GNDA.n4755 GNDA.n4644 3.4105
R12409 GNDA.n4751 GNDA.n4750 3.4105
R12410 GNDA.n4749 GNDA.n4748 3.4105
R12411 GNDA.n4747 GNDA.n4746 3.4105
R12412 GNDA.n4745 GNDA.n4646 3.4105
R12413 GNDA.n4741 GNDA.n4740 3.4105
R12414 GNDA.n4739 GNDA.n4738 3.4105
R12415 GNDA.n4737 GNDA.n4736 3.4105
R12416 GNDA.n4735 GNDA.n4648 3.4105
R12417 GNDA.n4731 GNDA.n4730 3.4105
R12418 GNDA.n4729 GNDA.n4728 3.4105
R12419 GNDA.n4727 GNDA.n4726 3.4105
R12420 GNDA.n4725 GNDA.n4650 3.4105
R12421 GNDA.n4721 GNDA.n4720 3.4105
R12422 GNDA.n4719 GNDA.n4718 3.4105
R12423 GNDA.n4717 GNDA.n4716 3.4105
R12424 GNDA.n4715 GNDA.n4652 3.4105
R12425 GNDA.n4711 GNDA.n4710 3.4105
R12426 GNDA.n4709 GNDA.n4708 3.4105
R12427 GNDA.n4707 GNDA.n4706 3.4105
R12428 GNDA.n4705 GNDA.n4654 3.4105
R12429 GNDA.n4701 GNDA.n4700 3.4105
R12430 GNDA.n4699 GNDA.n4698 3.4105
R12431 GNDA.n4697 GNDA.n4696 3.4105
R12432 GNDA.n4695 GNDA.n4656 3.4105
R12433 GNDA.n4691 GNDA.n4690 3.4105
R12434 GNDA.n4689 GNDA.n4688 3.4105
R12435 GNDA.n4687 GNDA.n4686 3.4105
R12436 GNDA.n4685 GNDA.n4658 3.4105
R12437 GNDA.n4681 GNDA.n4680 3.4105
R12438 GNDA.n4679 GNDA.n4678 3.4105
R12439 GNDA.n4677 GNDA.n4676 3.4105
R12440 GNDA.n4675 GNDA.n4660 3.4105
R12441 GNDA.n4671 GNDA.n4670 3.4105
R12442 GNDA.n4669 GNDA.n4668 3.4105
R12443 GNDA.n4667 GNDA.n4666 3.4105
R12444 GNDA.n4665 GNDA.n4662 3.4105
R12445 GNDA.n1598 GNDA.n1597 3.4105
R12446 GNDA.n4777 GNDA.n4776 3.4105
R12447 GNDA.n5663 GNDA.n5662 3.4105
R12448 GNDA.n5798 GNDA.n5797 3.4105
R12449 GNDA.n5796 GNDA.n5795 3.4105
R12450 GNDA.n5794 GNDA.n5793 3.4105
R12451 GNDA.n5792 GNDA.n5665 3.4105
R12452 GNDA.n5788 GNDA.n5787 3.4105
R12453 GNDA.n5786 GNDA.n5785 3.4105
R12454 GNDA.n5784 GNDA.n5783 3.4105
R12455 GNDA.n5782 GNDA.n5667 3.4105
R12456 GNDA.n5778 GNDA.n5777 3.4105
R12457 GNDA.n5776 GNDA.n5775 3.4105
R12458 GNDA.n5774 GNDA.n5773 3.4105
R12459 GNDA.n5772 GNDA.n5669 3.4105
R12460 GNDA.n5768 GNDA.n5767 3.4105
R12461 GNDA.n5766 GNDA.n5765 3.4105
R12462 GNDA.n5764 GNDA.n5763 3.4105
R12463 GNDA.n5762 GNDA.n5671 3.4105
R12464 GNDA.n5758 GNDA.n5757 3.4105
R12465 GNDA.n5756 GNDA.n5755 3.4105
R12466 GNDA.n5754 GNDA.n5753 3.4105
R12467 GNDA.n5752 GNDA.n5673 3.4105
R12468 GNDA.n5748 GNDA.n5747 3.4105
R12469 GNDA.n5746 GNDA.n5745 3.4105
R12470 GNDA.n5744 GNDA.n5743 3.4105
R12471 GNDA.n5742 GNDA.n5675 3.4105
R12472 GNDA.n5738 GNDA.n5737 3.4105
R12473 GNDA.n5736 GNDA.n5735 3.4105
R12474 GNDA.n5734 GNDA.n5733 3.4105
R12475 GNDA.n5732 GNDA.n5677 3.4105
R12476 GNDA.n5728 GNDA.n5727 3.4105
R12477 GNDA.n5726 GNDA.n5725 3.4105
R12478 GNDA.n5724 GNDA.n5723 3.4105
R12479 GNDA.n5722 GNDA.n5679 3.4105
R12480 GNDA.n5718 GNDA.n5717 3.4105
R12481 GNDA.n5716 GNDA.n5715 3.4105
R12482 GNDA.n5714 GNDA.n5713 3.4105
R12483 GNDA.n5712 GNDA.n5681 3.4105
R12484 GNDA.n5708 GNDA.n5707 3.4105
R12485 GNDA.n5706 GNDA.n5705 3.4105
R12486 GNDA.n5704 GNDA.n5703 3.4105
R12487 GNDA.n5702 GNDA.n5683 3.4105
R12488 GNDA.n5698 GNDA.n5697 3.4105
R12489 GNDA.n5696 GNDA.n5695 3.4105
R12490 GNDA.n5694 GNDA.n5693 3.4105
R12491 GNDA.n5692 GNDA.n5685 3.4105
R12492 GNDA.n5688 GNDA.n5687 3.4105
R12493 GNDA.n5686 GNDA.n4972 3.4105
R12494 GNDA.n2652 GNDA.n2651 3.4105
R12495 GNDA.n2788 GNDA.n2787 3.4105
R12496 GNDA.n2786 GNDA.n2785 3.4105
R12497 GNDA.n2784 GNDA.n2656 3.4105
R12498 GNDA.n2655 GNDA.n2654 3.4105
R12499 GNDA.n2780 GNDA.n2779 3.4105
R12500 GNDA.n2778 GNDA.n2777 3.4105
R12501 GNDA.n2776 GNDA.n2660 3.4105
R12502 GNDA.n2659 GNDA.n2658 3.4105
R12503 GNDA.n2772 GNDA.n2771 3.4105
R12504 GNDA.n2770 GNDA.n2769 3.4105
R12505 GNDA.n2768 GNDA.n2664 3.4105
R12506 GNDA.n2663 GNDA.n2662 3.4105
R12507 GNDA.n2764 GNDA.n2763 3.4105
R12508 GNDA.n2762 GNDA.n2761 3.4105
R12509 GNDA.n2760 GNDA.n2668 3.4105
R12510 GNDA.n2667 GNDA.n2666 3.4105
R12511 GNDA.n2756 GNDA.n2755 3.4105
R12512 GNDA.n2754 GNDA.n2753 3.4105
R12513 GNDA.n2752 GNDA.n2672 3.4105
R12514 GNDA.n2671 GNDA.n2670 3.4105
R12515 GNDA.n2748 GNDA.n2747 3.4105
R12516 GNDA.n2746 GNDA.n2745 3.4105
R12517 GNDA.n2744 GNDA.n2676 3.4105
R12518 GNDA.n2675 GNDA.n2674 3.4105
R12519 GNDA.n2740 GNDA.n2739 3.4105
R12520 GNDA.n2738 GNDA.n2737 3.4105
R12521 GNDA.n2736 GNDA.n2680 3.4105
R12522 GNDA.n2679 GNDA.n2678 3.4105
R12523 GNDA.n2732 GNDA.n2731 3.4105
R12524 GNDA.n2730 GNDA.n2729 3.4105
R12525 GNDA.n2728 GNDA.n2684 3.4105
R12526 GNDA.n2683 GNDA.n2682 3.4105
R12527 GNDA.n2724 GNDA.n2723 3.4105
R12528 GNDA.n2722 GNDA.n2721 3.4105
R12529 GNDA.n2720 GNDA.n2688 3.4105
R12530 GNDA.n2687 GNDA.n2686 3.4105
R12531 GNDA.n2716 GNDA.n2715 3.4105
R12532 GNDA.n2714 GNDA.n2713 3.4105
R12533 GNDA.n2712 GNDA.n2692 3.4105
R12534 GNDA.n2691 GNDA.n2690 3.4105
R12535 GNDA.n2708 GNDA.n2707 3.4105
R12536 GNDA.n2706 GNDA.n2705 3.4105
R12537 GNDA.n2704 GNDA.n2696 3.4105
R12538 GNDA.n2695 GNDA.n2694 3.4105
R12539 GNDA.n2700 GNDA.n2699 3.4105
R12540 GNDA.n2698 GNDA.n2462 3.4105
R12541 GNDA.n5945 GNDA.n5944 3.4105
R12542 GNDA.n6076 GNDA.n6075 3.4105
R12543 GNDA.n6074 GNDA.n6073 3.4105
R12544 GNDA.n6072 GNDA.n6071 3.4105
R12545 GNDA.n6070 GNDA.n5947 3.4105
R12546 GNDA.n6066 GNDA.n6065 3.4105
R12547 GNDA.n6064 GNDA.n6063 3.4105
R12548 GNDA.n6062 GNDA.n6061 3.4105
R12549 GNDA.n6060 GNDA.n5949 3.4105
R12550 GNDA.n6056 GNDA.n6055 3.4105
R12551 GNDA.n6054 GNDA.n6053 3.4105
R12552 GNDA.n6052 GNDA.n6051 3.4105
R12553 GNDA.n6050 GNDA.n5951 3.4105
R12554 GNDA.n6046 GNDA.n6045 3.4105
R12555 GNDA.n6044 GNDA.n6043 3.4105
R12556 GNDA.n6042 GNDA.n6041 3.4105
R12557 GNDA.n6040 GNDA.n5953 3.4105
R12558 GNDA.n6036 GNDA.n6035 3.4105
R12559 GNDA.n6034 GNDA.n6033 3.4105
R12560 GNDA.n6032 GNDA.n6031 3.4105
R12561 GNDA.n6030 GNDA.n5955 3.4105
R12562 GNDA.n6026 GNDA.n6025 3.4105
R12563 GNDA.n6024 GNDA.n6023 3.4105
R12564 GNDA.n6022 GNDA.n6021 3.4105
R12565 GNDA.n6020 GNDA.n5957 3.4105
R12566 GNDA.n6016 GNDA.n6015 3.4105
R12567 GNDA.n6014 GNDA.n6013 3.4105
R12568 GNDA.n6012 GNDA.n6011 3.4105
R12569 GNDA.n6010 GNDA.n5959 3.4105
R12570 GNDA.n6006 GNDA.n6005 3.4105
R12571 GNDA.n6004 GNDA.n6003 3.4105
R12572 GNDA.n6002 GNDA.n6001 3.4105
R12573 GNDA.n6000 GNDA.n5961 3.4105
R12574 GNDA.n5996 GNDA.n5995 3.4105
R12575 GNDA.n5994 GNDA.n5993 3.4105
R12576 GNDA.n5992 GNDA.n5991 3.4105
R12577 GNDA.n5990 GNDA.n5963 3.4105
R12578 GNDA.n5986 GNDA.n5985 3.4105
R12579 GNDA.n5984 GNDA.n5983 3.4105
R12580 GNDA.n5982 GNDA.n5981 3.4105
R12581 GNDA.n5980 GNDA.n5965 3.4105
R12582 GNDA.n5976 GNDA.n5975 3.4105
R12583 GNDA.n5974 GNDA.n5973 3.4105
R12584 GNDA.n5972 GNDA.n5971 3.4105
R12585 GNDA.n5970 GNDA.n5967 3.4105
R12586 GNDA.n1370 GNDA.n1369 3.4105
R12587 GNDA.n6082 GNDA.n6081 3.4105
R12588 GNDA.n1516 GNDA.n1469 3.4105
R12589 GNDA.n1518 GNDA.n1468 3.4105
R12590 GNDA.n1519 GNDA.n1467 3.4105
R12591 GNDA.n1521 GNDA.n1466 3.4105
R12592 GNDA.n1522 GNDA.n1465 3.4105
R12593 GNDA.n1524 GNDA.n1464 3.4105
R12594 GNDA.n1525 GNDA.n1463 3.4105
R12595 GNDA.n1527 GNDA.n1462 3.4105
R12596 GNDA.n1528 GNDA.n1461 3.4105
R12597 GNDA.n1530 GNDA.n1460 3.4105
R12598 GNDA.n1531 GNDA.n1459 3.4105
R12599 GNDA.n1533 GNDA.n1458 3.4105
R12600 GNDA.n1534 GNDA.n1457 3.4105
R12601 GNDA.n1536 GNDA.n1456 3.4105
R12602 GNDA.n1537 GNDA.n1455 3.4105
R12603 GNDA.n1539 GNDA.n1454 3.4105
R12604 GNDA.n1540 GNDA.n1453 3.4105
R12605 GNDA.n1542 GNDA.n1452 3.4105
R12606 GNDA.n1543 GNDA.n1451 3.4105
R12607 GNDA.n1545 GNDA.n1450 3.4105
R12608 GNDA.n1546 GNDA.n1449 3.4105
R12609 GNDA.n1548 GNDA.n1448 3.4105
R12610 GNDA.n1549 GNDA.n1447 3.4105
R12611 GNDA.n1551 GNDA.n1446 3.4105
R12612 GNDA.n1552 GNDA.n1445 3.4105
R12613 GNDA.n1554 GNDA.n1444 3.4105
R12614 GNDA.n1555 GNDA.n1443 3.4105
R12615 GNDA.n1557 GNDA.n1442 3.4105
R12616 GNDA.n1558 GNDA.n1441 3.4105
R12617 GNDA.n1560 GNDA.n1440 3.4105
R12618 GNDA.n1561 GNDA.n1439 3.4105
R12619 GNDA.n1563 GNDA.n1438 3.4105
R12620 GNDA.n1564 GNDA.n1437 3.4105
R12621 GNDA.n1566 GNDA.n1436 3.4105
R12622 GNDA.n1567 GNDA.n1435 3.4105
R12623 GNDA.n1569 GNDA.n1434 3.4105
R12624 GNDA.n1570 GNDA.n1433 3.4105
R12625 GNDA.n1572 GNDA.n1432 3.4105
R12626 GNDA.n1573 GNDA.n1431 3.4105
R12627 GNDA.n1575 GNDA.n1430 3.4105
R12628 GNDA.n1576 GNDA.n1429 3.4105
R12629 GNDA.n1578 GNDA.n1428 3.4105
R12630 GNDA.n1579 GNDA.n1427 3.4105
R12631 GNDA.n1581 GNDA.n1426 3.4105
R12632 GNDA.n1582 GNDA.n1425 3.4105
R12633 GNDA.n1584 GNDA.n1424 3.4105
R12634 GNDA.n1586 GNDA.n1585 3.4105
R12635 GNDA.n3611 GNDA.n3610 3.4105
R12636 GNDA.n3747 GNDA.n3746 3.4105
R12637 GNDA.n3745 GNDA.n3744 3.4105
R12638 GNDA.n3743 GNDA.n3742 3.4105
R12639 GNDA.n3741 GNDA.n3613 3.4105
R12640 GNDA.n3737 GNDA.n3736 3.4105
R12641 GNDA.n3735 GNDA.n3734 3.4105
R12642 GNDA.n3733 GNDA.n3732 3.4105
R12643 GNDA.n3731 GNDA.n3615 3.4105
R12644 GNDA.n3727 GNDA.n3726 3.4105
R12645 GNDA.n3725 GNDA.n3724 3.4105
R12646 GNDA.n3723 GNDA.n3722 3.4105
R12647 GNDA.n3721 GNDA.n3617 3.4105
R12648 GNDA.n3717 GNDA.n3716 3.4105
R12649 GNDA.n3715 GNDA.n3714 3.4105
R12650 GNDA.n3713 GNDA.n3712 3.4105
R12651 GNDA.n3711 GNDA.n3619 3.4105
R12652 GNDA.n3707 GNDA.n3706 3.4105
R12653 GNDA.n3705 GNDA.n3704 3.4105
R12654 GNDA.n3703 GNDA.n3702 3.4105
R12655 GNDA.n3701 GNDA.n3621 3.4105
R12656 GNDA.n3697 GNDA.n3696 3.4105
R12657 GNDA.n3695 GNDA.n3694 3.4105
R12658 GNDA.n3693 GNDA.n3692 3.4105
R12659 GNDA.n3691 GNDA.n3623 3.4105
R12660 GNDA.n3687 GNDA.n3686 3.4105
R12661 GNDA.n3685 GNDA.n3684 3.4105
R12662 GNDA.n3683 GNDA.n3682 3.4105
R12663 GNDA.n3681 GNDA.n3625 3.4105
R12664 GNDA.n3677 GNDA.n3676 3.4105
R12665 GNDA.n3675 GNDA.n3674 3.4105
R12666 GNDA.n3673 GNDA.n3672 3.4105
R12667 GNDA.n3671 GNDA.n3627 3.4105
R12668 GNDA.n3667 GNDA.n3666 3.4105
R12669 GNDA.n3665 GNDA.n3664 3.4105
R12670 GNDA.n3663 GNDA.n3662 3.4105
R12671 GNDA.n3661 GNDA.n3629 3.4105
R12672 GNDA.n3657 GNDA.n3656 3.4105
R12673 GNDA.n3655 GNDA.n3654 3.4105
R12674 GNDA.n3653 GNDA.n3652 3.4105
R12675 GNDA.n3651 GNDA.n3631 3.4105
R12676 GNDA.n3647 GNDA.n3646 3.4105
R12677 GNDA.n3645 GNDA.n3644 3.4105
R12678 GNDA.n3643 GNDA.n3642 3.4105
R12679 GNDA.n3641 GNDA.n3633 3.4105
R12680 GNDA.n3637 GNDA.n3636 3.4105
R12681 GNDA.n3635 GNDA.n3586 3.4105
R12682 GNDA.n3388 GNDA.n3341 3.4105
R12683 GNDA.n3390 GNDA.n3340 3.4105
R12684 GNDA.n3391 GNDA.n3339 3.4105
R12685 GNDA.n3393 GNDA.n3338 3.4105
R12686 GNDA.n3394 GNDA.n3337 3.4105
R12687 GNDA.n3396 GNDA.n3336 3.4105
R12688 GNDA.n3397 GNDA.n3335 3.4105
R12689 GNDA.n3399 GNDA.n3334 3.4105
R12690 GNDA.n3400 GNDA.n3333 3.4105
R12691 GNDA.n3402 GNDA.n3332 3.4105
R12692 GNDA.n3403 GNDA.n3331 3.4105
R12693 GNDA.n3405 GNDA.n3330 3.4105
R12694 GNDA.n3406 GNDA.n3329 3.4105
R12695 GNDA.n3408 GNDA.n3328 3.4105
R12696 GNDA.n3409 GNDA.n3327 3.4105
R12697 GNDA.n3411 GNDA.n3326 3.4105
R12698 GNDA.n3412 GNDA.n3325 3.4105
R12699 GNDA.n3414 GNDA.n3324 3.4105
R12700 GNDA.n3415 GNDA.n3323 3.4105
R12701 GNDA.n3417 GNDA.n3322 3.4105
R12702 GNDA.n3418 GNDA.n3321 3.4105
R12703 GNDA.n3420 GNDA.n3320 3.4105
R12704 GNDA.n3421 GNDA.n3319 3.4105
R12705 GNDA.n3423 GNDA.n3318 3.4105
R12706 GNDA.n3424 GNDA.n3317 3.4105
R12707 GNDA.n3426 GNDA.n3316 3.4105
R12708 GNDA.n3427 GNDA.n3315 3.4105
R12709 GNDA.n3429 GNDA.n3314 3.4105
R12710 GNDA.n3430 GNDA.n3313 3.4105
R12711 GNDA.n3432 GNDA.n3312 3.4105
R12712 GNDA.n3433 GNDA.n3311 3.4105
R12713 GNDA.n3435 GNDA.n3310 3.4105
R12714 GNDA.n3436 GNDA.n3309 3.4105
R12715 GNDA.n3438 GNDA.n3308 3.4105
R12716 GNDA.n3439 GNDA.n3307 3.4105
R12717 GNDA.n3441 GNDA.n3306 3.4105
R12718 GNDA.n3442 GNDA.n3305 3.4105
R12719 GNDA.n3444 GNDA.n3304 3.4105
R12720 GNDA.n3445 GNDA.n3303 3.4105
R12721 GNDA.n3447 GNDA.n3302 3.4105
R12722 GNDA.n3448 GNDA.n3301 3.4105
R12723 GNDA.n3450 GNDA.n3300 3.4105
R12724 GNDA.n3451 GNDA.n3299 3.4105
R12725 GNDA.n3453 GNDA.n3298 3.4105
R12726 GNDA.n3454 GNDA.n3297 3.4105
R12727 GNDA.n3456 GNDA.n3296 3.4105
R12728 GNDA.n3458 GNDA.n3457 3.4105
R12729 GNDA.n5096 GNDA.n5095 3.4105
R12730 GNDA.n5227 GNDA.n5226 3.4105
R12731 GNDA.n5225 GNDA.n5224 3.4105
R12732 GNDA.n5223 GNDA.n5222 3.4105
R12733 GNDA.n5221 GNDA.n5098 3.4105
R12734 GNDA.n5217 GNDA.n5216 3.4105
R12735 GNDA.n5215 GNDA.n5214 3.4105
R12736 GNDA.n5213 GNDA.n5212 3.4105
R12737 GNDA.n5211 GNDA.n5100 3.4105
R12738 GNDA.n5207 GNDA.n5206 3.4105
R12739 GNDA.n5205 GNDA.n5204 3.4105
R12740 GNDA.n5203 GNDA.n5202 3.4105
R12741 GNDA.n5201 GNDA.n5102 3.4105
R12742 GNDA.n5197 GNDA.n5196 3.4105
R12743 GNDA.n5195 GNDA.n5194 3.4105
R12744 GNDA.n5193 GNDA.n5192 3.4105
R12745 GNDA.n5191 GNDA.n5104 3.4105
R12746 GNDA.n5187 GNDA.n5186 3.4105
R12747 GNDA.n5185 GNDA.n5184 3.4105
R12748 GNDA.n5183 GNDA.n5182 3.4105
R12749 GNDA.n5181 GNDA.n5106 3.4105
R12750 GNDA.n5177 GNDA.n5176 3.4105
R12751 GNDA.n5175 GNDA.n5174 3.4105
R12752 GNDA.n5173 GNDA.n5172 3.4105
R12753 GNDA.n5171 GNDA.n5108 3.4105
R12754 GNDA.n5167 GNDA.n5166 3.4105
R12755 GNDA.n5165 GNDA.n5164 3.4105
R12756 GNDA.n5163 GNDA.n5162 3.4105
R12757 GNDA.n5161 GNDA.n5110 3.4105
R12758 GNDA.n5157 GNDA.n5156 3.4105
R12759 GNDA.n5155 GNDA.n5154 3.4105
R12760 GNDA.n5153 GNDA.n5152 3.4105
R12761 GNDA.n5151 GNDA.n5112 3.4105
R12762 GNDA.n5147 GNDA.n5146 3.4105
R12763 GNDA.n5145 GNDA.n5144 3.4105
R12764 GNDA.n5143 GNDA.n5142 3.4105
R12765 GNDA.n5141 GNDA.n5114 3.4105
R12766 GNDA.n5137 GNDA.n5136 3.4105
R12767 GNDA.n5135 GNDA.n5134 3.4105
R12768 GNDA.n5133 GNDA.n5132 3.4105
R12769 GNDA.n5131 GNDA.n5116 3.4105
R12770 GNDA.n5127 GNDA.n5126 3.4105
R12771 GNDA.n5125 GNDA.n5124 3.4105
R12772 GNDA.n5123 GNDA.n5122 3.4105
R12773 GNDA.n5121 GNDA.n5118 3.4105
R12774 GNDA.n5071 GNDA.n5070 3.4105
R12775 GNDA.n5233 GNDA.n5232 3.4105
R12776 GNDA.n5328 GNDA.n5281 3.4105
R12777 GNDA.n5330 GNDA.n5280 3.4105
R12778 GNDA.n5331 GNDA.n5279 3.4105
R12779 GNDA.n5333 GNDA.n5278 3.4105
R12780 GNDA.n5334 GNDA.n5277 3.4105
R12781 GNDA.n5336 GNDA.n5276 3.4105
R12782 GNDA.n5337 GNDA.n5275 3.4105
R12783 GNDA.n5339 GNDA.n5274 3.4105
R12784 GNDA.n5340 GNDA.n5273 3.4105
R12785 GNDA.n5342 GNDA.n5272 3.4105
R12786 GNDA.n5343 GNDA.n5271 3.4105
R12787 GNDA.n5345 GNDA.n5270 3.4105
R12788 GNDA.n5346 GNDA.n5269 3.4105
R12789 GNDA.n5348 GNDA.n5268 3.4105
R12790 GNDA.n5349 GNDA.n5267 3.4105
R12791 GNDA.n5351 GNDA.n5266 3.4105
R12792 GNDA.n5352 GNDA.n5265 3.4105
R12793 GNDA.n5354 GNDA.n5264 3.4105
R12794 GNDA.n5355 GNDA.n5263 3.4105
R12795 GNDA.n5357 GNDA.n5262 3.4105
R12796 GNDA.n5358 GNDA.n5261 3.4105
R12797 GNDA.n5360 GNDA.n5260 3.4105
R12798 GNDA.n5361 GNDA.n5259 3.4105
R12799 GNDA.n5363 GNDA.n5258 3.4105
R12800 GNDA.n5364 GNDA.n5257 3.4105
R12801 GNDA.n5366 GNDA.n5256 3.4105
R12802 GNDA.n5367 GNDA.n5255 3.4105
R12803 GNDA.n5369 GNDA.n5254 3.4105
R12804 GNDA.n5370 GNDA.n5253 3.4105
R12805 GNDA.n5372 GNDA.n5252 3.4105
R12806 GNDA.n5373 GNDA.n5251 3.4105
R12807 GNDA.n5375 GNDA.n5250 3.4105
R12808 GNDA.n5376 GNDA.n5249 3.4105
R12809 GNDA.n5378 GNDA.n5248 3.4105
R12810 GNDA.n5379 GNDA.n5247 3.4105
R12811 GNDA.n5381 GNDA.n5246 3.4105
R12812 GNDA.n5382 GNDA.n5245 3.4105
R12813 GNDA.n5384 GNDA.n5244 3.4105
R12814 GNDA.n5385 GNDA.n5243 3.4105
R12815 GNDA.n5387 GNDA.n5242 3.4105
R12816 GNDA.n5388 GNDA.n5241 3.4105
R12817 GNDA.n5390 GNDA.n5240 3.4105
R12818 GNDA.n5391 GNDA.n5239 3.4105
R12819 GNDA.n5393 GNDA.n5238 3.4105
R12820 GNDA.n5394 GNDA.n5237 3.4105
R12821 GNDA.n5396 GNDA.n5236 3.4105
R12822 GNDA.n5398 GNDA.n5397 3.4105
R12823 GNDA.n5046 GNDA.n5045 3.4105
R12824 GNDA.n5515 GNDA.n5514 3.4105
R12825 GNDA.n5513 GNDA.n5512 3.4105
R12826 GNDA.n5511 GNDA.n5510 3.4105
R12827 GNDA.n5509 GNDA.n5048 3.4105
R12828 GNDA.n5505 GNDA.n5504 3.4105
R12829 GNDA.n5503 GNDA.n5502 3.4105
R12830 GNDA.n5501 GNDA.n5500 3.4105
R12831 GNDA.n5499 GNDA.n5050 3.4105
R12832 GNDA.n5495 GNDA.n5494 3.4105
R12833 GNDA.n5493 GNDA.n5492 3.4105
R12834 GNDA.n5491 GNDA.n5490 3.4105
R12835 GNDA.n5489 GNDA.n5052 3.4105
R12836 GNDA.n5485 GNDA.n5484 3.4105
R12837 GNDA.n5483 GNDA.n5482 3.4105
R12838 GNDA.n5481 GNDA.n5480 3.4105
R12839 GNDA.n5479 GNDA.n5054 3.4105
R12840 GNDA.n5475 GNDA.n5474 3.4105
R12841 GNDA.n5473 GNDA.n5472 3.4105
R12842 GNDA.n5471 GNDA.n5470 3.4105
R12843 GNDA.n5469 GNDA.n5056 3.4105
R12844 GNDA.n5465 GNDA.n5464 3.4105
R12845 GNDA.n5463 GNDA.n5462 3.4105
R12846 GNDA.n5461 GNDA.n5460 3.4105
R12847 GNDA.n5459 GNDA.n5058 3.4105
R12848 GNDA.n5455 GNDA.n5454 3.4105
R12849 GNDA.n5453 GNDA.n5452 3.4105
R12850 GNDA.n5451 GNDA.n5450 3.4105
R12851 GNDA.n5449 GNDA.n5060 3.4105
R12852 GNDA.n5445 GNDA.n5444 3.4105
R12853 GNDA.n5443 GNDA.n5442 3.4105
R12854 GNDA.n5441 GNDA.n5440 3.4105
R12855 GNDA.n5439 GNDA.n5062 3.4105
R12856 GNDA.n5435 GNDA.n5434 3.4105
R12857 GNDA.n5433 GNDA.n5432 3.4105
R12858 GNDA.n5431 GNDA.n5430 3.4105
R12859 GNDA.n5429 GNDA.n5064 3.4105
R12860 GNDA.n5425 GNDA.n5424 3.4105
R12861 GNDA.n5423 GNDA.n5422 3.4105
R12862 GNDA.n5421 GNDA.n5420 3.4105
R12863 GNDA.n5419 GNDA.n5066 3.4105
R12864 GNDA.n5415 GNDA.n5414 3.4105
R12865 GNDA.n5413 GNDA.n5412 3.4105
R12866 GNDA.n5411 GNDA.n5410 3.4105
R12867 GNDA.n5409 GNDA.n5068 3.4105
R12868 GNDA.n5405 GNDA.n5404 3.4105
R12869 GNDA.n5403 GNDA.n5020 3.4105
R12870 GNDA.n5521 GNDA.n5520 3.4105
R12871 GNDA.n5657 GNDA.n5656 3.4105
R12872 GNDA.n5655 GNDA.n5654 3.4105
R12873 GNDA.n5653 GNDA.n5652 3.4105
R12874 GNDA.n5651 GNDA.n5523 3.4105
R12875 GNDA.n5647 GNDA.n5646 3.4105
R12876 GNDA.n5645 GNDA.n5644 3.4105
R12877 GNDA.n5643 GNDA.n5642 3.4105
R12878 GNDA.n5641 GNDA.n5525 3.4105
R12879 GNDA.n5637 GNDA.n5636 3.4105
R12880 GNDA.n5635 GNDA.n5634 3.4105
R12881 GNDA.n5633 GNDA.n5632 3.4105
R12882 GNDA.n5631 GNDA.n5527 3.4105
R12883 GNDA.n5627 GNDA.n5626 3.4105
R12884 GNDA.n5625 GNDA.n5624 3.4105
R12885 GNDA.n5623 GNDA.n5622 3.4105
R12886 GNDA.n5621 GNDA.n5529 3.4105
R12887 GNDA.n5617 GNDA.n5616 3.4105
R12888 GNDA.n5615 GNDA.n5614 3.4105
R12889 GNDA.n5613 GNDA.n5612 3.4105
R12890 GNDA.n5611 GNDA.n5531 3.4105
R12891 GNDA.n5607 GNDA.n5606 3.4105
R12892 GNDA.n5605 GNDA.n5604 3.4105
R12893 GNDA.n5603 GNDA.n5602 3.4105
R12894 GNDA.n5601 GNDA.n5533 3.4105
R12895 GNDA.n5597 GNDA.n5596 3.4105
R12896 GNDA.n5595 GNDA.n5594 3.4105
R12897 GNDA.n5593 GNDA.n5592 3.4105
R12898 GNDA.n5591 GNDA.n5535 3.4105
R12899 GNDA.n5587 GNDA.n5586 3.4105
R12900 GNDA.n5585 GNDA.n5584 3.4105
R12901 GNDA.n5583 GNDA.n5582 3.4105
R12902 GNDA.n5581 GNDA.n5537 3.4105
R12903 GNDA.n5577 GNDA.n5576 3.4105
R12904 GNDA.n5575 GNDA.n5574 3.4105
R12905 GNDA.n5573 GNDA.n5572 3.4105
R12906 GNDA.n5571 GNDA.n5539 3.4105
R12907 GNDA.n5567 GNDA.n5566 3.4105
R12908 GNDA.n5565 GNDA.n5564 3.4105
R12909 GNDA.n5563 GNDA.n5562 3.4105
R12910 GNDA.n5561 GNDA.n5541 3.4105
R12911 GNDA.n5557 GNDA.n5556 3.4105
R12912 GNDA.n5555 GNDA.n5554 3.4105
R12913 GNDA.n5553 GNDA.n5552 3.4105
R12914 GNDA.n5551 GNDA.n5543 3.4105
R12915 GNDA.n5547 GNDA.n5546 3.4105
R12916 GNDA.n5545 GNDA.n4996 3.4105
R12917 GNDA.n5804 GNDA.n5803 3.4105
R12918 GNDA.n5939 GNDA.n5938 3.4105
R12919 GNDA.n5937 GNDA.n5936 3.4105
R12920 GNDA.n5935 GNDA.n5934 3.4105
R12921 GNDA.n5933 GNDA.n5806 3.4105
R12922 GNDA.n5929 GNDA.n5928 3.4105
R12923 GNDA.n5927 GNDA.n5926 3.4105
R12924 GNDA.n5925 GNDA.n5924 3.4105
R12925 GNDA.n5923 GNDA.n5808 3.4105
R12926 GNDA.n5919 GNDA.n5918 3.4105
R12927 GNDA.n5917 GNDA.n5916 3.4105
R12928 GNDA.n5915 GNDA.n5914 3.4105
R12929 GNDA.n5913 GNDA.n5810 3.4105
R12930 GNDA.n5909 GNDA.n5908 3.4105
R12931 GNDA.n5907 GNDA.n5906 3.4105
R12932 GNDA.n5905 GNDA.n5904 3.4105
R12933 GNDA.n5903 GNDA.n5812 3.4105
R12934 GNDA.n5899 GNDA.n5898 3.4105
R12935 GNDA.n5897 GNDA.n5896 3.4105
R12936 GNDA.n5895 GNDA.n5894 3.4105
R12937 GNDA.n5893 GNDA.n5814 3.4105
R12938 GNDA.n5889 GNDA.n5888 3.4105
R12939 GNDA.n5887 GNDA.n5886 3.4105
R12940 GNDA.n5885 GNDA.n5884 3.4105
R12941 GNDA.n5883 GNDA.n5816 3.4105
R12942 GNDA.n5879 GNDA.n5878 3.4105
R12943 GNDA.n5877 GNDA.n5876 3.4105
R12944 GNDA.n5875 GNDA.n5874 3.4105
R12945 GNDA.n5873 GNDA.n5818 3.4105
R12946 GNDA.n5869 GNDA.n5868 3.4105
R12947 GNDA.n5867 GNDA.n5866 3.4105
R12948 GNDA.n5865 GNDA.n5864 3.4105
R12949 GNDA.n5863 GNDA.n5820 3.4105
R12950 GNDA.n5859 GNDA.n5858 3.4105
R12951 GNDA.n5857 GNDA.n5856 3.4105
R12952 GNDA.n5855 GNDA.n5854 3.4105
R12953 GNDA.n5853 GNDA.n5822 3.4105
R12954 GNDA.n5849 GNDA.n5848 3.4105
R12955 GNDA.n5847 GNDA.n5846 3.4105
R12956 GNDA.n5845 GNDA.n5844 3.4105
R12957 GNDA.n5843 GNDA.n5824 3.4105
R12958 GNDA.n5839 GNDA.n5838 3.4105
R12959 GNDA.n5837 GNDA.n5836 3.4105
R12960 GNDA.n5835 GNDA.n5834 3.4105
R12961 GNDA.n5833 GNDA.n5826 3.4105
R12962 GNDA.n5829 GNDA.n5828 3.4105
R12963 GNDA.n5827 GNDA.n4948 3.4105
R12964 GNDA.n1397 GNDA.n1396 3.4105
R12965 GNDA.n4920 GNDA.n4919 3.4105
R12966 GNDA.n4918 GNDA.n4917 3.4105
R12967 GNDA.n4916 GNDA.n4915 3.4105
R12968 GNDA.n4914 GNDA.n1399 3.4105
R12969 GNDA.n4910 GNDA.n4909 3.4105
R12970 GNDA.n4908 GNDA.n4907 3.4105
R12971 GNDA.n4906 GNDA.n4905 3.4105
R12972 GNDA.n4904 GNDA.n1401 3.4105
R12973 GNDA.n4900 GNDA.n4899 3.4105
R12974 GNDA.n4898 GNDA.n4897 3.4105
R12975 GNDA.n4896 GNDA.n4895 3.4105
R12976 GNDA.n4894 GNDA.n1403 3.4105
R12977 GNDA.n4890 GNDA.n4889 3.4105
R12978 GNDA.n4888 GNDA.n4887 3.4105
R12979 GNDA.n4886 GNDA.n4885 3.4105
R12980 GNDA.n4884 GNDA.n1405 3.4105
R12981 GNDA.n4880 GNDA.n4879 3.4105
R12982 GNDA.n4878 GNDA.n4877 3.4105
R12983 GNDA.n4876 GNDA.n4875 3.4105
R12984 GNDA.n4874 GNDA.n1407 3.4105
R12985 GNDA.n4870 GNDA.n4869 3.4105
R12986 GNDA.n4868 GNDA.n4867 3.4105
R12987 GNDA.n4866 GNDA.n4865 3.4105
R12988 GNDA.n4864 GNDA.n1409 3.4105
R12989 GNDA.n4860 GNDA.n4859 3.4105
R12990 GNDA.n4858 GNDA.n4857 3.4105
R12991 GNDA.n4856 GNDA.n4855 3.4105
R12992 GNDA.n4854 GNDA.n1411 3.4105
R12993 GNDA.n4850 GNDA.n4849 3.4105
R12994 GNDA.n4848 GNDA.n4847 3.4105
R12995 GNDA.n4846 GNDA.n4845 3.4105
R12996 GNDA.n4844 GNDA.n1413 3.4105
R12997 GNDA.n4840 GNDA.n4839 3.4105
R12998 GNDA.n4838 GNDA.n4837 3.4105
R12999 GNDA.n4836 GNDA.n4835 3.4105
R13000 GNDA.n4834 GNDA.n1415 3.4105
R13001 GNDA.n4830 GNDA.n4829 3.4105
R13002 GNDA.n4828 GNDA.n4827 3.4105
R13003 GNDA.n4826 GNDA.n4825 3.4105
R13004 GNDA.n4824 GNDA.n1417 3.4105
R13005 GNDA.n4820 GNDA.n4819 3.4105
R13006 GNDA.n4818 GNDA.n4817 3.4105
R13007 GNDA.n4816 GNDA.n4815 3.4105
R13008 GNDA.n4814 GNDA.n1419 3.4105
R13009 GNDA.n4810 GNDA.n4809 3.4105
R13010 GNDA.n4808 GNDA.n1372 3.4105
R13011 GNDA.n4498 GNDA.n4497 3.4105
R13012 GNDA.n4634 GNDA.n4633 3.4105
R13013 GNDA.n4632 GNDA.n4631 3.4105
R13014 GNDA.n4630 GNDA.n4629 3.4105
R13015 GNDA.n4628 GNDA.n4500 3.4105
R13016 GNDA.n4624 GNDA.n4623 3.4105
R13017 GNDA.n4622 GNDA.n4621 3.4105
R13018 GNDA.n4620 GNDA.n4619 3.4105
R13019 GNDA.n4618 GNDA.n4502 3.4105
R13020 GNDA.n4614 GNDA.n4613 3.4105
R13021 GNDA.n4612 GNDA.n4611 3.4105
R13022 GNDA.n4610 GNDA.n4609 3.4105
R13023 GNDA.n4608 GNDA.n4504 3.4105
R13024 GNDA.n4604 GNDA.n4603 3.4105
R13025 GNDA.n4602 GNDA.n4601 3.4105
R13026 GNDA.n4600 GNDA.n4599 3.4105
R13027 GNDA.n4598 GNDA.n4506 3.4105
R13028 GNDA.n4594 GNDA.n4593 3.4105
R13029 GNDA.n4592 GNDA.n4591 3.4105
R13030 GNDA.n4590 GNDA.n4589 3.4105
R13031 GNDA.n4588 GNDA.n4508 3.4105
R13032 GNDA.n4584 GNDA.n4583 3.4105
R13033 GNDA.n4582 GNDA.n4581 3.4105
R13034 GNDA.n4580 GNDA.n4579 3.4105
R13035 GNDA.n4578 GNDA.n4510 3.4105
R13036 GNDA.n4574 GNDA.n4573 3.4105
R13037 GNDA.n4572 GNDA.n4571 3.4105
R13038 GNDA.n4570 GNDA.n4569 3.4105
R13039 GNDA.n4568 GNDA.n4512 3.4105
R13040 GNDA.n4564 GNDA.n4563 3.4105
R13041 GNDA.n4562 GNDA.n4561 3.4105
R13042 GNDA.n4560 GNDA.n4559 3.4105
R13043 GNDA.n4558 GNDA.n4514 3.4105
R13044 GNDA.n4554 GNDA.n4553 3.4105
R13045 GNDA.n4552 GNDA.n4551 3.4105
R13046 GNDA.n4550 GNDA.n4549 3.4105
R13047 GNDA.n4548 GNDA.n4516 3.4105
R13048 GNDA.n4544 GNDA.n4543 3.4105
R13049 GNDA.n4542 GNDA.n4541 3.4105
R13050 GNDA.n4540 GNDA.n4539 3.4105
R13051 GNDA.n4538 GNDA.n4518 3.4105
R13052 GNDA.n4534 GNDA.n4533 3.4105
R13053 GNDA.n4532 GNDA.n4531 3.4105
R13054 GNDA.n4530 GNDA.n4529 3.4105
R13055 GNDA.n4528 GNDA.n4520 3.4105
R13056 GNDA.n4524 GNDA.n4523 3.4105
R13057 GNDA.n4522 GNDA.n4473 3.4105
R13058 GNDA.n4309 GNDA.n4308 3.4105
R13059 GNDA.n4445 GNDA.n4444 3.4105
R13060 GNDA.n4443 GNDA.n4442 3.4105
R13061 GNDA.n4441 GNDA.n4440 3.4105
R13062 GNDA.n4439 GNDA.n4311 3.4105
R13063 GNDA.n4435 GNDA.n4434 3.4105
R13064 GNDA.n4433 GNDA.n4432 3.4105
R13065 GNDA.n4431 GNDA.n4430 3.4105
R13066 GNDA.n4429 GNDA.n4313 3.4105
R13067 GNDA.n4425 GNDA.n4424 3.4105
R13068 GNDA.n4423 GNDA.n4422 3.4105
R13069 GNDA.n4421 GNDA.n4420 3.4105
R13070 GNDA.n4419 GNDA.n4315 3.4105
R13071 GNDA.n4415 GNDA.n4414 3.4105
R13072 GNDA.n4413 GNDA.n4412 3.4105
R13073 GNDA.n4411 GNDA.n4410 3.4105
R13074 GNDA.n4409 GNDA.n4317 3.4105
R13075 GNDA.n4405 GNDA.n4404 3.4105
R13076 GNDA.n4403 GNDA.n4402 3.4105
R13077 GNDA.n4401 GNDA.n4400 3.4105
R13078 GNDA.n4399 GNDA.n4319 3.4105
R13079 GNDA.n4395 GNDA.n4394 3.4105
R13080 GNDA.n4393 GNDA.n4392 3.4105
R13081 GNDA.n4391 GNDA.n4390 3.4105
R13082 GNDA.n4389 GNDA.n4321 3.4105
R13083 GNDA.n4385 GNDA.n4384 3.4105
R13084 GNDA.n4383 GNDA.n4382 3.4105
R13085 GNDA.n4381 GNDA.n4380 3.4105
R13086 GNDA.n4379 GNDA.n4323 3.4105
R13087 GNDA.n4375 GNDA.n4374 3.4105
R13088 GNDA.n4373 GNDA.n4372 3.4105
R13089 GNDA.n4371 GNDA.n4370 3.4105
R13090 GNDA.n4369 GNDA.n4325 3.4105
R13091 GNDA.n4365 GNDA.n4364 3.4105
R13092 GNDA.n4363 GNDA.n4362 3.4105
R13093 GNDA.n4361 GNDA.n4360 3.4105
R13094 GNDA.n4359 GNDA.n4327 3.4105
R13095 GNDA.n4355 GNDA.n4354 3.4105
R13096 GNDA.n4353 GNDA.n4352 3.4105
R13097 GNDA.n4351 GNDA.n4350 3.4105
R13098 GNDA.n4349 GNDA.n4329 3.4105
R13099 GNDA.n4345 GNDA.n4344 3.4105
R13100 GNDA.n4343 GNDA.n4342 3.4105
R13101 GNDA.n4341 GNDA.n4340 3.4105
R13102 GNDA.n4339 GNDA.n4331 3.4105
R13103 GNDA.n4335 GNDA.n4334 3.4105
R13104 GNDA.n4333 GNDA.n4284 3.4105
R13105 GNDA.n1625 GNDA.n1624 3.4105
R13106 GNDA.n4279 GNDA.n4278 3.4105
R13107 GNDA.n4277 GNDA.n4276 3.4105
R13108 GNDA.n4275 GNDA.n4274 3.4105
R13109 GNDA.n4273 GNDA.n1627 3.4105
R13110 GNDA.n4269 GNDA.n4268 3.4105
R13111 GNDA.n4267 GNDA.n4266 3.4105
R13112 GNDA.n4265 GNDA.n4264 3.4105
R13113 GNDA.n4263 GNDA.n1629 3.4105
R13114 GNDA.n4259 GNDA.n4258 3.4105
R13115 GNDA.n4257 GNDA.n4256 3.4105
R13116 GNDA.n4255 GNDA.n4254 3.4105
R13117 GNDA.n4253 GNDA.n1631 3.4105
R13118 GNDA.n4249 GNDA.n4248 3.4105
R13119 GNDA.n4247 GNDA.n4246 3.4105
R13120 GNDA.n4245 GNDA.n4244 3.4105
R13121 GNDA.n4243 GNDA.n1633 3.4105
R13122 GNDA.n4239 GNDA.n4238 3.4105
R13123 GNDA.n4237 GNDA.n4236 3.4105
R13124 GNDA.n4235 GNDA.n4234 3.4105
R13125 GNDA.n4233 GNDA.n1635 3.4105
R13126 GNDA.n4229 GNDA.n4228 3.4105
R13127 GNDA.n4227 GNDA.n4226 3.4105
R13128 GNDA.n4225 GNDA.n4224 3.4105
R13129 GNDA.n4223 GNDA.n1637 3.4105
R13130 GNDA.n4219 GNDA.n4218 3.4105
R13131 GNDA.n4217 GNDA.n4216 3.4105
R13132 GNDA.n4215 GNDA.n4214 3.4105
R13133 GNDA.n4213 GNDA.n1639 3.4105
R13134 GNDA.n4209 GNDA.n4208 3.4105
R13135 GNDA.n4207 GNDA.n4206 3.4105
R13136 GNDA.n4205 GNDA.n4204 3.4105
R13137 GNDA.n4203 GNDA.n1641 3.4105
R13138 GNDA.n4199 GNDA.n4198 3.4105
R13139 GNDA.n4197 GNDA.n4196 3.4105
R13140 GNDA.n4195 GNDA.n4194 3.4105
R13141 GNDA.n4193 GNDA.n1643 3.4105
R13142 GNDA.n4189 GNDA.n4188 3.4105
R13143 GNDA.n4187 GNDA.n4186 3.4105
R13144 GNDA.n4185 GNDA.n4184 3.4105
R13145 GNDA.n4183 GNDA.n1645 3.4105
R13146 GNDA.n4179 GNDA.n4178 3.4105
R13147 GNDA.n4177 GNDA.n4176 3.4105
R13148 GNDA.n4175 GNDA.n4174 3.4105
R13149 GNDA.n4173 GNDA.n1647 3.4105
R13150 GNDA.n4169 GNDA.n4168 3.4105
R13151 GNDA.n4167 GNDA.n1600 3.4105
R13152 GNDA.n1742 GNDA.n1695 3.4105
R13153 GNDA.n1744 GNDA.n1694 3.4105
R13154 GNDA.n1745 GNDA.n1693 3.4105
R13155 GNDA.n1747 GNDA.n1692 3.4105
R13156 GNDA.n1748 GNDA.n1691 3.4105
R13157 GNDA.n1750 GNDA.n1690 3.4105
R13158 GNDA.n1751 GNDA.n1689 3.4105
R13159 GNDA.n1753 GNDA.n1688 3.4105
R13160 GNDA.n1754 GNDA.n1687 3.4105
R13161 GNDA.n1756 GNDA.n1686 3.4105
R13162 GNDA.n1757 GNDA.n1685 3.4105
R13163 GNDA.n1759 GNDA.n1684 3.4105
R13164 GNDA.n1760 GNDA.n1683 3.4105
R13165 GNDA.n1762 GNDA.n1682 3.4105
R13166 GNDA.n1763 GNDA.n1681 3.4105
R13167 GNDA.n1765 GNDA.n1680 3.4105
R13168 GNDA.n1766 GNDA.n1679 3.4105
R13169 GNDA.n1768 GNDA.n1678 3.4105
R13170 GNDA.n1769 GNDA.n1677 3.4105
R13171 GNDA.n1771 GNDA.n1676 3.4105
R13172 GNDA.n1772 GNDA.n1675 3.4105
R13173 GNDA.n1774 GNDA.n1674 3.4105
R13174 GNDA.n1775 GNDA.n1673 3.4105
R13175 GNDA.n1777 GNDA.n1672 3.4105
R13176 GNDA.n1778 GNDA.n1671 3.4105
R13177 GNDA.n1780 GNDA.n1670 3.4105
R13178 GNDA.n1781 GNDA.n1669 3.4105
R13179 GNDA.n1783 GNDA.n1668 3.4105
R13180 GNDA.n1784 GNDA.n1667 3.4105
R13181 GNDA.n1786 GNDA.n1666 3.4105
R13182 GNDA.n1787 GNDA.n1665 3.4105
R13183 GNDA.n1789 GNDA.n1664 3.4105
R13184 GNDA.n1790 GNDA.n1663 3.4105
R13185 GNDA.n1792 GNDA.n1662 3.4105
R13186 GNDA.n1793 GNDA.n1661 3.4105
R13187 GNDA.n1795 GNDA.n1660 3.4105
R13188 GNDA.n1796 GNDA.n1659 3.4105
R13189 GNDA.n1798 GNDA.n1658 3.4105
R13190 GNDA.n1799 GNDA.n1657 3.4105
R13191 GNDA.n1801 GNDA.n1656 3.4105
R13192 GNDA.n1802 GNDA.n1655 3.4105
R13193 GNDA.n1804 GNDA.n1654 3.4105
R13194 GNDA.n1805 GNDA.n1653 3.4105
R13195 GNDA.n1807 GNDA.n1652 3.4105
R13196 GNDA.n1808 GNDA.n1651 3.4105
R13197 GNDA.n1810 GNDA.n1650 3.4105
R13198 GNDA.n1812 GNDA.n1811 3.4105
R13199 GNDA.n3800 GNDA.n3799 3.4105
R13200 GNDA.n3936 GNDA.n3935 3.4105
R13201 GNDA.n3934 GNDA.n3933 3.4105
R13202 GNDA.n3932 GNDA.n3931 3.4105
R13203 GNDA.n3930 GNDA.n3802 3.4105
R13204 GNDA.n3926 GNDA.n3925 3.4105
R13205 GNDA.n3924 GNDA.n3923 3.4105
R13206 GNDA.n3922 GNDA.n3921 3.4105
R13207 GNDA.n3920 GNDA.n3804 3.4105
R13208 GNDA.n3916 GNDA.n3915 3.4105
R13209 GNDA.n3914 GNDA.n3913 3.4105
R13210 GNDA.n3912 GNDA.n3911 3.4105
R13211 GNDA.n3910 GNDA.n3806 3.4105
R13212 GNDA.n3906 GNDA.n3905 3.4105
R13213 GNDA.n3904 GNDA.n3903 3.4105
R13214 GNDA.n3902 GNDA.n3901 3.4105
R13215 GNDA.n3900 GNDA.n3808 3.4105
R13216 GNDA.n3896 GNDA.n3895 3.4105
R13217 GNDA.n3894 GNDA.n3893 3.4105
R13218 GNDA.n3892 GNDA.n3891 3.4105
R13219 GNDA.n3890 GNDA.n3810 3.4105
R13220 GNDA.n3886 GNDA.n3885 3.4105
R13221 GNDA.n3884 GNDA.n3883 3.4105
R13222 GNDA.n3882 GNDA.n3881 3.4105
R13223 GNDA.n3880 GNDA.n3812 3.4105
R13224 GNDA.n3876 GNDA.n3875 3.4105
R13225 GNDA.n3874 GNDA.n3873 3.4105
R13226 GNDA.n3872 GNDA.n3871 3.4105
R13227 GNDA.n3870 GNDA.n3814 3.4105
R13228 GNDA.n3866 GNDA.n3865 3.4105
R13229 GNDA.n3864 GNDA.n3863 3.4105
R13230 GNDA.n3862 GNDA.n3861 3.4105
R13231 GNDA.n3860 GNDA.n3816 3.4105
R13232 GNDA.n3856 GNDA.n3855 3.4105
R13233 GNDA.n3854 GNDA.n3853 3.4105
R13234 GNDA.n3852 GNDA.n3851 3.4105
R13235 GNDA.n3850 GNDA.n3818 3.4105
R13236 GNDA.n3846 GNDA.n3845 3.4105
R13237 GNDA.n3844 GNDA.n3843 3.4105
R13238 GNDA.n3842 GNDA.n3841 3.4105
R13239 GNDA.n3840 GNDA.n3820 3.4105
R13240 GNDA.n3836 GNDA.n3835 3.4105
R13241 GNDA.n3834 GNDA.n3833 3.4105
R13242 GNDA.n3832 GNDA.n3831 3.4105
R13243 GNDA.n3830 GNDA.n3822 3.4105
R13244 GNDA.n3826 GNDA.n3825 3.4105
R13245 GNDA.n3824 GNDA.n3775 3.4105
R13246 GNDA.n3942 GNDA.n3941 3.4105
R13247 GNDA.n4073 GNDA.n4072 3.4105
R13248 GNDA.n4071 GNDA.n4070 3.4105
R13249 GNDA.n4069 GNDA.n4068 3.4105
R13250 GNDA.n4067 GNDA.n3944 3.4105
R13251 GNDA.n4063 GNDA.n4062 3.4105
R13252 GNDA.n4061 GNDA.n4060 3.4105
R13253 GNDA.n4059 GNDA.n4058 3.4105
R13254 GNDA.n4057 GNDA.n3946 3.4105
R13255 GNDA.n4053 GNDA.n4052 3.4105
R13256 GNDA.n4051 GNDA.n4050 3.4105
R13257 GNDA.n4049 GNDA.n4048 3.4105
R13258 GNDA.n4047 GNDA.n3948 3.4105
R13259 GNDA.n4043 GNDA.n4042 3.4105
R13260 GNDA.n4041 GNDA.n4040 3.4105
R13261 GNDA.n4039 GNDA.n4038 3.4105
R13262 GNDA.n4037 GNDA.n3950 3.4105
R13263 GNDA.n4033 GNDA.n4032 3.4105
R13264 GNDA.n4031 GNDA.n4030 3.4105
R13265 GNDA.n4029 GNDA.n4028 3.4105
R13266 GNDA.n4027 GNDA.n3952 3.4105
R13267 GNDA.n4023 GNDA.n4022 3.4105
R13268 GNDA.n4021 GNDA.n4020 3.4105
R13269 GNDA.n4019 GNDA.n4018 3.4105
R13270 GNDA.n4017 GNDA.n3954 3.4105
R13271 GNDA.n4013 GNDA.n4012 3.4105
R13272 GNDA.n4011 GNDA.n4010 3.4105
R13273 GNDA.n4009 GNDA.n4008 3.4105
R13274 GNDA.n4007 GNDA.n3956 3.4105
R13275 GNDA.n4003 GNDA.n4002 3.4105
R13276 GNDA.n4001 GNDA.n4000 3.4105
R13277 GNDA.n3999 GNDA.n3998 3.4105
R13278 GNDA.n3997 GNDA.n3958 3.4105
R13279 GNDA.n3993 GNDA.n3992 3.4105
R13280 GNDA.n3991 GNDA.n3990 3.4105
R13281 GNDA.n3989 GNDA.n3988 3.4105
R13282 GNDA.n3987 GNDA.n3960 3.4105
R13283 GNDA.n3983 GNDA.n3982 3.4105
R13284 GNDA.n3981 GNDA.n3980 3.4105
R13285 GNDA.n3979 GNDA.n3978 3.4105
R13286 GNDA.n3977 GNDA.n3962 3.4105
R13287 GNDA.n3973 GNDA.n3972 3.4105
R13288 GNDA.n3971 GNDA.n3970 3.4105
R13289 GNDA.n3969 GNDA.n3968 3.4105
R13290 GNDA.n3967 GNDA.n3964 3.4105
R13291 GNDA.n1837 GNDA.n1836 3.4105
R13292 GNDA.n4079 GNDA.n4078 3.4105
R13293 GNDA.n1864 GNDA.n1863 3.4105
R13294 GNDA.n3581 GNDA.n3580 3.4105
R13295 GNDA.n3579 GNDA.n3578 3.4105
R13296 GNDA.n3577 GNDA.n3576 3.4105
R13297 GNDA.n3575 GNDA.n1866 3.4105
R13298 GNDA.n3571 GNDA.n3570 3.4105
R13299 GNDA.n3569 GNDA.n3568 3.4105
R13300 GNDA.n3567 GNDA.n3566 3.4105
R13301 GNDA.n3565 GNDA.n1868 3.4105
R13302 GNDA.n3561 GNDA.n3560 3.4105
R13303 GNDA.n3559 GNDA.n3558 3.4105
R13304 GNDA.n3557 GNDA.n3556 3.4105
R13305 GNDA.n3555 GNDA.n1870 3.4105
R13306 GNDA.n3551 GNDA.n3550 3.4105
R13307 GNDA.n3549 GNDA.n3548 3.4105
R13308 GNDA.n3547 GNDA.n3546 3.4105
R13309 GNDA.n3545 GNDA.n1872 3.4105
R13310 GNDA.n3541 GNDA.n3540 3.4105
R13311 GNDA.n3539 GNDA.n3538 3.4105
R13312 GNDA.n3537 GNDA.n3536 3.4105
R13313 GNDA.n3535 GNDA.n1874 3.4105
R13314 GNDA.n3531 GNDA.n3530 3.4105
R13315 GNDA.n3529 GNDA.n3528 3.4105
R13316 GNDA.n3527 GNDA.n3526 3.4105
R13317 GNDA.n3525 GNDA.n1876 3.4105
R13318 GNDA.n3521 GNDA.n3520 3.4105
R13319 GNDA.n3519 GNDA.n3518 3.4105
R13320 GNDA.n3517 GNDA.n3516 3.4105
R13321 GNDA.n3515 GNDA.n1878 3.4105
R13322 GNDA.n3511 GNDA.n3510 3.4105
R13323 GNDA.n3509 GNDA.n3508 3.4105
R13324 GNDA.n3507 GNDA.n3506 3.4105
R13325 GNDA.n3505 GNDA.n1880 3.4105
R13326 GNDA.n3501 GNDA.n3500 3.4105
R13327 GNDA.n3499 GNDA.n3498 3.4105
R13328 GNDA.n3497 GNDA.n3496 3.4105
R13329 GNDA.n3495 GNDA.n1882 3.4105
R13330 GNDA.n3491 GNDA.n3490 3.4105
R13331 GNDA.n3489 GNDA.n3488 3.4105
R13332 GNDA.n3487 GNDA.n3486 3.4105
R13333 GNDA.n3485 GNDA.n1884 3.4105
R13334 GNDA.n3481 GNDA.n3480 3.4105
R13335 GNDA.n3479 GNDA.n3478 3.4105
R13336 GNDA.n3477 GNDA.n3476 3.4105
R13337 GNDA.n3475 GNDA.n1886 3.4105
R13338 GNDA.n3471 GNDA.n3470 3.4105
R13339 GNDA.n3469 GNDA.n1839 3.4105
R13340 GNDA.n2511 GNDA.n2510 3.4105
R13341 GNDA.n2646 GNDA.n2645 3.4105
R13342 GNDA.n2644 GNDA.n2643 3.4105
R13343 GNDA.n2642 GNDA.n2641 3.4105
R13344 GNDA.n2640 GNDA.n2513 3.4105
R13345 GNDA.n2636 GNDA.n2635 3.4105
R13346 GNDA.n2634 GNDA.n2633 3.4105
R13347 GNDA.n2632 GNDA.n2631 3.4105
R13348 GNDA.n2630 GNDA.n2515 3.4105
R13349 GNDA.n2626 GNDA.n2625 3.4105
R13350 GNDA.n2624 GNDA.n2623 3.4105
R13351 GNDA.n2622 GNDA.n2621 3.4105
R13352 GNDA.n2620 GNDA.n2517 3.4105
R13353 GNDA.n2616 GNDA.n2615 3.4105
R13354 GNDA.n2614 GNDA.n2613 3.4105
R13355 GNDA.n2612 GNDA.n2611 3.4105
R13356 GNDA.n2610 GNDA.n2519 3.4105
R13357 GNDA.n2606 GNDA.n2605 3.4105
R13358 GNDA.n2604 GNDA.n2603 3.4105
R13359 GNDA.n2602 GNDA.n2601 3.4105
R13360 GNDA.n2600 GNDA.n2521 3.4105
R13361 GNDA.n2596 GNDA.n2595 3.4105
R13362 GNDA.n2594 GNDA.n2593 3.4105
R13363 GNDA.n2592 GNDA.n2591 3.4105
R13364 GNDA.n2590 GNDA.n2523 3.4105
R13365 GNDA.n2586 GNDA.n2585 3.4105
R13366 GNDA.n2584 GNDA.n2583 3.4105
R13367 GNDA.n2582 GNDA.n2581 3.4105
R13368 GNDA.n2580 GNDA.n2525 3.4105
R13369 GNDA.n2576 GNDA.n2575 3.4105
R13370 GNDA.n2574 GNDA.n2573 3.4105
R13371 GNDA.n2572 GNDA.n2571 3.4105
R13372 GNDA.n2570 GNDA.n2527 3.4105
R13373 GNDA.n2566 GNDA.n2565 3.4105
R13374 GNDA.n2564 GNDA.n2563 3.4105
R13375 GNDA.n2562 GNDA.n2561 3.4105
R13376 GNDA.n2560 GNDA.n2529 3.4105
R13377 GNDA.n2556 GNDA.n2555 3.4105
R13378 GNDA.n2554 GNDA.n2553 3.4105
R13379 GNDA.n2552 GNDA.n2551 3.4105
R13380 GNDA.n2550 GNDA.n2531 3.4105
R13381 GNDA.n2546 GNDA.n2545 3.4105
R13382 GNDA.n2544 GNDA.n2543 3.4105
R13383 GNDA.n2542 GNDA.n2541 3.4105
R13384 GNDA.n2540 GNDA.n2533 3.4105
R13385 GNDA.n2536 GNDA.n2535 3.4105
R13386 GNDA.n2534 GNDA.n2486 3.4105
R13387 GNDA.n2794 GNDA.n2793 3.4105
R13388 GNDA.n2929 GNDA.n2928 3.4105
R13389 GNDA.n2927 GNDA.n2926 3.4105
R13390 GNDA.n2925 GNDA.n2924 3.4105
R13391 GNDA.n2923 GNDA.n2796 3.4105
R13392 GNDA.n2919 GNDA.n2918 3.4105
R13393 GNDA.n2917 GNDA.n2916 3.4105
R13394 GNDA.n2915 GNDA.n2914 3.4105
R13395 GNDA.n2913 GNDA.n2798 3.4105
R13396 GNDA.n2909 GNDA.n2908 3.4105
R13397 GNDA.n2907 GNDA.n2906 3.4105
R13398 GNDA.n2905 GNDA.n2904 3.4105
R13399 GNDA.n2903 GNDA.n2800 3.4105
R13400 GNDA.n2899 GNDA.n2898 3.4105
R13401 GNDA.n2897 GNDA.n2896 3.4105
R13402 GNDA.n2895 GNDA.n2894 3.4105
R13403 GNDA.n2893 GNDA.n2802 3.4105
R13404 GNDA.n2889 GNDA.n2888 3.4105
R13405 GNDA.n2887 GNDA.n2886 3.4105
R13406 GNDA.n2885 GNDA.n2884 3.4105
R13407 GNDA.n2883 GNDA.n2804 3.4105
R13408 GNDA.n2879 GNDA.n2878 3.4105
R13409 GNDA.n2877 GNDA.n2876 3.4105
R13410 GNDA.n2875 GNDA.n2874 3.4105
R13411 GNDA.n2873 GNDA.n2806 3.4105
R13412 GNDA.n2869 GNDA.n2868 3.4105
R13413 GNDA.n2867 GNDA.n2866 3.4105
R13414 GNDA.n2865 GNDA.n2864 3.4105
R13415 GNDA.n2863 GNDA.n2808 3.4105
R13416 GNDA.n2859 GNDA.n2858 3.4105
R13417 GNDA.n2857 GNDA.n2856 3.4105
R13418 GNDA.n2855 GNDA.n2854 3.4105
R13419 GNDA.n2853 GNDA.n2810 3.4105
R13420 GNDA.n2849 GNDA.n2848 3.4105
R13421 GNDA.n2847 GNDA.n2846 3.4105
R13422 GNDA.n2845 GNDA.n2844 3.4105
R13423 GNDA.n2843 GNDA.n2812 3.4105
R13424 GNDA.n2839 GNDA.n2838 3.4105
R13425 GNDA.n2837 GNDA.n2836 3.4105
R13426 GNDA.n2835 GNDA.n2834 3.4105
R13427 GNDA.n2833 GNDA.n2814 3.4105
R13428 GNDA.n2829 GNDA.n2828 3.4105
R13429 GNDA.n2827 GNDA.n2826 3.4105
R13430 GNDA.n2825 GNDA.n2824 3.4105
R13431 GNDA.n2823 GNDA.n2816 3.4105
R13432 GNDA.n2819 GNDA.n2818 3.4105
R13433 GNDA.n2817 GNDA.n2438 3.4105
R13434 GNDA.n2935 GNDA.n2934 3.4105
R13435 GNDA.n3070 GNDA.n3069 3.4105
R13436 GNDA.n3068 GNDA.n3067 3.4105
R13437 GNDA.n3066 GNDA.n3065 3.4105
R13438 GNDA.n3064 GNDA.n2937 3.4105
R13439 GNDA.n3060 GNDA.n3059 3.4105
R13440 GNDA.n3058 GNDA.n3057 3.4105
R13441 GNDA.n3056 GNDA.n3055 3.4105
R13442 GNDA.n3054 GNDA.n2939 3.4105
R13443 GNDA.n3050 GNDA.n3049 3.4105
R13444 GNDA.n3048 GNDA.n3047 3.4105
R13445 GNDA.n3046 GNDA.n3045 3.4105
R13446 GNDA.n3044 GNDA.n2941 3.4105
R13447 GNDA.n3040 GNDA.n3039 3.4105
R13448 GNDA.n3038 GNDA.n3037 3.4105
R13449 GNDA.n3036 GNDA.n3035 3.4105
R13450 GNDA.n3034 GNDA.n2943 3.4105
R13451 GNDA.n3030 GNDA.n3029 3.4105
R13452 GNDA.n3028 GNDA.n3027 3.4105
R13453 GNDA.n3026 GNDA.n3025 3.4105
R13454 GNDA.n3024 GNDA.n2945 3.4105
R13455 GNDA.n3020 GNDA.n3019 3.4105
R13456 GNDA.n3018 GNDA.n3017 3.4105
R13457 GNDA.n3016 GNDA.n3015 3.4105
R13458 GNDA.n3014 GNDA.n2947 3.4105
R13459 GNDA.n3010 GNDA.n3009 3.4105
R13460 GNDA.n3008 GNDA.n3007 3.4105
R13461 GNDA.n3006 GNDA.n3005 3.4105
R13462 GNDA.n3004 GNDA.n2949 3.4105
R13463 GNDA.n3000 GNDA.n2999 3.4105
R13464 GNDA.n2998 GNDA.n2997 3.4105
R13465 GNDA.n2996 GNDA.n2995 3.4105
R13466 GNDA.n2994 GNDA.n2951 3.4105
R13467 GNDA.n2990 GNDA.n2989 3.4105
R13468 GNDA.n2988 GNDA.n2987 3.4105
R13469 GNDA.n2986 GNDA.n2985 3.4105
R13470 GNDA.n2984 GNDA.n2953 3.4105
R13471 GNDA.n2980 GNDA.n2979 3.4105
R13472 GNDA.n2978 GNDA.n2977 3.4105
R13473 GNDA.n2976 GNDA.n2975 3.4105
R13474 GNDA.n2974 GNDA.n2955 3.4105
R13475 GNDA.n2970 GNDA.n2969 3.4105
R13476 GNDA.n2968 GNDA.n2967 3.4105
R13477 GNDA.n2966 GNDA.n2965 3.4105
R13478 GNDA.n2964 GNDA.n2957 3.4105
R13479 GNDA.n2960 GNDA.n2959 3.4105
R13480 GNDA.n2958 GNDA.n2414 3.4105
R13481 GNDA.n3076 GNDA.n3075 3.4105
R13482 GNDA.n3211 GNDA.n3210 3.4105
R13483 GNDA.n3209 GNDA.n3208 3.4105
R13484 GNDA.n3207 GNDA.n3206 3.4105
R13485 GNDA.n3205 GNDA.n3078 3.4105
R13486 GNDA.n3201 GNDA.n3200 3.4105
R13487 GNDA.n3199 GNDA.n3198 3.4105
R13488 GNDA.n3197 GNDA.n3196 3.4105
R13489 GNDA.n3195 GNDA.n3080 3.4105
R13490 GNDA.n3191 GNDA.n3190 3.4105
R13491 GNDA.n3189 GNDA.n3188 3.4105
R13492 GNDA.n3187 GNDA.n3186 3.4105
R13493 GNDA.n3185 GNDA.n3082 3.4105
R13494 GNDA.n3181 GNDA.n3180 3.4105
R13495 GNDA.n3179 GNDA.n3178 3.4105
R13496 GNDA.n3177 GNDA.n3176 3.4105
R13497 GNDA.n3175 GNDA.n3084 3.4105
R13498 GNDA.n3171 GNDA.n3170 3.4105
R13499 GNDA.n3169 GNDA.n3168 3.4105
R13500 GNDA.n3167 GNDA.n3166 3.4105
R13501 GNDA.n3165 GNDA.n3086 3.4105
R13502 GNDA.n3161 GNDA.n3160 3.4105
R13503 GNDA.n3159 GNDA.n3158 3.4105
R13504 GNDA.n3157 GNDA.n3156 3.4105
R13505 GNDA.n3155 GNDA.n3088 3.4105
R13506 GNDA.n3151 GNDA.n3150 3.4105
R13507 GNDA.n3149 GNDA.n3148 3.4105
R13508 GNDA.n3147 GNDA.n3146 3.4105
R13509 GNDA.n3145 GNDA.n3090 3.4105
R13510 GNDA.n3141 GNDA.n3140 3.4105
R13511 GNDA.n3139 GNDA.n3138 3.4105
R13512 GNDA.n3137 GNDA.n3136 3.4105
R13513 GNDA.n3135 GNDA.n3092 3.4105
R13514 GNDA.n3131 GNDA.n3130 3.4105
R13515 GNDA.n3129 GNDA.n3128 3.4105
R13516 GNDA.n3127 GNDA.n3126 3.4105
R13517 GNDA.n3125 GNDA.n3094 3.4105
R13518 GNDA.n3121 GNDA.n3120 3.4105
R13519 GNDA.n3119 GNDA.n3118 3.4105
R13520 GNDA.n3117 GNDA.n3116 3.4105
R13521 GNDA.n3115 GNDA.n3096 3.4105
R13522 GNDA.n3111 GNDA.n3110 3.4105
R13523 GNDA.n3109 GNDA.n3108 3.4105
R13524 GNDA.n3107 GNDA.n3106 3.4105
R13525 GNDA.n3105 GNDA.n3098 3.4105
R13526 GNDA.n3101 GNDA.n3100 3.4105
R13527 GNDA.n3099 GNDA.n2390 3.4105
R13528 GNDA.n3215 GNDA.n2390 3.4105
R13529 GNDA.n3215 GNDA.n3214 3.4105
R13530 GNDA.n3074 GNDA.n2414 3.4105
R13531 GNDA.n3074 GNDA.n3073 3.4105
R13532 GNDA.n2933 GNDA.n2438 3.4105
R13533 GNDA.n2933 GNDA.n2932 3.4105
R13534 GNDA.n2650 GNDA.n2486 3.4105
R13535 GNDA.n2650 GNDA.n2649 3.4105
R13536 GNDA.n3585 GNDA.n1839 3.4105
R13537 GNDA.n3585 GNDA.n3584 3.4105
R13538 GNDA.n4078 GNDA.n4077 3.4105
R13539 GNDA.n4077 GNDA.n4076 3.4105
R13540 GNDA.n3940 GNDA.n3775 3.4105
R13541 GNDA.n3940 GNDA.n3939 3.4105
R13542 GNDA.n1811 GNDA.n1599 3.4105
R13543 GNDA.n1741 GNDA.n1599 3.4105
R13544 GNDA.n4283 GNDA.n1600 3.4105
R13545 GNDA.n4283 GNDA.n4282 3.4105
R13546 GNDA.n4449 GNDA.n4284 3.4105
R13547 GNDA.n4449 GNDA.n4448 3.4105
R13548 GNDA.n4638 GNDA.n4473 3.4105
R13549 GNDA.n4638 GNDA.n4637 3.4105
R13550 GNDA.n4924 GNDA.n1372 3.4105
R13551 GNDA.n4924 GNDA.n4923 3.4105
R13552 GNDA.n5943 GNDA.n4948 3.4105
R13553 GNDA.n5943 GNDA.n5942 3.4105
R13554 GNDA.n5661 GNDA.n4996 3.4105
R13555 GNDA.n5661 GNDA.n5660 3.4105
R13556 GNDA.n5519 GNDA.n5020 3.4105
R13557 GNDA.n5519 GNDA.n5518 3.4105
R13558 GNDA.n5397 GNDA.n5044 3.4105
R13559 GNDA.n5327 GNDA.n5044 3.4105
R13560 GNDA.n5232 GNDA.n5231 3.4105
R13561 GNDA.n5231 GNDA.n5230 3.4105
R13562 GNDA.n3457 GNDA.n1838 3.4105
R13563 GNDA.n3387 GNDA.n1838 3.4105
R13564 GNDA.n3751 GNDA.n3586 3.4105
R13565 GNDA.n3751 GNDA.n3750 3.4105
R13566 GNDA.n1585 GNDA.n1371 3.4105
R13567 GNDA.n1515 GNDA.n1371 3.4105
R13568 GNDA.n6081 GNDA.n6080 3.4105
R13569 GNDA.n6080 GNDA.n6079 3.4105
R13570 GNDA.n2792 GNDA.n2462 3.4105
R13571 GNDA.n2792 GNDA.n2791 3.4105
R13572 GNDA.n5802 GNDA.n4972 3.4105
R13573 GNDA.n5802 GNDA.n5801 3.4105
R13574 GNDA.n4776 GNDA.n4775 3.4105
R13575 GNDA.n4775 GNDA.n4774 3.4105
R13576 GNDA.n3219 GNDA.n1950 3.4105
R13577 GNDA.n3220 GNDA.n1949 3.4105
R13578 GNDA.n3221 GNDA.n1948 3.4105
R13579 GNDA.n2387 GNDA.n1946 3.4105
R13580 GNDA.n3225 GNDA.n1945 3.4105
R13581 GNDA.n3226 GNDA.n1944 3.4105
R13582 GNDA.n3227 GNDA.n1943 3.4105
R13583 GNDA.n2384 GNDA.n1941 3.4105
R13584 GNDA.n3231 GNDA.n1940 3.4105
R13585 GNDA.n3232 GNDA.n1939 3.4105
R13586 GNDA.n3233 GNDA.n1938 3.4105
R13587 GNDA.n2381 GNDA.n1936 3.4105
R13588 GNDA.n3237 GNDA.n1935 3.4105
R13589 GNDA.n3238 GNDA.n1934 3.4105
R13590 GNDA.n3239 GNDA.n1933 3.4105
R13591 GNDA.n2378 GNDA.n1931 3.4105
R13592 GNDA.n3243 GNDA.n1930 3.4105
R13593 GNDA.n3244 GNDA.n1929 3.4105
R13594 GNDA.n3245 GNDA.n1928 3.4105
R13595 GNDA.n2375 GNDA.n1926 3.4105
R13596 GNDA.n3249 GNDA.n1925 3.4105
R13597 GNDA.n3250 GNDA.n1924 3.4105
R13598 GNDA.n3251 GNDA.n1923 3.4105
R13599 GNDA.n2372 GNDA.n1921 3.4105
R13600 GNDA.n3255 GNDA.n1920 3.4105
R13601 GNDA.n3256 GNDA.n1919 3.4105
R13602 GNDA.n3257 GNDA.n1918 3.4105
R13603 GNDA.n2369 GNDA.n1916 3.4105
R13604 GNDA.n3261 GNDA.n1915 3.4105
R13605 GNDA.n3262 GNDA.n1914 3.4105
R13606 GNDA.n3263 GNDA.n1913 3.4105
R13607 GNDA.n2366 GNDA.n1911 3.4105
R13608 GNDA.n3267 GNDA.n1910 3.4105
R13609 GNDA.n3268 GNDA.n1909 3.4105
R13610 GNDA.n3269 GNDA.n1908 3.4105
R13611 GNDA.n2363 GNDA.n1906 3.4105
R13612 GNDA.n3273 GNDA.n1905 3.4105
R13613 GNDA.n3274 GNDA.n1904 3.4105
R13614 GNDA.n3275 GNDA.n1903 3.4105
R13615 GNDA.n2360 GNDA.n1901 3.4105
R13616 GNDA.n3279 GNDA.n1900 3.4105
R13617 GNDA.n3280 GNDA.n1899 3.4105
R13618 GNDA.n3281 GNDA.n1898 3.4105
R13619 GNDA.n2357 GNDA.n1896 3.4105
R13620 GNDA.n3285 GNDA.n1895 3.4105
R13621 GNDA.n3286 GNDA.n1894 3.4105
R13622 GNDA.n360 GNDA.n359 3.4105
R13623 GNDA.n6444 GNDA.n6443 3.4105
R13624 GNDA.n6311 GNDA.n6310 3.4105
R13625 GNDA.n6439 GNDA.n6438 3.4105
R13626 GNDA.n6437 GNDA.n6436 3.4105
R13627 GNDA.n6435 GNDA.n6315 3.4105
R13628 GNDA.n6314 GNDA.n6313 3.4105
R13629 GNDA.n6431 GNDA.n6430 3.4105
R13630 GNDA.n6429 GNDA.n6428 3.4105
R13631 GNDA.n6427 GNDA.n6319 3.4105
R13632 GNDA.n6318 GNDA.n6317 3.4105
R13633 GNDA.n6423 GNDA.n6422 3.4105
R13634 GNDA.n6421 GNDA.n6420 3.4105
R13635 GNDA.n6419 GNDA.n6323 3.4105
R13636 GNDA.n6322 GNDA.n6321 3.4105
R13637 GNDA.n6415 GNDA.n6414 3.4105
R13638 GNDA.n6413 GNDA.n6412 3.4105
R13639 GNDA.n6411 GNDA.n6327 3.4105
R13640 GNDA.n6326 GNDA.n6325 3.4105
R13641 GNDA.n6407 GNDA.n6406 3.4105
R13642 GNDA.n6405 GNDA.n6404 3.4105
R13643 GNDA.n6403 GNDA.n6331 3.4105
R13644 GNDA.n6330 GNDA.n6329 3.4105
R13645 GNDA.n6399 GNDA.n6398 3.4105
R13646 GNDA.n6397 GNDA.n6396 3.4105
R13647 GNDA.n6395 GNDA.n6335 3.4105
R13648 GNDA.n6334 GNDA.n6333 3.4105
R13649 GNDA.n6391 GNDA.n6390 3.4105
R13650 GNDA.n6389 GNDA.n6388 3.4105
R13651 GNDA.n6387 GNDA.n6339 3.4105
R13652 GNDA.n6338 GNDA.n6337 3.4105
R13653 GNDA.n6383 GNDA.n6382 3.4105
R13654 GNDA.n6381 GNDA.n6380 3.4105
R13655 GNDA.n6379 GNDA.n6343 3.4105
R13656 GNDA.n6342 GNDA.n6341 3.4105
R13657 GNDA.n6375 GNDA.n6374 3.4105
R13658 GNDA.n6373 GNDA.n6372 3.4105
R13659 GNDA.n6371 GNDA.n6347 3.4105
R13660 GNDA.n6346 GNDA.n6345 3.4105
R13661 GNDA.n6367 GNDA.n6366 3.4105
R13662 GNDA.n6365 GNDA.n6364 3.4105
R13663 GNDA.n6363 GNDA.n6351 3.4105
R13664 GNDA.n6350 GNDA.n6349 3.4105
R13665 GNDA.n6359 GNDA.n6358 3.4105
R13666 GNDA.n6357 GNDA.n6356 3.4105
R13667 GNDA.n6355 GNDA.n6354 3.4105
R13668 GNDA.n6617 GNDA.n6616 3.4105
R13669 GNDA.n387 GNDA.n386 3.4105
R13670 GNDA.n521 GNDA.n520 3.4105
R13671 GNDA.n519 GNDA.n518 3.4105
R13672 GNDA.n517 GNDA.n516 3.4105
R13673 GNDA.n515 GNDA.n389 3.4105
R13674 GNDA.n511 GNDA.n510 3.4105
R13675 GNDA.n509 GNDA.n508 3.4105
R13676 GNDA.n507 GNDA.n506 3.4105
R13677 GNDA.n505 GNDA.n391 3.4105
R13678 GNDA.n501 GNDA.n500 3.4105
R13679 GNDA.n499 GNDA.n498 3.4105
R13680 GNDA.n497 GNDA.n496 3.4105
R13681 GNDA.n495 GNDA.n393 3.4105
R13682 GNDA.n491 GNDA.n490 3.4105
R13683 GNDA.n489 GNDA.n488 3.4105
R13684 GNDA.n487 GNDA.n486 3.4105
R13685 GNDA.n485 GNDA.n395 3.4105
R13686 GNDA.n481 GNDA.n480 3.4105
R13687 GNDA.n479 GNDA.n478 3.4105
R13688 GNDA.n477 GNDA.n476 3.4105
R13689 GNDA.n475 GNDA.n397 3.4105
R13690 GNDA.n471 GNDA.n470 3.4105
R13691 GNDA.n469 GNDA.n468 3.4105
R13692 GNDA.n467 GNDA.n466 3.4105
R13693 GNDA.n465 GNDA.n399 3.4105
R13694 GNDA.n461 GNDA.n460 3.4105
R13695 GNDA.n459 GNDA.n458 3.4105
R13696 GNDA.n457 GNDA.n456 3.4105
R13697 GNDA.n455 GNDA.n401 3.4105
R13698 GNDA.n451 GNDA.n450 3.4105
R13699 GNDA.n449 GNDA.n448 3.4105
R13700 GNDA.n447 GNDA.n446 3.4105
R13701 GNDA.n445 GNDA.n403 3.4105
R13702 GNDA.n441 GNDA.n440 3.4105
R13703 GNDA.n439 GNDA.n438 3.4105
R13704 GNDA.n437 GNDA.n436 3.4105
R13705 GNDA.n435 GNDA.n405 3.4105
R13706 GNDA.n431 GNDA.n430 3.4105
R13707 GNDA.n429 GNDA.n428 3.4105
R13708 GNDA.n427 GNDA.n426 3.4105
R13709 GNDA.n425 GNDA.n407 3.4105
R13710 GNDA.n421 GNDA.n420 3.4105
R13711 GNDA.n419 GNDA.n418 3.4105
R13712 GNDA.n417 GNDA.n416 3.4105
R13713 GNDA.n415 GNDA.n409 3.4105
R13714 GNDA.n411 GNDA.n410 3.4105
R13715 GNDA.n6285 GNDA.n6284 3.4105
R13716 GNDA.n6286 GNDA.n362 3.4105
R13717 GNDA.n6286 GNDA.n6285 3.4105
R13718 GNDA.n6615 GNDA.n6287 3.4105
R13719 GNDA.n6616 GNDA.n6615 3.4105
R13720 GNDA.n2163 GNDA.n361 3.4105
R13721 GNDA.n2163 GNDA.n2134 3.4105
R13722 GNDA.n2226 GNDA.n2163 3.4105
R13723 GNDA.n2224 GNDA.n2181 3.4105
R13724 GNDA.n2226 GNDA.n2181 3.4105
R13725 GNDA.n2224 GNDA.n2149 3.4105
R13726 GNDA.n2149 GNDA.n2119 3.4105
R13727 GNDA.n2149 GNDA.n2121 3.4105
R13728 GNDA.n2149 GNDA.n2118 3.4105
R13729 GNDA.n2149 GNDA.n2122 3.4105
R13730 GNDA.n2149 GNDA.n2117 3.4105
R13731 GNDA.n2149 GNDA.n2123 3.4105
R13732 GNDA.n2149 GNDA.n2116 3.4105
R13733 GNDA.n2149 GNDA.n2124 3.4105
R13734 GNDA.n2149 GNDA.n2115 3.4105
R13735 GNDA.n2149 GNDA.n2125 3.4105
R13736 GNDA.n2149 GNDA.n2114 3.4105
R13737 GNDA.n2149 GNDA.n2126 3.4105
R13738 GNDA.n2149 GNDA.n2113 3.4105
R13739 GNDA.n2149 GNDA.n2127 3.4105
R13740 GNDA.n2149 GNDA.n2112 3.4105
R13741 GNDA.n2149 GNDA.n2128 3.4105
R13742 GNDA.n2149 GNDA.n2111 3.4105
R13743 GNDA.n2149 GNDA.n2129 3.4105
R13744 GNDA.n2149 GNDA.n2110 3.4105
R13745 GNDA.n2149 GNDA.n2130 3.4105
R13746 GNDA.n2149 GNDA.n2109 3.4105
R13747 GNDA.n2149 GNDA.n2131 3.4105
R13748 GNDA.n2149 GNDA.n2108 3.4105
R13749 GNDA.n2149 GNDA.n2132 3.4105
R13750 GNDA.n2149 GNDA.n2107 3.4105
R13751 GNDA.n2149 GNDA.n2133 3.4105
R13752 GNDA.n2149 GNDA.n2106 3.4105
R13753 GNDA.n2149 GNDA.n2134 3.4105
R13754 GNDA.n2226 GNDA.n2149 3.4105
R13755 GNDA.n2224 GNDA.n2184 3.4105
R13756 GNDA.n2184 GNDA.n2119 3.4105
R13757 GNDA.n2184 GNDA.n2121 3.4105
R13758 GNDA.n2184 GNDA.n2118 3.4105
R13759 GNDA.n2184 GNDA.n2122 3.4105
R13760 GNDA.n2184 GNDA.n2117 3.4105
R13761 GNDA.n2184 GNDA.n2123 3.4105
R13762 GNDA.n2184 GNDA.n2116 3.4105
R13763 GNDA.n2184 GNDA.n2124 3.4105
R13764 GNDA.n2184 GNDA.n2115 3.4105
R13765 GNDA.n2184 GNDA.n2125 3.4105
R13766 GNDA.n2184 GNDA.n2114 3.4105
R13767 GNDA.n2184 GNDA.n2126 3.4105
R13768 GNDA.n2184 GNDA.n2113 3.4105
R13769 GNDA.n2184 GNDA.n2127 3.4105
R13770 GNDA.n2184 GNDA.n2112 3.4105
R13771 GNDA.n2184 GNDA.n2128 3.4105
R13772 GNDA.n2184 GNDA.n2111 3.4105
R13773 GNDA.n2184 GNDA.n2129 3.4105
R13774 GNDA.n2184 GNDA.n2110 3.4105
R13775 GNDA.n2184 GNDA.n2130 3.4105
R13776 GNDA.n2184 GNDA.n2109 3.4105
R13777 GNDA.n2184 GNDA.n2131 3.4105
R13778 GNDA.n2184 GNDA.n2108 3.4105
R13779 GNDA.n2184 GNDA.n2132 3.4105
R13780 GNDA.n2184 GNDA.n2107 3.4105
R13781 GNDA.n2184 GNDA.n2133 3.4105
R13782 GNDA.n2184 GNDA.n2106 3.4105
R13783 GNDA.n2184 GNDA.n2134 3.4105
R13784 GNDA.n2226 GNDA.n2184 3.4105
R13785 GNDA.n2224 GNDA.n2148 3.4105
R13786 GNDA.n2148 GNDA.n2119 3.4105
R13787 GNDA.n2148 GNDA.n2121 3.4105
R13788 GNDA.n2148 GNDA.n2118 3.4105
R13789 GNDA.n2148 GNDA.n2122 3.4105
R13790 GNDA.n2148 GNDA.n2117 3.4105
R13791 GNDA.n2148 GNDA.n2123 3.4105
R13792 GNDA.n2148 GNDA.n2116 3.4105
R13793 GNDA.n2148 GNDA.n2124 3.4105
R13794 GNDA.n2148 GNDA.n2115 3.4105
R13795 GNDA.n2148 GNDA.n2125 3.4105
R13796 GNDA.n2148 GNDA.n2114 3.4105
R13797 GNDA.n2148 GNDA.n2126 3.4105
R13798 GNDA.n2148 GNDA.n2113 3.4105
R13799 GNDA.n2148 GNDA.n2127 3.4105
R13800 GNDA.n2148 GNDA.n2112 3.4105
R13801 GNDA.n2148 GNDA.n2128 3.4105
R13802 GNDA.n2148 GNDA.n2111 3.4105
R13803 GNDA.n2148 GNDA.n2129 3.4105
R13804 GNDA.n2148 GNDA.n2110 3.4105
R13805 GNDA.n2148 GNDA.n2130 3.4105
R13806 GNDA.n2148 GNDA.n2109 3.4105
R13807 GNDA.n2148 GNDA.n2131 3.4105
R13808 GNDA.n2148 GNDA.n2108 3.4105
R13809 GNDA.n2148 GNDA.n2132 3.4105
R13810 GNDA.n2148 GNDA.n2107 3.4105
R13811 GNDA.n2148 GNDA.n2133 3.4105
R13812 GNDA.n2148 GNDA.n2106 3.4105
R13813 GNDA.n2148 GNDA.n2134 3.4105
R13814 GNDA.n2226 GNDA.n2148 3.4105
R13815 GNDA.n2224 GNDA.n2187 3.4105
R13816 GNDA.n2187 GNDA.n2119 3.4105
R13817 GNDA.n2187 GNDA.n2121 3.4105
R13818 GNDA.n2187 GNDA.n2118 3.4105
R13819 GNDA.n2187 GNDA.n2122 3.4105
R13820 GNDA.n2187 GNDA.n2117 3.4105
R13821 GNDA.n2187 GNDA.n2123 3.4105
R13822 GNDA.n2187 GNDA.n2116 3.4105
R13823 GNDA.n2187 GNDA.n2124 3.4105
R13824 GNDA.n2187 GNDA.n2115 3.4105
R13825 GNDA.n2187 GNDA.n2125 3.4105
R13826 GNDA.n2187 GNDA.n2114 3.4105
R13827 GNDA.n2187 GNDA.n2126 3.4105
R13828 GNDA.n2187 GNDA.n2113 3.4105
R13829 GNDA.n2187 GNDA.n2127 3.4105
R13830 GNDA.n2187 GNDA.n2112 3.4105
R13831 GNDA.n2187 GNDA.n2128 3.4105
R13832 GNDA.n2187 GNDA.n2111 3.4105
R13833 GNDA.n2187 GNDA.n2129 3.4105
R13834 GNDA.n2187 GNDA.n2110 3.4105
R13835 GNDA.n2187 GNDA.n2130 3.4105
R13836 GNDA.n2187 GNDA.n2109 3.4105
R13837 GNDA.n2187 GNDA.n2131 3.4105
R13838 GNDA.n2187 GNDA.n2108 3.4105
R13839 GNDA.n2187 GNDA.n2132 3.4105
R13840 GNDA.n2187 GNDA.n2107 3.4105
R13841 GNDA.n2187 GNDA.n2133 3.4105
R13842 GNDA.n2187 GNDA.n2106 3.4105
R13843 GNDA.n2187 GNDA.n2134 3.4105
R13844 GNDA.n2226 GNDA.n2187 3.4105
R13845 GNDA.n2224 GNDA.n2147 3.4105
R13846 GNDA.n2147 GNDA.n2119 3.4105
R13847 GNDA.n2147 GNDA.n2121 3.4105
R13848 GNDA.n2147 GNDA.n2118 3.4105
R13849 GNDA.n2147 GNDA.n2122 3.4105
R13850 GNDA.n2147 GNDA.n2117 3.4105
R13851 GNDA.n2147 GNDA.n2123 3.4105
R13852 GNDA.n2147 GNDA.n2116 3.4105
R13853 GNDA.n2147 GNDA.n2124 3.4105
R13854 GNDA.n2147 GNDA.n2115 3.4105
R13855 GNDA.n2147 GNDA.n2125 3.4105
R13856 GNDA.n2147 GNDA.n2114 3.4105
R13857 GNDA.n2147 GNDA.n2126 3.4105
R13858 GNDA.n2147 GNDA.n2113 3.4105
R13859 GNDA.n2147 GNDA.n2127 3.4105
R13860 GNDA.n2147 GNDA.n2112 3.4105
R13861 GNDA.n2147 GNDA.n2128 3.4105
R13862 GNDA.n2147 GNDA.n2111 3.4105
R13863 GNDA.n2147 GNDA.n2129 3.4105
R13864 GNDA.n2147 GNDA.n2110 3.4105
R13865 GNDA.n2147 GNDA.n2130 3.4105
R13866 GNDA.n2147 GNDA.n2109 3.4105
R13867 GNDA.n2147 GNDA.n2131 3.4105
R13868 GNDA.n2147 GNDA.n2108 3.4105
R13869 GNDA.n2147 GNDA.n2132 3.4105
R13870 GNDA.n2147 GNDA.n2107 3.4105
R13871 GNDA.n2147 GNDA.n2133 3.4105
R13872 GNDA.n2147 GNDA.n2106 3.4105
R13873 GNDA.n2147 GNDA.n2134 3.4105
R13874 GNDA.n2226 GNDA.n2147 3.4105
R13875 GNDA.n2224 GNDA.n2190 3.4105
R13876 GNDA.n2190 GNDA.n2119 3.4105
R13877 GNDA.n2190 GNDA.n2121 3.4105
R13878 GNDA.n2190 GNDA.n2118 3.4105
R13879 GNDA.n2190 GNDA.n2122 3.4105
R13880 GNDA.n2190 GNDA.n2117 3.4105
R13881 GNDA.n2190 GNDA.n2123 3.4105
R13882 GNDA.n2190 GNDA.n2116 3.4105
R13883 GNDA.n2190 GNDA.n2124 3.4105
R13884 GNDA.n2190 GNDA.n2115 3.4105
R13885 GNDA.n2190 GNDA.n2125 3.4105
R13886 GNDA.n2190 GNDA.n2114 3.4105
R13887 GNDA.n2190 GNDA.n2126 3.4105
R13888 GNDA.n2190 GNDA.n2113 3.4105
R13889 GNDA.n2190 GNDA.n2127 3.4105
R13890 GNDA.n2190 GNDA.n2112 3.4105
R13891 GNDA.n2190 GNDA.n2128 3.4105
R13892 GNDA.n2190 GNDA.n2111 3.4105
R13893 GNDA.n2190 GNDA.n2129 3.4105
R13894 GNDA.n2190 GNDA.n2110 3.4105
R13895 GNDA.n2190 GNDA.n2130 3.4105
R13896 GNDA.n2190 GNDA.n2109 3.4105
R13897 GNDA.n2190 GNDA.n2131 3.4105
R13898 GNDA.n2190 GNDA.n2108 3.4105
R13899 GNDA.n2190 GNDA.n2132 3.4105
R13900 GNDA.n2190 GNDA.n2107 3.4105
R13901 GNDA.n2190 GNDA.n2133 3.4105
R13902 GNDA.n2190 GNDA.n2106 3.4105
R13903 GNDA.n2190 GNDA.n2134 3.4105
R13904 GNDA.n2226 GNDA.n2190 3.4105
R13905 GNDA.n2224 GNDA.n2146 3.4105
R13906 GNDA.n2146 GNDA.n2119 3.4105
R13907 GNDA.n2146 GNDA.n2121 3.4105
R13908 GNDA.n2146 GNDA.n2118 3.4105
R13909 GNDA.n2146 GNDA.n2122 3.4105
R13910 GNDA.n2146 GNDA.n2117 3.4105
R13911 GNDA.n2146 GNDA.n2123 3.4105
R13912 GNDA.n2146 GNDA.n2116 3.4105
R13913 GNDA.n2146 GNDA.n2124 3.4105
R13914 GNDA.n2146 GNDA.n2115 3.4105
R13915 GNDA.n2146 GNDA.n2125 3.4105
R13916 GNDA.n2146 GNDA.n2114 3.4105
R13917 GNDA.n2146 GNDA.n2126 3.4105
R13918 GNDA.n2146 GNDA.n2113 3.4105
R13919 GNDA.n2146 GNDA.n2127 3.4105
R13920 GNDA.n2146 GNDA.n2112 3.4105
R13921 GNDA.n2146 GNDA.n2128 3.4105
R13922 GNDA.n2146 GNDA.n2111 3.4105
R13923 GNDA.n2146 GNDA.n2129 3.4105
R13924 GNDA.n2146 GNDA.n2110 3.4105
R13925 GNDA.n2146 GNDA.n2130 3.4105
R13926 GNDA.n2146 GNDA.n2109 3.4105
R13927 GNDA.n2146 GNDA.n2131 3.4105
R13928 GNDA.n2146 GNDA.n2108 3.4105
R13929 GNDA.n2146 GNDA.n2132 3.4105
R13930 GNDA.n2146 GNDA.n2107 3.4105
R13931 GNDA.n2146 GNDA.n2133 3.4105
R13932 GNDA.n2146 GNDA.n2106 3.4105
R13933 GNDA.n2146 GNDA.n2134 3.4105
R13934 GNDA.n2226 GNDA.n2146 3.4105
R13935 GNDA.n2224 GNDA.n2193 3.4105
R13936 GNDA.n2193 GNDA.n2119 3.4105
R13937 GNDA.n2193 GNDA.n2121 3.4105
R13938 GNDA.n2193 GNDA.n2118 3.4105
R13939 GNDA.n2193 GNDA.n2122 3.4105
R13940 GNDA.n2193 GNDA.n2117 3.4105
R13941 GNDA.n2193 GNDA.n2123 3.4105
R13942 GNDA.n2193 GNDA.n2116 3.4105
R13943 GNDA.n2193 GNDA.n2124 3.4105
R13944 GNDA.n2193 GNDA.n2115 3.4105
R13945 GNDA.n2193 GNDA.n2125 3.4105
R13946 GNDA.n2193 GNDA.n2114 3.4105
R13947 GNDA.n2193 GNDA.n2126 3.4105
R13948 GNDA.n2193 GNDA.n2113 3.4105
R13949 GNDA.n2193 GNDA.n2127 3.4105
R13950 GNDA.n2193 GNDA.n2112 3.4105
R13951 GNDA.n2193 GNDA.n2128 3.4105
R13952 GNDA.n2193 GNDA.n2111 3.4105
R13953 GNDA.n2193 GNDA.n2129 3.4105
R13954 GNDA.n2193 GNDA.n2110 3.4105
R13955 GNDA.n2193 GNDA.n2130 3.4105
R13956 GNDA.n2193 GNDA.n2109 3.4105
R13957 GNDA.n2193 GNDA.n2131 3.4105
R13958 GNDA.n2193 GNDA.n2108 3.4105
R13959 GNDA.n2193 GNDA.n2132 3.4105
R13960 GNDA.n2193 GNDA.n2107 3.4105
R13961 GNDA.n2193 GNDA.n2133 3.4105
R13962 GNDA.n2193 GNDA.n2106 3.4105
R13963 GNDA.n2193 GNDA.n2134 3.4105
R13964 GNDA.n2226 GNDA.n2193 3.4105
R13965 GNDA.n2224 GNDA.n2145 3.4105
R13966 GNDA.n2145 GNDA.n2119 3.4105
R13967 GNDA.n2145 GNDA.n2121 3.4105
R13968 GNDA.n2145 GNDA.n2118 3.4105
R13969 GNDA.n2145 GNDA.n2122 3.4105
R13970 GNDA.n2145 GNDA.n2117 3.4105
R13971 GNDA.n2145 GNDA.n2123 3.4105
R13972 GNDA.n2145 GNDA.n2116 3.4105
R13973 GNDA.n2145 GNDA.n2124 3.4105
R13974 GNDA.n2145 GNDA.n2115 3.4105
R13975 GNDA.n2145 GNDA.n2125 3.4105
R13976 GNDA.n2145 GNDA.n2114 3.4105
R13977 GNDA.n2145 GNDA.n2126 3.4105
R13978 GNDA.n2145 GNDA.n2113 3.4105
R13979 GNDA.n2145 GNDA.n2127 3.4105
R13980 GNDA.n2145 GNDA.n2112 3.4105
R13981 GNDA.n2145 GNDA.n2128 3.4105
R13982 GNDA.n2145 GNDA.n2111 3.4105
R13983 GNDA.n2145 GNDA.n2129 3.4105
R13984 GNDA.n2145 GNDA.n2110 3.4105
R13985 GNDA.n2145 GNDA.n2130 3.4105
R13986 GNDA.n2145 GNDA.n2109 3.4105
R13987 GNDA.n2145 GNDA.n2131 3.4105
R13988 GNDA.n2145 GNDA.n2108 3.4105
R13989 GNDA.n2145 GNDA.n2132 3.4105
R13990 GNDA.n2145 GNDA.n2107 3.4105
R13991 GNDA.n2145 GNDA.n2133 3.4105
R13992 GNDA.n2145 GNDA.n2106 3.4105
R13993 GNDA.n2145 GNDA.n2134 3.4105
R13994 GNDA.n2226 GNDA.n2145 3.4105
R13995 GNDA.n2224 GNDA.n2196 3.4105
R13996 GNDA.n2196 GNDA.n2119 3.4105
R13997 GNDA.n2196 GNDA.n2121 3.4105
R13998 GNDA.n2196 GNDA.n2118 3.4105
R13999 GNDA.n2196 GNDA.n2122 3.4105
R14000 GNDA.n2196 GNDA.n2117 3.4105
R14001 GNDA.n2196 GNDA.n2123 3.4105
R14002 GNDA.n2196 GNDA.n2116 3.4105
R14003 GNDA.n2196 GNDA.n2124 3.4105
R14004 GNDA.n2196 GNDA.n2115 3.4105
R14005 GNDA.n2196 GNDA.n2125 3.4105
R14006 GNDA.n2196 GNDA.n2114 3.4105
R14007 GNDA.n2196 GNDA.n2126 3.4105
R14008 GNDA.n2196 GNDA.n2113 3.4105
R14009 GNDA.n2196 GNDA.n2127 3.4105
R14010 GNDA.n2196 GNDA.n2112 3.4105
R14011 GNDA.n2196 GNDA.n2128 3.4105
R14012 GNDA.n2196 GNDA.n2111 3.4105
R14013 GNDA.n2196 GNDA.n2129 3.4105
R14014 GNDA.n2196 GNDA.n2110 3.4105
R14015 GNDA.n2196 GNDA.n2130 3.4105
R14016 GNDA.n2196 GNDA.n2109 3.4105
R14017 GNDA.n2196 GNDA.n2131 3.4105
R14018 GNDA.n2196 GNDA.n2108 3.4105
R14019 GNDA.n2196 GNDA.n2132 3.4105
R14020 GNDA.n2196 GNDA.n2107 3.4105
R14021 GNDA.n2196 GNDA.n2133 3.4105
R14022 GNDA.n2196 GNDA.n2106 3.4105
R14023 GNDA.n2196 GNDA.n2134 3.4105
R14024 GNDA.n2226 GNDA.n2196 3.4105
R14025 GNDA.n2224 GNDA.n2144 3.4105
R14026 GNDA.n2144 GNDA.n2119 3.4105
R14027 GNDA.n2144 GNDA.n2121 3.4105
R14028 GNDA.n2144 GNDA.n2118 3.4105
R14029 GNDA.n2144 GNDA.n2122 3.4105
R14030 GNDA.n2144 GNDA.n2117 3.4105
R14031 GNDA.n2144 GNDA.n2123 3.4105
R14032 GNDA.n2144 GNDA.n2116 3.4105
R14033 GNDA.n2144 GNDA.n2124 3.4105
R14034 GNDA.n2144 GNDA.n2115 3.4105
R14035 GNDA.n2144 GNDA.n2125 3.4105
R14036 GNDA.n2144 GNDA.n2114 3.4105
R14037 GNDA.n2144 GNDA.n2126 3.4105
R14038 GNDA.n2144 GNDA.n2113 3.4105
R14039 GNDA.n2144 GNDA.n2127 3.4105
R14040 GNDA.n2144 GNDA.n2112 3.4105
R14041 GNDA.n2144 GNDA.n2128 3.4105
R14042 GNDA.n2144 GNDA.n2111 3.4105
R14043 GNDA.n2144 GNDA.n2129 3.4105
R14044 GNDA.n2144 GNDA.n2110 3.4105
R14045 GNDA.n2144 GNDA.n2130 3.4105
R14046 GNDA.n2144 GNDA.n2109 3.4105
R14047 GNDA.n2144 GNDA.n2131 3.4105
R14048 GNDA.n2144 GNDA.n2108 3.4105
R14049 GNDA.n2144 GNDA.n2132 3.4105
R14050 GNDA.n2144 GNDA.n2107 3.4105
R14051 GNDA.n2144 GNDA.n2133 3.4105
R14052 GNDA.n2144 GNDA.n2106 3.4105
R14053 GNDA.n2144 GNDA.n2134 3.4105
R14054 GNDA.n2226 GNDA.n2144 3.4105
R14055 GNDA.n2224 GNDA.n2199 3.4105
R14056 GNDA.n2199 GNDA.n2119 3.4105
R14057 GNDA.n2199 GNDA.n2121 3.4105
R14058 GNDA.n2199 GNDA.n2118 3.4105
R14059 GNDA.n2199 GNDA.n2122 3.4105
R14060 GNDA.n2199 GNDA.n2117 3.4105
R14061 GNDA.n2199 GNDA.n2123 3.4105
R14062 GNDA.n2199 GNDA.n2116 3.4105
R14063 GNDA.n2199 GNDA.n2124 3.4105
R14064 GNDA.n2199 GNDA.n2115 3.4105
R14065 GNDA.n2199 GNDA.n2125 3.4105
R14066 GNDA.n2199 GNDA.n2114 3.4105
R14067 GNDA.n2199 GNDA.n2126 3.4105
R14068 GNDA.n2199 GNDA.n2113 3.4105
R14069 GNDA.n2199 GNDA.n2127 3.4105
R14070 GNDA.n2199 GNDA.n2112 3.4105
R14071 GNDA.n2199 GNDA.n2128 3.4105
R14072 GNDA.n2199 GNDA.n2111 3.4105
R14073 GNDA.n2199 GNDA.n2129 3.4105
R14074 GNDA.n2199 GNDA.n2110 3.4105
R14075 GNDA.n2199 GNDA.n2130 3.4105
R14076 GNDA.n2199 GNDA.n2109 3.4105
R14077 GNDA.n2199 GNDA.n2131 3.4105
R14078 GNDA.n2199 GNDA.n2108 3.4105
R14079 GNDA.n2199 GNDA.n2132 3.4105
R14080 GNDA.n2199 GNDA.n2107 3.4105
R14081 GNDA.n2199 GNDA.n2133 3.4105
R14082 GNDA.n2199 GNDA.n2106 3.4105
R14083 GNDA.n2199 GNDA.n2134 3.4105
R14084 GNDA.n2226 GNDA.n2199 3.4105
R14085 GNDA.n2224 GNDA.n2143 3.4105
R14086 GNDA.n2143 GNDA.n2119 3.4105
R14087 GNDA.n2143 GNDA.n2121 3.4105
R14088 GNDA.n2143 GNDA.n2118 3.4105
R14089 GNDA.n2143 GNDA.n2122 3.4105
R14090 GNDA.n2143 GNDA.n2117 3.4105
R14091 GNDA.n2143 GNDA.n2123 3.4105
R14092 GNDA.n2143 GNDA.n2116 3.4105
R14093 GNDA.n2143 GNDA.n2124 3.4105
R14094 GNDA.n2143 GNDA.n2115 3.4105
R14095 GNDA.n2143 GNDA.n2125 3.4105
R14096 GNDA.n2143 GNDA.n2114 3.4105
R14097 GNDA.n2143 GNDA.n2126 3.4105
R14098 GNDA.n2143 GNDA.n2113 3.4105
R14099 GNDA.n2143 GNDA.n2127 3.4105
R14100 GNDA.n2143 GNDA.n2112 3.4105
R14101 GNDA.n2143 GNDA.n2128 3.4105
R14102 GNDA.n2143 GNDA.n2111 3.4105
R14103 GNDA.n2143 GNDA.n2129 3.4105
R14104 GNDA.n2143 GNDA.n2110 3.4105
R14105 GNDA.n2143 GNDA.n2130 3.4105
R14106 GNDA.n2143 GNDA.n2109 3.4105
R14107 GNDA.n2143 GNDA.n2131 3.4105
R14108 GNDA.n2143 GNDA.n2108 3.4105
R14109 GNDA.n2143 GNDA.n2132 3.4105
R14110 GNDA.n2143 GNDA.n2107 3.4105
R14111 GNDA.n2143 GNDA.n2133 3.4105
R14112 GNDA.n2143 GNDA.n2106 3.4105
R14113 GNDA.n2143 GNDA.n2134 3.4105
R14114 GNDA.n2226 GNDA.n2143 3.4105
R14115 GNDA.n2224 GNDA.n2202 3.4105
R14116 GNDA.n2202 GNDA.n2119 3.4105
R14117 GNDA.n2202 GNDA.n2121 3.4105
R14118 GNDA.n2202 GNDA.n2118 3.4105
R14119 GNDA.n2202 GNDA.n2122 3.4105
R14120 GNDA.n2202 GNDA.n2117 3.4105
R14121 GNDA.n2202 GNDA.n2123 3.4105
R14122 GNDA.n2202 GNDA.n2116 3.4105
R14123 GNDA.n2202 GNDA.n2124 3.4105
R14124 GNDA.n2202 GNDA.n2115 3.4105
R14125 GNDA.n2202 GNDA.n2125 3.4105
R14126 GNDA.n2202 GNDA.n2114 3.4105
R14127 GNDA.n2202 GNDA.n2126 3.4105
R14128 GNDA.n2202 GNDA.n2113 3.4105
R14129 GNDA.n2202 GNDA.n2127 3.4105
R14130 GNDA.n2202 GNDA.n2112 3.4105
R14131 GNDA.n2202 GNDA.n2128 3.4105
R14132 GNDA.n2202 GNDA.n2111 3.4105
R14133 GNDA.n2202 GNDA.n2129 3.4105
R14134 GNDA.n2202 GNDA.n2110 3.4105
R14135 GNDA.n2202 GNDA.n2130 3.4105
R14136 GNDA.n2202 GNDA.n2109 3.4105
R14137 GNDA.n2202 GNDA.n2131 3.4105
R14138 GNDA.n2202 GNDA.n2108 3.4105
R14139 GNDA.n2202 GNDA.n2132 3.4105
R14140 GNDA.n2202 GNDA.n2107 3.4105
R14141 GNDA.n2202 GNDA.n2133 3.4105
R14142 GNDA.n2202 GNDA.n2106 3.4105
R14143 GNDA.n2202 GNDA.n2134 3.4105
R14144 GNDA.n2226 GNDA.n2202 3.4105
R14145 GNDA.n2224 GNDA.n2142 3.4105
R14146 GNDA.n2142 GNDA.n2119 3.4105
R14147 GNDA.n2142 GNDA.n2121 3.4105
R14148 GNDA.n2142 GNDA.n2118 3.4105
R14149 GNDA.n2142 GNDA.n2122 3.4105
R14150 GNDA.n2142 GNDA.n2117 3.4105
R14151 GNDA.n2142 GNDA.n2123 3.4105
R14152 GNDA.n2142 GNDA.n2116 3.4105
R14153 GNDA.n2142 GNDA.n2124 3.4105
R14154 GNDA.n2142 GNDA.n2115 3.4105
R14155 GNDA.n2142 GNDA.n2125 3.4105
R14156 GNDA.n2142 GNDA.n2114 3.4105
R14157 GNDA.n2142 GNDA.n2126 3.4105
R14158 GNDA.n2142 GNDA.n2113 3.4105
R14159 GNDA.n2142 GNDA.n2127 3.4105
R14160 GNDA.n2142 GNDA.n2112 3.4105
R14161 GNDA.n2142 GNDA.n2128 3.4105
R14162 GNDA.n2142 GNDA.n2111 3.4105
R14163 GNDA.n2142 GNDA.n2129 3.4105
R14164 GNDA.n2142 GNDA.n2110 3.4105
R14165 GNDA.n2142 GNDA.n2130 3.4105
R14166 GNDA.n2142 GNDA.n2109 3.4105
R14167 GNDA.n2142 GNDA.n2131 3.4105
R14168 GNDA.n2142 GNDA.n2108 3.4105
R14169 GNDA.n2142 GNDA.n2132 3.4105
R14170 GNDA.n2142 GNDA.n2107 3.4105
R14171 GNDA.n2142 GNDA.n2133 3.4105
R14172 GNDA.n2142 GNDA.n2106 3.4105
R14173 GNDA.n2142 GNDA.n2134 3.4105
R14174 GNDA.n2226 GNDA.n2142 3.4105
R14175 GNDA.n2224 GNDA.n2205 3.4105
R14176 GNDA.n2205 GNDA.n2119 3.4105
R14177 GNDA.n2205 GNDA.n2121 3.4105
R14178 GNDA.n2205 GNDA.n2118 3.4105
R14179 GNDA.n2205 GNDA.n2122 3.4105
R14180 GNDA.n2205 GNDA.n2117 3.4105
R14181 GNDA.n2205 GNDA.n2123 3.4105
R14182 GNDA.n2205 GNDA.n2116 3.4105
R14183 GNDA.n2205 GNDA.n2124 3.4105
R14184 GNDA.n2205 GNDA.n2115 3.4105
R14185 GNDA.n2205 GNDA.n2125 3.4105
R14186 GNDA.n2205 GNDA.n2114 3.4105
R14187 GNDA.n2205 GNDA.n2126 3.4105
R14188 GNDA.n2205 GNDA.n2113 3.4105
R14189 GNDA.n2205 GNDA.n2127 3.4105
R14190 GNDA.n2205 GNDA.n2112 3.4105
R14191 GNDA.n2205 GNDA.n2128 3.4105
R14192 GNDA.n2205 GNDA.n2111 3.4105
R14193 GNDA.n2205 GNDA.n2129 3.4105
R14194 GNDA.n2205 GNDA.n2110 3.4105
R14195 GNDA.n2205 GNDA.n2130 3.4105
R14196 GNDA.n2205 GNDA.n2109 3.4105
R14197 GNDA.n2205 GNDA.n2131 3.4105
R14198 GNDA.n2205 GNDA.n2108 3.4105
R14199 GNDA.n2205 GNDA.n2132 3.4105
R14200 GNDA.n2205 GNDA.n2107 3.4105
R14201 GNDA.n2205 GNDA.n2133 3.4105
R14202 GNDA.n2205 GNDA.n2106 3.4105
R14203 GNDA.n2205 GNDA.n2134 3.4105
R14204 GNDA.n2226 GNDA.n2205 3.4105
R14205 GNDA.n2224 GNDA.n2141 3.4105
R14206 GNDA.n2141 GNDA.n2119 3.4105
R14207 GNDA.n2141 GNDA.n2121 3.4105
R14208 GNDA.n2141 GNDA.n2118 3.4105
R14209 GNDA.n2141 GNDA.n2122 3.4105
R14210 GNDA.n2141 GNDA.n2117 3.4105
R14211 GNDA.n2141 GNDA.n2123 3.4105
R14212 GNDA.n2141 GNDA.n2116 3.4105
R14213 GNDA.n2141 GNDA.n2124 3.4105
R14214 GNDA.n2141 GNDA.n2115 3.4105
R14215 GNDA.n2141 GNDA.n2125 3.4105
R14216 GNDA.n2141 GNDA.n2114 3.4105
R14217 GNDA.n2141 GNDA.n2126 3.4105
R14218 GNDA.n2141 GNDA.n2113 3.4105
R14219 GNDA.n2141 GNDA.n2127 3.4105
R14220 GNDA.n2141 GNDA.n2112 3.4105
R14221 GNDA.n2141 GNDA.n2128 3.4105
R14222 GNDA.n2141 GNDA.n2111 3.4105
R14223 GNDA.n2141 GNDA.n2129 3.4105
R14224 GNDA.n2141 GNDA.n2110 3.4105
R14225 GNDA.n2141 GNDA.n2130 3.4105
R14226 GNDA.n2141 GNDA.n2109 3.4105
R14227 GNDA.n2141 GNDA.n2131 3.4105
R14228 GNDA.n2141 GNDA.n2108 3.4105
R14229 GNDA.n2141 GNDA.n2132 3.4105
R14230 GNDA.n2141 GNDA.n2107 3.4105
R14231 GNDA.n2141 GNDA.n2133 3.4105
R14232 GNDA.n2141 GNDA.n2106 3.4105
R14233 GNDA.n2141 GNDA.n2134 3.4105
R14234 GNDA.n2226 GNDA.n2141 3.4105
R14235 GNDA.n2224 GNDA.n2208 3.4105
R14236 GNDA.n2208 GNDA.n2119 3.4105
R14237 GNDA.n2208 GNDA.n2121 3.4105
R14238 GNDA.n2208 GNDA.n2118 3.4105
R14239 GNDA.n2208 GNDA.n2122 3.4105
R14240 GNDA.n2208 GNDA.n2117 3.4105
R14241 GNDA.n2208 GNDA.n2123 3.4105
R14242 GNDA.n2208 GNDA.n2116 3.4105
R14243 GNDA.n2208 GNDA.n2124 3.4105
R14244 GNDA.n2208 GNDA.n2115 3.4105
R14245 GNDA.n2208 GNDA.n2125 3.4105
R14246 GNDA.n2208 GNDA.n2114 3.4105
R14247 GNDA.n2208 GNDA.n2126 3.4105
R14248 GNDA.n2208 GNDA.n2113 3.4105
R14249 GNDA.n2208 GNDA.n2127 3.4105
R14250 GNDA.n2208 GNDA.n2112 3.4105
R14251 GNDA.n2208 GNDA.n2128 3.4105
R14252 GNDA.n2208 GNDA.n2111 3.4105
R14253 GNDA.n2208 GNDA.n2129 3.4105
R14254 GNDA.n2208 GNDA.n2110 3.4105
R14255 GNDA.n2208 GNDA.n2130 3.4105
R14256 GNDA.n2208 GNDA.n2109 3.4105
R14257 GNDA.n2208 GNDA.n2131 3.4105
R14258 GNDA.n2208 GNDA.n2108 3.4105
R14259 GNDA.n2208 GNDA.n2132 3.4105
R14260 GNDA.n2208 GNDA.n2107 3.4105
R14261 GNDA.n2208 GNDA.n2133 3.4105
R14262 GNDA.n2208 GNDA.n2106 3.4105
R14263 GNDA.n2208 GNDA.n2134 3.4105
R14264 GNDA.n2226 GNDA.n2208 3.4105
R14265 GNDA.n2224 GNDA.n2140 3.4105
R14266 GNDA.n2140 GNDA.n2119 3.4105
R14267 GNDA.n2140 GNDA.n2121 3.4105
R14268 GNDA.n2140 GNDA.n2118 3.4105
R14269 GNDA.n2140 GNDA.n2122 3.4105
R14270 GNDA.n2140 GNDA.n2117 3.4105
R14271 GNDA.n2140 GNDA.n2123 3.4105
R14272 GNDA.n2140 GNDA.n2116 3.4105
R14273 GNDA.n2140 GNDA.n2124 3.4105
R14274 GNDA.n2140 GNDA.n2115 3.4105
R14275 GNDA.n2140 GNDA.n2125 3.4105
R14276 GNDA.n2140 GNDA.n2114 3.4105
R14277 GNDA.n2140 GNDA.n2126 3.4105
R14278 GNDA.n2140 GNDA.n2113 3.4105
R14279 GNDA.n2140 GNDA.n2127 3.4105
R14280 GNDA.n2140 GNDA.n2112 3.4105
R14281 GNDA.n2140 GNDA.n2128 3.4105
R14282 GNDA.n2140 GNDA.n2111 3.4105
R14283 GNDA.n2140 GNDA.n2129 3.4105
R14284 GNDA.n2140 GNDA.n2110 3.4105
R14285 GNDA.n2140 GNDA.n2130 3.4105
R14286 GNDA.n2140 GNDA.n2109 3.4105
R14287 GNDA.n2140 GNDA.n2131 3.4105
R14288 GNDA.n2140 GNDA.n2108 3.4105
R14289 GNDA.n2140 GNDA.n2132 3.4105
R14290 GNDA.n2140 GNDA.n2107 3.4105
R14291 GNDA.n2140 GNDA.n2133 3.4105
R14292 GNDA.n2140 GNDA.n2106 3.4105
R14293 GNDA.n2140 GNDA.n2134 3.4105
R14294 GNDA.n2226 GNDA.n2140 3.4105
R14295 GNDA.n2224 GNDA.n2211 3.4105
R14296 GNDA.n2211 GNDA.n2119 3.4105
R14297 GNDA.n2211 GNDA.n2121 3.4105
R14298 GNDA.n2211 GNDA.n2118 3.4105
R14299 GNDA.n2211 GNDA.n2122 3.4105
R14300 GNDA.n2211 GNDA.n2117 3.4105
R14301 GNDA.n2211 GNDA.n2123 3.4105
R14302 GNDA.n2211 GNDA.n2116 3.4105
R14303 GNDA.n2211 GNDA.n2124 3.4105
R14304 GNDA.n2211 GNDA.n2115 3.4105
R14305 GNDA.n2211 GNDA.n2125 3.4105
R14306 GNDA.n2211 GNDA.n2114 3.4105
R14307 GNDA.n2211 GNDA.n2126 3.4105
R14308 GNDA.n2211 GNDA.n2113 3.4105
R14309 GNDA.n2211 GNDA.n2127 3.4105
R14310 GNDA.n2211 GNDA.n2112 3.4105
R14311 GNDA.n2211 GNDA.n2128 3.4105
R14312 GNDA.n2211 GNDA.n2111 3.4105
R14313 GNDA.n2211 GNDA.n2129 3.4105
R14314 GNDA.n2211 GNDA.n2110 3.4105
R14315 GNDA.n2211 GNDA.n2130 3.4105
R14316 GNDA.n2211 GNDA.n2109 3.4105
R14317 GNDA.n2211 GNDA.n2131 3.4105
R14318 GNDA.n2211 GNDA.n2108 3.4105
R14319 GNDA.n2211 GNDA.n2132 3.4105
R14320 GNDA.n2211 GNDA.n2107 3.4105
R14321 GNDA.n2211 GNDA.n2133 3.4105
R14322 GNDA.n2211 GNDA.n2106 3.4105
R14323 GNDA.n2211 GNDA.n2134 3.4105
R14324 GNDA.n2226 GNDA.n2211 3.4105
R14325 GNDA.n2224 GNDA.n2139 3.4105
R14326 GNDA.n2139 GNDA.n2119 3.4105
R14327 GNDA.n2139 GNDA.n2121 3.4105
R14328 GNDA.n2139 GNDA.n2118 3.4105
R14329 GNDA.n2139 GNDA.n2122 3.4105
R14330 GNDA.n2139 GNDA.n2117 3.4105
R14331 GNDA.n2139 GNDA.n2123 3.4105
R14332 GNDA.n2139 GNDA.n2116 3.4105
R14333 GNDA.n2139 GNDA.n2124 3.4105
R14334 GNDA.n2139 GNDA.n2115 3.4105
R14335 GNDA.n2139 GNDA.n2125 3.4105
R14336 GNDA.n2139 GNDA.n2114 3.4105
R14337 GNDA.n2139 GNDA.n2126 3.4105
R14338 GNDA.n2139 GNDA.n2113 3.4105
R14339 GNDA.n2139 GNDA.n2127 3.4105
R14340 GNDA.n2139 GNDA.n2112 3.4105
R14341 GNDA.n2139 GNDA.n2128 3.4105
R14342 GNDA.n2139 GNDA.n2111 3.4105
R14343 GNDA.n2139 GNDA.n2129 3.4105
R14344 GNDA.n2139 GNDA.n2110 3.4105
R14345 GNDA.n2139 GNDA.n2130 3.4105
R14346 GNDA.n2139 GNDA.n2109 3.4105
R14347 GNDA.n2139 GNDA.n2131 3.4105
R14348 GNDA.n2139 GNDA.n2108 3.4105
R14349 GNDA.n2139 GNDA.n2132 3.4105
R14350 GNDA.n2139 GNDA.n2107 3.4105
R14351 GNDA.n2139 GNDA.n2133 3.4105
R14352 GNDA.n2139 GNDA.n2106 3.4105
R14353 GNDA.n2139 GNDA.n2134 3.4105
R14354 GNDA.n2226 GNDA.n2139 3.4105
R14355 GNDA.n2224 GNDA.n2214 3.4105
R14356 GNDA.n2214 GNDA.n2119 3.4105
R14357 GNDA.n2214 GNDA.n2121 3.4105
R14358 GNDA.n2214 GNDA.n2118 3.4105
R14359 GNDA.n2214 GNDA.n2122 3.4105
R14360 GNDA.n2214 GNDA.n2117 3.4105
R14361 GNDA.n2214 GNDA.n2123 3.4105
R14362 GNDA.n2214 GNDA.n2116 3.4105
R14363 GNDA.n2214 GNDA.n2124 3.4105
R14364 GNDA.n2214 GNDA.n2115 3.4105
R14365 GNDA.n2214 GNDA.n2125 3.4105
R14366 GNDA.n2214 GNDA.n2114 3.4105
R14367 GNDA.n2214 GNDA.n2126 3.4105
R14368 GNDA.n2214 GNDA.n2113 3.4105
R14369 GNDA.n2214 GNDA.n2127 3.4105
R14370 GNDA.n2214 GNDA.n2112 3.4105
R14371 GNDA.n2214 GNDA.n2128 3.4105
R14372 GNDA.n2214 GNDA.n2111 3.4105
R14373 GNDA.n2214 GNDA.n2129 3.4105
R14374 GNDA.n2214 GNDA.n2110 3.4105
R14375 GNDA.n2214 GNDA.n2130 3.4105
R14376 GNDA.n2214 GNDA.n2109 3.4105
R14377 GNDA.n2214 GNDA.n2131 3.4105
R14378 GNDA.n2214 GNDA.n2108 3.4105
R14379 GNDA.n2214 GNDA.n2132 3.4105
R14380 GNDA.n2214 GNDA.n2107 3.4105
R14381 GNDA.n2214 GNDA.n2133 3.4105
R14382 GNDA.n2214 GNDA.n2106 3.4105
R14383 GNDA.n2214 GNDA.n2134 3.4105
R14384 GNDA.n2226 GNDA.n2214 3.4105
R14385 GNDA.n2224 GNDA.n2138 3.4105
R14386 GNDA.n2138 GNDA.n2119 3.4105
R14387 GNDA.n2138 GNDA.n2121 3.4105
R14388 GNDA.n2138 GNDA.n2118 3.4105
R14389 GNDA.n2138 GNDA.n2122 3.4105
R14390 GNDA.n2138 GNDA.n2117 3.4105
R14391 GNDA.n2138 GNDA.n2123 3.4105
R14392 GNDA.n2138 GNDA.n2116 3.4105
R14393 GNDA.n2138 GNDA.n2124 3.4105
R14394 GNDA.n2138 GNDA.n2115 3.4105
R14395 GNDA.n2138 GNDA.n2125 3.4105
R14396 GNDA.n2138 GNDA.n2114 3.4105
R14397 GNDA.n2138 GNDA.n2126 3.4105
R14398 GNDA.n2138 GNDA.n2113 3.4105
R14399 GNDA.n2138 GNDA.n2127 3.4105
R14400 GNDA.n2138 GNDA.n2112 3.4105
R14401 GNDA.n2138 GNDA.n2128 3.4105
R14402 GNDA.n2138 GNDA.n2111 3.4105
R14403 GNDA.n2138 GNDA.n2129 3.4105
R14404 GNDA.n2138 GNDA.n2110 3.4105
R14405 GNDA.n2138 GNDA.n2130 3.4105
R14406 GNDA.n2138 GNDA.n2109 3.4105
R14407 GNDA.n2138 GNDA.n2131 3.4105
R14408 GNDA.n2138 GNDA.n2108 3.4105
R14409 GNDA.n2138 GNDA.n2132 3.4105
R14410 GNDA.n2138 GNDA.n2107 3.4105
R14411 GNDA.n2138 GNDA.n2133 3.4105
R14412 GNDA.n2138 GNDA.n2106 3.4105
R14413 GNDA.n2138 GNDA.n2134 3.4105
R14414 GNDA.n2226 GNDA.n2138 3.4105
R14415 GNDA.n2224 GNDA.n2217 3.4105
R14416 GNDA.n2217 GNDA.n2119 3.4105
R14417 GNDA.n2217 GNDA.n2121 3.4105
R14418 GNDA.n2217 GNDA.n2118 3.4105
R14419 GNDA.n2217 GNDA.n2122 3.4105
R14420 GNDA.n2217 GNDA.n2117 3.4105
R14421 GNDA.n2217 GNDA.n2123 3.4105
R14422 GNDA.n2217 GNDA.n2116 3.4105
R14423 GNDA.n2217 GNDA.n2124 3.4105
R14424 GNDA.n2217 GNDA.n2115 3.4105
R14425 GNDA.n2217 GNDA.n2125 3.4105
R14426 GNDA.n2217 GNDA.n2114 3.4105
R14427 GNDA.n2217 GNDA.n2126 3.4105
R14428 GNDA.n2217 GNDA.n2113 3.4105
R14429 GNDA.n2217 GNDA.n2127 3.4105
R14430 GNDA.n2217 GNDA.n2112 3.4105
R14431 GNDA.n2217 GNDA.n2128 3.4105
R14432 GNDA.n2217 GNDA.n2111 3.4105
R14433 GNDA.n2217 GNDA.n2129 3.4105
R14434 GNDA.n2217 GNDA.n2110 3.4105
R14435 GNDA.n2217 GNDA.n2130 3.4105
R14436 GNDA.n2217 GNDA.n2109 3.4105
R14437 GNDA.n2217 GNDA.n2131 3.4105
R14438 GNDA.n2217 GNDA.n2108 3.4105
R14439 GNDA.n2217 GNDA.n2132 3.4105
R14440 GNDA.n2217 GNDA.n2107 3.4105
R14441 GNDA.n2217 GNDA.n2133 3.4105
R14442 GNDA.n2217 GNDA.n2106 3.4105
R14443 GNDA.n2217 GNDA.n2134 3.4105
R14444 GNDA.n2226 GNDA.n2217 3.4105
R14445 GNDA.n2224 GNDA.n2137 3.4105
R14446 GNDA.n2137 GNDA.n2119 3.4105
R14447 GNDA.n2137 GNDA.n2121 3.4105
R14448 GNDA.n2137 GNDA.n2118 3.4105
R14449 GNDA.n2137 GNDA.n2122 3.4105
R14450 GNDA.n2137 GNDA.n2117 3.4105
R14451 GNDA.n2137 GNDA.n2123 3.4105
R14452 GNDA.n2137 GNDA.n2116 3.4105
R14453 GNDA.n2137 GNDA.n2124 3.4105
R14454 GNDA.n2137 GNDA.n2115 3.4105
R14455 GNDA.n2137 GNDA.n2125 3.4105
R14456 GNDA.n2137 GNDA.n2114 3.4105
R14457 GNDA.n2137 GNDA.n2126 3.4105
R14458 GNDA.n2137 GNDA.n2113 3.4105
R14459 GNDA.n2137 GNDA.n2127 3.4105
R14460 GNDA.n2137 GNDA.n2112 3.4105
R14461 GNDA.n2137 GNDA.n2128 3.4105
R14462 GNDA.n2137 GNDA.n2111 3.4105
R14463 GNDA.n2137 GNDA.n2129 3.4105
R14464 GNDA.n2137 GNDA.n2110 3.4105
R14465 GNDA.n2137 GNDA.n2130 3.4105
R14466 GNDA.n2137 GNDA.n2109 3.4105
R14467 GNDA.n2137 GNDA.n2131 3.4105
R14468 GNDA.n2137 GNDA.n2108 3.4105
R14469 GNDA.n2137 GNDA.n2132 3.4105
R14470 GNDA.n2137 GNDA.n2107 3.4105
R14471 GNDA.n2137 GNDA.n2133 3.4105
R14472 GNDA.n2137 GNDA.n2106 3.4105
R14473 GNDA.n2137 GNDA.n2134 3.4105
R14474 GNDA.n2226 GNDA.n2137 3.4105
R14475 GNDA.n2224 GNDA.n2220 3.4105
R14476 GNDA.n2220 GNDA.n2119 3.4105
R14477 GNDA.n2220 GNDA.n2121 3.4105
R14478 GNDA.n2220 GNDA.n2118 3.4105
R14479 GNDA.n2220 GNDA.n2122 3.4105
R14480 GNDA.n2220 GNDA.n2117 3.4105
R14481 GNDA.n2220 GNDA.n2123 3.4105
R14482 GNDA.n2220 GNDA.n2116 3.4105
R14483 GNDA.n2220 GNDA.n2124 3.4105
R14484 GNDA.n2220 GNDA.n2115 3.4105
R14485 GNDA.n2220 GNDA.n2125 3.4105
R14486 GNDA.n2220 GNDA.n2114 3.4105
R14487 GNDA.n2220 GNDA.n2126 3.4105
R14488 GNDA.n2220 GNDA.n2113 3.4105
R14489 GNDA.n2220 GNDA.n2127 3.4105
R14490 GNDA.n2220 GNDA.n2112 3.4105
R14491 GNDA.n2220 GNDA.n2128 3.4105
R14492 GNDA.n2220 GNDA.n2111 3.4105
R14493 GNDA.n2220 GNDA.n2129 3.4105
R14494 GNDA.n2220 GNDA.n2110 3.4105
R14495 GNDA.n2220 GNDA.n2130 3.4105
R14496 GNDA.n2220 GNDA.n2109 3.4105
R14497 GNDA.n2220 GNDA.n2131 3.4105
R14498 GNDA.n2220 GNDA.n2108 3.4105
R14499 GNDA.n2220 GNDA.n2132 3.4105
R14500 GNDA.n2220 GNDA.n2107 3.4105
R14501 GNDA.n2220 GNDA.n2133 3.4105
R14502 GNDA.n2220 GNDA.n2106 3.4105
R14503 GNDA.n2220 GNDA.n2134 3.4105
R14504 GNDA.n2226 GNDA.n2220 3.4105
R14505 GNDA.n2224 GNDA.n2136 3.4105
R14506 GNDA.n2136 GNDA.n2119 3.4105
R14507 GNDA.n2136 GNDA.n2121 3.4105
R14508 GNDA.n2136 GNDA.n2118 3.4105
R14509 GNDA.n2136 GNDA.n2122 3.4105
R14510 GNDA.n2136 GNDA.n2117 3.4105
R14511 GNDA.n2136 GNDA.n2123 3.4105
R14512 GNDA.n2136 GNDA.n2116 3.4105
R14513 GNDA.n2136 GNDA.n2124 3.4105
R14514 GNDA.n2136 GNDA.n2115 3.4105
R14515 GNDA.n2136 GNDA.n2125 3.4105
R14516 GNDA.n2136 GNDA.n2114 3.4105
R14517 GNDA.n2136 GNDA.n2126 3.4105
R14518 GNDA.n2136 GNDA.n2113 3.4105
R14519 GNDA.n2136 GNDA.n2127 3.4105
R14520 GNDA.n2136 GNDA.n2112 3.4105
R14521 GNDA.n2136 GNDA.n2128 3.4105
R14522 GNDA.n2136 GNDA.n2111 3.4105
R14523 GNDA.n2136 GNDA.n2129 3.4105
R14524 GNDA.n2136 GNDA.n2110 3.4105
R14525 GNDA.n2136 GNDA.n2130 3.4105
R14526 GNDA.n2136 GNDA.n2109 3.4105
R14527 GNDA.n2136 GNDA.n2131 3.4105
R14528 GNDA.n2136 GNDA.n2108 3.4105
R14529 GNDA.n2136 GNDA.n2132 3.4105
R14530 GNDA.n2136 GNDA.n2107 3.4105
R14531 GNDA.n2136 GNDA.n2133 3.4105
R14532 GNDA.n2136 GNDA.n2106 3.4105
R14533 GNDA.n2136 GNDA.n2134 3.4105
R14534 GNDA.n2226 GNDA.n2136 3.4105
R14535 GNDA.n2225 GNDA.n2224 3.4105
R14536 GNDA.n2225 GNDA.n2119 3.4105
R14537 GNDA.n2225 GNDA.n2121 3.4105
R14538 GNDA.n2225 GNDA.n2118 3.4105
R14539 GNDA.n2225 GNDA.n2122 3.4105
R14540 GNDA.n2225 GNDA.n2117 3.4105
R14541 GNDA.n2225 GNDA.n2123 3.4105
R14542 GNDA.n2225 GNDA.n2116 3.4105
R14543 GNDA.n2225 GNDA.n2124 3.4105
R14544 GNDA.n2225 GNDA.n2115 3.4105
R14545 GNDA.n2225 GNDA.n2125 3.4105
R14546 GNDA.n2225 GNDA.n2114 3.4105
R14547 GNDA.n2225 GNDA.n2126 3.4105
R14548 GNDA.n2225 GNDA.n2113 3.4105
R14549 GNDA.n2225 GNDA.n2127 3.4105
R14550 GNDA.n2225 GNDA.n2112 3.4105
R14551 GNDA.n2225 GNDA.n2128 3.4105
R14552 GNDA.n2225 GNDA.n2111 3.4105
R14553 GNDA.n2225 GNDA.n2129 3.4105
R14554 GNDA.n2225 GNDA.n2110 3.4105
R14555 GNDA.n2225 GNDA.n2130 3.4105
R14556 GNDA.n2225 GNDA.n2109 3.4105
R14557 GNDA.n2225 GNDA.n2131 3.4105
R14558 GNDA.n2225 GNDA.n2108 3.4105
R14559 GNDA.n2225 GNDA.n2132 3.4105
R14560 GNDA.n2225 GNDA.n2107 3.4105
R14561 GNDA.n2225 GNDA.n2133 3.4105
R14562 GNDA.n2225 GNDA.n2106 3.4105
R14563 GNDA.n2225 GNDA.n2134 3.4105
R14564 GNDA.n2226 GNDA.n2225 3.4105
R14565 GNDA.n2224 GNDA.n2135 3.4105
R14566 GNDA.n2135 GNDA.n2119 3.4105
R14567 GNDA.n2135 GNDA.n2121 3.4105
R14568 GNDA.n2135 GNDA.n2118 3.4105
R14569 GNDA.n2135 GNDA.n2122 3.4105
R14570 GNDA.n2135 GNDA.n2117 3.4105
R14571 GNDA.n2135 GNDA.n2123 3.4105
R14572 GNDA.n2135 GNDA.n2116 3.4105
R14573 GNDA.n2135 GNDA.n2124 3.4105
R14574 GNDA.n2135 GNDA.n2115 3.4105
R14575 GNDA.n2135 GNDA.n2125 3.4105
R14576 GNDA.n2135 GNDA.n2114 3.4105
R14577 GNDA.n2135 GNDA.n2126 3.4105
R14578 GNDA.n2135 GNDA.n2113 3.4105
R14579 GNDA.n2135 GNDA.n2127 3.4105
R14580 GNDA.n2135 GNDA.n2112 3.4105
R14581 GNDA.n2135 GNDA.n2128 3.4105
R14582 GNDA.n2135 GNDA.n2111 3.4105
R14583 GNDA.n2135 GNDA.n2129 3.4105
R14584 GNDA.n2135 GNDA.n2110 3.4105
R14585 GNDA.n2135 GNDA.n2130 3.4105
R14586 GNDA.n2135 GNDA.n2109 3.4105
R14587 GNDA.n2135 GNDA.n2131 3.4105
R14588 GNDA.n2135 GNDA.n2108 3.4105
R14589 GNDA.n2135 GNDA.n2132 3.4105
R14590 GNDA.n2135 GNDA.n2107 3.4105
R14591 GNDA.n2135 GNDA.n2133 3.4105
R14592 GNDA.n2135 GNDA.n2106 3.4105
R14593 GNDA.n2135 GNDA.n2134 3.4105
R14594 GNDA.n2226 GNDA.n2135 3.4105
R14595 GNDA.n2227 GNDA.n2119 3.4105
R14596 GNDA.n2227 GNDA.n2121 3.4105
R14597 GNDA.n2227 GNDA.n2118 3.4105
R14598 GNDA.n2227 GNDA.n2122 3.4105
R14599 GNDA.n2227 GNDA.n2117 3.4105
R14600 GNDA.n2227 GNDA.n2123 3.4105
R14601 GNDA.n2227 GNDA.n2116 3.4105
R14602 GNDA.n2227 GNDA.n2124 3.4105
R14603 GNDA.n2227 GNDA.n2115 3.4105
R14604 GNDA.n2227 GNDA.n2125 3.4105
R14605 GNDA.n2227 GNDA.n2114 3.4105
R14606 GNDA.n2227 GNDA.n2126 3.4105
R14607 GNDA.n2227 GNDA.n2113 3.4105
R14608 GNDA.n2227 GNDA.n2127 3.4105
R14609 GNDA.n2227 GNDA.n2112 3.4105
R14610 GNDA.n2227 GNDA.n2128 3.4105
R14611 GNDA.n2227 GNDA.n2111 3.4105
R14612 GNDA.n2227 GNDA.n2129 3.4105
R14613 GNDA.n2227 GNDA.n2110 3.4105
R14614 GNDA.n2227 GNDA.n2130 3.4105
R14615 GNDA.n2227 GNDA.n2109 3.4105
R14616 GNDA.n2227 GNDA.n2131 3.4105
R14617 GNDA.n2227 GNDA.n2108 3.4105
R14618 GNDA.n2227 GNDA.n2132 3.4105
R14619 GNDA.n2227 GNDA.n2107 3.4105
R14620 GNDA.n2227 GNDA.n2133 3.4105
R14621 GNDA.n2227 GNDA.n2106 3.4105
R14622 GNDA.n2227 GNDA.n2134 3.4105
R14623 GNDA.n2227 GNDA.n2226 3.4105
R14624 GNDA.n2356 GNDA.n2249 3.4105
R14625 GNDA.n2352 GNDA.n2249 3.4105
R14626 GNDA.n2354 GNDA.n2249 3.4105
R14627 GNDA.n2353 GNDA.n2352 3.4105
R14628 GNDA.n2354 GNDA.n2353 3.4105
R14629 GNDA.n2356 GNDA.n1966 3.4105
R14630 GNDA.n2280 GNDA.n1966 3.4105
R14631 GNDA.n2278 GNDA.n1966 3.4105
R14632 GNDA.n2282 GNDA.n1966 3.4105
R14633 GNDA.n2277 GNDA.n1966 3.4105
R14634 GNDA.n2284 GNDA.n1966 3.4105
R14635 GNDA.n2276 GNDA.n1966 3.4105
R14636 GNDA.n2286 GNDA.n1966 3.4105
R14637 GNDA.n2275 GNDA.n1966 3.4105
R14638 GNDA.n2288 GNDA.n1966 3.4105
R14639 GNDA.n2274 GNDA.n1966 3.4105
R14640 GNDA.n2290 GNDA.n1966 3.4105
R14641 GNDA.n2273 GNDA.n1966 3.4105
R14642 GNDA.n2292 GNDA.n1966 3.4105
R14643 GNDA.n2272 GNDA.n1966 3.4105
R14644 GNDA.n2294 GNDA.n1966 3.4105
R14645 GNDA.n2271 GNDA.n1966 3.4105
R14646 GNDA.n2296 GNDA.n1966 3.4105
R14647 GNDA.n2270 GNDA.n1966 3.4105
R14648 GNDA.n2298 GNDA.n1966 3.4105
R14649 GNDA.n2269 GNDA.n1966 3.4105
R14650 GNDA.n2300 GNDA.n1966 3.4105
R14651 GNDA.n2268 GNDA.n1966 3.4105
R14652 GNDA.n2302 GNDA.n1966 3.4105
R14653 GNDA.n2267 GNDA.n1966 3.4105
R14654 GNDA.n2304 GNDA.n1966 3.4105
R14655 GNDA.n2266 GNDA.n1966 3.4105
R14656 GNDA.n2305 GNDA.n1966 3.4105
R14657 GNDA.n2352 GNDA.n1966 3.4105
R14658 GNDA.n2354 GNDA.n1966 3.4105
R14659 GNDA.n2356 GNDA.n2250 3.4105
R14660 GNDA.n2280 GNDA.n2250 3.4105
R14661 GNDA.n2278 GNDA.n2250 3.4105
R14662 GNDA.n2282 GNDA.n2250 3.4105
R14663 GNDA.n2277 GNDA.n2250 3.4105
R14664 GNDA.n2284 GNDA.n2250 3.4105
R14665 GNDA.n2276 GNDA.n2250 3.4105
R14666 GNDA.n2286 GNDA.n2250 3.4105
R14667 GNDA.n2275 GNDA.n2250 3.4105
R14668 GNDA.n2288 GNDA.n2250 3.4105
R14669 GNDA.n2274 GNDA.n2250 3.4105
R14670 GNDA.n2290 GNDA.n2250 3.4105
R14671 GNDA.n2273 GNDA.n2250 3.4105
R14672 GNDA.n2292 GNDA.n2250 3.4105
R14673 GNDA.n2272 GNDA.n2250 3.4105
R14674 GNDA.n2294 GNDA.n2250 3.4105
R14675 GNDA.n2271 GNDA.n2250 3.4105
R14676 GNDA.n2296 GNDA.n2250 3.4105
R14677 GNDA.n2270 GNDA.n2250 3.4105
R14678 GNDA.n2298 GNDA.n2250 3.4105
R14679 GNDA.n2269 GNDA.n2250 3.4105
R14680 GNDA.n2300 GNDA.n2250 3.4105
R14681 GNDA.n2268 GNDA.n2250 3.4105
R14682 GNDA.n2302 GNDA.n2250 3.4105
R14683 GNDA.n2267 GNDA.n2250 3.4105
R14684 GNDA.n2304 GNDA.n2250 3.4105
R14685 GNDA.n2266 GNDA.n2250 3.4105
R14686 GNDA.n2305 GNDA.n2250 3.4105
R14687 GNDA.n2352 GNDA.n2250 3.4105
R14688 GNDA.n2354 GNDA.n2250 3.4105
R14689 GNDA.n2356 GNDA.n1965 3.4105
R14690 GNDA.n2280 GNDA.n1965 3.4105
R14691 GNDA.n2278 GNDA.n1965 3.4105
R14692 GNDA.n2282 GNDA.n1965 3.4105
R14693 GNDA.n2277 GNDA.n1965 3.4105
R14694 GNDA.n2284 GNDA.n1965 3.4105
R14695 GNDA.n2276 GNDA.n1965 3.4105
R14696 GNDA.n2286 GNDA.n1965 3.4105
R14697 GNDA.n2275 GNDA.n1965 3.4105
R14698 GNDA.n2288 GNDA.n1965 3.4105
R14699 GNDA.n2274 GNDA.n1965 3.4105
R14700 GNDA.n2290 GNDA.n1965 3.4105
R14701 GNDA.n2273 GNDA.n1965 3.4105
R14702 GNDA.n2292 GNDA.n1965 3.4105
R14703 GNDA.n2272 GNDA.n1965 3.4105
R14704 GNDA.n2294 GNDA.n1965 3.4105
R14705 GNDA.n2271 GNDA.n1965 3.4105
R14706 GNDA.n2296 GNDA.n1965 3.4105
R14707 GNDA.n2270 GNDA.n1965 3.4105
R14708 GNDA.n2298 GNDA.n1965 3.4105
R14709 GNDA.n2269 GNDA.n1965 3.4105
R14710 GNDA.n2300 GNDA.n1965 3.4105
R14711 GNDA.n2268 GNDA.n1965 3.4105
R14712 GNDA.n2302 GNDA.n1965 3.4105
R14713 GNDA.n2267 GNDA.n1965 3.4105
R14714 GNDA.n2304 GNDA.n1965 3.4105
R14715 GNDA.n2266 GNDA.n1965 3.4105
R14716 GNDA.n2305 GNDA.n1965 3.4105
R14717 GNDA.n2352 GNDA.n1965 3.4105
R14718 GNDA.n2354 GNDA.n1965 3.4105
R14719 GNDA.n2356 GNDA.n2251 3.4105
R14720 GNDA.n2280 GNDA.n2251 3.4105
R14721 GNDA.n2278 GNDA.n2251 3.4105
R14722 GNDA.n2282 GNDA.n2251 3.4105
R14723 GNDA.n2277 GNDA.n2251 3.4105
R14724 GNDA.n2284 GNDA.n2251 3.4105
R14725 GNDA.n2276 GNDA.n2251 3.4105
R14726 GNDA.n2286 GNDA.n2251 3.4105
R14727 GNDA.n2275 GNDA.n2251 3.4105
R14728 GNDA.n2288 GNDA.n2251 3.4105
R14729 GNDA.n2274 GNDA.n2251 3.4105
R14730 GNDA.n2290 GNDA.n2251 3.4105
R14731 GNDA.n2273 GNDA.n2251 3.4105
R14732 GNDA.n2292 GNDA.n2251 3.4105
R14733 GNDA.n2272 GNDA.n2251 3.4105
R14734 GNDA.n2294 GNDA.n2251 3.4105
R14735 GNDA.n2271 GNDA.n2251 3.4105
R14736 GNDA.n2296 GNDA.n2251 3.4105
R14737 GNDA.n2270 GNDA.n2251 3.4105
R14738 GNDA.n2298 GNDA.n2251 3.4105
R14739 GNDA.n2269 GNDA.n2251 3.4105
R14740 GNDA.n2300 GNDA.n2251 3.4105
R14741 GNDA.n2268 GNDA.n2251 3.4105
R14742 GNDA.n2302 GNDA.n2251 3.4105
R14743 GNDA.n2267 GNDA.n2251 3.4105
R14744 GNDA.n2304 GNDA.n2251 3.4105
R14745 GNDA.n2266 GNDA.n2251 3.4105
R14746 GNDA.n2305 GNDA.n2251 3.4105
R14747 GNDA.n2352 GNDA.n2251 3.4105
R14748 GNDA.n2354 GNDA.n2251 3.4105
R14749 GNDA.n2356 GNDA.n1964 3.4105
R14750 GNDA.n2280 GNDA.n1964 3.4105
R14751 GNDA.n2278 GNDA.n1964 3.4105
R14752 GNDA.n2282 GNDA.n1964 3.4105
R14753 GNDA.n2277 GNDA.n1964 3.4105
R14754 GNDA.n2284 GNDA.n1964 3.4105
R14755 GNDA.n2276 GNDA.n1964 3.4105
R14756 GNDA.n2286 GNDA.n1964 3.4105
R14757 GNDA.n2275 GNDA.n1964 3.4105
R14758 GNDA.n2288 GNDA.n1964 3.4105
R14759 GNDA.n2274 GNDA.n1964 3.4105
R14760 GNDA.n2290 GNDA.n1964 3.4105
R14761 GNDA.n2273 GNDA.n1964 3.4105
R14762 GNDA.n2292 GNDA.n1964 3.4105
R14763 GNDA.n2272 GNDA.n1964 3.4105
R14764 GNDA.n2294 GNDA.n1964 3.4105
R14765 GNDA.n2271 GNDA.n1964 3.4105
R14766 GNDA.n2296 GNDA.n1964 3.4105
R14767 GNDA.n2270 GNDA.n1964 3.4105
R14768 GNDA.n2298 GNDA.n1964 3.4105
R14769 GNDA.n2269 GNDA.n1964 3.4105
R14770 GNDA.n2300 GNDA.n1964 3.4105
R14771 GNDA.n2268 GNDA.n1964 3.4105
R14772 GNDA.n2302 GNDA.n1964 3.4105
R14773 GNDA.n2267 GNDA.n1964 3.4105
R14774 GNDA.n2304 GNDA.n1964 3.4105
R14775 GNDA.n2266 GNDA.n1964 3.4105
R14776 GNDA.n2305 GNDA.n1964 3.4105
R14777 GNDA.n2352 GNDA.n1964 3.4105
R14778 GNDA.n2354 GNDA.n1964 3.4105
R14779 GNDA.n2356 GNDA.n2252 3.4105
R14780 GNDA.n2280 GNDA.n2252 3.4105
R14781 GNDA.n2278 GNDA.n2252 3.4105
R14782 GNDA.n2282 GNDA.n2252 3.4105
R14783 GNDA.n2277 GNDA.n2252 3.4105
R14784 GNDA.n2284 GNDA.n2252 3.4105
R14785 GNDA.n2276 GNDA.n2252 3.4105
R14786 GNDA.n2286 GNDA.n2252 3.4105
R14787 GNDA.n2275 GNDA.n2252 3.4105
R14788 GNDA.n2288 GNDA.n2252 3.4105
R14789 GNDA.n2274 GNDA.n2252 3.4105
R14790 GNDA.n2290 GNDA.n2252 3.4105
R14791 GNDA.n2273 GNDA.n2252 3.4105
R14792 GNDA.n2292 GNDA.n2252 3.4105
R14793 GNDA.n2272 GNDA.n2252 3.4105
R14794 GNDA.n2294 GNDA.n2252 3.4105
R14795 GNDA.n2271 GNDA.n2252 3.4105
R14796 GNDA.n2296 GNDA.n2252 3.4105
R14797 GNDA.n2270 GNDA.n2252 3.4105
R14798 GNDA.n2298 GNDA.n2252 3.4105
R14799 GNDA.n2269 GNDA.n2252 3.4105
R14800 GNDA.n2300 GNDA.n2252 3.4105
R14801 GNDA.n2268 GNDA.n2252 3.4105
R14802 GNDA.n2302 GNDA.n2252 3.4105
R14803 GNDA.n2267 GNDA.n2252 3.4105
R14804 GNDA.n2304 GNDA.n2252 3.4105
R14805 GNDA.n2266 GNDA.n2252 3.4105
R14806 GNDA.n2305 GNDA.n2252 3.4105
R14807 GNDA.n2352 GNDA.n2252 3.4105
R14808 GNDA.n2354 GNDA.n2252 3.4105
R14809 GNDA.n2356 GNDA.n1963 3.4105
R14810 GNDA.n2280 GNDA.n1963 3.4105
R14811 GNDA.n2278 GNDA.n1963 3.4105
R14812 GNDA.n2282 GNDA.n1963 3.4105
R14813 GNDA.n2277 GNDA.n1963 3.4105
R14814 GNDA.n2284 GNDA.n1963 3.4105
R14815 GNDA.n2276 GNDA.n1963 3.4105
R14816 GNDA.n2286 GNDA.n1963 3.4105
R14817 GNDA.n2275 GNDA.n1963 3.4105
R14818 GNDA.n2288 GNDA.n1963 3.4105
R14819 GNDA.n2274 GNDA.n1963 3.4105
R14820 GNDA.n2290 GNDA.n1963 3.4105
R14821 GNDA.n2273 GNDA.n1963 3.4105
R14822 GNDA.n2292 GNDA.n1963 3.4105
R14823 GNDA.n2272 GNDA.n1963 3.4105
R14824 GNDA.n2294 GNDA.n1963 3.4105
R14825 GNDA.n2271 GNDA.n1963 3.4105
R14826 GNDA.n2296 GNDA.n1963 3.4105
R14827 GNDA.n2270 GNDA.n1963 3.4105
R14828 GNDA.n2298 GNDA.n1963 3.4105
R14829 GNDA.n2269 GNDA.n1963 3.4105
R14830 GNDA.n2300 GNDA.n1963 3.4105
R14831 GNDA.n2268 GNDA.n1963 3.4105
R14832 GNDA.n2302 GNDA.n1963 3.4105
R14833 GNDA.n2267 GNDA.n1963 3.4105
R14834 GNDA.n2304 GNDA.n1963 3.4105
R14835 GNDA.n2266 GNDA.n1963 3.4105
R14836 GNDA.n2305 GNDA.n1963 3.4105
R14837 GNDA.n2352 GNDA.n1963 3.4105
R14838 GNDA.n2354 GNDA.n1963 3.4105
R14839 GNDA.n2356 GNDA.n2253 3.4105
R14840 GNDA.n2280 GNDA.n2253 3.4105
R14841 GNDA.n2278 GNDA.n2253 3.4105
R14842 GNDA.n2282 GNDA.n2253 3.4105
R14843 GNDA.n2277 GNDA.n2253 3.4105
R14844 GNDA.n2284 GNDA.n2253 3.4105
R14845 GNDA.n2276 GNDA.n2253 3.4105
R14846 GNDA.n2286 GNDA.n2253 3.4105
R14847 GNDA.n2275 GNDA.n2253 3.4105
R14848 GNDA.n2288 GNDA.n2253 3.4105
R14849 GNDA.n2274 GNDA.n2253 3.4105
R14850 GNDA.n2290 GNDA.n2253 3.4105
R14851 GNDA.n2273 GNDA.n2253 3.4105
R14852 GNDA.n2292 GNDA.n2253 3.4105
R14853 GNDA.n2272 GNDA.n2253 3.4105
R14854 GNDA.n2294 GNDA.n2253 3.4105
R14855 GNDA.n2271 GNDA.n2253 3.4105
R14856 GNDA.n2296 GNDA.n2253 3.4105
R14857 GNDA.n2270 GNDA.n2253 3.4105
R14858 GNDA.n2298 GNDA.n2253 3.4105
R14859 GNDA.n2269 GNDA.n2253 3.4105
R14860 GNDA.n2300 GNDA.n2253 3.4105
R14861 GNDA.n2268 GNDA.n2253 3.4105
R14862 GNDA.n2302 GNDA.n2253 3.4105
R14863 GNDA.n2267 GNDA.n2253 3.4105
R14864 GNDA.n2304 GNDA.n2253 3.4105
R14865 GNDA.n2266 GNDA.n2253 3.4105
R14866 GNDA.n2305 GNDA.n2253 3.4105
R14867 GNDA.n2352 GNDA.n2253 3.4105
R14868 GNDA.n2354 GNDA.n2253 3.4105
R14869 GNDA.n2356 GNDA.n1962 3.4105
R14870 GNDA.n2280 GNDA.n1962 3.4105
R14871 GNDA.n2278 GNDA.n1962 3.4105
R14872 GNDA.n2282 GNDA.n1962 3.4105
R14873 GNDA.n2277 GNDA.n1962 3.4105
R14874 GNDA.n2284 GNDA.n1962 3.4105
R14875 GNDA.n2276 GNDA.n1962 3.4105
R14876 GNDA.n2286 GNDA.n1962 3.4105
R14877 GNDA.n2275 GNDA.n1962 3.4105
R14878 GNDA.n2288 GNDA.n1962 3.4105
R14879 GNDA.n2274 GNDA.n1962 3.4105
R14880 GNDA.n2290 GNDA.n1962 3.4105
R14881 GNDA.n2273 GNDA.n1962 3.4105
R14882 GNDA.n2292 GNDA.n1962 3.4105
R14883 GNDA.n2272 GNDA.n1962 3.4105
R14884 GNDA.n2294 GNDA.n1962 3.4105
R14885 GNDA.n2271 GNDA.n1962 3.4105
R14886 GNDA.n2296 GNDA.n1962 3.4105
R14887 GNDA.n2270 GNDA.n1962 3.4105
R14888 GNDA.n2298 GNDA.n1962 3.4105
R14889 GNDA.n2269 GNDA.n1962 3.4105
R14890 GNDA.n2300 GNDA.n1962 3.4105
R14891 GNDA.n2268 GNDA.n1962 3.4105
R14892 GNDA.n2302 GNDA.n1962 3.4105
R14893 GNDA.n2267 GNDA.n1962 3.4105
R14894 GNDA.n2304 GNDA.n1962 3.4105
R14895 GNDA.n2266 GNDA.n1962 3.4105
R14896 GNDA.n2305 GNDA.n1962 3.4105
R14897 GNDA.n2352 GNDA.n1962 3.4105
R14898 GNDA.n2354 GNDA.n1962 3.4105
R14899 GNDA.n2356 GNDA.n2254 3.4105
R14900 GNDA.n2280 GNDA.n2254 3.4105
R14901 GNDA.n2278 GNDA.n2254 3.4105
R14902 GNDA.n2282 GNDA.n2254 3.4105
R14903 GNDA.n2277 GNDA.n2254 3.4105
R14904 GNDA.n2284 GNDA.n2254 3.4105
R14905 GNDA.n2276 GNDA.n2254 3.4105
R14906 GNDA.n2286 GNDA.n2254 3.4105
R14907 GNDA.n2275 GNDA.n2254 3.4105
R14908 GNDA.n2288 GNDA.n2254 3.4105
R14909 GNDA.n2274 GNDA.n2254 3.4105
R14910 GNDA.n2290 GNDA.n2254 3.4105
R14911 GNDA.n2273 GNDA.n2254 3.4105
R14912 GNDA.n2292 GNDA.n2254 3.4105
R14913 GNDA.n2272 GNDA.n2254 3.4105
R14914 GNDA.n2294 GNDA.n2254 3.4105
R14915 GNDA.n2271 GNDA.n2254 3.4105
R14916 GNDA.n2296 GNDA.n2254 3.4105
R14917 GNDA.n2270 GNDA.n2254 3.4105
R14918 GNDA.n2298 GNDA.n2254 3.4105
R14919 GNDA.n2269 GNDA.n2254 3.4105
R14920 GNDA.n2300 GNDA.n2254 3.4105
R14921 GNDA.n2268 GNDA.n2254 3.4105
R14922 GNDA.n2302 GNDA.n2254 3.4105
R14923 GNDA.n2267 GNDA.n2254 3.4105
R14924 GNDA.n2304 GNDA.n2254 3.4105
R14925 GNDA.n2266 GNDA.n2254 3.4105
R14926 GNDA.n2305 GNDA.n2254 3.4105
R14927 GNDA.n2352 GNDA.n2254 3.4105
R14928 GNDA.n2354 GNDA.n2254 3.4105
R14929 GNDA.n2356 GNDA.n1961 3.4105
R14930 GNDA.n2280 GNDA.n1961 3.4105
R14931 GNDA.n2278 GNDA.n1961 3.4105
R14932 GNDA.n2282 GNDA.n1961 3.4105
R14933 GNDA.n2277 GNDA.n1961 3.4105
R14934 GNDA.n2284 GNDA.n1961 3.4105
R14935 GNDA.n2276 GNDA.n1961 3.4105
R14936 GNDA.n2286 GNDA.n1961 3.4105
R14937 GNDA.n2275 GNDA.n1961 3.4105
R14938 GNDA.n2288 GNDA.n1961 3.4105
R14939 GNDA.n2274 GNDA.n1961 3.4105
R14940 GNDA.n2290 GNDA.n1961 3.4105
R14941 GNDA.n2273 GNDA.n1961 3.4105
R14942 GNDA.n2292 GNDA.n1961 3.4105
R14943 GNDA.n2272 GNDA.n1961 3.4105
R14944 GNDA.n2294 GNDA.n1961 3.4105
R14945 GNDA.n2271 GNDA.n1961 3.4105
R14946 GNDA.n2296 GNDA.n1961 3.4105
R14947 GNDA.n2270 GNDA.n1961 3.4105
R14948 GNDA.n2298 GNDA.n1961 3.4105
R14949 GNDA.n2269 GNDA.n1961 3.4105
R14950 GNDA.n2300 GNDA.n1961 3.4105
R14951 GNDA.n2268 GNDA.n1961 3.4105
R14952 GNDA.n2302 GNDA.n1961 3.4105
R14953 GNDA.n2267 GNDA.n1961 3.4105
R14954 GNDA.n2304 GNDA.n1961 3.4105
R14955 GNDA.n2266 GNDA.n1961 3.4105
R14956 GNDA.n2305 GNDA.n1961 3.4105
R14957 GNDA.n2352 GNDA.n1961 3.4105
R14958 GNDA.n2354 GNDA.n1961 3.4105
R14959 GNDA.n2356 GNDA.n2255 3.4105
R14960 GNDA.n2280 GNDA.n2255 3.4105
R14961 GNDA.n2278 GNDA.n2255 3.4105
R14962 GNDA.n2282 GNDA.n2255 3.4105
R14963 GNDA.n2277 GNDA.n2255 3.4105
R14964 GNDA.n2284 GNDA.n2255 3.4105
R14965 GNDA.n2276 GNDA.n2255 3.4105
R14966 GNDA.n2286 GNDA.n2255 3.4105
R14967 GNDA.n2275 GNDA.n2255 3.4105
R14968 GNDA.n2288 GNDA.n2255 3.4105
R14969 GNDA.n2274 GNDA.n2255 3.4105
R14970 GNDA.n2290 GNDA.n2255 3.4105
R14971 GNDA.n2273 GNDA.n2255 3.4105
R14972 GNDA.n2292 GNDA.n2255 3.4105
R14973 GNDA.n2272 GNDA.n2255 3.4105
R14974 GNDA.n2294 GNDA.n2255 3.4105
R14975 GNDA.n2271 GNDA.n2255 3.4105
R14976 GNDA.n2296 GNDA.n2255 3.4105
R14977 GNDA.n2270 GNDA.n2255 3.4105
R14978 GNDA.n2298 GNDA.n2255 3.4105
R14979 GNDA.n2269 GNDA.n2255 3.4105
R14980 GNDA.n2300 GNDA.n2255 3.4105
R14981 GNDA.n2268 GNDA.n2255 3.4105
R14982 GNDA.n2302 GNDA.n2255 3.4105
R14983 GNDA.n2267 GNDA.n2255 3.4105
R14984 GNDA.n2304 GNDA.n2255 3.4105
R14985 GNDA.n2266 GNDA.n2255 3.4105
R14986 GNDA.n2305 GNDA.n2255 3.4105
R14987 GNDA.n2352 GNDA.n2255 3.4105
R14988 GNDA.n2354 GNDA.n2255 3.4105
R14989 GNDA.n2356 GNDA.n1960 3.4105
R14990 GNDA.n2280 GNDA.n1960 3.4105
R14991 GNDA.n2278 GNDA.n1960 3.4105
R14992 GNDA.n2282 GNDA.n1960 3.4105
R14993 GNDA.n2277 GNDA.n1960 3.4105
R14994 GNDA.n2284 GNDA.n1960 3.4105
R14995 GNDA.n2276 GNDA.n1960 3.4105
R14996 GNDA.n2286 GNDA.n1960 3.4105
R14997 GNDA.n2275 GNDA.n1960 3.4105
R14998 GNDA.n2288 GNDA.n1960 3.4105
R14999 GNDA.n2274 GNDA.n1960 3.4105
R15000 GNDA.n2290 GNDA.n1960 3.4105
R15001 GNDA.n2273 GNDA.n1960 3.4105
R15002 GNDA.n2292 GNDA.n1960 3.4105
R15003 GNDA.n2272 GNDA.n1960 3.4105
R15004 GNDA.n2294 GNDA.n1960 3.4105
R15005 GNDA.n2271 GNDA.n1960 3.4105
R15006 GNDA.n2296 GNDA.n1960 3.4105
R15007 GNDA.n2270 GNDA.n1960 3.4105
R15008 GNDA.n2298 GNDA.n1960 3.4105
R15009 GNDA.n2269 GNDA.n1960 3.4105
R15010 GNDA.n2300 GNDA.n1960 3.4105
R15011 GNDA.n2268 GNDA.n1960 3.4105
R15012 GNDA.n2302 GNDA.n1960 3.4105
R15013 GNDA.n2267 GNDA.n1960 3.4105
R15014 GNDA.n2304 GNDA.n1960 3.4105
R15015 GNDA.n2266 GNDA.n1960 3.4105
R15016 GNDA.n2305 GNDA.n1960 3.4105
R15017 GNDA.n2352 GNDA.n1960 3.4105
R15018 GNDA.n2354 GNDA.n1960 3.4105
R15019 GNDA.n2356 GNDA.n2256 3.4105
R15020 GNDA.n2280 GNDA.n2256 3.4105
R15021 GNDA.n2278 GNDA.n2256 3.4105
R15022 GNDA.n2282 GNDA.n2256 3.4105
R15023 GNDA.n2277 GNDA.n2256 3.4105
R15024 GNDA.n2284 GNDA.n2256 3.4105
R15025 GNDA.n2276 GNDA.n2256 3.4105
R15026 GNDA.n2286 GNDA.n2256 3.4105
R15027 GNDA.n2275 GNDA.n2256 3.4105
R15028 GNDA.n2288 GNDA.n2256 3.4105
R15029 GNDA.n2274 GNDA.n2256 3.4105
R15030 GNDA.n2290 GNDA.n2256 3.4105
R15031 GNDA.n2273 GNDA.n2256 3.4105
R15032 GNDA.n2292 GNDA.n2256 3.4105
R15033 GNDA.n2272 GNDA.n2256 3.4105
R15034 GNDA.n2294 GNDA.n2256 3.4105
R15035 GNDA.n2271 GNDA.n2256 3.4105
R15036 GNDA.n2296 GNDA.n2256 3.4105
R15037 GNDA.n2270 GNDA.n2256 3.4105
R15038 GNDA.n2298 GNDA.n2256 3.4105
R15039 GNDA.n2269 GNDA.n2256 3.4105
R15040 GNDA.n2300 GNDA.n2256 3.4105
R15041 GNDA.n2268 GNDA.n2256 3.4105
R15042 GNDA.n2302 GNDA.n2256 3.4105
R15043 GNDA.n2267 GNDA.n2256 3.4105
R15044 GNDA.n2304 GNDA.n2256 3.4105
R15045 GNDA.n2266 GNDA.n2256 3.4105
R15046 GNDA.n2305 GNDA.n2256 3.4105
R15047 GNDA.n2352 GNDA.n2256 3.4105
R15048 GNDA.n2354 GNDA.n2256 3.4105
R15049 GNDA.n2356 GNDA.n1959 3.4105
R15050 GNDA.n2280 GNDA.n1959 3.4105
R15051 GNDA.n2278 GNDA.n1959 3.4105
R15052 GNDA.n2282 GNDA.n1959 3.4105
R15053 GNDA.n2277 GNDA.n1959 3.4105
R15054 GNDA.n2284 GNDA.n1959 3.4105
R15055 GNDA.n2276 GNDA.n1959 3.4105
R15056 GNDA.n2286 GNDA.n1959 3.4105
R15057 GNDA.n2275 GNDA.n1959 3.4105
R15058 GNDA.n2288 GNDA.n1959 3.4105
R15059 GNDA.n2274 GNDA.n1959 3.4105
R15060 GNDA.n2290 GNDA.n1959 3.4105
R15061 GNDA.n2273 GNDA.n1959 3.4105
R15062 GNDA.n2292 GNDA.n1959 3.4105
R15063 GNDA.n2272 GNDA.n1959 3.4105
R15064 GNDA.n2294 GNDA.n1959 3.4105
R15065 GNDA.n2271 GNDA.n1959 3.4105
R15066 GNDA.n2296 GNDA.n1959 3.4105
R15067 GNDA.n2270 GNDA.n1959 3.4105
R15068 GNDA.n2298 GNDA.n1959 3.4105
R15069 GNDA.n2269 GNDA.n1959 3.4105
R15070 GNDA.n2300 GNDA.n1959 3.4105
R15071 GNDA.n2268 GNDA.n1959 3.4105
R15072 GNDA.n2302 GNDA.n1959 3.4105
R15073 GNDA.n2267 GNDA.n1959 3.4105
R15074 GNDA.n2304 GNDA.n1959 3.4105
R15075 GNDA.n2266 GNDA.n1959 3.4105
R15076 GNDA.n2305 GNDA.n1959 3.4105
R15077 GNDA.n2352 GNDA.n1959 3.4105
R15078 GNDA.n2354 GNDA.n1959 3.4105
R15079 GNDA.n2356 GNDA.n2257 3.4105
R15080 GNDA.n2280 GNDA.n2257 3.4105
R15081 GNDA.n2278 GNDA.n2257 3.4105
R15082 GNDA.n2282 GNDA.n2257 3.4105
R15083 GNDA.n2277 GNDA.n2257 3.4105
R15084 GNDA.n2284 GNDA.n2257 3.4105
R15085 GNDA.n2276 GNDA.n2257 3.4105
R15086 GNDA.n2286 GNDA.n2257 3.4105
R15087 GNDA.n2275 GNDA.n2257 3.4105
R15088 GNDA.n2288 GNDA.n2257 3.4105
R15089 GNDA.n2274 GNDA.n2257 3.4105
R15090 GNDA.n2290 GNDA.n2257 3.4105
R15091 GNDA.n2273 GNDA.n2257 3.4105
R15092 GNDA.n2292 GNDA.n2257 3.4105
R15093 GNDA.n2272 GNDA.n2257 3.4105
R15094 GNDA.n2294 GNDA.n2257 3.4105
R15095 GNDA.n2271 GNDA.n2257 3.4105
R15096 GNDA.n2296 GNDA.n2257 3.4105
R15097 GNDA.n2270 GNDA.n2257 3.4105
R15098 GNDA.n2298 GNDA.n2257 3.4105
R15099 GNDA.n2269 GNDA.n2257 3.4105
R15100 GNDA.n2300 GNDA.n2257 3.4105
R15101 GNDA.n2268 GNDA.n2257 3.4105
R15102 GNDA.n2302 GNDA.n2257 3.4105
R15103 GNDA.n2267 GNDA.n2257 3.4105
R15104 GNDA.n2304 GNDA.n2257 3.4105
R15105 GNDA.n2266 GNDA.n2257 3.4105
R15106 GNDA.n2305 GNDA.n2257 3.4105
R15107 GNDA.n2352 GNDA.n2257 3.4105
R15108 GNDA.n2354 GNDA.n2257 3.4105
R15109 GNDA.n2356 GNDA.n1958 3.4105
R15110 GNDA.n2280 GNDA.n1958 3.4105
R15111 GNDA.n2278 GNDA.n1958 3.4105
R15112 GNDA.n2282 GNDA.n1958 3.4105
R15113 GNDA.n2277 GNDA.n1958 3.4105
R15114 GNDA.n2284 GNDA.n1958 3.4105
R15115 GNDA.n2276 GNDA.n1958 3.4105
R15116 GNDA.n2286 GNDA.n1958 3.4105
R15117 GNDA.n2275 GNDA.n1958 3.4105
R15118 GNDA.n2288 GNDA.n1958 3.4105
R15119 GNDA.n2274 GNDA.n1958 3.4105
R15120 GNDA.n2290 GNDA.n1958 3.4105
R15121 GNDA.n2273 GNDA.n1958 3.4105
R15122 GNDA.n2292 GNDA.n1958 3.4105
R15123 GNDA.n2272 GNDA.n1958 3.4105
R15124 GNDA.n2294 GNDA.n1958 3.4105
R15125 GNDA.n2271 GNDA.n1958 3.4105
R15126 GNDA.n2296 GNDA.n1958 3.4105
R15127 GNDA.n2270 GNDA.n1958 3.4105
R15128 GNDA.n2298 GNDA.n1958 3.4105
R15129 GNDA.n2269 GNDA.n1958 3.4105
R15130 GNDA.n2300 GNDA.n1958 3.4105
R15131 GNDA.n2268 GNDA.n1958 3.4105
R15132 GNDA.n2302 GNDA.n1958 3.4105
R15133 GNDA.n2267 GNDA.n1958 3.4105
R15134 GNDA.n2304 GNDA.n1958 3.4105
R15135 GNDA.n2266 GNDA.n1958 3.4105
R15136 GNDA.n2305 GNDA.n1958 3.4105
R15137 GNDA.n2352 GNDA.n1958 3.4105
R15138 GNDA.n2354 GNDA.n1958 3.4105
R15139 GNDA.n2356 GNDA.n2258 3.4105
R15140 GNDA.n2280 GNDA.n2258 3.4105
R15141 GNDA.n2278 GNDA.n2258 3.4105
R15142 GNDA.n2282 GNDA.n2258 3.4105
R15143 GNDA.n2277 GNDA.n2258 3.4105
R15144 GNDA.n2284 GNDA.n2258 3.4105
R15145 GNDA.n2276 GNDA.n2258 3.4105
R15146 GNDA.n2286 GNDA.n2258 3.4105
R15147 GNDA.n2275 GNDA.n2258 3.4105
R15148 GNDA.n2288 GNDA.n2258 3.4105
R15149 GNDA.n2274 GNDA.n2258 3.4105
R15150 GNDA.n2290 GNDA.n2258 3.4105
R15151 GNDA.n2273 GNDA.n2258 3.4105
R15152 GNDA.n2292 GNDA.n2258 3.4105
R15153 GNDA.n2272 GNDA.n2258 3.4105
R15154 GNDA.n2294 GNDA.n2258 3.4105
R15155 GNDA.n2271 GNDA.n2258 3.4105
R15156 GNDA.n2296 GNDA.n2258 3.4105
R15157 GNDA.n2270 GNDA.n2258 3.4105
R15158 GNDA.n2298 GNDA.n2258 3.4105
R15159 GNDA.n2269 GNDA.n2258 3.4105
R15160 GNDA.n2300 GNDA.n2258 3.4105
R15161 GNDA.n2268 GNDA.n2258 3.4105
R15162 GNDA.n2302 GNDA.n2258 3.4105
R15163 GNDA.n2267 GNDA.n2258 3.4105
R15164 GNDA.n2304 GNDA.n2258 3.4105
R15165 GNDA.n2266 GNDA.n2258 3.4105
R15166 GNDA.n2305 GNDA.n2258 3.4105
R15167 GNDA.n2352 GNDA.n2258 3.4105
R15168 GNDA.n2354 GNDA.n2258 3.4105
R15169 GNDA.n2356 GNDA.n1957 3.4105
R15170 GNDA.n2280 GNDA.n1957 3.4105
R15171 GNDA.n2278 GNDA.n1957 3.4105
R15172 GNDA.n2282 GNDA.n1957 3.4105
R15173 GNDA.n2277 GNDA.n1957 3.4105
R15174 GNDA.n2284 GNDA.n1957 3.4105
R15175 GNDA.n2276 GNDA.n1957 3.4105
R15176 GNDA.n2286 GNDA.n1957 3.4105
R15177 GNDA.n2275 GNDA.n1957 3.4105
R15178 GNDA.n2288 GNDA.n1957 3.4105
R15179 GNDA.n2274 GNDA.n1957 3.4105
R15180 GNDA.n2290 GNDA.n1957 3.4105
R15181 GNDA.n2273 GNDA.n1957 3.4105
R15182 GNDA.n2292 GNDA.n1957 3.4105
R15183 GNDA.n2272 GNDA.n1957 3.4105
R15184 GNDA.n2294 GNDA.n1957 3.4105
R15185 GNDA.n2271 GNDA.n1957 3.4105
R15186 GNDA.n2296 GNDA.n1957 3.4105
R15187 GNDA.n2270 GNDA.n1957 3.4105
R15188 GNDA.n2298 GNDA.n1957 3.4105
R15189 GNDA.n2269 GNDA.n1957 3.4105
R15190 GNDA.n2300 GNDA.n1957 3.4105
R15191 GNDA.n2268 GNDA.n1957 3.4105
R15192 GNDA.n2302 GNDA.n1957 3.4105
R15193 GNDA.n2267 GNDA.n1957 3.4105
R15194 GNDA.n2304 GNDA.n1957 3.4105
R15195 GNDA.n2266 GNDA.n1957 3.4105
R15196 GNDA.n2305 GNDA.n1957 3.4105
R15197 GNDA.n2352 GNDA.n1957 3.4105
R15198 GNDA.n2354 GNDA.n1957 3.4105
R15199 GNDA.n2356 GNDA.n2259 3.4105
R15200 GNDA.n2280 GNDA.n2259 3.4105
R15201 GNDA.n2278 GNDA.n2259 3.4105
R15202 GNDA.n2282 GNDA.n2259 3.4105
R15203 GNDA.n2277 GNDA.n2259 3.4105
R15204 GNDA.n2284 GNDA.n2259 3.4105
R15205 GNDA.n2276 GNDA.n2259 3.4105
R15206 GNDA.n2286 GNDA.n2259 3.4105
R15207 GNDA.n2275 GNDA.n2259 3.4105
R15208 GNDA.n2288 GNDA.n2259 3.4105
R15209 GNDA.n2274 GNDA.n2259 3.4105
R15210 GNDA.n2290 GNDA.n2259 3.4105
R15211 GNDA.n2273 GNDA.n2259 3.4105
R15212 GNDA.n2292 GNDA.n2259 3.4105
R15213 GNDA.n2272 GNDA.n2259 3.4105
R15214 GNDA.n2294 GNDA.n2259 3.4105
R15215 GNDA.n2271 GNDA.n2259 3.4105
R15216 GNDA.n2296 GNDA.n2259 3.4105
R15217 GNDA.n2270 GNDA.n2259 3.4105
R15218 GNDA.n2298 GNDA.n2259 3.4105
R15219 GNDA.n2269 GNDA.n2259 3.4105
R15220 GNDA.n2300 GNDA.n2259 3.4105
R15221 GNDA.n2268 GNDA.n2259 3.4105
R15222 GNDA.n2302 GNDA.n2259 3.4105
R15223 GNDA.n2267 GNDA.n2259 3.4105
R15224 GNDA.n2304 GNDA.n2259 3.4105
R15225 GNDA.n2266 GNDA.n2259 3.4105
R15226 GNDA.n2305 GNDA.n2259 3.4105
R15227 GNDA.n2352 GNDA.n2259 3.4105
R15228 GNDA.n2354 GNDA.n2259 3.4105
R15229 GNDA.n2356 GNDA.n1956 3.4105
R15230 GNDA.n2280 GNDA.n1956 3.4105
R15231 GNDA.n2278 GNDA.n1956 3.4105
R15232 GNDA.n2282 GNDA.n1956 3.4105
R15233 GNDA.n2277 GNDA.n1956 3.4105
R15234 GNDA.n2284 GNDA.n1956 3.4105
R15235 GNDA.n2276 GNDA.n1956 3.4105
R15236 GNDA.n2286 GNDA.n1956 3.4105
R15237 GNDA.n2275 GNDA.n1956 3.4105
R15238 GNDA.n2288 GNDA.n1956 3.4105
R15239 GNDA.n2274 GNDA.n1956 3.4105
R15240 GNDA.n2290 GNDA.n1956 3.4105
R15241 GNDA.n2273 GNDA.n1956 3.4105
R15242 GNDA.n2292 GNDA.n1956 3.4105
R15243 GNDA.n2272 GNDA.n1956 3.4105
R15244 GNDA.n2294 GNDA.n1956 3.4105
R15245 GNDA.n2271 GNDA.n1956 3.4105
R15246 GNDA.n2296 GNDA.n1956 3.4105
R15247 GNDA.n2270 GNDA.n1956 3.4105
R15248 GNDA.n2298 GNDA.n1956 3.4105
R15249 GNDA.n2269 GNDA.n1956 3.4105
R15250 GNDA.n2300 GNDA.n1956 3.4105
R15251 GNDA.n2268 GNDA.n1956 3.4105
R15252 GNDA.n2302 GNDA.n1956 3.4105
R15253 GNDA.n2267 GNDA.n1956 3.4105
R15254 GNDA.n2304 GNDA.n1956 3.4105
R15255 GNDA.n2266 GNDA.n1956 3.4105
R15256 GNDA.n2305 GNDA.n1956 3.4105
R15257 GNDA.n2352 GNDA.n1956 3.4105
R15258 GNDA.n2354 GNDA.n1956 3.4105
R15259 GNDA.n2356 GNDA.n2260 3.4105
R15260 GNDA.n2280 GNDA.n2260 3.4105
R15261 GNDA.n2278 GNDA.n2260 3.4105
R15262 GNDA.n2282 GNDA.n2260 3.4105
R15263 GNDA.n2277 GNDA.n2260 3.4105
R15264 GNDA.n2284 GNDA.n2260 3.4105
R15265 GNDA.n2276 GNDA.n2260 3.4105
R15266 GNDA.n2286 GNDA.n2260 3.4105
R15267 GNDA.n2275 GNDA.n2260 3.4105
R15268 GNDA.n2288 GNDA.n2260 3.4105
R15269 GNDA.n2274 GNDA.n2260 3.4105
R15270 GNDA.n2290 GNDA.n2260 3.4105
R15271 GNDA.n2273 GNDA.n2260 3.4105
R15272 GNDA.n2292 GNDA.n2260 3.4105
R15273 GNDA.n2272 GNDA.n2260 3.4105
R15274 GNDA.n2294 GNDA.n2260 3.4105
R15275 GNDA.n2271 GNDA.n2260 3.4105
R15276 GNDA.n2296 GNDA.n2260 3.4105
R15277 GNDA.n2270 GNDA.n2260 3.4105
R15278 GNDA.n2298 GNDA.n2260 3.4105
R15279 GNDA.n2269 GNDA.n2260 3.4105
R15280 GNDA.n2300 GNDA.n2260 3.4105
R15281 GNDA.n2268 GNDA.n2260 3.4105
R15282 GNDA.n2302 GNDA.n2260 3.4105
R15283 GNDA.n2267 GNDA.n2260 3.4105
R15284 GNDA.n2304 GNDA.n2260 3.4105
R15285 GNDA.n2266 GNDA.n2260 3.4105
R15286 GNDA.n2305 GNDA.n2260 3.4105
R15287 GNDA.n2352 GNDA.n2260 3.4105
R15288 GNDA.n2354 GNDA.n2260 3.4105
R15289 GNDA.n2356 GNDA.n1955 3.4105
R15290 GNDA.n2280 GNDA.n1955 3.4105
R15291 GNDA.n2278 GNDA.n1955 3.4105
R15292 GNDA.n2282 GNDA.n1955 3.4105
R15293 GNDA.n2277 GNDA.n1955 3.4105
R15294 GNDA.n2284 GNDA.n1955 3.4105
R15295 GNDA.n2276 GNDA.n1955 3.4105
R15296 GNDA.n2286 GNDA.n1955 3.4105
R15297 GNDA.n2275 GNDA.n1955 3.4105
R15298 GNDA.n2288 GNDA.n1955 3.4105
R15299 GNDA.n2274 GNDA.n1955 3.4105
R15300 GNDA.n2290 GNDA.n1955 3.4105
R15301 GNDA.n2273 GNDA.n1955 3.4105
R15302 GNDA.n2292 GNDA.n1955 3.4105
R15303 GNDA.n2272 GNDA.n1955 3.4105
R15304 GNDA.n2294 GNDA.n1955 3.4105
R15305 GNDA.n2271 GNDA.n1955 3.4105
R15306 GNDA.n2296 GNDA.n1955 3.4105
R15307 GNDA.n2270 GNDA.n1955 3.4105
R15308 GNDA.n2298 GNDA.n1955 3.4105
R15309 GNDA.n2269 GNDA.n1955 3.4105
R15310 GNDA.n2300 GNDA.n1955 3.4105
R15311 GNDA.n2268 GNDA.n1955 3.4105
R15312 GNDA.n2302 GNDA.n1955 3.4105
R15313 GNDA.n2267 GNDA.n1955 3.4105
R15314 GNDA.n2304 GNDA.n1955 3.4105
R15315 GNDA.n2266 GNDA.n1955 3.4105
R15316 GNDA.n2305 GNDA.n1955 3.4105
R15317 GNDA.n2352 GNDA.n1955 3.4105
R15318 GNDA.n2354 GNDA.n1955 3.4105
R15319 GNDA.n2356 GNDA.n2261 3.4105
R15320 GNDA.n2280 GNDA.n2261 3.4105
R15321 GNDA.n2278 GNDA.n2261 3.4105
R15322 GNDA.n2282 GNDA.n2261 3.4105
R15323 GNDA.n2277 GNDA.n2261 3.4105
R15324 GNDA.n2284 GNDA.n2261 3.4105
R15325 GNDA.n2276 GNDA.n2261 3.4105
R15326 GNDA.n2286 GNDA.n2261 3.4105
R15327 GNDA.n2275 GNDA.n2261 3.4105
R15328 GNDA.n2288 GNDA.n2261 3.4105
R15329 GNDA.n2274 GNDA.n2261 3.4105
R15330 GNDA.n2290 GNDA.n2261 3.4105
R15331 GNDA.n2273 GNDA.n2261 3.4105
R15332 GNDA.n2292 GNDA.n2261 3.4105
R15333 GNDA.n2272 GNDA.n2261 3.4105
R15334 GNDA.n2294 GNDA.n2261 3.4105
R15335 GNDA.n2271 GNDA.n2261 3.4105
R15336 GNDA.n2296 GNDA.n2261 3.4105
R15337 GNDA.n2270 GNDA.n2261 3.4105
R15338 GNDA.n2298 GNDA.n2261 3.4105
R15339 GNDA.n2269 GNDA.n2261 3.4105
R15340 GNDA.n2300 GNDA.n2261 3.4105
R15341 GNDA.n2268 GNDA.n2261 3.4105
R15342 GNDA.n2302 GNDA.n2261 3.4105
R15343 GNDA.n2267 GNDA.n2261 3.4105
R15344 GNDA.n2304 GNDA.n2261 3.4105
R15345 GNDA.n2266 GNDA.n2261 3.4105
R15346 GNDA.n2305 GNDA.n2261 3.4105
R15347 GNDA.n2352 GNDA.n2261 3.4105
R15348 GNDA.n2354 GNDA.n2261 3.4105
R15349 GNDA.n2356 GNDA.n1954 3.4105
R15350 GNDA.n2280 GNDA.n1954 3.4105
R15351 GNDA.n2278 GNDA.n1954 3.4105
R15352 GNDA.n2282 GNDA.n1954 3.4105
R15353 GNDA.n2277 GNDA.n1954 3.4105
R15354 GNDA.n2284 GNDA.n1954 3.4105
R15355 GNDA.n2276 GNDA.n1954 3.4105
R15356 GNDA.n2286 GNDA.n1954 3.4105
R15357 GNDA.n2275 GNDA.n1954 3.4105
R15358 GNDA.n2288 GNDA.n1954 3.4105
R15359 GNDA.n2274 GNDA.n1954 3.4105
R15360 GNDA.n2290 GNDA.n1954 3.4105
R15361 GNDA.n2273 GNDA.n1954 3.4105
R15362 GNDA.n2292 GNDA.n1954 3.4105
R15363 GNDA.n2272 GNDA.n1954 3.4105
R15364 GNDA.n2294 GNDA.n1954 3.4105
R15365 GNDA.n2271 GNDA.n1954 3.4105
R15366 GNDA.n2296 GNDA.n1954 3.4105
R15367 GNDA.n2270 GNDA.n1954 3.4105
R15368 GNDA.n2298 GNDA.n1954 3.4105
R15369 GNDA.n2269 GNDA.n1954 3.4105
R15370 GNDA.n2300 GNDA.n1954 3.4105
R15371 GNDA.n2268 GNDA.n1954 3.4105
R15372 GNDA.n2302 GNDA.n1954 3.4105
R15373 GNDA.n2267 GNDA.n1954 3.4105
R15374 GNDA.n2304 GNDA.n1954 3.4105
R15375 GNDA.n2266 GNDA.n1954 3.4105
R15376 GNDA.n2305 GNDA.n1954 3.4105
R15377 GNDA.n2352 GNDA.n1954 3.4105
R15378 GNDA.n2354 GNDA.n1954 3.4105
R15379 GNDA.n2356 GNDA.n2262 3.4105
R15380 GNDA.n2280 GNDA.n2262 3.4105
R15381 GNDA.n2278 GNDA.n2262 3.4105
R15382 GNDA.n2282 GNDA.n2262 3.4105
R15383 GNDA.n2277 GNDA.n2262 3.4105
R15384 GNDA.n2284 GNDA.n2262 3.4105
R15385 GNDA.n2276 GNDA.n2262 3.4105
R15386 GNDA.n2286 GNDA.n2262 3.4105
R15387 GNDA.n2275 GNDA.n2262 3.4105
R15388 GNDA.n2288 GNDA.n2262 3.4105
R15389 GNDA.n2274 GNDA.n2262 3.4105
R15390 GNDA.n2290 GNDA.n2262 3.4105
R15391 GNDA.n2273 GNDA.n2262 3.4105
R15392 GNDA.n2292 GNDA.n2262 3.4105
R15393 GNDA.n2272 GNDA.n2262 3.4105
R15394 GNDA.n2294 GNDA.n2262 3.4105
R15395 GNDA.n2271 GNDA.n2262 3.4105
R15396 GNDA.n2296 GNDA.n2262 3.4105
R15397 GNDA.n2270 GNDA.n2262 3.4105
R15398 GNDA.n2298 GNDA.n2262 3.4105
R15399 GNDA.n2269 GNDA.n2262 3.4105
R15400 GNDA.n2300 GNDA.n2262 3.4105
R15401 GNDA.n2268 GNDA.n2262 3.4105
R15402 GNDA.n2302 GNDA.n2262 3.4105
R15403 GNDA.n2267 GNDA.n2262 3.4105
R15404 GNDA.n2304 GNDA.n2262 3.4105
R15405 GNDA.n2266 GNDA.n2262 3.4105
R15406 GNDA.n2305 GNDA.n2262 3.4105
R15407 GNDA.n2352 GNDA.n2262 3.4105
R15408 GNDA.n2354 GNDA.n2262 3.4105
R15409 GNDA.n2356 GNDA.n1953 3.4105
R15410 GNDA.n2280 GNDA.n1953 3.4105
R15411 GNDA.n2278 GNDA.n1953 3.4105
R15412 GNDA.n2282 GNDA.n1953 3.4105
R15413 GNDA.n2277 GNDA.n1953 3.4105
R15414 GNDA.n2284 GNDA.n1953 3.4105
R15415 GNDA.n2276 GNDA.n1953 3.4105
R15416 GNDA.n2286 GNDA.n1953 3.4105
R15417 GNDA.n2275 GNDA.n1953 3.4105
R15418 GNDA.n2288 GNDA.n1953 3.4105
R15419 GNDA.n2274 GNDA.n1953 3.4105
R15420 GNDA.n2290 GNDA.n1953 3.4105
R15421 GNDA.n2273 GNDA.n1953 3.4105
R15422 GNDA.n2292 GNDA.n1953 3.4105
R15423 GNDA.n2272 GNDA.n1953 3.4105
R15424 GNDA.n2294 GNDA.n1953 3.4105
R15425 GNDA.n2271 GNDA.n1953 3.4105
R15426 GNDA.n2296 GNDA.n1953 3.4105
R15427 GNDA.n2270 GNDA.n1953 3.4105
R15428 GNDA.n2298 GNDA.n1953 3.4105
R15429 GNDA.n2269 GNDA.n1953 3.4105
R15430 GNDA.n2300 GNDA.n1953 3.4105
R15431 GNDA.n2268 GNDA.n1953 3.4105
R15432 GNDA.n2302 GNDA.n1953 3.4105
R15433 GNDA.n2267 GNDA.n1953 3.4105
R15434 GNDA.n2304 GNDA.n1953 3.4105
R15435 GNDA.n2266 GNDA.n1953 3.4105
R15436 GNDA.n2305 GNDA.n1953 3.4105
R15437 GNDA.n2352 GNDA.n1953 3.4105
R15438 GNDA.n2354 GNDA.n1953 3.4105
R15439 GNDA.n2356 GNDA.n2263 3.4105
R15440 GNDA.n2280 GNDA.n2263 3.4105
R15441 GNDA.n2278 GNDA.n2263 3.4105
R15442 GNDA.n2282 GNDA.n2263 3.4105
R15443 GNDA.n2277 GNDA.n2263 3.4105
R15444 GNDA.n2284 GNDA.n2263 3.4105
R15445 GNDA.n2276 GNDA.n2263 3.4105
R15446 GNDA.n2286 GNDA.n2263 3.4105
R15447 GNDA.n2275 GNDA.n2263 3.4105
R15448 GNDA.n2288 GNDA.n2263 3.4105
R15449 GNDA.n2274 GNDA.n2263 3.4105
R15450 GNDA.n2290 GNDA.n2263 3.4105
R15451 GNDA.n2273 GNDA.n2263 3.4105
R15452 GNDA.n2292 GNDA.n2263 3.4105
R15453 GNDA.n2272 GNDA.n2263 3.4105
R15454 GNDA.n2294 GNDA.n2263 3.4105
R15455 GNDA.n2271 GNDA.n2263 3.4105
R15456 GNDA.n2296 GNDA.n2263 3.4105
R15457 GNDA.n2270 GNDA.n2263 3.4105
R15458 GNDA.n2298 GNDA.n2263 3.4105
R15459 GNDA.n2269 GNDA.n2263 3.4105
R15460 GNDA.n2300 GNDA.n2263 3.4105
R15461 GNDA.n2268 GNDA.n2263 3.4105
R15462 GNDA.n2302 GNDA.n2263 3.4105
R15463 GNDA.n2267 GNDA.n2263 3.4105
R15464 GNDA.n2304 GNDA.n2263 3.4105
R15465 GNDA.n2266 GNDA.n2263 3.4105
R15466 GNDA.n2305 GNDA.n2263 3.4105
R15467 GNDA.n2352 GNDA.n2263 3.4105
R15468 GNDA.n2354 GNDA.n2263 3.4105
R15469 GNDA.n2356 GNDA.n1952 3.4105
R15470 GNDA.n2280 GNDA.n1952 3.4105
R15471 GNDA.n2278 GNDA.n1952 3.4105
R15472 GNDA.n2282 GNDA.n1952 3.4105
R15473 GNDA.n2277 GNDA.n1952 3.4105
R15474 GNDA.n2284 GNDA.n1952 3.4105
R15475 GNDA.n2276 GNDA.n1952 3.4105
R15476 GNDA.n2286 GNDA.n1952 3.4105
R15477 GNDA.n2275 GNDA.n1952 3.4105
R15478 GNDA.n2288 GNDA.n1952 3.4105
R15479 GNDA.n2274 GNDA.n1952 3.4105
R15480 GNDA.n2290 GNDA.n1952 3.4105
R15481 GNDA.n2273 GNDA.n1952 3.4105
R15482 GNDA.n2292 GNDA.n1952 3.4105
R15483 GNDA.n2272 GNDA.n1952 3.4105
R15484 GNDA.n2294 GNDA.n1952 3.4105
R15485 GNDA.n2271 GNDA.n1952 3.4105
R15486 GNDA.n2296 GNDA.n1952 3.4105
R15487 GNDA.n2270 GNDA.n1952 3.4105
R15488 GNDA.n2298 GNDA.n1952 3.4105
R15489 GNDA.n2269 GNDA.n1952 3.4105
R15490 GNDA.n2300 GNDA.n1952 3.4105
R15491 GNDA.n2268 GNDA.n1952 3.4105
R15492 GNDA.n2302 GNDA.n1952 3.4105
R15493 GNDA.n2267 GNDA.n1952 3.4105
R15494 GNDA.n2304 GNDA.n1952 3.4105
R15495 GNDA.n2266 GNDA.n1952 3.4105
R15496 GNDA.n2305 GNDA.n1952 3.4105
R15497 GNDA.n2352 GNDA.n1952 3.4105
R15498 GNDA.n2354 GNDA.n1952 3.4105
R15499 GNDA.n2356 GNDA.n2355 3.4105
R15500 GNDA.n2355 GNDA.n2280 3.4105
R15501 GNDA.n2355 GNDA.n2278 3.4105
R15502 GNDA.n2355 GNDA.n2282 3.4105
R15503 GNDA.n2355 GNDA.n2277 3.4105
R15504 GNDA.n2355 GNDA.n2284 3.4105
R15505 GNDA.n2355 GNDA.n2276 3.4105
R15506 GNDA.n2355 GNDA.n2286 3.4105
R15507 GNDA.n2355 GNDA.n2275 3.4105
R15508 GNDA.n2355 GNDA.n2288 3.4105
R15509 GNDA.n2355 GNDA.n2274 3.4105
R15510 GNDA.n2355 GNDA.n2290 3.4105
R15511 GNDA.n2355 GNDA.n2273 3.4105
R15512 GNDA.n2355 GNDA.n2292 3.4105
R15513 GNDA.n2355 GNDA.n2272 3.4105
R15514 GNDA.n2355 GNDA.n2294 3.4105
R15515 GNDA.n2355 GNDA.n2271 3.4105
R15516 GNDA.n2355 GNDA.n2296 3.4105
R15517 GNDA.n2355 GNDA.n2270 3.4105
R15518 GNDA.n2355 GNDA.n2298 3.4105
R15519 GNDA.n2355 GNDA.n2269 3.4105
R15520 GNDA.n2355 GNDA.n2300 3.4105
R15521 GNDA.n2355 GNDA.n2268 3.4105
R15522 GNDA.n2355 GNDA.n2302 3.4105
R15523 GNDA.n2355 GNDA.n2267 3.4105
R15524 GNDA.n2355 GNDA.n2304 3.4105
R15525 GNDA.n2355 GNDA.n2266 3.4105
R15526 GNDA.n2355 GNDA.n2305 3.4105
R15527 GNDA.n2355 GNDA.n2354 3.4105
R15528 GNDA.n2243 GNDA.n1981 3.4105
R15529 GNDA.n2026 GNDA.n1981 3.4105
R15530 GNDA.n2026 GNDA.n1980 3.4105
R15531 GNDA.n2245 GNDA.n2026 3.4105
R15532 GNDA.n2247 GNDA.n2026 3.4105
R15533 GNDA.n2012 GNDA.n1981 3.4105
R15534 GNDA.n2012 GNDA.n1983 3.4105
R15535 GNDA.n2012 GNDA.n1979 3.4105
R15536 GNDA.n2012 GNDA.n1984 3.4105
R15537 GNDA.n2012 GNDA.n1978 3.4105
R15538 GNDA.n2012 GNDA.n1985 3.4105
R15539 GNDA.n2012 GNDA.n1977 3.4105
R15540 GNDA.n2012 GNDA.n1986 3.4105
R15541 GNDA.n2012 GNDA.n1976 3.4105
R15542 GNDA.n2012 GNDA.n1987 3.4105
R15543 GNDA.n2012 GNDA.n1975 3.4105
R15544 GNDA.n2012 GNDA.n1988 3.4105
R15545 GNDA.n2012 GNDA.n1974 3.4105
R15546 GNDA.n2012 GNDA.n1989 3.4105
R15547 GNDA.n2012 GNDA.n1973 3.4105
R15548 GNDA.n2012 GNDA.n1990 3.4105
R15549 GNDA.n2012 GNDA.n1972 3.4105
R15550 GNDA.n2012 GNDA.n1991 3.4105
R15551 GNDA.n2012 GNDA.n1971 3.4105
R15552 GNDA.n2012 GNDA.n1992 3.4105
R15553 GNDA.n2012 GNDA.n1970 3.4105
R15554 GNDA.n2012 GNDA.n1993 3.4105
R15555 GNDA.n2012 GNDA.n1969 3.4105
R15556 GNDA.n2012 GNDA.n1994 3.4105
R15557 GNDA.n2012 GNDA.n1968 3.4105
R15558 GNDA.n2012 GNDA.n1995 3.4105
R15559 GNDA.n2245 GNDA.n2012 3.4105
R15560 GNDA.n2247 GNDA.n2012 3.4105
R15561 GNDA.n2028 GNDA.n1980 3.4105
R15562 GNDA.n2028 GNDA.n1983 3.4105
R15563 GNDA.n2028 GNDA.n1979 3.4105
R15564 GNDA.n2028 GNDA.n1984 3.4105
R15565 GNDA.n2028 GNDA.n1978 3.4105
R15566 GNDA.n2028 GNDA.n1985 3.4105
R15567 GNDA.n2028 GNDA.n1977 3.4105
R15568 GNDA.n2028 GNDA.n1986 3.4105
R15569 GNDA.n2028 GNDA.n1976 3.4105
R15570 GNDA.n2028 GNDA.n1987 3.4105
R15571 GNDA.n2028 GNDA.n1975 3.4105
R15572 GNDA.n2028 GNDA.n1988 3.4105
R15573 GNDA.n2028 GNDA.n1974 3.4105
R15574 GNDA.n2028 GNDA.n1989 3.4105
R15575 GNDA.n2028 GNDA.n1973 3.4105
R15576 GNDA.n2028 GNDA.n1990 3.4105
R15577 GNDA.n2028 GNDA.n1972 3.4105
R15578 GNDA.n2028 GNDA.n1991 3.4105
R15579 GNDA.n2028 GNDA.n1971 3.4105
R15580 GNDA.n2028 GNDA.n1992 3.4105
R15581 GNDA.n2028 GNDA.n1970 3.4105
R15582 GNDA.n2028 GNDA.n1993 3.4105
R15583 GNDA.n2028 GNDA.n1969 3.4105
R15584 GNDA.n2028 GNDA.n1994 3.4105
R15585 GNDA.n2028 GNDA.n1968 3.4105
R15586 GNDA.n2028 GNDA.n1995 3.4105
R15587 GNDA.n2245 GNDA.n2028 3.4105
R15588 GNDA.n2247 GNDA.n2028 3.4105
R15589 GNDA.n2010 GNDA.n1981 3.4105
R15590 GNDA.n2010 GNDA.n1982 3.4105
R15591 GNDA.n2010 GNDA.n1980 3.4105
R15592 GNDA.n2010 GNDA.n1983 3.4105
R15593 GNDA.n2010 GNDA.n1979 3.4105
R15594 GNDA.n2010 GNDA.n1984 3.4105
R15595 GNDA.n2010 GNDA.n1978 3.4105
R15596 GNDA.n2010 GNDA.n1985 3.4105
R15597 GNDA.n2010 GNDA.n1977 3.4105
R15598 GNDA.n2010 GNDA.n1986 3.4105
R15599 GNDA.n2010 GNDA.n1976 3.4105
R15600 GNDA.n2010 GNDA.n1987 3.4105
R15601 GNDA.n2010 GNDA.n1975 3.4105
R15602 GNDA.n2010 GNDA.n1988 3.4105
R15603 GNDA.n2010 GNDA.n1974 3.4105
R15604 GNDA.n2010 GNDA.n1989 3.4105
R15605 GNDA.n2010 GNDA.n1973 3.4105
R15606 GNDA.n2010 GNDA.n1990 3.4105
R15607 GNDA.n2010 GNDA.n1972 3.4105
R15608 GNDA.n2010 GNDA.n1991 3.4105
R15609 GNDA.n2010 GNDA.n1971 3.4105
R15610 GNDA.n2010 GNDA.n1992 3.4105
R15611 GNDA.n2010 GNDA.n1970 3.4105
R15612 GNDA.n2010 GNDA.n1993 3.4105
R15613 GNDA.n2010 GNDA.n1969 3.4105
R15614 GNDA.n2010 GNDA.n1994 3.4105
R15615 GNDA.n2010 GNDA.n1968 3.4105
R15616 GNDA.n2010 GNDA.n1995 3.4105
R15617 GNDA.n2245 GNDA.n2010 3.4105
R15618 GNDA.n2247 GNDA.n2010 3.4105
R15619 GNDA.n2029 GNDA.n1981 3.4105
R15620 GNDA.n2029 GNDA.n1982 3.4105
R15621 GNDA.n2029 GNDA.n1980 3.4105
R15622 GNDA.n2029 GNDA.n1983 3.4105
R15623 GNDA.n2029 GNDA.n1979 3.4105
R15624 GNDA.n2029 GNDA.n1984 3.4105
R15625 GNDA.n2029 GNDA.n1978 3.4105
R15626 GNDA.n2029 GNDA.n1985 3.4105
R15627 GNDA.n2029 GNDA.n1977 3.4105
R15628 GNDA.n2029 GNDA.n1986 3.4105
R15629 GNDA.n2029 GNDA.n1976 3.4105
R15630 GNDA.n2029 GNDA.n1987 3.4105
R15631 GNDA.n2029 GNDA.n1975 3.4105
R15632 GNDA.n2029 GNDA.n1988 3.4105
R15633 GNDA.n2029 GNDA.n1974 3.4105
R15634 GNDA.n2029 GNDA.n1989 3.4105
R15635 GNDA.n2029 GNDA.n1973 3.4105
R15636 GNDA.n2029 GNDA.n1990 3.4105
R15637 GNDA.n2029 GNDA.n1972 3.4105
R15638 GNDA.n2029 GNDA.n1991 3.4105
R15639 GNDA.n2029 GNDA.n1971 3.4105
R15640 GNDA.n2029 GNDA.n1992 3.4105
R15641 GNDA.n2029 GNDA.n1970 3.4105
R15642 GNDA.n2029 GNDA.n1993 3.4105
R15643 GNDA.n2029 GNDA.n1969 3.4105
R15644 GNDA.n2029 GNDA.n1994 3.4105
R15645 GNDA.n2029 GNDA.n1968 3.4105
R15646 GNDA.n2029 GNDA.n1995 3.4105
R15647 GNDA.n2245 GNDA.n2029 3.4105
R15648 GNDA.n2247 GNDA.n2029 3.4105
R15649 GNDA.n2009 GNDA.n1981 3.4105
R15650 GNDA.n2009 GNDA.n1982 3.4105
R15651 GNDA.n2009 GNDA.n1980 3.4105
R15652 GNDA.n2009 GNDA.n1983 3.4105
R15653 GNDA.n2009 GNDA.n1979 3.4105
R15654 GNDA.n2009 GNDA.n1984 3.4105
R15655 GNDA.n2009 GNDA.n1978 3.4105
R15656 GNDA.n2009 GNDA.n1985 3.4105
R15657 GNDA.n2009 GNDA.n1977 3.4105
R15658 GNDA.n2009 GNDA.n1986 3.4105
R15659 GNDA.n2009 GNDA.n1976 3.4105
R15660 GNDA.n2009 GNDA.n1987 3.4105
R15661 GNDA.n2009 GNDA.n1975 3.4105
R15662 GNDA.n2009 GNDA.n1988 3.4105
R15663 GNDA.n2009 GNDA.n1974 3.4105
R15664 GNDA.n2009 GNDA.n1989 3.4105
R15665 GNDA.n2009 GNDA.n1973 3.4105
R15666 GNDA.n2009 GNDA.n1990 3.4105
R15667 GNDA.n2009 GNDA.n1972 3.4105
R15668 GNDA.n2009 GNDA.n1991 3.4105
R15669 GNDA.n2009 GNDA.n1971 3.4105
R15670 GNDA.n2009 GNDA.n1992 3.4105
R15671 GNDA.n2009 GNDA.n1970 3.4105
R15672 GNDA.n2009 GNDA.n1993 3.4105
R15673 GNDA.n2009 GNDA.n1969 3.4105
R15674 GNDA.n2009 GNDA.n1994 3.4105
R15675 GNDA.n2009 GNDA.n1968 3.4105
R15676 GNDA.n2009 GNDA.n1995 3.4105
R15677 GNDA.n2245 GNDA.n2009 3.4105
R15678 GNDA.n2247 GNDA.n2009 3.4105
R15679 GNDA.n2030 GNDA.n1981 3.4105
R15680 GNDA.n2030 GNDA.n1982 3.4105
R15681 GNDA.n2030 GNDA.n1980 3.4105
R15682 GNDA.n2030 GNDA.n1983 3.4105
R15683 GNDA.n2030 GNDA.n1979 3.4105
R15684 GNDA.n2030 GNDA.n1984 3.4105
R15685 GNDA.n2030 GNDA.n1978 3.4105
R15686 GNDA.n2030 GNDA.n1985 3.4105
R15687 GNDA.n2030 GNDA.n1977 3.4105
R15688 GNDA.n2030 GNDA.n1986 3.4105
R15689 GNDA.n2030 GNDA.n1976 3.4105
R15690 GNDA.n2030 GNDA.n1987 3.4105
R15691 GNDA.n2030 GNDA.n1975 3.4105
R15692 GNDA.n2030 GNDA.n1988 3.4105
R15693 GNDA.n2030 GNDA.n1974 3.4105
R15694 GNDA.n2030 GNDA.n1989 3.4105
R15695 GNDA.n2030 GNDA.n1973 3.4105
R15696 GNDA.n2030 GNDA.n1990 3.4105
R15697 GNDA.n2030 GNDA.n1972 3.4105
R15698 GNDA.n2030 GNDA.n1991 3.4105
R15699 GNDA.n2030 GNDA.n1971 3.4105
R15700 GNDA.n2030 GNDA.n1992 3.4105
R15701 GNDA.n2030 GNDA.n1970 3.4105
R15702 GNDA.n2030 GNDA.n1993 3.4105
R15703 GNDA.n2030 GNDA.n1969 3.4105
R15704 GNDA.n2030 GNDA.n1994 3.4105
R15705 GNDA.n2030 GNDA.n1968 3.4105
R15706 GNDA.n2030 GNDA.n1995 3.4105
R15707 GNDA.n2245 GNDA.n2030 3.4105
R15708 GNDA.n2247 GNDA.n2030 3.4105
R15709 GNDA.n2008 GNDA.n1981 3.4105
R15710 GNDA.n2008 GNDA.n1982 3.4105
R15711 GNDA.n2008 GNDA.n1980 3.4105
R15712 GNDA.n2008 GNDA.n1983 3.4105
R15713 GNDA.n2008 GNDA.n1979 3.4105
R15714 GNDA.n2008 GNDA.n1984 3.4105
R15715 GNDA.n2008 GNDA.n1978 3.4105
R15716 GNDA.n2008 GNDA.n1985 3.4105
R15717 GNDA.n2008 GNDA.n1977 3.4105
R15718 GNDA.n2008 GNDA.n1986 3.4105
R15719 GNDA.n2008 GNDA.n1976 3.4105
R15720 GNDA.n2008 GNDA.n1987 3.4105
R15721 GNDA.n2008 GNDA.n1975 3.4105
R15722 GNDA.n2008 GNDA.n1988 3.4105
R15723 GNDA.n2008 GNDA.n1974 3.4105
R15724 GNDA.n2008 GNDA.n1989 3.4105
R15725 GNDA.n2008 GNDA.n1973 3.4105
R15726 GNDA.n2008 GNDA.n1990 3.4105
R15727 GNDA.n2008 GNDA.n1972 3.4105
R15728 GNDA.n2008 GNDA.n1991 3.4105
R15729 GNDA.n2008 GNDA.n1971 3.4105
R15730 GNDA.n2008 GNDA.n1992 3.4105
R15731 GNDA.n2008 GNDA.n1970 3.4105
R15732 GNDA.n2008 GNDA.n1993 3.4105
R15733 GNDA.n2008 GNDA.n1969 3.4105
R15734 GNDA.n2008 GNDA.n1994 3.4105
R15735 GNDA.n2008 GNDA.n1968 3.4105
R15736 GNDA.n2008 GNDA.n1995 3.4105
R15737 GNDA.n2245 GNDA.n2008 3.4105
R15738 GNDA.n2247 GNDA.n2008 3.4105
R15739 GNDA.n2031 GNDA.n1981 3.4105
R15740 GNDA.n2031 GNDA.n1982 3.4105
R15741 GNDA.n2031 GNDA.n1980 3.4105
R15742 GNDA.n2031 GNDA.n1983 3.4105
R15743 GNDA.n2031 GNDA.n1979 3.4105
R15744 GNDA.n2031 GNDA.n1984 3.4105
R15745 GNDA.n2031 GNDA.n1978 3.4105
R15746 GNDA.n2031 GNDA.n1985 3.4105
R15747 GNDA.n2031 GNDA.n1977 3.4105
R15748 GNDA.n2031 GNDA.n1986 3.4105
R15749 GNDA.n2031 GNDA.n1976 3.4105
R15750 GNDA.n2031 GNDA.n1987 3.4105
R15751 GNDA.n2031 GNDA.n1975 3.4105
R15752 GNDA.n2031 GNDA.n1988 3.4105
R15753 GNDA.n2031 GNDA.n1974 3.4105
R15754 GNDA.n2031 GNDA.n1989 3.4105
R15755 GNDA.n2031 GNDA.n1973 3.4105
R15756 GNDA.n2031 GNDA.n1990 3.4105
R15757 GNDA.n2031 GNDA.n1972 3.4105
R15758 GNDA.n2031 GNDA.n1991 3.4105
R15759 GNDA.n2031 GNDA.n1971 3.4105
R15760 GNDA.n2031 GNDA.n1992 3.4105
R15761 GNDA.n2031 GNDA.n1970 3.4105
R15762 GNDA.n2031 GNDA.n1993 3.4105
R15763 GNDA.n2031 GNDA.n1969 3.4105
R15764 GNDA.n2031 GNDA.n1994 3.4105
R15765 GNDA.n2031 GNDA.n1968 3.4105
R15766 GNDA.n2031 GNDA.n1995 3.4105
R15767 GNDA.n2245 GNDA.n2031 3.4105
R15768 GNDA.n2247 GNDA.n2031 3.4105
R15769 GNDA.n2007 GNDA.n1981 3.4105
R15770 GNDA.n2007 GNDA.n1982 3.4105
R15771 GNDA.n2007 GNDA.n1980 3.4105
R15772 GNDA.n2007 GNDA.n1983 3.4105
R15773 GNDA.n2007 GNDA.n1979 3.4105
R15774 GNDA.n2007 GNDA.n1984 3.4105
R15775 GNDA.n2007 GNDA.n1978 3.4105
R15776 GNDA.n2007 GNDA.n1985 3.4105
R15777 GNDA.n2007 GNDA.n1977 3.4105
R15778 GNDA.n2007 GNDA.n1986 3.4105
R15779 GNDA.n2007 GNDA.n1976 3.4105
R15780 GNDA.n2007 GNDA.n1987 3.4105
R15781 GNDA.n2007 GNDA.n1975 3.4105
R15782 GNDA.n2007 GNDA.n1988 3.4105
R15783 GNDA.n2007 GNDA.n1974 3.4105
R15784 GNDA.n2007 GNDA.n1989 3.4105
R15785 GNDA.n2007 GNDA.n1973 3.4105
R15786 GNDA.n2007 GNDA.n1990 3.4105
R15787 GNDA.n2007 GNDA.n1972 3.4105
R15788 GNDA.n2007 GNDA.n1991 3.4105
R15789 GNDA.n2007 GNDA.n1971 3.4105
R15790 GNDA.n2007 GNDA.n1992 3.4105
R15791 GNDA.n2007 GNDA.n1970 3.4105
R15792 GNDA.n2007 GNDA.n1993 3.4105
R15793 GNDA.n2007 GNDA.n1969 3.4105
R15794 GNDA.n2007 GNDA.n1994 3.4105
R15795 GNDA.n2007 GNDA.n1968 3.4105
R15796 GNDA.n2007 GNDA.n1995 3.4105
R15797 GNDA.n2245 GNDA.n2007 3.4105
R15798 GNDA.n2247 GNDA.n2007 3.4105
R15799 GNDA.n2032 GNDA.n1981 3.4105
R15800 GNDA.n2032 GNDA.n1982 3.4105
R15801 GNDA.n2032 GNDA.n1980 3.4105
R15802 GNDA.n2032 GNDA.n1983 3.4105
R15803 GNDA.n2032 GNDA.n1979 3.4105
R15804 GNDA.n2032 GNDA.n1984 3.4105
R15805 GNDA.n2032 GNDA.n1978 3.4105
R15806 GNDA.n2032 GNDA.n1985 3.4105
R15807 GNDA.n2032 GNDA.n1977 3.4105
R15808 GNDA.n2032 GNDA.n1986 3.4105
R15809 GNDA.n2032 GNDA.n1976 3.4105
R15810 GNDA.n2032 GNDA.n1987 3.4105
R15811 GNDA.n2032 GNDA.n1975 3.4105
R15812 GNDA.n2032 GNDA.n1988 3.4105
R15813 GNDA.n2032 GNDA.n1974 3.4105
R15814 GNDA.n2032 GNDA.n1989 3.4105
R15815 GNDA.n2032 GNDA.n1973 3.4105
R15816 GNDA.n2032 GNDA.n1990 3.4105
R15817 GNDA.n2032 GNDA.n1972 3.4105
R15818 GNDA.n2032 GNDA.n1991 3.4105
R15819 GNDA.n2032 GNDA.n1971 3.4105
R15820 GNDA.n2032 GNDA.n1992 3.4105
R15821 GNDA.n2032 GNDA.n1970 3.4105
R15822 GNDA.n2032 GNDA.n1993 3.4105
R15823 GNDA.n2032 GNDA.n1969 3.4105
R15824 GNDA.n2032 GNDA.n1994 3.4105
R15825 GNDA.n2032 GNDA.n1968 3.4105
R15826 GNDA.n2032 GNDA.n1995 3.4105
R15827 GNDA.n2245 GNDA.n2032 3.4105
R15828 GNDA.n2247 GNDA.n2032 3.4105
R15829 GNDA.n2006 GNDA.n1981 3.4105
R15830 GNDA.n2006 GNDA.n1982 3.4105
R15831 GNDA.n2006 GNDA.n1980 3.4105
R15832 GNDA.n2006 GNDA.n1983 3.4105
R15833 GNDA.n2006 GNDA.n1979 3.4105
R15834 GNDA.n2006 GNDA.n1984 3.4105
R15835 GNDA.n2006 GNDA.n1978 3.4105
R15836 GNDA.n2006 GNDA.n1985 3.4105
R15837 GNDA.n2006 GNDA.n1977 3.4105
R15838 GNDA.n2006 GNDA.n1986 3.4105
R15839 GNDA.n2006 GNDA.n1976 3.4105
R15840 GNDA.n2006 GNDA.n1987 3.4105
R15841 GNDA.n2006 GNDA.n1975 3.4105
R15842 GNDA.n2006 GNDA.n1988 3.4105
R15843 GNDA.n2006 GNDA.n1974 3.4105
R15844 GNDA.n2006 GNDA.n1989 3.4105
R15845 GNDA.n2006 GNDA.n1973 3.4105
R15846 GNDA.n2006 GNDA.n1990 3.4105
R15847 GNDA.n2006 GNDA.n1972 3.4105
R15848 GNDA.n2006 GNDA.n1991 3.4105
R15849 GNDA.n2006 GNDA.n1971 3.4105
R15850 GNDA.n2006 GNDA.n1992 3.4105
R15851 GNDA.n2006 GNDA.n1970 3.4105
R15852 GNDA.n2006 GNDA.n1993 3.4105
R15853 GNDA.n2006 GNDA.n1969 3.4105
R15854 GNDA.n2006 GNDA.n1994 3.4105
R15855 GNDA.n2006 GNDA.n1968 3.4105
R15856 GNDA.n2006 GNDA.n1995 3.4105
R15857 GNDA.n2245 GNDA.n2006 3.4105
R15858 GNDA.n2247 GNDA.n2006 3.4105
R15859 GNDA.n2033 GNDA.n1981 3.4105
R15860 GNDA.n2033 GNDA.n1982 3.4105
R15861 GNDA.n2033 GNDA.n1980 3.4105
R15862 GNDA.n2033 GNDA.n1983 3.4105
R15863 GNDA.n2033 GNDA.n1979 3.4105
R15864 GNDA.n2033 GNDA.n1984 3.4105
R15865 GNDA.n2033 GNDA.n1978 3.4105
R15866 GNDA.n2033 GNDA.n1985 3.4105
R15867 GNDA.n2033 GNDA.n1977 3.4105
R15868 GNDA.n2033 GNDA.n1986 3.4105
R15869 GNDA.n2033 GNDA.n1976 3.4105
R15870 GNDA.n2033 GNDA.n1987 3.4105
R15871 GNDA.n2033 GNDA.n1975 3.4105
R15872 GNDA.n2033 GNDA.n1988 3.4105
R15873 GNDA.n2033 GNDA.n1974 3.4105
R15874 GNDA.n2033 GNDA.n1989 3.4105
R15875 GNDA.n2033 GNDA.n1973 3.4105
R15876 GNDA.n2033 GNDA.n1990 3.4105
R15877 GNDA.n2033 GNDA.n1972 3.4105
R15878 GNDA.n2033 GNDA.n1991 3.4105
R15879 GNDA.n2033 GNDA.n1971 3.4105
R15880 GNDA.n2033 GNDA.n1992 3.4105
R15881 GNDA.n2033 GNDA.n1970 3.4105
R15882 GNDA.n2033 GNDA.n1993 3.4105
R15883 GNDA.n2033 GNDA.n1969 3.4105
R15884 GNDA.n2033 GNDA.n1994 3.4105
R15885 GNDA.n2033 GNDA.n1968 3.4105
R15886 GNDA.n2033 GNDA.n1995 3.4105
R15887 GNDA.n2245 GNDA.n2033 3.4105
R15888 GNDA.n2247 GNDA.n2033 3.4105
R15889 GNDA.n2005 GNDA.n1981 3.4105
R15890 GNDA.n2005 GNDA.n1982 3.4105
R15891 GNDA.n2005 GNDA.n1980 3.4105
R15892 GNDA.n2005 GNDA.n1983 3.4105
R15893 GNDA.n2005 GNDA.n1979 3.4105
R15894 GNDA.n2005 GNDA.n1984 3.4105
R15895 GNDA.n2005 GNDA.n1978 3.4105
R15896 GNDA.n2005 GNDA.n1985 3.4105
R15897 GNDA.n2005 GNDA.n1977 3.4105
R15898 GNDA.n2005 GNDA.n1986 3.4105
R15899 GNDA.n2005 GNDA.n1976 3.4105
R15900 GNDA.n2005 GNDA.n1987 3.4105
R15901 GNDA.n2005 GNDA.n1975 3.4105
R15902 GNDA.n2005 GNDA.n1988 3.4105
R15903 GNDA.n2005 GNDA.n1974 3.4105
R15904 GNDA.n2005 GNDA.n1989 3.4105
R15905 GNDA.n2005 GNDA.n1973 3.4105
R15906 GNDA.n2005 GNDA.n1990 3.4105
R15907 GNDA.n2005 GNDA.n1972 3.4105
R15908 GNDA.n2005 GNDA.n1991 3.4105
R15909 GNDA.n2005 GNDA.n1971 3.4105
R15910 GNDA.n2005 GNDA.n1992 3.4105
R15911 GNDA.n2005 GNDA.n1970 3.4105
R15912 GNDA.n2005 GNDA.n1993 3.4105
R15913 GNDA.n2005 GNDA.n1969 3.4105
R15914 GNDA.n2005 GNDA.n1994 3.4105
R15915 GNDA.n2005 GNDA.n1968 3.4105
R15916 GNDA.n2005 GNDA.n1995 3.4105
R15917 GNDA.n2245 GNDA.n2005 3.4105
R15918 GNDA.n2247 GNDA.n2005 3.4105
R15919 GNDA.n2034 GNDA.n1981 3.4105
R15920 GNDA.n2034 GNDA.n1982 3.4105
R15921 GNDA.n2034 GNDA.n1980 3.4105
R15922 GNDA.n2034 GNDA.n1983 3.4105
R15923 GNDA.n2034 GNDA.n1979 3.4105
R15924 GNDA.n2034 GNDA.n1984 3.4105
R15925 GNDA.n2034 GNDA.n1978 3.4105
R15926 GNDA.n2034 GNDA.n1985 3.4105
R15927 GNDA.n2034 GNDA.n1977 3.4105
R15928 GNDA.n2034 GNDA.n1986 3.4105
R15929 GNDA.n2034 GNDA.n1976 3.4105
R15930 GNDA.n2034 GNDA.n1987 3.4105
R15931 GNDA.n2034 GNDA.n1975 3.4105
R15932 GNDA.n2034 GNDA.n1988 3.4105
R15933 GNDA.n2034 GNDA.n1974 3.4105
R15934 GNDA.n2034 GNDA.n1989 3.4105
R15935 GNDA.n2034 GNDA.n1973 3.4105
R15936 GNDA.n2034 GNDA.n1990 3.4105
R15937 GNDA.n2034 GNDA.n1972 3.4105
R15938 GNDA.n2034 GNDA.n1991 3.4105
R15939 GNDA.n2034 GNDA.n1971 3.4105
R15940 GNDA.n2034 GNDA.n1992 3.4105
R15941 GNDA.n2034 GNDA.n1970 3.4105
R15942 GNDA.n2034 GNDA.n1993 3.4105
R15943 GNDA.n2034 GNDA.n1969 3.4105
R15944 GNDA.n2034 GNDA.n1994 3.4105
R15945 GNDA.n2034 GNDA.n1968 3.4105
R15946 GNDA.n2034 GNDA.n1995 3.4105
R15947 GNDA.n2245 GNDA.n2034 3.4105
R15948 GNDA.n2247 GNDA.n2034 3.4105
R15949 GNDA.n2004 GNDA.n1981 3.4105
R15950 GNDA.n2004 GNDA.n1982 3.4105
R15951 GNDA.n2004 GNDA.n1980 3.4105
R15952 GNDA.n2004 GNDA.n1983 3.4105
R15953 GNDA.n2004 GNDA.n1979 3.4105
R15954 GNDA.n2004 GNDA.n1984 3.4105
R15955 GNDA.n2004 GNDA.n1978 3.4105
R15956 GNDA.n2004 GNDA.n1985 3.4105
R15957 GNDA.n2004 GNDA.n1977 3.4105
R15958 GNDA.n2004 GNDA.n1986 3.4105
R15959 GNDA.n2004 GNDA.n1976 3.4105
R15960 GNDA.n2004 GNDA.n1987 3.4105
R15961 GNDA.n2004 GNDA.n1975 3.4105
R15962 GNDA.n2004 GNDA.n1988 3.4105
R15963 GNDA.n2004 GNDA.n1974 3.4105
R15964 GNDA.n2004 GNDA.n1989 3.4105
R15965 GNDA.n2004 GNDA.n1973 3.4105
R15966 GNDA.n2004 GNDA.n1990 3.4105
R15967 GNDA.n2004 GNDA.n1972 3.4105
R15968 GNDA.n2004 GNDA.n1991 3.4105
R15969 GNDA.n2004 GNDA.n1971 3.4105
R15970 GNDA.n2004 GNDA.n1992 3.4105
R15971 GNDA.n2004 GNDA.n1970 3.4105
R15972 GNDA.n2004 GNDA.n1993 3.4105
R15973 GNDA.n2004 GNDA.n1969 3.4105
R15974 GNDA.n2004 GNDA.n1994 3.4105
R15975 GNDA.n2004 GNDA.n1968 3.4105
R15976 GNDA.n2004 GNDA.n1995 3.4105
R15977 GNDA.n2245 GNDA.n2004 3.4105
R15978 GNDA.n2247 GNDA.n2004 3.4105
R15979 GNDA.n2035 GNDA.n1981 3.4105
R15980 GNDA.n2035 GNDA.n1982 3.4105
R15981 GNDA.n2035 GNDA.n1980 3.4105
R15982 GNDA.n2035 GNDA.n1983 3.4105
R15983 GNDA.n2035 GNDA.n1979 3.4105
R15984 GNDA.n2035 GNDA.n1984 3.4105
R15985 GNDA.n2035 GNDA.n1978 3.4105
R15986 GNDA.n2035 GNDA.n1985 3.4105
R15987 GNDA.n2035 GNDA.n1977 3.4105
R15988 GNDA.n2035 GNDA.n1986 3.4105
R15989 GNDA.n2035 GNDA.n1976 3.4105
R15990 GNDA.n2035 GNDA.n1987 3.4105
R15991 GNDA.n2035 GNDA.n1975 3.4105
R15992 GNDA.n2035 GNDA.n1988 3.4105
R15993 GNDA.n2035 GNDA.n1974 3.4105
R15994 GNDA.n2035 GNDA.n1989 3.4105
R15995 GNDA.n2035 GNDA.n1973 3.4105
R15996 GNDA.n2035 GNDA.n1990 3.4105
R15997 GNDA.n2035 GNDA.n1972 3.4105
R15998 GNDA.n2035 GNDA.n1991 3.4105
R15999 GNDA.n2035 GNDA.n1971 3.4105
R16000 GNDA.n2035 GNDA.n1992 3.4105
R16001 GNDA.n2035 GNDA.n1970 3.4105
R16002 GNDA.n2035 GNDA.n1993 3.4105
R16003 GNDA.n2035 GNDA.n1969 3.4105
R16004 GNDA.n2035 GNDA.n1994 3.4105
R16005 GNDA.n2035 GNDA.n1968 3.4105
R16006 GNDA.n2035 GNDA.n1995 3.4105
R16007 GNDA.n2245 GNDA.n2035 3.4105
R16008 GNDA.n2247 GNDA.n2035 3.4105
R16009 GNDA.n2003 GNDA.n1981 3.4105
R16010 GNDA.n2003 GNDA.n1982 3.4105
R16011 GNDA.n2003 GNDA.n1980 3.4105
R16012 GNDA.n2003 GNDA.n1983 3.4105
R16013 GNDA.n2003 GNDA.n1979 3.4105
R16014 GNDA.n2003 GNDA.n1984 3.4105
R16015 GNDA.n2003 GNDA.n1978 3.4105
R16016 GNDA.n2003 GNDA.n1985 3.4105
R16017 GNDA.n2003 GNDA.n1977 3.4105
R16018 GNDA.n2003 GNDA.n1986 3.4105
R16019 GNDA.n2003 GNDA.n1976 3.4105
R16020 GNDA.n2003 GNDA.n1987 3.4105
R16021 GNDA.n2003 GNDA.n1975 3.4105
R16022 GNDA.n2003 GNDA.n1988 3.4105
R16023 GNDA.n2003 GNDA.n1974 3.4105
R16024 GNDA.n2003 GNDA.n1989 3.4105
R16025 GNDA.n2003 GNDA.n1973 3.4105
R16026 GNDA.n2003 GNDA.n1990 3.4105
R16027 GNDA.n2003 GNDA.n1972 3.4105
R16028 GNDA.n2003 GNDA.n1991 3.4105
R16029 GNDA.n2003 GNDA.n1971 3.4105
R16030 GNDA.n2003 GNDA.n1992 3.4105
R16031 GNDA.n2003 GNDA.n1970 3.4105
R16032 GNDA.n2003 GNDA.n1993 3.4105
R16033 GNDA.n2003 GNDA.n1969 3.4105
R16034 GNDA.n2003 GNDA.n1994 3.4105
R16035 GNDA.n2003 GNDA.n1968 3.4105
R16036 GNDA.n2003 GNDA.n1995 3.4105
R16037 GNDA.n2245 GNDA.n2003 3.4105
R16038 GNDA.n2247 GNDA.n2003 3.4105
R16039 GNDA.n2036 GNDA.n1981 3.4105
R16040 GNDA.n2036 GNDA.n1982 3.4105
R16041 GNDA.n2036 GNDA.n1980 3.4105
R16042 GNDA.n2036 GNDA.n1983 3.4105
R16043 GNDA.n2036 GNDA.n1979 3.4105
R16044 GNDA.n2036 GNDA.n1984 3.4105
R16045 GNDA.n2036 GNDA.n1978 3.4105
R16046 GNDA.n2036 GNDA.n1985 3.4105
R16047 GNDA.n2036 GNDA.n1977 3.4105
R16048 GNDA.n2036 GNDA.n1986 3.4105
R16049 GNDA.n2036 GNDA.n1976 3.4105
R16050 GNDA.n2036 GNDA.n1987 3.4105
R16051 GNDA.n2036 GNDA.n1975 3.4105
R16052 GNDA.n2036 GNDA.n1988 3.4105
R16053 GNDA.n2036 GNDA.n1974 3.4105
R16054 GNDA.n2036 GNDA.n1989 3.4105
R16055 GNDA.n2036 GNDA.n1973 3.4105
R16056 GNDA.n2036 GNDA.n1990 3.4105
R16057 GNDA.n2036 GNDA.n1972 3.4105
R16058 GNDA.n2036 GNDA.n1991 3.4105
R16059 GNDA.n2036 GNDA.n1971 3.4105
R16060 GNDA.n2036 GNDA.n1992 3.4105
R16061 GNDA.n2036 GNDA.n1970 3.4105
R16062 GNDA.n2036 GNDA.n1993 3.4105
R16063 GNDA.n2036 GNDA.n1969 3.4105
R16064 GNDA.n2036 GNDA.n1994 3.4105
R16065 GNDA.n2036 GNDA.n1968 3.4105
R16066 GNDA.n2036 GNDA.n1995 3.4105
R16067 GNDA.n2245 GNDA.n2036 3.4105
R16068 GNDA.n2247 GNDA.n2036 3.4105
R16069 GNDA.n2002 GNDA.n1981 3.4105
R16070 GNDA.n2002 GNDA.n1982 3.4105
R16071 GNDA.n2002 GNDA.n1980 3.4105
R16072 GNDA.n2002 GNDA.n1983 3.4105
R16073 GNDA.n2002 GNDA.n1979 3.4105
R16074 GNDA.n2002 GNDA.n1984 3.4105
R16075 GNDA.n2002 GNDA.n1978 3.4105
R16076 GNDA.n2002 GNDA.n1985 3.4105
R16077 GNDA.n2002 GNDA.n1977 3.4105
R16078 GNDA.n2002 GNDA.n1986 3.4105
R16079 GNDA.n2002 GNDA.n1976 3.4105
R16080 GNDA.n2002 GNDA.n1987 3.4105
R16081 GNDA.n2002 GNDA.n1975 3.4105
R16082 GNDA.n2002 GNDA.n1988 3.4105
R16083 GNDA.n2002 GNDA.n1974 3.4105
R16084 GNDA.n2002 GNDA.n1989 3.4105
R16085 GNDA.n2002 GNDA.n1973 3.4105
R16086 GNDA.n2002 GNDA.n1990 3.4105
R16087 GNDA.n2002 GNDA.n1972 3.4105
R16088 GNDA.n2002 GNDA.n1991 3.4105
R16089 GNDA.n2002 GNDA.n1971 3.4105
R16090 GNDA.n2002 GNDA.n1992 3.4105
R16091 GNDA.n2002 GNDA.n1970 3.4105
R16092 GNDA.n2002 GNDA.n1993 3.4105
R16093 GNDA.n2002 GNDA.n1969 3.4105
R16094 GNDA.n2002 GNDA.n1994 3.4105
R16095 GNDA.n2002 GNDA.n1968 3.4105
R16096 GNDA.n2002 GNDA.n1995 3.4105
R16097 GNDA.n2245 GNDA.n2002 3.4105
R16098 GNDA.n2247 GNDA.n2002 3.4105
R16099 GNDA.n2037 GNDA.n1981 3.4105
R16100 GNDA.n2037 GNDA.n1982 3.4105
R16101 GNDA.n2037 GNDA.n1980 3.4105
R16102 GNDA.n2037 GNDA.n1983 3.4105
R16103 GNDA.n2037 GNDA.n1979 3.4105
R16104 GNDA.n2037 GNDA.n1984 3.4105
R16105 GNDA.n2037 GNDA.n1978 3.4105
R16106 GNDA.n2037 GNDA.n1985 3.4105
R16107 GNDA.n2037 GNDA.n1977 3.4105
R16108 GNDA.n2037 GNDA.n1986 3.4105
R16109 GNDA.n2037 GNDA.n1976 3.4105
R16110 GNDA.n2037 GNDA.n1987 3.4105
R16111 GNDA.n2037 GNDA.n1975 3.4105
R16112 GNDA.n2037 GNDA.n1988 3.4105
R16113 GNDA.n2037 GNDA.n1974 3.4105
R16114 GNDA.n2037 GNDA.n1989 3.4105
R16115 GNDA.n2037 GNDA.n1973 3.4105
R16116 GNDA.n2037 GNDA.n1990 3.4105
R16117 GNDA.n2037 GNDA.n1972 3.4105
R16118 GNDA.n2037 GNDA.n1991 3.4105
R16119 GNDA.n2037 GNDA.n1971 3.4105
R16120 GNDA.n2037 GNDA.n1992 3.4105
R16121 GNDA.n2037 GNDA.n1970 3.4105
R16122 GNDA.n2037 GNDA.n1993 3.4105
R16123 GNDA.n2037 GNDA.n1969 3.4105
R16124 GNDA.n2037 GNDA.n1994 3.4105
R16125 GNDA.n2037 GNDA.n1968 3.4105
R16126 GNDA.n2037 GNDA.n1995 3.4105
R16127 GNDA.n2245 GNDA.n2037 3.4105
R16128 GNDA.n2247 GNDA.n2037 3.4105
R16129 GNDA.n2001 GNDA.n1981 3.4105
R16130 GNDA.n2001 GNDA.n1982 3.4105
R16131 GNDA.n2001 GNDA.n1980 3.4105
R16132 GNDA.n2001 GNDA.n1983 3.4105
R16133 GNDA.n2001 GNDA.n1979 3.4105
R16134 GNDA.n2001 GNDA.n1984 3.4105
R16135 GNDA.n2001 GNDA.n1978 3.4105
R16136 GNDA.n2001 GNDA.n1985 3.4105
R16137 GNDA.n2001 GNDA.n1977 3.4105
R16138 GNDA.n2001 GNDA.n1986 3.4105
R16139 GNDA.n2001 GNDA.n1976 3.4105
R16140 GNDA.n2001 GNDA.n1987 3.4105
R16141 GNDA.n2001 GNDA.n1975 3.4105
R16142 GNDA.n2001 GNDA.n1988 3.4105
R16143 GNDA.n2001 GNDA.n1974 3.4105
R16144 GNDA.n2001 GNDA.n1989 3.4105
R16145 GNDA.n2001 GNDA.n1973 3.4105
R16146 GNDA.n2001 GNDA.n1990 3.4105
R16147 GNDA.n2001 GNDA.n1972 3.4105
R16148 GNDA.n2001 GNDA.n1991 3.4105
R16149 GNDA.n2001 GNDA.n1971 3.4105
R16150 GNDA.n2001 GNDA.n1992 3.4105
R16151 GNDA.n2001 GNDA.n1970 3.4105
R16152 GNDA.n2001 GNDA.n1993 3.4105
R16153 GNDA.n2001 GNDA.n1969 3.4105
R16154 GNDA.n2001 GNDA.n1994 3.4105
R16155 GNDA.n2001 GNDA.n1968 3.4105
R16156 GNDA.n2001 GNDA.n1995 3.4105
R16157 GNDA.n2245 GNDA.n2001 3.4105
R16158 GNDA.n2247 GNDA.n2001 3.4105
R16159 GNDA.n2038 GNDA.n1981 3.4105
R16160 GNDA.n2038 GNDA.n1982 3.4105
R16161 GNDA.n2038 GNDA.n1980 3.4105
R16162 GNDA.n2038 GNDA.n1983 3.4105
R16163 GNDA.n2038 GNDA.n1979 3.4105
R16164 GNDA.n2038 GNDA.n1984 3.4105
R16165 GNDA.n2038 GNDA.n1978 3.4105
R16166 GNDA.n2038 GNDA.n1985 3.4105
R16167 GNDA.n2038 GNDA.n1977 3.4105
R16168 GNDA.n2038 GNDA.n1986 3.4105
R16169 GNDA.n2038 GNDA.n1976 3.4105
R16170 GNDA.n2038 GNDA.n1987 3.4105
R16171 GNDA.n2038 GNDA.n1975 3.4105
R16172 GNDA.n2038 GNDA.n1988 3.4105
R16173 GNDA.n2038 GNDA.n1974 3.4105
R16174 GNDA.n2038 GNDA.n1989 3.4105
R16175 GNDA.n2038 GNDA.n1973 3.4105
R16176 GNDA.n2038 GNDA.n1990 3.4105
R16177 GNDA.n2038 GNDA.n1972 3.4105
R16178 GNDA.n2038 GNDA.n1991 3.4105
R16179 GNDA.n2038 GNDA.n1971 3.4105
R16180 GNDA.n2038 GNDA.n1992 3.4105
R16181 GNDA.n2038 GNDA.n1970 3.4105
R16182 GNDA.n2038 GNDA.n1993 3.4105
R16183 GNDA.n2038 GNDA.n1969 3.4105
R16184 GNDA.n2038 GNDA.n1994 3.4105
R16185 GNDA.n2038 GNDA.n1968 3.4105
R16186 GNDA.n2038 GNDA.n1995 3.4105
R16187 GNDA.n2245 GNDA.n2038 3.4105
R16188 GNDA.n2247 GNDA.n2038 3.4105
R16189 GNDA.n2000 GNDA.n1981 3.4105
R16190 GNDA.n2000 GNDA.n1982 3.4105
R16191 GNDA.n2000 GNDA.n1980 3.4105
R16192 GNDA.n2000 GNDA.n1983 3.4105
R16193 GNDA.n2000 GNDA.n1979 3.4105
R16194 GNDA.n2000 GNDA.n1984 3.4105
R16195 GNDA.n2000 GNDA.n1978 3.4105
R16196 GNDA.n2000 GNDA.n1985 3.4105
R16197 GNDA.n2000 GNDA.n1977 3.4105
R16198 GNDA.n2000 GNDA.n1986 3.4105
R16199 GNDA.n2000 GNDA.n1976 3.4105
R16200 GNDA.n2000 GNDA.n1987 3.4105
R16201 GNDA.n2000 GNDA.n1975 3.4105
R16202 GNDA.n2000 GNDA.n1988 3.4105
R16203 GNDA.n2000 GNDA.n1974 3.4105
R16204 GNDA.n2000 GNDA.n1989 3.4105
R16205 GNDA.n2000 GNDA.n1973 3.4105
R16206 GNDA.n2000 GNDA.n1990 3.4105
R16207 GNDA.n2000 GNDA.n1972 3.4105
R16208 GNDA.n2000 GNDA.n1991 3.4105
R16209 GNDA.n2000 GNDA.n1971 3.4105
R16210 GNDA.n2000 GNDA.n1992 3.4105
R16211 GNDA.n2000 GNDA.n1970 3.4105
R16212 GNDA.n2000 GNDA.n1993 3.4105
R16213 GNDA.n2000 GNDA.n1969 3.4105
R16214 GNDA.n2000 GNDA.n1994 3.4105
R16215 GNDA.n2000 GNDA.n1968 3.4105
R16216 GNDA.n2000 GNDA.n1995 3.4105
R16217 GNDA.n2245 GNDA.n2000 3.4105
R16218 GNDA.n2247 GNDA.n2000 3.4105
R16219 GNDA.n2039 GNDA.n1981 3.4105
R16220 GNDA.n2039 GNDA.n1982 3.4105
R16221 GNDA.n2039 GNDA.n1980 3.4105
R16222 GNDA.n2039 GNDA.n1983 3.4105
R16223 GNDA.n2039 GNDA.n1979 3.4105
R16224 GNDA.n2039 GNDA.n1984 3.4105
R16225 GNDA.n2039 GNDA.n1978 3.4105
R16226 GNDA.n2039 GNDA.n1985 3.4105
R16227 GNDA.n2039 GNDA.n1977 3.4105
R16228 GNDA.n2039 GNDA.n1986 3.4105
R16229 GNDA.n2039 GNDA.n1976 3.4105
R16230 GNDA.n2039 GNDA.n1987 3.4105
R16231 GNDA.n2039 GNDA.n1975 3.4105
R16232 GNDA.n2039 GNDA.n1988 3.4105
R16233 GNDA.n2039 GNDA.n1974 3.4105
R16234 GNDA.n2039 GNDA.n1989 3.4105
R16235 GNDA.n2039 GNDA.n1973 3.4105
R16236 GNDA.n2039 GNDA.n1990 3.4105
R16237 GNDA.n2039 GNDA.n1972 3.4105
R16238 GNDA.n2039 GNDA.n1991 3.4105
R16239 GNDA.n2039 GNDA.n1971 3.4105
R16240 GNDA.n2039 GNDA.n1992 3.4105
R16241 GNDA.n2039 GNDA.n1970 3.4105
R16242 GNDA.n2039 GNDA.n1993 3.4105
R16243 GNDA.n2039 GNDA.n1969 3.4105
R16244 GNDA.n2039 GNDA.n1994 3.4105
R16245 GNDA.n2039 GNDA.n1968 3.4105
R16246 GNDA.n2039 GNDA.n1995 3.4105
R16247 GNDA.n2245 GNDA.n2039 3.4105
R16248 GNDA.n2247 GNDA.n2039 3.4105
R16249 GNDA.n1999 GNDA.n1981 3.4105
R16250 GNDA.n1999 GNDA.n1982 3.4105
R16251 GNDA.n1999 GNDA.n1980 3.4105
R16252 GNDA.n1999 GNDA.n1983 3.4105
R16253 GNDA.n1999 GNDA.n1979 3.4105
R16254 GNDA.n1999 GNDA.n1984 3.4105
R16255 GNDA.n1999 GNDA.n1978 3.4105
R16256 GNDA.n1999 GNDA.n1985 3.4105
R16257 GNDA.n1999 GNDA.n1977 3.4105
R16258 GNDA.n1999 GNDA.n1986 3.4105
R16259 GNDA.n1999 GNDA.n1976 3.4105
R16260 GNDA.n1999 GNDA.n1987 3.4105
R16261 GNDA.n1999 GNDA.n1975 3.4105
R16262 GNDA.n1999 GNDA.n1988 3.4105
R16263 GNDA.n1999 GNDA.n1974 3.4105
R16264 GNDA.n1999 GNDA.n1989 3.4105
R16265 GNDA.n1999 GNDA.n1973 3.4105
R16266 GNDA.n1999 GNDA.n1990 3.4105
R16267 GNDA.n1999 GNDA.n1972 3.4105
R16268 GNDA.n1999 GNDA.n1991 3.4105
R16269 GNDA.n1999 GNDA.n1971 3.4105
R16270 GNDA.n1999 GNDA.n1992 3.4105
R16271 GNDA.n1999 GNDA.n1970 3.4105
R16272 GNDA.n1999 GNDA.n1993 3.4105
R16273 GNDA.n1999 GNDA.n1969 3.4105
R16274 GNDA.n1999 GNDA.n1994 3.4105
R16275 GNDA.n1999 GNDA.n1968 3.4105
R16276 GNDA.n1999 GNDA.n1995 3.4105
R16277 GNDA.n2245 GNDA.n1999 3.4105
R16278 GNDA.n2247 GNDA.n1999 3.4105
R16279 GNDA.n2040 GNDA.n1981 3.4105
R16280 GNDA.n2040 GNDA.n1982 3.4105
R16281 GNDA.n2040 GNDA.n1980 3.4105
R16282 GNDA.n2040 GNDA.n1983 3.4105
R16283 GNDA.n2040 GNDA.n1979 3.4105
R16284 GNDA.n2040 GNDA.n1984 3.4105
R16285 GNDA.n2040 GNDA.n1978 3.4105
R16286 GNDA.n2040 GNDA.n1985 3.4105
R16287 GNDA.n2040 GNDA.n1977 3.4105
R16288 GNDA.n2040 GNDA.n1986 3.4105
R16289 GNDA.n2040 GNDA.n1976 3.4105
R16290 GNDA.n2040 GNDA.n1987 3.4105
R16291 GNDA.n2040 GNDA.n1975 3.4105
R16292 GNDA.n2040 GNDA.n1988 3.4105
R16293 GNDA.n2040 GNDA.n1974 3.4105
R16294 GNDA.n2040 GNDA.n1989 3.4105
R16295 GNDA.n2040 GNDA.n1973 3.4105
R16296 GNDA.n2040 GNDA.n1990 3.4105
R16297 GNDA.n2040 GNDA.n1972 3.4105
R16298 GNDA.n2040 GNDA.n1991 3.4105
R16299 GNDA.n2040 GNDA.n1971 3.4105
R16300 GNDA.n2040 GNDA.n1992 3.4105
R16301 GNDA.n2040 GNDA.n1970 3.4105
R16302 GNDA.n2040 GNDA.n1993 3.4105
R16303 GNDA.n2040 GNDA.n1969 3.4105
R16304 GNDA.n2040 GNDA.n1994 3.4105
R16305 GNDA.n2040 GNDA.n1968 3.4105
R16306 GNDA.n2040 GNDA.n1995 3.4105
R16307 GNDA.n2245 GNDA.n2040 3.4105
R16308 GNDA.n2247 GNDA.n2040 3.4105
R16309 GNDA.n1998 GNDA.n1981 3.4105
R16310 GNDA.n1998 GNDA.n1982 3.4105
R16311 GNDA.n1998 GNDA.n1980 3.4105
R16312 GNDA.n1998 GNDA.n1983 3.4105
R16313 GNDA.n1998 GNDA.n1979 3.4105
R16314 GNDA.n1998 GNDA.n1984 3.4105
R16315 GNDA.n1998 GNDA.n1978 3.4105
R16316 GNDA.n1998 GNDA.n1985 3.4105
R16317 GNDA.n1998 GNDA.n1977 3.4105
R16318 GNDA.n1998 GNDA.n1986 3.4105
R16319 GNDA.n1998 GNDA.n1976 3.4105
R16320 GNDA.n1998 GNDA.n1987 3.4105
R16321 GNDA.n1998 GNDA.n1975 3.4105
R16322 GNDA.n1998 GNDA.n1988 3.4105
R16323 GNDA.n1998 GNDA.n1974 3.4105
R16324 GNDA.n1998 GNDA.n1989 3.4105
R16325 GNDA.n1998 GNDA.n1973 3.4105
R16326 GNDA.n1998 GNDA.n1990 3.4105
R16327 GNDA.n1998 GNDA.n1972 3.4105
R16328 GNDA.n1998 GNDA.n1991 3.4105
R16329 GNDA.n1998 GNDA.n1971 3.4105
R16330 GNDA.n1998 GNDA.n1992 3.4105
R16331 GNDA.n1998 GNDA.n1970 3.4105
R16332 GNDA.n1998 GNDA.n1993 3.4105
R16333 GNDA.n1998 GNDA.n1969 3.4105
R16334 GNDA.n1998 GNDA.n1994 3.4105
R16335 GNDA.n1998 GNDA.n1968 3.4105
R16336 GNDA.n1998 GNDA.n1995 3.4105
R16337 GNDA.n2245 GNDA.n1998 3.4105
R16338 GNDA.n2247 GNDA.n1998 3.4105
R16339 GNDA.n2246 GNDA.n1981 3.4105
R16340 GNDA.n2246 GNDA.n1982 3.4105
R16341 GNDA.n2246 GNDA.n1980 3.4105
R16342 GNDA.n2246 GNDA.n1983 3.4105
R16343 GNDA.n2246 GNDA.n1979 3.4105
R16344 GNDA.n2246 GNDA.n1984 3.4105
R16345 GNDA.n2246 GNDA.n1978 3.4105
R16346 GNDA.n2246 GNDA.n1985 3.4105
R16347 GNDA.n2246 GNDA.n1977 3.4105
R16348 GNDA.n2246 GNDA.n1986 3.4105
R16349 GNDA.n2246 GNDA.n1976 3.4105
R16350 GNDA.n2246 GNDA.n1987 3.4105
R16351 GNDA.n2246 GNDA.n1975 3.4105
R16352 GNDA.n2246 GNDA.n1988 3.4105
R16353 GNDA.n2246 GNDA.n1974 3.4105
R16354 GNDA.n2246 GNDA.n1989 3.4105
R16355 GNDA.n2246 GNDA.n1973 3.4105
R16356 GNDA.n2246 GNDA.n1990 3.4105
R16357 GNDA.n2246 GNDA.n1972 3.4105
R16358 GNDA.n2246 GNDA.n1991 3.4105
R16359 GNDA.n2246 GNDA.n1971 3.4105
R16360 GNDA.n2246 GNDA.n1992 3.4105
R16361 GNDA.n2246 GNDA.n1970 3.4105
R16362 GNDA.n2246 GNDA.n1993 3.4105
R16363 GNDA.n2246 GNDA.n1969 3.4105
R16364 GNDA.n2246 GNDA.n1994 3.4105
R16365 GNDA.n2246 GNDA.n1968 3.4105
R16366 GNDA.n2246 GNDA.n1995 3.4105
R16367 GNDA.n2246 GNDA.n2245 3.4105
R16368 GNDA.n2247 GNDA.n2246 3.4105
R16369 GNDA.n1997 GNDA.n1981 3.4105
R16370 GNDA.n1997 GNDA.n1982 3.4105
R16371 GNDA.n1997 GNDA.n1980 3.4105
R16372 GNDA.n1997 GNDA.n1983 3.4105
R16373 GNDA.n1997 GNDA.n1979 3.4105
R16374 GNDA.n1997 GNDA.n1984 3.4105
R16375 GNDA.n1997 GNDA.n1978 3.4105
R16376 GNDA.n1997 GNDA.n1985 3.4105
R16377 GNDA.n1997 GNDA.n1977 3.4105
R16378 GNDA.n1997 GNDA.n1986 3.4105
R16379 GNDA.n1997 GNDA.n1976 3.4105
R16380 GNDA.n1997 GNDA.n1987 3.4105
R16381 GNDA.n1997 GNDA.n1975 3.4105
R16382 GNDA.n1997 GNDA.n1988 3.4105
R16383 GNDA.n1997 GNDA.n1974 3.4105
R16384 GNDA.n1997 GNDA.n1989 3.4105
R16385 GNDA.n1997 GNDA.n1973 3.4105
R16386 GNDA.n1997 GNDA.n1990 3.4105
R16387 GNDA.n1997 GNDA.n1972 3.4105
R16388 GNDA.n1997 GNDA.n1991 3.4105
R16389 GNDA.n1997 GNDA.n1971 3.4105
R16390 GNDA.n1997 GNDA.n1992 3.4105
R16391 GNDA.n1997 GNDA.n1970 3.4105
R16392 GNDA.n1997 GNDA.n1993 3.4105
R16393 GNDA.n1997 GNDA.n1969 3.4105
R16394 GNDA.n1997 GNDA.n1994 3.4105
R16395 GNDA.n1997 GNDA.n1968 3.4105
R16396 GNDA.n1997 GNDA.n1995 3.4105
R16397 GNDA.n2245 GNDA.n1997 3.4105
R16398 GNDA.n2247 GNDA.n1997 3.4105
R16399 GNDA.n2248 GNDA.n1981 3.4105
R16400 GNDA.n2248 GNDA.n1982 3.4105
R16401 GNDA.n2248 GNDA.n1980 3.4105
R16402 GNDA.n2248 GNDA.n1983 3.4105
R16403 GNDA.n2248 GNDA.n1979 3.4105
R16404 GNDA.n2248 GNDA.n1984 3.4105
R16405 GNDA.n2248 GNDA.n1978 3.4105
R16406 GNDA.n2248 GNDA.n1985 3.4105
R16407 GNDA.n2248 GNDA.n1977 3.4105
R16408 GNDA.n2248 GNDA.n1986 3.4105
R16409 GNDA.n2248 GNDA.n1976 3.4105
R16410 GNDA.n2248 GNDA.n1987 3.4105
R16411 GNDA.n2248 GNDA.n1975 3.4105
R16412 GNDA.n2248 GNDA.n1988 3.4105
R16413 GNDA.n2248 GNDA.n1974 3.4105
R16414 GNDA.n2248 GNDA.n1989 3.4105
R16415 GNDA.n2248 GNDA.n1973 3.4105
R16416 GNDA.n2248 GNDA.n1990 3.4105
R16417 GNDA.n2248 GNDA.n1972 3.4105
R16418 GNDA.n2248 GNDA.n1991 3.4105
R16419 GNDA.n2248 GNDA.n1971 3.4105
R16420 GNDA.n2248 GNDA.n1992 3.4105
R16421 GNDA.n2248 GNDA.n1970 3.4105
R16422 GNDA.n2248 GNDA.n1993 3.4105
R16423 GNDA.n2248 GNDA.n1969 3.4105
R16424 GNDA.n2248 GNDA.n1994 3.4105
R16425 GNDA.n2248 GNDA.n1968 3.4105
R16426 GNDA.n2248 GNDA.n1995 3.4105
R16427 GNDA.n2248 GNDA.n2247 3.4105
R16428 GNDA.n4117 GNDA.n4116 3.39217
R16429 GNDA.n4113 GNDA.n1815 3.39217
R16430 GNDA.n4783 GNDA.n4782 3.39217
R16431 GNDA.n4128 GNDA.n4127 3.39217
R16432 GNDA.n1051 GNDA.n1049 3.32293
R16433 GNDA.n6192 GNDA.n599 3.32293
R16434 GNDA.t62 GNDA.n1331 3.32293
R16435 GNDA.t88 GNDA.n541 3.32293
R16436 GNDA.n4094 GNDA.n1831 3.313
R16437 GNDA.n4792 GNDA.n1349 3.313
R16438 GNDA.n4788 GNDA.n1590 3.13621
R16439 GNDA.n4788 GNDA.n4787 3.13621
R16440 GNDA.n4134 GNDA.n4131 3.13621
R16441 GNDA.n4135 GNDA.n4134 3.13621
R16442 GNDA.n6233 GNDA.n6232 2.86505
R16443 GNDA.n6234 GNDA.n6233 2.86505
R16444 GNDA.n6238 GNDA.n6236 2.86505
R16445 GNDA.n6241 GNDA.n6236 2.86505
R16446 GNDA.n6237 GNDA.n6234 2.86505
R16447 GNDA.n6241 GNDA.n6240 2.86505
R16448 GNDA.n6243 GNDA.n6232 2.86505
R16449 GNDA.n6238 GNDA.n6237 2.86505
R16450 GNDA.n954 GNDA.n952 2.86505
R16451 GNDA.n956 GNDA.n954 2.86505
R16452 GNDA.n956 GNDA.n955 2.86505
R16453 GNDA.n952 GNDA.n950 2.86505
R16454 GNDA.n1308 GNDA.n568 2.6629
R16455 GNDA.n6196 GNDA.n6195 2.6629
R16456 GNDA.n6226 GNDA.n6225 2.6629
R16457 GNDA.n7111 GNDA.n7110 2.6629
R16458 GNDA.n655 GNDA.n654 2.6629
R16459 GNDA.n782 GNDA.n781 2.6629
R16460 GNDA.n7040 GNDA.n7039 2.6629
R16461 GNDA.n6953 GNDA.n161 2.6629
R16462 GNDA.n7319 GNDA.n7318 2.6629
R16463 GNDA.n7232 GNDA.n82 2.6629
R16464 GNDA.n6896 GNDA.n6895 2.6629
R16465 GNDA.n6804 GNDA.n56 2.6629
R16466 GNDA.n1056 GNDA.n922 2.6629
R16467 GNDA.n6198 GNDA.n6197 2.6629
R16468 GNDA.n7226 GNDA.n7225 2.6629
R16469 GNDA.n6225 GNDA.n568 2.4581
R16470 GNDA.n1340 GNDA.n636 2.4581
R16471 GNDA.n6197 GNDA.n6196 2.4581
R16472 GNDA.n6226 GNDA.n567 2.4581
R16473 GNDA.n7111 GNDA.n161 2.4581
R16474 GNDA.n654 GNDA.n187 2.4581
R16475 GNDA.n781 GNDA.n655 2.4581
R16476 GNDA.n819 GNDA.n818 2.4581
R16477 GNDA.n6954 GNDA.n6953 2.4581
R16478 GNDA.n7319 GNDA.n56 2.4581
R16479 GNDA.n7233 GNDA.n7232 2.4581
R16480 GNDA.n6805 GNDA.n6804 2.4581
R16481 GNDA.n6199 GNDA.n6198 2.4581
R16482 GNDA.n7226 GNDA.n82 2.4581
R16483 GNDA.n7159 GNDA.n7158 2.4581
R16484 GNDA.n6353 GNDA.n6352 2.39683
R16485 GNDA.n413 GNDA.n412 2.39683
R16486 GNDA.n5400 GNDA.n5399 2.3951
R16487 GNDA.n5402 GNDA.n5401 2.3951
R16488 GNDA.n5544 GNDA.n1362 2.3951
R16489 GNDA.n6086 GNDA.n1363 2.3951
R16490 GNDA.n4807 GNDA.n4806 2.3951
R16491 GNDA.n4521 GNDA.n1592 2.3951
R16492 GNDA.n4332 GNDA.n1591 2.3951
R16493 GNDA.n4166 GNDA.n4165 2.3951
R16494 GNDA.n4164 GNDA.n1813 2.3951
R16495 GNDA.n3823 GNDA.n1814 2.3951
R16496 GNDA.n4081 GNDA.n4080 2.3951
R16497 GNDA.n3468 GNDA.n3467 2.3951
R16498 GNDA.n3293 GNDA.n1887 2.3951
R16499 GNDA.n3291 GNDA.n1889 2.3951
R16500 GNDA.n3290 GNDA.n1890 2.3951
R16501 GNDA.n3289 GNDA.n1891 2.3951
R16502 GNDA.n4773 GNDA.n4772 2.30736
R16503 GNDA.n5800 GNDA.n5799 2.30736
R16504 GNDA.n6078 GNDA.n6077 2.30736
R16505 GNDA.n1514 GNDA.n1513 2.30736
R16506 GNDA.n3749 GNDA.n3748 2.30736
R16507 GNDA.n3386 GNDA.n3385 2.30736
R16508 GNDA.n5229 GNDA.n5228 2.30736
R16509 GNDA.n5326 GNDA.n5325 2.30736
R16510 GNDA.n5517 GNDA.n5516 2.30736
R16511 GNDA.n5659 GNDA.n5658 2.30736
R16512 GNDA.n5941 GNDA.n5940 2.30736
R16513 GNDA.n4922 GNDA.n4921 2.30736
R16514 GNDA.n4636 GNDA.n4635 2.30736
R16515 GNDA.n4447 GNDA.n4446 2.30736
R16516 GNDA.n4281 GNDA.n4280 2.30736
R16517 GNDA.n1740 GNDA.n1739 2.30736
R16518 GNDA.n3938 GNDA.n3937 2.30736
R16519 GNDA.n4075 GNDA.n4074 2.30736
R16520 GNDA.n3583 GNDA.n3582 2.30736
R16521 GNDA.n2648 GNDA.n2647 2.30736
R16522 GNDA.n2931 GNDA.n2930 2.30736
R16523 GNDA.n3072 GNDA.n3071 2.30736
R16524 GNDA.n3213 GNDA.n3212 2.30736
R16525 GNDA.n3218 GNDA.n1947 2.30736
R16526 GNDA.n2790 GNDA.n2789 2.30736
R16527 GNDA.n1588 GNDA.n1422 2.251
R16528 GNDA.n3460 GNDA.n3294 2.251
R16529 GNDA.n4082 GNDA.n1832 2.251
R16530 GNDA.n6085 GNDA.n6084 2.251
R16531 GNDA.n4115 GNDA.n4114 2.2505
R16532 GNDA.n4162 GNDA.n4139 2.19633
R16533 GNDA.n4120 GNDA.n4119 2.19633
R16534 GNDA.n4125 GNDA.n4124 2.19633
R16535 GNDA.n329 GNDA.n56 2.18124
R16536 GNDA.n7115 GNDA.n161 2.18124
R16537 GNDA.n6197 GNDA.n587 2.18124
R16538 GNDA.n6651 GNDA.n82 2.18124
R16539 GNDA.n901 GNDA.n655 2.18124
R16540 GNDA.n6225 GNDA.n569 2.18124
R16541 GNDA.n636 GNDA.n546 2.1509
R16542 GNDA.n620 GNDA.n567 2.1509
R16543 GNDA.n7046 GNDA.n187 2.1509
R16544 GNDA.n818 GNDA.n817 2.1509
R16545 GNDA.n6972 GNDA.n6954 2.1509
R16546 GNDA.n7251 GNDA.n7233 2.1509
R16547 GNDA.n6831 GNDA.n6805 2.1509
R16548 GNDA.n6200 GNDA.n6199 2.1509
R16549 GNDA.n7169 GNDA.n7159 2.1509
R16550 GNDA.n1309 GNDA.n1308 2.13383
R16551 GNDA.n6195 GNDA.n595 2.13383
R16552 GNDA.n7110 GNDA.n165 2.13383
R16553 GNDA.n6895 GNDA.n6782 2.13383
R16554 GNDA.n782 GNDA.n780 2.13383
R16555 GNDA.n7039 GNDA.n6926 2.13383
R16556 GNDA.n7318 GNDA.n57 2.13383
R16557 GNDA.n1037 GNDA.n922 2.13383
R16558 GNDA.n7225 GNDA.n7224 2.13383
R16559 GNDA.n1366 GNDA.n1365 2.09414
R16560 GNDA.n4801 GNDA.n4800 2.09414
R16561 GNDA.n4086 GNDA.n4085 2.09414
R16562 GNDA.n3462 GNDA.n3461 2.09414
R16563 GNDA.n134 GNDA.n56 2.08643
R16564 GNDA.n163 GNDA.n161 2.08643
R16565 GNDA.n6197 GNDA.n584 2.08643
R16566 GNDA.n84 GNDA.n82 2.08643
R16567 GNDA.n904 GNDA.n655 2.08643
R16568 GNDA.n6225 GNDA.n6224 2.08643
R16569 GNDA.n1308 GNDA.n1307 1.9461
R16570 GNDA.n6195 GNDA.n6194 1.9461
R16571 GNDA.n7110 GNDA.n7109 1.9461
R16572 GNDA.n783 GNDA.n782 1.9461
R16573 GNDA.n7039 GNDA.n7038 1.9461
R16574 GNDA.n7318 GNDA.n7317 1.9461
R16575 GNDA.n6895 GNDA.n6894 1.9461
R16576 GNDA.n924 GNDA.n922 1.9461
R16577 GNDA.n7225 GNDA.n22 1.9461
R16578 GNDA.n6092 GNDA.n6091 1.93383
R16579 GNDA.n4797 GNDA.n4796 1.93383
R16580 GNDA.n4093 GNDA.n4092 1.93383
R16581 GNDA.n4097 GNDA.n4096 1.93383
R16582 GNDA.n1595 GNDA.n1594 1.91062
R16583 GNDA.n6620 GNDA.n6619 1.90675
R16584 GNDA.t107 GNDA.t93 1.83536
R16585 GNDA.n4129 GNDA.t45 1.83536
R16586 GNDA.n4785 GNDA.t832 1.83536
R16587 GNDA.n4784 GNDA.t101 1.83536
R16588 GNDA.t853 GNDA.t139 1.83536
R16589 GNDA.n4791 GNDA.n1589 1.7505
R16590 GNDA.n2165 GNDA.n2164 1.70567
R16591 GNDA.n2182 GNDA.n2164 1.70567
R16592 GNDA.n2185 GNDA.n2164 1.70567
R16593 GNDA.n2188 GNDA.n2164 1.70567
R16594 GNDA.n2191 GNDA.n2164 1.70567
R16595 GNDA.n2194 GNDA.n2164 1.70567
R16596 GNDA.n2197 GNDA.n2164 1.70567
R16597 GNDA.n2200 GNDA.n2164 1.70567
R16598 GNDA.n2203 GNDA.n2164 1.70567
R16599 GNDA.n2206 GNDA.n2164 1.70567
R16600 GNDA.n2209 GNDA.n2164 1.70567
R16601 GNDA.n2212 GNDA.n2164 1.70567
R16602 GNDA.n2215 GNDA.n2164 1.70567
R16603 GNDA.n2218 GNDA.n2164 1.70567
R16604 GNDA.n2221 GNDA.n2164 1.70567
R16605 GNDA.n2164 GNDA.n2105 1.70567
R16606 GNDA.n2321 GNDA.n2320 1.70567
R16607 GNDA.n2320 GNDA.n2306 1.70567
R16608 GNDA.n2320 GNDA.n2307 1.70567
R16609 GNDA.n2320 GNDA.n2308 1.70567
R16610 GNDA.n2320 GNDA.n2309 1.70567
R16611 GNDA.n2320 GNDA.n2310 1.70567
R16612 GNDA.n2320 GNDA.n2311 1.70567
R16613 GNDA.n2320 GNDA.n2312 1.70567
R16614 GNDA.n2320 GNDA.n2313 1.70567
R16615 GNDA.n2320 GNDA.n2314 1.70567
R16616 GNDA.n2320 GNDA.n2315 1.70567
R16617 GNDA.n2320 GNDA.n2316 1.70567
R16618 GNDA.n2320 GNDA.n2317 1.70567
R16619 GNDA.n2320 GNDA.n2318 1.70567
R16620 GNDA.n2320 GNDA.n2319 1.70567
R16621 GNDA.n2320 GNDA.n2264 1.70567
R16622 GNDA.n2242 GNDA.n1982 1.70567
R16623 GNDA.n2072 GNDA.n2059 1.70567
R16624 GNDA.n2072 GNDA.n2060 1.70567
R16625 GNDA.n2072 GNDA.n2061 1.70567
R16626 GNDA.n2072 GNDA.n2062 1.70567
R16627 GNDA.n2072 GNDA.n2063 1.70567
R16628 GNDA.n2072 GNDA.n2064 1.70567
R16629 GNDA.n2072 GNDA.n2065 1.70567
R16630 GNDA.n2072 GNDA.n2066 1.70567
R16631 GNDA.n2072 GNDA.n2067 1.70567
R16632 GNDA.n2072 GNDA.n2068 1.70567
R16633 GNDA.n2072 GNDA.n2069 1.70567
R16634 GNDA.n2072 GNDA.n2070 1.70567
R16635 GNDA.n2072 GNDA.n2071 1.70567
R16636 GNDA.n2072 GNDA.n2041 1.70567
R16637 GNDA.n2072 GNDA.n1967 1.70567
R16638 GNDA.n2223 GNDA.n2163 1.70565
R16639 GNDA.n2163 GNDA.n2161 1.70565
R16640 GNDA.n2163 GNDA.n2159 1.70565
R16641 GNDA.n2163 GNDA.n2157 1.70565
R16642 GNDA.n2163 GNDA.n2155 1.70565
R16643 GNDA.n2163 GNDA.n2153 1.70565
R16644 GNDA.n2163 GNDA.n2151 1.70565
R16645 GNDA.n2181 GNDA.n2177 1.70565
R16646 GNDA.n2181 GNDA.n2176 1.70565
R16647 GNDA.n2181 GNDA.n2173 1.70565
R16648 GNDA.n2181 GNDA.n2172 1.70565
R16649 GNDA.n2181 GNDA.n2169 1.70565
R16650 GNDA.n2181 GNDA.n2168 1.70565
R16651 GNDA.n2227 GNDA.n2120 1.70565
R16652 GNDA.n2279 GNDA.n2249 1.70565
R16653 GNDA.n2283 GNDA.n2249 1.70565
R16654 GNDA.n2287 GNDA.n2249 1.70565
R16655 GNDA.n2291 GNDA.n2249 1.70565
R16656 GNDA.n2295 GNDA.n2249 1.70565
R16657 GNDA.n2299 GNDA.n2249 1.70565
R16658 GNDA.n2303 GNDA.n2249 1.70565
R16659 GNDA.n2353 GNDA.n1951 1.70565
R16660 GNDA.n2353 GNDA.n2349 1.70565
R16661 GNDA.n2353 GNDA.n2348 1.70565
R16662 GNDA.n2353 GNDA.n2345 1.70565
R16663 GNDA.n2353 GNDA.n2344 1.70565
R16664 GNDA.n2353 GNDA.n2341 1.70565
R16665 GNDA.n2353 GNDA.n2340 1.70565
R16666 GNDA.n2243 GNDA.n2239 1.70565
R16667 GNDA.n2243 GNDA.n2238 1.70565
R16668 GNDA.n2243 GNDA.n2235 1.70565
R16669 GNDA.n2243 GNDA.n2234 1.70565
R16670 GNDA.n2243 GNDA.n2231 1.70565
R16671 GNDA.n2243 GNDA.n2230 1.70565
R16672 GNDA.n2243 GNDA.n2013 1.70565
R16673 GNDA.n2026 GNDA.n2024 1.70565
R16674 GNDA.n2026 GNDA.n2022 1.70565
R16675 GNDA.n2026 GNDA.n2020 1.70565
R16676 GNDA.n2026 GNDA.n2018 1.70565
R16677 GNDA.n2026 GNDA.n2016 1.70565
R16678 GNDA.n2026 GNDA.n2014 1.70565
R16679 GNDA.n2012 GNDA.n2011 1.70565
R16680 GNDA.n2028 GNDA.n2027 1.70565
R16681 GNDA.n2248 GNDA.n1996 1.70565
R16682 GNDA.n2163 GNDA.n2162 1.70563
R16683 GNDA.n2163 GNDA.n2158 1.70563
R16684 GNDA.n2163 GNDA.n2154 1.70563
R16685 GNDA.n2163 GNDA.n2150 1.70563
R16686 GNDA.n2181 GNDA.n2179 1.70563
R16687 GNDA.n2181 GNDA.n2178 1.70563
R16688 GNDA.n2181 GNDA.n2175 1.70563
R16689 GNDA.n2181 GNDA.n2174 1.70563
R16690 GNDA.n2181 GNDA.n2171 1.70563
R16691 GNDA.n2181 GNDA.n2170 1.70563
R16692 GNDA.n2181 GNDA.n2167 1.70563
R16693 GNDA.n2181 GNDA.n2166 1.70563
R16694 GNDA.n2180 GNDA.n361 1.70563
R16695 GNDA.n2186 GNDA.n361 1.70563
R16696 GNDA.n2192 GNDA.n361 1.70563
R16697 GNDA.n2198 GNDA.n361 1.70563
R16698 GNDA.n2204 GNDA.n361 1.70563
R16699 GNDA.n2210 GNDA.n361 1.70563
R16700 GNDA.n2216 GNDA.n361 1.70563
R16701 GNDA.n2222 GNDA.n361 1.70563
R16702 GNDA.n2281 GNDA.n2249 1.70563
R16703 GNDA.n2289 GNDA.n2249 1.70563
R16704 GNDA.n2297 GNDA.n2249 1.70563
R16705 GNDA.n2336 GNDA.n2249 1.70563
R16706 GNDA.n2353 GNDA.n2351 1.70563
R16707 GNDA.n2353 GNDA.n2350 1.70563
R16708 GNDA.n2353 GNDA.n2347 1.70563
R16709 GNDA.n2353 GNDA.n2346 1.70563
R16710 GNDA.n2353 GNDA.n2343 1.70563
R16711 GNDA.n2353 GNDA.n2342 1.70563
R16712 GNDA.n2353 GNDA.n2339 1.70563
R16713 GNDA.n2338 GNDA.n2337 1.70563
R16714 GNDA.n2337 GNDA.n2334 1.70563
R16715 GNDA.n2337 GNDA.n2332 1.70563
R16716 GNDA.n2337 GNDA.n2330 1.70563
R16717 GNDA.n2337 GNDA.n2328 1.70563
R16718 GNDA.n2337 GNDA.n2326 1.70563
R16719 GNDA.n2337 GNDA.n2324 1.70563
R16720 GNDA.n2337 GNDA.n2322 1.70563
R16721 GNDA.n2355 GNDA.n2265 1.70563
R16722 GNDA.n2243 GNDA.n2241 1.70563
R16723 GNDA.n2243 GNDA.n2240 1.70563
R16724 GNDA.n2243 GNDA.n2237 1.70563
R16725 GNDA.n2243 GNDA.n2236 1.70563
R16726 GNDA.n2243 GNDA.n2233 1.70563
R16727 GNDA.n2243 GNDA.n2232 1.70563
R16728 GNDA.n2243 GNDA.n2229 1.70563
R16729 GNDA.n2244 GNDA.n2243 1.70563
R16730 GNDA.n2026 GNDA.n2025 1.70563
R16731 GNDA.n2026 GNDA.n2021 1.70563
R16732 GNDA.n2026 GNDA.n2017 1.70563
R16733 GNDA.n2058 GNDA.n2026 1.70563
R16734 GNDA.n2056 GNDA.n2055 1.70563
R16735 GNDA.n2056 GNDA.n2053 1.70563
R16736 GNDA.n2056 GNDA.n2051 1.70563
R16737 GNDA.n2056 GNDA.n2049 1.70563
R16738 GNDA.n2056 GNDA.n2047 1.70563
R16739 GNDA.n2056 GNDA.n2045 1.70563
R16740 GNDA.n2056 GNDA.n2043 1.70563
R16741 GNDA.n2057 GNDA.n2056 1.70563
R16742 GNDA.n2163 GNDA.n2160 1.70556
R16743 GNDA.n2163 GNDA.n2156 1.70556
R16744 GNDA.n2163 GNDA.n2152 1.70556
R16745 GNDA.n2183 GNDA.n361 1.70556
R16746 GNDA.n2189 GNDA.n361 1.70556
R16747 GNDA.n2195 GNDA.n361 1.70556
R16748 GNDA.n2201 GNDA.n361 1.70556
R16749 GNDA.n2207 GNDA.n361 1.70556
R16750 GNDA.n2213 GNDA.n361 1.70556
R16751 GNDA.n2219 GNDA.n361 1.70556
R16752 GNDA.n2285 GNDA.n2249 1.70556
R16753 GNDA.n2293 GNDA.n2249 1.70556
R16754 GNDA.n2301 GNDA.n2249 1.70556
R16755 GNDA.n2337 GNDA.n2335 1.70556
R16756 GNDA.n2337 GNDA.n2333 1.70556
R16757 GNDA.n2337 GNDA.n2331 1.70556
R16758 GNDA.n2337 GNDA.n2329 1.70556
R16759 GNDA.n2337 GNDA.n2327 1.70556
R16760 GNDA.n2337 GNDA.n2325 1.70556
R16761 GNDA.n2337 GNDA.n2323 1.70556
R16762 GNDA.n2026 GNDA.n2023 1.70556
R16763 GNDA.n2026 GNDA.n2019 1.70556
R16764 GNDA.n2026 GNDA.n2015 1.70556
R16765 GNDA.n2056 GNDA.n2054 1.70556
R16766 GNDA.n2056 GNDA.n2052 1.70556
R16767 GNDA.n2056 GNDA.n2050 1.70556
R16768 GNDA.n2056 GNDA.n2048 1.70556
R16769 GNDA.n2056 GNDA.n2046 1.70556
R16770 GNDA.n2056 GNDA.n2044 1.70556
R16771 GNDA.n2056 GNDA.n2042 1.70556
R16772 GNDA.n3215 GNDA.n2411 1.69433
R16773 GNDA.n3215 GNDA.n2408 1.69433
R16774 GNDA.n3215 GNDA.n2405 1.69433
R16775 GNDA.n3215 GNDA.n2402 1.69433
R16776 GNDA.n3215 GNDA.n2399 1.69433
R16777 GNDA.n3215 GNDA.n2396 1.69433
R16778 GNDA.n3215 GNDA.n2393 1.69433
R16779 GNDA.n3074 GNDA.n2435 1.69433
R16780 GNDA.n3074 GNDA.n2432 1.69433
R16781 GNDA.n3074 GNDA.n2429 1.69433
R16782 GNDA.n3074 GNDA.n2426 1.69433
R16783 GNDA.n3074 GNDA.n2423 1.69433
R16784 GNDA.n3074 GNDA.n2420 1.69433
R16785 GNDA.n3074 GNDA.n2417 1.69433
R16786 GNDA.n2933 GNDA.n2459 1.69433
R16787 GNDA.n2933 GNDA.n2456 1.69433
R16788 GNDA.n2933 GNDA.n2453 1.69433
R16789 GNDA.n2933 GNDA.n2450 1.69433
R16790 GNDA.n2933 GNDA.n2447 1.69433
R16791 GNDA.n2933 GNDA.n2444 1.69433
R16792 GNDA.n2933 GNDA.n2441 1.69433
R16793 GNDA.n2650 GNDA.n2507 1.69433
R16794 GNDA.n2650 GNDA.n2504 1.69433
R16795 GNDA.n2650 GNDA.n2501 1.69433
R16796 GNDA.n2650 GNDA.n2498 1.69433
R16797 GNDA.n2650 GNDA.n2495 1.69433
R16798 GNDA.n2650 GNDA.n2492 1.69433
R16799 GNDA.n2650 GNDA.n2489 1.69433
R16800 GNDA.n3585 GNDA.n1860 1.69433
R16801 GNDA.n3585 GNDA.n1857 1.69433
R16802 GNDA.n3585 GNDA.n1854 1.69433
R16803 GNDA.n3585 GNDA.n1851 1.69433
R16804 GNDA.n3585 GNDA.n1848 1.69433
R16805 GNDA.n3585 GNDA.n1845 1.69433
R16806 GNDA.n3585 GNDA.n1842 1.69433
R16807 GNDA.n4077 GNDA.n3772 1.69433
R16808 GNDA.n4077 GNDA.n3769 1.69433
R16809 GNDA.n4077 GNDA.n3766 1.69433
R16810 GNDA.n4077 GNDA.n3763 1.69433
R16811 GNDA.n4077 GNDA.n3760 1.69433
R16812 GNDA.n4077 GNDA.n3757 1.69433
R16813 GNDA.n4077 GNDA.n3754 1.69433
R16814 GNDA.n3940 GNDA.n3796 1.69433
R16815 GNDA.n3940 GNDA.n3793 1.69433
R16816 GNDA.n3940 GNDA.n3790 1.69433
R16817 GNDA.n3940 GNDA.n3787 1.69433
R16818 GNDA.n3940 GNDA.n3784 1.69433
R16819 GNDA.n3940 GNDA.n3781 1.69433
R16820 GNDA.n3940 GNDA.n3778 1.69433
R16821 GNDA.n1749 GNDA.n1599 1.69433
R16822 GNDA.n1758 GNDA.n1599 1.69433
R16823 GNDA.n1767 GNDA.n1599 1.69433
R16824 GNDA.n1776 GNDA.n1599 1.69433
R16825 GNDA.n1785 GNDA.n1599 1.69433
R16826 GNDA.n1794 GNDA.n1599 1.69433
R16827 GNDA.n1803 GNDA.n1599 1.69433
R16828 GNDA.n4283 GNDA.n1621 1.69433
R16829 GNDA.n4283 GNDA.n1618 1.69433
R16830 GNDA.n4283 GNDA.n1615 1.69433
R16831 GNDA.n4283 GNDA.n1612 1.69433
R16832 GNDA.n4283 GNDA.n1609 1.69433
R16833 GNDA.n4283 GNDA.n1606 1.69433
R16834 GNDA.n4283 GNDA.n1603 1.69433
R16835 GNDA.n4449 GNDA.n4305 1.69433
R16836 GNDA.n4449 GNDA.n4302 1.69433
R16837 GNDA.n4449 GNDA.n4299 1.69433
R16838 GNDA.n4449 GNDA.n4296 1.69433
R16839 GNDA.n4449 GNDA.n4293 1.69433
R16840 GNDA.n4449 GNDA.n4290 1.69433
R16841 GNDA.n4449 GNDA.n4287 1.69433
R16842 GNDA.n4638 GNDA.n4494 1.69433
R16843 GNDA.n4638 GNDA.n4491 1.69433
R16844 GNDA.n4638 GNDA.n4488 1.69433
R16845 GNDA.n4638 GNDA.n4485 1.69433
R16846 GNDA.n4638 GNDA.n4482 1.69433
R16847 GNDA.n4638 GNDA.n4479 1.69433
R16848 GNDA.n4638 GNDA.n4476 1.69433
R16849 GNDA.n4924 GNDA.n1393 1.69433
R16850 GNDA.n4924 GNDA.n1390 1.69433
R16851 GNDA.n4924 GNDA.n1387 1.69433
R16852 GNDA.n4924 GNDA.n1384 1.69433
R16853 GNDA.n4924 GNDA.n1381 1.69433
R16854 GNDA.n4924 GNDA.n1378 1.69433
R16855 GNDA.n4924 GNDA.n1375 1.69433
R16856 GNDA.n5943 GNDA.n4969 1.69433
R16857 GNDA.n5943 GNDA.n4966 1.69433
R16858 GNDA.n5943 GNDA.n4963 1.69433
R16859 GNDA.n5943 GNDA.n4960 1.69433
R16860 GNDA.n5943 GNDA.n4957 1.69433
R16861 GNDA.n5943 GNDA.n4954 1.69433
R16862 GNDA.n5943 GNDA.n4951 1.69433
R16863 GNDA.n5661 GNDA.n5017 1.69433
R16864 GNDA.n5661 GNDA.n5014 1.69433
R16865 GNDA.n5661 GNDA.n5011 1.69433
R16866 GNDA.n5661 GNDA.n5008 1.69433
R16867 GNDA.n5661 GNDA.n5005 1.69433
R16868 GNDA.n5661 GNDA.n5002 1.69433
R16869 GNDA.n5661 GNDA.n4999 1.69433
R16870 GNDA.n5519 GNDA.n5041 1.69433
R16871 GNDA.n5519 GNDA.n5038 1.69433
R16872 GNDA.n5519 GNDA.n5035 1.69433
R16873 GNDA.n5519 GNDA.n5032 1.69433
R16874 GNDA.n5519 GNDA.n5029 1.69433
R16875 GNDA.n5519 GNDA.n5026 1.69433
R16876 GNDA.n5519 GNDA.n5023 1.69433
R16877 GNDA.n5335 GNDA.n5044 1.69433
R16878 GNDA.n5344 GNDA.n5044 1.69433
R16879 GNDA.n5353 GNDA.n5044 1.69433
R16880 GNDA.n5362 GNDA.n5044 1.69433
R16881 GNDA.n5371 GNDA.n5044 1.69433
R16882 GNDA.n5380 GNDA.n5044 1.69433
R16883 GNDA.n5389 GNDA.n5044 1.69433
R16884 GNDA.n5231 GNDA.n5092 1.69433
R16885 GNDA.n5231 GNDA.n5089 1.69433
R16886 GNDA.n5231 GNDA.n5086 1.69433
R16887 GNDA.n5231 GNDA.n5083 1.69433
R16888 GNDA.n5231 GNDA.n5080 1.69433
R16889 GNDA.n5231 GNDA.n5077 1.69433
R16890 GNDA.n5231 GNDA.n5074 1.69433
R16891 GNDA.n3395 GNDA.n1838 1.69433
R16892 GNDA.n3404 GNDA.n1838 1.69433
R16893 GNDA.n3413 GNDA.n1838 1.69433
R16894 GNDA.n3422 GNDA.n1838 1.69433
R16895 GNDA.n3431 GNDA.n1838 1.69433
R16896 GNDA.n3440 GNDA.n1838 1.69433
R16897 GNDA.n3449 GNDA.n1838 1.69433
R16898 GNDA.n3751 GNDA.n3607 1.69433
R16899 GNDA.n3751 GNDA.n3604 1.69433
R16900 GNDA.n3751 GNDA.n3601 1.69433
R16901 GNDA.n3751 GNDA.n3598 1.69433
R16902 GNDA.n3751 GNDA.n3595 1.69433
R16903 GNDA.n3751 GNDA.n3592 1.69433
R16904 GNDA.n3751 GNDA.n3589 1.69433
R16905 GNDA.n1523 GNDA.n1371 1.69433
R16906 GNDA.n1532 GNDA.n1371 1.69433
R16907 GNDA.n1541 GNDA.n1371 1.69433
R16908 GNDA.n1550 GNDA.n1371 1.69433
R16909 GNDA.n1559 GNDA.n1371 1.69433
R16910 GNDA.n1568 GNDA.n1371 1.69433
R16911 GNDA.n1577 GNDA.n1371 1.69433
R16912 GNDA.n6080 GNDA.n4945 1.69433
R16913 GNDA.n6080 GNDA.n4942 1.69433
R16914 GNDA.n6080 GNDA.n4939 1.69433
R16915 GNDA.n6080 GNDA.n4936 1.69433
R16916 GNDA.n6080 GNDA.n4933 1.69433
R16917 GNDA.n6080 GNDA.n4930 1.69433
R16918 GNDA.n6080 GNDA.n4927 1.69433
R16919 GNDA.n2792 GNDA.n2483 1.69433
R16920 GNDA.n2792 GNDA.n2480 1.69433
R16921 GNDA.n2792 GNDA.n2477 1.69433
R16922 GNDA.n2792 GNDA.n2474 1.69433
R16923 GNDA.n2792 GNDA.n2471 1.69433
R16924 GNDA.n2792 GNDA.n2468 1.69433
R16925 GNDA.n2792 GNDA.n2465 1.69433
R16926 GNDA.n5802 GNDA.n4993 1.69433
R16927 GNDA.n5802 GNDA.n4990 1.69433
R16928 GNDA.n5802 GNDA.n4987 1.69433
R16929 GNDA.n5802 GNDA.n4984 1.69433
R16930 GNDA.n5802 GNDA.n4981 1.69433
R16931 GNDA.n5802 GNDA.n4978 1.69433
R16932 GNDA.n5802 GNDA.n4975 1.69433
R16933 GNDA.n4775 GNDA.n4470 1.69433
R16934 GNDA.n4775 GNDA.n4467 1.69433
R16935 GNDA.n4775 GNDA.n4464 1.69433
R16936 GNDA.n4775 GNDA.n4461 1.69433
R16937 GNDA.n4775 GNDA.n4458 1.69433
R16938 GNDA.n4775 GNDA.n4455 1.69433
R16939 GNDA.n4775 GNDA.n4452 1.69433
R16940 GNDA.n6286 GNDA.n383 1.69433
R16941 GNDA.n6286 GNDA.n380 1.69433
R16942 GNDA.n6286 GNDA.n377 1.69433
R16943 GNDA.n6286 GNDA.n374 1.69433
R16944 GNDA.n6286 GNDA.n371 1.69433
R16945 GNDA.n6286 GNDA.n368 1.69433
R16946 GNDA.n6286 GNDA.n365 1.69433
R16947 GNDA.n6615 GNDA.n6308 1.69433
R16948 GNDA.n6615 GNDA.n6305 1.69433
R16949 GNDA.n6615 GNDA.n6302 1.69433
R16950 GNDA.n6615 GNDA.n6299 1.69433
R16951 GNDA.n6615 GNDA.n6296 1.69433
R16952 GNDA.n6615 GNDA.n6293 1.69433
R16953 GNDA.n6615 GNDA.n6290 1.69433
R16954 GNDA.n3216 GNDA.n2388 1.69337
R16955 GNDA.n3216 GNDA.n2386 1.69337
R16956 GNDA.n3216 GNDA.n2383 1.69337
R16957 GNDA.n3216 GNDA.n2382 1.69337
R16958 GNDA.n3216 GNDA.n2379 1.69337
R16959 GNDA.n3216 GNDA.n2377 1.69337
R16960 GNDA.n3216 GNDA.n2374 1.69337
R16961 GNDA.n3216 GNDA.n2373 1.69337
R16962 GNDA.n3216 GNDA.n2370 1.69337
R16963 GNDA.n3216 GNDA.n2368 1.69337
R16964 GNDA.n3216 GNDA.n2365 1.69337
R16965 GNDA.n3216 GNDA.n2364 1.69337
R16966 GNDA.n3216 GNDA.n2361 1.69337
R16967 GNDA.n3216 GNDA.n2359 1.69337
R16968 GNDA.n3216 GNDA.n1893 1.69337
R16969 GNDA.n3217 GNDA.n3216 1.69337
R16970 GNDA.n3215 GNDA.n2413 1.6924
R16971 GNDA.n3215 GNDA.n2412 1.6924
R16972 GNDA.n3215 GNDA.n2410 1.6924
R16973 GNDA.n3215 GNDA.n2409 1.6924
R16974 GNDA.n3215 GNDA.n2407 1.6924
R16975 GNDA.n3215 GNDA.n2406 1.6924
R16976 GNDA.n3215 GNDA.n2404 1.6924
R16977 GNDA.n3215 GNDA.n2403 1.6924
R16978 GNDA.n3215 GNDA.n2401 1.6924
R16979 GNDA.n3215 GNDA.n2400 1.6924
R16980 GNDA.n3215 GNDA.n2398 1.6924
R16981 GNDA.n3215 GNDA.n2397 1.6924
R16982 GNDA.n3215 GNDA.n2395 1.6924
R16983 GNDA.n3215 GNDA.n2394 1.6924
R16984 GNDA.n3215 GNDA.n2392 1.6924
R16985 GNDA.n3215 GNDA.n2391 1.6924
R16986 GNDA.n3074 GNDA.n2437 1.6924
R16987 GNDA.n3074 GNDA.n2436 1.6924
R16988 GNDA.n3074 GNDA.n2434 1.6924
R16989 GNDA.n3074 GNDA.n2433 1.6924
R16990 GNDA.n3074 GNDA.n2431 1.6924
R16991 GNDA.n3074 GNDA.n2430 1.6924
R16992 GNDA.n3074 GNDA.n2428 1.6924
R16993 GNDA.n3074 GNDA.n2427 1.6924
R16994 GNDA.n3074 GNDA.n2425 1.6924
R16995 GNDA.n3074 GNDA.n2424 1.6924
R16996 GNDA.n3074 GNDA.n2422 1.6924
R16997 GNDA.n3074 GNDA.n2421 1.6924
R16998 GNDA.n3074 GNDA.n2419 1.6924
R16999 GNDA.n3074 GNDA.n2418 1.6924
R17000 GNDA.n3074 GNDA.n2416 1.6924
R17001 GNDA.n3074 GNDA.n2415 1.6924
R17002 GNDA.n2933 GNDA.n2461 1.6924
R17003 GNDA.n2933 GNDA.n2460 1.6924
R17004 GNDA.n2933 GNDA.n2458 1.6924
R17005 GNDA.n2933 GNDA.n2457 1.6924
R17006 GNDA.n2933 GNDA.n2455 1.6924
R17007 GNDA.n2933 GNDA.n2454 1.6924
R17008 GNDA.n2933 GNDA.n2452 1.6924
R17009 GNDA.n2933 GNDA.n2451 1.6924
R17010 GNDA.n2933 GNDA.n2449 1.6924
R17011 GNDA.n2933 GNDA.n2448 1.6924
R17012 GNDA.n2933 GNDA.n2446 1.6924
R17013 GNDA.n2933 GNDA.n2445 1.6924
R17014 GNDA.n2933 GNDA.n2443 1.6924
R17015 GNDA.n2933 GNDA.n2442 1.6924
R17016 GNDA.n2933 GNDA.n2440 1.6924
R17017 GNDA.n2933 GNDA.n2439 1.6924
R17018 GNDA.n2650 GNDA.n2509 1.6924
R17019 GNDA.n2650 GNDA.n2508 1.6924
R17020 GNDA.n2650 GNDA.n2506 1.6924
R17021 GNDA.n2650 GNDA.n2505 1.6924
R17022 GNDA.n2650 GNDA.n2503 1.6924
R17023 GNDA.n2650 GNDA.n2502 1.6924
R17024 GNDA.n2650 GNDA.n2500 1.6924
R17025 GNDA.n2650 GNDA.n2499 1.6924
R17026 GNDA.n2650 GNDA.n2497 1.6924
R17027 GNDA.n2650 GNDA.n2496 1.6924
R17028 GNDA.n2650 GNDA.n2494 1.6924
R17029 GNDA.n2650 GNDA.n2493 1.6924
R17030 GNDA.n2650 GNDA.n2491 1.6924
R17031 GNDA.n2650 GNDA.n2490 1.6924
R17032 GNDA.n2650 GNDA.n2488 1.6924
R17033 GNDA.n2650 GNDA.n2487 1.6924
R17034 GNDA.n3585 GNDA.n1862 1.6924
R17035 GNDA.n3585 GNDA.n1861 1.6924
R17036 GNDA.n3585 GNDA.n1859 1.6924
R17037 GNDA.n3585 GNDA.n1858 1.6924
R17038 GNDA.n3585 GNDA.n1856 1.6924
R17039 GNDA.n3585 GNDA.n1855 1.6924
R17040 GNDA.n3585 GNDA.n1853 1.6924
R17041 GNDA.n3585 GNDA.n1852 1.6924
R17042 GNDA.n3585 GNDA.n1850 1.6924
R17043 GNDA.n3585 GNDA.n1849 1.6924
R17044 GNDA.n3585 GNDA.n1847 1.6924
R17045 GNDA.n3585 GNDA.n1846 1.6924
R17046 GNDA.n3585 GNDA.n1844 1.6924
R17047 GNDA.n3585 GNDA.n1843 1.6924
R17048 GNDA.n3585 GNDA.n1841 1.6924
R17049 GNDA.n3585 GNDA.n1840 1.6924
R17050 GNDA.n4077 GNDA.n3774 1.6924
R17051 GNDA.n4077 GNDA.n3773 1.6924
R17052 GNDA.n4077 GNDA.n3771 1.6924
R17053 GNDA.n4077 GNDA.n3770 1.6924
R17054 GNDA.n4077 GNDA.n3768 1.6924
R17055 GNDA.n4077 GNDA.n3767 1.6924
R17056 GNDA.n4077 GNDA.n3765 1.6924
R17057 GNDA.n4077 GNDA.n3764 1.6924
R17058 GNDA.n4077 GNDA.n3762 1.6924
R17059 GNDA.n4077 GNDA.n3761 1.6924
R17060 GNDA.n4077 GNDA.n3759 1.6924
R17061 GNDA.n4077 GNDA.n3758 1.6924
R17062 GNDA.n4077 GNDA.n3756 1.6924
R17063 GNDA.n4077 GNDA.n3755 1.6924
R17064 GNDA.n4077 GNDA.n3753 1.6924
R17065 GNDA.n4077 GNDA.n3752 1.6924
R17066 GNDA.n3940 GNDA.n3798 1.6924
R17067 GNDA.n3940 GNDA.n3797 1.6924
R17068 GNDA.n3940 GNDA.n3795 1.6924
R17069 GNDA.n3940 GNDA.n3794 1.6924
R17070 GNDA.n3940 GNDA.n3792 1.6924
R17071 GNDA.n3940 GNDA.n3791 1.6924
R17072 GNDA.n3940 GNDA.n3789 1.6924
R17073 GNDA.n3940 GNDA.n3788 1.6924
R17074 GNDA.n3940 GNDA.n3786 1.6924
R17075 GNDA.n3940 GNDA.n3785 1.6924
R17076 GNDA.n3940 GNDA.n3783 1.6924
R17077 GNDA.n3940 GNDA.n3782 1.6924
R17078 GNDA.n3940 GNDA.n3780 1.6924
R17079 GNDA.n3940 GNDA.n3779 1.6924
R17080 GNDA.n3940 GNDA.n3777 1.6924
R17081 GNDA.n3940 GNDA.n3776 1.6924
R17082 GNDA.n1743 GNDA.n1599 1.6924
R17083 GNDA.n1746 GNDA.n1599 1.6924
R17084 GNDA.n1752 GNDA.n1599 1.6924
R17085 GNDA.n1755 GNDA.n1599 1.6924
R17086 GNDA.n1761 GNDA.n1599 1.6924
R17087 GNDA.n1764 GNDA.n1599 1.6924
R17088 GNDA.n1770 GNDA.n1599 1.6924
R17089 GNDA.n1773 GNDA.n1599 1.6924
R17090 GNDA.n1779 GNDA.n1599 1.6924
R17091 GNDA.n1782 GNDA.n1599 1.6924
R17092 GNDA.n1788 GNDA.n1599 1.6924
R17093 GNDA.n1791 GNDA.n1599 1.6924
R17094 GNDA.n1797 GNDA.n1599 1.6924
R17095 GNDA.n1800 GNDA.n1599 1.6924
R17096 GNDA.n1806 GNDA.n1599 1.6924
R17097 GNDA.n1809 GNDA.n1599 1.6924
R17098 GNDA.n4283 GNDA.n1623 1.6924
R17099 GNDA.n4283 GNDA.n1622 1.6924
R17100 GNDA.n4283 GNDA.n1620 1.6924
R17101 GNDA.n4283 GNDA.n1619 1.6924
R17102 GNDA.n4283 GNDA.n1617 1.6924
R17103 GNDA.n4283 GNDA.n1616 1.6924
R17104 GNDA.n4283 GNDA.n1614 1.6924
R17105 GNDA.n4283 GNDA.n1613 1.6924
R17106 GNDA.n4283 GNDA.n1611 1.6924
R17107 GNDA.n4283 GNDA.n1610 1.6924
R17108 GNDA.n4283 GNDA.n1608 1.6924
R17109 GNDA.n4283 GNDA.n1607 1.6924
R17110 GNDA.n4283 GNDA.n1605 1.6924
R17111 GNDA.n4283 GNDA.n1604 1.6924
R17112 GNDA.n4283 GNDA.n1602 1.6924
R17113 GNDA.n4283 GNDA.n1601 1.6924
R17114 GNDA.n4449 GNDA.n4307 1.6924
R17115 GNDA.n4449 GNDA.n4306 1.6924
R17116 GNDA.n4449 GNDA.n4304 1.6924
R17117 GNDA.n4449 GNDA.n4303 1.6924
R17118 GNDA.n4449 GNDA.n4301 1.6924
R17119 GNDA.n4449 GNDA.n4300 1.6924
R17120 GNDA.n4449 GNDA.n4298 1.6924
R17121 GNDA.n4449 GNDA.n4297 1.6924
R17122 GNDA.n4449 GNDA.n4295 1.6924
R17123 GNDA.n4449 GNDA.n4294 1.6924
R17124 GNDA.n4449 GNDA.n4292 1.6924
R17125 GNDA.n4449 GNDA.n4291 1.6924
R17126 GNDA.n4449 GNDA.n4289 1.6924
R17127 GNDA.n4449 GNDA.n4288 1.6924
R17128 GNDA.n4449 GNDA.n4286 1.6924
R17129 GNDA.n4449 GNDA.n4285 1.6924
R17130 GNDA.n4638 GNDA.n4496 1.6924
R17131 GNDA.n4638 GNDA.n4495 1.6924
R17132 GNDA.n4638 GNDA.n4493 1.6924
R17133 GNDA.n4638 GNDA.n4492 1.6924
R17134 GNDA.n4638 GNDA.n4490 1.6924
R17135 GNDA.n4638 GNDA.n4489 1.6924
R17136 GNDA.n4638 GNDA.n4487 1.6924
R17137 GNDA.n4638 GNDA.n4486 1.6924
R17138 GNDA.n4638 GNDA.n4484 1.6924
R17139 GNDA.n4638 GNDA.n4483 1.6924
R17140 GNDA.n4638 GNDA.n4481 1.6924
R17141 GNDA.n4638 GNDA.n4480 1.6924
R17142 GNDA.n4638 GNDA.n4478 1.6924
R17143 GNDA.n4638 GNDA.n4477 1.6924
R17144 GNDA.n4638 GNDA.n4475 1.6924
R17145 GNDA.n4638 GNDA.n4474 1.6924
R17146 GNDA.n4924 GNDA.n1395 1.6924
R17147 GNDA.n4924 GNDA.n1394 1.6924
R17148 GNDA.n4924 GNDA.n1392 1.6924
R17149 GNDA.n4924 GNDA.n1391 1.6924
R17150 GNDA.n4924 GNDA.n1389 1.6924
R17151 GNDA.n4924 GNDA.n1388 1.6924
R17152 GNDA.n4924 GNDA.n1386 1.6924
R17153 GNDA.n4924 GNDA.n1385 1.6924
R17154 GNDA.n4924 GNDA.n1383 1.6924
R17155 GNDA.n4924 GNDA.n1382 1.6924
R17156 GNDA.n4924 GNDA.n1380 1.6924
R17157 GNDA.n4924 GNDA.n1379 1.6924
R17158 GNDA.n4924 GNDA.n1377 1.6924
R17159 GNDA.n4924 GNDA.n1376 1.6924
R17160 GNDA.n4924 GNDA.n1374 1.6924
R17161 GNDA.n4924 GNDA.n1373 1.6924
R17162 GNDA.n5943 GNDA.n4971 1.6924
R17163 GNDA.n5943 GNDA.n4970 1.6924
R17164 GNDA.n5943 GNDA.n4968 1.6924
R17165 GNDA.n5943 GNDA.n4967 1.6924
R17166 GNDA.n5943 GNDA.n4965 1.6924
R17167 GNDA.n5943 GNDA.n4964 1.6924
R17168 GNDA.n5943 GNDA.n4962 1.6924
R17169 GNDA.n5943 GNDA.n4961 1.6924
R17170 GNDA.n5943 GNDA.n4959 1.6924
R17171 GNDA.n5943 GNDA.n4958 1.6924
R17172 GNDA.n5943 GNDA.n4956 1.6924
R17173 GNDA.n5943 GNDA.n4955 1.6924
R17174 GNDA.n5943 GNDA.n4953 1.6924
R17175 GNDA.n5943 GNDA.n4952 1.6924
R17176 GNDA.n5943 GNDA.n4950 1.6924
R17177 GNDA.n5943 GNDA.n4949 1.6924
R17178 GNDA.n5661 GNDA.n5019 1.6924
R17179 GNDA.n5661 GNDA.n5018 1.6924
R17180 GNDA.n5661 GNDA.n5016 1.6924
R17181 GNDA.n5661 GNDA.n5015 1.6924
R17182 GNDA.n5661 GNDA.n5013 1.6924
R17183 GNDA.n5661 GNDA.n5012 1.6924
R17184 GNDA.n5661 GNDA.n5010 1.6924
R17185 GNDA.n5661 GNDA.n5009 1.6924
R17186 GNDA.n5661 GNDA.n5007 1.6924
R17187 GNDA.n5661 GNDA.n5006 1.6924
R17188 GNDA.n5661 GNDA.n5004 1.6924
R17189 GNDA.n5661 GNDA.n5003 1.6924
R17190 GNDA.n5661 GNDA.n5001 1.6924
R17191 GNDA.n5661 GNDA.n5000 1.6924
R17192 GNDA.n5661 GNDA.n4998 1.6924
R17193 GNDA.n5661 GNDA.n4997 1.6924
R17194 GNDA.n5519 GNDA.n5043 1.6924
R17195 GNDA.n5519 GNDA.n5042 1.6924
R17196 GNDA.n5519 GNDA.n5040 1.6924
R17197 GNDA.n5519 GNDA.n5039 1.6924
R17198 GNDA.n5519 GNDA.n5037 1.6924
R17199 GNDA.n5519 GNDA.n5036 1.6924
R17200 GNDA.n5519 GNDA.n5034 1.6924
R17201 GNDA.n5519 GNDA.n5033 1.6924
R17202 GNDA.n5519 GNDA.n5031 1.6924
R17203 GNDA.n5519 GNDA.n5030 1.6924
R17204 GNDA.n5519 GNDA.n5028 1.6924
R17205 GNDA.n5519 GNDA.n5027 1.6924
R17206 GNDA.n5519 GNDA.n5025 1.6924
R17207 GNDA.n5519 GNDA.n5024 1.6924
R17208 GNDA.n5519 GNDA.n5022 1.6924
R17209 GNDA.n5519 GNDA.n5021 1.6924
R17210 GNDA.n5329 GNDA.n5044 1.6924
R17211 GNDA.n5332 GNDA.n5044 1.6924
R17212 GNDA.n5338 GNDA.n5044 1.6924
R17213 GNDA.n5341 GNDA.n5044 1.6924
R17214 GNDA.n5347 GNDA.n5044 1.6924
R17215 GNDA.n5350 GNDA.n5044 1.6924
R17216 GNDA.n5356 GNDA.n5044 1.6924
R17217 GNDA.n5359 GNDA.n5044 1.6924
R17218 GNDA.n5365 GNDA.n5044 1.6924
R17219 GNDA.n5368 GNDA.n5044 1.6924
R17220 GNDA.n5374 GNDA.n5044 1.6924
R17221 GNDA.n5377 GNDA.n5044 1.6924
R17222 GNDA.n5383 GNDA.n5044 1.6924
R17223 GNDA.n5386 GNDA.n5044 1.6924
R17224 GNDA.n5392 GNDA.n5044 1.6924
R17225 GNDA.n5395 GNDA.n5044 1.6924
R17226 GNDA.n5231 GNDA.n5094 1.6924
R17227 GNDA.n5231 GNDA.n5093 1.6924
R17228 GNDA.n5231 GNDA.n5091 1.6924
R17229 GNDA.n5231 GNDA.n5090 1.6924
R17230 GNDA.n5231 GNDA.n5088 1.6924
R17231 GNDA.n5231 GNDA.n5087 1.6924
R17232 GNDA.n5231 GNDA.n5085 1.6924
R17233 GNDA.n5231 GNDA.n5084 1.6924
R17234 GNDA.n5231 GNDA.n5082 1.6924
R17235 GNDA.n5231 GNDA.n5081 1.6924
R17236 GNDA.n5231 GNDA.n5079 1.6924
R17237 GNDA.n5231 GNDA.n5078 1.6924
R17238 GNDA.n5231 GNDA.n5076 1.6924
R17239 GNDA.n5231 GNDA.n5075 1.6924
R17240 GNDA.n5231 GNDA.n5073 1.6924
R17241 GNDA.n5231 GNDA.n5072 1.6924
R17242 GNDA.n3389 GNDA.n1838 1.6924
R17243 GNDA.n3392 GNDA.n1838 1.6924
R17244 GNDA.n3398 GNDA.n1838 1.6924
R17245 GNDA.n3401 GNDA.n1838 1.6924
R17246 GNDA.n3407 GNDA.n1838 1.6924
R17247 GNDA.n3410 GNDA.n1838 1.6924
R17248 GNDA.n3416 GNDA.n1838 1.6924
R17249 GNDA.n3419 GNDA.n1838 1.6924
R17250 GNDA.n3425 GNDA.n1838 1.6924
R17251 GNDA.n3428 GNDA.n1838 1.6924
R17252 GNDA.n3434 GNDA.n1838 1.6924
R17253 GNDA.n3437 GNDA.n1838 1.6924
R17254 GNDA.n3443 GNDA.n1838 1.6924
R17255 GNDA.n3446 GNDA.n1838 1.6924
R17256 GNDA.n3452 GNDA.n1838 1.6924
R17257 GNDA.n3455 GNDA.n1838 1.6924
R17258 GNDA.n3751 GNDA.n3609 1.6924
R17259 GNDA.n3751 GNDA.n3608 1.6924
R17260 GNDA.n3751 GNDA.n3606 1.6924
R17261 GNDA.n3751 GNDA.n3605 1.6924
R17262 GNDA.n3751 GNDA.n3603 1.6924
R17263 GNDA.n3751 GNDA.n3602 1.6924
R17264 GNDA.n3751 GNDA.n3600 1.6924
R17265 GNDA.n3751 GNDA.n3599 1.6924
R17266 GNDA.n3751 GNDA.n3597 1.6924
R17267 GNDA.n3751 GNDA.n3596 1.6924
R17268 GNDA.n3751 GNDA.n3594 1.6924
R17269 GNDA.n3751 GNDA.n3593 1.6924
R17270 GNDA.n3751 GNDA.n3591 1.6924
R17271 GNDA.n3751 GNDA.n3590 1.6924
R17272 GNDA.n3751 GNDA.n3588 1.6924
R17273 GNDA.n3751 GNDA.n3587 1.6924
R17274 GNDA.n1517 GNDA.n1371 1.6924
R17275 GNDA.n1520 GNDA.n1371 1.6924
R17276 GNDA.n1526 GNDA.n1371 1.6924
R17277 GNDA.n1529 GNDA.n1371 1.6924
R17278 GNDA.n1535 GNDA.n1371 1.6924
R17279 GNDA.n1538 GNDA.n1371 1.6924
R17280 GNDA.n1544 GNDA.n1371 1.6924
R17281 GNDA.n1547 GNDA.n1371 1.6924
R17282 GNDA.n1553 GNDA.n1371 1.6924
R17283 GNDA.n1556 GNDA.n1371 1.6924
R17284 GNDA.n1562 GNDA.n1371 1.6924
R17285 GNDA.n1565 GNDA.n1371 1.6924
R17286 GNDA.n1571 GNDA.n1371 1.6924
R17287 GNDA.n1574 GNDA.n1371 1.6924
R17288 GNDA.n1580 GNDA.n1371 1.6924
R17289 GNDA.n1583 GNDA.n1371 1.6924
R17290 GNDA.n6080 GNDA.n4947 1.6924
R17291 GNDA.n6080 GNDA.n4946 1.6924
R17292 GNDA.n6080 GNDA.n4944 1.6924
R17293 GNDA.n6080 GNDA.n4943 1.6924
R17294 GNDA.n6080 GNDA.n4941 1.6924
R17295 GNDA.n6080 GNDA.n4940 1.6924
R17296 GNDA.n6080 GNDA.n4938 1.6924
R17297 GNDA.n6080 GNDA.n4937 1.6924
R17298 GNDA.n6080 GNDA.n4935 1.6924
R17299 GNDA.n6080 GNDA.n4934 1.6924
R17300 GNDA.n6080 GNDA.n4932 1.6924
R17301 GNDA.n6080 GNDA.n4931 1.6924
R17302 GNDA.n6080 GNDA.n4929 1.6924
R17303 GNDA.n6080 GNDA.n4928 1.6924
R17304 GNDA.n6080 GNDA.n4926 1.6924
R17305 GNDA.n6080 GNDA.n4925 1.6924
R17306 GNDA.n2792 GNDA.n2485 1.6924
R17307 GNDA.n2792 GNDA.n2484 1.6924
R17308 GNDA.n2792 GNDA.n2482 1.6924
R17309 GNDA.n2792 GNDA.n2481 1.6924
R17310 GNDA.n2792 GNDA.n2479 1.6924
R17311 GNDA.n2792 GNDA.n2478 1.6924
R17312 GNDA.n2792 GNDA.n2476 1.6924
R17313 GNDA.n2792 GNDA.n2475 1.6924
R17314 GNDA.n2792 GNDA.n2473 1.6924
R17315 GNDA.n2792 GNDA.n2472 1.6924
R17316 GNDA.n2792 GNDA.n2470 1.6924
R17317 GNDA.n2792 GNDA.n2469 1.6924
R17318 GNDA.n2792 GNDA.n2467 1.6924
R17319 GNDA.n2792 GNDA.n2466 1.6924
R17320 GNDA.n2792 GNDA.n2464 1.6924
R17321 GNDA.n2792 GNDA.n2463 1.6924
R17322 GNDA.n5802 GNDA.n4995 1.6924
R17323 GNDA.n5802 GNDA.n4994 1.6924
R17324 GNDA.n5802 GNDA.n4992 1.6924
R17325 GNDA.n5802 GNDA.n4991 1.6924
R17326 GNDA.n5802 GNDA.n4989 1.6924
R17327 GNDA.n5802 GNDA.n4988 1.6924
R17328 GNDA.n5802 GNDA.n4986 1.6924
R17329 GNDA.n5802 GNDA.n4985 1.6924
R17330 GNDA.n5802 GNDA.n4983 1.6924
R17331 GNDA.n5802 GNDA.n4982 1.6924
R17332 GNDA.n5802 GNDA.n4980 1.6924
R17333 GNDA.n5802 GNDA.n4979 1.6924
R17334 GNDA.n5802 GNDA.n4977 1.6924
R17335 GNDA.n5802 GNDA.n4976 1.6924
R17336 GNDA.n5802 GNDA.n4974 1.6924
R17337 GNDA.n5802 GNDA.n4973 1.6924
R17338 GNDA.n4775 GNDA.n4472 1.6924
R17339 GNDA.n4775 GNDA.n4471 1.6924
R17340 GNDA.n4775 GNDA.n4469 1.6924
R17341 GNDA.n4775 GNDA.n4468 1.6924
R17342 GNDA.n4775 GNDA.n4466 1.6924
R17343 GNDA.n4775 GNDA.n4465 1.6924
R17344 GNDA.n4775 GNDA.n4463 1.6924
R17345 GNDA.n4775 GNDA.n4462 1.6924
R17346 GNDA.n4775 GNDA.n4460 1.6924
R17347 GNDA.n4775 GNDA.n4459 1.6924
R17348 GNDA.n4775 GNDA.n4457 1.6924
R17349 GNDA.n4775 GNDA.n4456 1.6924
R17350 GNDA.n4775 GNDA.n4454 1.6924
R17351 GNDA.n4775 GNDA.n4453 1.6924
R17352 GNDA.n4775 GNDA.n4451 1.6924
R17353 GNDA.n4775 GNDA.n4450 1.6924
R17354 GNDA.n6286 GNDA.n385 1.6924
R17355 GNDA.n6286 GNDA.n384 1.6924
R17356 GNDA.n6286 GNDA.n382 1.6924
R17357 GNDA.n6286 GNDA.n381 1.6924
R17358 GNDA.n6286 GNDA.n379 1.6924
R17359 GNDA.n6286 GNDA.n378 1.6924
R17360 GNDA.n6286 GNDA.n376 1.6924
R17361 GNDA.n6286 GNDA.n375 1.6924
R17362 GNDA.n6286 GNDA.n373 1.6924
R17363 GNDA.n6286 GNDA.n372 1.6924
R17364 GNDA.n6286 GNDA.n370 1.6924
R17365 GNDA.n6286 GNDA.n369 1.6924
R17366 GNDA.n6286 GNDA.n367 1.6924
R17367 GNDA.n6286 GNDA.n366 1.6924
R17368 GNDA.n6286 GNDA.n364 1.6924
R17369 GNDA.n6286 GNDA.n363 1.6924
R17370 GNDA.n6615 GNDA.n6445 1.6924
R17371 GNDA.n6615 GNDA.n6309 1.6924
R17372 GNDA.n6615 GNDA.n6307 1.6924
R17373 GNDA.n6615 GNDA.n6306 1.6924
R17374 GNDA.n6615 GNDA.n6304 1.6924
R17375 GNDA.n6615 GNDA.n6303 1.6924
R17376 GNDA.n6615 GNDA.n6301 1.6924
R17377 GNDA.n6615 GNDA.n6300 1.6924
R17378 GNDA.n6615 GNDA.n6298 1.6924
R17379 GNDA.n6615 GNDA.n6297 1.6924
R17380 GNDA.n6615 GNDA.n6295 1.6924
R17381 GNDA.n6615 GNDA.n6294 1.6924
R17382 GNDA.n6615 GNDA.n6292 1.6924
R17383 GNDA.n6615 GNDA.n6291 1.6924
R17384 GNDA.n6615 GNDA.n6289 1.6924
R17385 GNDA.n6615 GNDA.n6288 1.6924
R17386 GNDA.n3216 GNDA.n2389 1.6924
R17387 GNDA.n3216 GNDA.n2385 1.6924
R17388 GNDA.n3216 GNDA.n2380 1.6924
R17389 GNDA.n3216 GNDA.n2376 1.6924
R17390 GNDA.n3216 GNDA.n2371 1.6924
R17391 GNDA.n3216 GNDA.n2367 1.6924
R17392 GNDA.n3216 GNDA.n2362 1.6924
R17393 GNDA.n3216 GNDA.n2358 1.6924
R17394 GNDA.t743 GNDA.t34 1.57352
R17395 GNDA.n1339 GNDA.n1338 1.47392
R17396 GNDA.n824 GNDA.n823 1.47392
R17397 GNDA.n6925 GNDA.n229 1.47392
R17398 GNDA.n6902 GNDA.n6899 1.47392
R17399 GNDA.n1058 GNDA.n1057 1.47392
R17400 GNDA.n7148 GNDA.n87 1.47392
R17401 GNDA.n6088 GNDA.n6087 1.44719
R17402 GNDA.n4780 GNDA.n4779 1.44719
R17403 GNDA.n3292 GNDA.n1888 1.44719
R17404 GNDA.t469 GNDA.n105 1.37214
R17405 GNDA.n3290 GNDA.n3289 1.08947
R17406 GNDA.n3291 GNDA.n3290 1.08947
R17407 GNDA.n3292 GNDA.n3291 1.08947
R17408 GNDA.n4081 GNDA.n1814 1.08947
R17409 GNDA.n4165 GNDA.n4164 1.08947
R17410 GNDA.n6087 GNDA.n6086 1.08947
R17411 GNDA.n5401 GNDA.n1362 1.08947
R17412 GNDA.n5401 GNDA.n5400 1.08947
R17413 GNDA.n6087 GNDA.n1362 1.08947
R17414 GNDA.n4780 GNDA.n1592 1.08947
R17415 GNDA.n3293 GNDA.n3292 1.08947
R17416 GNDA.n3294 GNDA.n3293 1.03004
R17417 GNDA.n1592 GNDA.n1422 1.03004
R17418 GNDA.n4082 GNDA.n4081 1.02968
R17419 GNDA.n6086 GNDA.n6085 1.02968
R17420 GNDA.n4779 GNDA.n4778 0.948417
R17421 GNDA.n6088 GNDA.n1361 0.948417
R17422 GNDA.n2697 GNDA.n1888 0.948417
R17423 GNDA.n6084 GNDA.n6083 0.927583
R17424 GNDA.n1588 GNDA.n1587 0.927583
R17425 GNDA.n3634 GNDA.n1832 0.927583
R17426 GNDA.n3460 GNDA.n3459 0.927583
R17427 GNDA.n1329 GNDA.n1241 0.8197
R17428 GNDA.n1328 GNDA.n1242 0.8197
R17429 GNDA.n1324 GNDA.n1323 0.8197
R17430 GNDA.n1318 GNDA.n1315 0.8197
R17431 GNDA.n6250 GNDA.n6249 0.8197
R17432 GNDA.n549 GNDA.n548 0.8197
R17433 GNDA.n6258 GNDA.n545 0.8197
R17434 GNDA.n6257 GNDA.n546 0.8197
R17435 GNDA.n601 GNDA.n596 0.8197
R17436 GNDA.n6188 GNDA.n602 0.8197
R17437 GNDA.n6187 GNDA.n603 0.8197
R17438 GNDA.n6110 GNDA.n6106 0.8197
R17439 GNDA.n6119 GNDA.n6117 0.8197
R17440 GNDA.n6118 GNDA.n623 0.8197
R17441 GNDA.n6127 GNDA.n6126 0.8197
R17442 GNDA.n621 GNDA.n620 0.8197
R17443 GNDA.n7106 GNDA.n166 0.8197
R17444 GNDA.n7105 GNDA.n168 0.8197
R17445 GNDA.n219 GNDA.n201 0.8197
R17446 GNDA.n218 GNDA.n216 0.8197
R17447 GNDA.n212 GNDA.n211 0.8197
R17448 GNDA.n208 GNDA.n204 0.8197
R17449 GNDA.n207 GNDA.n188 0.8197
R17450 GNDA.n7047 GNDA.n7046 0.8197
R17451 GNDA.n808 GNDA.n807 0.8197
R17452 GNDA.n804 GNDA.n803 0.8197
R17453 GNDA.n800 GNDA.n784 0.8197
R17454 GNDA.n799 GNDA.n796 0.8197
R17455 GNDA.n792 GNDA.n789 0.8197
R17456 GNDA.n786 GNDA.n708 0.8197
R17457 GNDA.n814 GNDA.n813 0.8197
R17458 GNDA.n817 GNDA.n707 0.8197
R17459 GNDA.n7037 GNDA.n6928 0.8197
R17460 GNDA.n7034 GNDA.n7033 0.8197
R17461 GNDA.n7030 GNDA.n6931 0.8197
R17462 GNDA.n7029 GNDA.n6932 0.8197
R17463 GNDA.n6964 GNDA.n6961 0.8197
R17464 GNDA.n6965 GNDA.n6955 0.8197
R17465 GNDA.n6969 GNDA.n6968 0.8197
R17466 GNDA.n6973 GNDA.n6972 0.8197
R17467 GNDA.n7316 GNDA.n59 0.8197
R17468 GNDA.n7313 GNDA.n7312 0.8197
R17469 GNDA.n7309 GNDA.n62 0.8197
R17470 GNDA.n7308 GNDA.n63 0.8197
R17471 GNDA.n7243 GNDA.n7240 0.8197
R17472 GNDA.n7244 GNDA.n7234 0.8197
R17473 GNDA.n7248 GNDA.n7247 0.8197
R17474 GNDA.n7252 GNDA.n7251 0.8197
R17475 GNDA.n6891 GNDA.n6783 0.8197
R17476 GNDA.n6890 GNDA.n6784 0.8197
R17477 GNDA.n6810 GNDA.n6807 0.8197
R17478 GNDA.n6813 GNDA.n6812 0.8197
R17479 GNDA.n6823 GNDA.n6820 0.8197
R17480 GNDA.n6824 GNDA.n6806 0.8197
R17481 GNDA.n6828 GNDA.n6827 0.8197
R17482 GNDA.n6832 GNDA.n6831 0.8197
R17483 GNDA.n1041 GNDA.n1040 0.8197
R17484 GNDA.n1047 GNDA.n929 0.8197
R17485 GNDA.n1046 GNDA.n930 0.8197
R17486 GNDA.n966 GNDA.n965 0.8197
R17487 GNDA.n972 GNDA.n964 0.8197
R17488 GNDA.n980 GNDA.n946 0.8197
R17489 GNDA.n982 GNDA.n981 0.8197
R17490 GNDA.n6200 GNDA.n593 0.8197
R17491 GNDA.n7326 GNDA.n7325 0.8197
R17492 GNDA.n32 GNDA.n23 0.8197
R17493 GNDA.n39 GNDA.n33 0.8197
R17494 GNDA.n38 GNDA.n35 0.8197
R17495 GNDA.n7331 GNDA.n1 0.8197
R17496 GNDA.n7163 GNDA.n7160 0.8197
R17497 GNDA.n7166 GNDA.n7165 0.8197
R17498 GNDA.n7170 GNDA.n7169 0.8197
R17499 GNDA.n4164 GNDA.n4163 0.794805
R17500 GNDA.n4781 GNDA.n4780 0.77918
R17501 GNDA.n1648 GNDA.n1591 0.71668
R17502 GNDA.n3466 GNDA.n3464 0.65675
R17503 GNDA.n4083 GNDA.n1834 0.65675
R17504 GNDA.n4805 GNDA.n4803 0.65675
R17505 GNDA.n1421 GNDA.n1364 0.65675
R17506 GNDA.n6615 GNDA.n6614 0.626041
R17507 GNDA.n1317 GNDA 0.5637
R17508 GNDA.n6112 GNDA 0.5637
R17509 GNDA.n215 GNDA 0.5637
R17510 GNDA GNDA.n785 0.5637
R17511 GNDA GNDA.n6956 0.5637
R17512 GNDA GNDA.n7235 0.5637
R17513 GNDA.n6817 GNDA 0.5637
R17514 GNDA.n967 GNDA 0.5637
R17515 GNDA.n34 GNDA 0.5637
R17516 GNDA.n4161 GNDA.n4159 0.563
R17517 GNDA.n4159 GNDA.n4157 0.563
R17518 GNDA.n4157 GNDA.n4155 0.563
R17519 GNDA.n4155 GNDA.n4153 0.563
R17520 GNDA.n4153 GNDA.n4151 0.563
R17521 GNDA.n4151 GNDA.n4149 0.563
R17522 GNDA.n4149 GNDA.n4147 0.563
R17523 GNDA.n4147 GNDA.n4145 0.563
R17524 GNDA.n4145 GNDA.n4143 0.563
R17525 GNDA.n4143 GNDA.n4141 0.563
R17526 GNDA.n1354 GNDA.n1352 0.563
R17527 GNDA.n1356 GNDA.n1354 0.563
R17528 GNDA.n1358 GNDA.n1356 0.563
R17529 GNDA.n1360 GNDA.n1358 0.563
R17530 GNDA.n1829 GNDA.n1827 0.563
R17531 GNDA.n1827 GNDA.n1825 0.563
R17532 GNDA.n1825 GNDA.n1823 0.563
R17533 GNDA.n1823 GNDA.n1821 0.563
R17534 GNDA.n1821 GNDA.n1819 0.563
R17535 GNDA.n4123 GNDA.n4121 0.563
R17536 GNDA.n4165 GNDA.n1648 0.373287
R17537 GNDA.n6447 GNDA.n6446 0.3295
R17538 GNDA.n6448 GNDA.n6447 0.3295
R17539 GNDA.n6452 GNDA.n6448 0.3295
R17540 GNDA.n6452 GNDA.n6451 0.3295
R17541 GNDA.n6451 GNDA.n6450 0.3295
R17542 GNDA.n6450 GNDA.n6449 0.3295
R17543 GNDA.n6454 GNDA.n6453 0.3295
R17544 GNDA.n6455 GNDA.n6454 0.3295
R17545 GNDA.n6459 GNDA.n6455 0.3295
R17546 GNDA.n6459 GNDA.n6458 0.3295
R17547 GNDA.n6458 GNDA.n6457 0.3295
R17548 GNDA.n6457 GNDA.n6456 0.3295
R17549 GNDA.n6461 GNDA.n6460 0.3295
R17550 GNDA.n6462 GNDA.n6461 0.3295
R17551 GNDA.n6466 GNDA.n6462 0.3295
R17552 GNDA.n6466 GNDA.n6465 0.3295
R17553 GNDA.n6465 GNDA.n6464 0.3295
R17554 GNDA.n6464 GNDA.n6463 0.3295
R17555 GNDA.n6468 GNDA.n6467 0.3295
R17556 GNDA.n6469 GNDA.n6468 0.3295
R17557 GNDA.n6473 GNDA.n6469 0.3295
R17558 GNDA.n6473 GNDA.n6472 0.3295
R17559 GNDA.n6472 GNDA.n6471 0.3295
R17560 GNDA.n6471 GNDA.n6470 0.3295
R17561 GNDA.n6475 GNDA.n6474 0.3295
R17562 GNDA.n6476 GNDA.n6475 0.3295
R17563 GNDA.n6480 GNDA.n6476 0.3295
R17564 GNDA.n6480 GNDA.n6479 0.3295
R17565 GNDA.n6479 GNDA.n6478 0.3295
R17566 GNDA.n6478 GNDA.n6477 0.3295
R17567 GNDA.n6482 GNDA.n6481 0.3295
R17568 GNDA.n6483 GNDA.n6482 0.3295
R17569 GNDA.n6487 GNDA.n6483 0.3295
R17570 GNDA.n6487 GNDA.n6486 0.3295
R17571 GNDA.n6486 GNDA.n6485 0.3295
R17572 GNDA.n6485 GNDA.n6484 0.3295
R17573 GNDA.n6489 GNDA.n6488 0.3295
R17574 GNDA.n6490 GNDA.n6489 0.3295
R17575 GNDA.n6494 GNDA.n6490 0.3295
R17576 GNDA.n6494 GNDA.n6493 0.3295
R17577 GNDA.n6493 GNDA.n6492 0.3295
R17578 GNDA.n6492 GNDA.n6491 0.3295
R17579 GNDA.n6496 GNDA.n6495 0.3295
R17580 GNDA.n6497 GNDA.n6496 0.3295
R17581 GNDA.n6501 GNDA.n6497 0.3295
R17582 GNDA.n6501 GNDA.n6500 0.3295
R17583 GNDA.n6500 GNDA.n6499 0.3295
R17584 GNDA.n6499 GNDA.n6498 0.3295
R17585 GNDA.n6503 GNDA.n6502 0.3295
R17586 GNDA.n6504 GNDA.n6503 0.3295
R17587 GNDA.n6508 GNDA.n6504 0.3295
R17588 GNDA.n6508 GNDA.n6507 0.3295
R17589 GNDA.n6507 GNDA.n6506 0.3295
R17590 GNDA.n6506 GNDA.n6505 0.3295
R17591 GNDA.n6510 GNDA.n6509 0.3295
R17592 GNDA.n6511 GNDA.n6510 0.3295
R17593 GNDA.n6515 GNDA.n6511 0.3295
R17594 GNDA.n6515 GNDA.n6514 0.3295
R17595 GNDA.n6514 GNDA.n6513 0.3295
R17596 GNDA.n6513 GNDA.n6512 0.3295
R17597 GNDA.n6517 GNDA.n6516 0.3295
R17598 GNDA.n6518 GNDA.n6517 0.3295
R17599 GNDA.n6522 GNDA.n6518 0.3295
R17600 GNDA.n6522 GNDA.n6521 0.3295
R17601 GNDA.n6521 GNDA.n6520 0.3295
R17602 GNDA.n6520 GNDA.n6519 0.3295
R17603 GNDA.n6524 GNDA.n6523 0.3295
R17604 GNDA.n6525 GNDA.n6524 0.3295
R17605 GNDA.n6529 GNDA.n6525 0.3295
R17606 GNDA.n6529 GNDA.n6528 0.3295
R17607 GNDA.n6528 GNDA.n6527 0.3295
R17608 GNDA.n6527 GNDA.n6526 0.3295
R17609 GNDA.n6531 GNDA.n6530 0.3295
R17610 GNDA.n6532 GNDA.n6531 0.3295
R17611 GNDA.n6536 GNDA.n6532 0.3295
R17612 GNDA.n6536 GNDA.n6535 0.3295
R17613 GNDA.n6535 GNDA.n6534 0.3295
R17614 GNDA.n6534 GNDA.n6533 0.3295
R17615 GNDA.n6538 GNDA.n6537 0.3295
R17616 GNDA.n6539 GNDA.n6538 0.3295
R17617 GNDA.n6543 GNDA.n6539 0.3295
R17618 GNDA.n6543 GNDA.n6542 0.3295
R17619 GNDA.n6542 GNDA.n6541 0.3295
R17620 GNDA.n6541 GNDA.n6540 0.3295
R17621 GNDA.n6545 GNDA.n6544 0.3295
R17622 GNDA.n6546 GNDA.n6545 0.3295
R17623 GNDA.n6550 GNDA.n6546 0.3295
R17624 GNDA.n6550 GNDA.n6549 0.3295
R17625 GNDA.n6549 GNDA.n6548 0.3295
R17626 GNDA.n6548 GNDA.n6547 0.3295
R17627 GNDA.n6552 GNDA.n6551 0.3295
R17628 GNDA.n6553 GNDA.n6552 0.3295
R17629 GNDA.n6557 GNDA.n6553 0.3295
R17630 GNDA.n6557 GNDA.n6556 0.3295
R17631 GNDA.n6556 GNDA.n6555 0.3295
R17632 GNDA.n6555 GNDA.n6554 0.3295
R17633 GNDA.n6559 GNDA.n6558 0.3295
R17634 GNDA.n6560 GNDA.n6559 0.3295
R17635 GNDA.n6564 GNDA.n6560 0.3295
R17636 GNDA.n6564 GNDA.n6563 0.3295
R17637 GNDA.n6563 GNDA.n6562 0.3295
R17638 GNDA.n6562 GNDA.n6561 0.3295
R17639 GNDA.n6566 GNDA.n6565 0.3295
R17640 GNDA.n6567 GNDA.n6566 0.3295
R17641 GNDA.n6571 GNDA.n6567 0.3295
R17642 GNDA.n6571 GNDA.n6570 0.3295
R17643 GNDA.n6570 GNDA.n6569 0.3295
R17644 GNDA.n6569 GNDA.n6568 0.3295
R17645 GNDA.n6573 GNDA.n6572 0.3295
R17646 GNDA.n6574 GNDA.n6573 0.3295
R17647 GNDA.n6578 GNDA.n6574 0.3295
R17648 GNDA.n6578 GNDA.n6577 0.3295
R17649 GNDA.n6577 GNDA.n6576 0.3295
R17650 GNDA.n6576 GNDA.n6575 0.3295
R17651 GNDA.n6580 GNDA.n6579 0.3295
R17652 GNDA.n6581 GNDA.n6580 0.3295
R17653 GNDA.n6585 GNDA.n6581 0.3295
R17654 GNDA.n6585 GNDA.n6584 0.3295
R17655 GNDA.n6584 GNDA.n6583 0.3295
R17656 GNDA.n6583 GNDA.n6582 0.3295
R17657 GNDA.n6587 GNDA.n6586 0.3295
R17658 GNDA.n6588 GNDA.n6587 0.3295
R17659 GNDA.n6592 GNDA.n6588 0.3295
R17660 GNDA.n6592 GNDA.n6591 0.3295
R17661 GNDA.n6591 GNDA.n6590 0.3295
R17662 GNDA.n6590 GNDA.n6589 0.3295
R17663 GNDA.n6594 GNDA.n6593 0.3295
R17664 GNDA.n6595 GNDA.n6594 0.3295
R17665 GNDA.n6599 GNDA.n6595 0.3295
R17666 GNDA.n6599 GNDA.n6598 0.3295
R17667 GNDA.n6598 GNDA.n6597 0.3295
R17668 GNDA.n6597 GNDA.n6596 0.3295
R17669 GNDA.n6601 GNDA.n6600 0.3295
R17670 GNDA.n6602 GNDA.n6601 0.3295
R17671 GNDA.n6606 GNDA.n6602 0.3295
R17672 GNDA.n6606 GNDA.n6605 0.3295
R17673 GNDA.n6605 GNDA.n6604 0.3295
R17674 GNDA.n6604 GNDA.n6603 0.3295
R17675 GNDA.n6614 GNDA.n6613 0.3295
R17676 GNDA.n6613 GNDA.n6612 0.3295
R17677 GNDA.n6612 GNDA.n6611 0.3295
R17678 GNDA.n6611 GNDA.n6610 0.3295
R17679 GNDA.n6610 GNDA.n6609 0.3295
R17680 GNDA.n6609 GNDA.n6608 0.3295
R17681 GNDA.n6608 GNDA.n6607 0.3295
R17682 GNDA.n3467 GNDA.n1834 0.310787
R17683 GNDA.n4781 GNDA.n1591 0.310787
R17684 GNDA.n4806 GNDA.n1421 0.310787
R17685 GNDA.n3467 GNDA.n3466 0.31043
R17686 GNDA.n4806 GNDA.n4805 0.31043
R17687 GNDA.n4163 GNDA.n1814 0.295162
R17688 GNDA.n6459 GNDA.n6452 0.2825
R17689 GNDA.n6466 GNDA.n6459 0.2825
R17690 GNDA.n6473 GNDA.n6466 0.2825
R17691 GNDA.n6480 GNDA.n6473 0.2825
R17692 GNDA.n6487 GNDA.n6480 0.2825
R17693 GNDA.n6494 GNDA.n6487 0.2825
R17694 GNDA.n6501 GNDA.n6494 0.2825
R17695 GNDA.n6508 GNDA.n6501 0.2825
R17696 GNDA.n6515 GNDA.n6508 0.2825
R17697 GNDA.n6522 GNDA.n6515 0.2825
R17698 GNDA.n6529 GNDA.n6522 0.2825
R17699 GNDA.n6536 GNDA.n6529 0.2825
R17700 GNDA.n6543 GNDA.n6536 0.2825
R17701 GNDA.n6550 GNDA.n6543 0.2825
R17702 GNDA.n6557 GNDA.n6550 0.2825
R17703 GNDA.n6564 GNDA.n6557 0.2825
R17704 GNDA.n6571 GNDA.n6564 0.2825
R17705 GNDA.n6578 GNDA.n6571 0.2825
R17706 GNDA.n6585 GNDA.n6578 0.2825
R17707 GNDA.n6592 GNDA.n6585 0.2825
R17708 GNDA.n6599 GNDA.n6592 0.2825
R17709 GNDA.n6606 GNDA.n6599 0.2825
R17710 GNDA.n6610 GNDA.n6606 0.2825
R17711 GNDA.n6922 GNDA.n105 0.270774
R17712 GNDA GNDA.n1316 0.2565
R17713 GNDA GNDA.n6111 0.2565
R17714 GNDA.n203 GNDA 0.2565
R17715 GNDA.n793 GNDA 0.2565
R17716 GNDA.n6959 GNDA 0.2565
R17717 GNDA.n7238 GNDA 0.2565
R17718 GNDA GNDA.n6816 0.2565
R17719 GNDA.n973 GNDA 0.2565
R17720 GNDA GNDA.n0 0.2565
R17721 GNDA.n6277 GNDA.n6276 0.214042
R17722 GNDA.n4790 GNDA.n4788 0.208833
R17723 GNDA.n4134 GNDA.n4133 0.208833
R17724 GNDA.n3464 GNDA.n3294 0.186811
R17725 GNDA.n4083 GNDA.n4082 0.186811
R17726 GNDA.n4803 GNDA.n1422 0.186811
R17727 GNDA.n6085 GNDA.n1364 0.186811
R17728 GNDA.t404 GNDA.t570 0.1603
R17729 GNDA.t274 GNDA.t404 0.1603
R17730 GNDA.t342 GNDA.t274 0.1603
R17731 GNDA.t416 GNDA.t342 0.1603
R17732 GNDA.t285 GNDA.t416 0.1603
R17733 GNDA.t352 GNDA.t285 0.1603
R17734 GNDA.t223 GNDA.t352 0.1603
R17735 GNDA.t577 GNDA.t725 0.1603
R17736 GNDA.t412 GNDA.t577 0.1603
R17737 GNDA.t515 GNDA.t412 0.1603
R17738 GNDA.t588 GNDA.t515 0.1603
R17739 GNDA.t423 GNDA.t588 0.1603
R17740 GNDA.t525 GNDA.t423 0.1603
R17741 GNDA.t362 GNDA.t525 0.1603
R17742 GNDA.t208 GNDA.t296 0.1603
R17743 GNDA.t338 GNDA.t208 0.1603
R17744 GNDA.t505 GNDA.t338 0.1603
R17745 GNDA.t403 GNDA.t505 0.1603
R17746 GNDA.t568 GNDA.t403 0.1603
R17747 GNDA.t714 GNDA.t568 0.1603
R17748 GNDA.t632 GNDA.t714 0.1603
R17749 GNDA.t424 GNDA.t589 0.1603
R17750 GNDA.t294 GNDA.t424 0.1603
R17751 GNDA.t364 GNDA.t294 0.1603
R17752 GNDA.t436 GNDA.t364 0.1603
R17753 GNDA.t306 GNDA.t436 0.1603
R17754 GNDA.t376 GNDA.t306 0.1603
R17755 GNDA.t245 GNDA.t376 0.1603
R17756 GNDA.t619 GNDA.t702 0.1603
R17757 GNDA.t220 GNDA.t619 0.1603
R17758 GNDA.t350 GNDA.t220 0.1603
R17759 GNDA.t284 GNDA.t350 0.1603
R17760 GNDA.t413 GNDA.t284 0.1603
R17761 GNDA.t579 GNDA.t413 0.1603
R17762 GNDA.t496 GNDA.t579 0.1603
R17763 GNDA.t595 GNDA.t197 0.1603
R17764 GNDA.t433 GNDA.t595 0.1603
R17765 GNDA.t534 GNDA.t433 0.1603
R17766 GNDA.t607 GNDA.t534 0.1603
R17767 GNDA.t443 GNDA.t607 0.1603
R17768 GNDA.t545 GNDA.t443 0.1603
R17769 GNDA.t384 GNDA.t545 0.1603
R17770 GNDA.t231 GNDA.t456 0.1603
R17771 GNDA.t359 GNDA.t231 0.1603
R17772 GNDA.t522 GNDA.t359 0.1603
R17773 GNDA.t422 GNDA.t522 0.1603
R17774 GNDA.t585 GNDA.t422 0.1603
R17775 GNDA.t188 GNDA.t585 0.1603
R17776 GNDA.t652 GNDA.t188 0.1603
R17777 GNDA.t205 GNDA.t336 0.1603
R17778 GNDA.t602 GNDA.t205 0.1603
R17779 GNDA.t689 GNDA.t602 0.1603
R17780 GNDA.t218 GNDA.t689 0.1603
R17781 GNDA.t614 GNDA.t218 0.1603
R17782 GNDA.t700 GNDA.t614 0.1603
R17783 GNDA.t552 GNDA.t700 0.1603
R17784 GNDA.t370 GNDA.t477 0.1603
R17785 GNDA.t529 GNDA.t370 0.1603
R17786 GNDA.t677 GNDA.t529 0.1603
R17787 GNDA.t593 GNDA.t677 0.1603
R17788 GNDA.t193 GNDA.t593 0.1603
R17789 GNDA.t327 GNDA.t193 0.1603
R17790 GNDA.t259 GNDA.t327 0.1603
R17791 GNDA.t615 GNDA.t219 0.1603
R17792 GNDA.t476 GNDA.t615 0.1603
R17793 GNDA.t554 GNDA.t476 0.1603
R17794 GNDA.t631 GNDA.t554 0.1603
R17795 GNDA.t736 GNDA.t631 0.1603
R17796 GNDA.t565 GNDA.t736 0.1603
R17797 GNDA.t401 GNDA.t565 0.1603
R17798 GNDA.t250 GNDA.t320 0.1603
R17799 GNDA.t382 GNDA.t250 0.1603
R17800 GNDA.t543 GNDA.t382 0.1603
R17801 GNDA.t441 GNDA.t543 0.1603
R17802 GNDA.t604 GNDA.t441 0.1603
R17803 GNDA.t204 GNDA.t604 0.1603
R17804 GNDA.t667 GNDA.t204 0.1603
R17805 GNDA.t228 GNDA.t358 0.1603
R17806 GNDA.t628 GNDA.t228 0.1603
R17807 GNDA.t709 GNDA.t628 0.1603
R17808 GNDA.t242 GNDA.t709 0.1603
R17809 GNDA.t639 GNDA.t242 0.1603
R17810 GNDA.t721 GNDA.t639 0.1603
R17811 GNDA.t575 GNDA.t721 0.1603
R17812 GNDA.t387 GNDA.t492 0.1603
R17813 GNDA.t550 GNDA.t387 0.1603
R17814 GNDA.t698 GNDA.t550 0.1603
R17815 GNDA.t613 GNDA.t698 0.1603
R17816 GNDA.t215 GNDA.t613 0.1603
R17817 GNDA.t347 GNDA.t215 0.1603
R17818 GNDA.t279 GNDA.t347 0.1603
R17819 GNDA.t344 GNDA.t509 0.1603
R17820 GNDA.t211 GNDA.t344 0.1603
R17821 GNDA.t301 GNDA.t211 0.1603
R17822 GNDA.t354 GNDA.t301 0.1603
R17823 GNDA.t225 GNDA.t354 0.1603
R17824 GNDA.t453 GNDA.t225 0.1603
R17825 GNDA.t705 GNDA.t453 0.1603
R17826 GNDA.t538 GNDA.t626 0.1603
R17827 GNDA.t684 GNDA.t538 0.1603
R17828 GNDA.t288 GNDA.t684 0.1603
R17829 GNDA.t201 GNDA.t288 0.1603
R17830 GNDA.t332 GNDA.t201 0.1603
R17831 GNDA.t499 GNDA.t332 0.1603
R17832 GNDA.t398 GNDA.t499 0.1603
R17833 GNDA.t226 GNDA.t357 0.1603
R17834 GNDA.t624 GNDA.t226 0.1603
R17835 GNDA.t708 GNDA.t624 0.1603
R17836 GNDA.t237 GNDA.t708 0.1603
R17837 GNDA.t638 GNDA.t237 0.1603
R17838 GNDA.t717 GNDA.t638 0.1603
R17839 GNDA.t571 GNDA.t717 0.1603
R17840 GNDA.t468 GNDA.t489 0.1603
R17841 GNDA.t549 GNDA.t468 0.1603
R17842 GNDA.t696 GNDA.t549 0.1603
R17843 GNDA.t611 GNDA.t696 0.1603
R17844 GNDA.t214 GNDA.t611 0.1603
R17845 GNDA.t343 GNDA.t214 0.1603
R17846 GNDA.t277 GNDA.t343 0.1603
R17847 GNDA.t365 GNDA.t527 0.1603
R17848 GNDA.t234 GNDA.t365 0.1603
R17849 GNDA.t461 GNDA.t234 0.1603
R17850 GNDA.t377 GNDA.t461 0.1603
R17851 GNDA.t246 GNDA.t377 0.1603
R17852 GNDA.t313 GNDA.t246 0.1603
R17853 GNDA.t726 GNDA.t313 0.1603
R17854 GNDA.t557 GNDA.t645 0.1603
R17855 GNDA.t703 GNDA.t557 0.1603
R17856 GNDA.t449 GNDA.t703 0.1603
R17857 GNDA.t222 GNDA.t449 0.1603
R17858 GNDA.t351 GNDA.t222 0.1603
R17859 GNDA.t516 GNDA.t351 0.1603
R17860 GNDA.t415 GNDA.t516 0.1603
R17861 GNDA.t535 GNDA.t682 0.1603
R17862 GNDA.t373 GNDA.t535 0.1603
R17863 GNDA.t732 GNDA.t373 0.1603
R17864 GNDA.t546 GNDA.t732 0.1603
R17865 GNDA.t385 GNDA.t546 0.1603
R17866 GNDA.t485 GNDA.t385 0.1603
R17867 GNDA.t321 GNDA.t485 0.1603
R17868 GNDA.t712 GNDA.t255 0.1603
R17869 GNDA.t457 GNDA.t712 0.1603
R17870 GNDA.t472 GNDA.t457 0.1603
R17871 GNDA.t361 GNDA.t472 0.1603
R17872 GNDA.t524 GNDA.t361 0.1603
R17873 GNDA.t672 GNDA.t524 0.1603
R17874 GNDA.t587 GNDA.t672 0.1603
R17875 GNDA.t690 GNDA.t293 0.1603
R17876 GNDA.t542 GNDA.t690 0.1603
R17877 GNDA.t634 GNDA.t542 0.1603
R17878 GNDA.t699 GNDA.t634 0.1603
R17879 GNDA.t553 GNDA.t699 0.1603
R17880 GNDA.t642 GNDA.t553 0.1603
R17881 GNDA.t493 GNDA.t642 0.1603
R17882 GNDA.t309 GNDA.t393 0.1603
R17883 GNDA.t479 GNDA.t309 0.1603
R17884 GNDA.t618 GNDA.t479 0.1603
R17885 GNDA.t532 GNDA.t618 0.1603
R17886 GNDA.t680 GNDA.t532 0.1603
R17887 GNDA.t282 GNDA.t680 0.1603
R17888 GNDA.t195 GNDA.t282 0.1603
R17889 GNDA.t555 GNDA.t701 0.1603
R17890 GNDA.t391 GNDA.t555 0.1603
R17891 GNDA.t495 GNDA.t391 0.1603
R17892 GNDA.t567 GNDA.t495 0.1603
R17893 GNDA.t402 GNDA.t567 0.1603
R17894 GNDA.t503 GNDA.t402 0.1603
R17895 GNDA.t337 GNDA.t503 0.1603
R17896 GNDA.t186 GNDA.t272 0.1603
R17897 GNDA.t319 GNDA.t186 0.1603
R17898 GNDA.t484 GNDA.t319 0.1603
R17899 GNDA.t383 GNDA.t484 0.1603
R17900 GNDA.t544 GNDA.t383 0.1603
R17901 GNDA.t691 GNDA.t544 0.1603
R17902 GNDA.t606 GNDA.t691 0.1603
R17903 GNDA.t710 GNDA.t455 0.1603
R17904 GNDA.t563 GNDA.t710 0.1603
R17905 GNDA.t651 GNDA.t563 0.1603
R17906 GNDA.t722 GNDA.t651 0.1603
R17907 GNDA.t576 GNDA.t722 0.1603
R17908 GNDA.t660 GNDA.t576 0.1603
R17909 GNDA.t512 GNDA.t660 0.1603
R17910 GNDA.t325 GNDA.t411 0.1603
R17911 GNDA.t491 GNDA.t325 0.1603
R17912 GNDA.t641 GNDA.t491 0.1603
R17913 GNDA.t551 GNDA.t641 0.1603
R17914 GNDA.t697 GNDA.t551 0.1603
R17915 GNDA.t304 GNDA.t697 0.1603
R17916 GNDA.t217 GNDA.t304 0.1603
R17917 GNDA.t463 GNDA.t475 0.1603
R17918 GNDA.t716 GNDA.t463 0.1603
R17919 GNDA.t258 GNDA.t716 0.1603
R17920 GNDA.t316 GNDA.t258 0.1603
R17921 GNDA.t183 GNDA.t316 0.1603
R17922 GNDA.t268 GNDA.t183 0.1603
R17923 GNDA.t666 GNDA.t268 0.1603
R17924 GNDA.t501 GNDA.t583 0.1603
R17925 GNDA.t648 GNDA.t501 0.1603
R17926 GNDA.t249 GNDA.t648 0.1603
R17927 GNDA.t707 GNDA.t249 0.1603
R17928 GNDA.t452 GNDA.t707 0.1603
R17929 GNDA.t440 GNDA.t452 0.1603
R17930 GNDA.t356 GNDA.t440 0.1603
R17931 GNDA.t184 GNDA.t318 0.1603
R17932 GNDA.t582 GNDA.t184 0.1603
R17933 GNDA.t669 GNDA.t582 0.1603
R17934 GNDA.t192 GNDA.t669 0.1603
R17935 GNDA.t592 GNDA.t192 0.1603
R17936 GNDA.t676 GNDA.t592 0.1603
R17937 GNDA.t528 GNDA.t676 0.1603
R17938 GNDA.t346 GNDA.t432 0.1603
R17939 GNDA.t510 GNDA.t346 0.1603
R17940 GNDA.t657 GNDA.t510 0.1603
R17941 GNDA.t573 GNDA.t657 0.1603
R17942 GNDA.t719 GNDA.t573 0.1603
R17943 GNDA.t462 GNDA.t719 0.1603
R17944 GNDA.t239 GNDA.t462 0.1603
R17945 GNDA.t324 GNDA.t490 0.1603
R17946 GNDA.t191 GNDA.t324 0.1603
R17947 GNDA.t280 GNDA.t191 0.1603
R17948 GNDA.t335 GNDA.t280 0.1603
R17949 GNDA.t202 GNDA.t335 0.1603
R17950 GNDA.t290 GNDA.t202 0.1603
R17951 GNDA.t687 GNDA.t290 0.1603
R17952 GNDA.t517 GNDA.t601 0.1603
R17953 GNDA.t664 GNDA.t517 0.1603
R17954 GNDA.t266 GNDA.t664 0.1603
R17955 GNDA.t727 GNDA.t266 0.1603
R17956 GNDA.t314 GNDA.t727 0.1603
R17957 GNDA.t734 GNDA.t314 0.1603
R17958 GNDA.t378 GNDA.t734 0.1603
R17959 GNDA.t497 GNDA.t646 0.1603
R17960 GNDA.t330 GNDA.t497 0.1603
R17961 GNDA.t417 GNDA.t330 0.1603
R17962 GNDA.t507 GNDA.t417 0.1603
R17963 GNDA.t341 GNDA.t507 0.1603
R17964 GNDA.t427 GNDA.t341 0.1603
R17965 GNDA.t298 GNDA.t427 0.1603
R17966 GNDA.t674 GNDA.t213 0.1603
R17967 GNDA.t276 GNDA.t674 0.1603
R17968 GNDA.t407 GNDA.t276 0.1603
R17969 GNDA.t323 GNDA.t407 0.1603
R17970 GNDA.t487 GNDA.t323 0.1603
R17971 GNDA.t636 GNDA.t487 0.1603
R17972 GNDA.t547 GNDA.t636 0.1603
R17973 GNDA.t340 GNDA.t508 0.1603
R17974 GNDA.t210 GNDA.t340 0.1603
R17975 GNDA.t300 GNDA.t210 0.1603
R17976 GNDA.t353 GNDA.t300 0.1603
R17977 GNDA.t224 GNDA.t353 0.1603
R17978 GNDA.t450 GNDA.t224 0.1603
R17979 GNDA.t704 GNDA.t450 0.1603
R17980 GNDA.t537 GNDA.t625 0.1603
R17981 GNDA.t683 GNDA.t537 0.1603
R17982 GNDA.t287 GNDA.t683 0.1603
R17983 GNDA.t200 GNDA.t287 0.1603
R17984 GNDA.t331 GNDA.t200 0.1603
R17985 GNDA.t498 GNDA.t331 0.1603
R17986 GNDA.t395 GNDA.t498 0.1603
R17987 GNDA.t514 GNDA.t663 0.1603
R17988 GNDA.t349 GNDA.t514 0.1603
R17989 GNDA.t437 GNDA.t349 0.1603
R17990 GNDA.t526 GNDA.t437 0.1603
R17991 GNDA.t363 GNDA.t526 0.1603
R17992 GNDA.t473 GNDA.t363 0.1603
R17993 GNDA.t459 GNDA.t473 0.1603
R17994 GNDA.t692 GNDA.t235 0.1603
R17995 GNDA.t295 GNDA.t692 0.1603
R17996 GNDA.t425 GNDA.t295 0.1603
R17997 GNDA.t339 GNDA.t425 0.1603
R17998 GNDA.t504 GNDA.t339 0.1603
R17999 GNDA.t654 GNDA.t504 0.1603
R18000 GNDA.t566 GNDA.t654 0.1603
R18001 GNDA.t671 GNDA.t273 0.1603
R18002 GNDA.t521 GNDA.t671 0.1603
R18003 GNDA.t608 GNDA.t521 0.1603
R18004 GNDA.t681 GNDA.t608 0.1603
R18005 GNDA.t533 GNDA.t681 0.1603
R18006 GNDA.t620 GNDA.t533 0.1603
R18007 GNDA.t481 GNDA.t620 0.1603
R18008 GNDA.t305 GNDA.t374 0.1603
R18009 GNDA.t434 GNDA.t305 0.1603
R18010 GNDA.t596 GNDA.t434 0.1603
R18011 GNDA.t513 GNDA.t596 0.1603
R18012 GNDA.t661 GNDA.t513 0.1603
R18013 GNDA.t263 GNDA.t661 0.1603
R18014 GNDA.t724 GNDA.t263 0.1603
R18015 GNDA.t260 GNDA.t390 0.1603
R18016 GNDA.t656 GNDA.t260 0.1603
R18017 GNDA.t196 GNDA.t656 0.1603
R18018 GNDA.t269 GNDA.t196 0.1603
R18019 GNDA.t668 GNDA.t269 0.1603
R18020 GNDA.t206 GNDA.t668 0.1603
R18021 GNDA.t603 GNDA.t206 0.1603
R18022 GNDA.t420 GNDA.t520 0.1603
R18023 GNDA.t584 GNDA.t420 0.1603
R18024 GNDA.t185 GNDA.t584 0.1603
R18025 GNDA.t649 GNDA.t185 0.1603
R18026 GNDA.t251 GNDA.t649 0.1603
R18027 GNDA.t381 GNDA.t251 0.1603
R18028 GNDA.t454 GNDA.t381 0.1603
R18029 GNDA.t670 GNDA.t271 0.1603
R18030 GNDA.t519 GNDA.t670 0.1603
R18031 GNDA.t605 GNDA.t519 0.1603
R18032 GNDA.t679 GNDA.t605 0.1603
R18033 GNDA.t531 GNDA.t679 0.1603
R18034 GNDA.t616 GNDA.t531 0.1603
R18035 GNDA.t478 GNDA.t616 0.1603
R18036 GNDA.t303 GNDA.t371 0.1603
R18037 GNDA.t431 GNDA.t303 0.1603
R18038 GNDA.t594 GNDA.t431 0.1603
R18039 GNDA.t511 GNDA.t594 0.1603
R18040 GNDA.t659 GNDA.t511 0.1603
R18041 GNDA.t261 GNDA.t659 0.1603
R18042 GNDA.t720 GNDA.t261 0.1603
R18043 GNDA.t281 GNDA.t410 0.1603
R18044 GNDA.t675 GNDA.t281 0.1603
R18045 GNDA.t216 GNDA.t675 0.1603
R18046 GNDA.t292 GNDA.t216 0.1603
R18047 GNDA.t688 GNDA.t292 0.1603
R18048 GNDA.t229 GNDA.t688 0.1603
R18049 GNDA.t629 GNDA.t229 0.1603
R18050 GNDA.t439 GNDA.t540 0.1603
R18051 GNDA.t600 GNDA.t439 0.1603
R18052 GNDA.t203 GNDA.t600 0.1603
R18053 GNDA.t665 GNDA.t203 0.1603
R18054 GNDA.t267 GNDA.t665 0.1603
R18055 GNDA.t399 GNDA.t267 0.1603
R18056 GNDA.t315 GNDA.t399 0.1603
R18057 GNDA.t419 GNDA.t581 0.1603
R18058 GNDA.t286 GNDA.t419 0.1603
R18059 GNDA.t355 GNDA.t286 0.1603
R18060 GNDA.t428 GNDA.t355 0.1603
R18061 GNDA.t299 GNDA.t428 0.1603
R18062 GNDA.t367 GNDA.t299 0.1603
R18063 GNDA.t238 GNDA.t367 0.1603
R18064 GNDA.t612 GNDA.t695 0.1603
R18065 GNDA.t212 GNDA.t612 0.1603
R18066 GNDA.t345 GNDA.t212 0.1603
R18067 GNDA.t278 GNDA.t345 0.1603
R18068 GNDA.t406 GNDA.t278 0.1603
R18069 GNDA.t572 GNDA.t406 0.1603
R18070 GNDA.t488 GNDA.t572 0.1603
R18071 GNDA.t302 GNDA.t430 0.1603
R18072 GNDA.t694 GNDA.t302 0.1603
R18073 GNDA.t241 GNDA.t694 0.1603
R18074 GNDA.t451 GNDA.t241 0.1603
R18075 GNDA.t706 GNDA.t451 0.1603
R18076 GNDA.t248 GNDA.t706 0.1603
R18077 GNDA.t647 GNDA.t248 0.1603
R18078 GNDA.t733 GNDA.t562 0.1603
R18079 GNDA.t627 GNDA.t733 0.1603
R18080 GNDA.t227 GNDA.t627 0.1603
R18081 GNDA.t686 GNDA.t227 0.1603
R18082 GNDA.t289 GNDA.t686 0.1603
R18083 GNDA.t418 GNDA.t289 0.1603
R18084 GNDA.t334 GNDA.t418 0.1603
R18085 GNDA.t438 GNDA.t599 0.1603
R18086 GNDA.t448 GNDA.t438 0.1603
R18087 GNDA.t379 GNDA.t448 0.1603
R18088 GNDA.t474 GNDA.t379 0.1603
R18089 GNDA.t460 GNDA.t474 0.1603
R18090 GNDA.t386 GNDA.t460 0.1603
R18091 GNDA.t256 GNDA.t386 0.1603
R18092 GNDA.t635 GNDA.t715 0.1603
R18093 GNDA.t236 GNDA.t635 0.1603
R18094 GNDA.t366 GNDA.t236 0.1603
R18095 GNDA.t297 GNDA.t366 0.1603
R18096 GNDA.t426 GNDA.t297 0.1603
R18097 GNDA.t590 GNDA.t426 0.1603
R18098 GNDA.t506 GNDA.t590 0.1603
R18099 GNDA.t609 GNDA.t209 0.1603
R18100 GNDA.t444 GNDA.t609 0.1603
R18101 GNDA.t548 GNDA.t444 0.1603
R18102 GNDA.t621 GNDA.t548 0.1603
R18103 GNDA.t730 GNDA.t621 0.1603
R18104 GNDA.t559 GNDA.t730 0.1603
R18105 GNDA.t394 GNDA.t559 0.1603
R18106 GNDA.t244 GNDA.t312 0.1603
R18107 GNDA.t375 GNDA.t244 0.1603
R18108 GNDA.t536 GNDA.t375 0.1603
R18109 GNDA.t435 GNDA.t536 0.1603
R18110 GNDA.t598 GNDA.t435 0.1603
R18111 GNDA.t198 GNDA.t598 0.1603
R18112 GNDA.t662 GNDA.t198 0.1603
R18113 GNDA.t731 GNDA.t623 0.1603
R18114 GNDA.t311 GNDA.t731 0.1603
R18115 GNDA.t397 GNDA.t311 0.1603
R18116 GNDA.t486 GNDA.t397 0.1603
R18117 GNDA.t322 GNDA.t486 0.1603
R18118 GNDA.t405 GNDA.t322 0.1603
R18119 GNDA.t275 GNDA.t405 0.1603
R18120 GNDA.t653 GNDA.t190 0.1603
R18121 GNDA.t254 GNDA.t653 0.1603
R18122 GNDA.t467 GNDA.t254 0.1603
R18123 GNDA.t458 GNDA.t467 0.1603
R18124 GNDA.t471 GNDA.t458 0.1603
R18125 GNDA.t610 GNDA.t471 0.1603
R18126 GNDA.t523 GNDA.t610 0.1603
R18127 GNDA.t633 GNDA.t233 0.1603
R18128 GNDA.t483 GNDA.t633 0.1603
R18129 GNDA.t569 GNDA.t483 0.1603
R18130 GNDA.t644 GNDA.t569 0.1603
R18131 GNDA.t494 GNDA.t644 0.1603
R18132 GNDA.t578 GNDA.t494 0.1603
R18133 GNDA.t414 GNDA.t578 0.1603
R18134 GNDA.t262 GNDA.t329 0.1603
R18135 GNDA.t392 GNDA.t262 0.1603
R18136 GNDA.t556 GNDA.t392 0.1603
R18137 GNDA.t480 GNDA.t556 0.1603
R18138 GNDA.t617 GNDA.t480 0.1603
R18139 GNDA.t221 GNDA.t617 0.1603
R18140 GNDA.t678 GNDA.t221 0.1603
R18141 GNDA.t243 GNDA.t372 0.1603
R18142 GNDA.t640 GNDA.t243 0.1603
R18143 GNDA.t723 GNDA.t640 0.1603
R18144 GNDA.t253 GNDA.t723 0.1603
R18145 GNDA.t650 GNDA.t253 0.1603
R18146 GNDA.t187 GNDA.t650 0.1603
R18147 GNDA.t586 GNDA.t187 0.1603
R18148 GNDA.t400 GNDA.t502 0.1603
R18149 GNDA.t564 GNDA.t400 0.1603
R18150 GNDA.t711 GNDA.t564 0.1603
R18151 GNDA.t630 GNDA.t711 0.1603
R18152 GNDA.t230 GNDA.t630 0.1603
R18153 GNDA.t360 GNDA.t230 0.1603
R18154 GNDA.t291 GNDA.t360 0.1603
R18155 GNDA.t380 GNDA.t541 0.1603
R18156 GNDA.t247 GNDA.t380 0.1603
R18157 GNDA.t317 GNDA.t247 0.1603
R18158 GNDA.t389 GNDA.t317 0.1603
R18159 GNDA.t257 GNDA.t389 0.1603
R18160 GNDA.t326 GNDA.t257 0.1603
R18161 GNDA.t194 GNDA.t326 0.1603
R18162 GNDA.t574 GNDA.t658 0.1603
R18163 GNDA.t718 GNDA.t574 0.1603
R18164 GNDA.t307 GNDA.t718 0.1603
R18165 GNDA.t240 GNDA.t307 0.1603
R18166 GNDA.t368 GNDA.t240 0.1603
R18167 GNDA.t530 GNDA.t368 0.1603
R18168 GNDA.t429 GNDA.t530 0.1603
R18169 GNDA.t558 GNDA.t482 0.1603
R18170 GNDA.t396 GNDA.t558 0.1603
R18171 GNDA.t264 GNDA.t396 0.1603
R18172 GNDA.t333 GNDA.t264 0.1603
R18173 GNDA.t199 GNDA.t333 0.1603
R18174 GNDA.t597 GNDA.t199 0.1603
R18175 GNDA.t685 GNDA.t597 0.1603
R18176 GNDA.t421 GNDA.n2073 0.159278
R18177 GNDA.t283 GNDA.n2074 0.159278
R18178 GNDA.t673 GNDA.n2075 0.159278
R18179 GNDA.t265 GNDA.n2076 0.159278
R18180 GNDA.t655 GNDA.n2077 0.159278
R18181 GNDA.t500 GNDA.n2078 0.159278
R18182 GNDA.t637 GNDA.n2079 0.159278
R18183 GNDA.t735 GNDA.n2080 0.159278
R18184 GNDA.t308 GNDA.n2081 0.159278
R18185 GNDA.t442 GNDA.n2082 0.159278
R18186 GNDA.t310 GNDA.n2083 0.159278
R18187 GNDA.t713 GNDA.n2084 0.159278
R18188 GNDA.t560 GNDA.n2085 0.159278
R18189 GNDA.t693 GNDA.n2086 0.159278
R18190 GNDA.t539 GNDA.n2087 0.159278
R18191 GNDA.t369 GNDA.n2088 0.159278
R18192 GNDA.t518 GNDA.n2089 0.159278
R18193 GNDA.t348 GNDA.n2090 0.159278
R18194 GNDA.t207 GNDA.n2091 0.159278
R18195 GNDA.t328 GNDA.n2092 0.159278
R18196 GNDA.t189 GNDA.n2093 0.159278
R18197 GNDA.t580 GNDA.n2094 0.159278
R18198 GNDA.t408 GNDA.n2095 0.159278
R18199 GNDA.t561 GNDA.n2096 0.159278
R18200 GNDA.t409 GNDA.n2097 0.159278
R18201 GNDA.t270 GNDA.n2098 0.159278
R18202 GNDA.t388 GNDA.n2099 0.159278
R18203 GNDA.t252 GNDA.n2100 0.159278
R18204 GNDA.t643 GNDA.n2101 0.159278
R18205 GNDA.t232 GNDA.n2102 0.159278
R18206 GNDA.t622 GNDA.n2103 0.159278
R18207 GNDA.n6272 GNDA.n6271 0.15675
R18208 GNDA.n6268 GNDA.n6267 0.15675
R18209 GNDA.n4662 GNDA.n1597 0.146333
R18210 GNDA.n4667 GNDA.n4662 0.146333
R18211 GNDA.n4668 GNDA.n4667 0.146333
R18212 GNDA.n4678 GNDA.n4677 0.146333
R18213 GNDA.n4681 GNDA.n4678 0.146333
R18214 GNDA.n4681 GNDA.n4658 0.146333
R18215 GNDA.n4691 GNDA.n4656 0.146333
R18216 GNDA.n4697 GNDA.n4656 0.146333
R18217 GNDA.n4698 GNDA.n4697 0.146333
R18218 GNDA.n4708 GNDA.n4707 0.146333
R18219 GNDA.n4711 GNDA.n4708 0.146333
R18220 GNDA.n4711 GNDA.n4652 0.146333
R18221 GNDA.n4721 GNDA.n4650 0.146333
R18222 GNDA.n4727 GNDA.n4650 0.146333
R18223 GNDA.n4728 GNDA.n4727 0.146333
R18224 GNDA.n4738 GNDA.n4737 0.146333
R18225 GNDA.n4741 GNDA.n4738 0.146333
R18226 GNDA.n4741 GNDA.n4646 0.146333
R18227 GNDA.n4751 GNDA.n4644 0.146333
R18228 GNDA.n4757 GNDA.n4644 0.146333
R18229 GNDA.n4758 GNDA.n4757 0.146333
R18230 GNDA.n4768 GNDA.n4767 0.146333
R18231 GNDA.n4771 GNDA.n4768 0.146333
R18232 GNDA.n4771 GNDA.n4640 0.146333
R18233 GNDA.n5688 GNDA.n5685 0.146333
R18234 GNDA.n5694 GNDA.n5685 0.146333
R18235 GNDA.n5695 GNDA.n5694 0.146333
R18236 GNDA.n5705 GNDA.n5704 0.146333
R18237 GNDA.n5708 GNDA.n5705 0.146333
R18238 GNDA.n5708 GNDA.n5681 0.146333
R18239 GNDA.n5718 GNDA.n5679 0.146333
R18240 GNDA.n5724 GNDA.n5679 0.146333
R18241 GNDA.n5725 GNDA.n5724 0.146333
R18242 GNDA.n5735 GNDA.n5734 0.146333
R18243 GNDA.n5738 GNDA.n5735 0.146333
R18244 GNDA.n5738 GNDA.n5675 0.146333
R18245 GNDA.n5748 GNDA.n5673 0.146333
R18246 GNDA.n5754 GNDA.n5673 0.146333
R18247 GNDA.n5755 GNDA.n5754 0.146333
R18248 GNDA.n5765 GNDA.n5764 0.146333
R18249 GNDA.n5768 GNDA.n5765 0.146333
R18250 GNDA.n5768 GNDA.n5669 0.146333
R18251 GNDA.n5778 GNDA.n5667 0.146333
R18252 GNDA.n5784 GNDA.n5667 0.146333
R18253 GNDA.n5785 GNDA.n5784 0.146333
R18254 GNDA.n5795 GNDA.n5794 0.146333
R18255 GNDA.n5798 GNDA.n5795 0.146333
R18256 GNDA.n5798 GNDA.n5663 0.146333
R18257 GNDA.n2700 GNDA.n2694 0.146333
R18258 GNDA.n2704 GNDA.n2694 0.146333
R18259 GNDA.n2705 GNDA.n2704 0.146333
R18260 GNDA.n2713 GNDA.n2712 0.146333
R18261 GNDA.n2716 GNDA.n2713 0.146333
R18262 GNDA.n2716 GNDA.n2686 0.146333
R18263 GNDA.n2724 GNDA.n2682 0.146333
R18264 GNDA.n2728 GNDA.n2682 0.146333
R18265 GNDA.n2729 GNDA.n2728 0.146333
R18266 GNDA.n2737 GNDA.n2736 0.146333
R18267 GNDA.n2740 GNDA.n2737 0.146333
R18268 GNDA.n2740 GNDA.n2674 0.146333
R18269 GNDA.n2748 GNDA.n2670 0.146333
R18270 GNDA.n2752 GNDA.n2670 0.146333
R18271 GNDA.n2753 GNDA.n2752 0.146333
R18272 GNDA.n2761 GNDA.n2760 0.146333
R18273 GNDA.n2764 GNDA.n2761 0.146333
R18274 GNDA.n2764 GNDA.n2662 0.146333
R18275 GNDA.n2772 GNDA.n2658 0.146333
R18276 GNDA.n2776 GNDA.n2658 0.146333
R18277 GNDA.n2777 GNDA.n2776 0.146333
R18278 GNDA.n2785 GNDA.n2784 0.146333
R18279 GNDA.n2788 GNDA.n2785 0.146333
R18280 GNDA.n2788 GNDA.n2652 0.146333
R18281 GNDA.n5967 GNDA.n1369 0.146333
R18282 GNDA.n5972 GNDA.n5967 0.146333
R18283 GNDA.n5973 GNDA.n5972 0.146333
R18284 GNDA.n5983 GNDA.n5982 0.146333
R18285 GNDA.n5986 GNDA.n5983 0.146333
R18286 GNDA.n5986 GNDA.n5963 0.146333
R18287 GNDA.n5996 GNDA.n5961 0.146333
R18288 GNDA.n6002 GNDA.n5961 0.146333
R18289 GNDA.n6003 GNDA.n6002 0.146333
R18290 GNDA.n6013 GNDA.n6012 0.146333
R18291 GNDA.n6016 GNDA.n6013 0.146333
R18292 GNDA.n6016 GNDA.n5957 0.146333
R18293 GNDA.n6026 GNDA.n5955 0.146333
R18294 GNDA.n6032 GNDA.n5955 0.146333
R18295 GNDA.n6033 GNDA.n6032 0.146333
R18296 GNDA.n6043 GNDA.n6042 0.146333
R18297 GNDA.n6046 GNDA.n6043 0.146333
R18298 GNDA.n6046 GNDA.n5951 0.146333
R18299 GNDA.n6056 GNDA.n5949 0.146333
R18300 GNDA.n6062 GNDA.n5949 0.146333
R18301 GNDA.n6063 GNDA.n6062 0.146333
R18302 GNDA.n6073 GNDA.n6072 0.146333
R18303 GNDA.n6076 GNDA.n6073 0.146333
R18304 GNDA.n6076 GNDA.n5945 0.146333
R18305 GNDA.n1425 GNDA.n1424 0.146333
R18306 GNDA.n1426 GNDA.n1425 0.146333
R18307 GNDA.n1427 GNDA.n1426 0.146333
R18308 GNDA.n1431 GNDA.n1430 0.146333
R18309 GNDA.n1432 GNDA.n1431 0.146333
R18310 GNDA.n1433 GNDA.n1432 0.146333
R18311 GNDA.n1437 GNDA.n1436 0.146333
R18312 GNDA.n1438 GNDA.n1437 0.146333
R18313 GNDA.n1439 GNDA.n1438 0.146333
R18314 GNDA.n1443 GNDA.n1442 0.146333
R18315 GNDA.n1444 GNDA.n1443 0.146333
R18316 GNDA.n1445 GNDA.n1444 0.146333
R18317 GNDA.n1449 GNDA.n1448 0.146333
R18318 GNDA.n1450 GNDA.n1449 0.146333
R18319 GNDA.n1451 GNDA.n1450 0.146333
R18320 GNDA.n1455 GNDA.n1454 0.146333
R18321 GNDA.n1456 GNDA.n1455 0.146333
R18322 GNDA.n1457 GNDA.n1456 0.146333
R18323 GNDA.n1461 GNDA.n1460 0.146333
R18324 GNDA.n1462 GNDA.n1461 0.146333
R18325 GNDA.n1463 GNDA.n1462 0.146333
R18326 GNDA.n1467 GNDA.n1466 0.146333
R18327 GNDA.n1468 GNDA.n1467 0.146333
R18328 GNDA.n1469 GNDA.n1468 0.146333
R18329 GNDA.n3637 GNDA.n3633 0.146333
R18330 GNDA.n3643 GNDA.n3633 0.146333
R18331 GNDA.n3644 GNDA.n3643 0.146333
R18332 GNDA.n3654 GNDA.n3653 0.146333
R18333 GNDA.n3657 GNDA.n3654 0.146333
R18334 GNDA.n3657 GNDA.n3629 0.146333
R18335 GNDA.n3667 GNDA.n3627 0.146333
R18336 GNDA.n3673 GNDA.n3627 0.146333
R18337 GNDA.n3674 GNDA.n3673 0.146333
R18338 GNDA.n3684 GNDA.n3683 0.146333
R18339 GNDA.n3687 GNDA.n3684 0.146333
R18340 GNDA.n3687 GNDA.n3623 0.146333
R18341 GNDA.n3697 GNDA.n3621 0.146333
R18342 GNDA.n3703 GNDA.n3621 0.146333
R18343 GNDA.n3704 GNDA.n3703 0.146333
R18344 GNDA.n3714 GNDA.n3713 0.146333
R18345 GNDA.n3717 GNDA.n3714 0.146333
R18346 GNDA.n3717 GNDA.n3617 0.146333
R18347 GNDA.n3727 GNDA.n3615 0.146333
R18348 GNDA.n3733 GNDA.n3615 0.146333
R18349 GNDA.n3734 GNDA.n3733 0.146333
R18350 GNDA.n3744 GNDA.n3743 0.146333
R18351 GNDA.n3747 GNDA.n3744 0.146333
R18352 GNDA.n3747 GNDA.n3611 0.146333
R18353 GNDA.n3297 GNDA.n3296 0.146333
R18354 GNDA.n3298 GNDA.n3297 0.146333
R18355 GNDA.n3299 GNDA.n3298 0.146333
R18356 GNDA.n3303 GNDA.n3302 0.146333
R18357 GNDA.n3304 GNDA.n3303 0.146333
R18358 GNDA.n3305 GNDA.n3304 0.146333
R18359 GNDA.n3309 GNDA.n3308 0.146333
R18360 GNDA.n3310 GNDA.n3309 0.146333
R18361 GNDA.n3311 GNDA.n3310 0.146333
R18362 GNDA.n3315 GNDA.n3314 0.146333
R18363 GNDA.n3316 GNDA.n3315 0.146333
R18364 GNDA.n3317 GNDA.n3316 0.146333
R18365 GNDA.n3321 GNDA.n3320 0.146333
R18366 GNDA.n3322 GNDA.n3321 0.146333
R18367 GNDA.n3323 GNDA.n3322 0.146333
R18368 GNDA.n3327 GNDA.n3326 0.146333
R18369 GNDA.n3328 GNDA.n3327 0.146333
R18370 GNDA.n3329 GNDA.n3328 0.146333
R18371 GNDA.n3333 GNDA.n3332 0.146333
R18372 GNDA.n3334 GNDA.n3333 0.146333
R18373 GNDA.n3335 GNDA.n3334 0.146333
R18374 GNDA.n3339 GNDA.n3338 0.146333
R18375 GNDA.n3340 GNDA.n3339 0.146333
R18376 GNDA.n3341 GNDA.n3340 0.146333
R18377 GNDA.n5118 GNDA.n5070 0.146333
R18378 GNDA.n5123 GNDA.n5118 0.146333
R18379 GNDA.n5124 GNDA.n5123 0.146333
R18380 GNDA.n5134 GNDA.n5133 0.146333
R18381 GNDA.n5137 GNDA.n5134 0.146333
R18382 GNDA.n5137 GNDA.n5114 0.146333
R18383 GNDA.n5147 GNDA.n5112 0.146333
R18384 GNDA.n5153 GNDA.n5112 0.146333
R18385 GNDA.n5154 GNDA.n5153 0.146333
R18386 GNDA.n5164 GNDA.n5163 0.146333
R18387 GNDA.n5167 GNDA.n5164 0.146333
R18388 GNDA.n5167 GNDA.n5108 0.146333
R18389 GNDA.n5177 GNDA.n5106 0.146333
R18390 GNDA.n5183 GNDA.n5106 0.146333
R18391 GNDA.n5184 GNDA.n5183 0.146333
R18392 GNDA.n5194 GNDA.n5193 0.146333
R18393 GNDA.n5197 GNDA.n5194 0.146333
R18394 GNDA.n5197 GNDA.n5102 0.146333
R18395 GNDA.n5207 GNDA.n5100 0.146333
R18396 GNDA.n5213 GNDA.n5100 0.146333
R18397 GNDA.n5214 GNDA.n5213 0.146333
R18398 GNDA.n5224 GNDA.n5223 0.146333
R18399 GNDA.n5227 GNDA.n5224 0.146333
R18400 GNDA.n5227 GNDA.n5096 0.146333
R18401 GNDA.n5237 GNDA.n5236 0.146333
R18402 GNDA.n5238 GNDA.n5237 0.146333
R18403 GNDA.n5239 GNDA.n5238 0.146333
R18404 GNDA.n5243 GNDA.n5242 0.146333
R18405 GNDA.n5244 GNDA.n5243 0.146333
R18406 GNDA.n5245 GNDA.n5244 0.146333
R18407 GNDA.n5249 GNDA.n5248 0.146333
R18408 GNDA.n5250 GNDA.n5249 0.146333
R18409 GNDA.n5251 GNDA.n5250 0.146333
R18410 GNDA.n5255 GNDA.n5254 0.146333
R18411 GNDA.n5256 GNDA.n5255 0.146333
R18412 GNDA.n5257 GNDA.n5256 0.146333
R18413 GNDA.n5261 GNDA.n5260 0.146333
R18414 GNDA.n5262 GNDA.n5261 0.146333
R18415 GNDA.n5263 GNDA.n5262 0.146333
R18416 GNDA.n5267 GNDA.n5266 0.146333
R18417 GNDA.n5268 GNDA.n5267 0.146333
R18418 GNDA.n5269 GNDA.n5268 0.146333
R18419 GNDA.n5273 GNDA.n5272 0.146333
R18420 GNDA.n5274 GNDA.n5273 0.146333
R18421 GNDA.n5275 GNDA.n5274 0.146333
R18422 GNDA.n5279 GNDA.n5278 0.146333
R18423 GNDA.n5280 GNDA.n5279 0.146333
R18424 GNDA.n5281 GNDA.n5280 0.146333
R18425 GNDA.n5405 GNDA.n5068 0.146333
R18426 GNDA.n5411 GNDA.n5068 0.146333
R18427 GNDA.n5412 GNDA.n5411 0.146333
R18428 GNDA.n5422 GNDA.n5421 0.146333
R18429 GNDA.n5425 GNDA.n5422 0.146333
R18430 GNDA.n5425 GNDA.n5064 0.146333
R18431 GNDA.n5435 GNDA.n5062 0.146333
R18432 GNDA.n5441 GNDA.n5062 0.146333
R18433 GNDA.n5442 GNDA.n5441 0.146333
R18434 GNDA.n5452 GNDA.n5451 0.146333
R18435 GNDA.n5455 GNDA.n5452 0.146333
R18436 GNDA.n5455 GNDA.n5058 0.146333
R18437 GNDA.n5465 GNDA.n5056 0.146333
R18438 GNDA.n5471 GNDA.n5056 0.146333
R18439 GNDA.n5472 GNDA.n5471 0.146333
R18440 GNDA.n5482 GNDA.n5481 0.146333
R18441 GNDA.n5485 GNDA.n5482 0.146333
R18442 GNDA.n5485 GNDA.n5052 0.146333
R18443 GNDA.n5495 GNDA.n5050 0.146333
R18444 GNDA.n5501 GNDA.n5050 0.146333
R18445 GNDA.n5502 GNDA.n5501 0.146333
R18446 GNDA.n5512 GNDA.n5511 0.146333
R18447 GNDA.n5515 GNDA.n5512 0.146333
R18448 GNDA.n5515 GNDA.n5046 0.146333
R18449 GNDA.n5547 GNDA.n5543 0.146333
R18450 GNDA.n5553 GNDA.n5543 0.146333
R18451 GNDA.n5554 GNDA.n5553 0.146333
R18452 GNDA.n5564 GNDA.n5563 0.146333
R18453 GNDA.n5567 GNDA.n5564 0.146333
R18454 GNDA.n5567 GNDA.n5539 0.146333
R18455 GNDA.n5577 GNDA.n5537 0.146333
R18456 GNDA.n5583 GNDA.n5537 0.146333
R18457 GNDA.n5584 GNDA.n5583 0.146333
R18458 GNDA.n5594 GNDA.n5593 0.146333
R18459 GNDA.n5597 GNDA.n5594 0.146333
R18460 GNDA.n5597 GNDA.n5533 0.146333
R18461 GNDA.n5607 GNDA.n5531 0.146333
R18462 GNDA.n5613 GNDA.n5531 0.146333
R18463 GNDA.n5614 GNDA.n5613 0.146333
R18464 GNDA.n5624 GNDA.n5623 0.146333
R18465 GNDA.n5627 GNDA.n5624 0.146333
R18466 GNDA.n5627 GNDA.n5527 0.146333
R18467 GNDA.n5637 GNDA.n5525 0.146333
R18468 GNDA.n5643 GNDA.n5525 0.146333
R18469 GNDA.n5644 GNDA.n5643 0.146333
R18470 GNDA.n5654 GNDA.n5653 0.146333
R18471 GNDA.n5657 GNDA.n5654 0.146333
R18472 GNDA.n5657 GNDA.n5521 0.146333
R18473 GNDA.n5829 GNDA.n5826 0.146333
R18474 GNDA.n5835 GNDA.n5826 0.146333
R18475 GNDA.n5836 GNDA.n5835 0.146333
R18476 GNDA.n5846 GNDA.n5845 0.146333
R18477 GNDA.n5849 GNDA.n5846 0.146333
R18478 GNDA.n5849 GNDA.n5822 0.146333
R18479 GNDA.n5859 GNDA.n5820 0.146333
R18480 GNDA.n5865 GNDA.n5820 0.146333
R18481 GNDA.n5866 GNDA.n5865 0.146333
R18482 GNDA.n5876 GNDA.n5875 0.146333
R18483 GNDA.n5879 GNDA.n5876 0.146333
R18484 GNDA.n5879 GNDA.n5816 0.146333
R18485 GNDA.n5889 GNDA.n5814 0.146333
R18486 GNDA.n5895 GNDA.n5814 0.146333
R18487 GNDA.n5896 GNDA.n5895 0.146333
R18488 GNDA.n5906 GNDA.n5905 0.146333
R18489 GNDA.n5909 GNDA.n5906 0.146333
R18490 GNDA.n5909 GNDA.n5810 0.146333
R18491 GNDA.n5919 GNDA.n5808 0.146333
R18492 GNDA.n5925 GNDA.n5808 0.146333
R18493 GNDA.n5926 GNDA.n5925 0.146333
R18494 GNDA.n5936 GNDA.n5935 0.146333
R18495 GNDA.n5939 GNDA.n5936 0.146333
R18496 GNDA.n5939 GNDA.n5804 0.146333
R18497 GNDA.n4810 GNDA.n1419 0.146333
R18498 GNDA.n4816 GNDA.n1419 0.146333
R18499 GNDA.n4817 GNDA.n4816 0.146333
R18500 GNDA.n4827 GNDA.n4826 0.146333
R18501 GNDA.n4830 GNDA.n4827 0.146333
R18502 GNDA.n4830 GNDA.n1415 0.146333
R18503 GNDA.n4840 GNDA.n1413 0.146333
R18504 GNDA.n4846 GNDA.n1413 0.146333
R18505 GNDA.n4847 GNDA.n4846 0.146333
R18506 GNDA.n4857 GNDA.n4856 0.146333
R18507 GNDA.n4860 GNDA.n4857 0.146333
R18508 GNDA.n4860 GNDA.n1409 0.146333
R18509 GNDA.n4870 GNDA.n1407 0.146333
R18510 GNDA.n4876 GNDA.n1407 0.146333
R18511 GNDA.n4877 GNDA.n4876 0.146333
R18512 GNDA.n4887 GNDA.n4886 0.146333
R18513 GNDA.n4890 GNDA.n4887 0.146333
R18514 GNDA.n4890 GNDA.n1403 0.146333
R18515 GNDA.n4900 GNDA.n1401 0.146333
R18516 GNDA.n4906 GNDA.n1401 0.146333
R18517 GNDA.n4907 GNDA.n4906 0.146333
R18518 GNDA.n4917 GNDA.n4916 0.146333
R18519 GNDA.n4920 GNDA.n4917 0.146333
R18520 GNDA.n4920 GNDA.n1397 0.146333
R18521 GNDA.n4524 GNDA.n4520 0.146333
R18522 GNDA.n4530 GNDA.n4520 0.146333
R18523 GNDA.n4531 GNDA.n4530 0.146333
R18524 GNDA.n4541 GNDA.n4540 0.146333
R18525 GNDA.n4544 GNDA.n4541 0.146333
R18526 GNDA.n4544 GNDA.n4516 0.146333
R18527 GNDA.n4554 GNDA.n4514 0.146333
R18528 GNDA.n4560 GNDA.n4514 0.146333
R18529 GNDA.n4561 GNDA.n4560 0.146333
R18530 GNDA.n4571 GNDA.n4570 0.146333
R18531 GNDA.n4574 GNDA.n4571 0.146333
R18532 GNDA.n4574 GNDA.n4510 0.146333
R18533 GNDA.n4584 GNDA.n4508 0.146333
R18534 GNDA.n4590 GNDA.n4508 0.146333
R18535 GNDA.n4591 GNDA.n4590 0.146333
R18536 GNDA.n4601 GNDA.n4600 0.146333
R18537 GNDA.n4604 GNDA.n4601 0.146333
R18538 GNDA.n4604 GNDA.n4504 0.146333
R18539 GNDA.n4614 GNDA.n4502 0.146333
R18540 GNDA.n4620 GNDA.n4502 0.146333
R18541 GNDA.n4621 GNDA.n4620 0.146333
R18542 GNDA.n4631 GNDA.n4630 0.146333
R18543 GNDA.n4634 GNDA.n4631 0.146333
R18544 GNDA.n4634 GNDA.n4498 0.146333
R18545 GNDA.n4335 GNDA.n4331 0.146333
R18546 GNDA.n4341 GNDA.n4331 0.146333
R18547 GNDA.n4342 GNDA.n4341 0.146333
R18548 GNDA.n4352 GNDA.n4351 0.146333
R18549 GNDA.n4355 GNDA.n4352 0.146333
R18550 GNDA.n4355 GNDA.n4327 0.146333
R18551 GNDA.n4365 GNDA.n4325 0.146333
R18552 GNDA.n4371 GNDA.n4325 0.146333
R18553 GNDA.n4372 GNDA.n4371 0.146333
R18554 GNDA.n4382 GNDA.n4381 0.146333
R18555 GNDA.n4385 GNDA.n4382 0.146333
R18556 GNDA.n4385 GNDA.n4321 0.146333
R18557 GNDA.n4395 GNDA.n4319 0.146333
R18558 GNDA.n4401 GNDA.n4319 0.146333
R18559 GNDA.n4402 GNDA.n4401 0.146333
R18560 GNDA.n4412 GNDA.n4411 0.146333
R18561 GNDA.n4415 GNDA.n4412 0.146333
R18562 GNDA.n4415 GNDA.n4315 0.146333
R18563 GNDA.n4425 GNDA.n4313 0.146333
R18564 GNDA.n4431 GNDA.n4313 0.146333
R18565 GNDA.n4432 GNDA.n4431 0.146333
R18566 GNDA.n4442 GNDA.n4441 0.146333
R18567 GNDA.n4445 GNDA.n4442 0.146333
R18568 GNDA.n4445 GNDA.n4309 0.146333
R18569 GNDA.n4169 GNDA.n1647 0.146333
R18570 GNDA.n4175 GNDA.n1647 0.146333
R18571 GNDA.n4176 GNDA.n4175 0.146333
R18572 GNDA.n4186 GNDA.n4185 0.146333
R18573 GNDA.n4189 GNDA.n4186 0.146333
R18574 GNDA.n4189 GNDA.n1643 0.146333
R18575 GNDA.n4199 GNDA.n1641 0.146333
R18576 GNDA.n4205 GNDA.n1641 0.146333
R18577 GNDA.n4206 GNDA.n4205 0.146333
R18578 GNDA.n4216 GNDA.n4215 0.146333
R18579 GNDA.n4219 GNDA.n4216 0.146333
R18580 GNDA.n4219 GNDA.n1637 0.146333
R18581 GNDA.n4229 GNDA.n1635 0.146333
R18582 GNDA.n4235 GNDA.n1635 0.146333
R18583 GNDA.n4236 GNDA.n4235 0.146333
R18584 GNDA.n4246 GNDA.n4245 0.146333
R18585 GNDA.n4249 GNDA.n4246 0.146333
R18586 GNDA.n4249 GNDA.n1631 0.146333
R18587 GNDA.n4259 GNDA.n1629 0.146333
R18588 GNDA.n4265 GNDA.n1629 0.146333
R18589 GNDA.n4266 GNDA.n4265 0.146333
R18590 GNDA.n4276 GNDA.n4275 0.146333
R18591 GNDA.n4279 GNDA.n4276 0.146333
R18592 GNDA.n4279 GNDA.n1625 0.146333
R18593 GNDA.n1651 GNDA.n1650 0.146333
R18594 GNDA.n1652 GNDA.n1651 0.146333
R18595 GNDA.n1653 GNDA.n1652 0.146333
R18596 GNDA.n1657 GNDA.n1656 0.146333
R18597 GNDA.n1658 GNDA.n1657 0.146333
R18598 GNDA.n1659 GNDA.n1658 0.146333
R18599 GNDA.n1663 GNDA.n1662 0.146333
R18600 GNDA.n1664 GNDA.n1663 0.146333
R18601 GNDA.n1665 GNDA.n1664 0.146333
R18602 GNDA.n1669 GNDA.n1668 0.146333
R18603 GNDA.n1670 GNDA.n1669 0.146333
R18604 GNDA.n1671 GNDA.n1670 0.146333
R18605 GNDA.n1675 GNDA.n1674 0.146333
R18606 GNDA.n1676 GNDA.n1675 0.146333
R18607 GNDA.n1677 GNDA.n1676 0.146333
R18608 GNDA.n1681 GNDA.n1680 0.146333
R18609 GNDA.n1682 GNDA.n1681 0.146333
R18610 GNDA.n1683 GNDA.n1682 0.146333
R18611 GNDA.n1687 GNDA.n1686 0.146333
R18612 GNDA.n1688 GNDA.n1687 0.146333
R18613 GNDA.n1689 GNDA.n1688 0.146333
R18614 GNDA.n1693 GNDA.n1692 0.146333
R18615 GNDA.n1694 GNDA.n1693 0.146333
R18616 GNDA.n1695 GNDA.n1694 0.146333
R18617 GNDA.n3826 GNDA.n3822 0.146333
R18618 GNDA.n3832 GNDA.n3822 0.146333
R18619 GNDA.n3833 GNDA.n3832 0.146333
R18620 GNDA.n3843 GNDA.n3842 0.146333
R18621 GNDA.n3846 GNDA.n3843 0.146333
R18622 GNDA.n3846 GNDA.n3818 0.146333
R18623 GNDA.n3856 GNDA.n3816 0.146333
R18624 GNDA.n3862 GNDA.n3816 0.146333
R18625 GNDA.n3863 GNDA.n3862 0.146333
R18626 GNDA.n3873 GNDA.n3872 0.146333
R18627 GNDA.n3876 GNDA.n3873 0.146333
R18628 GNDA.n3876 GNDA.n3812 0.146333
R18629 GNDA.n3886 GNDA.n3810 0.146333
R18630 GNDA.n3892 GNDA.n3810 0.146333
R18631 GNDA.n3893 GNDA.n3892 0.146333
R18632 GNDA.n3903 GNDA.n3902 0.146333
R18633 GNDA.n3906 GNDA.n3903 0.146333
R18634 GNDA.n3906 GNDA.n3806 0.146333
R18635 GNDA.n3916 GNDA.n3804 0.146333
R18636 GNDA.n3922 GNDA.n3804 0.146333
R18637 GNDA.n3923 GNDA.n3922 0.146333
R18638 GNDA.n3933 GNDA.n3932 0.146333
R18639 GNDA.n3936 GNDA.n3933 0.146333
R18640 GNDA.n3936 GNDA.n3800 0.146333
R18641 GNDA.n3964 GNDA.n1836 0.146333
R18642 GNDA.n3969 GNDA.n3964 0.146333
R18643 GNDA.n3970 GNDA.n3969 0.146333
R18644 GNDA.n3980 GNDA.n3979 0.146333
R18645 GNDA.n3983 GNDA.n3980 0.146333
R18646 GNDA.n3983 GNDA.n3960 0.146333
R18647 GNDA.n3993 GNDA.n3958 0.146333
R18648 GNDA.n3999 GNDA.n3958 0.146333
R18649 GNDA.n4000 GNDA.n3999 0.146333
R18650 GNDA.n4010 GNDA.n4009 0.146333
R18651 GNDA.n4013 GNDA.n4010 0.146333
R18652 GNDA.n4013 GNDA.n3954 0.146333
R18653 GNDA.n4023 GNDA.n3952 0.146333
R18654 GNDA.n4029 GNDA.n3952 0.146333
R18655 GNDA.n4030 GNDA.n4029 0.146333
R18656 GNDA.n4040 GNDA.n4039 0.146333
R18657 GNDA.n4043 GNDA.n4040 0.146333
R18658 GNDA.n4043 GNDA.n3948 0.146333
R18659 GNDA.n4053 GNDA.n3946 0.146333
R18660 GNDA.n4059 GNDA.n3946 0.146333
R18661 GNDA.n4060 GNDA.n4059 0.146333
R18662 GNDA.n4070 GNDA.n4069 0.146333
R18663 GNDA.n4073 GNDA.n4070 0.146333
R18664 GNDA.n4073 GNDA.n3942 0.146333
R18665 GNDA.n3471 GNDA.n1886 0.146333
R18666 GNDA.n3477 GNDA.n1886 0.146333
R18667 GNDA.n3478 GNDA.n3477 0.146333
R18668 GNDA.n3488 GNDA.n3487 0.146333
R18669 GNDA.n3491 GNDA.n3488 0.146333
R18670 GNDA.n3491 GNDA.n1882 0.146333
R18671 GNDA.n3501 GNDA.n1880 0.146333
R18672 GNDA.n3507 GNDA.n1880 0.146333
R18673 GNDA.n3508 GNDA.n3507 0.146333
R18674 GNDA.n3518 GNDA.n3517 0.146333
R18675 GNDA.n3521 GNDA.n3518 0.146333
R18676 GNDA.n3521 GNDA.n1876 0.146333
R18677 GNDA.n3531 GNDA.n1874 0.146333
R18678 GNDA.n3537 GNDA.n1874 0.146333
R18679 GNDA.n3538 GNDA.n3537 0.146333
R18680 GNDA.n3548 GNDA.n3547 0.146333
R18681 GNDA.n3551 GNDA.n3548 0.146333
R18682 GNDA.n3551 GNDA.n1870 0.146333
R18683 GNDA.n3561 GNDA.n1868 0.146333
R18684 GNDA.n3567 GNDA.n1868 0.146333
R18685 GNDA.n3568 GNDA.n3567 0.146333
R18686 GNDA.n3578 GNDA.n3577 0.146333
R18687 GNDA.n3581 GNDA.n3578 0.146333
R18688 GNDA.n3581 GNDA.n1864 0.146333
R18689 GNDA.n2536 GNDA.n2533 0.146333
R18690 GNDA.n2542 GNDA.n2533 0.146333
R18691 GNDA.n2543 GNDA.n2542 0.146333
R18692 GNDA.n2553 GNDA.n2552 0.146333
R18693 GNDA.n2556 GNDA.n2553 0.146333
R18694 GNDA.n2556 GNDA.n2529 0.146333
R18695 GNDA.n2566 GNDA.n2527 0.146333
R18696 GNDA.n2572 GNDA.n2527 0.146333
R18697 GNDA.n2573 GNDA.n2572 0.146333
R18698 GNDA.n2583 GNDA.n2582 0.146333
R18699 GNDA.n2586 GNDA.n2583 0.146333
R18700 GNDA.n2586 GNDA.n2523 0.146333
R18701 GNDA.n2596 GNDA.n2521 0.146333
R18702 GNDA.n2602 GNDA.n2521 0.146333
R18703 GNDA.n2603 GNDA.n2602 0.146333
R18704 GNDA.n2613 GNDA.n2612 0.146333
R18705 GNDA.n2616 GNDA.n2613 0.146333
R18706 GNDA.n2616 GNDA.n2517 0.146333
R18707 GNDA.n2626 GNDA.n2515 0.146333
R18708 GNDA.n2632 GNDA.n2515 0.146333
R18709 GNDA.n2633 GNDA.n2632 0.146333
R18710 GNDA.n2643 GNDA.n2642 0.146333
R18711 GNDA.n2646 GNDA.n2643 0.146333
R18712 GNDA.n2646 GNDA.n2511 0.146333
R18713 GNDA.n2819 GNDA.n2816 0.146333
R18714 GNDA.n2825 GNDA.n2816 0.146333
R18715 GNDA.n2826 GNDA.n2825 0.146333
R18716 GNDA.n2836 GNDA.n2835 0.146333
R18717 GNDA.n2839 GNDA.n2836 0.146333
R18718 GNDA.n2839 GNDA.n2812 0.146333
R18719 GNDA.n2849 GNDA.n2810 0.146333
R18720 GNDA.n2855 GNDA.n2810 0.146333
R18721 GNDA.n2856 GNDA.n2855 0.146333
R18722 GNDA.n2866 GNDA.n2865 0.146333
R18723 GNDA.n2869 GNDA.n2866 0.146333
R18724 GNDA.n2869 GNDA.n2806 0.146333
R18725 GNDA.n2879 GNDA.n2804 0.146333
R18726 GNDA.n2885 GNDA.n2804 0.146333
R18727 GNDA.n2886 GNDA.n2885 0.146333
R18728 GNDA.n2896 GNDA.n2895 0.146333
R18729 GNDA.n2899 GNDA.n2896 0.146333
R18730 GNDA.n2899 GNDA.n2800 0.146333
R18731 GNDA.n2909 GNDA.n2798 0.146333
R18732 GNDA.n2915 GNDA.n2798 0.146333
R18733 GNDA.n2916 GNDA.n2915 0.146333
R18734 GNDA.n2926 GNDA.n2925 0.146333
R18735 GNDA.n2929 GNDA.n2926 0.146333
R18736 GNDA.n2929 GNDA.n2794 0.146333
R18737 GNDA.n2960 GNDA.n2957 0.146333
R18738 GNDA.n2966 GNDA.n2957 0.146333
R18739 GNDA.n2967 GNDA.n2966 0.146333
R18740 GNDA.n2977 GNDA.n2976 0.146333
R18741 GNDA.n2980 GNDA.n2977 0.146333
R18742 GNDA.n2980 GNDA.n2953 0.146333
R18743 GNDA.n2990 GNDA.n2951 0.146333
R18744 GNDA.n2996 GNDA.n2951 0.146333
R18745 GNDA.n2997 GNDA.n2996 0.146333
R18746 GNDA.n3007 GNDA.n3006 0.146333
R18747 GNDA.n3010 GNDA.n3007 0.146333
R18748 GNDA.n3010 GNDA.n2947 0.146333
R18749 GNDA.n3020 GNDA.n2945 0.146333
R18750 GNDA.n3026 GNDA.n2945 0.146333
R18751 GNDA.n3027 GNDA.n3026 0.146333
R18752 GNDA.n3037 GNDA.n3036 0.146333
R18753 GNDA.n3040 GNDA.n3037 0.146333
R18754 GNDA.n3040 GNDA.n2941 0.146333
R18755 GNDA.n3050 GNDA.n2939 0.146333
R18756 GNDA.n3056 GNDA.n2939 0.146333
R18757 GNDA.n3057 GNDA.n3056 0.146333
R18758 GNDA.n3067 GNDA.n3066 0.146333
R18759 GNDA.n3070 GNDA.n3067 0.146333
R18760 GNDA.n3070 GNDA.n2935 0.146333
R18761 GNDA.n3101 GNDA.n3098 0.146333
R18762 GNDA.n3107 GNDA.n3098 0.146333
R18763 GNDA.n3108 GNDA.n3107 0.146333
R18764 GNDA.n3118 GNDA.n3117 0.146333
R18765 GNDA.n3121 GNDA.n3118 0.146333
R18766 GNDA.n3121 GNDA.n3094 0.146333
R18767 GNDA.n3131 GNDA.n3092 0.146333
R18768 GNDA.n3137 GNDA.n3092 0.146333
R18769 GNDA.n3138 GNDA.n3137 0.146333
R18770 GNDA.n3148 GNDA.n3147 0.146333
R18771 GNDA.n3151 GNDA.n3148 0.146333
R18772 GNDA.n3151 GNDA.n3088 0.146333
R18773 GNDA.n3161 GNDA.n3086 0.146333
R18774 GNDA.n3167 GNDA.n3086 0.146333
R18775 GNDA.n3168 GNDA.n3167 0.146333
R18776 GNDA.n3178 GNDA.n3177 0.146333
R18777 GNDA.n3181 GNDA.n3178 0.146333
R18778 GNDA.n3181 GNDA.n3082 0.146333
R18779 GNDA.n3191 GNDA.n3080 0.146333
R18780 GNDA.n3197 GNDA.n3080 0.146333
R18781 GNDA.n3198 GNDA.n3197 0.146333
R18782 GNDA.n3208 GNDA.n3207 0.146333
R18783 GNDA.n3211 GNDA.n3208 0.146333
R18784 GNDA.n3211 GNDA.n3076 0.146333
R18785 GNDA.n3286 GNDA.n3285 0.146333
R18786 GNDA.n3285 GNDA.n1896 0.146333
R18787 GNDA.n3281 GNDA.n1896 0.146333
R18788 GNDA.n3275 GNDA.n1901 0.146333
R18789 GNDA.n3275 GNDA.n3274 0.146333
R18790 GNDA.n3274 GNDA.n3273 0.146333
R18791 GNDA.n3268 GNDA.n3267 0.146333
R18792 GNDA.n3267 GNDA.n1911 0.146333
R18793 GNDA.n3263 GNDA.n1911 0.146333
R18794 GNDA.n3257 GNDA.n1916 0.146333
R18795 GNDA.n3257 GNDA.n3256 0.146333
R18796 GNDA.n3256 GNDA.n3255 0.146333
R18797 GNDA.n3250 GNDA.n3249 0.146333
R18798 GNDA.n3249 GNDA.n1926 0.146333
R18799 GNDA.n3245 GNDA.n1926 0.146333
R18800 GNDA.n3239 GNDA.n1931 0.146333
R18801 GNDA.n3239 GNDA.n3238 0.146333
R18802 GNDA.n3238 GNDA.n3237 0.146333
R18803 GNDA.n3232 GNDA.n3231 0.146333
R18804 GNDA.n3231 GNDA.n1941 0.146333
R18805 GNDA.n3227 GNDA.n1941 0.146333
R18806 GNDA.n3221 GNDA.n1946 0.146333
R18807 GNDA.n3221 GNDA.n3220 0.146333
R18808 GNDA.n3220 GNDA.n3219 0.146333
R18809 GNDA.n6356 GNDA.n6355 0.146333
R18810 GNDA.n6359 GNDA.n6356 0.146333
R18811 GNDA.n6359 GNDA.n6349 0.146333
R18812 GNDA.n6367 GNDA.n6345 0.146333
R18813 GNDA.n6371 GNDA.n6345 0.146333
R18814 GNDA.n6372 GNDA.n6371 0.146333
R18815 GNDA.n6380 GNDA.n6379 0.146333
R18816 GNDA.n6383 GNDA.n6380 0.146333
R18817 GNDA.n6383 GNDA.n6337 0.146333
R18818 GNDA.n6391 GNDA.n6333 0.146333
R18819 GNDA.n6395 GNDA.n6333 0.146333
R18820 GNDA.n6396 GNDA.n6395 0.146333
R18821 GNDA.n6404 GNDA.n6403 0.146333
R18822 GNDA.n6407 GNDA.n6404 0.146333
R18823 GNDA.n6407 GNDA.n6325 0.146333
R18824 GNDA.n6415 GNDA.n6321 0.146333
R18825 GNDA.n6419 GNDA.n6321 0.146333
R18826 GNDA.n6420 GNDA.n6419 0.146333
R18827 GNDA.n6428 GNDA.n6427 0.146333
R18828 GNDA.n6431 GNDA.n6428 0.146333
R18829 GNDA.n6431 GNDA.n6313 0.146333
R18830 GNDA.n6439 GNDA.n6311 0.146333
R18831 GNDA.n6443 GNDA.n6311 0.146333
R18832 GNDA.n6443 GNDA.n359 0.146333
R18833 GNDA.n6360 GNDA.n6352 0.146333
R18834 GNDA.n6361 GNDA.n6360 0.146333
R18835 GNDA.n6369 GNDA.n6368 0.146333
R18836 GNDA.n6370 GNDA.n6369 0.146333
R18837 GNDA.n6370 GNDA.n6344 0.146333
R18838 GNDA.n6378 GNDA.n6340 0.146333
R18839 GNDA.n6384 GNDA.n6340 0.146333
R18840 GNDA.n6385 GNDA.n6384 0.146333
R18841 GNDA.n6393 GNDA.n6392 0.146333
R18842 GNDA.n6394 GNDA.n6393 0.146333
R18843 GNDA.n6394 GNDA.n6332 0.146333
R18844 GNDA.n6402 GNDA.n6328 0.146333
R18845 GNDA.n6408 GNDA.n6328 0.146333
R18846 GNDA.n6409 GNDA.n6408 0.146333
R18847 GNDA.n6417 GNDA.n6416 0.146333
R18848 GNDA.n6418 GNDA.n6417 0.146333
R18849 GNDA.n6418 GNDA.n6320 0.146333
R18850 GNDA.n6426 GNDA.n6316 0.146333
R18851 GNDA.n6432 GNDA.n6316 0.146333
R18852 GNDA.n6433 GNDA.n6432 0.146333
R18853 GNDA.n6441 GNDA.n6440 0.146333
R18854 GNDA.n6442 GNDA.n6441 0.146333
R18855 GNDA.n6442 GNDA.n358 0.146333
R18856 GNDA.n414 GNDA.n413 0.146333
R18857 GNDA.n414 GNDA.n408 0.146333
R18858 GNDA.n424 GNDA.n406 0.146333
R18859 GNDA.n432 GNDA.n406 0.146333
R18860 GNDA.n433 GNDA.n432 0.146333
R18861 GNDA.n443 GNDA.n442 0.146333
R18862 GNDA.n444 GNDA.n443 0.146333
R18863 GNDA.n444 GNDA.n402 0.146333
R18864 GNDA.n454 GNDA.n400 0.146333
R18865 GNDA.n462 GNDA.n400 0.146333
R18866 GNDA.n463 GNDA.n462 0.146333
R18867 GNDA.n473 GNDA.n472 0.146333
R18868 GNDA.n474 GNDA.n473 0.146333
R18869 GNDA.n474 GNDA.n396 0.146333
R18870 GNDA.n484 GNDA.n394 0.146333
R18871 GNDA.n492 GNDA.n394 0.146333
R18872 GNDA.n493 GNDA.n492 0.146333
R18873 GNDA.n503 GNDA.n502 0.146333
R18874 GNDA.n504 GNDA.n503 0.146333
R18875 GNDA.n504 GNDA.n390 0.146333
R18876 GNDA.n514 GNDA.n388 0.146333
R18877 GNDA.n522 GNDA.n388 0.146333
R18878 GNDA.n523 GNDA.n522 0.146333
R18879 GNDA.n411 GNDA.n409 0.146333
R18880 GNDA.n417 GNDA.n409 0.146333
R18881 GNDA.n418 GNDA.n417 0.146333
R18882 GNDA.n428 GNDA.n427 0.146333
R18883 GNDA.n431 GNDA.n428 0.146333
R18884 GNDA.n431 GNDA.n405 0.146333
R18885 GNDA.n441 GNDA.n403 0.146333
R18886 GNDA.n447 GNDA.n403 0.146333
R18887 GNDA.n448 GNDA.n447 0.146333
R18888 GNDA.n458 GNDA.n457 0.146333
R18889 GNDA.n461 GNDA.n458 0.146333
R18890 GNDA.n461 GNDA.n399 0.146333
R18891 GNDA.n471 GNDA.n397 0.146333
R18892 GNDA.n477 GNDA.n397 0.146333
R18893 GNDA.n478 GNDA.n477 0.146333
R18894 GNDA.n488 GNDA.n487 0.146333
R18895 GNDA.n491 GNDA.n488 0.146333
R18896 GNDA.n491 GNDA.n393 0.146333
R18897 GNDA.n501 GNDA.n391 0.146333
R18898 GNDA.n507 GNDA.n391 0.146333
R18899 GNDA.n508 GNDA.n507 0.146333
R18900 GNDA.n518 GNDA.n517 0.146333
R18901 GNDA.n521 GNDA.n518 0.146333
R18902 GNDA.n521 GNDA.n387 0.146333
R18903 GNDA.n2104 GNDA.t223 0.1368
R18904 GNDA.n2103 GNDA.t362 0.1368
R18905 GNDA.n2103 GNDA.t632 0.1368
R18906 GNDA.n2102 GNDA.t245 0.1368
R18907 GNDA.n2102 GNDA.t496 0.1368
R18908 GNDA.n2101 GNDA.t384 0.1368
R18909 GNDA.n2101 GNDA.t652 0.1368
R18910 GNDA.n2100 GNDA.t552 0.1368
R18911 GNDA.n2100 GNDA.t259 0.1368
R18912 GNDA.n2099 GNDA.t401 0.1368
R18913 GNDA.n2099 GNDA.t667 0.1368
R18914 GNDA.n2098 GNDA.t575 0.1368
R18915 GNDA.n2098 GNDA.t279 0.1368
R18916 GNDA.n2097 GNDA.t705 0.1368
R18917 GNDA.n2097 GNDA.t398 0.1368
R18918 GNDA.n2096 GNDA.t571 0.1368
R18919 GNDA.n2096 GNDA.t277 0.1368
R18920 GNDA.n2095 GNDA.t726 0.1368
R18921 GNDA.n2095 GNDA.t415 0.1368
R18922 GNDA.n2094 GNDA.t321 0.1368
R18923 GNDA.n2094 GNDA.t587 0.1368
R18924 GNDA.n2093 GNDA.t493 0.1368
R18925 GNDA.n2093 GNDA.t195 0.1368
R18926 GNDA.n2092 GNDA.t337 0.1368
R18927 GNDA.n2092 GNDA.t606 0.1368
R18928 GNDA.n2091 GNDA.t512 0.1368
R18929 GNDA.n2091 GNDA.t217 0.1368
R18930 GNDA.n2090 GNDA.t666 0.1368
R18931 GNDA.n2090 GNDA.t356 0.1368
R18932 GNDA.n2089 GNDA.t528 0.1368
R18933 GNDA.n2089 GNDA.t239 0.1368
R18934 GNDA.n2088 GNDA.t687 0.1368
R18935 GNDA.n2088 GNDA.t378 0.1368
R18936 GNDA.n2087 GNDA.t298 0.1368
R18937 GNDA.n2087 GNDA.t547 0.1368
R18938 GNDA.n2086 GNDA.t704 0.1368
R18939 GNDA.n2086 GNDA.t395 0.1368
R18940 GNDA.n2085 GNDA.t459 0.1368
R18941 GNDA.n2085 GNDA.t566 0.1368
R18942 GNDA.n2084 GNDA.t481 0.1368
R18943 GNDA.n2084 GNDA.t724 0.1368
R18944 GNDA.n2083 GNDA.t603 0.1368
R18945 GNDA.n2083 GNDA.t454 0.1368
R18946 GNDA.n2082 GNDA.t478 0.1368
R18947 GNDA.n2082 GNDA.t720 0.1368
R18948 GNDA.n2081 GNDA.t629 0.1368
R18949 GNDA.n2081 GNDA.t315 0.1368
R18950 GNDA.n2080 GNDA.t238 0.1368
R18951 GNDA.n2080 GNDA.t488 0.1368
R18952 GNDA.n2079 GNDA.t647 0.1368
R18953 GNDA.n2079 GNDA.t334 0.1368
R18954 GNDA.n2078 GNDA.t256 0.1368
R18955 GNDA.n2078 GNDA.t506 0.1368
R18956 GNDA.n2077 GNDA.t394 0.1368
R18957 GNDA.n2077 GNDA.t662 0.1368
R18958 GNDA.n2076 GNDA.t275 0.1368
R18959 GNDA.n2076 GNDA.t523 0.1368
R18960 GNDA.n2075 GNDA.t414 0.1368
R18961 GNDA.n2075 GNDA.t678 0.1368
R18962 GNDA.n2074 GNDA.t586 0.1368
R18963 GNDA.n2074 GNDA.t291 0.1368
R18964 GNDA.n2073 GNDA.t194 0.1368
R18965 GNDA.n2073 GNDA.t429 0.1368
R18966 GNDA.t482 GNDA.n2104 0.1368
R18967 GNDA.n2228 GNDA.t685 0.1368
R18968 GNDA.n4777 GNDA.n1597 0.135917
R18969 GNDA.n4671 GNDA.n4668 0.135917
R18970 GNDA.n4677 GNDA.n4660 0.135917
R18971 GNDA.n4687 GNDA.n4658 0.135917
R18972 GNDA.n4691 GNDA.n4688 0.135917
R18973 GNDA.n4701 GNDA.n4698 0.135917
R18974 GNDA.n4707 GNDA.n4654 0.135917
R18975 GNDA.n4717 GNDA.n4652 0.135917
R18976 GNDA.n4721 GNDA.n4718 0.135917
R18977 GNDA.n4731 GNDA.n4728 0.135917
R18978 GNDA.n4737 GNDA.n4648 0.135917
R18979 GNDA.n4747 GNDA.n4646 0.135917
R18980 GNDA.n4751 GNDA.n4748 0.135917
R18981 GNDA.n4761 GNDA.n4758 0.135917
R18982 GNDA.n4767 GNDA.n4642 0.135917
R18983 GNDA.n5688 GNDA.n5686 0.135917
R18984 GNDA.n5698 GNDA.n5695 0.135917
R18985 GNDA.n5704 GNDA.n5683 0.135917
R18986 GNDA.n5714 GNDA.n5681 0.135917
R18987 GNDA.n5718 GNDA.n5715 0.135917
R18988 GNDA.n5728 GNDA.n5725 0.135917
R18989 GNDA.n5734 GNDA.n5677 0.135917
R18990 GNDA.n5744 GNDA.n5675 0.135917
R18991 GNDA.n5748 GNDA.n5745 0.135917
R18992 GNDA.n5758 GNDA.n5755 0.135917
R18993 GNDA.n5764 GNDA.n5671 0.135917
R18994 GNDA.n5774 GNDA.n5669 0.135917
R18995 GNDA.n5778 GNDA.n5775 0.135917
R18996 GNDA.n5788 GNDA.n5785 0.135917
R18997 GNDA.n5794 GNDA.n5665 0.135917
R18998 GNDA.n2700 GNDA.n2698 0.135917
R18999 GNDA.n2708 GNDA.n2705 0.135917
R19000 GNDA.n2712 GNDA.n2690 0.135917
R19001 GNDA.n2720 GNDA.n2686 0.135917
R19002 GNDA.n2724 GNDA.n2721 0.135917
R19003 GNDA.n2732 GNDA.n2729 0.135917
R19004 GNDA.n2736 GNDA.n2678 0.135917
R19005 GNDA.n2744 GNDA.n2674 0.135917
R19006 GNDA.n2748 GNDA.n2745 0.135917
R19007 GNDA.n2756 GNDA.n2753 0.135917
R19008 GNDA.n2760 GNDA.n2666 0.135917
R19009 GNDA.n2768 GNDA.n2662 0.135917
R19010 GNDA.n2772 GNDA.n2769 0.135917
R19011 GNDA.n2780 GNDA.n2777 0.135917
R19012 GNDA.n2784 GNDA.n2654 0.135917
R19013 GNDA.n6082 GNDA.n1369 0.135917
R19014 GNDA.n5976 GNDA.n5973 0.135917
R19015 GNDA.n5982 GNDA.n5965 0.135917
R19016 GNDA.n5992 GNDA.n5963 0.135917
R19017 GNDA.n5996 GNDA.n5993 0.135917
R19018 GNDA.n6006 GNDA.n6003 0.135917
R19019 GNDA.n6012 GNDA.n5959 0.135917
R19020 GNDA.n6022 GNDA.n5957 0.135917
R19021 GNDA.n6026 GNDA.n6023 0.135917
R19022 GNDA.n6036 GNDA.n6033 0.135917
R19023 GNDA.n6042 GNDA.n5953 0.135917
R19024 GNDA.n6052 GNDA.n5951 0.135917
R19025 GNDA.n6056 GNDA.n6053 0.135917
R19026 GNDA.n6066 GNDA.n6063 0.135917
R19027 GNDA.n6072 GNDA.n5947 0.135917
R19028 GNDA.n1586 GNDA.n1424 0.135917
R19029 GNDA.n1428 GNDA.n1427 0.135917
R19030 GNDA.n1430 GNDA.n1429 0.135917
R19031 GNDA.n1434 GNDA.n1433 0.135917
R19032 GNDA.n1436 GNDA.n1435 0.135917
R19033 GNDA.n1440 GNDA.n1439 0.135917
R19034 GNDA.n1442 GNDA.n1441 0.135917
R19035 GNDA.n1446 GNDA.n1445 0.135917
R19036 GNDA.n1448 GNDA.n1447 0.135917
R19037 GNDA.n1452 GNDA.n1451 0.135917
R19038 GNDA.n1454 GNDA.n1453 0.135917
R19039 GNDA.n1458 GNDA.n1457 0.135917
R19040 GNDA.n1460 GNDA.n1459 0.135917
R19041 GNDA.n1464 GNDA.n1463 0.135917
R19042 GNDA.n1466 GNDA.n1465 0.135917
R19043 GNDA.n3637 GNDA.n3635 0.135917
R19044 GNDA.n3647 GNDA.n3644 0.135917
R19045 GNDA.n3653 GNDA.n3631 0.135917
R19046 GNDA.n3663 GNDA.n3629 0.135917
R19047 GNDA.n3667 GNDA.n3664 0.135917
R19048 GNDA.n3677 GNDA.n3674 0.135917
R19049 GNDA.n3683 GNDA.n3625 0.135917
R19050 GNDA.n3693 GNDA.n3623 0.135917
R19051 GNDA.n3697 GNDA.n3694 0.135917
R19052 GNDA.n3707 GNDA.n3704 0.135917
R19053 GNDA.n3713 GNDA.n3619 0.135917
R19054 GNDA.n3723 GNDA.n3617 0.135917
R19055 GNDA.n3727 GNDA.n3724 0.135917
R19056 GNDA.n3737 GNDA.n3734 0.135917
R19057 GNDA.n3743 GNDA.n3613 0.135917
R19058 GNDA.n3458 GNDA.n3296 0.135917
R19059 GNDA.n3300 GNDA.n3299 0.135917
R19060 GNDA.n3302 GNDA.n3301 0.135917
R19061 GNDA.n3306 GNDA.n3305 0.135917
R19062 GNDA.n3308 GNDA.n3307 0.135917
R19063 GNDA.n3312 GNDA.n3311 0.135917
R19064 GNDA.n3314 GNDA.n3313 0.135917
R19065 GNDA.n3318 GNDA.n3317 0.135917
R19066 GNDA.n3320 GNDA.n3319 0.135917
R19067 GNDA.n3324 GNDA.n3323 0.135917
R19068 GNDA.n3326 GNDA.n3325 0.135917
R19069 GNDA.n3330 GNDA.n3329 0.135917
R19070 GNDA.n3332 GNDA.n3331 0.135917
R19071 GNDA.n3336 GNDA.n3335 0.135917
R19072 GNDA.n3338 GNDA.n3337 0.135917
R19073 GNDA.n5233 GNDA.n5070 0.135917
R19074 GNDA.n5127 GNDA.n5124 0.135917
R19075 GNDA.n5133 GNDA.n5116 0.135917
R19076 GNDA.n5143 GNDA.n5114 0.135917
R19077 GNDA.n5147 GNDA.n5144 0.135917
R19078 GNDA.n5157 GNDA.n5154 0.135917
R19079 GNDA.n5163 GNDA.n5110 0.135917
R19080 GNDA.n5173 GNDA.n5108 0.135917
R19081 GNDA.n5177 GNDA.n5174 0.135917
R19082 GNDA.n5187 GNDA.n5184 0.135917
R19083 GNDA.n5193 GNDA.n5104 0.135917
R19084 GNDA.n5203 GNDA.n5102 0.135917
R19085 GNDA.n5207 GNDA.n5204 0.135917
R19086 GNDA.n5217 GNDA.n5214 0.135917
R19087 GNDA.n5223 GNDA.n5098 0.135917
R19088 GNDA.n5398 GNDA.n5236 0.135917
R19089 GNDA.n5240 GNDA.n5239 0.135917
R19090 GNDA.n5242 GNDA.n5241 0.135917
R19091 GNDA.n5246 GNDA.n5245 0.135917
R19092 GNDA.n5248 GNDA.n5247 0.135917
R19093 GNDA.n5252 GNDA.n5251 0.135917
R19094 GNDA.n5254 GNDA.n5253 0.135917
R19095 GNDA.n5258 GNDA.n5257 0.135917
R19096 GNDA.n5260 GNDA.n5259 0.135917
R19097 GNDA.n5264 GNDA.n5263 0.135917
R19098 GNDA.n5266 GNDA.n5265 0.135917
R19099 GNDA.n5270 GNDA.n5269 0.135917
R19100 GNDA.n5272 GNDA.n5271 0.135917
R19101 GNDA.n5276 GNDA.n5275 0.135917
R19102 GNDA.n5278 GNDA.n5277 0.135917
R19103 GNDA.n5405 GNDA.n5403 0.135917
R19104 GNDA.n5415 GNDA.n5412 0.135917
R19105 GNDA.n5421 GNDA.n5066 0.135917
R19106 GNDA.n5431 GNDA.n5064 0.135917
R19107 GNDA.n5435 GNDA.n5432 0.135917
R19108 GNDA.n5445 GNDA.n5442 0.135917
R19109 GNDA.n5451 GNDA.n5060 0.135917
R19110 GNDA.n5461 GNDA.n5058 0.135917
R19111 GNDA.n5465 GNDA.n5462 0.135917
R19112 GNDA.n5475 GNDA.n5472 0.135917
R19113 GNDA.n5481 GNDA.n5054 0.135917
R19114 GNDA.n5491 GNDA.n5052 0.135917
R19115 GNDA.n5495 GNDA.n5492 0.135917
R19116 GNDA.n5505 GNDA.n5502 0.135917
R19117 GNDA.n5511 GNDA.n5048 0.135917
R19118 GNDA.n5547 GNDA.n5545 0.135917
R19119 GNDA.n5557 GNDA.n5554 0.135917
R19120 GNDA.n5563 GNDA.n5541 0.135917
R19121 GNDA.n5573 GNDA.n5539 0.135917
R19122 GNDA.n5577 GNDA.n5574 0.135917
R19123 GNDA.n5587 GNDA.n5584 0.135917
R19124 GNDA.n5593 GNDA.n5535 0.135917
R19125 GNDA.n5603 GNDA.n5533 0.135917
R19126 GNDA.n5607 GNDA.n5604 0.135917
R19127 GNDA.n5617 GNDA.n5614 0.135917
R19128 GNDA.n5623 GNDA.n5529 0.135917
R19129 GNDA.n5633 GNDA.n5527 0.135917
R19130 GNDA.n5637 GNDA.n5634 0.135917
R19131 GNDA.n5647 GNDA.n5644 0.135917
R19132 GNDA.n5653 GNDA.n5523 0.135917
R19133 GNDA.n5829 GNDA.n5827 0.135917
R19134 GNDA.n5839 GNDA.n5836 0.135917
R19135 GNDA.n5845 GNDA.n5824 0.135917
R19136 GNDA.n5855 GNDA.n5822 0.135917
R19137 GNDA.n5859 GNDA.n5856 0.135917
R19138 GNDA.n5869 GNDA.n5866 0.135917
R19139 GNDA.n5875 GNDA.n5818 0.135917
R19140 GNDA.n5885 GNDA.n5816 0.135917
R19141 GNDA.n5889 GNDA.n5886 0.135917
R19142 GNDA.n5899 GNDA.n5896 0.135917
R19143 GNDA.n5905 GNDA.n5812 0.135917
R19144 GNDA.n5915 GNDA.n5810 0.135917
R19145 GNDA.n5919 GNDA.n5916 0.135917
R19146 GNDA.n5929 GNDA.n5926 0.135917
R19147 GNDA.n5935 GNDA.n5806 0.135917
R19148 GNDA.n4810 GNDA.n4808 0.135917
R19149 GNDA.n4820 GNDA.n4817 0.135917
R19150 GNDA.n4826 GNDA.n1417 0.135917
R19151 GNDA.n4836 GNDA.n1415 0.135917
R19152 GNDA.n4840 GNDA.n4837 0.135917
R19153 GNDA.n4850 GNDA.n4847 0.135917
R19154 GNDA.n4856 GNDA.n1411 0.135917
R19155 GNDA.n4866 GNDA.n1409 0.135917
R19156 GNDA.n4870 GNDA.n4867 0.135917
R19157 GNDA.n4880 GNDA.n4877 0.135917
R19158 GNDA.n4886 GNDA.n1405 0.135917
R19159 GNDA.n4896 GNDA.n1403 0.135917
R19160 GNDA.n4900 GNDA.n4897 0.135917
R19161 GNDA.n4910 GNDA.n4907 0.135917
R19162 GNDA.n4916 GNDA.n1399 0.135917
R19163 GNDA.n4524 GNDA.n4522 0.135917
R19164 GNDA.n4534 GNDA.n4531 0.135917
R19165 GNDA.n4540 GNDA.n4518 0.135917
R19166 GNDA.n4550 GNDA.n4516 0.135917
R19167 GNDA.n4554 GNDA.n4551 0.135917
R19168 GNDA.n4564 GNDA.n4561 0.135917
R19169 GNDA.n4570 GNDA.n4512 0.135917
R19170 GNDA.n4580 GNDA.n4510 0.135917
R19171 GNDA.n4584 GNDA.n4581 0.135917
R19172 GNDA.n4594 GNDA.n4591 0.135917
R19173 GNDA.n4600 GNDA.n4506 0.135917
R19174 GNDA.n4610 GNDA.n4504 0.135917
R19175 GNDA.n4614 GNDA.n4611 0.135917
R19176 GNDA.n4624 GNDA.n4621 0.135917
R19177 GNDA.n4630 GNDA.n4500 0.135917
R19178 GNDA.n4335 GNDA.n4333 0.135917
R19179 GNDA.n4345 GNDA.n4342 0.135917
R19180 GNDA.n4351 GNDA.n4329 0.135917
R19181 GNDA.n4361 GNDA.n4327 0.135917
R19182 GNDA.n4365 GNDA.n4362 0.135917
R19183 GNDA.n4375 GNDA.n4372 0.135917
R19184 GNDA.n4381 GNDA.n4323 0.135917
R19185 GNDA.n4391 GNDA.n4321 0.135917
R19186 GNDA.n4395 GNDA.n4392 0.135917
R19187 GNDA.n4405 GNDA.n4402 0.135917
R19188 GNDA.n4411 GNDA.n4317 0.135917
R19189 GNDA.n4421 GNDA.n4315 0.135917
R19190 GNDA.n4425 GNDA.n4422 0.135917
R19191 GNDA.n4435 GNDA.n4432 0.135917
R19192 GNDA.n4441 GNDA.n4311 0.135917
R19193 GNDA.n4169 GNDA.n4167 0.135917
R19194 GNDA.n4179 GNDA.n4176 0.135917
R19195 GNDA.n4185 GNDA.n1645 0.135917
R19196 GNDA.n4195 GNDA.n1643 0.135917
R19197 GNDA.n4199 GNDA.n4196 0.135917
R19198 GNDA.n4209 GNDA.n4206 0.135917
R19199 GNDA.n4215 GNDA.n1639 0.135917
R19200 GNDA.n4225 GNDA.n1637 0.135917
R19201 GNDA.n4229 GNDA.n4226 0.135917
R19202 GNDA.n4239 GNDA.n4236 0.135917
R19203 GNDA.n4245 GNDA.n1633 0.135917
R19204 GNDA.n4255 GNDA.n1631 0.135917
R19205 GNDA.n4259 GNDA.n4256 0.135917
R19206 GNDA.n4269 GNDA.n4266 0.135917
R19207 GNDA.n4275 GNDA.n1627 0.135917
R19208 GNDA.n1812 GNDA.n1650 0.135917
R19209 GNDA.n1654 GNDA.n1653 0.135917
R19210 GNDA.n1656 GNDA.n1655 0.135917
R19211 GNDA.n1660 GNDA.n1659 0.135917
R19212 GNDA.n1662 GNDA.n1661 0.135917
R19213 GNDA.n1666 GNDA.n1665 0.135917
R19214 GNDA.n1668 GNDA.n1667 0.135917
R19215 GNDA.n1672 GNDA.n1671 0.135917
R19216 GNDA.n1674 GNDA.n1673 0.135917
R19217 GNDA.n1678 GNDA.n1677 0.135917
R19218 GNDA.n1680 GNDA.n1679 0.135917
R19219 GNDA.n1684 GNDA.n1683 0.135917
R19220 GNDA.n1686 GNDA.n1685 0.135917
R19221 GNDA.n1690 GNDA.n1689 0.135917
R19222 GNDA.n1692 GNDA.n1691 0.135917
R19223 GNDA.n3826 GNDA.n3824 0.135917
R19224 GNDA.n3836 GNDA.n3833 0.135917
R19225 GNDA.n3842 GNDA.n3820 0.135917
R19226 GNDA.n3852 GNDA.n3818 0.135917
R19227 GNDA.n3856 GNDA.n3853 0.135917
R19228 GNDA.n3866 GNDA.n3863 0.135917
R19229 GNDA.n3872 GNDA.n3814 0.135917
R19230 GNDA.n3882 GNDA.n3812 0.135917
R19231 GNDA.n3886 GNDA.n3883 0.135917
R19232 GNDA.n3896 GNDA.n3893 0.135917
R19233 GNDA.n3902 GNDA.n3808 0.135917
R19234 GNDA.n3912 GNDA.n3806 0.135917
R19235 GNDA.n3916 GNDA.n3913 0.135917
R19236 GNDA.n3926 GNDA.n3923 0.135917
R19237 GNDA.n3932 GNDA.n3802 0.135917
R19238 GNDA.n4079 GNDA.n1836 0.135917
R19239 GNDA.n3973 GNDA.n3970 0.135917
R19240 GNDA.n3979 GNDA.n3962 0.135917
R19241 GNDA.n3989 GNDA.n3960 0.135917
R19242 GNDA.n3993 GNDA.n3990 0.135917
R19243 GNDA.n4003 GNDA.n4000 0.135917
R19244 GNDA.n4009 GNDA.n3956 0.135917
R19245 GNDA.n4019 GNDA.n3954 0.135917
R19246 GNDA.n4023 GNDA.n4020 0.135917
R19247 GNDA.n4033 GNDA.n4030 0.135917
R19248 GNDA.n4039 GNDA.n3950 0.135917
R19249 GNDA.n4049 GNDA.n3948 0.135917
R19250 GNDA.n4053 GNDA.n4050 0.135917
R19251 GNDA.n4063 GNDA.n4060 0.135917
R19252 GNDA.n4069 GNDA.n3944 0.135917
R19253 GNDA.n3471 GNDA.n3469 0.135917
R19254 GNDA.n3481 GNDA.n3478 0.135917
R19255 GNDA.n3487 GNDA.n1884 0.135917
R19256 GNDA.n3497 GNDA.n1882 0.135917
R19257 GNDA.n3501 GNDA.n3498 0.135917
R19258 GNDA.n3511 GNDA.n3508 0.135917
R19259 GNDA.n3517 GNDA.n1878 0.135917
R19260 GNDA.n3527 GNDA.n1876 0.135917
R19261 GNDA.n3531 GNDA.n3528 0.135917
R19262 GNDA.n3541 GNDA.n3538 0.135917
R19263 GNDA.n3547 GNDA.n1872 0.135917
R19264 GNDA.n3557 GNDA.n1870 0.135917
R19265 GNDA.n3561 GNDA.n3558 0.135917
R19266 GNDA.n3571 GNDA.n3568 0.135917
R19267 GNDA.n3577 GNDA.n1866 0.135917
R19268 GNDA.n2536 GNDA.n2534 0.135917
R19269 GNDA.n2546 GNDA.n2543 0.135917
R19270 GNDA.n2552 GNDA.n2531 0.135917
R19271 GNDA.n2562 GNDA.n2529 0.135917
R19272 GNDA.n2566 GNDA.n2563 0.135917
R19273 GNDA.n2576 GNDA.n2573 0.135917
R19274 GNDA.n2582 GNDA.n2525 0.135917
R19275 GNDA.n2592 GNDA.n2523 0.135917
R19276 GNDA.n2596 GNDA.n2593 0.135917
R19277 GNDA.n2606 GNDA.n2603 0.135917
R19278 GNDA.n2612 GNDA.n2519 0.135917
R19279 GNDA.n2622 GNDA.n2517 0.135917
R19280 GNDA.n2626 GNDA.n2623 0.135917
R19281 GNDA.n2636 GNDA.n2633 0.135917
R19282 GNDA.n2642 GNDA.n2513 0.135917
R19283 GNDA.n2819 GNDA.n2817 0.135917
R19284 GNDA.n2829 GNDA.n2826 0.135917
R19285 GNDA.n2835 GNDA.n2814 0.135917
R19286 GNDA.n2845 GNDA.n2812 0.135917
R19287 GNDA.n2849 GNDA.n2846 0.135917
R19288 GNDA.n2859 GNDA.n2856 0.135917
R19289 GNDA.n2865 GNDA.n2808 0.135917
R19290 GNDA.n2875 GNDA.n2806 0.135917
R19291 GNDA.n2879 GNDA.n2876 0.135917
R19292 GNDA.n2889 GNDA.n2886 0.135917
R19293 GNDA.n2895 GNDA.n2802 0.135917
R19294 GNDA.n2905 GNDA.n2800 0.135917
R19295 GNDA.n2909 GNDA.n2906 0.135917
R19296 GNDA.n2919 GNDA.n2916 0.135917
R19297 GNDA.n2925 GNDA.n2796 0.135917
R19298 GNDA.n2960 GNDA.n2958 0.135917
R19299 GNDA.n2970 GNDA.n2967 0.135917
R19300 GNDA.n2976 GNDA.n2955 0.135917
R19301 GNDA.n2986 GNDA.n2953 0.135917
R19302 GNDA.n2990 GNDA.n2987 0.135917
R19303 GNDA.n3000 GNDA.n2997 0.135917
R19304 GNDA.n3006 GNDA.n2949 0.135917
R19305 GNDA.n3016 GNDA.n2947 0.135917
R19306 GNDA.n3020 GNDA.n3017 0.135917
R19307 GNDA.n3030 GNDA.n3027 0.135917
R19308 GNDA.n3036 GNDA.n2943 0.135917
R19309 GNDA.n3046 GNDA.n2941 0.135917
R19310 GNDA.n3050 GNDA.n3047 0.135917
R19311 GNDA.n3060 GNDA.n3057 0.135917
R19312 GNDA.n3066 GNDA.n2937 0.135917
R19313 GNDA.n3101 GNDA.n3099 0.135917
R19314 GNDA.n3111 GNDA.n3108 0.135917
R19315 GNDA.n3117 GNDA.n3096 0.135917
R19316 GNDA.n3127 GNDA.n3094 0.135917
R19317 GNDA.n3131 GNDA.n3128 0.135917
R19318 GNDA.n3141 GNDA.n3138 0.135917
R19319 GNDA.n3147 GNDA.n3090 0.135917
R19320 GNDA.n3157 GNDA.n3088 0.135917
R19321 GNDA.n3161 GNDA.n3158 0.135917
R19322 GNDA.n3171 GNDA.n3168 0.135917
R19323 GNDA.n3177 GNDA.n3084 0.135917
R19324 GNDA.n3187 GNDA.n3082 0.135917
R19325 GNDA.n3191 GNDA.n3188 0.135917
R19326 GNDA.n3201 GNDA.n3198 0.135917
R19327 GNDA.n3207 GNDA.n3078 0.135917
R19328 GNDA.n3287 GNDA.n3286 0.135917
R19329 GNDA.n3281 GNDA.n3280 0.135917
R19330 GNDA.n3279 GNDA.n1901 0.135917
R19331 GNDA.n3273 GNDA.n1906 0.135917
R19332 GNDA.n3269 GNDA.n3268 0.135917
R19333 GNDA.n3263 GNDA.n3262 0.135917
R19334 GNDA.n3261 GNDA.n1916 0.135917
R19335 GNDA.n3255 GNDA.n1921 0.135917
R19336 GNDA.n3251 GNDA.n3250 0.135917
R19337 GNDA.n3245 GNDA.n3244 0.135917
R19338 GNDA.n3243 GNDA.n1931 0.135917
R19339 GNDA.n3237 GNDA.n1936 0.135917
R19340 GNDA.n3233 GNDA.n3232 0.135917
R19341 GNDA.n3227 GNDA.n3226 0.135917
R19342 GNDA.n3225 GNDA.n1946 0.135917
R19343 GNDA.n6363 GNDA.n6349 0.135917
R19344 GNDA.n6367 GNDA.n6364 0.135917
R19345 GNDA.n6375 GNDA.n6372 0.135917
R19346 GNDA.n6379 GNDA.n6341 0.135917
R19347 GNDA.n6387 GNDA.n6337 0.135917
R19348 GNDA.n6391 GNDA.n6388 0.135917
R19349 GNDA.n6399 GNDA.n6396 0.135917
R19350 GNDA.n6403 GNDA.n6329 0.135917
R19351 GNDA.n6411 GNDA.n6325 0.135917
R19352 GNDA.n6415 GNDA.n6412 0.135917
R19353 GNDA.n6423 GNDA.n6420 0.135917
R19354 GNDA.n6427 GNDA.n6317 0.135917
R19355 GNDA.n6435 GNDA.n6313 0.135917
R19356 GNDA.n6439 GNDA.n6436 0.135917
R19357 GNDA.n6617 GNDA.n359 0.135917
R19358 GNDA.n6362 GNDA.n6361 0.135917
R19359 GNDA.n6368 GNDA.n6348 0.135917
R19360 GNDA.n6376 GNDA.n6344 0.135917
R19361 GNDA.n6378 GNDA.n6377 0.135917
R19362 GNDA.n6386 GNDA.n6385 0.135917
R19363 GNDA.n6392 GNDA.n6336 0.135917
R19364 GNDA.n6400 GNDA.n6332 0.135917
R19365 GNDA.n6402 GNDA.n6401 0.135917
R19366 GNDA.n6410 GNDA.n6409 0.135917
R19367 GNDA.n6416 GNDA.n6324 0.135917
R19368 GNDA.n6424 GNDA.n6320 0.135917
R19369 GNDA.n6426 GNDA.n6425 0.135917
R19370 GNDA.n6434 GNDA.n6433 0.135917
R19371 GNDA.n6440 GNDA.n6312 0.135917
R19372 GNDA.n6618 GNDA.n358 0.135917
R19373 GNDA.n422 GNDA.n408 0.135917
R19374 GNDA.n424 GNDA.n423 0.135917
R19375 GNDA.n434 GNDA.n433 0.135917
R19376 GNDA.n442 GNDA.n404 0.135917
R19377 GNDA.n452 GNDA.n402 0.135917
R19378 GNDA.n454 GNDA.n453 0.135917
R19379 GNDA.n464 GNDA.n463 0.135917
R19380 GNDA.n472 GNDA.n398 0.135917
R19381 GNDA.n482 GNDA.n396 0.135917
R19382 GNDA.n484 GNDA.n483 0.135917
R19383 GNDA.n494 GNDA.n493 0.135917
R19384 GNDA.n502 GNDA.n392 0.135917
R19385 GNDA.n512 GNDA.n390 0.135917
R19386 GNDA.n514 GNDA.n513 0.135917
R19387 GNDA.n6283 GNDA.n523 0.135917
R19388 GNDA.n421 GNDA.n418 0.135917
R19389 GNDA.n427 GNDA.n407 0.135917
R19390 GNDA.n437 GNDA.n405 0.135917
R19391 GNDA.n441 GNDA.n438 0.135917
R19392 GNDA.n451 GNDA.n448 0.135917
R19393 GNDA.n457 GNDA.n401 0.135917
R19394 GNDA.n467 GNDA.n399 0.135917
R19395 GNDA.n471 GNDA.n468 0.135917
R19396 GNDA.n481 GNDA.n478 0.135917
R19397 GNDA.n487 GNDA.n395 0.135917
R19398 GNDA.n497 GNDA.n393 0.135917
R19399 GNDA.n501 GNDA.n498 0.135917
R19400 GNDA.n511 GNDA.n508 0.135917
R19401 GNDA.n517 GNDA.n389 0.135917
R19402 GNDA.n6284 GNDA.n387 0.135917
R19403 GNDA.n4671 GNDA.n4660 0.1255
R19404 GNDA.n4688 GNDA.n4687 0.1255
R19405 GNDA.n4701 GNDA.n4654 0.1255
R19406 GNDA.n4718 GNDA.n4717 0.1255
R19407 GNDA.n4731 GNDA.n4648 0.1255
R19408 GNDA.n4748 GNDA.n4747 0.1255
R19409 GNDA.n4761 GNDA.n4642 0.1255
R19410 GNDA.n5698 GNDA.n5683 0.1255
R19411 GNDA.n5715 GNDA.n5714 0.1255
R19412 GNDA.n5728 GNDA.n5677 0.1255
R19413 GNDA.n5745 GNDA.n5744 0.1255
R19414 GNDA.n5758 GNDA.n5671 0.1255
R19415 GNDA.n5775 GNDA.n5774 0.1255
R19416 GNDA.n5788 GNDA.n5665 0.1255
R19417 GNDA.n2708 GNDA.n2690 0.1255
R19418 GNDA.n2721 GNDA.n2720 0.1255
R19419 GNDA.n2732 GNDA.n2678 0.1255
R19420 GNDA.n2745 GNDA.n2744 0.1255
R19421 GNDA.n2756 GNDA.n2666 0.1255
R19422 GNDA.n2769 GNDA.n2768 0.1255
R19423 GNDA.n2780 GNDA.n2654 0.1255
R19424 GNDA.n6084 GNDA.n1367 0.1255
R19425 GNDA.n5976 GNDA.n5965 0.1255
R19426 GNDA.n5993 GNDA.n5992 0.1255
R19427 GNDA.n6006 GNDA.n5959 0.1255
R19428 GNDA.n6023 GNDA.n6022 0.1255
R19429 GNDA.n6036 GNDA.n5953 0.1255
R19430 GNDA.n6053 GNDA.n6052 0.1255
R19431 GNDA.n6066 GNDA.n5947 0.1255
R19432 GNDA.n4802 GNDA.n1588 0.1255
R19433 GNDA.n1429 GNDA.n1428 0.1255
R19434 GNDA.n1435 GNDA.n1434 0.1255
R19435 GNDA.n1441 GNDA.n1440 0.1255
R19436 GNDA.n1447 GNDA.n1446 0.1255
R19437 GNDA.n1453 GNDA.n1452 0.1255
R19438 GNDA.n1459 GNDA.n1458 0.1255
R19439 GNDA.n1465 GNDA.n1464 0.1255
R19440 GNDA.n4084 GNDA.n1832 0.1255
R19441 GNDA.n3647 GNDA.n3631 0.1255
R19442 GNDA.n3664 GNDA.n3663 0.1255
R19443 GNDA.n3677 GNDA.n3625 0.1255
R19444 GNDA.n3694 GNDA.n3693 0.1255
R19445 GNDA.n3707 GNDA.n3619 0.1255
R19446 GNDA.n3724 GNDA.n3723 0.1255
R19447 GNDA.n3737 GNDA.n3613 0.1255
R19448 GNDA.n3463 GNDA.n3460 0.1255
R19449 GNDA.n3301 GNDA.n3300 0.1255
R19450 GNDA.n3307 GNDA.n3306 0.1255
R19451 GNDA.n3313 GNDA.n3312 0.1255
R19452 GNDA.n3319 GNDA.n3318 0.1255
R19453 GNDA.n3325 GNDA.n3324 0.1255
R19454 GNDA.n3331 GNDA.n3330 0.1255
R19455 GNDA.n3337 GNDA.n3336 0.1255
R19456 GNDA.n5127 GNDA.n5116 0.1255
R19457 GNDA.n5144 GNDA.n5143 0.1255
R19458 GNDA.n5157 GNDA.n5110 0.1255
R19459 GNDA.n5174 GNDA.n5173 0.1255
R19460 GNDA.n5187 GNDA.n5104 0.1255
R19461 GNDA.n5204 GNDA.n5203 0.1255
R19462 GNDA.n5217 GNDA.n5098 0.1255
R19463 GNDA.n5241 GNDA.n5240 0.1255
R19464 GNDA.n5247 GNDA.n5246 0.1255
R19465 GNDA.n5253 GNDA.n5252 0.1255
R19466 GNDA.n5259 GNDA.n5258 0.1255
R19467 GNDA.n5265 GNDA.n5264 0.1255
R19468 GNDA.n5271 GNDA.n5270 0.1255
R19469 GNDA.n5277 GNDA.n5276 0.1255
R19470 GNDA.n5415 GNDA.n5066 0.1255
R19471 GNDA.n5432 GNDA.n5431 0.1255
R19472 GNDA.n5445 GNDA.n5060 0.1255
R19473 GNDA.n5462 GNDA.n5461 0.1255
R19474 GNDA.n5475 GNDA.n5054 0.1255
R19475 GNDA.n5492 GNDA.n5491 0.1255
R19476 GNDA.n5505 GNDA.n5048 0.1255
R19477 GNDA.n5557 GNDA.n5541 0.1255
R19478 GNDA.n5574 GNDA.n5573 0.1255
R19479 GNDA.n5587 GNDA.n5535 0.1255
R19480 GNDA.n5604 GNDA.n5603 0.1255
R19481 GNDA.n5617 GNDA.n5529 0.1255
R19482 GNDA.n5634 GNDA.n5633 0.1255
R19483 GNDA.n5647 GNDA.n5523 0.1255
R19484 GNDA.n5839 GNDA.n5824 0.1255
R19485 GNDA.n5856 GNDA.n5855 0.1255
R19486 GNDA.n5869 GNDA.n5818 0.1255
R19487 GNDA.n5886 GNDA.n5885 0.1255
R19488 GNDA.n5899 GNDA.n5812 0.1255
R19489 GNDA.n5916 GNDA.n5915 0.1255
R19490 GNDA.n5929 GNDA.n5806 0.1255
R19491 GNDA.n4820 GNDA.n1417 0.1255
R19492 GNDA.n4837 GNDA.n4836 0.1255
R19493 GNDA.n4850 GNDA.n1411 0.1255
R19494 GNDA.n4867 GNDA.n4866 0.1255
R19495 GNDA.n4880 GNDA.n1405 0.1255
R19496 GNDA.n4897 GNDA.n4896 0.1255
R19497 GNDA.n4910 GNDA.n1399 0.1255
R19498 GNDA.n4534 GNDA.n4518 0.1255
R19499 GNDA.n4551 GNDA.n4550 0.1255
R19500 GNDA.n4564 GNDA.n4512 0.1255
R19501 GNDA.n4581 GNDA.n4580 0.1255
R19502 GNDA.n4594 GNDA.n4506 0.1255
R19503 GNDA.n4611 GNDA.n4610 0.1255
R19504 GNDA.n4624 GNDA.n4500 0.1255
R19505 GNDA.n4345 GNDA.n4329 0.1255
R19506 GNDA.n4362 GNDA.n4361 0.1255
R19507 GNDA.n4375 GNDA.n4323 0.1255
R19508 GNDA.n4392 GNDA.n4391 0.1255
R19509 GNDA.n4405 GNDA.n4317 0.1255
R19510 GNDA.n4422 GNDA.n4421 0.1255
R19511 GNDA.n4435 GNDA.n4311 0.1255
R19512 GNDA.n4179 GNDA.n1645 0.1255
R19513 GNDA.n4196 GNDA.n4195 0.1255
R19514 GNDA.n4209 GNDA.n1639 0.1255
R19515 GNDA.n4226 GNDA.n4225 0.1255
R19516 GNDA.n4239 GNDA.n1633 0.1255
R19517 GNDA.n4256 GNDA.n4255 0.1255
R19518 GNDA.n4269 GNDA.n1627 0.1255
R19519 GNDA.n1655 GNDA.n1654 0.1255
R19520 GNDA.n1661 GNDA.n1660 0.1255
R19521 GNDA.n1667 GNDA.n1666 0.1255
R19522 GNDA.n1673 GNDA.n1672 0.1255
R19523 GNDA.n1679 GNDA.n1678 0.1255
R19524 GNDA.n1685 GNDA.n1684 0.1255
R19525 GNDA.n1691 GNDA.n1690 0.1255
R19526 GNDA.n3836 GNDA.n3820 0.1255
R19527 GNDA.n3853 GNDA.n3852 0.1255
R19528 GNDA.n3866 GNDA.n3814 0.1255
R19529 GNDA.n3883 GNDA.n3882 0.1255
R19530 GNDA.n3896 GNDA.n3808 0.1255
R19531 GNDA.n3913 GNDA.n3912 0.1255
R19532 GNDA.n3926 GNDA.n3802 0.1255
R19533 GNDA.n3973 GNDA.n3962 0.1255
R19534 GNDA.n3990 GNDA.n3989 0.1255
R19535 GNDA.n4003 GNDA.n3956 0.1255
R19536 GNDA.n4020 GNDA.n4019 0.1255
R19537 GNDA.n4033 GNDA.n3950 0.1255
R19538 GNDA.n4050 GNDA.n4049 0.1255
R19539 GNDA.n4063 GNDA.n3944 0.1255
R19540 GNDA.n3481 GNDA.n1884 0.1255
R19541 GNDA.n3498 GNDA.n3497 0.1255
R19542 GNDA.n3511 GNDA.n1878 0.1255
R19543 GNDA.n3528 GNDA.n3527 0.1255
R19544 GNDA.n3541 GNDA.n1872 0.1255
R19545 GNDA.n3558 GNDA.n3557 0.1255
R19546 GNDA.n3571 GNDA.n1866 0.1255
R19547 GNDA.n2546 GNDA.n2531 0.1255
R19548 GNDA.n2563 GNDA.n2562 0.1255
R19549 GNDA.n2576 GNDA.n2525 0.1255
R19550 GNDA.n2593 GNDA.n2592 0.1255
R19551 GNDA.n2606 GNDA.n2519 0.1255
R19552 GNDA.n2623 GNDA.n2622 0.1255
R19553 GNDA.n2636 GNDA.n2513 0.1255
R19554 GNDA.n2829 GNDA.n2814 0.1255
R19555 GNDA.n2846 GNDA.n2845 0.1255
R19556 GNDA.n2859 GNDA.n2808 0.1255
R19557 GNDA.n2876 GNDA.n2875 0.1255
R19558 GNDA.n2889 GNDA.n2802 0.1255
R19559 GNDA.n2906 GNDA.n2905 0.1255
R19560 GNDA.n2919 GNDA.n2796 0.1255
R19561 GNDA.n2970 GNDA.n2955 0.1255
R19562 GNDA.n2987 GNDA.n2986 0.1255
R19563 GNDA.n3000 GNDA.n2949 0.1255
R19564 GNDA.n3017 GNDA.n3016 0.1255
R19565 GNDA.n3030 GNDA.n2943 0.1255
R19566 GNDA.n3047 GNDA.n3046 0.1255
R19567 GNDA.n3060 GNDA.n2937 0.1255
R19568 GNDA.n3111 GNDA.n3096 0.1255
R19569 GNDA.n3128 GNDA.n3127 0.1255
R19570 GNDA.n3141 GNDA.n3090 0.1255
R19571 GNDA.n3158 GNDA.n3157 0.1255
R19572 GNDA.n3171 GNDA.n3084 0.1255
R19573 GNDA.n3188 GNDA.n3187 0.1255
R19574 GNDA.n3201 GNDA.n3078 0.1255
R19575 GNDA.n3280 GNDA.n3279 0.1255
R19576 GNDA.n3269 GNDA.n1906 0.1255
R19577 GNDA.n3262 GNDA.n3261 0.1255
R19578 GNDA.n3251 GNDA.n1921 0.1255
R19579 GNDA.n3244 GNDA.n3243 0.1255
R19580 GNDA.n3233 GNDA.n1936 0.1255
R19581 GNDA.n3226 GNDA.n3225 0.1255
R19582 GNDA.n6364 GNDA.n6363 0.1255
R19583 GNDA.n6375 GNDA.n6341 0.1255
R19584 GNDA.n6388 GNDA.n6387 0.1255
R19585 GNDA.n6399 GNDA.n6329 0.1255
R19586 GNDA.n6412 GNDA.n6411 0.1255
R19587 GNDA.n6423 GNDA.n6317 0.1255
R19588 GNDA.n6436 GNDA.n6435 0.1255
R19589 GNDA.n6362 GNDA.n6348 0.1255
R19590 GNDA.n6377 GNDA.n6376 0.1255
R19591 GNDA.n6386 GNDA.n6336 0.1255
R19592 GNDA.n6401 GNDA.n6400 0.1255
R19593 GNDA.n6410 GNDA.n6324 0.1255
R19594 GNDA.n6425 GNDA.n6424 0.1255
R19595 GNDA.n6434 GNDA.n6312 0.1255
R19596 GNDA.n423 GNDA.n422 0.1255
R19597 GNDA.n434 GNDA.n404 0.1255
R19598 GNDA.n453 GNDA.n452 0.1255
R19599 GNDA.n464 GNDA.n398 0.1255
R19600 GNDA.n483 GNDA.n482 0.1255
R19601 GNDA.n494 GNDA.n392 0.1255
R19602 GNDA.n513 GNDA.n512 0.1255
R19603 GNDA.n421 GNDA.n407 0.1255
R19604 GNDA.n438 GNDA.n437 0.1255
R19605 GNDA.n451 GNDA.n401 0.1255
R19606 GNDA.n468 GNDA.n467 0.1255
R19607 GNDA.n481 GNDA.n395 0.1255
R19608 GNDA.n498 GNDA.n497 0.1255
R19609 GNDA.n511 GNDA.n389 0.1255
R19610 GNDA.n6286 GNDA.n361 0.119909
R19611 GNDA.n2243 GNDA.n2228 0.115503
R19612 GNDA.n1367 GNDA.n1366 0.115083
R19613 GNDA.n4802 GNDA.n4801 0.115083
R19614 GNDA.n4085 GNDA.n4084 0.115083
R19615 GNDA.n3463 GNDA.n3462 0.115083
R19616 GNDA.n6280 GNDA.n6279 0.115083
R19617 GNDA.n6279 GNDA.n6278 0.115083
R19618 GNDA.n6276 GNDA.n6275 0.115083
R19619 GNDA.n6275 GNDA.n6274 0.115083
R19620 GNDA.n6274 GNDA.n6273 0.115083
R19621 GNDA.n6273 GNDA.n6272 0.115083
R19622 GNDA.n6271 GNDA.n6270 0.115083
R19623 GNDA.n6270 GNDA.n6269 0.115083
R19624 GNDA.n6269 GNDA.n6268 0.115083
R19625 GNDA.n6267 GNDA.n6266 0.115083
R19626 GNDA.n6266 GNDA.n6265 0.115083
R19627 GNDA.n6265 GNDA.n6264 0.115083
R19628 GNDA.n2249 GNDA.n2248 0.108012
R19629 GNDA.n3216 GNDA.n2356 0.090975
R19630 GNDA.n4663 GNDA.n1596 0.0734167
R19631 GNDA.n4664 GNDA.n4663 0.0734167
R19632 GNDA.n4664 GNDA.n4661 0.0734167
R19633 GNDA.n4674 GNDA.n4659 0.0734167
R19634 GNDA.n4682 GNDA.n4659 0.0734167
R19635 GNDA.n4683 GNDA.n4682 0.0734167
R19636 GNDA.n4693 GNDA.n4692 0.0734167
R19637 GNDA.n4694 GNDA.n4693 0.0734167
R19638 GNDA.n4694 GNDA.n4655 0.0734167
R19639 GNDA.n4704 GNDA.n4653 0.0734167
R19640 GNDA.n4712 GNDA.n4653 0.0734167
R19641 GNDA.n4713 GNDA.n4712 0.0734167
R19642 GNDA.n4723 GNDA.n4722 0.0734167
R19643 GNDA.n4724 GNDA.n4723 0.0734167
R19644 GNDA.n4724 GNDA.n4649 0.0734167
R19645 GNDA.n4734 GNDA.n4647 0.0734167
R19646 GNDA.n4742 GNDA.n4647 0.0734167
R19647 GNDA.n4743 GNDA.n4742 0.0734167
R19648 GNDA.n4753 GNDA.n4752 0.0734167
R19649 GNDA.n4754 GNDA.n4753 0.0734167
R19650 GNDA.n4754 GNDA.n4643 0.0734167
R19651 GNDA.n4764 GNDA.n4641 0.0734167
R19652 GNDA.n4772 GNDA.n4641 0.0734167
R19653 GNDA.n5690 GNDA.n5689 0.0734167
R19654 GNDA.n5691 GNDA.n5690 0.0734167
R19655 GNDA.n5691 GNDA.n5684 0.0734167
R19656 GNDA.n5701 GNDA.n5682 0.0734167
R19657 GNDA.n5709 GNDA.n5682 0.0734167
R19658 GNDA.n5710 GNDA.n5709 0.0734167
R19659 GNDA.n5720 GNDA.n5719 0.0734167
R19660 GNDA.n5721 GNDA.n5720 0.0734167
R19661 GNDA.n5721 GNDA.n5678 0.0734167
R19662 GNDA.n5731 GNDA.n5676 0.0734167
R19663 GNDA.n5739 GNDA.n5676 0.0734167
R19664 GNDA.n5740 GNDA.n5739 0.0734167
R19665 GNDA.n5750 GNDA.n5749 0.0734167
R19666 GNDA.n5751 GNDA.n5750 0.0734167
R19667 GNDA.n5751 GNDA.n5672 0.0734167
R19668 GNDA.n5761 GNDA.n5670 0.0734167
R19669 GNDA.n5769 GNDA.n5670 0.0734167
R19670 GNDA.n5770 GNDA.n5769 0.0734167
R19671 GNDA.n5780 GNDA.n5779 0.0734167
R19672 GNDA.n5781 GNDA.n5780 0.0734167
R19673 GNDA.n5781 GNDA.n5666 0.0734167
R19674 GNDA.n5791 GNDA.n5664 0.0734167
R19675 GNDA.n5799 GNDA.n5664 0.0734167
R19676 GNDA.n5968 GNDA.n1368 0.0734167
R19677 GNDA.n5969 GNDA.n5968 0.0734167
R19678 GNDA.n5969 GNDA.n5966 0.0734167
R19679 GNDA.n5979 GNDA.n5964 0.0734167
R19680 GNDA.n5987 GNDA.n5964 0.0734167
R19681 GNDA.n5988 GNDA.n5987 0.0734167
R19682 GNDA.n5998 GNDA.n5997 0.0734167
R19683 GNDA.n5999 GNDA.n5998 0.0734167
R19684 GNDA.n5999 GNDA.n5960 0.0734167
R19685 GNDA.n6009 GNDA.n5958 0.0734167
R19686 GNDA.n6017 GNDA.n5958 0.0734167
R19687 GNDA.n6018 GNDA.n6017 0.0734167
R19688 GNDA.n6028 GNDA.n6027 0.0734167
R19689 GNDA.n6029 GNDA.n6028 0.0734167
R19690 GNDA.n6029 GNDA.n5954 0.0734167
R19691 GNDA.n6039 GNDA.n5952 0.0734167
R19692 GNDA.n6047 GNDA.n5952 0.0734167
R19693 GNDA.n6048 GNDA.n6047 0.0734167
R19694 GNDA.n6058 GNDA.n6057 0.0734167
R19695 GNDA.n6059 GNDA.n6058 0.0734167
R19696 GNDA.n6059 GNDA.n5948 0.0734167
R19697 GNDA.n6069 GNDA.n5946 0.0734167
R19698 GNDA.n6077 GNDA.n5946 0.0734167
R19699 GNDA.n1470 GNDA.n1423 0.0734167
R19700 GNDA.n1471 GNDA.n1470 0.0734167
R19701 GNDA.n1472 GNDA.n1471 0.0734167
R19702 GNDA.n1476 GNDA.n1475 0.0734167
R19703 GNDA.n1477 GNDA.n1476 0.0734167
R19704 GNDA.n1478 GNDA.n1477 0.0734167
R19705 GNDA.n1482 GNDA.n1481 0.0734167
R19706 GNDA.n1483 GNDA.n1482 0.0734167
R19707 GNDA.n1484 GNDA.n1483 0.0734167
R19708 GNDA.n1488 GNDA.n1487 0.0734167
R19709 GNDA.n1489 GNDA.n1488 0.0734167
R19710 GNDA.n1490 GNDA.n1489 0.0734167
R19711 GNDA.n1494 GNDA.n1493 0.0734167
R19712 GNDA.n1495 GNDA.n1494 0.0734167
R19713 GNDA.n1496 GNDA.n1495 0.0734167
R19714 GNDA.n1500 GNDA.n1499 0.0734167
R19715 GNDA.n1501 GNDA.n1500 0.0734167
R19716 GNDA.n1502 GNDA.n1501 0.0734167
R19717 GNDA.n1506 GNDA.n1505 0.0734167
R19718 GNDA.n1507 GNDA.n1506 0.0734167
R19719 GNDA.n1508 GNDA.n1507 0.0734167
R19720 GNDA.n1512 GNDA.n1511 0.0734167
R19721 GNDA.n1513 GNDA.n1512 0.0734167
R19722 GNDA.n3639 GNDA.n3638 0.0734167
R19723 GNDA.n3640 GNDA.n3639 0.0734167
R19724 GNDA.n3640 GNDA.n3632 0.0734167
R19725 GNDA.n3650 GNDA.n3630 0.0734167
R19726 GNDA.n3658 GNDA.n3630 0.0734167
R19727 GNDA.n3659 GNDA.n3658 0.0734167
R19728 GNDA.n3669 GNDA.n3668 0.0734167
R19729 GNDA.n3670 GNDA.n3669 0.0734167
R19730 GNDA.n3670 GNDA.n3626 0.0734167
R19731 GNDA.n3680 GNDA.n3624 0.0734167
R19732 GNDA.n3688 GNDA.n3624 0.0734167
R19733 GNDA.n3689 GNDA.n3688 0.0734167
R19734 GNDA.n3699 GNDA.n3698 0.0734167
R19735 GNDA.n3700 GNDA.n3699 0.0734167
R19736 GNDA.n3700 GNDA.n3620 0.0734167
R19737 GNDA.n3710 GNDA.n3618 0.0734167
R19738 GNDA.n3718 GNDA.n3618 0.0734167
R19739 GNDA.n3719 GNDA.n3718 0.0734167
R19740 GNDA.n3729 GNDA.n3728 0.0734167
R19741 GNDA.n3730 GNDA.n3729 0.0734167
R19742 GNDA.n3730 GNDA.n3614 0.0734167
R19743 GNDA.n3740 GNDA.n3612 0.0734167
R19744 GNDA.n3748 GNDA.n3612 0.0734167
R19745 GNDA.n3342 GNDA.n3295 0.0734167
R19746 GNDA.n3343 GNDA.n3342 0.0734167
R19747 GNDA.n3344 GNDA.n3343 0.0734167
R19748 GNDA.n3348 GNDA.n3347 0.0734167
R19749 GNDA.n3349 GNDA.n3348 0.0734167
R19750 GNDA.n3350 GNDA.n3349 0.0734167
R19751 GNDA.n3354 GNDA.n3353 0.0734167
R19752 GNDA.n3355 GNDA.n3354 0.0734167
R19753 GNDA.n3356 GNDA.n3355 0.0734167
R19754 GNDA.n3360 GNDA.n3359 0.0734167
R19755 GNDA.n3361 GNDA.n3360 0.0734167
R19756 GNDA.n3362 GNDA.n3361 0.0734167
R19757 GNDA.n3366 GNDA.n3365 0.0734167
R19758 GNDA.n3367 GNDA.n3366 0.0734167
R19759 GNDA.n3368 GNDA.n3367 0.0734167
R19760 GNDA.n3372 GNDA.n3371 0.0734167
R19761 GNDA.n3373 GNDA.n3372 0.0734167
R19762 GNDA.n3374 GNDA.n3373 0.0734167
R19763 GNDA.n3378 GNDA.n3377 0.0734167
R19764 GNDA.n3379 GNDA.n3378 0.0734167
R19765 GNDA.n3380 GNDA.n3379 0.0734167
R19766 GNDA.n3384 GNDA.n3383 0.0734167
R19767 GNDA.n3385 GNDA.n3384 0.0734167
R19768 GNDA.n5119 GNDA.n5069 0.0734167
R19769 GNDA.n5120 GNDA.n5119 0.0734167
R19770 GNDA.n5120 GNDA.n5117 0.0734167
R19771 GNDA.n5130 GNDA.n5115 0.0734167
R19772 GNDA.n5138 GNDA.n5115 0.0734167
R19773 GNDA.n5139 GNDA.n5138 0.0734167
R19774 GNDA.n5149 GNDA.n5148 0.0734167
R19775 GNDA.n5150 GNDA.n5149 0.0734167
R19776 GNDA.n5150 GNDA.n5111 0.0734167
R19777 GNDA.n5160 GNDA.n5109 0.0734167
R19778 GNDA.n5168 GNDA.n5109 0.0734167
R19779 GNDA.n5169 GNDA.n5168 0.0734167
R19780 GNDA.n5179 GNDA.n5178 0.0734167
R19781 GNDA.n5180 GNDA.n5179 0.0734167
R19782 GNDA.n5180 GNDA.n5105 0.0734167
R19783 GNDA.n5190 GNDA.n5103 0.0734167
R19784 GNDA.n5198 GNDA.n5103 0.0734167
R19785 GNDA.n5199 GNDA.n5198 0.0734167
R19786 GNDA.n5209 GNDA.n5208 0.0734167
R19787 GNDA.n5210 GNDA.n5209 0.0734167
R19788 GNDA.n5210 GNDA.n5099 0.0734167
R19789 GNDA.n5220 GNDA.n5097 0.0734167
R19790 GNDA.n5228 GNDA.n5097 0.0734167
R19791 GNDA.n5282 GNDA.n5235 0.0734167
R19792 GNDA.n5283 GNDA.n5282 0.0734167
R19793 GNDA.n5284 GNDA.n5283 0.0734167
R19794 GNDA.n5288 GNDA.n5287 0.0734167
R19795 GNDA.n5289 GNDA.n5288 0.0734167
R19796 GNDA.n5290 GNDA.n5289 0.0734167
R19797 GNDA.n5294 GNDA.n5293 0.0734167
R19798 GNDA.n5295 GNDA.n5294 0.0734167
R19799 GNDA.n5296 GNDA.n5295 0.0734167
R19800 GNDA.n5300 GNDA.n5299 0.0734167
R19801 GNDA.n5301 GNDA.n5300 0.0734167
R19802 GNDA.n5302 GNDA.n5301 0.0734167
R19803 GNDA.n5306 GNDA.n5305 0.0734167
R19804 GNDA.n5307 GNDA.n5306 0.0734167
R19805 GNDA.n5308 GNDA.n5307 0.0734167
R19806 GNDA.n5312 GNDA.n5311 0.0734167
R19807 GNDA.n5313 GNDA.n5312 0.0734167
R19808 GNDA.n5314 GNDA.n5313 0.0734167
R19809 GNDA.n5318 GNDA.n5317 0.0734167
R19810 GNDA.n5319 GNDA.n5318 0.0734167
R19811 GNDA.n5320 GNDA.n5319 0.0734167
R19812 GNDA.n5324 GNDA.n5323 0.0734167
R19813 GNDA.n5325 GNDA.n5324 0.0734167
R19814 GNDA.n5407 GNDA.n5406 0.0734167
R19815 GNDA.n5408 GNDA.n5407 0.0734167
R19816 GNDA.n5408 GNDA.n5067 0.0734167
R19817 GNDA.n5418 GNDA.n5065 0.0734167
R19818 GNDA.n5426 GNDA.n5065 0.0734167
R19819 GNDA.n5427 GNDA.n5426 0.0734167
R19820 GNDA.n5437 GNDA.n5436 0.0734167
R19821 GNDA.n5438 GNDA.n5437 0.0734167
R19822 GNDA.n5438 GNDA.n5061 0.0734167
R19823 GNDA.n5448 GNDA.n5059 0.0734167
R19824 GNDA.n5456 GNDA.n5059 0.0734167
R19825 GNDA.n5457 GNDA.n5456 0.0734167
R19826 GNDA.n5467 GNDA.n5466 0.0734167
R19827 GNDA.n5468 GNDA.n5467 0.0734167
R19828 GNDA.n5468 GNDA.n5055 0.0734167
R19829 GNDA.n5478 GNDA.n5053 0.0734167
R19830 GNDA.n5486 GNDA.n5053 0.0734167
R19831 GNDA.n5487 GNDA.n5486 0.0734167
R19832 GNDA.n5497 GNDA.n5496 0.0734167
R19833 GNDA.n5498 GNDA.n5497 0.0734167
R19834 GNDA.n5498 GNDA.n5049 0.0734167
R19835 GNDA.n5508 GNDA.n5047 0.0734167
R19836 GNDA.n5516 GNDA.n5047 0.0734167
R19837 GNDA.n5549 GNDA.n5548 0.0734167
R19838 GNDA.n5550 GNDA.n5549 0.0734167
R19839 GNDA.n5550 GNDA.n5542 0.0734167
R19840 GNDA.n5560 GNDA.n5540 0.0734167
R19841 GNDA.n5568 GNDA.n5540 0.0734167
R19842 GNDA.n5569 GNDA.n5568 0.0734167
R19843 GNDA.n5579 GNDA.n5578 0.0734167
R19844 GNDA.n5580 GNDA.n5579 0.0734167
R19845 GNDA.n5580 GNDA.n5536 0.0734167
R19846 GNDA.n5590 GNDA.n5534 0.0734167
R19847 GNDA.n5598 GNDA.n5534 0.0734167
R19848 GNDA.n5599 GNDA.n5598 0.0734167
R19849 GNDA.n5609 GNDA.n5608 0.0734167
R19850 GNDA.n5610 GNDA.n5609 0.0734167
R19851 GNDA.n5610 GNDA.n5530 0.0734167
R19852 GNDA.n5620 GNDA.n5528 0.0734167
R19853 GNDA.n5628 GNDA.n5528 0.0734167
R19854 GNDA.n5629 GNDA.n5628 0.0734167
R19855 GNDA.n5639 GNDA.n5638 0.0734167
R19856 GNDA.n5640 GNDA.n5639 0.0734167
R19857 GNDA.n5640 GNDA.n5524 0.0734167
R19858 GNDA.n5650 GNDA.n5522 0.0734167
R19859 GNDA.n5658 GNDA.n5522 0.0734167
R19860 GNDA.n5831 GNDA.n5830 0.0734167
R19861 GNDA.n5832 GNDA.n5831 0.0734167
R19862 GNDA.n5832 GNDA.n5825 0.0734167
R19863 GNDA.n5842 GNDA.n5823 0.0734167
R19864 GNDA.n5850 GNDA.n5823 0.0734167
R19865 GNDA.n5851 GNDA.n5850 0.0734167
R19866 GNDA.n5861 GNDA.n5860 0.0734167
R19867 GNDA.n5862 GNDA.n5861 0.0734167
R19868 GNDA.n5862 GNDA.n5819 0.0734167
R19869 GNDA.n5872 GNDA.n5817 0.0734167
R19870 GNDA.n5880 GNDA.n5817 0.0734167
R19871 GNDA.n5881 GNDA.n5880 0.0734167
R19872 GNDA.n5891 GNDA.n5890 0.0734167
R19873 GNDA.n5892 GNDA.n5891 0.0734167
R19874 GNDA.n5892 GNDA.n5813 0.0734167
R19875 GNDA.n5902 GNDA.n5811 0.0734167
R19876 GNDA.n5910 GNDA.n5811 0.0734167
R19877 GNDA.n5911 GNDA.n5910 0.0734167
R19878 GNDA.n5921 GNDA.n5920 0.0734167
R19879 GNDA.n5922 GNDA.n5921 0.0734167
R19880 GNDA.n5922 GNDA.n5807 0.0734167
R19881 GNDA.n5932 GNDA.n5805 0.0734167
R19882 GNDA.n5940 GNDA.n5805 0.0734167
R19883 GNDA.n4812 GNDA.n4811 0.0734167
R19884 GNDA.n4813 GNDA.n4812 0.0734167
R19885 GNDA.n4813 GNDA.n1418 0.0734167
R19886 GNDA.n4823 GNDA.n1416 0.0734167
R19887 GNDA.n4831 GNDA.n1416 0.0734167
R19888 GNDA.n4832 GNDA.n4831 0.0734167
R19889 GNDA.n4842 GNDA.n4841 0.0734167
R19890 GNDA.n4843 GNDA.n4842 0.0734167
R19891 GNDA.n4843 GNDA.n1412 0.0734167
R19892 GNDA.n4853 GNDA.n1410 0.0734167
R19893 GNDA.n4861 GNDA.n1410 0.0734167
R19894 GNDA.n4862 GNDA.n4861 0.0734167
R19895 GNDA.n4872 GNDA.n4871 0.0734167
R19896 GNDA.n4873 GNDA.n4872 0.0734167
R19897 GNDA.n4873 GNDA.n1406 0.0734167
R19898 GNDA.n4883 GNDA.n1404 0.0734167
R19899 GNDA.n4891 GNDA.n1404 0.0734167
R19900 GNDA.n4892 GNDA.n4891 0.0734167
R19901 GNDA.n4902 GNDA.n4901 0.0734167
R19902 GNDA.n4903 GNDA.n4902 0.0734167
R19903 GNDA.n4903 GNDA.n1400 0.0734167
R19904 GNDA.n4913 GNDA.n1398 0.0734167
R19905 GNDA.n4921 GNDA.n1398 0.0734167
R19906 GNDA.n4526 GNDA.n4525 0.0734167
R19907 GNDA.n4527 GNDA.n4526 0.0734167
R19908 GNDA.n4527 GNDA.n4519 0.0734167
R19909 GNDA.n4537 GNDA.n4517 0.0734167
R19910 GNDA.n4545 GNDA.n4517 0.0734167
R19911 GNDA.n4546 GNDA.n4545 0.0734167
R19912 GNDA.n4556 GNDA.n4555 0.0734167
R19913 GNDA.n4557 GNDA.n4556 0.0734167
R19914 GNDA.n4557 GNDA.n4513 0.0734167
R19915 GNDA.n4567 GNDA.n4511 0.0734167
R19916 GNDA.n4575 GNDA.n4511 0.0734167
R19917 GNDA.n4576 GNDA.n4575 0.0734167
R19918 GNDA.n4586 GNDA.n4585 0.0734167
R19919 GNDA.n4587 GNDA.n4586 0.0734167
R19920 GNDA.n4587 GNDA.n4507 0.0734167
R19921 GNDA.n4597 GNDA.n4505 0.0734167
R19922 GNDA.n4605 GNDA.n4505 0.0734167
R19923 GNDA.n4606 GNDA.n4605 0.0734167
R19924 GNDA.n4616 GNDA.n4615 0.0734167
R19925 GNDA.n4617 GNDA.n4616 0.0734167
R19926 GNDA.n4617 GNDA.n4501 0.0734167
R19927 GNDA.n4627 GNDA.n4499 0.0734167
R19928 GNDA.n4635 GNDA.n4499 0.0734167
R19929 GNDA.n4337 GNDA.n4336 0.0734167
R19930 GNDA.n4338 GNDA.n4337 0.0734167
R19931 GNDA.n4338 GNDA.n4330 0.0734167
R19932 GNDA.n4348 GNDA.n4328 0.0734167
R19933 GNDA.n4356 GNDA.n4328 0.0734167
R19934 GNDA.n4357 GNDA.n4356 0.0734167
R19935 GNDA.n4367 GNDA.n4366 0.0734167
R19936 GNDA.n4368 GNDA.n4367 0.0734167
R19937 GNDA.n4368 GNDA.n4324 0.0734167
R19938 GNDA.n4378 GNDA.n4322 0.0734167
R19939 GNDA.n4386 GNDA.n4322 0.0734167
R19940 GNDA.n4387 GNDA.n4386 0.0734167
R19941 GNDA.n4397 GNDA.n4396 0.0734167
R19942 GNDA.n4398 GNDA.n4397 0.0734167
R19943 GNDA.n4398 GNDA.n4318 0.0734167
R19944 GNDA.n4408 GNDA.n4316 0.0734167
R19945 GNDA.n4416 GNDA.n4316 0.0734167
R19946 GNDA.n4417 GNDA.n4416 0.0734167
R19947 GNDA.n4427 GNDA.n4426 0.0734167
R19948 GNDA.n4428 GNDA.n4427 0.0734167
R19949 GNDA.n4428 GNDA.n4312 0.0734167
R19950 GNDA.n4438 GNDA.n4310 0.0734167
R19951 GNDA.n4446 GNDA.n4310 0.0734167
R19952 GNDA.n4171 GNDA.n4170 0.0734167
R19953 GNDA.n4172 GNDA.n4171 0.0734167
R19954 GNDA.n4172 GNDA.n1646 0.0734167
R19955 GNDA.n4182 GNDA.n1644 0.0734167
R19956 GNDA.n4190 GNDA.n1644 0.0734167
R19957 GNDA.n4191 GNDA.n4190 0.0734167
R19958 GNDA.n4201 GNDA.n4200 0.0734167
R19959 GNDA.n4202 GNDA.n4201 0.0734167
R19960 GNDA.n4202 GNDA.n1640 0.0734167
R19961 GNDA.n4212 GNDA.n1638 0.0734167
R19962 GNDA.n4220 GNDA.n1638 0.0734167
R19963 GNDA.n4221 GNDA.n4220 0.0734167
R19964 GNDA.n4231 GNDA.n4230 0.0734167
R19965 GNDA.n4232 GNDA.n4231 0.0734167
R19966 GNDA.n4232 GNDA.n1634 0.0734167
R19967 GNDA.n4242 GNDA.n1632 0.0734167
R19968 GNDA.n4250 GNDA.n1632 0.0734167
R19969 GNDA.n4251 GNDA.n4250 0.0734167
R19970 GNDA.n4261 GNDA.n4260 0.0734167
R19971 GNDA.n4262 GNDA.n4261 0.0734167
R19972 GNDA.n4262 GNDA.n1628 0.0734167
R19973 GNDA.n4272 GNDA.n1626 0.0734167
R19974 GNDA.n4280 GNDA.n1626 0.0734167
R19975 GNDA.n1696 GNDA.n1649 0.0734167
R19976 GNDA.n1697 GNDA.n1696 0.0734167
R19977 GNDA.n1698 GNDA.n1697 0.0734167
R19978 GNDA.n1702 GNDA.n1701 0.0734167
R19979 GNDA.n1703 GNDA.n1702 0.0734167
R19980 GNDA.n1704 GNDA.n1703 0.0734167
R19981 GNDA.n1708 GNDA.n1707 0.0734167
R19982 GNDA.n1709 GNDA.n1708 0.0734167
R19983 GNDA.n1710 GNDA.n1709 0.0734167
R19984 GNDA.n1714 GNDA.n1713 0.0734167
R19985 GNDA.n1715 GNDA.n1714 0.0734167
R19986 GNDA.n1716 GNDA.n1715 0.0734167
R19987 GNDA.n1720 GNDA.n1719 0.0734167
R19988 GNDA.n1721 GNDA.n1720 0.0734167
R19989 GNDA.n1722 GNDA.n1721 0.0734167
R19990 GNDA.n1726 GNDA.n1725 0.0734167
R19991 GNDA.n1727 GNDA.n1726 0.0734167
R19992 GNDA.n1728 GNDA.n1727 0.0734167
R19993 GNDA.n1732 GNDA.n1731 0.0734167
R19994 GNDA.n1733 GNDA.n1732 0.0734167
R19995 GNDA.n1734 GNDA.n1733 0.0734167
R19996 GNDA.n1738 GNDA.n1737 0.0734167
R19997 GNDA.n1739 GNDA.n1738 0.0734167
R19998 GNDA.n3828 GNDA.n3827 0.0734167
R19999 GNDA.n3829 GNDA.n3828 0.0734167
R20000 GNDA.n3829 GNDA.n3821 0.0734167
R20001 GNDA.n3839 GNDA.n3819 0.0734167
R20002 GNDA.n3847 GNDA.n3819 0.0734167
R20003 GNDA.n3848 GNDA.n3847 0.0734167
R20004 GNDA.n3858 GNDA.n3857 0.0734167
R20005 GNDA.n3859 GNDA.n3858 0.0734167
R20006 GNDA.n3859 GNDA.n3815 0.0734167
R20007 GNDA.n3869 GNDA.n3813 0.0734167
R20008 GNDA.n3877 GNDA.n3813 0.0734167
R20009 GNDA.n3878 GNDA.n3877 0.0734167
R20010 GNDA.n3888 GNDA.n3887 0.0734167
R20011 GNDA.n3889 GNDA.n3888 0.0734167
R20012 GNDA.n3889 GNDA.n3809 0.0734167
R20013 GNDA.n3899 GNDA.n3807 0.0734167
R20014 GNDA.n3907 GNDA.n3807 0.0734167
R20015 GNDA.n3908 GNDA.n3907 0.0734167
R20016 GNDA.n3918 GNDA.n3917 0.0734167
R20017 GNDA.n3919 GNDA.n3918 0.0734167
R20018 GNDA.n3919 GNDA.n3803 0.0734167
R20019 GNDA.n3929 GNDA.n3801 0.0734167
R20020 GNDA.n3937 GNDA.n3801 0.0734167
R20021 GNDA.n3965 GNDA.n1835 0.0734167
R20022 GNDA.n3966 GNDA.n3965 0.0734167
R20023 GNDA.n3966 GNDA.n3963 0.0734167
R20024 GNDA.n3976 GNDA.n3961 0.0734167
R20025 GNDA.n3984 GNDA.n3961 0.0734167
R20026 GNDA.n3985 GNDA.n3984 0.0734167
R20027 GNDA.n3995 GNDA.n3994 0.0734167
R20028 GNDA.n3996 GNDA.n3995 0.0734167
R20029 GNDA.n3996 GNDA.n3957 0.0734167
R20030 GNDA.n4006 GNDA.n3955 0.0734167
R20031 GNDA.n4014 GNDA.n3955 0.0734167
R20032 GNDA.n4015 GNDA.n4014 0.0734167
R20033 GNDA.n4025 GNDA.n4024 0.0734167
R20034 GNDA.n4026 GNDA.n4025 0.0734167
R20035 GNDA.n4026 GNDA.n3951 0.0734167
R20036 GNDA.n4036 GNDA.n3949 0.0734167
R20037 GNDA.n4044 GNDA.n3949 0.0734167
R20038 GNDA.n4045 GNDA.n4044 0.0734167
R20039 GNDA.n4055 GNDA.n4054 0.0734167
R20040 GNDA.n4056 GNDA.n4055 0.0734167
R20041 GNDA.n4056 GNDA.n3945 0.0734167
R20042 GNDA.n4066 GNDA.n3943 0.0734167
R20043 GNDA.n4074 GNDA.n3943 0.0734167
R20044 GNDA.n3473 GNDA.n3472 0.0734167
R20045 GNDA.n3474 GNDA.n3473 0.0734167
R20046 GNDA.n3474 GNDA.n1885 0.0734167
R20047 GNDA.n3484 GNDA.n1883 0.0734167
R20048 GNDA.n3492 GNDA.n1883 0.0734167
R20049 GNDA.n3493 GNDA.n3492 0.0734167
R20050 GNDA.n3503 GNDA.n3502 0.0734167
R20051 GNDA.n3504 GNDA.n3503 0.0734167
R20052 GNDA.n3504 GNDA.n1879 0.0734167
R20053 GNDA.n3514 GNDA.n1877 0.0734167
R20054 GNDA.n3522 GNDA.n1877 0.0734167
R20055 GNDA.n3523 GNDA.n3522 0.0734167
R20056 GNDA.n3533 GNDA.n3532 0.0734167
R20057 GNDA.n3534 GNDA.n3533 0.0734167
R20058 GNDA.n3534 GNDA.n1873 0.0734167
R20059 GNDA.n3544 GNDA.n1871 0.0734167
R20060 GNDA.n3552 GNDA.n1871 0.0734167
R20061 GNDA.n3553 GNDA.n3552 0.0734167
R20062 GNDA.n3563 GNDA.n3562 0.0734167
R20063 GNDA.n3564 GNDA.n3563 0.0734167
R20064 GNDA.n3564 GNDA.n1867 0.0734167
R20065 GNDA.n3574 GNDA.n1865 0.0734167
R20066 GNDA.n3582 GNDA.n1865 0.0734167
R20067 GNDA.n2538 GNDA.n2537 0.0734167
R20068 GNDA.n2539 GNDA.n2538 0.0734167
R20069 GNDA.n2539 GNDA.n2532 0.0734167
R20070 GNDA.n2549 GNDA.n2530 0.0734167
R20071 GNDA.n2557 GNDA.n2530 0.0734167
R20072 GNDA.n2558 GNDA.n2557 0.0734167
R20073 GNDA.n2568 GNDA.n2567 0.0734167
R20074 GNDA.n2569 GNDA.n2568 0.0734167
R20075 GNDA.n2569 GNDA.n2526 0.0734167
R20076 GNDA.n2579 GNDA.n2524 0.0734167
R20077 GNDA.n2587 GNDA.n2524 0.0734167
R20078 GNDA.n2588 GNDA.n2587 0.0734167
R20079 GNDA.n2598 GNDA.n2597 0.0734167
R20080 GNDA.n2599 GNDA.n2598 0.0734167
R20081 GNDA.n2599 GNDA.n2520 0.0734167
R20082 GNDA.n2609 GNDA.n2518 0.0734167
R20083 GNDA.n2617 GNDA.n2518 0.0734167
R20084 GNDA.n2618 GNDA.n2617 0.0734167
R20085 GNDA.n2628 GNDA.n2627 0.0734167
R20086 GNDA.n2629 GNDA.n2628 0.0734167
R20087 GNDA.n2629 GNDA.n2514 0.0734167
R20088 GNDA.n2639 GNDA.n2512 0.0734167
R20089 GNDA.n2647 GNDA.n2512 0.0734167
R20090 GNDA.n2821 GNDA.n2820 0.0734167
R20091 GNDA.n2822 GNDA.n2821 0.0734167
R20092 GNDA.n2822 GNDA.n2815 0.0734167
R20093 GNDA.n2832 GNDA.n2813 0.0734167
R20094 GNDA.n2840 GNDA.n2813 0.0734167
R20095 GNDA.n2841 GNDA.n2840 0.0734167
R20096 GNDA.n2851 GNDA.n2850 0.0734167
R20097 GNDA.n2852 GNDA.n2851 0.0734167
R20098 GNDA.n2852 GNDA.n2809 0.0734167
R20099 GNDA.n2862 GNDA.n2807 0.0734167
R20100 GNDA.n2870 GNDA.n2807 0.0734167
R20101 GNDA.n2871 GNDA.n2870 0.0734167
R20102 GNDA.n2881 GNDA.n2880 0.0734167
R20103 GNDA.n2882 GNDA.n2881 0.0734167
R20104 GNDA.n2882 GNDA.n2803 0.0734167
R20105 GNDA.n2892 GNDA.n2801 0.0734167
R20106 GNDA.n2900 GNDA.n2801 0.0734167
R20107 GNDA.n2901 GNDA.n2900 0.0734167
R20108 GNDA.n2911 GNDA.n2910 0.0734167
R20109 GNDA.n2912 GNDA.n2911 0.0734167
R20110 GNDA.n2912 GNDA.n2797 0.0734167
R20111 GNDA.n2922 GNDA.n2795 0.0734167
R20112 GNDA.n2930 GNDA.n2795 0.0734167
R20113 GNDA.n2962 GNDA.n2961 0.0734167
R20114 GNDA.n2963 GNDA.n2962 0.0734167
R20115 GNDA.n2963 GNDA.n2956 0.0734167
R20116 GNDA.n2973 GNDA.n2954 0.0734167
R20117 GNDA.n2981 GNDA.n2954 0.0734167
R20118 GNDA.n2982 GNDA.n2981 0.0734167
R20119 GNDA.n2992 GNDA.n2991 0.0734167
R20120 GNDA.n2993 GNDA.n2992 0.0734167
R20121 GNDA.n2993 GNDA.n2950 0.0734167
R20122 GNDA.n3003 GNDA.n2948 0.0734167
R20123 GNDA.n3011 GNDA.n2948 0.0734167
R20124 GNDA.n3012 GNDA.n3011 0.0734167
R20125 GNDA.n3022 GNDA.n3021 0.0734167
R20126 GNDA.n3023 GNDA.n3022 0.0734167
R20127 GNDA.n3023 GNDA.n2944 0.0734167
R20128 GNDA.n3033 GNDA.n2942 0.0734167
R20129 GNDA.n3041 GNDA.n2942 0.0734167
R20130 GNDA.n3042 GNDA.n3041 0.0734167
R20131 GNDA.n3052 GNDA.n3051 0.0734167
R20132 GNDA.n3053 GNDA.n3052 0.0734167
R20133 GNDA.n3053 GNDA.n2938 0.0734167
R20134 GNDA.n3063 GNDA.n2936 0.0734167
R20135 GNDA.n3071 GNDA.n2936 0.0734167
R20136 GNDA.n3103 GNDA.n3102 0.0734167
R20137 GNDA.n3104 GNDA.n3103 0.0734167
R20138 GNDA.n3104 GNDA.n3097 0.0734167
R20139 GNDA.n3114 GNDA.n3095 0.0734167
R20140 GNDA.n3122 GNDA.n3095 0.0734167
R20141 GNDA.n3123 GNDA.n3122 0.0734167
R20142 GNDA.n3133 GNDA.n3132 0.0734167
R20143 GNDA.n3134 GNDA.n3133 0.0734167
R20144 GNDA.n3134 GNDA.n3091 0.0734167
R20145 GNDA.n3144 GNDA.n3089 0.0734167
R20146 GNDA.n3152 GNDA.n3089 0.0734167
R20147 GNDA.n3153 GNDA.n3152 0.0734167
R20148 GNDA.n3163 GNDA.n3162 0.0734167
R20149 GNDA.n3164 GNDA.n3163 0.0734167
R20150 GNDA.n3164 GNDA.n3085 0.0734167
R20151 GNDA.n3174 GNDA.n3083 0.0734167
R20152 GNDA.n3182 GNDA.n3083 0.0734167
R20153 GNDA.n3183 GNDA.n3182 0.0734167
R20154 GNDA.n3193 GNDA.n3192 0.0734167
R20155 GNDA.n3194 GNDA.n3193 0.0734167
R20156 GNDA.n3194 GNDA.n3079 0.0734167
R20157 GNDA.n3204 GNDA.n3077 0.0734167
R20158 GNDA.n3212 GNDA.n3077 0.0734167
R20159 GNDA.n3284 GNDA.n1892 0.0734167
R20160 GNDA.n3284 GNDA.n3283 0.0734167
R20161 GNDA.n3283 GNDA.n3282 0.0734167
R20162 GNDA.n3277 GNDA.n3276 0.0734167
R20163 GNDA.n3276 GNDA.n1902 0.0734167
R20164 GNDA.n3272 GNDA.n1902 0.0734167
R20165 GNDA.n3266 GNDA.n1907 0.0734167
R20166 GNDA.n3266 GNDA.n3265 0.0734167
R20167 GNDA.n3265 GNDA.n3264 0.0734167
R20168 GNDA.n3259 GNDA.n3258 0.0734167
R20169 GNDA.n3258 GNDA.n1917 0.0734167
R20170 GNDA.n3254 GNDA.n1917 0.0734167
R20171 GNDA.n3248 GNDA.n1922 0.0734167
R20172 GNDA.n3248 GNDA.n3247 0.0734167
R20173 GNDA.n3247 GNDA.n3246 0.0734167
R20174 GNDA.n3241 GNDA.n3240 0.0734167
R20175 GNDA.n3240 GNDA.n1932 0.0734167
R20176 GNDA.n3236 GNDA.n1932 0.0734167
R20177 GNDA.n3230 GNDA.n1937 0.0734167
R20178 GNDA.n3230 GNDA.n3229 0.0734167
R20179 GNDA.n3229 GNDA.n3228 0.0734167
R20180 GNDA.n3223 GNDA.n3222 0.0734167
R20181 GNDA.n3222 GNDA.n1947 0.0734167
R20182 GNDA.n2702 GNDA.n2701 0.0734167
R20183 GNDA.n2703 GNDA.n2702 0.0734167
R20184 GNDA.n2703 GNDA.n2693 0.0734167
R20185 GNDA.n2711 GNDA.n2689 0.0734167
R20186 GNDA.n2717 GNDA.n2689 0.0734167
R20187 GNDA.n2718 GNDA.n2717 0.0734167
R20188 GNDA.n2726 GNDA.n2725 0.0734167
R20189 GNDA.n2727 GNDA.n2726 0.0734167
R20190 GNDA.n2727 GNDA.n2681 0.0734167
R20191 GNDA.n2735 GNDA.n2677 0.0734167
R20192 GNDA.n2741 GNDA.n2677 0.0734167
R20193 GNDA.n2742 GNDA.n2741 0.0734167
R20194 GNDA.n2750 GNDA.n2749 0.0734167
R20195 GNDA.n2751 GNDA.n2750 0.0734167
R20196 GNDA.n2751 GNDA.n2669 0.0734167
R20197 GNDA.n2759 GNDA.n2665 0.0734167
R20198 GNDA.n2765 GNDA.n2665 0.0734167
R20199 GNDA.n2766 GNDA.n2765 0.0734167
R20200 GNDA.n2774 GNDA.n2773 0.0734167
R20201 GNDA.n2775 GNDA.n2774 0.0734167
R20202 GNDA.n2775 GNDA.n2657 0.0734167
R20203 GNDA.n2783 GNDA.n2653 0.0734167
R20204 GNDA.n2789 GNDA.n2653 0.0734167
R20205 GNDA.n4778 GNDA.n1596 0.0682083
R20206 GNDA.n4672 GNDA.n4661 0.0682083
R20207 GNDA.n4674 GNDA.n4673 0.0682083
R20208 GNDA.n4684 GNDA.n4683 0.0682083
R20209 GNDA.n4692 GNDA.n4657 0.0682083
R20210 GNDA.n4702 GNDA.n4655 0.0682083
R20211 GNDA.n4704 GNDA.n4703 0.0682083
R20212 GNDA.n4714 GNDA.n4713 0.0682083
R20213 GNDA.n4722 GNDA.n4651 0.0682083
R20214 GNDA.n4732 GNDA.n4649 0.0682083
R20215 GNDA.n4734 GNDA.n4733 0.0682083
R20216 GNDA.n4744 GNDA.n4743 0.0682083
R20217 GNDA.n4752 GNDA.n4645 0.0682083
R20218 GNDA.n4762 GNDA.n4643 0.0682083
R20219 GNDA.n4764 GNDA.n4763 0.0682083
R20220 GNDA.n5689 GNDA.n1361 0.0682083
R20221 GNDA.n5699 GNDA.n5684 0.0682083
R20222 GNDA.n5701 GNDA.n5700 0.0682083
R20223 GNDA.n5711 GNDA.n5710 0.0682083
R20224 GNDA.n5719 GNDA.n5680 0.0682083
R20225 GNDA.n5729 GNDA.n5678 0.0682083
R20226 GNDA.n5731 GNDA.n5730 0.0682083
R20227 GNDA.n5741 GNDA.n5740 0.0682083
R20228 GNDA.n5749 GNDA.n5674 0.0682083
R20229 GNDA.n5759 GNDA.n5672 0.0682083
R20230 GNDA.n5761 GNDA.n5760 0.0682083
R20231 GNDA.n5771 GNDA.n5770 0.0682083
R20232 GNDA.n5779 GNDA.n5668 0.0682083
R20233 GNDA.n5789 GNDA.n5666 0.0682083
R20234 GNDA.n5791 GNDA.n5790 0.0682083
R20235 GNDA.n6083 GNDA.n1368 0.0682083
R20236 GNDA.n5977 GNDA.n5966 0.0682083
R20237 GNDA.n5979 GNDA.n5978 0.0682083
R20238 GNDA.n5989 GNDA.n5988 0.0682083
R20239 GNDA.n5997 GNDA.n5962 0.0682083
R20240 GNDA.n6007 GNDA.n5960 0.0682083
R20241 GNDA.n6009 GNDA.n6008 0.0682083
R20242 GNDA.n6019 GNDA.n6018 0.0682083
R20243 GNDA.n6027 GNDA.n5956 0.0682083
R20244 GNDA.n6037 GNDA.n5954 0.0682083
R20245 GNDA.n6039 GNDA.n6038 0.0682083
R20246 GNDA.n6049 GNDA.n6048 0.0682083
R20247 GNDA.n6057 GNDA.n5950 0.0682083
R20248 GNDA.n6067 GNDA.n5948 0.0682083
R20249 GNDA.n6069 GNDA.n6068 0.0682083
R20250 GNDA.n1587 GNDA.n1423 0.0682083
R20251 GNDA.n1473 GNDA.n1472 0.0682083
R20252 GNDA.n1475 GNDA.n1474 0.0682083
R20253 GNDA.n1479 GNDA.n1478 0.0682083
R20254 GNDA.n1481 GNDA.n1480 0.0682083
R20255 GNDA.n1485 GNDA.n1484 0.0682083
R20256 GNDA.n1487 GNDA.n1486 0.0682083
R20257 GNDA.n1491 GNDA.n1490 0.0682083
R20258 GNDA.n1493 GNDA.n1492 0.0682083
R20259 GNDA.n1497 GNDA.n1496 0.0682083
R20260 GNDA.n1499 GNDA.n1498 0.0682083
R20261 GNDA.n1503 GNDA.n1502 0.0682083
R20262 GNDA.n1505 GNDA.n1504 0.0682083
R20263 GNDA.n1509 GNDA.n1508 0.0682083
R20264 GNDA.n1511 GNDA.n1510 0.0682083
R20265 GNDA.n3638 GNDA.n3634 0.0682083
R20266 GNDA.n3648 GNDA.n3632 0.0682083
R20267 GNDA.n3650 GNDA.n3649 0.0682083
R20268 GNDA.n3660 GNDA.n3659 0.0682083
R20269 GNDA.n3668 GNDA.n3628 0.0682083
R20270 GNDA.n3678 GNDA.n3626 0.0682083
R20271 GNDA.n3680 GNDA.n3679 0.0682083
R20272 GNDA.n3690 GNDA.n3689 0.0682083
R20273 GNDA.n3698 GNDA.n3622 0.0682083
R20274 GNDA.n3708 GNDA.n3620 0.0682083
R20275 GNDA.n3710 GNDA.n3709 0.0682083
R20276 GNDA.n3720 GNDA.n3719 0.0682083
R20277 GNDA.n3728 GNDA.n3616 0.0682083
R20278 GNDA.n3738 GNDA.n3614 0.0682083
R20279 GNDA.n3740 GNDA.n3739 0.0682083
R20280 GNDA.n3459 GNDA.n3295 0.0682083
R20281 GNDA.n3345 GNDA.n3344 0.0682083
R20282 GNDA.n3347 GNDA.n3346 0.0682083
R20283 GNDA.n3351 GNDA.n3350 0.0682083
R20284 GNDA.n3353 GNDA.n3352 0.0682083
R20285 GNDA.n3357 GNDA.n3356 0.0682083
R20286 GNDA.n3359 GNDA.n3358 0.0682083
R20287 GNDA.n3363 GNDA.n3362 0.0682083
R20288 GNDA.n3365 GNDA.n3364 0.0682083
R20289 GNDA.n3369 GNDA.n3368 0.0682083
R20290 GNDA.n3371 GNDA.n3370 0.0682083
R20291 GNDA.n3375 GNDA.n3374 0.0682083
R20292 GNDA.n3377 GNDA.n3376 0.0682083
R20293 GNDA.n3381 GNDA.n3380 0.0682083
R20294 GNDA.n3383 GNDA.n3382 0.0682083
R20295 GNDA.n5234 GNDA.n5069 0.0682083
R20296 GNDA.n5128 GNDA.n5117 0.0682083
R20297 GNDA.n5130 GNDA.n5129 0.0682083
R20298 GNDA.n5140 GNDA.n5139 0.0682083
R20299 GNDA.n5148 GNDA.n5113 0.0682083
R20300 GNDA.n5158 GNDA.n5111 0.0682083
R20301 GNDA.n5160 GNDA.n5159 0.0682083
R20302 GNDA.n5170 GNDA.n5169 0.0682083
R20303 GNDA.n5178 GNDA.n5107 0.0682083
R20304 GNDA.n5188 GNDA.n5105 0.0682083
R20305 GNDA.n5190 GNDA.n5189 0.0682083
R20306 GNDA.n5200 GNDA.n5199 0.0682083
R20307 GNDA.n5208 GNDA.n5101 0.0682083
R20308 GNDA.n5218 GNDA.n5099 0.0682083
R20309 GNDA.n5220 GNDA.n5219 0.0682083
R20310 GNDA.n5399 GNDA.n5235 0.0682083
R20311 GNDA.n5285 GNDA.n5284 0.0682083
R20312 GNDA.n5287 GNDA.n5286 0.0682083
R20313 GNDA.n5291 GNDA.n5290 0.0682083
R20314 GNDA.n5293 GNDA.n5292 0.0682083
R20315 GNDA.n5297 GNDA.n5296 0.0682083
R20316 GNDA.n5299 GNDA.n5298 0.0682083
R20317 GNDA.n5303 GNDA.n5302 0.0682083
R20318 GNDA.n5305 GNDA.n5304 0.0682083
R20319 GNDA.n5309 GNDA.n5308 0.0682083
R20320 GNDA.n5311 GNDA.n5310 0.0682083
R20321 GNDA.n5315 GNDA.n5314 0.0682083
R20322 GNDA.n5317 GNDA.n5316 0.0682083
R20323 GNDA.n5321 GNDA.n5320 0.0682083
R20324 GNDA.n5323 GNDA.n5322 0.0682083
R20325 GNDA.n5406 GNDA.n5402 0.0682083
R20326 GNDA.n5416 GNDA.n5067 0.0682083
R20327 GNDA.n5418 GNDA.n5417 0.0682083
R20328 GNDA.n5428 GNDA.n5427 0.0682083
R20329 GNDA.n5436 GNDA.n5063 0.0682083
R20330 GNDA.n5446 GNDA.n5061 0.0682083
R20331 GNDA.n5448 GNDA.n5447 0.0682083
R20332 GNDA.n5458 GNDA.n5457 0.0682083
R20333 GNDA.n5466 GNDA.n5057 0.0682083
R20334 GNDA.n5476 GNDA.n5055 0.0682083
R20335 GNDA.n5478 GNDA.n5477 0.0682083
R20336 GNDA.n5488 GNDA.n5487 0.0682083
R20337 GNDA.n5496 GNDA.n5051 0.0682083
R20338 GNDA.n5506 GNDA.n5049 0.0682083
R20339 GNDA.n5508 GNDA.n5507 0.0682083
R20340 GNDA.n5548 GNDA.n5544 0.0682083
R20341 GNDA.n5558 GNDA.n5542 0.0682083
R20342 GNDA.n5560 GNDA.n5559 0.0682083
R20343 GNDA.n5570 GNDA.n5569 0.0682083
R20344 GNDA.n5578 GNDA.n5538 0.0682083
R20345 GNDA.n5588 GNDA.n5536 0.0682083
R20346 GNDA.n5590 GNDA.n5589 0.0682083
R20347 GNDA.n5600 GNDA.n5599 0.0682083
R20348 GNDA.n5608 GNDA.n5532 0.0682083
R20349 GNDA.n5618 GNDA.n5530 0.0682083
R20350 GNDA.n5620 GNDA.n5619 0.0682083
R20351 GNDA.n5630 GNDA.n5629 0.0682083
R20352 GNDA.n5638 GNDA.n5526 0.0682083
R20353 GNDA.n5648 GNDA.n5524 0.0682083
R20354 GNDA.n5650 GNDA.n5649 0.0682083
R20355 GNDA.n5830 GNDA.n1363 0.0682083
R20356 GNDA.n5840 GNDA.n5825 0.0682083
R20357 GNDA.n5842 GNDA.n5841 0.0682083
R20358 GNDA.n5852 GNDA.n5851 0.0682083
R20359 GNDA.n5860 GNDA.n5821 0.0682083
R20360 GNDA.n5870 GNDA.n5819 0.0682083
R20361 GNDA.n5872 GNDA.n5871 0.0682083
R20362 GNDA.n5882 GNDA.n5881 0.0682083
R20363 GNDA.n5890 GNDA.n5815 0.0682083
R20364 GNDA.n5900 GNDA.n5813 0.0682083
R20365 GNDA.n5902 GNDA.n5901 0.0682083
R20366 GNDA.n5912 GNDA.n5911 0.0682083
R20367 GNDA.n5920 GNDA.n5809 0.0682083
R20368 GNDA.n5930 GNDA.n5807 0.0682083
R20369 GNDA.n5932 GNDA.n5931 0.0682083
R20370 GNDA.n4811 GNDA.n4807 0.0682083
R20371 GNDA.n4821 GNDA.n1418 0.0682083
R20372 GNDA.n4823 GNDA.n4822 0.0682083
R20373 GNDA.n4833 GNDA.n4832 0.0682083
R20374 GNDA.n4841 GNDA.n1414 0.0682083
R20375 GNDA.n4851 GNDA.n1412 0.0682083
R20376 GNDA.n4853 GNDA.n4852 0.0682083
R20377 GNDA.n4863 GNDA.n4862 0.0682083
R20378 GNDA.n4871 GNDA.n1408 0.0682083
R20379 GNDA.n4881 GNDA.n1406 0.0682083
R20380 GNDA.n4883 GNDA.n4882 0.0682083
R20381 GNDA.n4893 GNDA.n4892 0.0682083
R20382 GNDA.n4901 GNDA.n1402 0.0682083
R20383 GNDA.n4911 GNDA.n1400 0.0682083
R20384 GNDA.n4913 GNDA.n4912 0.0682083
R20385 GNDA.n4525 GNDA.n4521 0.0682083
R20386 GNDA.n4535 GNDA.n4519 0.0682083
R20387 GNDA.n4537 GNDA.n4536 0.0682083
R20388 GNDA.n4547 GNDA.n4546 0.0682083
R20389 GNDA.n4555 GNDA.n4515 0.0682083
R20390 GNDA.n4565 GNDA.n4513 0.0682083
R20391 GNDA.n4567 GNDA.n4566 0.0682083
R20392 GNDA.n4577 GNDA.n4576 0.0682083
R20393 GNDA.n4585 GNDA.n4509 0.0682083
R20394 GNDA.n4595 GNDA.n4507 0.0682083
R20395 GNDA.n4597 GNDA.n4596 0.0682083
R20396 GNDA.n4607 GNDA.n4606 0.0682083
R20397 GNDA.n4615 GNDA.n4503 0.0682083
R20398 GNDA.n4625 GNDA.n4501 0.0682083
R20399 GNDA.n4627 GNDA.n4626 0.0682083
R20400 GNDA.n4336 GNDA.n4332 0.0682083
R20401 GNDA.n4346 GNDA.n4330 0.0682083
R20402 GNDA.n4348 GNDA.n4347 0.0682083
R20403 GNDA.n4358 GNDA.n4357 0.0682083
R20404 GNDA.n4366 GNDA.n4326 0.0682083
R20405 GNDA.n4376 GNDA.n4324 0.0682083
R20406 GNDA.n4378 GNDA.n4377 0.0682083
R20407 GNDA.n4388 GNDA.n4387 0.0682083
R20408 GNDA.n4396 GNDA.n4320 0.0682083
R20409 GNDA.n4406 GNDA.n4318 0.0682083
R20410 GNDA.n4408 GNDA.n4407 0.0682083
R20411 GNDA.n4418 GNDA.n4417 0.0682083
R20412 GNDA.n4426 GNDA.n4314 0.0682083
R20413 GNDA.n4436 GNDA.n4312 0.0682083
R20414 GNDA.n4438 GNDA.n4437 0.0682083
R20415 GNDA.n4170 GNDA.n4166 0.0682083
R20416 GNDA.n4180 GNDA.n1646 0.0682083
R20417 GNDA.n4182 GNDA.n4181 0.0682083
R20418 GNDA.n4192 GNDA.n4191 0.0682083
R20419 GNDA.n4200 GNDA.n1642 0.0682083
R20420 GNDA.n4210 GNDA.n1640 0.0682083
R20421 GNDA.n4212 GNDA.n4211 0.0682083
R20422 GNDA.n4222 GNDA.n4221 0.0682083
R20423 GNDA.n4230 GNDA.n1636 0.0682083
R20424 GNDA.n4240 GNDA.n1634 0.0682083
R20425 GNDA.n4242 GNDA.n4241 0.0682083
R20426 GNDA.n4252 GNDA.n4251 0.0682083
R20427 GNDA.n4260 GNDA.n1630 0.0682083
R20428 GNDA.n4270 GNDA.n1628 0.0682083
R20429 GNDA.n4272 GNDA.n4271 0.0682083
R20430 GNDA.n1813 GNDA.n1649 0.0682083
R20431 GNDA.n1699 GNDA.n1698 0.0682083
R20432 GNDA.n1701 GNDA.n1700 0.0682083
R20433 GNDA.n1705 GNDA.n1704 0.0682083
R20434 GNDA.n1707 GNDA.n1706 0.0682083
R20435 GNDA.n1711 GNDA.n1710 0.0682083
R20436 GNDA.n1713 GNDA.n1712 0.0682083
R20437 GNDA.n1717 GNDA.n1716 0.0682083
R20438 GNDA.n1719 GNDA.n1718 0.0682083
R20439 GNDA.n1723 GNDA.n1722 0.0682083
R20440 GNDA.n1725 GNDA.n1724 0.0682083
R20441 GNDA.n1729 GNDA.n1728 0.0682083
R20442 GNDA.n1731 GNDA.n1730 0.0682083
R20443 GNDA.n1735 GNDA.n1734 0.0682083
R20444 GNDA.n1737 GNDA.n1736 0.0682083
R20445 GNDA.n3827 GNDA.n3823 0.0682083
R20446 GNDA.n3837 GNDA.n3821 0.0682083
R20447 GNDA.n3839 GNDA.n3838 0.0682083
R20448 GNDA.n3849 GNDA.n3848 0.0682083
R20449 GNDA.n3857 GNDA.n3817 0.0682083
R20450 GNDA.n3867 GNDA.n3815 0.0682083
R20451 GNDA.n3869 GNDA.n3868 0.0682083
R20452 GNDA.n3879 GNDA.n3878 0.0682083
R20453 GNDA.n3887 GNDA.n3811 0.0682083
R20454 GNDA.n3897 GNDA.n3809 0.0682083
R20455 GNDA.n3899 GNDA.n3898 0.0682083
R20456 GNDA.n3909 GNDA.n3908 0.0682083
R20457 GNDA.n3917 GNDA.n3805 0.0682083
R20458 GNDA.n3927 GNDA.n3803 0.0682083
R20459 GNDA.n3929 GNDA.n3928 0.0682083
R20460 GNDA.n4080 GNDA.n1835 0.0682083
R20461 GNDA.n3974 GNDA.n3963 0.0682083
R20462 GNDA.n3976 GNDA.n3975 0.0682083
R20463 GNDA.n3986 GNDA.n3985 0.0682083
R20464 GNDA.n3994 GNDA.n3959 0.0682083
R20465 GNDA.n4004 GNDA.n3957 0.0682083
R20466 GNDA.n4006 GNDA.n4005 0.0682083
R20467 GNDA.n4016 GNDA.n4015 0.0682083
R20468 GNDA.n4024 GNDA.n3953 0.0682083
R20469 GNDA.n4034 GNDA.n3951 0.0682083
R20470 GNDA.n4036 GNDA.n4035 0.0682083
R20471 GNDA.n4046 GNDA.n4045 0.0682083
R20472 GNDA.n4054 GNDA.n3947 0.0682083
R20473 GNDA.n4064 GNDA.n3945 0.0682083
R20474 GNDA.n4066 GNDA.n4065 0.0682083
R20475 GNDA.n3472 GNDA.n3468 0.0682083
R20476 GNDA.n3482 GNDA.n1885 0.0682083
R20477 GNDA.n3484 GNDA.n3483 0.0682083
R20478 GNDA.n3494 GNDA.n3493 0.0682083
R20479 GNDA.n3502 GNDA.n1881 0.0682083
R20480 GNDA.n3512 GNDA.n1879 0.0682083
R20481 GNDA.n3514 GNDA.n3513 0.0682083
R20482 GNDA.n3524 GNDA.n3523 0.0682083
R20483 GNDA.n3532 GNDA.n1875 0.0682083
R20484 GNDA.n3542 GNDA.n1873 0.0682083
R20485 GNDA.n3544 GNDA.n3543 0.0682083
R20486 GNDA.n3554 GNDA.n3553 0.0682083
R20487 GNDA.n3562 GNDA.n1869 0.0682083
R20488 GNDA.n3572 GNDA.n1867 0.0682083
R20489 GNDA.n3574 GNDA.n3573 0.0682083
R20490 GNDA.n2537 GNDA.n1887 0.0682083
R20491 GNDA.n2547 GNDA.n2532 0.0682083
R20492 GNDA.n2549 GNDA.n2548 0.0682083
R20493 GNDA.n2559 GNDA.n2558 0.0682083
R20494 GNDA.n2567 GNDA.n2528 0.0682083
R20495 GNDA.n2577 GNDA.n2526 0.0682083
R20496 GNDA.n2579 GNDA.n2578 0.0682083
R20497 GNDA.n2589 GNDA.n2588 0.0682083
R20498 GNDA.n2597 GNDA.n2522 0.0682083
R20499 GNDA.n2607 GNDA.n2520 0.0682083
R20500 GNDA.n2609 GNDA.n2608 0.0682083
R20501 GNDA.n2619 GNDA.n2618 0.0682083
R20502 GNDA.n2627 GNDA.n2516 0.0682083
R20503 GNDA.n2637 GNDA.n2514 0.0682083
R20504 GNDA.n2639 GNDA.n2638 0.0682083
R20505 GNDA.n2820 GNDA.n1889 0.0682083
R20506 GNDA.n2830 GNDA.n2815 0.0682083
R20507 GNDA.n2832 GNDA.n2831 0.0682083
R20508 GNDA.n2842 GNDA.n2841 0.0682083
R20509 GNDA.n2850 GNDA.n2811 0.0682083
R20510 GNDA.n2860 GNDA.n2809 0.0682083
R20511 GNDA.n2862 GNDA.n2861 0.0682083
R20512 GNDA.n2872 GNDA.n2871 0.0682083
R20513 GNDA.n2880 GNDA.n2805 0.0682083
R20514 GNDA.n2890 GNDA.n2803 0.0682083
R20515 GNDA.n2892 GNDA.n2891 0.0682083
R20516 GNDA.n2902 GNDA.n2901 0.0682083
R20517 GNDA.n2910 GNDA.n2799 0.0682083
R20518 GNDA.n2920 GNDA.n2797 0.0682083
R20519 GNDA.n2922 GNDA.n2921 0.0682083
R20520 GNDA.n2961 GNDA.n1890 0.0682083
R20521 GNDA.n2971 GNDA.n2956 0.0682083
R20522 GNDA.n2973 GNDA.n2972 0.0682083
R20523 GNDA.n2983 GNDA.n2982 0.0682083
R20524 GNDA.n2991 GNDA.n2952 0.0682083
R20525 GNDA.n3001 GNDA.n2950 0.0682083
R20526 GNDA.n3003 GNDA.n3002 0.0682083
R20527 GNDA.n3013 GNDA.n3012 0.0682083
R20528 GNDA.n3021 GNDA.n2946 0.0682083
R20529 GNDA.n3031 GNDA.n2944 0.0682083
R20530 GNDA.n3033 GNDA.n3032 0.0682083
R20531 GNDA.n3043 GNDA.n3042 0.0682083
R20532 GNDA.n3051 GNDA.n2940 0.0682083
R20533 GNDA.n3061 GNDA.n2938 0.0682083
R20534 GNDA.n3063 GNDA.n3062 0.0682083
R20535 GNDA.n3102 GNDA.n1891 0.0682083
R20536 GNDA.n3112 GNDA.n3097 0.0682083
R20537 GNDA.n3114 GNDA.n3113 0.0682083
R20538 GNDA.n3124 GNDA.n3123 0.0682083
R20539 GNDA.n3132 GNDA.n3093 0.0682083
R20540 GNDA.n3142 GNDA.n3091 0.0682083
R20541 GNDA.n3144 GNDA.n3143 0.0682083
R20542 GNDA.n3154 GNDA.n3153 0.0682083
R20543 GNDA.n3162 GNDA.n3087 0.0682083
R20544 GNDA.n3172 GNDA.n3085 0.0682083
R20545 GNDA.n3174 GNDA.n3173 0.0682083
R20546 GNDA.n3184 GNDA.n3183 0.0682083
R20547 GNDA.n3192 GNDA.n3081 0.0682083
R20548 GNDA.n3202 GNDA.n3079 0.0682083
R20549 GNDA.n3204 GNDA.n3203 0.0682083
R20550 GNDA.n3288 GNDA.n1892 0.0682083
R20551 GNDA.n3282 GNDA.n1897 0.0682083
R20552 GNDA.n3278 GNDA.n3277 0.0682083
R20553 GNDA.n3272 GNDA.n3271 0.0682083
R20554 GNDA.n3270 GNDA.n1907 0.0682083
R20555 GNDA.n3264 GNDA.n1912 0.0682083
R20556 GNDA.n3260 GNDA.n3259 0.0682083
R20557 GNDA.n3254 GNDA.n3253 0.0682083
R20558 GNDA.n3252 GNDA.n1922 0.0682083
R20559 GNDA.n3246 GNDA.n1927 0.0682083
R20560 GNDA.n3242 GNDA.n3241 0.0682083
R20561 GNDA.n3236 GNDA.n3235 0.0682083
R20562 GNDA.n3234 GNDA.n1937 0.0682083
R20563 GNDA.n3228 GNDA.n1942 0.0682083
R20564 GNDA.n3224 GNDA.n3223 0.0682083
R20565 GNDA.n2701 GNDA.n2697 0.0682083
R20566 GNDA.n2709 GNDA.n2693 0.0682083
R20567 GNDA.n2711 GNDA.n2710 0.0682083
R20568 GNDA.n2719 GNDA.n2718 0.0682083
R20569 GNDA.n2725 GNDA.n2685 0.0682083
R20570 GNDA.n2733 GNDA.n2681 0.0682083
R20571 GNDA.n2735 GNDA.n2734 0.0682083
R20572 GNDA.n2743 GNDA.n2742 0.0682083
R20573 GNDA.n2749 GNDA.n2673 0.0682083
R20574 GNDA.n2757 GNDA.n2669 0.0682083
R20575 GNDA.n2759 GNDA.n2758 0.0682083
R20576 GNDA.n2767 GNDA.n2766 0.0682083
R20577 GNDA.n2773 GNDA.n2661 0.0682083
R20578 GNDA.n2781 GNDA.n2657 0.0682083
R20579 GNDA.n2783 GNDA.n2782 0.0682083
R20580 GNDA.n4773 GNDA.n4640 0.0672139
R20581 GNDA.n5800 GNDA.n5663 0.0672139
R20582 GNDA.n6078 GNDA.n5945 0.0672139
R20583 GNDA.n1514 GNDA.n1469 0.0672139
R20584 GNDA.n3749 GNDA.n3611 0.0672139
R20585 GNDA.n3386 GNDA.n3341 0.0672139
R20586 GNDA.n5229 GNDA.n5096 0.0672139
R20587 GNDA.n5326 GNDA.n5281 0.0672139
R20588 GNDA.n5517 GNDA.n5046 0.0672139
R20589 GNDA.n5659 GNDA.n5521 0.0672139
R20590 GNDA.n5941 GNDA.n5804 0.0672139
R20591 GNDA.n4922 GNDA.n1397 0.0672139
R20592 GNDA.n4636 GNDA.n4498 0.0672139
R20593 GNDA.n4447 GNDA.n4309 0.0672139
R20594 GNDA.n4281 GNDA.n1625 0.0672139
R20595 GNDA.n1740 GNDA.n1695 0.0672139
R20596 GNDA.n3938 GNDA.n3800 0.0672139
R20597 GNDA.n4075 GNDA.n3942 0.0672139
R20598 GNDA.n3583 GNDA.n1864 0.0672139
R20599 GNDA.n2648 GNDA.n2511 0.0672139
R20600 GNDA.n2931 GNDA.n2794 0.0672139
R20601 GNDA.n3072 GNDA.n2935 0.0672139
R20602 GNDA.n3213 GNDA.n3076 0.0672139
R20603 GNDA.n3219 GNDA.n3218 0.0672139
R20604 GNDA.n2790 GNDA.n2652 0.0672139
R20605 GNDA.n6355 GNDA.n6353 0.0667303
R20606 GNDA.n412 GNDA.n411 0.0667303
R20607 GNDA.n6615 GNDA.n6286 0.0646844
R20608 GNDA.n4673 GNDA.n4672 0.063
R20609 GNDA.n4684 GNDA.n4657 0.063
R20610 GNDA.n4703 GNDA.n4702 0.063
R20611 GNDA.n4714 GNDA.n4651 0.063
R20612 GNDA.n4733 GNDA.n4732 0.063
R20613 GNDA.n4744 GNDA.n4645 0.063
R20614 GNDA.n4763 GNDA.n4762 0.063
R20615 GNDA.n5700 GNDA.n5699 0.063
R20616 GNDA.n5711 GNDA.n5680 0.063
R20617 GNDA.n5730 GNDA.n5729 0.063
R20618 GNDA.n5741 GNDA.n5674 0.063
R20619 GNDA.n5760 GNDA.n5759 0.063
R20620 GNDA.n5771 GNDA.n5668 0.063
R20621 GNDA.n5790 GNDA.n5789 0.063
R20622 GNDA.n5978 GNDA.n5977 0.063
R20623 GNDA.n5989 GNDA.n5962 0.063
R20624 GNDA.n6008 GNDA.n6007 0.063
R20625 GNDA.n6019 GNDA.n5956 0.063
R20626 GNDA.n6038 GNDA.n6037 0.063
R20627 GNDA.n6049 GNDA.n5950 0.063
R20628 GNDA.n6068 GNDA.n6067 0.063
R20629 GNDA.n1474 GNDA.n1473 0.063
R20630 GNDA.n1480 GNDA.n1479 0.063
R20631 GNDA.n1486 GNDA.n1485 0.063
R20632 GNDA.n1492 GNDA.n1491 0.063
R20633 GNDA.n1498 GNDA.n1497 0.063
R20634 GNDA.n1504 GNDA.n1503 0.063
R20635 GNDA.n1510 GNDA.n1509 0.063
R20636 GNDA.n3649 GNDA.n3648 0.063
R20637 GNDA.n3660 GNDA.n3628 0.063
R20638 GNDA.n3679 GNDA.n3678 0.063
R20639 GNDA.n3690 GNDA.n3622 0.063
R20640 GNDA.n3709 GNDA.n3708 0.063
R20641 GNDA.n3720 GNDA.n3616 0.063
R20642 GNDA.n3739 GNDA.n3738 0.063
R20643 GNDA.n3346 GNDA.n3345 0.063
R20644 GNDA.n3352 GNDA.n3351 0.063
R20645 GNDA.n3358 GNDA.n3357 0.063
R20646 GNDA.n3364 GNDA.n3363 0.063
R20647 GNDA.n3370 GNDA.n3369 0.063
R20648 GNDA.n3376 GNDA.n3375 0.063
R20649 GNDA.n3382 GNDA.n3381 0.063
R20650 GNDA.n5129 GNDA.n5128 0.063
R20651 GNDA.n5140 GNDA.n5113 0.063
R20652 GNDA.n5159 GNDA.n5158 0.063
R20653 GNDA.n5170 GNDA.n5107 0.063
R20654 GNDA.n5189 GNDA.n5188 0.063
R20655 GNDA.n5200 GNDA.n5101 0.063
R20656 GNDA.n5219 GNDA.n5218 0.063
R20657 GNDA.n5286 GNDA.n5285 0.063
R20658 GNDA.n5292 GNDA.n5291 0.063
R20659 GNDA.n5298 GNDA.n5297 0.063
R20660 GNDA.n5304 GNDA.n5303 0.063
R20661 GNDA.n5310 GNDA.n5309 0.063
R20662 GNDA.n5316 GNDA.n5315 0.063
R20663 GNDA.n5322 GNDA.n5321 0.063
R20664 GNDA.n5417 GNDA.n5416 0.063
R20665 GNDA.n5428 GNDA.n5063 0.063
R20666 GNDA.n5447 GNDA.n5446 0.063
R20667 GNDA.n5458 GNDA.n5057 0.063
R20668 GNDA.n5477 GNDA.n5476 0.063
R20669 GNDA.n5488 GNDA.n5051 0.063
R20670 GNDA.n5507 GNDA.n5506 0.063
R20671 GNDA.n5559 GNDA.n5558 0.063
R20672 GNDA.n5570 GNDA.n5538 0.063
R20673 GNDA.n5589 GNDA.n5588 0.063
R20674 GNDA.n5600 GNDA.n5532 0.063
R20675 GNDA.n5619 GNDA.n5618 0.063
R20676 GNDA.n5630 GNDA.n5526 0.063
R20677 GNDA.n5649 GNDA.n5648 0.063
R20678 GNDA.n5841 GNDA.n5840 0.063
R20679 GNDA.n5852 GNDA.n5821 0.063
R20680 GNDA.n5871 GNDA.n5870 0.063
R20681 GNDA.n5882 GNDA.n5815 0.063
R20682 GNDA.n5901 GNDA.n5900 0.063
R20683 GNDA.n5912 GNDA.n5809 0.063
R20684 GNDA.n5931 GNDA.n5930 0.063
R20685 GNDA.n4822 GNDA.n4821 0.063
R20686 GNDA.n4833 GNDA.n1414 0.063
R20687 GNDA.n4852 GNDA.n4851 0.063
R20688 GNDA.n4863 GNDA.n1408 0.063
R20689 GNDA.n4882 GNDA.n4881 0.063
R20690 GNDA.n4893 GNDA.n1402 0.063
R20691 GNDA.n4912 GNDA.n4911 0.063
R20692 GNDA.n4536 GNDA.n4535 0.063
R20693 GNDA.n4547 GNDA.n4515 0.063
R20694 GNDA.n4566 GNDA.n4565 0.063
R20695 GNDA.n4577 GNDA.n4509 0.063
R20696 GNDA.n4596 GNDA.n4595 0.063
R20697 GNDA.n4607 GNDA.n4503 0.063
R20698 GNDA.n4626 GNDA.n4625 0.063
R20699 GNDA.n4347 GNDA.n4346 0.063
R20700 GNDA.n4358 GNDA.n4326 0.063
R20701 GNDA.n4377 GNDA.n4376 0.063
R20702 GNDA.n4388 GNDA.n4320 0.063
R20703 GNDA.n4407 GNDA.n4406 0.063
R20704 GNDA.n4418 GNDA.n4314 0.063
R20705 GNDA.n4437 GNDA.n4436 0.063
R20706 GNDA.n4181 GNDA.n4180 0.063
R20707 GNDA.n4192 GNDA.n1642 0.063
R20708 GNDA.n4211 GNDA.n4210 0.063
R20709 GNDA.n4222 GNDA.n1636 0.063
R20710 GNDA.n4241 GNDA.n4240 0.063
R20711 GNDA.n4252 GNDA.n1630 0.063
R20712 GNDA.n4271 GNDA.n4270 0.063
R20713 GNDA.n1700 GNDA.n1699 0.063
R20714 GNDA.n1706 GNDA.n1705 0.063
R20715 GNDA.n1712 GNDA.n1711 0.063
R20716 GNDA.n1718 GNDA.n1717 0.063
R20717 GNDA.n1724 GNDA.n1723 0.063
R20718 GNDA.n1730 GNDA.n1729 0.063
R20719 GNDA.n1736 GNDA.n1735 0.063
R20720 GNDA.n3838 GNDA.n3837 0.063
R20721 GNDA.n3849 GNDA.n3817 0.063
R20722 GNDA.n3868 GNDA.n3867 0.063
R20723 GNDA.n3879 GNDA.n3811 0.063
R20724 GNDA.n3898 GNDA.n3897 0.063
R20725 GNDA.n3909 GNDA.n3805 0.063
R20726 GNDA.n3928 GNDA.n3927 0.063
R20727 GNDA.n3975 GNDA.n3974 0.063
R20728 GNDA.n3986 GNDA.n3959 0.063
R20729 GNDA.n4005 GNDA.n4004 0.063
R20730 GNDA.n4016 GNDA.n3953 0.063
R20731 GNDA.n4035 GNDA.n4034 0.063
R20732 GNDA.n4046 GNDA.n3947 0.063
R20733 GNDA.n4065 GNDA.n4064 0.063
R20734 GNDA.n3483 GNDA.n3482 0.063
R20735 GNDA.n3494 GNDA.n1881 0.063
R20736 GNDA.n3513 GNDA.n3512 0.063
R20737 GNDA.n3524 GNDA.n1875 0.063
R20738 GNDA.n3543 GNDA.n3542 0.063
R20739 GNDA.n3554 GNDA.n1869 0.063
R20740 GNDA.n3573 GNDA.n3572 0.063
R20741 GNDA.n2548 GNDA.n2547 0.063
R20742 GNDA.n2559 GNDA.n2528 0.063
R20743 GNDA.n2578 GNDA.n2577 0.063
R20744 GNDA.n2589 GNDA.n2522 0.063
R20745 GNDA.n2608 GNDA.n2607 0.063
R20746 GNDA.n2619 GNDA.n2516 0.063
R20747 GNDA.n2638 GNDA.n2637 0.063
R20748 GNDA.n2831 GNDA.n2830 0.063
R20749 GNDA.n2842 GNDA.n2811 0.063
R20750 GNDA.n2861 GNDA.n2860 0.063
R20751 GNDA.n2872 GNDA.n2805 0.063
R20752 GNDA.n2891 GNDA.n2890 0.063
R20753 GNDA.n2902 GNDA.n2799 0.063
R20754 GNDA.n2921 GNDA.n2920 0.063
R20755 GNDA.n2972 GNDA.n2971 0.063
R20756 GNDA.n2983 GNDA.n2952 0.063
R20757 GNDA.n3002 GNDA.n3001 0.063
R20758 GNDA.n3013 GNDA.n2946 0.063
R20759 GNDA.n3032 GNDA.n3031 0.063
R20760 GNDA.n3043 GNDA.n2940 0.063
R20761 GNDA.n3062 GNDA.n3061 0.063
R20762 GNDA.n3113 GNDA.n3112 0.063
R20763 GNDA.n3124 GNDA.n3093 0.063
R20764 GNDA.n3143 GNDA.n3142 0.063
R20765 GNDA.n3154 GNDA.n3087 0.063
R20766 GNDA.n3173 GNDA.n3172 0.063
R20767 GNDA.n3184 GNDA.n3081 0.063
R20768 GNDA.n3203 GNDA.n3202 0.063
R20769 GNDA.n3278 GNDA.n1897 0.063
R20770 GNDA.n3271 GNDA.n3270 0.063
R20771 GNDA.n3260 GNDA.n1912 0.063
R20772 GNDA.n3253 GNDA.n3252 0.063
R20773 GNDA.n3242 GNDA.n1927 0.063
R20774 GNDA.n3235 GNDA.n3234 0.063
R20775 GNDA.n3224 GNDA.n1942 0.063
R20776 GNDA.n2710 GNDA.n2709 0.063
R20777 GNDA.n2719 GNDA.n2685 0.063
R20778 GNDA.n2734 GNDA.n2733 0.063
R20779 GNDA.n2743 GNDA.n2673 0.063
R20780 GNDA.n2758 GNDA.n2757 0.063
R20781 GNDA.n2767 GNDA.n2661 0.063
R20782 GNDA.n2782 GNDA.n2781 0.063
R20783 GNDA.n6278 GNDA.n6277 0.063
R20784 GNDA.n4666 GNDA.n4665 0.0553333
R20785 GNDA.n4680 GNDA.n4679 0.0553333
R20786 GNDA.n4696 GNDA.n4695 0.0553333
R20787 GNDA.n4710 GNDA.n4709 0.0553333
R20788 GNDA.n4726 GNDA.n4725 0.0553333
R20789 GNDA.n4740 GNDA.n4739 0.0553333
R20790 GNDA.n4756 GNDA.n4755 0.0553333
R20791 GNDA.n4770 GNDA.n4769 0.0553333
R20792 GNDA.n5693 GNDA.n5692 0.0553333
R20793 GNDA.n5707 GNDA.n5706 0.0553333
R20794 GNDA.n5723 GNDA.n5722 0.0553333
R20795 GNDA.n5737 GNDA.n5736 0.0553333
R20796 GNDA.n5753 GNDA.n5752 0.0553333
R20797 GNDA.n5767 GNDA.n5766 0.0553333
R20798 GNDA.n5783 GNDA.n5782 0.0553333
R20799 GNDA.n5797 GNDA.n5796 0.0553333
R20800 GNDA.n2696 GNDA.n2695 0.0553333
R20801 GNDA.n2715 GNDA.n2714 0.0553333
R20802 GNDA.n2684 GNDA.n2683 0.0553333
R20803 GNDA.n2739 GNDA.n2738 0.0553333
R20804 GNDA.n2672 GNDA.n2671 0.0553333
R20805 GNDA.n2763 GNDA.n2762 0.0553333
R20806 GNDA.n2660 GNDA.n2659 0.0553333
R20807 GNDA.n2787 GNDA.n2786 0.0553333
R20808 GNDA.n5971 GNDA.n5970 0.0553333
R20809 GNDA.n5985 GNDA.n5984 0.0553333
R20810 GNDA.n6001 GNDA.n6000 0.0553333
R20811 GNDA.n6015 GNDA.n6014 0.0553333
R20812 GNDA.n6031 GNDA.n6030 0.0553333
R20813 GNDA.n6045 GNDA.n6044 0.0553333
R20814 GNDA.n6061 GNDA.n6060 0.0553333
R20815 GNDA.n6075 GNDA.n6074 0.0553333
R20816 GNDA.n1582 GNDA.n1581 0.0553333
R20817 GNDA.n1573 GNDA.n1572 0.0553333
R20818 GNDA.n1564 GNDA.n1563 0.0553333
R20819 GNDA.n1555 GNDA.n1554 0.0553333
R20820 GNDA.n1546 GNDA.n1545 0.0553333
R20821 GNDA.n1537 GNDA.n1536 0.0553333
R20822 GNDA.n1528 GNDA.n1527 0.0553333
R20823 GNDA.n1519 GNDA.n1518 0.0553333
R20824 GNDA.n3642 GNDA.n3641 0.0553333
R20825 GNDA.n3656 GNDA.n3655 0.0553333
R20826 GNDA.n3672 GNDA.n3671 0.0553333
R20827 GNDA.n3686 GNDA.n3685 0.0553333
R20828 GNDA.n3702 GNDA.n3701 0.0553333
R20829 GNDA.n3716 GNDA.n3715 0.0553333
R20830 GNDA.n3732 GNDA.n3731 0.0553333
R20831 GNDA.n3746 GNDA.n3745 0.0553333
R20832 GNDA.n3454 GNDA.n3453 0.0553333
R20833 GNDA.n3445 GNDA.n3444 0.0553333
R20834 GNDA.n3436 GNDA.n3435 0.0553333
R20835 GNDA.n3427 GNDA.n3426 0.0553333
R20836 GNDA.n3418 GNDA.n3417 0.0553333
R20837 GNDA.n3409 GNDA.n3408 0.0553333
R20838 GNDA.n3400 GNDA.n3399 0.0553333
R20839 GNDA.n3391 GNDA.n3390 0.0553333
R20840 GNDA.n5122 GNDA.n5121 0.0553333
R20841 GNDA.n5136 GNDA.n5135 0.0553333
R20842 GNDA.n5152 GNDA.n5151 0.0553333
R20843 GNDA.n5166 GNDA.n5165 0.0553333
R20844 GNDA.n5182 GNDA.n5181 0.0553333
R20845 GNDA.n5196 GNDA.n5195 0.0553333
R20846 GNDA.n5212 GNDA.n5211 0.0553333
R20847 GNDA.n5226 GNDA.n5225 0.0553333
R20848 GNDA.n5394 GNDA.n5393 0.0553333
R20849 GNDA.n5385 GNDA.n5384 0.0553333
R20850 GNDA.n5376 GNDA.n5375 0.0553333
R20851 GNDA.n5367 GNDA.n5366 0.0553333
R20852 GNDA.n5358 GNDA.n5357 0.0553333
R20853 GNDA.n5349 GNDA.n5348 0.0553333
R20854 GNDA.n5340 GNDA.n5339 0.0553333
R20855 GNDA.n5331 GNDA.n5330 0.0553333
R20856 GNDA.n5410 GNDA.n5409 0.0553333
R20857 GNDA.n5424 GNDA.n5423 0.0553333
R20858 GNDA.n5440 GNDA.n5439 0.0553333
R20859 GNDA.n5454 GNDA.n5453 0.0553333
R20860 GNDA.n5470 GNDA.n5469 0.0553333
R20861 GNDA.n5484 GNDA.n5483 0.0553333
R20862 GNDA.n5500 GNDA.n5499 0.0553333
R20863 GNDA.n5514 GNDA.n5513 0.0553333
R20864 GNDA.n5552 GNDA.n5551 0.0553333
R20865 GNDA.n5566 GNDA.n5565 0.0553333
R20866 GNDA.n5582 GNDA.n5581 0.0553333
R20867 GNDA.n5596 GNDA.n5595 0.0553333
R20868 GNDA.n5612 GNDA.n5611 0.0553333
R20869 GNDA.n5626 GNDA.n5625 0.0553333
R20870 GNDA.n5642 GNDA.n5641 0.0553333
R20871 GNDA.n5656 GNDA.n5655 0.0553333
R20872 GNDA.n5834 GNDA.n5833 0.0553333
R20873 GNDA.n5848 GNDA.n5847 0.0553333
R20874 GNDA.n5864 GNDA.n5863 0.0553333
R20875 GNDA.n5878 GNDA.n5877 0.0553333
R20876 GNDA.n5894 GNDA.n5893 0.0553333
R20877 GNDA.n5908 GNDA.n5907 0.0553333
R20878 GNDA.n5924 GNDA.n5923 0.0553333
R20879 GNDA.n5938 GNDA.n5937 0.0553333
R20880 GNDA.n4815 GNDA.n4814 0.0553333
R20881 GNDA.n4829 GNDA.n4828 0.0553333
R20882 GNDA.n4845 GNDA.n4844 0.0553333
R20883 GNDA.n4859 GNDA.n4858 0.0553333
R20884 GNDA.n4875 GNDA.n4874 0.0553333
R20885 GNDA.n4889 GNDA.n4888 0.0553333
R20886 GNDA.n4905 GNDA.n4904 0.0553333
R20887 GNDA.n4919 GNDA.n4918 0.0553333
R20888 GNDA.n4529 GNDA.n4528 0.0553333
R20889 GNDA.n4543 GNDA.n4542 0.0553333
R20890 GNDA.n4559 GNDA.n4558 0.0553333
R20891 GNDA.n4573 GNDA.n4572 0.0553333
R20892 GNDA.n4589 GNDA.n4588 0.0553333
R20893 GNDA.n4603 GNDA.n4602 0.0553333
R20894 GNDA.n4619 GNDA.n4618 0.0553333
R20895 GNDA.n4633 GNDA.n4632 0.0553333
R20896 GNDA.n4340 GNDA.n4339 0.0553333
R20897 GNDA.n4354 GNDA.n4353 0.0553333
R20898 GNDA.n4370 GNDA.n4369 0.0553333
R20899 GNDA.n4384 GNDA.n4383 0.0553333
R20900 GNDA.n4400 GNDA.n4399 0.0553333
R20901 GNDA.n4414 GNDA.n4413 0.0553333
R20902 GNDA.n4430 GNDA.n4429 0.0553333
R20903 GNDA.n4444 GNDA.n4443 0.0553333
R20904 GNDA.n4174 GNDA.n4173 0.0553333
R20905 GNDA.n4188 GNDA.n4187 0.0553333
R20906 GNDA.n4204 GNDA.n4203 0.0553333
R20907 GNDA.n4218 GNDA.n4217 0.0553333
R20908 GNDA.n4234 GNDA.n4233 0.0553333
R20909 GNDA.n4248 GNDA.n4247 0.0553333
R20910 GNDA.n4264 GNDA.n4263 0.0553333
R20911 GNDA.n4278 GNDA.n4277 0.0553333
R20912 GNDA.n1808 GNDA.n1807 0.0553333
R20913 GNDA.n1799 GNDA.n1798 0.0553333
R20914 GNDA.n1790 GNDA.n1789 0.0553333
R20915 GNDA.n1781 GNDA.n1780 0.0553333
R20916 GNDA.n1772 GNDA.n1771 0.0553333
R20917 GNDA.n1763 GNDA.n1762 0.0553333
R20918 GNDA.n1754 GNDA.n1753 0.0553333
R20919 GNDA.n1745 GNDA.n1744 0.0553333
R20920 GNDA.n3831 GNDA.n3830 0.0553333
R20921 GNDA.n3845 GNDA.n3844 0.0553333
R20922 GNDA.n3861 GNDA.n3860 0.0553333
R20923 GNDA.n3875 GNDA.n3874 0.0553333
R20924 GNDA.n3891 GNDA.n3890 0.0553333
R20925 GNDA.n3905 GNDA.n3904 0.0553333
R20926 GNDA.n3921 GNDA.n3920 0.0553333
R20927 GNDA.n3935 GNDA.n3934 0.0553333
R20928 GNDA.n3968 GNDA.n3967 0.0553333
R20929 GNDA.n3982 GNDA.n3981 0.0553333
R20930 GNDA.n3998 GNDA.n3997 0.0553333
R20931 GNDA.n4012 GNDA.n4011 0.0553333
R20932 GNDA.n4028 GNDA.n4027 0.0553333
R20933 GNDA.n4042 GNDA.n4041 0.0553333
R20934 GNDA.n4058 GNDA.n4057 0.0553333
R20935 GNDA.n4072 GNDA.n4071 0.0553333
R20936 GNDA.n3476 GNDA.n3475 0.0553333
R20937 GNDA.n3490 GNDA.n3489 0.0553333
R20938 GNDA.n3506 GNDA.n3505 0.0553333
R20939 GNDA.n3520 GNDA.n3519 0.0553333
R20940 GNDA.n3536 GNDA.n3535 0.0553333
R20941 GNDA.n3550 GNDA.n3549 0.0553333
R20942 GNDA.n3566 GNDA.n3565 0.0553333
R20943 GNDA.n3580 GNDA.n3579 0.0553333
R20944 GNDA.n2541 GNDA.n2540 0.0553333
R20945 GNDA.n2555 GNDA.n2554 0.0553333
R20946 GNDA.n2571 GNDA.n2570 0.0553333
R20947 GNDA.n2585 GNDA.n2584 0.0553333
R20948 GNDA.n2601 GNDA.n2600 0.0553333
R20949 GNDA.n2615 GNDA.n2614 0.0553333
R20950 GNDA.n2631 GNDA.n2630 0.0553333
R20951 GNDA.n2645 GNDA.n2644 0.0553333
R20952 GNDA.n2824 GNDA.n2823 0.0553333
R20953 GNDA.n2838 GNDA.n2837 0.0553333
R20954 GNDA.n2854 GNDA.n2853 0.0553333
R20955 GNDA.n2868 GNDA.n2867 0.0553333
R20956 GNDA.n2884 GNDA.n2883 0.0553333
R20957 GNDA.n2898 GNDA.n2897 0.0553333
R20958 GNDA.n2914 GNDA.n2913 0.0553333
R20959 GNDA.n2928 GNDA.n2927 0.0553333
R20960 GNDA.n2965 GNDA.n2964 0.0553333
R20961 GNDA.n2979 GNDA.n2978 0.0553333
R20962 GNDA.n2995 GNDA.n2994 0.0553333
R20963 GNDA.n3009 GNDA.n3008 0.0553333
R20964 GNDA.n3025 GNDA.n3024 0.0553333
R20965 GNDA.n3039 GNDA.n3038 0.0553333
R20966 GNDA.n3055 GNDA.n3054 0.0553333
R20967 GNDA.n3069 GNDA.n3068 0.0553333
R20968 GNDA.n3106 GNDA.n3105 0.0553333
R20969 GNDA.n3120 GNDA.n3119 0.0553333
R20970 GNDA.n3136 GNDA.n3135 0.0553333
R20971 GNDA.n3150 GNDA.n3149 0.0553333
R20972 GNDA.n3166 GNDA.n3165 0.0553333
R20973 GNDA.n3180 GNDA.n3179 0.0553333
R20974 GNDA.n3196 GNDA.n3195 0.0553333
R20975 GNDA.n3210 GNDA.n3209 0.0553333
R20976 GNDA.n1895 GNDA.n1894 0.0553333
R20977 GNDA.n2357 GNDA.n1898 0.0553333
R20978 GNDA.n2360 GNDA.n1903 0.0553333
R20979 GNDA.n1905 GNDA.n1904 0.0553333
R20980 GNDA.n1910 GNDA.n1909 0.0553333
R20981 GNDA.n2366 GNDA.n1913 0.0553333
R20982 GNDA.n2369 GNDA.n1918 0.0553333
R20983 GNDA.n1920 GNDA.n1919 0.0553333
R20984 GNDA.n1925 GNDA.n1924 0.0553333
R20985 GNDA.n2375 GNDA.n1928 0.0553333
R20986 GNDA.n2378 GNDA.n1933 0.0553333
R20987 GNDA.n1935 GNDA.n1934 0.0553333
R20988 GNDA.n1940 GNDA.n1939 0.0553333
R20989 GNDA.n2384 GNDA.n1943 0.0553333
R20990 GNDA.n2387 GNDA.n1948 0.0553333
R20991 GNDA.n1950 GNDA.n1949 0.0553333
R20992 GNDA.n6358 GNDA.n6357 0.0553333
R20993 GNDA.n6347 GNDA.n6346 0.0553333
R20994 GNDA.n6382 GNDA.n6381 0.0553333
R20995 GNDA.n6335 GNDA.n6334 0.0553333
R20996 GNDA.n6406 GNDA.n6405 0.0553333
R20997 GNDA.n6323 GNDA.n6322 0.0553333
R20998 GNDA.n6430 GNDA.n6429 0.0553333
R20999 GNDA.n6444 GNDA.n6310 0.0553333
R21000 GNDA.n416 GNDA.n415 0.0553333
R21001 GNDA.n430 GNDA.n429 0.0553333
R21002 GNDA.n446 GNDA.n445 0.0553333
R21003 GNDA.n460 GNDA.n459 0.0553333
R21004 GNDA.n476 GNDA.n475 0.0553333
R21005 GNDA.n490 GNDA.n489 0.0553333
R21006 GNDA.n506 GNDA.n505 0.0553333
R21007 GNDA.n520 GNDA.n519 0.0553333
R21008 GNDA.n1316 GNDA 0.0517
R21009 GNDA.n6111 GNDA 0.0517
R21010 GNDA GNDA.n203 0.0517
R21011 GNDA.n793 GNDA 0.0517
R21012 GNDA GNDA.n6959 0.0517
R21013 GNDA GNDA.n7238 0.0517
R21014 GNDA.n6816 GNDA 0.0517
R21015 GNDA.n973 GNDA 0.0517
R21016 GNDA GNDA.n0 0.0517
R21017 GNDA.n4776 GNDA.n1598 0.0514167
R21018 GNDA.n4670 GNDA.n4669 0.0514167
R21019 GNDA.n4676 GNDA.n4675 0.0514167
R21020 GNDA.n4686 GNDA.n4685 0.0514167
R21021 GNDA.n4690 GNDA.n4689 0.0514167
R21022 GNDA.n4700 GNDA.n4699 0.0514167
R21023 GNDA.n4706 GNDA.n4705 0.0514167
R21024 GNDA.n4716 GNDA.n4715 0.0514167
R21025 GNDA.n4720 GNDA.n4719 0.0514167
R21026 GNDA.n4730 GNDA.n4729 0.0514167
R21027 GNDA.n4736 GNDA.n4735 0.0514167
R21028 GNDA.n4746 GNDA.n4745 0.0514167
R21029 GNDA.n4750 GNDA.n4749 0.0514167
R21030 GNDA.n4760 GNDA.n4759 0.0514167
R21031 GNDA.n4766 GNDA.n4765 0.0514167
R21032 GNDA.n4774 GNDA.n4639 0.0514167
R21033 GNDA.n5687 GNDA.n4972 0.0514167
R21034 GNDA.n5697 GNDA.n5696 0.0514167
R21035 GNDA.n5703 GNDA.n5702 0.0514167
R21036 GNDA.n5713 GNDA.n5712 0.0514167
R21037 GNDA.n5717 GNDA.n5716 0.0514167
R21038 GNDA.n5727 GNDA.n5726 0.0514167
R21039 GNDA.n5733 GNDA.n5732 0.0514167
R21040 GNDA.n5743 GNDA.n5742 0.0514167
R21041 GNDA.n5747 GNDA.n5746 0.0514167
R21042 GNDA.n5757 GNDA.n5756 0.0514167
R21043 GNDA.n5763 GNDA.n5762 0.0514167
R21044 GNDA.n5773 GNDA.n5772 0.0514167
R21045 GNDA.n5777 GNDA.n5776 0.0514167
R21046 GNDA.n5787 GNDA.n5786 0.0514167
R21047 GNDA.n5793 GNDA.n5792 0.0514167
R21048 GNDA.n5801 GNDA.n5662 0.0514167
R21049 GNDA.n2699 GNDA.n2462 0.0514167
R21050 GNDA.n2707 GNDA.n2706 0.0514167
R21051 GNDA.n2692 GNDA.n2691 0.0514167
R21052 GNDA.n2688 GNDA.n2687 0.0514167
R21053 GNDA.n2723 GNDA.n2722 0.0514167
R21054 GNDA.n2731 GNDA.n2730 0.0514167
R21055 GNDA.n2680 GNDA.n2679 0.0514167
R21056 GNDA.n2676 GNDA.n2675 0.0514167
R21057 GNDA.n2747 GNDA.n2746 0.0514167
R21058 GNDA.n2755 GNDA.n2754 0.0514167
R21059 GNDA.n2668 GNDA.n2667 0.0514167
R21060 GNDA.n2664 GNDA.n2663 0.0514167
R21061 GNDA.n2771 GNDA.n2770 0.0514167
R21062 GNDA.n2779 GNDA.n2778 0.0514167
R21063 GNDA.n2656 GNDA.n2655 0.0514167
R21064 GNDA.n2791 GNDA.n2651 0.0514167
R21065 GNDA.n6081 GNDA.n1370 0.0514167
R21066 GNDA.n5975 GNDA.n5974 0.0514167
R21067 GNDA.n5981 GNDA.n5980 0.0514167
R21068 GNDA.n5991 GNDA.n5990 0.0514167
R21069 GNDA.n5995 GNDA.n5994 0.0514167
R21070 GNDA.n6005 GNDA.n6004 0.0514167
R21071 GNDA.n6011 GNDA.n6010 0.0514167
R21072 GNDA.n6021 GNDA.n6020 0.0514167
R21073 GNDA.n6025 GNDA.n6024 0.0514167
R21074 GNDA.n6035 GNDA.n6034 0.0514167
R21075 GNDA.n6041 GNDA.n6040 0.0514167
R21076 GNDA.n6051 GNDA.n6050 0.0514167
R21077 GNDA.n6055 GNDA.n6054 0.0514167
R21078 GNDA.n6065 GNDA.n6064 0.0514167
R21079 GNDA.n6071 GNDA.n6070 0.0514167
R21080 GNDA.n6079 GNDA.n5944 0.0514167
R21081 GNDA.n1585 GNDA.n1584 0.0514167
R21082 GNDA.n1579 GNDA.n1578 0.0514167
R21083 GNDA.n1576 GNDA.n1575 0.0514167
R21084 GNDA.n1570 GNDA.n1569 0.0514167
R21085 GNDA.n1567 GNDA.n1566 0.0514167
R21086 GNDA.n1561 GNDA.n1560 0.0514167
R21087 GNDA.n1558 GNDA.n1557 0.0514167
R21088 GNDA.n1552 GNDA.n1551 0.0514167
R21089 GNDA.n1549 GNDA.n1548 0.0514167
R21090 GNDA.n1543 GNDA.n1542 0.0514167
R21091 GNDA.n1540 GNDA.n1539 0.0514167
R21092 GNDA.n1534 GNDA.n1533 0.0514167
R21093 GNDA.n1531 GNDA.n1530 0.0514167
R21094 GNDA.n1525 GNDA.n1524 0.0514167
R21095 GNDA.n1522 GNDA.n1521 0.0514167
R21096 GNDA.n1516 GNDA.n1515 0.0514167
R21097 GNDA.n3636 GNDA.n3586 0.0514167
R21098 GNDA.n3646 GNDA.n3645 0.0514167
R21099 GNDA.n3652 GNDA.n3651 0.0514167
R21100 GNDA.n3662 GNDA.n3661 0.0514167
R21101 GNDA.n3666 GNDA.n3665 0.0514167
R21102 GNDA.n3676 GNDA.n3675 0.0514167
R21103 GNDA.n3682 GNDA.n3681 0.0514167
R21104 GNDA.n3692 GNDA.n3691 0.0514167
R21105 GNDA.n3696 GNDA.n3695 0.0514167
R21106 GNDA.n3706 GNDA.n3705 0.0514167
R21107 GNDA.n3712 GNDA.n3711 0.0514167
R21108 GNDA.n3722 GNDA.n3721 0.0514167
R21109 GNDA.n3726 GNDA.n3725 0.0514167
R21110 GNDA.n3736 GNDA.n3735 0.0514167
R21111 GNDA.n3742 GNDA.n3741 0.0514167
R21112 GNDA.n3750 GNDA.n3610 0.0514167
R21113 GNDA.n3457 GNDA.n3456 0.0514167
R21114 GNDA.n3451 GNDA.n3450 0.0514167
R21115 GNDA.n3448 GNDA.n3447 0.0514167
R21116 GNDA.n3442 GNDA.n3441 0.0514167
R21117 GNDA.n3439 GNDA.n3438 0.0514167
R21118 GNDA.n3433 GNDA.n3432 0.0514167
R21119 GNDA.n3430 GNDA.n3429 0.0514167
R21120 GNDA.n3424 GNDA.n3423 0.0514167
R21121 GNDA.n3421 GNDA.n3420 0.0514167
R21122 GNDA.n3415 GNDA.n3414 0.0514167
R21123 GNDA.n3412 GNDA.n3411 0.0514167
R21124 GNDA.n3406 GNDA.n3405 0.0514167
R21125 GNDA.n3403 GNDA.n3402 0.0514167
R21126 GNDA.n3397 GNDA.n3396 0.0514167
R21127 GNDA.n3394 GNDA.n3393 0.0514167
R21128 GNDA.n3388 GNDA.n3387 0.0514167
R21129 GNDA.n5232 GNDA.n5071 0.0514167
R21130 GNDA.n5126 GNDA.n5125 0.0514167
R21131 GNDA.n5132 GNDA.n5131 0.0514167
R21132 GNDA.n5142 GNDA.n5141 0.0514167
R21133 GNDA.n5146 GNDA.n5145 0.0514167
R21134 GNDA.n5156 GNDA.n5155 0.0514167
R21135 GNDA.n5162 GNDA.n5161 0.0514167
R21136 GNDA.n5172 GNDA.n5171 0.0514167
R21137 GNDA.n5176 GNDA.n5175 0.0514167
R21138 GNDA.n5186 GNDA.n5185 0.0514167
R21139 GNDA.n5192 GNDA.n5191 0.0514167
R21140 GNDA.n5202 GNDA.n5201 0.0514167
R21141 GNDA.n5206 GNDA.n5205 0.0514167
R21142 GNDA.n5216 GNDA.n5215 0.0514167
R21143 GNDA.n5222 GNDA.n5221 0.0514167
R21144 GNDA.n5230 GNDA.n5095 0.0514167
R21145 GNDA.n5397 GNDA.n5396 0.0514167
R21146 GNDA.n5391 GNDA.n5390 0.0514167
R21147 GNDA.n5388 GNDA.n5387 0.0514167
R21148 GNDA.n5382 GNDA.n5381 0.0514167
R21149 GNDA.n5379 GNDA.n5378 0.0514167
R21150 GNDA.n5373 GNDA.n5372 0.0514167
R21151 GNDA.n5370 GNDA.n5369 0.0514167
R21152 GNDA.n5364 GNDA.n5363 0.0514167
R21153 GNDA.n5361 GNDA.n5360 0.0514167
R21154 GNDA.n5355 GNDA.n5354 0.0514167
R21155 GNDA.n5352 GNDA.n5351 0.0514167
R21156 GNDA.n5346 GNDA.n5345 0.0514167
R21157 GNDA.n5343 GNDA.n5342 0.0514167
R21158 GNDA.n5337 GNDA.n5336 0.0514167
R21159 GNDA.n5334 GNDA.n5333 0.0514167
R21160 GNDA.n5328 GNDA.n5327 0.0514167
R21161 GNDA.n5404 GNDA.n5020 0.0514167
R21162 GNDA.n5414 GNDA.n5413 0.0514167
R21163 GNDA.n5420 GNDA.n5419 0.0514167
R21164 GNDA.n5430 GNDA.n5429 0.0514167
R21165 GNDA.n5434 GNDA.n5433 0.0514167
R21166 GNDA.n5444 GNDA.n5443 0.0514167
R21167 GNDA.n5450 GNDA.n5449 0.0514167
R21168 GNDA.n5460 GNDA.n5459 0.0514167
R21169 GNDA.n5464 GNDA.n5463 0.0514167
R21170 GNDA.n5474 GNDA.n5473 0.0514167
R21171 GNDA.n5480 GNDA.n5479 0.0514167
R21172 GNDA.n5490 GNDA.n5489 0.0514167
R21173 GNDA.n5494 GNDA.n5493 0.0514167
R21174 GNDA.n5504 GNDA.n5503 0.0514167
R21175 GNDA.n5510 GNDA.n5509 0.0514167
R21176 GNDA.n5518 GNDA.n5045 0.0514167
R21177 GNDA.n5546 GNDA.n4996 0.0514167
R21178 GNDA.n5556 GNDA.n5555 0.0514167
R21179 GNDA.n5562 GNDA.n5561 0.0514167
R21180 GNDA.n5572 GNDA.n5571 0.0514167
R21181 GNDA.n5576 GNDA.n5575 0.0514167
R21182 GNDA.n5586 GNDA.n5585 0.0514167
R21183 GNDA.n5592 GNDA.n5591 0.0514167
R21184 GNDA.n5602 GNDA.n5601 0.0514167
R21185 GNDA.n5606 GNDA.n5605 0.0514167
R21186 GNDA.n5616 GNDA.n5615 0.0514167
R21187 GNDA.n5622 GNDA.n5621 0.0514167
R21188 GNDA.n5632 GNDA.n5631 0.0514167
R21189 GNDA.n5636 GNDA.n5635 0.0514167
R21190 GNDA.n5646 GNDA.n5645 0.0514167
R21191 GNDA.n5652 GNDA.n5651 0.0514167
R21192 GNDA.n5660 GNDA.n5520 0.0514167
R21193 GNDA.n5828 GNDA.n4948 0.0514167
R21194 GNDA.n5838 GNDA.n5837 0.0514167
R21195 GNDA.n5844 GNDA.n5843 0.0514167
R21196 GNDA.n5854 GNDA.n5853 0.0514167
R21197 GNDA.n5858 GNDA.n5857 0.0514167
R21198 GNDA.n5868 GNDA.n5867 0.0514167
R21199 GNDA.n5874 GNDA.n5873 0.0514167
R21200 GNDA.n5884 GNDA.n5883 0.0514167
R21201 GNDA.n5888 GNDA.n5887 0.0514167
R21202 GNDA.n5898 GNDA.n5897 0.0514167
R21203 GNDA.n5904 GNDA.n5903 0.0514167
R21204 GNDA.n5914 GNDA.n5913 0.0514167
R21205 GNDA.n5918 GNDA.n5917 0.0514167
R21206 GNDA.n5928 GNDA.n5927 0.0514167
R21207 GNDA.n5934 GNDA.n5933 0.0514167
R21208 GNDA.n5942 GNDA.n5803 0.0514167
R21209 GNDA.n4809 GNDA.n1372 0.0514167
R21210 GNDA.n4819 GNDA.n4818 0.0514167
R21211 GNDA.n4825 GNDA.n4824 0.0514167
R21212 GNDA.n4835 GNDA.n4834 0.0514167
R21213 GNDA.n4839 GNDA.n4838 0.0514167
R21214 GNDA.n4849 GNDA.n4848 0.0514167
R21215 GNDA.n4855 GNDA.n4854 0.0514167
R21216 GNDA.n4865 GNDA.n4864 0.0514167
R21217 GNDA.n4869 GNDA.n4868 0.0514167
R21218 GNDA.n4879 GNDA.n4878 0.0514167
R21219 GNDA.n4885 GNDA.n4884 0.0514167
R21220 GNDA.n4895 GNDA.n4894 0.0514167
R21221 GNDA.n4899 GNDA.n4898 0.0514167
R21222 GNDA.n4909 GNDA.n4908 0.0514167
R21223 GNDA.n4915 GNDA.n4914 0.0514167
R21224 GNDA.n4923 GNDA.n1396 0.0514167
R21225 GNDA.n4523 GNDA.n4473 0.0514167
R21226 GNDA.n4533 GNDA.n4532 0.0514167
R21227 GNDA.n4539 GNDA.n4538 0.0514167
R21228 GNDA.n4549 GNDA.n4548 0.0514167
R21229 GNDA.n4553 GNDA.n4552 0.0514167
R21230 GNDA.n4563 GNDA.n4562 0.0514167
R21231 GNDA.n4569 GNDA.n4568 0.0514167
R21232 GNDA.n4579 GNDA.n4578 0.0514167
R21233 GNDA.n4583 GNDA.n4582 0.0514167
R21234 GNDA.n4593 GNDA.n4592 0.0514167
R21235 GNDA.n4599 GNDA.n4598 0.0514167
R21236 GNDA.n4609 GNDA.n4608 0.0514167
R21237 GNDA.n4613 GNDA.n4612 0.0514167
R21238 GNDA.n4623 GNDA.n4622 0.0514167
R21239 GNDA.n4629 GNDA.n4628 0.0514167
R21240 GNDA.n4637 GNDA.n4497 0.0514167
R21241 GNDA.n4334 GNDA.n4284 0.0514167
R21242 GNDA.n4344 GNDA.n4343 0.0514167
R21243 GNDA.n4350 GNDA.n4349 0.0514167
R21244 GNDA.n4360 GNDA.n4359 0.0514167
R21245 GNDA.n4364 GNDA.n4363 0.0514167
R21246 GNDA.n4374 GNDA.n4373 0.0514167
R21247 GNDA.n4380 GNDA.n4379 0.0514167
R21248 GNDA.n4390 GNDA.n4389 0.0514167
R21249 GNDA.n4394 GNDA.n4393 0.0514167
R21250 GNDA.n4404 GNDA.n4403 0.0514167
R21251 GNDA.n4410 GNDA.n4409 0.0514167
R21252 GNDA.n4420 GNDA.n4419 0.0514167
R21253 GNDA.n4424 GNDA.n4423 0.0514167
R21254 GNDA.n4434 GNDA.n4433 0.0514167
R21255 GNDA.n4440 GNDA.n4439 0.0514167
R21256 GNDA.n4448 GNDA.n4308 0.0514167
R21257 GNDA.n4168 GNDA.n1600 0.0514167
R21258 GNDA.n4178 GNDA.n4177 0.0514167
R21259 GNDA.n4184 GNDA.n4183 0.0514167
R21260 GNDA.n4194 GNDA.n4193 0.0514167
R21261 GNDA.n4198 GNDA.n4197 0.0514167
R21262 GNDA.n4208 GNDA.n4207 0.0514167
R21263 GNDA.n4214 GNDA.n4213 0.0514167
R21264 GNDA.n4224 GNDA.n4223 0.0514167
R21265 GNDA.n4228 GNDA.n4227 0.0514167
R21266 GNDA.n4238 GNDA.n4237 0.0514167
R21267 GNDA.n4244 GNDA.n4243 0.0514167
R21268 GNDA.n4254 GNDA.n4253 0.0514167
R21269 GNDA.n4258 GNDA.n4257 0.0514167
R21270 GNDA.n4268 GNDA.n4267 0.0514167
R21271 GNDA.n4274 GNDA.n4273 0.0514167
R21272 GNDA.n4282 GNDA.n1624 0.0514167
R21273 GNDA.n1811 GNDA.n1810 0.0514167
R21274 GNDA.n1805 GNDA.n1804 0.0514167
R21275 GNDA.n1802 GNDA.n1801 0.0514167
R21276 GNDA.n1796 GNDA.n1795 0.0514167
R21277 GNDA.n1793 GNDA.n1792 0.0514167
R21278 GNDA.n1787 GNDA.n1786 0.0514167
R21279 GNDA.n1784 GNDA.n1783 0.0514167
R21280 GNDA.n1778 GNDA.n1777 0.0514167
R21281 GNDA.n1775 GNDA.n1774 0.0514167
R21282 GNDA.n1769 GNDA.n1768 0.0514167
R21283 GNDA.n1766 GNDA.n1765 0.0514167
R21284 GNDA.n1760 GNDA.n1759 0.0514167
R21285 GNDA.n1757 GNDA.n1756 0.0514167
R21286 GNDA.n1751 GNDA.n1750 0.0514167
R21287 GNDA.n1748 GNDA.n1747 0.0514167
R21288 GNDA.n1742 GNDA.n1741 0.0514167
R21289 GNDA.n3825 GNDA.n3775 0.0514167
R21290 GNDA.n3835 GNDA.n3834 0.0514167
R21291 GNDA.n3841 GNDA.n3840 0.0514167
R21292 GNDA.n3851 GNDA.n3850 0.0514167
R21293 GNDA.n3855 GNDA.n3854 0.0514167
R21294 GNDA.n3865 GNDA.n3864 0.0514167
R21295 GNDA.n3871 GNDA.n3870 0.0514167
R21296 GNDA.n3881 GNDA.n3880 0.0514167
R21297 GNDA.n3885 GNDA.n3884 0.0514167
R21298 GNDA.n3895 GNDA.n3894 0.0514167
R21299 GNDA.n3901 GNDA.n3900 0.0514167
R21300 GNDA.n3911 GNDA.n3910 0.0514167
R21301 GNDA.n3915 GNDA.n3914 0.0514167
R21302 GNDA.n3925 GNDA.n3924 0.0514167
R21303 GNDA.n3931 GNDA.n3930 0.0514167
R21304 GNDA.n3939 GNDA.n3799 0.0514167
R21305 GNDA.n4078 GNDA.n1837 0.0514167
R21306 GNDA.n3972 GNDA.n3971 0.0514167
R21307 GNDA.n3978 GNDA.n3977 0.0514167
R21308 GNDA.n3988 GNDA.n3987 0.0514167
R21309 GNDA.n3992 GNDA.n3991 0.0514167
R21310 GNDA.n4002 GNDA.n4001 0.0514167
R21311 GNDA.n4008 GNDA.n4007 0.0514167
R21312 GNDA.n4018 GNDA.n4017 0.0514167
R21313 GNDA.n4022 GNDA.n4021 0.0514167
R21314 GNDA.n4032 GNDA.n4031 0.0514167
R21315 GNDA.n4038 GNDA.n4037 0.0514167
R21316 GNDA.n4048 GNDA.n4047 0.0514167
R21317 GNDA.n4052 GNDA.n4051 0.0514167
R21318 GNDA.n4062 GNDA.n4061 0.0514167
R21319 GNDA.n4068 GNDA.n4067 0.0514167
R21320 GNDA.n4076 GNDA.n3941 0.0514167
R21321 GNDA.n3470 GNDA.n1839 0.0514167
R21322 GNDA.n3480 GNDA.n3479 0.0514167
R21323 GNDA.n3486 GNDA.n3485 0.0514167
R21324 GNDA.n3496 GNDA.n3495 0.0514167
R21325 GNDA.n3500 GNDA.n3499 0.0514167
R21326 GNDA.n3510 GNDA.n3509 0.0514167
R21327 GNDA.n3516 GNDA.n3515 0.0514167
R21328 GNDA.n3526 GNDA.n3525 0.0514167
R21329 GNDA.n3530 GNDA.n3529 0.0514167
R21330 GNDA.n3540 GNDA.n3539 0.0514167
R21331 GNDA.n3546 GNDA.n3545 0.0514167
R21332 GNDA.n3556 GNDA.n3555 0.0514167
R21333 GNDA.n3560 GNDA.n3559 0.0514167
R21334 GNDA.n3570 GNDA.n3569 0.0514167
R21335 GNDA.n3576 GNDA.n3575 0.0514167
R21336 GNDA.n3584 GNDA.n1863 0.0514167
R21337 GNDA.n2535 GNDA.n2486 0.0514167
R21338 GNDA.n2545 GNDA.n2544 0.0514167
R21339 GNDA.n2551 GNDA.n2550 0.0514167
R21340 GNDA.n2561 GNDA.n2560 0.0514167
R21341 GNDA.n2565 GNDA.n2564 0.0514167
R21342 GNDA.n2575 GNDA.n2574 0.0514167
R21343 GNDA.n2581 GNDA.n2580 0.0514167
R21344 GNDA.n2591 GNDA.n2590 0.0514167
R21345 GNDA.n2595 GNDA.n2594 0.0514167
R21346 GNDA.n2605 GNDA.n2604 0.0514167
R21347 GNDA.n2611 GNDA.n2610 0.0514167
R21348 GNDA.n2621 GNDA.n2620 0.0514167
R21349 GNDA.n2625 GNDA.n2624 0.0514167
R21350 GNDA.n2635 GNDA.n2634 0.0514167
R21351 GNDA.n2641 GNDA.n2640 0.0514167
R21352 GNDA.n2649 GNDA.n2510 0.0514167
R21353 GNDA.n2818 GNDA.n2438 0.0514167
R21354 GNDA.n2828 GNDA.n2827 0.0514167
R21355 GNDA.n2834 GNDA.n2833 0.0514167
R21356 GNDA.n2844 GNDA.n2843 0.0514167
R21357 GNDA.n2848 GNDA.n2847 0.0514167
R21358 GNDA.n2858 GNDA.n2857 0.0514167
R21359 GNDA.n2864 GNDA.n2863 0.0514167
R21360 GNDA.n2874 GNDA.n2873 0.0514167
R21361 GNDA.n2878 GNDA.n2877 0.0514167
R21362 GNDA.n2888 GNDA.n2887 0.0514167
R21363 GNDA.n2894 GNDA.n2893 0.0514167
R21364 GNDA.n2904 GNDA.n2903 0.0514167
R21365 GNDA.n2908 GNDA.n2907 0.0514167
R21366 GNDA.n2918 GNDA.n2917 0.0514167
R21367 GNDA.n2924 GNDA.n2923 0.0514167
R21368 GNDA.n2932 GNDA.n2793 0.0514167
R21369 GNDA.n2959 GNDA.n2414 0.0514167
R21370 GNDA.n2969 GNDA.n2968 0.0514167
R21371 GNDA.n2975 GNDA.n2974 0.0514167
R21372 GNDA.n2985 GNDA.n2984 0.0514167
R21373 GNDA.n2989 GNDA.n2988 0.0514167
R21374 GNDA.n2999 GNDA.n2998 0.0514167
R21375 GNDA.n3005 GNDA.n3004 0.0514167
R21376 GNDA.n3015 GNDA.n3014 0.0514167
R21377 GNDA.n3019 GNDA.n3018 0.0514167
R21378 GNDA.n3029 GNDA.n3028 0.0514167
R21379 GNDA.n3035 GNDA.n3034 0.0514167
R21380 GNDA.n3045 GNDA.n3044 0.0514167
R21381 GNDA.n3049 GNDA.n3048 0.0514167
R21382 GNDA.n3059 GNDA.n3058 0.0514167
R21383 GNDA.n3065 GNDA.n3064 0.0514167
R21384 GNDA.n3073 GNDA.n2934 0.0514167
R21385 GNDA.n3100 GNDA.n2390 0.0514167
R21386 GNDA.n3110 GNDA.n3109 0.0514167
R21387 GNDA.n3116 GNDA.n3115 0.0514167
R21388 GNDA.n3126 GNDA.n3125 0.0514167
R21389 GNDA.n3130 GNDA.n3129 0.0514167
R21390 GNDA.n3140 GNDA.n3139 0.0514167
R21391 GNDA.n3146 GNDA.n3145 0.0514167
R21392 GNDA.n3156 GNDA.n3155 0.0514167
R21393 GNDA.n3160 GNDA.n3159 0.0514167
R21394 GNDA.n3170 GNDA.n3169 0.0514167
R21395 GNDA.n3176 GNDA.n3175 0.0514167
R21396 GNDA.n3186 GNDA.n3185 0.0514167
R21397 GNDA.n3190 GNDA.n3189 0.0514167
R21398 GNDA.n3200 GNDA.n3199 0.0514167
R21399 GNDA.n3206 GNDA.n3205 0.0514167
R21400 GNDA.n3214 GNDA.n3075 0.0514167
R21401 GNDA.n6354 GNDA.n6287 0.0514167
R21402 GNDA.n6351 GNDA.n6350 0.0514167
R21403 GNDA.n6366 GNDA.n6365 0.0514167
R21404 GNDA.n6374 GNDA.n6373 0.0514167
R21405 GNDA.n6343 GNDA.n6342 0.0514167
R21406 GNDA.n6339 GNDA.n6338 0.0514167
R21407 GNDA.n6390 GNDA.n6389 0.0514167
R21408 GNDA.n6398 GNDA.n6397 0.0514167
R21409 GNDA.n6331 GNDA.n6330 0.0514167
R21410 GNDA.n6327 GNDA.n6326 0.0514167
R21411 GNDA.n6414 GNDA.n6413 0.0514167
R21412 GNDA.n6422 GNDA.n6421 0.0514167
R21413 GNDA.n6319 GNDA.n6318 0.0514167
R21414 GNDA.n6315 GNDA.n6314 0.0514167
R21415 GNDA.n6438 GNDA.n6437 0.0514167
R21416 GNDA.n6616 GNDA.n360 0.0514167
R21417 GNDA.n410 GNDA.n362 0.0514167
R21418 GNDA.n420 GNDA.n419 0.0514167
R21419 GNDA.n426 GNDA.n425 0.0514167
R21420 GNDA.n436 GNDA.n435 0.0514167
R21421 GNDA.n440 GNDA.n439 0.0514167
R21422 GNDA.n450 GNDA.n449 0.0514167
R21423 GNDA.n456 GNDA.n455 0.0514167
R21424 GNDA.n466 GNDA.n465 0.0514167
R21425 GNDA.n470 GNDA.n469 0.0514167
R21426 GNDA.n480 GNDA.n479 0.0514167
R21427 GNDA.n486 GNDA.n485 0.0514167
R21428 GNDA.n496 GNDA.n495 0.0514167
R21429 GNDA.n500 GNDA.n499 0.0514167
R21430 GNDA.n510 GNDA.n509 0.0514167
R21431 GNDA.n516 GNDA.n515 0.0514167
R21432 GNDA.n6285 GNDA.n386 0.0514167
R21433 GNDA.n1900 GNDA.n1899 0.0475
R21434 GNDA.n2363 GNDA.n1908 0.0475
R21435 GNDA.n1915 GNDA.n1914 0.0475
R21436 GNDA.n2372 GNDA.n1923 0.0475
R21437 GNDA.n1930 GNDA.n1929 0.0475
R21438 GNDA.n2381 GNDA.n1938 0.0475
R21439 GNDA.n1945 GNDA.n1944 0.0475
R21440 GNDA.n2247 GNDA 0.0414781
R21441 GNDA.n4665 GNDA.n4450 0.028198
R21442 GNDA.n4669 GNDA.n4451 0.028198
R21443 GNDA.n4679 GNDA.n4453 0.028198
R21444 GNDA.n4685 GNDA.n4454 0.028198
R21445 GNDA.n4695 GNDA.n4456 0.028198
R21446 GNDA.n4699 GNDA.n4457 0.028198
R21447 GNDA.n4709 GNDA.n4459 0.028198
R21448 GNDA.n4715 GNDA.n4460 0.028198
R21449 GNDA.n4725 GNDA.n4462 0.028198
R21450 GNDA.n4729 GNDA.n4463 0.028198
R21451 GNDA.n4739 GNDA.n4465 0.028198
R21452 GNDA.n4745 GNDA.n4466 0.028198
R21453 GNDA.n4755 GNDA.n4468 0.028198
R21454 GNDA.n4759 GNDA.n4469 0.028198
R21455 GNDA.n4769 GNDA.n4471 0.028198
R21456 GNDA.n4639 GNDA.n4472 0.028198
R21457 GNDA.n5692 GNDA.n4973 0.028198
R21458 GNDA.n5696 GNDA.n4974 0.028198
R21459 GNDA.n5706 GNDA.n4976 0.028198
R21460 GNDA.n5712 GNDA.n4977 0.028198
R21461 GNDA.n5722 GNDA.n4979 0.028198
R21462 GNDA.n5726 GNDA.n4980 0.028198
R21463 GNDA.n5736 GNDA.n4982 0.028198
R21464 GNDA.n5742 GNDA.n4983 0.028198
R21465 GNDA.n5752 GNDA.n4985 0.028198
R21466 GNDA.n5756 GNDA.n4986 0.028198
R21467 GNDA.n5766 GNDA.n4988 0.028198
R21468 GNDA.n5772 GNDA.n4989 0.028198
R21469 GNDA.n5782 GNDA.n4991 0.028198
R21470 GNDA.n5786 GNDA.n4992 0.028198
R21471 GNDA.n5796 GNDA.n4994 0.028198
R21472 GNDA.n5662 GNDA.n4995 0.028198
R21473 GNDA.n2695 GNDA.n2463 0.028198
R21474 GNDA.n2706 GNDA.n2464 0.028198
R21475 GNDA.n2714 GNDA.n2466 0.028198
R21476 GNDA.n2687 GNDA.n2467 0.028198
R21477 GNDA.n2683 GNDA.n2469 0.028198
R21478 GNDA.n2730 GNDA.n2470 0.028198
R21479 GNDA.n2738 GNDA.n2472 0.028198
R21480 GNDA.n2675 GNDA.n2473 0.028198
R21481 GNDA.n2671 GNDA.n2475 0.028198
R21482 GNDA.n2754 GNDA.n2476 0.028198
R21483 GNDA.n2762 GNDA.n2478 0.028198
R21484 GNDA.n2663 GNDA.n2479 0.028198
R21485 GNDA.n2659 GNDA.n2481 0.028198
R21486 GNDA.n2778 GNDA.n2482 0.028198
R21487 GNDA.n2786 GNDA.n2484 0.028198
R21488 GNDA.n2651 GNDA.n2485 0.028198
R21489 GNDA.n5970 GNDA.n4925 0.028198
R21490 GNDA.n5974 GNDA.n4926 0.028198
R21491 GNDA.n5984 GNDA.n4928 0.028198
R21492 GNDA.n5990 GNDA.n4929 0.028198
R21493 GNDA.n6000 GNDA.n4931 0.028198
R21494 GNDA.n6004 GNDA.n4932 0.028198
R21495 GNDA.n6014 GNDA.n4934 0.028198
R21496 GNDA.n6020 GNDA.n4935 0.028198
R21497 GNDA.n6030 GNDA.n4937 0.028198
R21498 GNDA.n6034 GNDA.n4938 0.028198
R21499 GNDA.n6044 GNDA.n4940 0.028198
R21500 GNDA.n6050 GNDA.n4941 0.028198
R21501 GNDA.n6060 GNDA.n4943 0.028198
R21502 GNDA.n6064 GNDA.n4944 0.028198
R21503 GNDA.n6074 GNDA.n4946 0.028198
R21504 GNDA.n5944 GNDA.n4947 0.028198
R21505 GNDA.n1583 GNDA.n1582 0.028198
R21506 GNDA.n1580 GNDA.n1579 0.028198
R21507 GNDA.n1574 GNDA.n1573 0.028198
R21508 GNDA.n1571 GNDA.n1570 0.028198
R21509 GNDA.n1565 GNDA.n1564 0.028198
R21510 GNDA.n1562 GNDA.n1561 0.028198
R21511 GNDA.n1556 GNDA.n1555 0.028198
R21512 GNDA.n1553 GNDA.n1552 0.028198
R21513 GNDA.n1547 GNDA.n1546 0.028198
R21514 GNDA.n1544 GNDA.n1543 0.028198
R21515 GNDA.n1538 GNDA.n1537 0.028198
R21516 GNDA.n1535 GNDA.n1534 0.028198
R21517 GNDA.n1529 GNDA.n1528 0.028198
R21518 GNDA.n1526 GNDA.n1525 0.028198
R21519 GNDA.n1520 GNDA.n1519 0.028198
R21520 GNDA.n1517 GNDA.n1516 0.028198
R21521 GNDA.n3641 GNDA.n3587 0.028198
R21522 GNDA.n3645 GNDA.n3588 0.028198
R21523 GNDA.n3655 GNDA.n3590 0.028198
R21524 GNDA.n3661 GNDA.n3591 0.028198
R21525 GNDA.n3671 GNDA.n3593 0.028198
R21526 GNDA.n3675 GNDA.n3594 0.028198
R21527 GNDA.n3685 GNDA.n3596 0.028198
R21528 GNDA.n3691 GNDA.n3597 0.028198
R21529 GNDA.n3701 GNDA.n3599 0.028198
R21530 GNDA.n3705 GNDA.n3600 0.028198
R21531 GNDA.n3715 GNDA.n3602 0.028198
R21532 GNDA.n3721 GNDA.n3603 0.028198
R21533 GNDA.n3731 GNDA.n3605 0.028198
R21534 GNDA.n3735 GNDA.n3606 0.028198
R21535 GNDA.n3745 GNDA.n3608 0.028198
R21536 GNDA.n3610 GNDA.n3609 0.028198
R21537 GNDA.n3455 GNDA.n3454 0.028198
R21538 GNDA.n3452 GNDA.n3451 0.028198
R21539 GNDA.n3446 GNDA.n3445 0.028198
R21540 GNDA.n3443 GNDA.n3442 0.028198
R21541 GNDA.n3437 GNDA.n3436 0.028198
R21542 GNDA.n3434 GNDA.n3433 0.028198
R21543 GNDA.n3428 GNDA.n3427 0.028198
R21544 GNDA.n3425 GNDA.n3424 0.028198
R21545 GNDA.n3419 GNDA.n3418 0.028198
R21546 GNDA.n3416 GNDA.n3415 0.028198
R21547 GNDA.n3410 GNDA.n3409 0.028198
R21548 GNDA.n3407 GNDA.n3406 0.028198
R21549 GNDA.n3401 GNDA.n3400 0.028198
R21550 GNDA.n3398 GNDA.n3397 0.028198
R21551 GNDA.n3392 GNDA.n3391 0.028198
R21552 GNDA.n3389 GNDA.n3388 0.028198
R21553 GNDA.n5121 GNDA.n5072 0.028198
R21554 GNDA.n5125 GNDA.n5073 0.028198
R21555 GNDA.n5135 GNDA.n5075 0.028198
R21556 GNDA.n5141 GNDA.n5076 0.028198
R21557 GNDA.n5151 GNDA.n5078 0.028198
R21558 GNDA.n5155 GNDA.n5079 0.028198
R21559 GNDA.n5165 GNDA.n5081 0.028198
R21560 GNDA.n5171 GNDA.n5082 0.028198
R21561 GNDA.n5181 GNDA.n5084 0.028198
R21562 GNDA.n5185 GNDA.n5085 0.028198
R21563 GNDA.n5195 GNDA.n5087 0.028198
R21564 GNDA.n5201 GNDA.n5088 0.028198
R21565 GNDA.n5211 GNDA.n5090 0.028198
R21566 GNDA.n5215 GNDA.n5091 0.028198
R21567 GNDA.n5225 GNDA.n5093 0.028198
R21568 GNDA.n5095 GNDA.n5094 0.028198
R21569 GNDA.n5395 GNDA.n5394 0.028198
R21570 GNDA.n5392 GNDA.n5391 0.028198
R21571 GNDA.n5386 GNDA.n5385 0.028198
R21572 GNDA.n5383 GNDA.n5382 0.028198
R21573 GNDA.n5377 GNDA.n5376 0.028198
R21574 GNDA.n5374 GNDA.n5373 0.028198
R21575 GNDA.n5368 GNDA.n5367 0.028198
R21576 GNDA.n5365 GNDA.n5364 0.028198
R21577 GNDA.n5359 GNDA.n5358 0.028198
R21578 GNDA.n5356 GNDA.n5355 0.028198
R21579 GNDA.n5350 GNDA.n5349 0.028198
R21580 GNDA.n5347 GNDA.n5346 0.028198
R21581 GNDA.n5341 GNDA.n5340 0.028198
R21582 GNDA.n5338 GNDA.n5337 0.028198
R21583 GNDA.n5332 GNDA.n5331 0.028198
R21584 GNDA.n5329 GNDA.n5328 0.028198
R21585 GNDA.n5409 GNDA.n5021 0.028198
R21586 GNDA.n5413 GNDA.n5022 0.028198
R21587 GNDA.n5423 GNDA.n5024 0.028198
R21588 GNDA.n5429 GNDA.n5025 0.028198
R21589 GNDA.n5439 GNDA.n5027 0.028198
R21590 GNDA.n5443 GNDA.n5028 0.028198
R21591 GNDA.n5453 GNDA.n5030 0.028198
R21592 GNDA.n5459 GNDA.n5031 0.028198
R21593 GNDA.n5469 GNDA.n5033 0.028198
R21594 GNDA.n5473 GNDA.n5034 0.028198
R21595 GNDA.n5483 GNDA.n5036 0.028198
R21596 GNDA.n5489 GNDA.n5037 0.028198
R21597 GNDA.n5499 GNDA.n5039 0.028198
R21598 GNDA.n5503 GNDA.n5040 0.028198
R21599 GNDA.n5513 GNDA.n5042 0.028198
R21600 GNDA.n5045 GNDA.n5043 0.028198
R21601 GNDA.n5551 GNDA.n4997 0.028198
R21602 GNDA.n5555 GNDA.n4998 0.028198
R21603 GNDA.n5565 GNDA.n5000 0.028198
R21604 GNDA.n5571 GNDA.n5001 0.028198
R21605 GNDA.n5581 GNDA.n5003 0.028198
R21606 GNDA.n5585 GNDA.n5004 0.028198
R21607 GNDA.n5595 GNDA.n5006 0.028198
R21608 GNDA.n5601 GNDA.n5007 0.028198
R21609 GNDA.n5611 GNDA.n5009 0.028198
R21610 GNDA.n5615 GNDA.n5010 0.028198
R21611 GNDA.n5625 GNDA.n5012 0.028198
R21612 GNDA.n5631 GNDA.n5013 0.028198
R21613 GNDA.n5641 GNDA.n5015 0.028198
R21614 GNDA.n5645 GNDA.n5016 0.028198
R21615 GNDA.n5655 GNDA.n5018 0.028198
R21616 GNDA.n5520 GNDA.n5019 0.028198
R21617 GNDA.n5833 GNDA.n4949 0.028198
R21618 GNDA.n5837 GNDA.n4950 0.028198
R21619 GNDA.n5847 GNDA.n4952 0.028198
R21620 GNDA.n5853 GNDA.n4953 0.028198
R21621 GNDA.n5863 GNDA.n4955 0.028198
R21622 GNDA.n5867 GNDA.n4956 0.028198
R21623 GNDA.n5877 GNDA.n4958 0.028198
R21624 GNDA.n5883 GNDA.n4959 0.028198
R21625 GNDA.n5893 GNDA.n4961 0.028198
R21626 GNDA.n5897 GNDA.n4962 0.028198
R21627 GNDA.n5907 GNDA.n4964 0.028198
R21628 GNDA.n5913 GNDA.n4965 0.028198
R21629 GNDA.n5923 GNDA.n4967 0.028198
R21630 GNDA.n5927 GNDA.n4968 0.028198
R21631 GNDA.n5937 GNDA.n4970 0.028198
R21632 GNDA.n5803 GNDA.n4971 0.028198
R21633 GNDA.n4814 GNDA.n1373 0.028198
R21634 GNDA.n4818 GNDA.n1374 0.028198
R21635 GNDA.n4828 GNDA.n1376 0.028198
R21636 GNDA.n4834 GNDA.n1377 0.028198
R21637 GNDA.n4844 GNDA.n1379 0.028198
R21638 GNDA.n4848 GNDA.n1380 0.028198
R21639 GNDA.n4858 GNDA.n1382 0.028198
R21640 GNDA.n4864 GNDA.n1383 0.028198
R21641 GNDA.n4874 GNDA.n1385 0.028198
R21642 GNDA.n4878 GNDA.n1386 0.028198
R21643 GNDA.n4888 GNDA.n1388 0.028198
R21644 GNDA.n4894 GNDA.n1389 0.028198
R21645 GNDA.n4904 GNDA.n1391 0.028198
R21646 GNDA.n4908 GNDA.n1392 0.028198
R21647 GNDA.n4918 GNDA.n1394 0.028198
R21648 GNDA.n1396 GNDA.n1395 0.028198
R21649 GNDA.n4528 GNDA.n4474 0.028198
R21650 GNDA.n4532 GNDA.n4475 0.028198
R21651 GNDA.n4542 GNDA.n4477 0.028198
R21652 GNDA.n4548 GNDA.n4478 0.028198
R21653 GNDA.n4558 GNDA.n4480 0.028198
R21654 GNDA.n4562 GNDA.n4481 0.028198
R21655 GNDA.n4572 GNDA.n4483 0.028198
R21656 GNDA.n4578 GNDA.n4484 0.028198
R21657 GNDA.n4588 GNDA.n4486 0.028198
R21658 GNDA.n4592 GNDA.n4487 0.028198
R21659 GNDA.n4602 GNDA.n4489 0.028198
R21660 GNDA.n4608 GNDA.n4490 0.028198
R21661 GNDA.n4618 GNDA.n4492 0.028198
R21662 GNDA.n4622 GNDA.n4493 0.028198
R21663 GNDA.n4632 GNDA.n4495 0.028198
R21664 GNDA.n4497 GNDA.n4496 0.028198
R21665 GNDA.n4339 GNDA.n4285 0.028198
R21666 GNDA.n4343 GNDA.n4286 0.028198
R21667 GNDA.n4353 GNDA.n4288 0.028198
R21668 GNDA.n4359 GNDA.n4289 0.028198
R21669 GNDA.n4369 GNDA.n4291 0.028198
R21670 GNDA.n4373 GNDA.n4292 0.028198
R21671 GNDA.n4383 GNDA.n4294 0.028198
R21672 GNDA.n4389 GNDA.n4295 0.028198
R21673 GNDA.n4399 GNDA.n4297 0.028198
R21674 GNDA.n4403 GNDA.n4298 0.028198
R21675 GNDA.n4413 GNDA.n4300 0.028198
R21676 GNDA.n4419 GNDA.n4301 0.028198
R21677 GNDA.n4429 GNDA.n4303 0.028198
R21678 GNDA.n4433 GNDA.n4304 0.028198
R21679 GNDA.n4443 GNDA.n4306 0.028198
R21680 GNDA.n4308 GNDA.n4307 0.028198
R21681 GNDA.n4173 GNDA.n1601 0.028198
R21682 GNDA.n4177 GNDA.n1602 0.028198
R21683 GNDA.n4187 GNDA.n1604 0.028198
R21684 GNDA.n4193 GNDA.n1605 0.028198
R21685 GNDA.n4203 GNDA.n1607 0.028198
R21686 GNDA.n4207 GNDA.n1608 0.028198
R21687 GNDA.n4217 GNDA.n1610 0.028198
R21688 GNDA.n4223 GNDA.n1611 0.028198
R21689 GNDA.n4233 GNDA.n1613 0.028198
R21690 GNDA.n4237 GNDA.n1614 0.028198
R21691 GNDA.n4247 GNDA.n1616 0.028198
R21692 GNDA.n4253 GNDA.n1617 0.028198
R21693 GNDA.n4263 GNDA.n1619 0.028198
R21694 GNDA.n4267 GNDA.n1620 0.028198
R21695 GNDA.n4277 GNDA.n1622 0.028198
R21696 GNDA.n1624 GNDA.n1623 0.028198
R21697 GNDA.n1809 GNDA.n1808 0.028198
R21698 GNDA.n1806 GNDA.n1805 0.028198
R21699 GNDA.n1800 GNDA.n1799 0.028198
R21700 GNDA.n1797 GNDA.n1796 0.028198
R21701 GNDA.n1791 GNDA.n1790 0.028198
R21702 GNDA.n1788 GNDA.n1787 0.028198
R21703 GNDA.n1782 GNDA.n1781 0.028198
R21704 GNDA.n1779 GNDA.n1778 0.028198
R21705 GNDA.n1773 GNDA.n1772 0.028198
R21706 GNDA.n1770 GNDA.n1769 0.028198
R21707 GNDA.n1764 GNDA.n1763 0.028198
R21708 GNDA.n1761 GNDA.n1760 0.028198
R21709 GNDA.n1755 GNDA.n1754 0.028198
R21710 GNDA.n1752 GNDA.n1751 0.028198
R21711 GNDA.n1746 GNDA.n1745 0.028198
R21712 GNDA.n1743 GNDA.n1742 0.028198
R21713 GNDA.n3830 GNDA.n3776 0.028198
R21714 GNDA.n3834 GNDA.n3777 0.028198
R21715 GNDA.n3844 GNDA.n3779 0.028198
R21716 GNDA.n3850 GNDA.n3780 0.028198
R21717 GNDA.n3860 GNDA.n3782 0.028198
R21718 GNDA.n3864 GNDA.n3783 0.028198
R21719 GNDA.n3874 GNDA.n3785 0.028198
R21720 GNDA.n3880 GNDA.n3786 0.028198
R21721 GNDA.n3890 GNDA.n3788 0.028198
R21722 GNDA.n3894 GNDA.n3789 0.028198
R21723 GNDA.n3904 GNDA.n3791 0.028198
R21724 GNDA.n3910 GNDA.n3792 0.028198
R21725 GNDA.n3920 GNDA.n3794 0.028198
R21726 GNDA.n3924 GNDA.n3795 0.028198
R21727 GNDA.n3934 GNDA.n3797 0.028198
R21728 GNDA.n3799 GNDA.n3798 0.028198
R21729 GNDA.n3967 GNDA.n3752 0.028198
R21730 GNDA.n3971 GNDA.n3753 0.028198
R21731 GNDA.n3981 GNDA.n3755 0.028198
R21732 GNDA.n3987 GNDA.n3756 0.028198
R21733 GNDA.n3997 GNDA.n3758 0.028198
R21734 GNDA.n4001 GNDA.n3759 0.028198
R21735 GNDA.n4011 GNDA.n3761 0.028198
R21736 GNDA.n4017 GNDA.n3762 0.028198
R21737 GNDA.n4027 GNDA.n3764 0.028198
R21738 GNDA.n4031 GNDA.n3765 0.028198
R21739 GNDA.n4041 GNDA.n3767 0.028198
R21740 GNDA.n4047 GNDA.n3768 0.028198
R21741 GNDA.n4057 GNDA.n3770 0.028198
R21742 GNDA.n4061 GNDA.n3771 0.028198
R21743 GNDA.n4071 GNDA.n3773 0.028198
R21744 GNDA.n3941 GNDA.n3774 0.028198
R21745 GNDA.n3475 GNDA.n1840 0.028198
R21746 GNDA.n3479 GNDA.n1841 0.028198
R21747 GNDA.n3489 GNDA.n1843 0.028198
R21748 GNDA.n3495 GNDA.n1844 0.028198
R21749 GNDA.n3505 GNDA.n1846 0.028198
R21750 GNDA.n3509 GNDA.n1847 0.028198
R21751 GNDA.n3519 GNDA.n1849 0.028198
R21752 GNDA.n3525 GNDA.n1850 0.028198
R21753 GNDA.n3535 GNDA.n1852 0.028198
R21754 GNDA.n3539 GNDA.n1853 0.028198
R21755 GNDA.n3549 GNDA.n1855 0.028198
R21756 GNDA.n3555 GNDA.n1856 0.028198
R21757 GNDA.n3565 GNDA.n1858 0.028198
R21758 GNDA.n3569 GNDA.n1859 0.028198
R21759 GNDA.n3579 GNDA.n1861 0.028198
R21760 GNDA.n1863 GNDA.n1862 0.028198
R21761 GNDA.n2540 GNDA.n2487 0.028198
R21762 GNDA.n2544 GNDA.n2488 0.028198
R21763 GNDA.n2554 GNDA.n2490 0.028198
R21764 GNDA.n2560 GNDA.n2491 0.028198
R21765 GNDA.n2570 GNDA.n2493 0.028198
R21766 GNDA.n2574 GNDA.n2494 0.028198
R21767 GNDA.n2584 GNDA.n2496 0.028198
R21768 GNDA.n2590 GNDA.n2497 0.028198
R21769 GNDA.n2600 GNDA.n2499 0.028198
R21770 GNDA.n2604 GNDA.n2500 0.028198
R21771 GNDA.n2614 GNDA.n2502 0.028198
R21772 GNDA.n2620 GNDA.n2503 0.028198
R21773 GNDA.n2630 GNDA.n2505 0.028198
R21774 GNDA.n2634 GNDA.n2506 0.028198
R21775 GNDA.n2644 GNDA.n2508 0.028198
R21776 GNDA.n2510 GNDA.n2509 0.028198
R21777 GNDA.n2823 GNDA.n2439 0.028198
R21778 GNDA.n2827 GNDA.n2440 0.028198
R21779 GNDA.n2837 GNDA.n2442 0.028198
R21780 GNDA.n2843 GNDA.n2443 0.028198
R21781 GNDA.n2853 GNDA.n2445 0.028198
R21782 GNDA.n2857 GNDA.n2446 0.028198
R21783 GNDA.n2867 GNDA.n2448 0.028198
R21784 GNDA.n2873 GNDA.n2449 0.028198
R21785 GNDA.n2883 GNDA.n2451 0.028198
R21786 GNDA.n2887 GNDA.n2452 0.028198
R21787 GNDA.n2897 GNDA.n2454 0.028198
R21788 GNDA.n2903 GNDA.n2455 0.028198
R21789 GNDA.n2913 GNDA.n2457 0.028198
R21790 GNDA.n2917 GNDA.n2458 0.028198
R21791 GNDA.n2927 GNDA.n2460 0.028198
R21792 GNDA.n2793 GNDA.n2461 0.028198
R21793 GNDA.n2964 GNDA.n2415 0.028198
R21794 GNDA.n2968 GNDA.n2416 0.028198
R21795 GNDA.n2978 GNDA.n2418 0.028198
R21796 GNDA.n2984 GNDA.n2419 0.028198
R21797 GNDA.n2994 GNDA.n2421 0.028198
R21798 GNDA.n2998 GNDA.n2422 0.028198
R21799 GNDA.n3008 GNDA.n2424 0.028198
R21800 GNDA.n3014 GNDA.n2425 0.028198
R21801 GNDA.n3024 GNDA.n2427 0.028198
R21802 GNDA.n3028 GNDA.n2428 0.028198
R21803 GNDA.n3038 GNDA.n2430 0.028198
R21804 GNDA.n3044 GNDA.n2431 0.028198
R21805 GNDA.n3054 GNDA.n2433 0.028198
R21806 GNDA.n3058 GNDA.n2434 0.028198
R21807 GNDA.n3068 GNDA.n2436 0.028198
R21808 GNDA.n2934 GNDA.n2437 0.028198
R21809 GNDA.n3105 GNDA.n2391 0.028198
R21810 GNDA.n3109 GNDA.n2392 0.028198
R21811 GNDA.n3119 GNDA.n2394 0.028198
R21812 GNDA.n3125 GNDA.n2395 0.028198
R21813 GNDA.n3135 GNDA.n2397 0.028198
R21814 GNDA.n3139 GNDA.n2398 0.028198
R21815 GNDA.n3149 GNDA.n2400 0.028198
R21816 GNDA.n3155 GNDA.n2401 0.028198
R21817 GNDA.n3165 GNDA.n2403 0.028198
R21818 GNDA.n3169 GNDA.n2404 0.028198
R21819 GNDA.n3179 GNDA.n2406 0.028198
R21820 GNDA.n3185 GNDA.n2407 0.028198
R21821 GNDA.n3195 GNDA.n2409 0.028198
R21822 GNDA.n3199 GNDA.n2410 0.028198
R21823 GNDA.n3209 GNDA.n2412 0.028198
R21824 GNDA.n3075 GNDA.n2413 0.028198
R21825 GNDA.n3210 GNDA.n2413 0.028198
R21826 GNDA.n3206 GNDA.n2412 0.028198
R21827 GNDA.n3196 GNDA.n2410 0.028198
R21828 GNDA.n3190 GNDA.n2409 0.028198
R21829 GNDA.n3180 GNDA.n2407 0.028198
R21830 GNDA.n3176 GNDA.n2406 0.028198
R21831 GNDA.n3166 GNDA.n2404 0.028198
R21832 GNDA.n3160 GNDA.n2403 0.028198
R21833 GNDA.n3150 GNDA.n2401 0.028198
R21834 GNDA.n3146 GNDA.n2400 0.028198
R21835 GNDA.n3136 GNDA.n2398 0.028198
R21836 GNDA.n3130 GNDA.n2397 0.028198
R21837 GNDA.n3120 GNDA.n2395 0.028198
R21838 GNDA.n3116 GNDA.n2394 0.028198
R21839 GNDA.n3106 GNDA.n2392 0.028198
R21840 GNDA.n3100 GNDA.n2391 0.028198
R21841 GNDA.n3069 GNDA.n2437 0.028198
R21842 GNDA.n3065 GNDA.n2436 0.028198
R21843 GNDA.n3055 GNDA.n2434 0.028198
R21844 GNDA.n3049 GNDA.n2433 0.028198
R21845 GNDA.n3039 GNDA.n2431 0.028198
R21846 GNDA.n3035 GNDA.n2430 0.028198
R21847 GNDA.n3025 GNDA.n2428 0.028198
R21848 GNDA.n3019 GNDA.n2427 0.028198
R21849 GNDA.n3009 GNDA.n2425 0.028198
R21850 GNDA.n3005 GNDA.n2424 0.028198
R21851 GNDA.n2995 GNDA.n2422 0.028198
R21852 GNDA.n2989 GNDA.n2421 0.028198
R21853 GNDA.n2979 GNDA.n2419 0.028198
R21854 GNDA.n2975 GNDA.n2418 0.028198
R21855 GNDA.n2965 GNDA.n2416 0.028198
R21856 GNDA.n2959 GNDA.n2415 0.028198
R21857 GNDA.n2928 GNDA.n2461 0.028198
R21858 GNDA.n2924 GNDA.n2460 0.028198
R21859 GNDA.n2914 GNDA.n2458 0.028198
R21860 GNDA.n2908 GNDA.n2457 0.028198
R21861 GNDA.n2898 GNDA.n2455 0.028198
R21862 GNDA.n2894 GNDA.n2454 0.028198
R21863 GNDA.n2884 GNDA.n2452 0.028198
R21864 GNDA.n2878 GNDA.n2451 0.028198
R21865 GNDA.n2868 GNDA.n2449 0.028198
R21866 GNDA.n2864 GNDA.n2448 0.028198
R21867 GNDA.n2854 GNDA.n2446 0.028198
R21868 GNDA.n2848 GNDA.n2445 0.028198
R21869 GNDA.n2838 GNDA.n2443 0.028198
R21870 GNDA.n2834 GNDA.n2442 0.028198
R21871 GNDA.n2824 GNDA.n2440 0.028198
R21872 GNDA.n2818 GNDA.n2439 0.028198
R21873 GNDA.n2645 GNDA.n2509 0.028198
R21874 GNDA.n2641 GNDA.n2508 0.028198
R21875 GNDA.n2631 GNDA.n2506 0.028198
R21876 GNDA.n2625 GNDA.n2505 0.028198
R21877 GNDA.n2615 GNDA.n2503 0.028198
R21878 GNDA.n2611 GNDA.n2502 0.028198
R21879 GNDA.n2601 GNDA.n2500 0.028198
R21880 GNDA.n2595 GNDA.n2499 0.028198
R21881 GNDA.n2585 GNDA.n2497 0.028198
R21882 GNDA.n2581 GNDA.n2496 0.028198
R21883 GNDA.n2571 GNDA.n2494 0.028198
R21884 GNDA.n2565 GNDA.n2493 0.028198
R21885 GNDA.n2555 GNDA.n2491 0.028198
R21886 GNDA.n2551 GNDA.n2490 0.028198
R21887 GNDA.n2541 GNDA.n2488 0.028198
R21888 GNDA.n2535 GNDA.n2487 0.028198
R21889 GNDA.n3580 GNDA.n1862 0.028198
R21890 GNDA.n3576 GNDA.n1861 0.028198
R21891 GNDA.n3566 GNDA.n1859 0.028198
R21892 GNDA.n3560 GNDA.n1858 0.028198
R21893 GNDA.n3550 GNDA.n1856 0.028198
R21894 GNDA.n3546 GNDA.n1855 0.028198
R21895 GNDA.n3536 GNDA.n1853 0.028198
R21896 GNDA.n3530 GNDA.n1852 0.028198
R21897 GNDA.n3520 GNDA.n1850 0.028198
R21898 GNDA.n3516 GNDA.n1849 0.028198
R21899 GNDA.n3506 GNDA.n1847 0.028198
R21900 GNDA.n3500 GNDA.n1846 0.028198
R21901 GNDA.n3490 GNDA.n1844 0.028198
R21902 GNDA.n3486 GNDA.n1843 0.028198
R21903 GNDA.n3476 GNDA.n1841 0.028198
R21904 GNDA.n3470 GNDA.n1840 0.028198
R21905 GNDA.n4072 GNDA.n3774 0.028198
R21906 GNDA.n4068 GNDA.n3773 0.028198
R21907 GNDA.n4058 GNDA.n3771 0.028198
R21908 GNDA.n4052 GNDA.n3770 0.028198
R21909 GNDA.n4042 GNDA.n3768 0.028198
R21910 GNDA.n4038 GNDA.n3767 0.028198
R21911 GNDA.n4028 GNDA.n3765 0.028198
R21912 GNDA.n4022 GNDA.n3764 0.028198
R21913 GNDA.n4012 GNDA.n3762 0.028198
R21914 GNDA.n4008 GNDA.n3761 0.028198
R21915 GNDA.n3998 GNDA.n3759 0.028198
R21916 GNDA.n3992 GNDA.n3758 0.028198
R21917 GNDA.n3982 GNDA.n3756 0.028198
R21918 GNDA.n3978 GNDA.n3755 0.028198
R21919 GNDA.n3968 GNDA.n3753 0.028198
R21920 GNDA.n3752 GNDA.n1837 0.028198
R21921 GNDA.n3935 GNDA.n3798 0.028198
R21922 GNDA.n3931 GNDA.n3797 0.028198
R21923 GNDA.n3921 GNDA.n3795 0.028198
R21924 GNDA.n3915 GNDA.n3794 0.028198
R21925 GNDA.n3905 GNDA.n3792 0.028198
R21926 GNDA.n3901 GNDA.n3791 0.028198
R21927 GNDA.n3891 GNDA.n3789 0.028198
R21928 GNDA.n3885 GNDA.n3788 0.028198
R21929 GNDA.n3875 GNDA.n3786 0.028198
R21930 GNDA.n3871 GNDA.n3785 0.028198
R21931 GNDA.n3861 GNDA.n3783 0.028198
R21932 GNDA.n3855 GNDA.n3782 0.028198
R21933 GNDA.n3845 GNDA.n3780 0.028198
R21934 GNDA.n3841 GNDA.n3779 0.028198
R21935 GNDA.n3831 GNDA.n3777 0.028198
R21936 GNDA.n3825 GNDA.n3776 0.028198
R21937 GNDA.n1744 GNDA.n1743 0.028198
R21938 GNDA.n1747 GNDA.n1746 0.028198
R21939 GNDA.n1753 GNDA.n1752 0.028198
R21940 GNDA.n1756 GNDA.n1755 0.028198
R21941 GNDA.n1762 GNDA.n1761 0.028198
R21942 GNDA.n1765 GNDA.n1764 0.028198
R21943 GNDA.n1771 GNDA.n1770 0.028198
R21944 GNDA.n1774 GNDA.n1773 0.028198
R21945 GNDA.n1780 GNDA.n1779 0.028198
R21946 GNDA.n1783 GNDA.n1782 0.028198
R21947 GNDA.n1789 GNDA.n1788 0.028198
R21948 GNDA.n1792 GNDA.n1791 0.028198
R21949 GNDA.n1798 GNDA.n1797 0.028198
R21950 GNDA.n1801 GNDA.n1800 0.028198
R21951 GNDA.n1807 GNDA.n1806 0.028198
R21952 GNDA.n1810 GNDA.n1809 0.028198
R21953 GNDA.n4278 GNDA.n1623 0.028198
R21954 GNDA.n4274 GNDA.n1622 0.028198
R21955 GNDA.n4264 GNDA.n1620 0.028198
R21956 GNDA.n4258 GNDA.n1619 0.028198
R21957 GNDA.n4248 GNDA.n1617 0.028198
R21958 GNDA.n4244 GNDA.n1616 0.028198
R21959 GNDA.n4234 GNDA.n1614 0.028198
R21960 GNDA.n4228 GNDA.n1613 0.028198
R21961 GNDA.n4218 GNDA.n1611 0.028198
R21962 GNDA.n4214 GNDA.n1610 0.028198
R21963 GNDA.n4204 GNDA.n1608 0.028198
R21964 GNDA.n4198 GNDA.n1607 0.028198
R21965 GNDA.n4188 GNDA.n1605 0.028198
R21966 GNDA.n4184 GNDA.n1604 0.028198
R21967 GNDA.n4174 GNDA.n1602 0.028198
R21968 GNDA.n4168 GNDA.n1601 0.028198
R21969 GNDA.n4444 GNDA.n4307 0.028198
R21970 GNDA.n4440 GNDA.n4306 0.028198
R21971 GNDA.n4430 GNDA.n4304 0.028198
R21972 GNDA.n4424 GNDA.n4303 0.028198
R21973 GNDA.n4414 GNDA.n4301 0.028198
R21974 GNDA.n4410 GNDA.n4300 0.028198
R21975 GNDA.n4400 GNDA.n4298 0.028198
R21976 GNDA.n4394 GNDA.n4297 0.028198
R21977 GNDA.n4384 GNDA.n4295 0.028198
R21978 GNDA.n4380 GNDA.n4294 0.028198
R21979 GNDA.n4370 GNDA.n4292 0.028198
R21980 GNDA.n4364 GNDA.n4291 0.028198
R21981 GNDA.n4354 GNDA.n4289 0.028198
R21982 GNDA.n4350 GNDA.n4288 0.028198
R21983 GNDA.n4340 GNDA.n4286 0.028198
R21984 GNDA.n4334 GNDA.n4285 0.028198
R21985 GNDA.n4633 GNDA.n4496 0.028198
R21986 GNDA.n4629 GNDA.n4495 0.028198
R21987 GNDA.n4619 GNDA.n4493 0.028198
R21988 GNDA.n4613 GNDA.n4492 0.028198
R21989 GNDA.n4603 GNDA.n4490 0.028198
R21990 GNDA.n4599 GNDA.n4489 0.028198
R21991 GNDA.n4589 GNDA.n4487 0.028198
R21992 GNDA.n4583 GNDA.n4486 0.028198
R21993 GNDA.n4573 GNDA.n4484 0.028198
R21994 GNDA.n4569 GNDA.n4483 0.028198
R21995 GNDA.n4559 GNDA.n4481 0.028198
R21996 GNDA.n4553 GNDA.n4480 0.028198
R21997 GNDA.n4543 GNDA.n4478 0.028198
R21998 GNDA.n4539 GNDA.n4477 0.028198
R21999 GNDA.n4529 GNDA.n4475 0.028198
R22000 GNDA.n4523 GNDA.n4474 0.028198
R22001 GNDA.n4919 GNDA.n1395 0.028198
R22002 GNDA.n4915 GNDA.n1394 0.028198
R22003 GNDA.n4905 GNDA.n1392 0.028198
R22004 GNDA.n4899 GNDA.n1391 0.028198
R22005 GNDA.n4889 GNDA.n1389 0.028198
R22006 GNDA.n4885 GNDA.n1388 0.028198
R22007 GNDA.n4875 GNDA.n1386 0.028198
R22008 GNDA.n4869 GNDA.n1385 0.028198
R22009 GNDA.n4859 GNDA.n1383 0.028198
R22010 GNDA.n4855 GNDA.n1382 0.028198
R22011 GNDA.n4845 GNDA.n1380 0.028198
R22012 GNDA.n4839 GNDA.n1379 0.028198
R22013 GNDA.n4829 GNDA.n1377 0.028198
R22014 GNDA.n4825 GNDA.n1376 0.028198
R22015 GNDA.n4815 GNDA.n1374 0.028198
R22016 GNDA.n4809 GNDA.n1373 0.028198
R22017 GNDA.n5938 GNDA.n4971 0.028198
R22018 GNDA.n5934 GNDA.n4970 0.028198
R22019 GNDA.n5924 GNDA.n4968 0.028198
R22020 GNDA.n5918 GNDA.n4967 0.028198
R22021 GNDA.n5908 GNDA.n4965 0.028198
R22022 GNDA.n5904 GNDA.n4964 0.028198
R22023 GNDA.n5894 GNDA.n4962 0.028198
R22024 GNDA.n5888 GNDA.n4961 0.028198
R22025 GNDA.n5878 GNDA.n4959 0.028198
R22026 GNDA.n5874 GNDA.n4958 0.028198
R22027 GNDA.n5864 GNDA.n4956 0.028198
R22028 GNDA.n5858 GNDA.n4955 0.028198
R22029 GNDA.n5848 GNDA.n4953 0.028198
R22030 GNDA.n5844 GNDA.n4952 0.028198
R22031 GNDA.n5834 GNDA.n4950 0.028198
R22032 GNDA.n5828 GNDA.n4949 0.028198
R22033 GNDA.n5656 GNDA.n5019 0.028198
R22034 GNDA.n5652 GNDA.n5018 0.028198
R22035 GNDA.n5642 GNDA.n5016 0.028198
R22036 GNDA.n5636 GNDA.n5015 0.028198
R22037 GNDA.n5626 GNDA.n5013 0.028198
R22038 GNDA.n5622 GNDA.n5012 0.028198
R22039 GNDA.n5612 GNDA.n5010 0.028198
R22040 GNDA.n5606 GNDA.n5009 0.028198
R22041 GNDA.n5596 GNDA.n5007 0.028198
R22042 GNDA.n5592 GNDA.n5006 0.028198
R22043 GNDA.n5582 GNDA.n5004 0.028198
R22044 GNDA.n5576 GNDA.n5003 0.028198
R22045 GNDA.n5566 GNDA.n5001 0.028198
R22046 GNDA.n5562 GNDA.n5000 0.028198
R22047 GNDA.n5552 GNDA.n4998 0.028198
R22048 GNDA.n5546 GNDA.n4997 0.028198
R22049 GNDA.n5514 GNDA.n5043 0.028198
R22050 GNDA.n5510 GNDA.n5042 0.028198
R22051 GNDA.n5500 GNDA.n5040 0.028198
R22052 GNDA.n5494 GNDA.n5039 0.028198
R22053 GNDA.n5484 GNDA.n5037 0.028198
R22054 GNDA.n5480 GNDA.n5036 0.028198
R22055 GNDA.n5470 GNDA.n5034 0.028198
R22056 GNDA.n5464 GNDA.n5033 0.028198
R22057 GNDA.n5454 GNDA.n5031 0.028198
R22058 GNDA.n5450 GNDA.n5030 0.028198
R22059 GNDA.n5440 GNDA.n5028 0.028198
R22060 GNDA.n5434 GNDA.n5027 0.028198
R22061 GNDA.n5424 GNDA.n5025 0.028198
R22062 GNDA.n5420 GNDA.n5024 0.028198
R22063 GNDA.n5410 GNDA.n5022 0.028198
R22064 GNDA.n5404 GNDA.n5021 0.028198
R22065 GNDA.n5330 GNDA.n5329 0.028198
R22066 GNDA.n5333 GNDA.n5332 0.028198
R22067 GNDA.n5339 GNDA.n5338 0.028198
R22068 GNDA.n5342 GNDA.n5341 0.028198
R22069 GNDA.n5348 GNDA.n5347 0.028198
R22070 GNDA.n5351 GNDA.n5350 0.028198
R22071 GNDA.n5357 GNDA.n5356 0.028198
R22072 GNDA.n5360 GNDA.n5359 0.028198
R22073 GNDA.n5366 GNDA.n5365 0.028198
R22074 GNDA.n5369 GNDA.n5368 0.028198
R22075 GNDA.n5375 GNDA.n5374 0.028198
R22076 GNDA.n5378 GNDA.n5377 0.028198
R22077 GNDA.n5384 GNDA.n5383 0.028198
R22078 GNDA.n5387 GNDA.n5386 0.028198
R22079 GNDA.n5393 GNDA.n5392 0.028198
R22080 GNDA.n5396 GNDA.n5395 0.028198
R22081 GNDA.n5226 GNDA.n5094 0.028198
R22082 GNDA.n5222 GNDA.n5093 0.028198
R22083 GNDA.n5212 GNDA.n5091 0.028198
R22084 GNDA.n5206 GNDA.n5090 0.028198
R22085 GNDA.n5196 GNDA.n5088 0.028198
R22086 GNDA.n5192 GNDA.n5087 0.028198
R22087 GNDA.n5182 GNDA.n5085 0.028198
R22088 GNDA.n5176 GNDA.n5084 0.028198
R22089 GNDA.n5166 GNDA.n5082 0.028198
R22090 GNDA.n5162 GNDA.n5081 0.028198
R22091 GNDA.n5152 GNDA.n5079 0.028198
R22092 GNDA.n5146 GNDA.n5078 0.028198
R22093 GNDA.n5136 GNDA.n5076 0.028198
R22094 GNDA.n5132 GNDA.n5075 0.028198
R22095 GNDA.n5122 GNDA.n5073 0.028198
R22096 GNDA.n5072 GNDA.n5071 0.028198
R22097 GNDA.n3390 GNDA.n3389 0.028198
R22098 GNDA.n3393 GNDA.n3392 0.028198
R22099 GNDA.n3399 GNDA.n3398 0.028198
R22100 GNDA.n3402 GNDA.n3401 0.028198
R22101 GNDA.n3408 GNDA.n3407 0.028198
R22102 GNDA.n3411 GNDA.n3410 0.028198
R22103 GNDA.n3417 GNDA.n3416 0.028198
R22104 GNDA.n3420 GNDA.n3419 0.028198
R22105 GNDA.n3426 GNDA.n3425 0.028198
R22106 GNDA.n3429 GNDA.n3428 0.028198
R22107 GNDA.n3435 GNDA.n3434 0.028198
R22108 GNDA.n3438 GNDA.n3437 0.028198
R22109 GNDA.n3444 GNDA.n3443 0.028198
R22110 GNDA.n3447 GNDA.n3446 0.028198
R22111 GNDA.n3453 GNDA.n3452 0.028198
R22112 GNDA.n3456 GNDA.n3455 0.028198
R22113 GNDA.n3746 GNDA.n3609 0.028198
R22114 GNDA.n3742 GNDA.n3608 0.028198
R22115 GNDA.n3732 GNDA.n3606 0.028198
R22116 GNDA.n3726 GNDA.n3605 0.028198
R22117 GNDA.n3716 GNDA.n3603 0.028198
R22118 GNDA.n3712 GNDA.n3602 0.028198
R22119 GNDA.n3702 GNDA.n3600 0.028198
R22120 GNDA.n3696 GNDA.n3599 0.028198
R22121 GNDA.n3686 GNDA.n3597 0.028198
R22122 GNDA.n3682 GNDA.n3596 0.028198
R22123 GNDA.n3672 GNDA.n3594 0.028198
R22124 GNDA.n3666 GNDA.n3593 0.028198
R22125 GNDA.n3656 GNDA.n3591 0.028198
R22126 GNDA.n3652 GNDA.n3590 0.028198
R22127 GNDA.n3642 GNDA.n3588 0.028198
R22128 GNDA.n3636 GNDA.n3587 0.028198
R22129 GNDA.n1518 GNDA.n1517 0.028198
R22130 GNDA.n1521 GNDA.n1520 0.028198
R22131 GNDA.n1527 GNDA.n1526 0.028198
R22132 GNDA.n1530 GNDA.n1529 0.028198
R22133 GNDA.n1536 GNDA.n1535 0.028198
R22134 GNDA.n1539 GNDA.n1538 0.028198
R22135 GNDA.n1545 GNDA.n1544 0.028198
R22136 GNDA.n1548 GNDA.n1547 0.028198
R22137 GNDA.n1554 GNDA.n1553 0.028198
R22138 GNDA.n1557 GNDA.n1556 0.028198
R22139 GNDA.n1563 GNDA.n1562 0.028198
R22140 GNDA.n1566 GNDA.n1565 0.028198
R22141 GNDA.n1572 GNDA.n1571 0.028198
R22142 GNDA.n1575 GNDA.n1574 0.028198
R22143 GNDA.n1581 GNDA.n1580 0.028198
R22144 GNDA.n1584 GNDA.n1583 0.028198
R22145 GNDA.n6075 GNDA.n4947 0.028198
R22146 GNDA.n6071 GNDA.n4946 0.028198
R22147 GNDA.n6061 GNDA.n4944 0.028198
R22148 GNDA.n6055 GNDA.n4943 0.028198
R22149 GNDA.n6045 GNDA.n4941 0.028198
R22150 GNDA.n6041 GNDA.n4940 0.028198
R22151 GNDA.n6031 GNDA.n4938 0.028198
R22152 GNDA.n6025 GNDA.n4937 0.028198
R22153 GNDA.n6015 GNDA.n4935 0.028198
R22154 GNDA.n6011 GNDA.n4934 0.028198
R22155 GNDA.n6001 GNDA.n4932 0.028198
R22156 GNDA.n5995 GNDA.n4931 0.028198
R22157 GNDA.n5985 GNDA.n4929 0.028198
R22158 GNDA.n5981 GNDA.n4928 0.028198
R22159 GNDA.n5971 GNDA.n4926 0.028198
R22160 GNDA.n4925 GNDA.n1370 0.028198
R22161 GNDA.n2787 GNDA.n2485 0.028198
R22162 GNDA.n2656 GNDA.n2484 0.028198
R22163 GNDA.n2660 GNDA.n2482 0.028198
R22164 GNDA.n2771 GNDA.n2481 0.028198
R22165 GNDA.n2763 GNDA.n2479 0.028198
R22166 GNDA.n2668 GNDA.n2478 0.028198
R22167 GNDA.n2672 GNDA.n2476 0.028198
R22168 GNDA.n2747 GNDA.n2475 0.028198
R22169 GNDA.n2739 GNDA.n2473 0.028198
R22170 GNDA.n2680 GNDA.n2472 0.028198
R22171 GNDA.n2684 GNDA.n2470 0.028198
R22172 GNDA.n2723 GNDA.n2469 0.028198
R22173 GNDA.n2715 GNDA.n2467 0.028198
R22174 GNDA.n2692 GNDA.n2466 0.028198
R22175 GNDA.n2696 GNDA.n2464 0.028198
R22176 GNDA.n2699 GNDA.n2463 0.028198
R22177 GNDA.n5797 GNDA.n4995 0.028198
R22178 GNDA.n5793 GNDA.n4994 0.028198
R22179 GNDA.n5783 GNDA.n4992 0.028198
R22180 GNDA.n5777 GNDA.n4991 0.028198
R22181 GNDA.n5767 GNDA.n4989 0.028198
R22182 GNDA.n5763 GNDA.n4988 0.028198
R22183 GNDA.n5753 GNDA.n4986 0.028198
R22184 GNDA.n5747 GNDA.n4985 0.028198
R22185 GNDA.n5737 GNDA.n4983 0.028198
R22186 GNDA.n5733 GNDA.n4982 0.028198
R22187 GNDA.n5723 GNDA.n4980 0.028198
R22188 GNDA.n5717 GNDA.n4979 0.028198
R22189 GNDA.n5707 GNDA.n4977 0.028198
R22190 GNDA.n5703 GNDA.n4976 0.028198
R22191 GNDA.n5693 GNDA.n4974 0.028198
R22192 GNDA.n5687 GNDA.n4973 0.028198
R22193 GNDA.n4770 GNDA.n4472 0.028198
R22194 GNDA.n4766 GNDA.n4471 0.028198
R22195 GNDA.n4756 GNDA.n4469 0.028198
R22196 GNDA.n4750 GNDA.n4468 0.028198
R22197 GNDA.n4740 GNDA.n4466 0.028198
R22198 GNDA.n4736 GNDA.n4465 0.028198
R22199 GNDA.n4726 GNDA.n4463 0.028198
R22200 GNDA.n4720 GNDA.n4462 0.028198
R22201 GNDA.n4710 GNDA.n4460 0.028198
R22202 GNDA.n4706 GNDA.n4459 0.028198
R22203 GNDA.n4696 GNDA.n4457 0.028198
R22204 GNDA.n4690 GNDA.n4456 0.028198
R22205 GNDA.n4680 GNDA.n4454 0.028198
R22206 GNDA.n4676 GNDA.n4453 0.028198
R22207 GNDA.n4666 GNDA.n4451 0.028198
R22208 GNDA.n4450 GNDA.n1598 0.028198
R22209 GNDA.n6357 GNDA.n6288 0.028198
R22210 GNDA.n6350 GNDA.n6289 0.028198
R22211 GNDA.n6346 GNDA.n6291 0.028198
R22212 GNDA.n6373 GNDA.n6292 0.028198
R22213 GNDA.n6381 GNDA.n6294 0.028198
R22214 GNDA.n6338 GNDA.n6295 0.028198
R22215 GNDA.n6334 GNDA.n6297 0.028198
R22216 GNDA.n6397 GNDA.n6298 0.028198
R22217 GNDA.n6405 GNDA.n6300 0.028198
R22218 GNDA.n6326 GNDA.n6301 0.028198
R22219 GNDA.n6322 GNDA.n6303 0.028198
R22220 GNDA.n6421 GNDA.n6304 0.028198
R22221 GNDA.n6429 GNDA.n6306 0.028198
R22222 GNDA.n6314 GNDA.n6307 0.028198
R22223 GNDA.n6310 GNDA.n6309 0.028198
R22224 GNDA.n6445 GNDA.n360 0.028198
R22225 GNDA.n415 GNDA.n363 0.028198
R22226 GNDA.n419 GNDA.n364 0.028198
R22227 GNDA.n429 GNDA.n366 0.028198
R22228 GNDA.n435 GNDA.n367 0.028198
R22229 GNDA.n445 GNDA.n369 0.028198
R22230 GNDA.n449 GNDA.n370 0.028198
R22231 GNDA.n459 GNDA.n372 0.028198
R22232 GNDA.n465 GNDA.n373 0.028198
R22233 GNDA.n475 GNDA.n375 0.028198
R22234 GNDA.n479 GNDA.n376 0.028198
R22235 GNDA.n489 GNDA.n378 0.028198
R22236 GNDA.n495 GNDA.n379 0.028198
R22237 GNDA.n505 GNDA.n381 0.028198
R22238 GNDA.n509 GNDA.n382 0.028198
R22239 GNDA.n519 GNDA.n384 0.028198
R22240 GNDA.n386 GNDA.n385 0.028198
R22241 GNDA.n520 GNDA.n385 0.028198
R22242 GNDA.n516 GNDA.n384 0.028198
R22243 GNDA.n506 GNDA.n382 0.028198
R22244 GNDA.n500 GNDA.n381 0.028198
R22245 GNDA.n490 GNDA.n379 0.028198
R22246 GNDA.n486 GNDA.n378 0.028198
R22247 GNDA.n476 GNDA.n376 0.028198
R22248 GNDA.n470 GNDA.n375 0.028198
R22249 GNDA.n460 GNDA.n373 0.028198
R22250 GNDA.n456 GNDA.n372 0.028198
R22251 GNDA.n446 GNDA.n370 0.028198
R22252 GNDA.n440 GNDA.n369 0.028198
R22253 GNDA.n430 GNDA.n367 0.028198
R22254 GNDA.n426 GNDA.n366 0.028198
R22255 GNDA.n416 GNDA.n364 0.028198
R22256 GNDA.n410 GNDA.n363 0.028198
R22257 GNDA.n6445 GNDA.n6444 0.028198
R22258 GNDA.n6438 GNDA.n6309 0.028198
R22259 GNDA.n6430 GNDA.n6307 0.028198
R22260 GNDA.n6319 GNDA.n6306 0.028198
R22261 GNDA.n6323 GNDA.n6304 0.028198
R22262 GNDA.n6414 GNDA.n6303 0.028198
R22263 GNDA.n6406 GNDA.n6301 0.028198
R22264 GNDA.n6331 GNDA.n6300 0.028198
R22265 GNDA.n6335 GNDA.n6298 0.028198
R22266 GNDA.n6390 GNDA.n6297 0.028198
R22267 GNDA.n6382 GNDA.n6295 0.028198
R22268 GNDA.n6343 GNDA.n6294 0.028198
R22269 GNDA.n6347 GNDA.n6292 0.028198
R22270 GNDA.n6366 GNDA.n6291 0.028198
R22271 GNDA.n6358 GNDA.n6289 0.028198
R22272 GNDA.n6354 GNDA.n6288 0.028198
R22273 GNDA.n2358 GNDA.n1895 0.028198
R22274 GNDA.n2362 GNDA.n1903 0.028198
R22275 GNDA.n2367 GNDA.n1910 0.028198
R22276 GNDA.n2371 GNDA.n1918 0.028198
R22277 GNDA.n2376 GNDA.n1925 0.028198
R22278 GNDA.n2380 GNDA.n1933 0.028198
R22279 GNDA.n2385 GNDA.n1940 0.028198
R22280 GNDA.n2389 GNDA.n1948 0.028198
R22281 GNDA.n2389 GNDA.n1949 0.028198
R22282 GNDA.n2385 GNDA.n2384 0.028198
R22283 GNDA.n2380 GNDA.n1934 0.028198
R22284 GNDA.n2376 GNDA.n2375 0.028198
R22285 GNDA.n2371 GNDA.n1919 0.028198
R22286 GNDA.n2367 GNDA.n2366 0.028198
R22287 GNDA.n2362 GNDA.n1904 0.028198
R22288 GNDA.n2358 GNDA.n2357 0.028198
R22289 GNDA.n2359 GNDA.n1898 0.0262697
R22290 GNDA.n2361 GNDA.n1900 0.0262697
R22291 GNDA.n2364 GNDA.n1905 0.0262697
R22292 GNDA.n2365 GNDA.n1908 0.0262697
R22293 GNDA.n2368 GNDA.n1913 0.0262697
R22294 GNDA.n2370 GNDA.n1915 0.0262697
R22295 GNDA.n2373 GNDA.n1920 0.0262697
R22296 GNDA.n2374 GNDA.n1923 0.0262697
R22297 GNDA.n2377 GNDA.n1928 0.0262697
R22298 GNDA.n2379 GNDA.n1930 0.0262697
R22299 GNDA.n2382 GNDA.n1935 0.0262697
R22300 GNDA.n2383 GNDA.n1938 0.0262697
R22301 GNDA.n2386 GNDA.n1943 0.0262697
R22302 GNDA.n2388 GNDA.n1945 0.0262697
R22303 GNDA.n3217 GNDA.n1950 0.0262697
R22304 GNDA.n2388 GNDA.n2387 0.0262697
R22305 GNDA.n2386 GNDA.n1944 0.0262697
R22306 GNDA.n2383 GNDA.n1939 0.0262697
R22307 GNDA.n2382 GNDA.n2381 0.0262697
R22308 GNDA.n2379 GNDA.n2378 0.0262697
R22309 GNDA.n2377 GNDA.n1929 0.0262697
R22310 GNDA.n2374 GNDA.n1924 0.0262697
R22311 GNDA.n2373 GNDA.n2372 0.0262697
R22312 GNDA.n2370 GNDA.n2369 0.0262697
R22313 GNDA.n2368 GNDA.n1914 0.0262697
R22314 GNDA.n2365 GNDA.n1909 0.0262697
R22315 GNDA.n2364 GNDA.n2363 0.0262697
R22316 GNDA.n2361 GNDA.n2360 0.0262697
R22317 GNDA.n2359 GNDA.n1899 0.0262697
R22318 GNDA.n1894 GNDA.n1893 0.0262697
R22319 GNDA.n4675 GNDA.n4452 0.0243392
R22320 GNDA.n4689 GNDA.n4455 0.0243392
R22321 GNDA.n4705 GNDA.n4458 0.0243392
R22322 GNDA.n4719 GNDA.n4461 0.0243392
R22323 GNDA.n4735 GNDA.n4464 0.0243392
R22324 GNDA.n4749 GNDA.n4467 0.0243392
R22325 GNDA.n4765 GNDA.n4470 0.0243392
R22326 GNDA.n5702 GNDA.n4975 0.0243392
R22327 GNDA.n5716 GNDA.n4978 0.0243392
R22328 GNDA.n5732 GNDA.n4981 0.0243392
R22329 GNDA.n5746 GNDA.n4984 0.0243392
R22330 GNDA.n5762 GNDA.n4987 0.0243392
R22331 GNDA.n5776 GNDA.n4990 0.0243392
R22332 GNDA.n5792 GNDA.n4993 0.0243392
R22333 GNDA.n2691 GNDA.n2465 0.0243392
R22334 GNDA.n2722 GNDA.n2468 0.0243392
R22335 GNDA.n2679 GNDA.n2471 0.0243392
R22336 GNDA.n2746 GNDA.n2474 0.0243392
R22337 GNDA.n2667 GNDA.n2477 0.0243392
R22338 GNDA.n2770 GNDA.n2480 0.0243392
R22339 GNDA.n2655 GNDA.n2483 0.0243392
R22340 GNDA.n5980 GNDA.n4927 0.0243392
R22341 GNDA.n5994 GNDA.n4930 0.0243392
R22342 GNDA.n6010 GNDA.n4933 0.0243392
R22343 GNDA.n6024 GNDA.n4936 0.0243392
R22344 GNDA.n6040 GNDA.n4939 0.0243392
R22345 GNDA.n6054 GNDA.n4942 0.0243392
R22346 GNDA.n6070 GNDA.n4945 0.0243392
R22347 GNDA.n1577 GNDA.n1576 0.0243392
R22348 GNDA.n1568 GNDA.n1567 0.0243392
R22349 GNDA.n1559 GNDA.n1558 0.0243392
R22350 GNDA.n1550 GNDA.n1549 0.0243392
R22351 GNDA.n1541 GNDA.n1540 0.0243392
R22352 GNDA.n1532 GNDA.n1531 0.0243392
R22353 GNDA.n1523 GNDA.n1522 0.0243392
R22354 GNDA.n3651 GNDA.n3589 0.0243392
R22355 GNDA.n3665 GNDA.n3592 0.0243392
R22356 GNDA.n3681 GNDA.n3595 0.0243392
R22357 GNDA.n3695 GNDA.n3598 0.0243392
R22358 GNDA.n3711 GNDA.n3601 0.0243392
R22359 GNDA.n3725 GNDA.n3604 0.0243392
R22360 GNDA.n3741 GNDA.n3607 0.0243392
R22361 GNDA.n3449 GNDA.n3448 0.0243392
R22362 GNDA.n3440 GNDA.n3439 0.0243392
R22363 GNDA.n3431 GNDA.n3430 0.0243392
R22364 GNDA.n3422 GNDA.n3421 0.0243392
R22365 GNDA.n3413 GNDA.n3412 0.0243392
R22366 GNDA.n3404 GNDA.n3403 0.0243392
R22367 GNDA.n3395 GNDA.n3394 0.0243392
R22368 GNDA.n5131 GNDA.n5074 0.0243392
R22369 GNDA.n5145 GNDA.n5077 0.0243392
R22370 GNDA.n5161 GNDA.n5080 0.0243392
R22371 GNDA.n5175 GNDA.n5083 0.0243392
R22372 GNDA.n5191 GNDA.n5086 0.0243392
R22373 GNDA.n5205 GNDA.n5089 0.0243392
R22374 GNDA.n5221 GNDA.n5092 0.0243392
R22375 GNDA.n5389 GNDA.n5388 0.0243392
R22376 GNDA.n5380 GNDA.n5379 0.0243392
R22377 GNDA.n5371 GNDA.n5370 0.0243392
R22378 GNDA.n5362 GNDA.n5361 0.0243392
R22379 GNDA.n5353 GNDA.n5352 0.0243392
R22380 GNDA.n5344 GNDA.n5343 0.0243392
R22381 GNDA.n5335 GNDA.n5334 0.0243392
R22382 GNDA.n5419 GNDA.n5023 0.0243392
R22383 GNDA.n5433 GNDA.n5026 0.0243392
R22384 GNDA.n5449 GNDA.n5029 0.0243392
R22385 GNDA.n5463 GNDA.n5032 0.0243392
R22386 GNDA.n5479 GNDA.n5035 0.0243392
R22387 GNDA.n5493 GNDA.n5038 0.0243392
R22388 GNDA.n5509 GNDA.n5041 0.0243392
R22389 GNDA.n5561 GNDA.n4999 0.0243392
R22390 GNDA.n5575 GNDA.n5002 0.0243392
R22391 GNDA.n5591 GNDA.n5005 0.0243392
R22392 GNDA.n5605 GNDA.n5008 0.0243392
R22393 GNDA.n5621 GNDA.n5011 0.0243392
R22394 GNDA.n5635 GNDA.n5014 0.0243392
R22395 GNDA.n5651 GNDA.n5017 0.0243392
R22396 GNDA.n5843 GNDA.n4951 0.0243392
R22397 GNDA.n5857 GNDA.n4954 0.0243392
R22398 GNDA.n5873 GNDA.n4957 0.0243392
R22399 GNDA.n5887 GNDA.n4960 0.0243392
R22400 GNDA.n5903 GNDA.n4963 0.0243392
R22401 GNDA.n5917 GNDA.n4966 0.0243392
R22402 GNDA.n5933 GNDA.n4969 0.0243392
R22403 GNDA.n4824 GNDA.n1375 0.0243392
R22404 GNDA.n4838 GNDA.n1378 0.0243392
R22405 GNDA.n4854 GNDA.n1381 0.0243392
R22406 GNDA.n4868 GNDA.n1384 0.0243392
R22407 GNDA.n4884 GNDA.n1387 0.0243392
R22408 GNDA.n4898 GNDA.n1390 0.0243392
R22409 GNDA.n4914 GNDA.n1393 0.0243392
R22410 GNDA.n4538 GNDA.n4476 0.0243392
R22411 GNDA.n4552 GNDA.n4479 0.0243392
R22412 GNDA.n4568 GNDA.n4482 0.0243392
R22413 GNDA.n4582 GNDA.n4485 0.0243392
R22414 GNDA.n4598 GNDA.n4488 0.0243392
R22415 GNDA.n4612 GNDA.n4491 0.0243392
R22416 GNDA.n4628 GNDA.n4494 0.0243392
R22417 GNDA.n4349 GNDA.n4287 0.0243392
R22418 GNDA.n4363 GNDA.n4290 0.0243392
R22419 GNDA.n4379 GNDA.n4293 0.0243392
R22420 GNDA.n4393 GNDA.n4296 0.0243392
R22421 GNDA.n4409 GNDA.n4299 0.0243392
R22422 GNDA.n4423 GNDA.n4302 0.0243392
R22423 GNDA.n4439 GNDA.n4305 0.0243392
R22424 GNDA.n4183 GNDA.n1603 0.0243392
R22425 GNDA.n4197 GNDA.n1606 0.0243392
R22426 GNDA.n4213 GNDA.n1609 0.0243392
R22427 GNDA.n4227 GNDA.n1612 0.0243392
R22428 GNDA.n4243 GNDA.n1615 0.0243392
R22429 GNDA.n4257 GNDA.n1618 0.0243392
R22430 GNDA.n4273 GNDA.n1621 0.0243392
R22431 GNDA.n1803 GNDA.n1802 0.0243392
R22432 GNDA.n1794 GNDA.n1793 0.0243392
R22433 GNDA.n1785 GNDA.n1784 0.0243392
R22434 GNDA.n1776 GNDA.n1775 0.0243392
R22435 GNDA.n1767 GNDA.n1766 0.0243392
R22436 GNDA.n1758 GNDA.n1757 0.0243392
R22437 GNDA.n1749 GNDA.n1748 0.0243392
R22438 GNDA.n3840 GNDA.n3778 0.0243392
R22439 GNDA.n3854 GNDA.n3781 0.0243392
R22440 GNDA.n3870 GNDA.n3784 0.0243392
R22441 GNDA.n3884 GNDA.n3787 0.0243392
R22442 GNDA.n3900 GNDA.n3790 0.0243392
R22443 GNDA.n3914 GNDA.n3793 0.0243392
R22444 GNDA.n3930 GNDA.n3796 0.0243392
R22445 GNDA.n3977 GNDA.n3754 0.0243392
R22446 GNDA.n3991 GNDA.n3757 0.0243392
R22447 GNDA.n4007 GNDA.n3760 0.0243392
R22448 GNDA.n4021 GNDA.n3763 0.0243392
R22449 GNDA.n4037 GNDA.n3766 0.0243392
R22450 GNDA.n4051 GNDA.n3769 0.0243392
R22451 GNDA.n4067 GNDA.n3772 0.0243392
R22452 GNDA.n3485 GNDA.n1842 0.0243392
R22453 GNDA.n3499 GNDA.n1845 0.0243392
R22454 GNDA.n3515 GNDA.n1848 0.0243392
R22455 GNDA.n3529 GNDA.n1851 0.0243392
R22456 GNDA.n3545 GNDA.n1854 0.0243392
R22457 GNDA.n3559 GNDA.n1857 0.0243392
R22458 GNDA.n3575 GNDA.n1860 0.0243392
R22459 GNDA.n2550 GNDA.n2489 0.0243392
R22460 GNDA.n2564 GNDA.n2492 0.0243392
R22461 GNDA.n2580 GNDA.n2495 0.0243392
R22462 GNDA.n2594 GNDA.n2498 0.0243392
R22463 GNDA.n2610 GNDA.n2501 0.0243392
R22464 GNDA.n2624 GNDA.n2504 0.0243392
R22465 GNDA.n2640 GNDA.n2507 0.0243392
R22466 GNDA.n2833 GNDA.n2441 0.0243392
R22467 GNDA.n2847 GNDA.n2444 0.0243392
R22468 GNDA.n2863 GNDA.n2447 0.0243392
R22469 GNDA.n2877 GNDA.n2450 0.0243392
R22470 GNDA.n2893 GNDA.n2453 0.0243392
R22471 GNDA.n2907 GNDA.n2456 0.0243392
R22472 GNDA.n2923 GNDA.n2459 0.0243392
R22473 GNDA.n2974 GNDA.n2417 0.0243392
R22474 GNDA.n2988 GNDA.n2420 0.0243392
R22475 GNDA.n3004 GNDA.n2423 0.0243392
R22476 GNDA.n3018 GNDA.n2426 0.0243392
R22477 GNDA.n3034 GNDA.n2429 0.0243392
R22478 GNDA.n3048 GNDA.n2432 0.0243392
R22479 GNDA.n3064 GNDA.n2435 0.0243392
R22480 GNDA.n3115 GNDA.n2393 0.0243392
R22481 GNDA.n3129 GNDA.n2396 0.0243392
R22482 GNDA.n3145 GNDA.n2399 0.0243392
R22483 GNDA.n3159 GNDA.n2402 0.0243392
R22484 GNDA.n3175 GNDA.n2405 0.0243392
R22485 GNDA.n3189 GNDA.n2408 0.0243392
R22486 GNDA.n3205 GNDA.n2411 0.0243392
R22487 GNDA.n3200 GNDA.n2411 0.0243392
R22488 GNDA.n3186 GNDA.n2408 0.0243392
R22489 GNDA.n3170 GNDA.n2405 0.0243392
R22490 GNDA.n3156 GNDA.n2402 0.0243392
R22491 GNDA.n3140 GNDA.n2399 0.0243392
R22492 GNDA.n3126 GNDA.n2396 0.0243392
R22493 GNDA.n3110 GNDA.n2393 0.0243392
R22494 GNDA.n3059 GNDA.n2435 0.0243392
R22495 GNDA.n3045 GNDA.n2432 0.0243392
R22496 GNDA.n3029 GNDA.n2429 0.0243392
R22497 GNDA.n3015 GNDA.n2426 0.0243392
R22498 GNDA.n2999 GNDA.n2423 0.0243392
R22499 GNDA.n2985 GNDA.n2420 0.0243392
R22500 GNDA.n2969 GNDA.n2417 0.0243392
R22501 GNDA.n2918 GNDA.n2459 0.0243392
R22502 GNDA.n2904 GNDA.n2456 0.0243392
R22503 GNDA.n2888 GNDA.n2453 0.0243392
R22504 GNDA.n2874 GNDA.n2450 0.0243392
R22505 GNDA.n2858 GNDA.n2447 0.0243392
R22506 GNDA.n2844 GNDA.n2444 0.0243392
R22507 GNDA.n2828 GNDA.n2441 0.0243392
R22508 GNDA.n2635 GNDA.n2507 0.0243392
R22509 GNDA.n2621 GNDA.n2504 0.0243392
R22510 GNDA.n2605 GNDA.n2501 0.0243392
R22511 GNDA.n2591 GNDA.n2498 0.0243392
R22512 GNDA.n2575 GNDA.n2495 0.0243392
R22513 GNDA.n2561 GNDA.n2492 0.0243392
R22514 GNDA.n2545 GNDA.n2489 0.0243392
R22515 GNDA.n3570 GNDA.n1860 0.0243392
R22516 GNDA.n3556 GNDA.n1857 0.0243392
R22517 GNDA.n3540 GNDA.n1854 0.0243392
R22518 GNDA.n3526 GNDA.n1851 0.0243392
R22519 GNDA.n3510 GNDA.n1848 0.0243392
R22520 GNDA.n3496 GNDA.n1845 0.0243392
R22521 GNDA.n3480 GNDA.n1842 0.0243392
R22522 GNDA.n4062 GNDA.n3772 0.0243392
R22523 GNDA.n4048 GNDA.n3769 0.0243392
R22524 GNDA.n4032 GNDA.n3766 0.0243392
R22525 GNDA.n4018 GNDA.n3763 0.0243392
R22526 GNDA.n4002 GNDA.n3760 0.0243392
R22527 GNDA.n3988 GNDA.n3757 0.0243392
R22528 GNDA.n3972 GNDA.n3754 0.0243392
R22529 GNDA.n3925 GNDA.n3796 0.0243392
R22530 GNDA.n3911 GNDA.n3793 0.0243392
R22531 GNDA.n3895 GNDA.n3790 0.0243392
R22532 GNDA.n3881 GNDA.n3787 0.0243392
R22533 GNDA.n3865 GNDA.n3784 0.0243392
R22534 GNDA.n3851 GNDA.n3781 0.0243392
R22535 GNDA.n3835 GNDA.n3778 0.0243392
R22536 GNDA.n1750 GNDA.n1749 0.0243392
R22537 GNDA.n1759 GNDA.n1758 0.0243392
R22538 GNDA.n1768 GNDA.n1767 0.0243392
R22539 GNDA.n1777 GNDA.n1776 0.0243392
R22540 GNDA.n1786 GNDA.n1785 0.0243392
R22541 GNDA.n1795 GNDA.n1794 0.0243392
R22542 GNDA.n1804 GNDA.n1803 0.0243392
R22543 GNDA.n4268 GNDA.n1621 0.0243392
R22544 GNDA.n4254 GNDA.n1618 0.0243392
R22545 GNDA.n4238 GNDA.n1615 0.0243392
R22546 GNDA.n4224 GNDA.n1612 0.0243392
R22547 GNDA.n4208 GNDA.n1609 0.0243392
R22548 GNDA.n4194 GNDA.n1606 0.0243392
R22549 GNDA.n4178 GNDA.n1603 0.0243392
R22550 GNDA.n4434 GNDA.n4305 0.0243392
R22551 GNDA.n4420 GNDA.n4302 0.0243392
R22552 GNDA.n4404 GNDA.n4299 0.0243392
R22553 GNDA.n4390 GNDA.n4296 0.0243392
R22554 GNDA.n4374 GNDA.n4293 0.0243392
R22555 GNDA.n4360 GNDA.n4290 0.0243392
R22556 GNDA.n4344 GNDA.n4287 0.0243392
R22557 GNDA.n4623 GNDA.n4494 0.0243392
R22558 GNDA.n4609 GNDA.n4491 0.0243392
R22559 GNDA.n4593 GNDA.n4488 0.0243392
R22560 GNDA.n4579 GNDA.n4485 0.0243392
R22561 GNDA.n4563 GNDA.n4482 0.0243392
R22562 GNDA.n4549 GNDA.n4479 0.0243392
R22563 GNDA.n4533 GNDA.n4476 0.0243392
R22564 GNDA.n4909 GNDA.n1393 0.0243392
R22565 GNDA.n4895 GNDA.n1390 0.0243392
R22566 GNDA.n4879 GNDA.n1387 0.0243392
R22567 GNDA.n4865 GNDA.n1384 0.0243392
R22568 GNDA.n4849 GNDA.n1381 0.0243392
R22569 GNDA.n4835 GNDA.n1378 0.0243392
R22570 GNDA.n4819 GNDA.n1375 0.0243392
R22571 GNDA.n5928 GNDA.n4969 0.0243392
R22572 GNDA.n5914 GNDA.n4966 0.0243392
R22573 GNDA.n5898 GNDA.n4963 0.0243392
R22574 GNDA.n5884 GNDA.n4960 0.0243392
R22575 GNDA.n5868 GNDA.n4957 0.0243392
R22576 GNDA.n5854 GNDA.n4954 0.0243392
R22577 GNDA.n5838 GNDA.n4951 0.0243392
R22578 GNDA.n5646 GNDA.n5017 0.0243392
R22579 GNDA.n5632 GNDA.n5014 0.0243392
R22580 GNDA.n5616 GNDA.n5011 0.0243392
R22581 GNDA.n5602 GNDA.n5008 0.0243392
R22582 GNDA.n5586 GNDA.n5005 0.0243392
R22583 GNDA.n5572 GNDA.n5002 0.0243392
R22584 GNDA.n5556 GNDA.n4999 0.0243392
R22585 GNDA.n5504 GNDA.n5041 0.0243392
R22586 GNDA.n5490 GNDA.n5038 0.0243392
R22587 GNDA.n5474 GNDA.n5035 0.0243392
R22588 GNDA.n5460 GNDA.n5032 0.0243392
R22589 GNDA.n5444 GNDA.n5029 0.0243392
R22590 GNDA.n5430 GNDA.n5026 0.0243392
R22591 GNDA.n5414 GNDA.n5023 0.0243392
R22592 GNDA.n5336 GNDA.n5335 0.0243392
R22593 GNDA.n5345 GNDA.n5344 0.0243392
R22594 GNDA.n5354 GNDA.n5353 0.0243392
R22595 GNDA.n5363 GNDA.n5362 0.0243392
R22596 GNDA.n5372 GNDA.n5371 0.0243392
R22597 GNDA.n5381 GNDA.n5380 0.0243392
R22598 GNDA.n5390 GNDA.n5389 0.0243392
R22599 GNDA.n5216 GNDA.n5092 0.0243392
R22600 GNDA.n5202 GNDA.n5089 0.0243392
R22601 GNDA.n5186 GNDA.n5086 0.0243392
R22602 GNDA.n5172 GNDA.n5083 0.0243392
R22603 GNDA.n5156 GNDA.n5080 0.0243392
R22604 GNDA.n5142 GNDA.n5077 0.0243392
R22605 GNDA.n5126 GNDA.n5074 0.0243392
R22606 GNDA.n3396 GNDA.n3395 0.0243392
R22607 GNDA.n3405 GNDA.n3404 0.0243392
R22608 GNDA.n3414 GNDA.n3413 0.0243392
R22609 GNDA.n3423 GNDA.n3422 0.0243392
R22610 GNDA.n3432 GNDA.n3431 0.0243392
R22611 GNDA.n3441 GNDA.n3440 0.0243392
R22612 GNDA.n3450 GNDA.n3449 0.0243392
R22613 GNDA.n3736 GNDA.n3607 0.0243392
R22614 GNDA.n3722 GNDA.n3604 0.0243392
R22615 GNDA.n3706 GNDA.n3601 0.0243392
R22616 GNDA.n3692 GNDA.n3598 0.0243392
R22617 GNDA.n3676 GNDA.n3595 0.0243392
R22618 GNDA.n3662 GNDA.n3592 0.0243392
R22619 GNDA.n3646 GNDA.n3589 0.0243392
R22620 GNDA.n1524 GNDA.n1523 0.0243392
R22621 GNDA.n1533 GNDA.n1532 0.0243392
R22622 GNDA.n1542 GNDA.n1541 0.0243392
R22623 GNDA.n1551 GNDA.n1550 0.0243392
R22624 GNDA.n1560 GNDA.n1559 0.0243392
R22625 GNDA.n1569 GNDA.n1568 0.0243392
R22626 GNDA.n1578 GNDA.n1577 0.0243392
R22627 GNDA.n6065 GNDA.n4945 0.0243392
R22628 GNDA.n6051 GNDA.n4942 0.0243392
R22629 GNDA.n6035 GNDA.n4939 0.0243392
R22630 GNDA.n6021 GNDA.n4936 0.0243392
R22631 GNDA.n6005 GNDA.n4933 0.0243392
R22632 GNDA.n5991 GNDA.n4930 0.0243392
R22633 GNDA.n5975 GNDA.n4927 0.0243392
R22634 GNDA.n2779 GNDA.n2483 0.0243392
R22635 GNDA.n2664 GNDA.n2480 0.0243392
R22636 GNDA.n2755 GNDA.n2477 0.0243392
R22637 GNDA.n2676 GNDA.n2474 0.0243392
R22638 GNDA.n2731 GNDA.n2471 0.0243392
R22639 GNDA.n2688 GNDA.n2468 0.0243392
R22640 GNDA.n2707 GNDA.n2465 0.0243392
R22641 GNDA.n5787 GNDA.n4993 0.0243392
R22642 GNDA.n5773 GNDA.n4990 0.0243392
R22643 GNDA.n5757 GNDA.n4987 0.0243392
R22644 GNDA.n5743 GNDA.n4984 0.0243392
R22645 GNDA.n5727 GNDA.n4981 0.0243392
R22646 GNDA.n5713 GNDA.n4978 0.0243392
R22647 GNDA.n5697 GNDA.n4975 0.0243392
R22648 GNDA.n4760 GNDA.n4470 0.0243392
R22649 GNDA.n4746 GNDA.n4467 0.0243392
R22650 GNDA.n4730 GNDA.n4464 0.0243392
R22651 GNDA.n4716 GNDA.n4461 0.0243392
R22652 GNDA.n4700 GNDA.n4458 0.0243392
R22653 GNDA.n4686 GNDA.n4455 0.0243392
R22654 GNDA.n4670 GNDA.n4452 0.0243392
R22655 GNDA.n6365 GNDA.n6290 0.0243392
R22656 GNDA.n6342 GNDA.n6293 0.0243392
R22657 GNDA.n6389 GNDA.n6296 0.0243392
R22658 GNDA.n6330 GNDA.n6299 0.0243392
R22659 GNDA.n6413 GNDA.n6302 0.0243392
R22660 GNDA.n6318 GNDA.n6305 0.0243392
R22661 GNDA.n6437 GNDA.n6308 0.0243392
R22662 GNDA.n425 GNDA.n365 0.0243392
R22663 GNDA.n439 GNDA.n368 0.0243392
R22664 GNDA.n455 GNDA.n371 0.0243392
R22665 GNDA.n469 GNDA.n374 0.0243392
R22666 GNDA.n485 GNDA.n377 0.0243392
R22667 GNDA.n499 GNDA.n380 0.0243392
R22668 GNDA.n515 GNDA.n383 0.0243392
R22669 GNDA.n510 GNDA.n383 0.0243392
R22670 GNDA.n496 GNDA.n380 0.0243392
R22671 GNDA.n480 GNDA.n377 0.0243392
R22672 GNDA.n466 GNDA.n374 0.0243392
R22673 GNDA.n450 GNDA.n371 0.0243392
R22674 GNDA.n436 GNDA.n368 0.0243392
R22675 GNDA.n420 GNDA.n365 0.0243392
R22676 GNDA.n6315 GNDA.n6308 0.0243392
R22677 GNDA.n6422 GNDA.n6305 0.0243392
R22678 GNDA.n6327 GNDA.n6302 0.0243392
R22679 GNDA.n6398 GNDA.n6299 0.0243392
R22680 GNDA.n6339 GNDA.n6296 0.0243392
R22681 GNDA.n6374 GNDA.n6293 0.0243392
R22682 GNDA.n6351 GNDA.n6290 0.0243392
R22683 GNDA.n2228 GNDA.n2227 0.00586094
R22684 GNDA.n3216 GNDA.n3215 0.00564062
R22685 GNDA.n3215 GNDA.n3074 0.00564062
R22686 GNDA.n3074 GNDA.n2933 0.00564062
R22687 GNDA.n2933 GNDA.n2792 0.00564062
R22688 GNDA.n2792 GNDA.n2650 0.00564062
R22689 GNDA.n2650 GNDA.n1838 0.00564062
R22690 GNDA.n3585 GNDA.n1838 0.00564062
R22691 GNDA.n3751 GNDA.n3585 0.00564062
R22692 GNDA.n4077 GNDA.n3751 0.00564062
R22693 GNDA.n4077 GNDA.n3940 0.00564062
R22694 GNDA.n3940 GNDA.n1599 0.00564062
R22695 GNDA.n4283 GNDA.n1599 0.00564062
R22696 GNDA.n4449 GNDA.n4283 0.00564062
R22697 GNDA.n4775 GNDA.n4449 0.00564062
R22698 GNDA.n4775 GNDA.n4638 0.00564062
R22699 GNDA.n4638 GNDA.n1371 0.00564062
R22700 GNDA.n4924 GNDA.n1371 0.00564062
R22701 GNDA.n6080 GNDA.n4924 0.00564062
R22702 GNDA.n6080 GNDA.n5943 0.00564062
R22703 GNDA.n5943 GNDA.n5802 0.00564062
R22704 GNDA.n5802 GNDA.n5661 0.00564062
R22705 GNDA.n5661 GNDA.n5519 0.00564062
R22706 GNDA.n5519 GNDA.n5044 0.00564062
R22707 GNDA.n5231 GNDA.n5044 0.00564062
R22708 GNDA.n2354 GNDA.n2320 0.00189531
R22709 GNDA.n2352 GNDA.n2320 0.00189531
R22710 GNDA.n2226 GNDA.n2164 0.00189531
R22711 GNDA.n2164 GNDA.n2134 0.00189531
R22712 GNDA.n2301 GNDA.n2267 0.00188102
R22713 GNDA.n2293 GNDA.n2271 0.00188102
R22714 GNDA.n2285 GNDA.n2275 0.00188102
R22715 GNDA.n2152 GNDA.n2108 0.00188102
R22716 GNDA.n2156 GNDA.n2112 0.00188102
R22717 GNDA.n2160 GNDA.n2116 0.00188102
R22718 GNDA.n2183 GNDA.n2148 0.00188102
R22719 GNDA.n2189 GNDA.n2146 0.00188102
R22720 GNDA.n2195 GNDA.n2144 0.00188102
R22721 GNDA.n2201 GNDA.n2142 0.00188102
R22722 GNDA.n2207 GNDA.n2140 0.00188102
R22723 GNDA.n2213 GNDA.n2138 0.00188102
R22724 GNDA.n2219 GNDA.n2136 0.00188102
R22725 GNDA.n2054 GNDA.n2010 0.00188102
R22726 GNDA.n2052 GNDA.n2008 0.00188102
R22727 GNDA.n2050 GNDA.n2006 0.00188102
R22728 GNDA.n2048 GNDA.n2004 0.00188102
R22729 GNDA.n2046 GNDA.n2002 0.00188102
R22730 GNDA.n2044 GNDA.n2000 0.00188102
R22731 GNDA.n2042 GNDA.n1998 0.00188102
R22732 GNDA.n2335 GNDA.n1965 0.00188102
R22733 GNDA.n2333 GNDA.n1963 0.00188102
R22734 GNDA.n2331 GNDA.n1961 0.00188102
R22735 GNDA.n2329 GNDA.n1959 0.00188102
R22736 GNDA.n2327 GNDA.n1957 0.00188102
R22737 GNDA.n2325 GNDA.n1955 0.00188102
R22738 GNDA.n2323 GNDA.n1953 0.00188102
R22739 GNDA.n2160 GNDA.n2123 0.00188102
R22740 GNDA.n2156 GNDA.n2127 0.00188102
R22741 GNDA.n2152 GNDA.n2131 0.00188102
R22742 GNDA.n2184 GNDA.n2183 0.00188102
R22743 GNDA.n2190 GNDA.n2189 0.00188102
R22744 GNDA.n2196 GNDA.n2195 0.00188102
R22745 GNDA.n2202 GNDA.n2201 0.00188102
R22746 GNDA.n2208 GNDA.n2207 0.00188102
R22747 GNDA.n2214 GNDA.n2213 0.00188102
R22748 GNDA.n2220 GNDA.n2219 0.00188102
R22749 GNDA.n2286 GNDA.n2285 0.00188102
R22750 GNDA.n2294 GNDA.n2293 0.00188102
R22751 GNDA.n2302 GNDA.n2301 0.00188102
R22752 GNDA.n2335 GNDA.n2250 0.00188102
R22753 GNDA.n2333 GNDA.n2252 0.00188102
R22754 GNDA.n2331 GNDA.n2254 0.00188102
R22755 GNDA.n2329 GNDA.n2256 0.00188102
R22756 GNDA.n2327 GNDA.n2258 0.00188102
R22757 GNDA.n2325 GNDA.n2260 0.00188102
R22758 GNDA.n2323 GNDA.n2262 0.00188102
R22759 GNDA.n2015 GNDA.n1969 0.00188102
R22760 GNDA.n2019 GNDA.n1973 0.00188102
R22761 GNDA.n2023 GNDA.n1977 0.00188102
R22762 GNDA.n2023 GNDA.n1985 0.00188102
R22763 GNDA.n2019 GNDA.n1989 0.00188102
R22764 GNDA.n2015 GNDA.n1993 0.00188102
R22765 GNDA.n2054 GNDA.n2028 0.00188102
R22766 GNDA.n2052 GNDA.n2030 0.00188102
R22767 GNDA.n2050 GNDA.n2032 0.00188102
R22768 GNDA.n2048 GNDA.n2034 0.00188102
R22769 GNDA.n2046 GNDA.n2036 0.00188102
R22770 GNDA.n2044 GNDA.n2038 0.00188102
R22771 GNDA.n2042 GNDA.n2040 0.00188102
R22772 GNDA.n2337 GNDA.n2265 0.00173422
R22773 GNDA.n2337 GNDA.n2336 0.00173422
R22774 GNDA.n2339 GNDA.n2266 0.00173422
R22775 GNDA.n2342 GNDA.n2269 0.00173422
R22776 GNDA.n2297 GNDA.n2269 0.00173422
R22777 GNDA.n2343 GNDA.n2270 0.00173422
R22778 GNDA.n2346 GNDA.n2273 0.00173422
R22779 GNDA.n2289 GNDA.n2273 0.00173422
R22780 GNDA.n2347 GNDA.n2274 0.00173422
R22781 GNDA.n2350 GNDA.n2277 0.00173422
R22782 GNDA.n2281 GNDA.n2277 0.00173422
R22783 GNDA.n2351 GNDA.n2278 0.00173422
R22784 GNDA.n2166 GNDA.n2106 0.00173422
R22785 GNDA.n2150 GNDA.n2106 0.00173422
R22786 GNDA.n2167 GNDA.n2107 0.00173422
R22787 GNDA.n2170 GNDA.n2110 0.00173422
R22788 GNDA.n2154 GNDA.n2110 0.00173422
R22789 GNDA.n2171 GNDA.n2111 0.00173422
R22790 GNDA.n2174 GNDA.n2114 0.00173422
R22791 GNDA.n2158 GNDA.n2114 0.00173422
R22792 GNDA.n2175 GNDA.n2115 0.00173422
R22793 GNDA.n2178 GNDA.n2118 0.00173422
R22794 GNDA.n2162 GNDA.n2118 0.00173422
R22795 GNDA.n2179 GNDA.n2119 0.00173422
R22796 GNDA.n2180 GNDA.n2149 0.00173422
R22797 GNDA.n2186 GNDA.n2147 0.00173422
R22798 GNDA.n2192 GNDA.n2145 0.00173422
R22799 GNDA.n2198 GNDA.n2143 0.00173422
R22800 GNDA.n2204 GNDA.n2141 0.00173422
R22801 GNDA.n2210 GNDA.n2139 0.00173422
R22802 GNDA.n2216 GNDA.n2137 0.00173422
R22803 GNDA.n2222 GNDA.n2135 0.00173422
R22804 GNDA.n2055 GNDA.n2012 0.00173422
R22805 GNDA.n2053 GNDA.n2009 0.00173422
R22806 GNDA.n2051 GNDA.n2007 0.00173422
R22807 GNDA.n2049 GNDA.n2005 0.00173422
R22808 GNDA.n2047 GNDA.n2003 0.00173422
R22809 GNDA.n2045 GNDA.n2001 0.00173422
R22810 GNDA.n2043 GNDA.n1999 0.00173422
R22811 GNDA.n2057 GNDA.n1997 0.00173422
R22812 GNDA.n2338 GNDA.n1966 0.00173422
R22813 GNDA.n2334 GNDA.n1964 0.00173422
R22814 GNDA.n2332 GNDA.n1962 0.00173422
R22815 GNDA.n2330 GNDA.n1960 0.00173422
R22816 GNDA.n2328 GNDA.n1958 0.00173422
R22817 GNDA.n2326 GNDA.n1956 0.00173422
R22818 GNDA.n2324 GNDA.n1954 0.00173422
R22819 GNDA.n2322 GNDA.n1952 0.00173422
R22820 GNDA.n2162 GNDA.n2121 0.00173422
R22821 GNDA.n2158 GNDA.n2125 0.00173422
R22822 GNDA.n2154 GNDA.n2129 0.00173422
R22823 GNDA.n2150 GNDA.n2133 0.00173422
R22824 GNDA.n2181 GNDA.n2180 0.00173422
R22825 GNDA.n2179 GNDA.n2121 0.00173422
R22826 GNDA.n2178 GNDA.n2122 0.00173422
R22827 GNDA.n2175 GNDA.n2125 0.00173422
R22828 GNDA.n2174 GNDA.n2126 0.00173422
R22829 GNDA.n2171 GNDA.n2129 0.00173422
R22830 GNDA.n2170 GNDA.n2130 0.00173422
R22831 GNDA.n2167 GNDA.n2133 0.00173422
R22832 GNDA.n2166 GNDA.n2134 0.00173422
R22833 GNDA.n2187 GNDA.n2186 0.00173422
R22834 GNDA.n2193 GNDA.n2192 0.00173422
R22835 GNDA.n2199 GNDA.n2198 0.00173422
R22836 GNDA.n2205 GNDA.n2204 0.00173422
R22837 GNDA.n2211 GNDA.n2210 0.00173422
R22838 GNDA.n2217 GNDA.n2216 0.00173422
R22839 GNDA.n2225 GNDA.n2222 0.00173422
R22840 GNDA.n2282 GNDA.n2281 0.00173422
R22841 GNDA.n2290 GNDA.n2289 0.00173422
R22842 GNDA.n2298 GNDA.n2297 0.00173422
R22843 GNDA.n2336 GNDA.n2305 0.00173422
R22844 GNDA.n2351 GNDA.n2282 0.00173422
R22845 GNDA.n2350 GNDA.n2284 0.00173422
R22846 GNDA.n2347 GNDA.n2290 0.00173422
R22847 GNDA.n2346 GNDA.n2292 0.00173422
R22848 GNDA.n2343 GNDA.n2298 0.00173422
R22849 GNDA.n2342 GNDA.n2300 0.00173422
R22850 GNDA.n2339 GNDA.n2305 0.00173422
R22851 GNDA.n2353 GNDA.n2338 0.00173422
R22852 GNDA.n2334 GNDA.n2251 0.00173422
R22853 GNDA.n2332 GNDA.n2253 0.00173422
R22854 GNDA.n2330 GNDA.n2255 0.00173422
R22855 GNDA.n2328 GNDA.n2257 0.00173422
R22856 GNDA.n2326 GNDA.n2259 0.00173422
R22857 GNDA.n2324 GNDA.n2261 0.00173422
R22858 GNDA.n2322 GNDA.n2263 0.00173422
R22859 GNDA.n2352 GNDA.n2265 0.00173422
R22860 GNDA.n2245 GNDA.n2244 0.00173422
R22861 GNDA.n2072 GNDA.n2058 0.00173422
R22862 GNDA.n2229 GNDA.n1995 0.00173422
R22863 GNDA.n2232 GNDA.n1992 0.00173422
R22864 GNDA.n2017 GNDA.n1971 0.00173422
R22865 GNDA.n2233 GNDA.n1991 0.00173422
R22866 GNDA.n2236 GNDA.n1988 0.00173422
R22867 GNDA.n2021 GNDA.n1975 0.00173422
R22868 GNDA.n2237 GNDA.n1987 0.00173422
R22869 GNDA.n2240 GNDA.n1984 0.00173422
R22870 GNDA.n2025 GNDA.n1979 0.00173422
R22871 GNDA.n2241 GNDA.n1983 0.00173422
R22872 GNDA.n2241 GNDA.n1980 0.00173422
R22873 GNDA.n2240 GNDA.n1979 0.00173422
R22874 GNDA.n2237 GNDA.n1976 0.00173422
R22875 GNDA.n2236 GNDA.n1975 0.00173422
R22876 GNDA.n2233 GNDA.n1972 0.00173422
R22877 GNDA.n2232 GNDA.n1971 0.00173422
R22878 GNDA.n2229 GNDA.n1968 0.00173422
R22879 GNDA.n2244 GNDA.n2072 0.00173422
R22880 GNDA.n2025 GNDA.n1983 0.00173422
R22881 GNDA.n2021 GNDA.n1987 0.00173422
R22882 GNDA.n2017 GNDA.n1991 0.00173422
R22883 GNDA.n2058 GNDA.n1995 0.00173422
R22884 GNDA.n2055 GNDA.n2026 0.00173422
R22885 GNDA.n2053 GNDA.n2029 0.00173422
R22886 GNDA.n2051 GNDA.n2031 0.00173422
R22887 GNDA.n2049 GNDA.n2033 0.00173422
R22888 GNDA.n2047 GNDA.n2035 0.00173422
R22889 GNDA.n2045 GNDA.n2037 0.00173422
R22890 GNDA.n2043 GNDA.n2039 0.00173422
R22891 GNDA.n2246 GNDA.n2057 0.00173422
R22892 GNDA.n2303 GNDA.n2266 0.00169751
R22893 GNDA.n2340 GNDA.n2267 0.00169751
R22894 GNDA.n2341 GNDA.n2268 0.00169751
R22895 GNDA.n2299 GNDA.n2268 0.00169751
R22896 GNDA.n2295 GNDA.n2270 0.00169751
R22897 GNDA.n2344 GNDA.n2271 0.00169751
R22898 GNDA.n2345 GNDA.n2272 0.00169751
R22899 GNDA.n2291 GNDA.n2272 0.00169751
R22900 GNDA.n2287 GNDA.n2274 0.00169751
R22901 GNDA.n2348 GNDA.n2275 0.00169751
R22902 GNDA.n2349 GNDA.n2276 0.00169751
R22903 GNDA.n2283 GNDA.n2276 0.00169751
R22904 GNDA.n2279 GNDA.n2278 0.00169751
R22905 GNDA.n2356 GNDA.n1951 0.00169751
R22906 GNDA.n2151 GNDA.n2107 0.00169751
R22907 GNDA.n2168 GNDA.n2108 0.00169751
R22908 GNDA.n2169 GNDA.n2109 0.00169751
R22909 GNDA.n2153 GNDA.n2109 0.00169751
R22910 GNDA.n2155 GNDA.n2111 0.00169751
R22911 GNDA.n2172 GNDA.n2112 0.00169751
R22912 GNDA.n2173 GNDA.n2113 0.00169751
R22913 GNDA.n2157 GNDA.n2113 0.00169751
R22914 GNDA.n2159 GNDA.n2115 0.00169751
R22915 GNDA.n2176 GNDA.n2116 0.00169751
R22916 GNDA.n2177 GNDA.n2117 0.00169751
R22917 GNDA.n2161 GNDA.n2117 0.00169751
R22918 GNDA.n2223 GNDA.n2119 0.00169751
R22919 GNDA.n2120 GNDA.n361 0.00169751
R22920 GNDA.n2224 GNDA.n2223 0.00169751
R22921 GNDA.n2161 GNDA.n2122 0.00169751
R22922 GNDA.n2159 GNDA.n2124 0.00169751
R22923 GNDA.n2157 GNDA.n2126 0.00169751
R22924 GNDA.n2155 GNDA.n2128 0.00169751
R22925 GNDA.n2153 GNDA.n2130 0.00169751
R22926 GNDA.n2151 GNDA.n2132 0.00169751
R22927 GNDA.n2177 GNDA.n2123 0.00169751
R22928 GNDA.n2176 GNDA.n2124 0.00169751
R22929 GNDA.n2173 GNDA.n2127 0.00169751
R22930 GNDA.n2172 GNDA.n2128 0.00169751
R22931 GNDA.n2169 GNDA.n2131 0.00169751
R22932 GNDA.n2168 GNDA.n2132 0.00169751
R22933 GNDA.n2224 GNDA.n2120 0.00169751
R22934 GNDA.n2280 GNDA.n2279 0.00169751
R22935 GNDA.n2284 GNDA.n2283 0.00169751
R22936 GNDA.n2288 GNDA.n2287 0.00169751
R22937 GNDA.n2292 GNDA.n2291 0.00169751
R22938 GNDA.n2296 GNDA.n2295 0.00169751
R22939 GNDA.n2300 GNDA.n2299 0.00169751
R22940 GNDA.n2304 GNDA.n2303 0.00169751
R22941 GNDA.n2280 GNDA.n1951 0.00169751
R22942 GNDA.n2349 GNDA.n2286 0.00169751
R22943 GNDA.n2348 GNDA.n2288 0.00169751
R22944 GNDA.n2345 GNDA.n2294 0.00169751
R22945 GNDA.n2344 GNDA.n2296 0.00169751
R22946 GNDA.n2341 GNDA.n2302 0.00169751
R22947 GNDA.n2340 GNDA.n2304 0.00169751
R22948 GNDA.n2247 GNDA.n2013 0.00169751
R22949 GNDA.n2245 GNDA.n1996 0.00169751
R22950 GNDA.n2014 GNDA.n1968 0.00169751
R22951 GNDA.n2230 GNDA.n1994 0.00169751
R22952 GNDA.n2231 GNDA.n1993 0.00169751
R22953 GNDA.n2016 GNDA.n1970 0.00169751
R22954 GNDA.n2018 GNDA.n1972 0.00169751
R22955 GNDA.n2234 GNDA.n1990 0.00169751
R22956 GNDA.n2235 GNDA.n1989 0.00169751
R22957 GNDA.n2020 GNDA.n1974 0.00169751
R22958 GNDA.n2022 GNDA.n1976 0.00169751
R22959 GNDA.n2238 GNDA.n1986 0.00169751
R22960 GNDA.n2239 GNDA.n1985 0.00169751
R22961 GNDA.n2024 GNDA.n1978 0.00169751
R22962 GNDA.n2011 GNDA.n1980 0.00169751
R22963 GNDA.n2027 GNDA.n1981 0.00169751
R22964 GNDA.n2239 GNDA.n1978 0.00169751
R22965 GNDA.n2238 GNDA.n1977 0.00169751
R22966 GNDA.n2235 GNDA.n1974 0.00169751
R22967 GNDA.n2234 GNDA.n1973 0.00169751
R22968 GNDA.n2231 GNDA.n1970 0.00169751
R22969 GNDA.n2230 GNDA.n1969 0.00169751
R22970 GNDA.n2056 GNDA.n2013 0.00169751
R22971 GNDA.n2024 GNDA.n1984 0.00169751
R22972 GNDA.n2022 GNDA.n1986 0.00169751
R22973 GNDA.n2020 GNDA.n1988 0.00169751
R22974 GNDA.n2018 GNDA.n1990 0.00169751
R22975 GNDA.n2016 GNDA.n1992 0.00169751
R22976 GNDA.n2014 GNDA.n1994 0.00169751
R22977 GNDA.n2011 GNDA.n1982 0.00169751
R22978 GNDA.n2027 GNDA.n1982 0.00169751
R22979 GNDA.n2056 GNDA.n1996 0.00169751
R22980 GNDA.n2181 GNDA.n2165 0.00166081
R22981 GNDA.n2184 GNDA.n2182 0.00166081
R22982 GNDA.n2187 GNDA.n2185 0.00166081
R22983 GNDA.n2190 GNDA.n2188 0.00166081
R22984 GNDA.n2193 GNDA.n2191 0.00166081
R22985 GNDA.n2196 GNDA.n2194 0.00166081
R22986 GNDA.n2199 GNDA.n2197 0.00166081
R22987 GNDA.n2202 GNDA.n2200 0.00166081
R22988 GNDA.n2205 GNDA.n2203 0.00166081
R22989 GNDA.n2208 GNDA.n2206 0.00166081
R22990 GNDA.n2211 GNDA.n2209 0.00166081
R22991 GNDA.n2214 GNDA.n2212 0.00166081
R22992 GNDA.n2217 GNDA.n2215 0.00166081
R22993 GNDA.n2220 GNDA.n2218 0.00166081
R22994 GNDA.n2225 GNDA.n2221 0.00166081
R22995 GNDA.n2227 GNDA.n2105 0.00166081
R22996 GNDA.n2242 GNDA.n2026 0.00166081
R22997 GNDA.n2059 GNDA.n2028 0.00166081
R22998 GNDA.n2060 GNDA.n2029 0.00166081
R22999 GNDA.n2061 GNDA.n2030 0.00166081
R23000 GNDA.n2062 GNDA.n2031 0.00166081
R23001 GNDA.n2063 GNDA.n2032 0.00166081
R23002 GNDA.n2064 GNDA.n2033 0.00166081
R23003 GNDA.n2065 GNDA.n2034 0.00166081
R23004 GNDA.n2066 GNDA.n2035 0.00166081
R23005 GNDA.n2067 GNDA.n2036 0.00166081
R23006 GNDA.n2068 GNDA.n2037 0.00166081
R23007 GNDA.n2069 GNDA.n2038 0.00166081
R23008 GNDA.n2070 GNDA.n2039 0.00166081
R23009 GNDA.n2071 GNDA.n2040 0.00166081
R23010 GNDA.n2246 GNDA.n2041 0.00166081
R23011 GNDA.n2248 GNDA.n1967 0.00166081
R23012 GNDA.n2353 GNDA.n2321 0.00166081
R23013 GNDA.n2306 GNDA.n2250 0.00166081
R23014 GNDA.n2307 GNDA.n2251 0.00166081
R23015 GNDA.n2308 GNDA.n2252 0.00166081
R23016 GNDA.n2309 GNDA.n2253 0.00166081
R23017 GNDA.n2310 GNDA.n2254 0.00166081
R23018 GNDA.n2311 GNDA.n2255 0.00166081
R23019 GNDA.n2312 GNDA.n2256 0.00166081
R23020 GNDA.n2313 GNDA.n2257 0.00166081
R23021 GNDA.n2314 GNDA.n2258 0.00166081
R23022 GNDA.n2315 GNDA.n2259 0.00166081
R23023 GNDA.n2316 GNDA.n2260 0.00166081
R23024 GNDA.n2317 GNDA.n2261 0.00166081
R23025 GNDA.n2318 GNDA.n2262 0.00166081
R23026 GNDA.n2319 GNDA.n2263 0.00166081
R23027 GNDA.n2355 GNDA.n2264 0.00166081
R23028 GNDA.n2165 GNDA.n2163 0.00166081
R23029 GNDA.n2182 GNDA.n2149 0.00166081
R23030 GNDA.n2185 GNDA.n2148 0.00166081
R23031 GNDA.n2188 GNDA.n2147 0.00166081
R23032 GNDA.n2191 GNDA.n2146 0.00166081
R23033 GNDA.n2194 GNDA.n2145 0.00166081
R23034 GNDA.n2197 GNDA.n2144 0.00166081
R23035 GNDA.n2200 GNDA.n2143 0.00166081
R23036 GNDA.n2203 GNDA.n2142 0.00166081
R23037 GNDA.n2206 GNDA.n2141 0.00166081
R23038 GNDA.n2209 GNDA.n2140 0.00166081
R23039 GNDA.n2212 GNDA.n2139 0.00166081
R23040 GNDA.n2215 GNDA.n2138 0.00166081
R23041 GNDA.n2218 GNDA.n2137 0.00166081
R23042 GNDA.n2221 GNDA.n2136 0.00166081
R23043 GNDA.n2135 GNDA.n2105 0.00166081
R23044 GNDA.n2321 GNDA.n2249 0.00166081
R23045 GNDA.n2306 GNDA.n1966 0.00166081
R23046 GNDA.n2307 GNDA.n1965 0.00166081
R23047 GNDA.n2308 GNDA.n1964 0.00166081
R23048 GNDA.n2309 GNDA.n1963 0.00166081
R23049 GNDA.n2310 GNDA.n1962 0.00166081
R23050 GNDA.n2311 GNDA.n1961 0.00166081
R23051 GNDA.n2312 GNDA.n1960 0.00166081
R23052 GNDA.n2313 GNDA.n1959 0.00166081
R23053 GNDA.n2314 GNDA.n1958 0.00166081
R23054 GNDA.n2315 GNDA.n1957 0.00166081
R23055 GNDA.n2316 GNDA.n1956 0.00166081
R23056 GNDA.n2317 GNDA.n1955 0.00166081
R23057 GNDA.n2318 GNDA.n1954 0.00166081
R23058 GNDA.n2319 GNDA.n1953 0.00166081
R23059 GNDA.n2264 GNDA.n1952 0.00166081
R23060 GNDA.n2243 GNDA.n2242 0.00166081
R23061 GNDA.n2059 GNDA.n2012 0.00166081
R23062 GNDA.n2060 GNDA.n2010 0.00166081
R23063 GNDA.n2061 GNDA.n2009 0.00166081
R23064 GNDA.n2062 GNDA.n2008 0.00166081
R23065 GNDA.n2063 GNDA.n2007 0.00166081
R23066 GNDA.n2064 GNDA.n2006 0.00166081
R23067 GNDA.n2065 GNDA.n2005 0.00166081
R23068 GNDA.n2066 GNDA.n2004 0.00166081
R23069 GNDA.n2067 GNDA.n2003 0.00166081
R23070 GNDA.n2068 GNDA.n2002 0.00166081
R23071 GNDA.n2069 GNDA.n2001 0.00166081
R23072 GNDA.n2070 GNDA.n2000 0.00166081
R23073 GNDA.n2071 GNDA.n1999 0.00166081
R23074 GNDA.n2041 GNDA.n1998 0.00166081
R23075 GNDA.n1997 GNDA.n1967 0.00166081
R23076 GNDA.n2073 GNDA.t591 0.00152174
R23077 GNDA.n2074 GNDA.t421 0.00152174
R23078 GNDA.n2075 GNDA.t283 0.00152174
R23079 GNDA.n2076 GNDA.t673 0.00152174
R23080 GNDA.n2077 GNDA.t265 0.00152174
R23081 GNDA.n2078 GNDA.t655 0.00152174
R23082 GNDA.n2079 GNDA.t500 0.00152174
R23083 GNDA.n2080 GNDA.t637 0.00152174
R23084 GNDA.n2081 GNDA.t735 0.00152174
R23085 GNDA.n2082 GNDA.t308 0.00152174
R23086 GNDA.n2083 GNDA.t442 0.00152174
R23087 GNDA.n2084 GNDA.t310 0.00152174
R23088 GNDA.n2085 GNDA.t713 0.00152174
R23089 GNDA.n2086 GNDA.t560 0.00152174
R23090 GNDA.n2087 GNDA.t693 0.00152174
R23091 GNDA.n2088 GNDA.t539 0.00152174
R23092 GNDA.n2089 GNDA.t369 0.00152174
R23093 GNDA.n2090 GNDA.t518 0.00152174
R23094 GNDA.n2091 GNDA.t348 0.00152174
R23095 GNDA.n2092 GNDA.t207 0.00152174
R23096 GNDA.n2093 GNDA.t328 0.00152174
R23097 GNDA.n2094 GNDA.t189 0.00152174
R23098 GNDA.n2095 GNDA.t580 0.00152174
R23099 GNDA.n2096 GNDA.t408 0.00152174
R23100 GNDA.n2097 GNDA.t561 0.00152174
R23101 GNDA.n2098 GNDA.t409 0.00152174
R23102 GNDA.n2099 GNDA.t270 0.00152174
R23103 GNDA.n2100 GNDA.t388 0.00152174
R23104 GNDA.n2101 GNDA.t252 0.00152174
R23105 GNDA.n2102 GNDA.t643 0.00152174
R23106 GNDA.n2103 GNDA.t232 0.00152174
R23107 GNDA.n2104 GNDA.t622 0.00152174
R23108 two_stage_opamp_dummy_magic_24_0.Vb1.n26 two_stage_opamp_dummy_magic_24_0.Vb1.n25 964.561
R23109 two_stage_opamp_dummy_magic_24_0.Vb1.n36 two_stage_opamp_dummy_magic_24_0.Vb1.n35 630.693
R23110 two_stage_opamp_dummy_magic_24_0.Vb1.n17 two_stage_opamp_dummy_magic_24_0.Vb1.t237 449.868
R23111 two_stage_opamp_dummy_magic_24_0.Vb1.n8 two_stage_opamp_dummy_magic_24_0.Vb1.t222 449.868
R23112 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.t220 449.868
R23113 two_stage_opamp_dummy_magic_24_0.Vb1.n35 two_stage_opamp_dummy_magic_24_0.Vb1.t231 273.134
R23114 two_stage_opamp_dummy_magic_24_0.Vb1.n26 two_stage_opamp_dummy_magic_24_0.Vb1.t238 273.134
R23115 two_stage_opamp_dummy_magic_24_0.Vb1.n25 two_stage_opamp_dummy_magic_24_0.Vb1.t236 273.134
R23116 two_stage_opamp_dummy_magic_24_0.Vb1.n24 two_stage_opamp_dummy_magic_24_0.Vb1.t247 273.134
R23117 two_stage_opamp_dummy_magic_24_0.Vb1.n23 two_stage_opamp_dummy_magic_24_0.Vb1.t235 273.134
R23118 two_stage_opamp_dummy_magic_24_0.Vb1.n22 two_stage_opamp_dummy_magic_24_0.Vb1.t245 273.134
R23119 two_stage_opamp_dummy_magic_24_0.Vb1.n21 two_stage_opamp_dummy_magic_24_0.Vb1.t232 273.134
R23120 two_stage_opamp_dummy_magic_24_0.Vb1.n20 two_stage_opamp_dummy_magic_24_0.Vb1.t246 273.134
R23121 two_stage_opamp_dummy_magic_24_0.Vb1.n19 two_stage_opamp_dummy_magic_24_0.Vb1.t233 273.134
R23122 two_stage_opamp_dummy_magic_24_0.Vb1.n18 two_stage_opamp_dummy_magic_24_0.Vb1.t244 273.134
R23123 two_stage_opamp_dummy_magic_24_0.Vb1.n17 two_stage_opamp_dummy_magic_24_0.Vb1.t230 273.134
R23124 two_stage_opamp_dummy_magic_24_0.Vb1.n34 two_stage_opamp_dummy_magic_24_0.Vb1.t243 273.134
R23125 two_stage_opamp_dummy_magic_24_0.Vb1.n33 two_stage_opamp_dummy_magic_24_0.Vb1.t229 273.134
R23126 two_stage_opamp_dummy_magic_24_0.Vb1.n32 two_stage_opamp_dummy_magic_24_0.Vb1.t242 273.134
R23127 two_stage_opamp_dummy_magic_24_0.Vb1.n31 two_stage_opamp_dummy_magic_24_0.Vb1.t228 273.134
R23128 two_stage_opamp_dummy_magic_24_0.Vb1.n30 two_stage_opamp_dummy_magic_24_0.Vb1.t239 273.134
R23129 two_stage_opamp_dummy_magic_24_0.Vb1.n29 two_stage_opamp_dummy_magic_24_0.Vb1.t234 273.134
R23130 two_stage_opamp_dummy_magic_24_0.Vb1.n28 two_stage_opamp_dummy_magic_24_0.Vb1.t240 273.134
R23131 two_stage_opamp_dummy_magic_24_0.Vb1.n27 two_stage_opamp_dummy_magic_24_0.Vb1.t248 273.134
R23132 two_stage_opamp_dummy_magic_24_0.Vb1.n8 two_stage_opamp_dummy_magic_24_0.Vb1.t226 273.134
R23133 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.t224 273.134
R23134 two_stage_opamp_dummy_magic_24_0.Vb1.n2 two_stage_opamp_dummy_magic_24_0.Vb1.n0 217.208
R23135 two_stage_opamp_dummy_magic_24_0.Vb1.n18 two_stage_opamp_dummy_magic_24_0.Vb1.n17 176.733
R23136 two_stage_opamp_dummy_magic_24_0.Vb1.n19 two_stage_opamp_dummy_magic_24_0.Vb1.n18 176.733
R23137 two_stage_opamp_dummy_magic_24_0.Vb1.n20 two_stage_opamp_dummy_magic_24_0.Vb1.n19 176.733
R23138 two_stage_opamp_dummy_magic_24_0.Vb1.n21 two_stage_opamp_dummy_magic_24_0.Vb1.n20 176.733
R23139 two_stage_opamp_dummy_magic_24_0.Vb1.n22 two_stage_opamp_dummy_magic_24_0.Vb1.n21 176.733
R23140 two_stage_opamp_dummy_magic_24_0.Vb1.n23 two_stage_opamp_dummy_magic_24_0.Vb1.n22 176.733
R23141 two_stage_opamp_dummy_magic_24_0.Vb1.n24 two_stage_opamp_dummy_magic_24_0.Vb1.n23 176.733
R23142 two_stage_opamp_dummy_magic_24_0.Vb1.n25 two_stage_opamp_dummy_magic_24_0.Vb1.n24 176.733
R23143 two_stage_opamp_dummy_magic_24_0.Vb1.n27 two_stage_opamp_dummy_magic_24_0.Vb1.n26 176.733
R23144 two_stage_opamp_dummy_magic_24_0.Vb1.n28 two_stage_opamp_dummy_magic_24_0.Vb1.n27 176.733
R23145 two_stage_opamp_dummy_magic_24_0.Vb1.n29 two_stage_opamp_dummy_magic_24_0.Vb1.n28 176.733
R23146 two_stage_opamp_dummy_magic_24_0.Vb1.n30 two_stage_opamp_dummy_magic_24_0.Vb1.n29 176.733
R23147 two_stage_opamp_dummy_magic_24_0.Vb1.n31 two_stage_opamp_dummy_magic_24_0.Vb1.n30 176.733
R23148 two_stage_opamp_dummy_magic_24_0.Vb1.n32 two_stage_opamp_dummy_magic_24_0.Vb1.n31 176.733
R23149 two_stage_opamp_dummy_magic_24_0.Vb1.n33 two_stage_opamp_dummy_magic_24_0.Vb1.n32 176.733
R23150 two_stage_opamp_dummy_magic_24_0.Vb1.n34 two_stage_opamp_dummy_magic_24_0.Vb1.n33 176.733
R23151 two_stage_opamp_dummy_magic_24_0.Vb1.n35 two_stage_opamp_dummy_magic_24_0.Vb1.n34 176.733
R23152 two_stage_opamp_dummy_magic_24_0.Vb1.n4 two_stage_opamp_dummy_magic_24_0.Vb1.t241 167.769
R23153 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.n9 161.3
R23154 bgr_11_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_24_0.Vb1.n36 58.6984
R23155 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.n5 49.3505
R23156 two_stage_opamp_dummy_magic_24_0.Vb1.n12 two_stage_opamp_dummy_magic_24_0.Vb1.n11 49.3505
R23157 two_stage_opamp_dummy_magic_24_0.Vb1.n15 two_stage_opamp_dummy_magic_24_0.Vb1.n14 49.3505
R23158 two_stage_opamp_dummy_magic_24_0.Vb1.n9 two_stage_opamp_dummy_magic_24_0.Vb1.n8 45.5227
R23159 two_stage_opamp_dummy_magic_24_0.Vb1.n9 two_stage_opamp_dummy_magic_24_0.Vb1.n7 45.5227
R23160 two_stage_opamp_dummy_magic_24_0.Vb1.n36 two_stage_opamp_dummy_magic_24_0.Vb1.n16 19.9172
R23161 two_stage_opamp_dummy_magic_24_0.Vb1.n0 two_stage_opamp_dummy_magic_24_0.Vb1.t1 19.7005
R23162 two_stage_opamp_dummy_magic_24_0.Vb1.n0 two_stage_opamp_dummy_magic_24_0.Vb1.t0 19.7005
R23163 two_stage_opamp_dummy_magic_24_0.Vb1.n5 two_stage_opamp_dummy_magic_24_0.Vb1.t219 16.0005
R23164 two_stage_opamp_dummy_magic_24_0.Vb1.n5 two_stage_opamp_dummy_magic_24_0.Vb1.t221 16.0005
R23165 two_stage_opamp_dummy_magic_24_0.Vb1.n11 two_stage_opamp_dummy_magic_24_0.Vb1.t225 16.0005
R23166 two_stage_opamp_dummy_magic_24_0.Vb1.n11 two_stage_opamp_dummy_magic_24_0.Vb1.t227 16.0005
R23167 two_stage_opamp_dummy_magic_24_0.Vb1.n14 two_stage_opamp_dummy_magic_24_0.Vb1.t223 16.0005
R23168 two_stage_opamp_dummy_magic_24_0.Vb1.n14 two_stage_opamp_dummy_magic_24_0.Vb1.t218 16.0005
R23169 two_stage_opamp_dummy_magic_24_0.Vb1.n2 two_stage_opamp_dummy_magic_24_0.Vb1.t212 11.2142
R23170 two_stage_opamp_dummy_magic_24_0.Vb1.n15 two_stage_opamp_dummy_magic_24_0.Vb1.n13 5.6255
R23171 two_stage_opamp_dummy_magic_24_0.Vb1.n13 two_stage_opamp_dummy_magic_24_0.Vb1.n6 5.6255
R23172 two_stage_opamp_dummy_magic_24_0.Vb1.n13 two_stage_opamp_dummy_magic_24_0.Vb1.n12 5.063
R23173 two_stage_opamp_dummy_magic_24_0.Vb1.n16 two_stage_opamp_dummy_magic_24_0.Vb1.n15 4.938
R23174 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.n4 4.938
R23175 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.n3 4.5005
R23176 bgr_11_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_24_0.Vb1.n2 1.03175
R23177 two_stage_opamp_dummy_magic_24_0.Vb1.n4 two_stage_opamp_dummy_magic_24_0.Vb1.n3 0.563
R23178 two_stage_opamp_dummy_magic_24_0.Vb1.n16 two_stage_opamp_dummy_magic_24_0.Vb1.n3 0.563
R23179 two_stage_opamp_dummy_magic_24_0.Vb1.n12 two_stage_opamp_dummy_magic_24_0.Vb1.n10 0.438
R23180 two_stage_opamp_dummy_magic_24_0.Vb1.t217 two_stage_opamp_dummy_magic_24_0.Vb1.n1 0.334609
R23181 two_stage_opamp_dummy_magic_24_0.Vb1.t215 two_stage_opamp_dummy_magic_24_0.Vb1.t156 0.1603
R23182 two_stage_opamp_dummy_magic_24_0.Vb1.t178 two_stage_opamp_dummy_magic_24_0.Vb1.t215 0.1603
R23183 two_stage_opamp_dummy_magic_24_0.Vb1.t18 two_stage_opamp_dummy_magic_24_0.Vb1.t178 0.1603
R23184 two_stage_opamp_dummy_magic_24_0.Vb1.t151 two_stage_opamp_dummy_magic_24_0.Vb1.t93 0.1603
R23185 two_stage_opamp_dummy_magic_24_0.Vb1.t117 two_stage_opamp_dummy_magic_24_0.Vb1.t151 0.1603
R23186 two_stage_opamp_dummy_magic_24_0.Vb1.t170 two_stage_opamp_dummy_magic_24_0.Vb1.t117 0.1603
R23187 two_stage_opamp_dummy_magic_24_0.Vb1.t211 two_stage_opamp_dummy_magic_24_0.Vb1.t155 0.1603
R23188 two_stage_opamp_dummy_magic_24_0.Vb1.t53 two_stage_opamp_dummy_magic_24_0.Vb1.t211 0.1603
R23189 two_stage_opamp_dummy_magic_24_0.Vb1.t20 two_stage_opamp_dummy_magic_24_0.Vb1.t53 0.1603
R23190 two_stage_opamp_dummy_magic_24_0.Vb1.t61 two_stage_opamp_dummy_magic_24_0.Vb1.t2 0.1603
R23191 two_stage_opamp_dummy_magic_24_0.Vb1.t23 two_stage_opamp_dummy_magic_24_0.Vb1.t61 0.1603
R23192 two_stage_opamp_dummy_magic_24_0.Vb1.t82 two_stage_opamp_dummy_magic_24_0.Vb1.t23 0.1603
R23193 two_stage_opamp_dummy_magic_24_0.Vb1.t120 two_stage_opamp_dummy_magic_24_0.Vb1.t63 0.1603
R23194 two_stage_opamp_dummy_magic_24_0.Vb1.t176 two_stage_opamp_dummy_magic_24_0.Vb1.t120 0.1603
R23195 two_stage_opamp_dummy_magic_24_0.Vb1.t144 two_stage_opamp_dummy_magic_24_0.Vb1.t176 0.1603
R23196 two_stage_opamp_dummy_magic_24_0.Vb1.t122 two_stage_opamp_dummy_magic_24_0.Vb1.t64 0.1603
R23197 two_stage_opamp_dummy_magic_24_0.Vb1.t85 two_stage_opamp_dummy_magic_24_0.Vb1.t122 0.1603
R23198 two_stage_opamp_dummy_magic_24_0.Vb1.t143 two_stage_opamp_dummy_magic_24_0.Vb1.t85 0.1603
R23199 two_stage_opamp_dummy_magic_24_0.Vb1.t180 two_stage_opamp_dummy_magic_24_0.Vb1.t123 0.1603
R23200 two_stage_opamp_dummy_magic_24_0.Vb1.t22 two_stage_opamp_dummy_magic_24_0.Vb1.t180 0.1603
R23201 two_stage_opamp_dummy_magic_24_0.Vb1.t206 two_stage_opamp_dummy_magic_24_0.Vb1.t22 0.1603
R23202 two_stage_opamp_dummy_magic_24_0.Vb1.t70 two_stage_opamp_dummy_magic_24_0.Vb1.t12 0.1603
R23203 two_stage_opamp_dummy_magic_24_0.Vb1.t31 two_stage_opamp_dummy_magic_24_0.Vb1.t70 0.1603
R23204 two_stage_opamp_dummy_magic_24_0.Vb1.t87 two_stage_opamp_dummy_magic_24_0.Vb1.t31 0.1603
R23205 two_stage_opamp_dummy_magic_24_0.Vb1.t127 two_stage_opamp_dummy_magic_24_0.Vb1.t72 0.1603
R23206 two_stage_opamp_dummy_magic_24_0.Vb1.t185 two_stage_opamp_dummy_magic_24_0.Vb1.t127 0.1603
R23207 two_stage_opamp_dummy_magic_24_0.Vb1.t149 two_stage_opamp_dummy_magic_24_0.Vb1.t185 0.1603
R23208 two_stage_opamp_dummy_magic_24_0.Vb1.t131 two_stage_opamp_dummy_magic_24_0.Vb1.t74 0.1603
R23209 two_stage_opamp_dummy_magic_24_0.Vb1.t96 two_stage_opamp_dummy_magic_24_0.Vb1.t131 0.1603
R23210 two_stage_opamp_dummy_magic_24_0.Vb1.t148 two_stage_opamp_dummy_magic_24_0.Vb1.t96 0.1603
R23211 two_stage_opamp_dummy_magic_24_0.Vb1.t187 two_stage_opamp_dummy_magic_24_0.Vb1.t132 0.1603
R23212 two_stage_opamp_dummy_magic_24_0.Vb1.t30 two_stage_opamp_dummy_magic_24_0.Vb1.t187 0.1603
R23213 two_stage_opamp_dummy_magic_24_0.Vb1.t213 two_stage_opamp_dummy_magic_24_0.Vb1.t30 0.1603
R23214 two_stage_opamp_dummy_magic_24_0.Vb1.t190 two_stage_opamp_dummy_magic_24_0.Vb1.t134 0.1603
R23215 two_stage_opamp_dummy_magic_24_0.Vb1.t158 two_stage_opamp_dummy_magic_24_0.Vb1.t190 0.1603
R23216 two_stage_opamp_dummy_magic_24_0.Vb1.t209 two_stage_opamp_dummy_magic_24_0.Vb1.t158 0.1603
R23217 two_stage_opamp_dummy_magic_24_0.Vb1.t32 two_stage_opamp_dummy_magic_24_0.Vb1.t191 0.1603
R23218 two_stage_opamp_dummy_magic_24_0.Vb1.t92 two_stage_opamp_dummy_magic_24_0.Vb1.t32 0.1603
R23219 two_stage_opamp_dummy_magic_24_0.Vb1.t60 two_stage_opamp_dummy_magic_24_0.Vb1.t92 0.1603
R23220 two_stage_opamp_dummy_magic_24_0.Vb1.t137 two_stage_opamp_dummy_magic_24_0.Vb1.t78 0.1603
R23221 two_stage_opamp_dummy_magic_24_0.Vb1.t102 two_stage_opamp_dummy_magic_24_0.Vb1.t137 0.1603
R23222 two_stage_opamp_dummy_magic_24_0.Vb1.t159 two_stage_opamp_dummy_magic_24_0.Vb1.t102 0.1603
R23223 two_stage_opamp_dummy_magic_24_0.Vb1.t196 two_stage_opamp_dummy_magic_24_0.Vb1.t139 0.1603
R23224 two_stage_opamp_dummy_magic_24_0.Vb1.t40 two_stage_opamp_dummy_magic_24_0.Vb1.t196 0.1603
R23225 two_stage_opamp_dummy_magic_24_0.Vb1.t8 two_stage_opamp_dummy_magic_24_0.Vb1.t40 0.1603
R23226 two_stage_opamp_dummy_magic_24_0.Vb1.t199 two_stage_opamp_dummy_magic_24_0.Vb1.t141 0.1603
R23227 two_stage_opamp_dummy_magic_24_0.Vb1.t165 two_stage_opamp_dummy_magic_24_0.Vb1.t199 0.1603
R23228 two_stage_opamp_dummy_magic_24_0.Vb1.t7 two_stage_opamp_dummy_magic_24_0.Vb1.t165 0.1603
R23229 two_stage_opamp_dummy_magic_24_0.Vb1.t44 two_stage_opamp_dummy_magic_24_0.Vb1.t201 0.1603
R23230 two_stage_opamp_dummy_magic_24_0.Vb1.t101 two_stage_opamp_dummy_magic_24_0.Vb1.t44 0.1603
R23231 two_stage_opamp_dummy_magic_24_0.Vb1.t68 two_stage_opamp_dummy_magic_24_0.Vb1.t101 0.1603
R23232 two_stage_opamp_dummy_magic_24_0.Vb1.t36 two_stage_opamp_dummy_magic_24_0.Vb1.t193 0.1603
R23233 two_stage_opamp_dummy_magic_24_0.Vb1.t4 two_stage_opamp_dummy_magic_24_0.Vb1.t36 0.1603
R23234 two_stage_opamp_dummy_magic_24_0.Vb1.t57 two_stage_opamp_dummy_magic_24_0.Vb1.t4 0.1603
R23235 two_stage_opamp_dummy_magic_24_0.Vb1.t95 two_stage_opamp_dummy_magic_24_0.Vb1.t38 0.1603
R23236 two_stage_opamp_dummy_magic_24_0.Vb1.t154 two_stage_opamp_dummy_magic_24_0.Vb1.t95 0.1603
R23237 two_stage_opamp_dummy_magic_24_0.Vb1.t119 two_stage_opamp_dummy_magic_24_0.Vb1.t154 0.1603
R23238 two_stage_opamp_dummy_magic_24_0.Vb1.t198 two_stage_opamp_dummy_magic_24_0.Vb1.t140 0.1603
R23239 two_stage_opamp_dummy_magic_24_0.Vb1.t164 two_stage_opamp_dummy_magic_24_0.Vb1.t198 0.1603
R23240 two_stage_opamp_dummy_magic_24_0.Vb1.t6 two_stage_opamp_dummy_magic_24_0.Vb1.t164 0.1603
R23241 two_stage_opamp_dummy_magic_24_0.Vb1.t42 two_stage_opamp_dummy_magic_24_0.Vb1.t200 0.1603
R23242 two_stage_opamp_dummy_magic_24_0.Vb1.t99 two_stage_opamp_dummy_magic_24_0.Vb1.t42 0.1603
R23243 two_stage_opamp_dummy_magic_24_0.Vb1.t67 two_stage_opamp_dummy_magic_24_0.Vb1.t99 0.1603
R23244 two_stage_opamp_dummy_magic_24_0.Vb1.t46 two_stage_opamp_dummy_magic_24_0.Vb1.t202 0.1603
R23245 two_stage_opamp_dummy_magic_24_0.Vb1.t11 two_stage_opamp_dummy_magic_24_0.Vb1.t46 0.1603
R23246 two_stage_opamp_dummy_magic_24_0.Vb1.t66 two_stage_opamp_dummy_magic_24_0.Vb1.t11 0.1603
R23247 two_stage_opamp_dummy_magic_24_0.Vb1.t103 two_stage_opamp_dummy_magic_24_0.Vb1.t47 0.1603
R23248 two_stage_opamp_dummy_magic_24_0.Vb1.t163 two_stage_opamp_dummy_magic_24_0.Vb1.t103 0.1603
R23249 two_stage_opamp_dummy_magic_24_0.Vb1.t128 two_stage_opamp_dummy_magic_24_0.Vb1.t163 0.1603
R23250 two_stage_opamp_dummy_magic_24_0.Vb1.t105 two_stage_opamp_dummy_magic_24_0.Vb1.t48 0.1603
R23251 two_stage_opamp_dummy_magic_24_0.Vb1.t73 two_stage_opamp_dummy_magic_24_0.Vb1.t105 0.1603
R23252 two_stage_opamp_dummy_magic_24_0.Vb1.t126 two_stage_opamp_dummy_magic_24_0.Vb1.t73 0.1603
R23253 two_stage_opamp_dummy_magic_24_0.Vb1.t166 two_stage_opamp_dummy_magic_24_0.Vb1.t106 0.1603
R23254 two_stage_opamp_dummy_magic_24_0.Vb1.t10 two_stage_opamp_dummy_magic_24_0.Vb1.t166 0.1603
R23255 two_stage_opamp_dummy_magic_24_0.Vb1.t188 two_stage_opamp_dummy_magic_24_0.Vb1.t10 0.1603
R23256 two_stage_opamp_dummy_magic_24_0.Vb1.t167 two_stage_opamp_dummy_magic_24_0.Vb1.t107 0.1603
R23257 two_stage_opamp_dummy_magic_24_0.Vb1.t133 two_stage_opamp_dummy_magic_24_0.Vb1.t167 0.1603
R23258 two_stage_opamp_dummy_magic_24_0.Vb1.t186 two_stage_opamp_dummy_magic_24_0.Vb1.t133 0.1603
R23259 two_stage_opamp_dummy_magic_24_0.Vb1.t13 two_stage_opamp_dummy_magic_24_0.Vb1.t168 0.1603
R23260 two_stage_opamp_dummy_magic_24_0.Vb1.t71 two_stage_opamp_dummy_magic_24_0.Vb1.t13 0.1603
R23261 two_stage_opamp_dummy_magic_24_0.Vb1.t33 two_stage_opamp_dummy_magic_24_0.Vb1.t71 0.1603
R23262 two_stage_opamp_dummy_magic_24_0.Vb1.t111 two_stage_opamp_dummy_magic_24_0.Vb1.t52 0.1603
R23263 two_stage_opamp_dummy_magic_24_0.Vb1.t79 two_stage_opamp_dummy_magic_24_0.Vb1.t111 0.1603
R23264 two_stage_opamp_dummy_magic_24_0.Vb1.t135 two_stage_opamp_dummy_magic_24_0.Vb1.t79 0.1603
R23265 two_stage_opamp_dummy_magic_24_0.Vb1.t169 two_stage_opamp_dummy_magic_24_0.Vb1.t113 0.1603
R23266 two_stage_opamp_dummy_magic_24_0.Vb1.t15 two_stage_opamp_dummy_magic_24_0.Vb1.t169 0.1603
R23267 two_stage_opamp_dummy_magic_24_0.Vb1.t195 two_stage_opamp_dummy_magic_24_0.Vb1.t15 0.1603
R23268 two_stage_opamp_dummy_magic_24_0.Vb1.t172 two_stage_opamp_dummy_magic_24_0.Vb1.t114 0.1603
R23269 two_stage_opamp_dummy_magic_24_0.Vb1.t142 two_stage_opamp_dummy_magic_24_0.Vb1.t172 0.1603
R23270 two_stage_opamp_dummy_magic_24_0.Vb1.t194 two_stage_opamp_dummy_magic_24_0.Vb1.t142 0.1603
R23271 two_stage_opamp_dummy_magic_24_0.Vb1.t17 two_stage_opamp_dummy_magic_24_0.Vb1.t173 0.1603
R23272 two_stage_opamp_dummy_magic_24_0.Vb1.t77 two_stage_opamp_dummy_magic_24_0.Vb1.t17 0.1603
R23273 two_stage_opamp_dummy_magic_24_0.Vb1.t43 two_stage_opamp_dummy_magic_24_0.Vb1.t77 0.1603
R23274 two_stage_opamp_dummy_magic_24_0.Vb1.t19 two_stage_opamp_dummy_magic_24_0.Vb1.t175 0.1603
R23275 two_stage_opamp_dummy_magic_24_0.Vb1.t203 two_stage_opamp_dummy_magic_24_0.Vb1.t19 0.1603
R23276 two_stage_opamp_dummy_magic_24_0.Vb1.t41 two_stage_opamp_dummy_magic_24_0.Vb1.t203 0.1603
R23277 two_stage_opamp_dummy_magic_24_0.Vb1.t80 two_stage_opamp_dummy_magic_24_0.Vb1.t21 0.1603
R23278 two_stage_opamp_dummy_magic_24_0.Vb1.t138 two_stage_opamp_dummy_magic_24_0.Vb1.t80 0.1603
R23279 two_stage_opamp_dummy_magic_24_0.Vb1.t104 two_stage_opamp_dummy_magic_24_0.Vb1.t138 0.1603
R23280 two_stage_opamp_dummy_magic_24_0.Vb1.t182 two_stage_opamp_dummy_magic_24_0.Vb1.t124 0.1603
R23281 two_stage_opamp_dummy_magic_24_0.Vb1.t146 two_stage_opamp_dummy_magic_24_0.Vb1.t182 0.1603
R23282 two_stage_opamp_dummy_magic_24_0.Vb1.t204 two_stage_opamp_dummy_magic_24_0.Vb1.t146 0.1603
R23283 two_stage_opamp_dummy_magic_24_0.Vb1.t24 two_stage_opamp_dummy_magic_24_0.Vb1.t183 0.1603
R23284 two_stage_opamp_dummy_magic_24_0.Vb1.t84 two_stage_opamp_dummy_magic_24_0.Vb1.t24 0.1603
R23285 two_stage_opamp_dummy_magic_24_0.Vb1.t50 two_stage_opamp_dummy_magic_24_0.Vb1.t84 0.1603
R23286 two_stage_opamp_dummy_magic_24_0.Vb1.t26 two_stage_opamp_dummy_magic_24_0.Vb1.t184 0.1603
R23287 two_stage_opamp_dummy_magic_24_0.Vb1.t208 two_stage_opamp_dummy_magic_24_0.Vb1.t26 0.1603
R23288 two_stage_opamp_dummy_magic_24_0.Vb1.t49 two_stage_opamp_dummy_magic_24_0.Vb1.t208 0.1603
R23289 two_stage_opamp_dummy_magic_24_0.Vb1.t86 two_stage_opamp_dummy_magic_24_0.Vb1.t27 0.1603
R23290 two_stage_opamp_dummy_magic_24_0.Vb1.t145 two_stage_opamp_dummy_magic_24_0.Vb1.t86 0.1603
R23291 two_stage_opamp_dummy_magic_24_0.Vb1.t109 two_stage_opamp_dummy_magic_24_0.Vb1.t145 0.1603
R23292 two_stage_opamp_dummy_magic_24_0.Vb1.t89 two_stage_opamp_dummy_magic_24_0.Vb1.t29 0.1603
R23293 two_stage_opamp_dummy_magic_24_0.Vb1.t54 two_stage_opamp_dummy_magic_24_0.Vb1.t89 0.1603
R23294 two_stage_opamp_dummy_magic_24_0.Vb1.t108 two_stage_opamp_dummy_magic_24_0.Vb1.t54 0.1603
R23295 two_stage_opamp_dummy_magic_24_0.Vb1.t147 two_stage_opamp_dummy_magic_24_0.Vb1.t90 0.1603
R23296 two_stage_opamp_dummy_magic_24_0.Vb1.t207 two_stage_opamp_dummy_magic_24_0.Vb1.t147 0.1603
R23297 two_stage_opamp_dummy_magic_24_0.Vb1.t171 two_stage_opamp_dummy_magic_24_0.Vb1.t207 0.1603
R23298 two_stage_opamp_dummy_magic_24_0.Vb1.t35 two_stage_opamp_dummy_magic_24_0.Vb1.t192 0.1603
R23299 two_stage_opamp_dummy_magic_24_0.Vb1.t3 two_stage_opamp_dummy_magic_24_0.Vb1.t35 0.1603
R23300 two_stage_opamp_dummy_magic_24_0.Vb1.t56 two_stage_opamp_dummy_magic_24_0.Vb1.t3 0.1603
R23301 two_stage_opamp_dummy_magic_24_0.Vb1.t94 two_stage_opamp_dummy_magic_24_0.Vb1.t37 0.1603
R23302 two_stage_opamp_dummy_magic_24_0.Vb1.t153 two_stage_opamp_dummy_magic_24_0.Vb1.t94 0.1603
R23303 two_stage_opamp_dummy_magic_24_0.Vb1.t118 two_stage_opamp_dummy_magic_24_0.Vb1.t153 0.1603
R23304 two_stage_opamp_dummy_magic_24_0.Vb1.t97 two_stage_opamp_dummy_magic_24_0.Vb1.t39 0.1603
R23305 two_stage_opamp_dummy_magic_24_0.Vb1.t65 two_stage_opamp_dummy_magic_24_0.Vb1.t97 0.1603
R23306 two_stage_opamp_dummy_magic_24_0.Vb1.t116 two_stage_opamp_dummy_magic_24_0.Vb1.t65 0.1603
R23307 two_stage_opamp_dummy_magic_24_0.Vb1.t157 two_stage_opamp_dummy_magic_24_0.Vb1.t98 0.1603
R23308 two_stage_opamp_dummy_magic_24_0.Vb1.t216 two_stage_opamp_dummy_magic_24_0.Vb1.t157 0.1603
R23309 two_stage_opamp_dummy_magic_24_0.Vb1.t179 two_stage_opamp_dummy_magic_24_0.Vb1.t216 0.1603
R23310 two_stage_opamp_dummy_magic_24_0.Vb1.t160 two_stage_opamp_dummy_magic_24_0.Vb1.t100 0.1603
R23311 two_stage_opamp_dummy_magic_24_0.Vb1.t125 two_stage_opamp_dummy_magic_24_0.Vb1.t160 0.1603
R23312 two_stage_opamp_dummy_magic_24_0.Vb1.t177 two_stage_opamp_dummy_magic_24_0.Vb1.t125 0.1603
R23313 two_stage_opamp_dummy_magic_24_0.Vb1.t5 two_stage_opamp_dummy_magic_24_0.Vb1.t161 0.1603
R23314 two_stage_opamp_dummy_magic_24_0.Vb1.t62 two_stage_opamp_dummy_magic_24_0.Vb1.t5 0.1603
R23315 two_stage_opamp_dummy_magic_24_0.Vb1.t25 two_stage_opamp_dummy_magic_24_0.Vb1.t62 0.1603
R23316 two_stage_opamp_dummy_magic_24_0.Vb1.t210 two_stage_opamp_dummy_magic_24_0.Vb1.t152 0.1603
R23317 two_stage_opamp_dummy_magic_24_0.Vb1.t174 two_stage_opamp_dummy_magic_24_0.Vb1.t210 0.1603
R23318 two_stage_opamp_dummy_magic_24_0.Vb1.t16 two_stage_opamp_dummy_magic_24_0.Vb1.t174 0.1603
R23319 two_stage_opamp_dummy_magic_24_0.Vb1.t212 two_stage_opamp_dummy_magic_24_0.Vb1.t55 0.1603
R23320 two_stage_opamp_dummy_magic_24_0.Vb1.t55 two_stage_opamp_dummy_magic_24_0.Vb1.t112 0.1603
R23321 two_stage_opamp_dummy_magic_24_0.Vb1.t112 two_stage_opamp_dummy_magic_24_0.Vb1.t81 0.1603
R23322 two_stage_opamp_dummy_magic_24_0.Vb1.t83 two_stage_opamp_dummy_magic_24_0.Vb1.t115 0.1603
R23323 two_stage_opamp_dummy_magic_24_0.Vb1.t115 two_stage_opamp_dummy_magic_24_0.Vb1.t58 0.1603
R23324 two_stage_opamp_dummy_magic_24_0.Vb1.t58 two_stage_opamp_dummy_magic_24_0.Vb1.t217 0.1603
R23325 two_stage_opamp_dummy_magic_24_0.Vb1.t91 two_stage_opamp_dummy_magic_24_0.Vb1.t28 0.159278
R23326 two_stage_opamp_dummy_magic_24_0.Vb1.t88 two_stage_opamp_dummy_magic_24_0.Vb1.t34 0.159278
R23327 two_stage_opamp_dummy_magic_24_0.Vb1.t34 two_stage_opamp_dummy_magic_24_0.Vb1.t189 0.159278
R23328 two_stage_opamp_dummy_magic_24_0.Vb1.t189 two_stage_opamp_dummy_magic_24_0.Vb1.t129 0.159278
R23329 two_stage_opamp_dummy_magic_24_0.Vb1.t129 two_stage_opamp_dummy_magic_24_0.Vb1.t181 0.159278
R23330 two_stage_opamp_dummy_magic_24_0.Vb1.t181 two_stage_opamp_dummy_magic_24_0.Vb1.t121 0.159278
R23331 two_stage_opamp_dummy_magic_24_0.Vb1.t121 two_stage_opamp_dummy_magic_24_0.Vb1.t59 0.159278
R23332 two_stage_opamp_dummy_magic_24_0.Vb1.t59 two_stage_opamp_dummy_magic_24_0.Vb1.t110 0.159278
R23333 two_stage_opamp_dummy_magic_24_0.Vb1.t110 two_stage_opamp_dummy_magic_24_0.Vb1.t51 0.159278
R23334 two_stage_opamp_dummy_magic_24_0.Vb1.t51 two_stage_opamp_dummy_magic_24_0.Vb1.t205 0.159278
R23335 two_stage_opamp_dummy_magic_24_0.Vb1.t205 two_stage_opamp_dummy_magic_24_0.Vb1.t45 0.159278
R23336 two_stage_opamp_dummy_magic_24_0.Vb1.t45 two_stage_opamp_dummy_magic_24_0.Vb1.t197 0.159278
R23337 two_stage_opamp_dummy_magic_24_0.Vb1.t197 two_stage_opamp_dummy_magic_24_0.Vb1.t136 0.159278
R23338 two_stage_opamp_dummy_magic_24_0.Vb1.t136 two_stage_opamp_dummy_magic_24_0.Vb1.t75 0.159278
R23339 two_stage_opamp_dummy_magic_24_0.Vb1.t75 two_stage_opamp_dummy_magic_24_0.Vb1.t130 0.159278
R23340 two_stage_opamp_dummy_magic_24_0.Vb1.t130 two_stage_opamp_dummy_magic_24_0.Vb1.t76 0.159278
R23341 two_stage_opamp_dummy_magic_24_0.Vb1.t76 two_stage_opamp_dummy_magic_24_0.Vb1.t14 0.159278
R23342 two_stage_opamp_dummy_magic_24_0.Vb1.t14 two_stage_opamp_dummy_magic_24_0.Vb1.t69 0.159278
R23343 two_stage_opamp_dummy_magic_24_0.Vb1.t69 two_stage_opamp_dummy_magic_24_0.Vb1.t9 0.159278
R23344 two_stage_opamp_dummy_magic_24_0.Vb1.t9 two_stage_opamp_dummy_magic_24_0.Vb1.t162 0.159278
R23345 two_stage_opamp_dummy_magic_24_0.Vb1.t162 two_stage_opamp_dummy_magic_24_0.Vb1.t214 0.159278
R23346 two_stage_opamp_dummy_magic_24_0.Vb1.t214 two_stage_opamp_dummy_magic_24_0.Vb1.t150 0.159278
R23347 two_stage_opamp_dummy_magic_24_0.Vb1.t150 two_stage_opamp_dummy_magic_24_0.Vb1.t91 0.159278
R23348 two_stage_opamp_dummy_magic_24_0.Vb1.t91 two_stage_opamp_dummy_magic_24_0.Vb1.t18 0.137822
R23349 two_stage_opamp_dummy_magic_24_0.Vb1.t150 two_stage_opamp_dummy_magic_24_0.Vb1.t144 0.137822
R23350 two_stage_opamp_dummy_magic_24_0.Vb1.t214 two_stage_opamp_dummy_magic_24_0.Vb1.t206 0.137822
R23351 two_stage_opamp_dummy_magic_24_0.Vb1.t162 two_stage_opamp_dummy_magic_24_0.Vb1.t149 0.137822
R23352 two_stage_opamp_dummy_magic_24_0.Vb1.t9 two_stage_opamp_dummy_magic_24_0.Vb1.t213 0.137822
R23353 two_stage_opamp_dummy_magic_24_0.Vb1.t69 two_stage_opamp_dummy_magic_24_0.Vb1.t60 0.137822
R23354 two_stage_opamp_dummy_magic_24_0.Vb1.t14 two_stage_opamp_dummy_magic_24_0.Vb1.t8 0.137822
R23355 two_stage_opamp_dummy_magic_24_0.Vb1.t76 two_stage_opamp_dummy_magic_24_0.Vb1.t68 0.137822
R23356 two_stage_opamp_dummy_magic_24_0.Vb1.t130 two_stage_opamp_dummy_magic_24_0.Vb1.t119 0.137822
R23357 two_stage_opamp_dummy_magic_24_0.Vb1.t75 two_stage_opamp_dummy_magic_24_0.Vb1.t67 0.137822
R23358 two_stage_opamp_dummy_magic_24_0.Vb1.t136 two_stage_opamp_dummy_magic_24_0.Vb1.t128 0.137822
R23359 two_stage_opamp_dummy_magic_24_0.Vb1.t197 two_stage_opamp_dummy_magic_24_0.Vb1.t188 0.137822
R23360 two_stage_opamp_dummy_magic_24_0.Vb1.t45 two_stage_opamp_dummy_magic_24_0.Vb1.t33 0.137822
R23361 two_stage_opamp_dummy_magic_24_0.Vb1.t205 two_stage_opamp_dummy_magic_24_0.Vb1.t195 0.137822
R23362 two_stage_opamp_dummy_magic_24_0.Vb1.t51 two_stage_opamp_dummy_magic_24_0.Vb1.t43 0.137822
R23363 two_stage_opamp_dummy_magic_24_0.Vb1.t110 two_stage_opamp_dummy_magic_24_0.Vb1.t104 0.137822
R23364 two_stage_opamp_dummy_magic_24_0.Vb1.t59 two_stage_opamp_dummy_magic_24_0.Vb1.t50 0.137822
R23365 two_stage_opamp_dummy_magic_24_0.Vb1.t121 two_stage_opamp_dummy_magic_24_0.Vb1.t109 0.137822
R23366 two_stage_opamp_dummy_magic_24_0.Vb1.t181 two_stage_opamp_dummy_magic_24_0.Vb1.t171 0.137822
R23367 two_stage_opamp_dummy_magic_24_0.Vb1.t129 two_stage_opamp_dummy_magic_24_0.Vb1.t118 0.137822
R23368 two_stage_opamp_dummy_magic_24_0.Vb1.t189 two_stage_opamp_dummy_magic_24_0.Vb1.t179 0.137822
R23369 two_stage_opamp_dummy_magic_24_0.Vb1.t34 two_stage_opamp_dummy_magic_24_0.Vb1.t25 0.137822
R23370 two_stage_opamp_dummy_magic_24_0.Vb1.t28 two_stage_opamp_dummy_magic_24_0.Vb1.t20 0.137822
R23371 two_stage_opamp_dummy_magic_24_0.Vb1.t28 two_stage_opamp_dummy_magic_24_0.Vb1.t170 0.1368
R23372 two_stage_opamp_dummy_magic_24_0.Vb1.t150 two_stage_opamp_dummy_magic_24_0.Vb1.t82 0.1368
R23373 two_stage_opamp_dummy_magic_24_0.Vb1.t214 two_stage_opamp_dummy_magic_24_0.Vb1.t143 0.1368
R23374 two_stage_opamp_dummy_magic_24_0.Vb1.t162 two_stage_opamp_dummy_magic_24_0.Vb1.t87 0.1368
R23375 two_stage_opamp_dummy_magic_24_0.Vb1.t9 two_stage_opamp_dummy_magic_24_0.Vb1.t148 0.1368
R23376 two_stage_opamp_dummy_magic_24_0.Vb1.t69 two_stage_opamp_dummy_magic_24_0.Vb1.t209 0.1368
R23377 two_stage_opamp_dummy_magic_24_0.Vb1.t14 two_stage_opamp_dummy_magic_24_0.Vb1.t159 0.1368
R23378 two_stage_opamp_dummy_magic_24_0.Vb1.t76 two_stage_opamp_dummy_magic_24_0.Vb1.t7 0.1368
R23379 two_stage_opamp_dummy_magic_24_0.Vb1.t130 two_stage_opamp_dummy_magic_24_0.Vb1.t57 0.1368
R23380 two_stage_opamp_dummy_magic_24_0.Vb1.t75 two_stage_opamp_dummy_magic_24_0.Vb1.t6 0.1368
R23381 two_stage_opamp_dummy_magic_24_0.Vb1.t136 two_stage_opamp_dummy_magic_24_0.Vb1.t66 0.1368
R23382 two_stage_opamp_dummy_magic_24_0.Vb1.t197 two_stage_opamp_dummy_magic_24_0.Vb1.t126 0.1368
R23383 two_stage_opamp_dummy_magic_24_0.Vb1.t45 two_stage_opamp_dummy_magic_24_0.Vb1.t186 0.1368
R23384 two_stage_opamp_dummy_magic_24_0.Vb1.t205 two_stage_opamp_dummy_magic_24_0.Vb1.t135 0.1368
R23385 two_stage_opamp_dummy_magic_24_0.Vb1.t51 two_stage_opamp_dummy_magic_24_0.Vb1.t194 0.1368
R23386 two_stage_opamp_dummy_magic_24_0.Vb1.t110 two_stage_opamp_dummy_magic_24_0.Vb1.t41 0.1368
R23387 two_stage_opamp_dummy_magic_24_0.Vb1.t59 two_stage_opamp_dummy_magic_24_0.Vb1.t204 0.1368
R23388 two_stage_opamp_dummy_magic_24_0.Vb1.t121 two_stage_opamp_dummy_magic_24_0.Vb1.t49 0.1368
R23389 two_stage_opamp_dummy_magic_24_0.Vb1.t181 two_stage_opamp_dummy_magic_24_0.Vb1.t108 0.1368
R23390 two_stage_opamp_dummy_magic_24_0.Vb1.t129 two_stage_opamp_dummy_magic_24_0.Vb1.t56 0.1368
R23391 two_stage_opamp_dummy_magic_24_0.Vb1.t189 two_stage_opamp_dummy_magic_24_0.Vb1.t116 0.1368
R23392 two_stage_opamp_dummy_magic_24_0.Vb1.t34 two_stage_opamp_dummy_magic_24_0.Vb1.t177 0.1368
R23393 two_stage_opamp_dummy_magic_24_0.Vb1.t88 two_stage_opamp_dummy_magic_24_0.Vb1.t16 0.1368
R23394 two_stage_opamp_dummy_magic_24_0.Vb1.t81 two_stage_opamp_dummy_magic_24_0.Vb1.t88 0.1368
R23395 two_stage_opamp_dummy_magic_24_0.Vb1.t91 two_stage_opamp_dummy_magic_24_0.Vb1.t83 0.1368
R23396 two_stage_opamp_dummy_magic_24_0.Vb3.n25 two_stage_opamp_dummy_magic_24_0.Vb3.t15 768.551
R23397 two_stage_opamp_dummy_magic_24_0.Vb3.n19 two_stage_opamp_dummy_magic_24_0.Vb3.t16 611.739
R23398 two_stage_opamp_dummy_magic_24_0.Vb3.n15 two_stage_opamp_dummy_magic_24_0.Vb3.t10 611.739
R23399 two_stage_opamp_dummy_magic_24_0.Vb3.n10 two_stage_opamp_dummy_magic_24_0.Vb3.t26 611.739
R23400 two_stage_opamp_dummy_magic_24_0.Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb3.t17 611.739
R23401 two_stage_opamp_dummy_magic_24_0.Vb3.n24 two_stage_opamp_dummy_magic_24_0.Vb3.n23 429.007
R23402 two_stage_opamp_dummy_magic_24_0.Vb3.n24 two_stage_opamp_dummy_magic_24_0.Vb3.n14 428.445
R23403 two_stage_opamp_dummy_magic_24_0.Vb3.n19 two_stage_opamp_dummy_magic_24_0.Vb3.t20 421.75
R23404 two_stage_opamp_dummy_magic_24_0.Vb3.n20 two_stage_opamp_dummy_magic_24_0.Vb3.t14 421.75
R23405 two_stage_opamp_dummy_magic_24_0.Vb3.n21 two_stage_opamp_dummy_magic_24_0.Vb3.t8 421.75
R23406 two_stage_opamp_dummy_magic_24_0.Vb3.n22 two_stage_opamp_dummy_magic_24_0.Vb3.t25 421.75
R23407 two_stage_opamp_dummy_magic_24_0.Vb3.n15 two_stage_opamp_dummy_magic_24_0.Vb3.t12 421.75
R23408 two_stage_opamp_dummy_magic_24_0.Vb3.n16 two_stage_opamp_dummy_magic_24_0.Vb3.t18 421.75
R23409 two_stage_opamp_dummy_magic_24_0.Vb3.n17 two_stage_opamp_dummy_magic_24_0.Vb3.t23 421.75
R23410 two_stage_opamp_dummy_magic_24_0.Vb3.n18 two_stage_opamp_dummy_magic_24_0.Vb3.t21 421.75
R23411 two_stage_opamp_dummy_magic_24_0.Vb3.n10 two_stage_opamp_dummy_magic_24_0.Vb3.t28 421.75
R23412 two_stage_opamp_dummy_magic_24_0.Vb3.n11 two_stage_opamp_dummy_magic_24_0.Vb3.t24 421.75
R23413 two_stage_opamp_dummy_magic_24_0.Vb3.n12 two_stage_opamp_dummy_magic_24_0.Vb3.t19 421.75
R23414 two_stage_opamp_dummy_magic_24_0.Vb3.n13 two_stage_opamp_dummy_magic_24_0.Vb3.t13 421.75
R23415 two_stage_opamp_dummy_magic_24_0.Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb3.t22 421.75
R23416 two_stage_opamp_dummy_magic_24_0.Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb3.t27 421.75
R23417 two_stage_opamp_dummy_magic_24_0.Vb3.n8 two_stage_opamp_dummy_magic_24_0.Vb3.t9 421.75
R23418 two_stage_opamp_dummy_magic_24_0.Vb3.n9 two_stage_opamp_dummy_magic_24_0.Vb3.t11 421.75
R23419 two_stage_opamp_dummy_magic_24_0.Vb3.n20 two_stage_opamp_dummy_magic_24_0.Vb3.n19 167.094
R23420 two_stage_opamp_dummy_magic_24_0.Vb3.n21 two_stage_opamp_dummy_magic_24_0.Vb3.n20 167.094
R23421 two_stage_opamp_dummy_magic_24_0.Vb3.n22 two_stage_opamp_dummy_magic_24_0.Vb3.n21 167.094
R23422 two_stage_opamp_dummy_magic_24_0.Vb3.n16 two_stage_opamp_dummy_magic_24_0.Vb3.n15 167.094
R23423 two_stage_opamp_dummy_magic_24_0.Vb3.n17 two_stage_opamp_dummy_magic_24_0.Vb3.n16 167.094
R23424 two_stage_opamp_dummy_magic_24_0.Vb3.n18 two_stage_opamp_dummy_magic_24_0.Vb3.n17 167.094
R23425 two_stage_opamp_dummy_magic_24_0.Vb3.n11 two_stage_opamp_dummy_magic_24_0.Vb3.n10 167.094
R23426 two_stage_opamp_dummy_magic_24_0.Vb3.n12 two_stage_opamp_dummy_magic_24_0.Vb3.n11 167.094
R23427 two_stage_opamp_dummy_magic_24_0.Vb3.n13 two_stage_opamp_dummy_magic_24_0.Vb3.n12 167.094
R23428 two_stage_opamp_dummy_magic_24_0.Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb3.n6 167.094
R23429 two_stage_opamp_dummy_magic_24_0.Vb3.n8 two_stage_opamp_dummy_magic_24_0.Vb3.n7 167.094
R23430 two_stage_opamp_dummy_magic_24_0.Vb3.n9 two_stage_opamp_dummy_magic_24_0.Vb3.n8 167.094
R23431 two_stage_opamp_dummy_magic_24_0.Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb3.n0 139.639
R23432 two_stage_opamp_dummy_magic_24_0.Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb3.n1 139.638
R23433 two_stage_opamp_dummy_magic_24_0.Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb3.n3 134.577
R23434 two_stage_opamp_dummy_magic_24_0.Vb3.n26 two_stage_opamp_dummy_magic_24_0.Vb3.n5 73.3151
R23435 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_24_0.Vb3.n26 69.5943
R23436 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_24_0.Vb3.n4 43.063
R23437 two_stage_opamp_dummy_magic_24_0.Vb3.n23 two_stage_opamp_dummy_magic_24_0.Vb3.n22 35.3472
R23438 two_stage_opamp_dummy_magic_24_0.Vb3.n23 two_stage_opamp_dummy_magic_24_0.Vb3.n18 35.3472
R23439 two_stage_opamp_dummy_magic_24_0.Vb3.n14 two_stage_opamp_dummy_magic_24_0.Vb3.n13 35.3472
R23440 two_stage_opamp_dummy_magic_24_0.Vb3.n14 two_stage_opamp_dummy_magic_24_0.Vb3.n9 35.3472
R23441 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.t1 24.0005
R23442 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.t7 24.0005
R23443 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.t0 24.0005
R23444 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.t5 24.0005
R23445 two_stage_opamp_dummy_magic_24_0.Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb3.t6 24.0005
R23446 two_stage_opamp_dummy_magic_24_0.Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb3.t3 24.0005
R23447 two_stage_opamp_dummy_magic_24_0.Vb3.n25 two_stage_opamp_dummy_magic_24_0.Vb3.n24 15.313
R23448 two_stage_opamp_dummy_magic_24_0.Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb3.t2 11.2576
R23449 two_stage_opamp_dummy_magic_24_0.Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb3.t4 11.2576
R23450 two_stage_opamp_dummy_magic_24_0.Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb3.n2 4.5005
R23451 two_stage_opamp_dummy_magic_24_0.Vb3.n26 two_stage_opamp_dummy_magic_24_0.Vb3.n25 1.21925
R23452 two_stage_opamp_dummy_magic_24_0.VD4.n14 two_stage_opamp_dummy_magic_24_0.VD4.t32 672.293
R23453 two_stage_opamp_dummy_magic_24_0.VD4.n29 two_stage_opamp_dummy_magic_24_0.VD4.t35 672.293
R23454 two_stage_opamp_dummy_magic_24_0.VD4.n28 two_stage_opamp_dummy_magic_24_0.VD4.t36 213.131
R23455 two_stage_opamp_dummy_magic_24_0.VD4.t33 two_stage_opamp_dummy_magic_24_0.VD4.n27 213.131
R23456 two_stage_opamp_dummy_magic_24_0.VD4.t36 two_stage_opamp_dummy_magic_24_0.VD4.t6 146.155
R23457 two_stage_opamp_dummy_magic_24_0.VD4.t6 two_stage_opamp_dummy_magic_24_0.VD4.t18 146.155
R23458 two_stage_opamp_dummy_magic_24_0.VD4.t18 two_stage_opamp_dummy_magic_24_0.VD4.t12 146.155
R23459 two_stage_opamp_dummy_magic_24_0.VD4.t12 two_stage_opamp_dummy_magic_24_0.VD4.t10 146.155
R23460 two_stage_opamp_dummy_magic_24_0.VD4.t10 two_stage_opamp_dummy_magic_24_0.VD4.t0 146.155
R23461 two_stage_opamp_dummy_magic_24_0.VD4.t0 two_stage_opamp_dummy_magic_24_0.VD4.t8 146.155
R23462 two_stage_opamp_dummy_magic_24_0.VD4.t8 two_stage_opamp_dummy_magic_24_0.VD4.t2 146.155
R23463 two_stage_opamp_dummy_magic_24_0.VD4.t2 two_stage_opamp_dummy_magic_24_0.VD4.t16 146.155
R23464 two_stage_opamp_dummy_magic_24_0.VD4.t16 two_stage_opamp_dummy_magic_24_0.VD4.t4 146.155
R23465 two_stage_opamp_dummy_magic_24_0.VD4.t4 two_stage_opamp_dummy_magic_24_0.VD4.t14 146.155
R23466 two_stage_opamp_dummy_magic_24_0.VD4.t14 two_stage_opamp_dummy_magic_24_0.VD4.t33 146.155
R23467 two_stage_opamp_dummy_magic_24_0.VD4.n28 two_stage_opamp_dummy_magic_24_0.VD4.t37 76.2576
R23468 two_stage_opamp_dummy_magic_24_0.VD4.n27 two_stage_opamp_dummy_magic_24_0.VD4.t34 76.2576
R23469 two_stage_opamp_dummy_magic_24_0.VD4.n26 two_stage_opamp_dummy_magic_24_0.VD4.n25 66.9922
R23470 two_stage_opamp_dummy_magic_24_0.VD4.n34 two_stage_opamp_dummy_magic_24_0.VD4.n24 66.9922
R23471 two_stage_opamp_dummy_magic_24_0.VD4.n39 two_stage_opamp_dummy_magic_24_0.VD4.n21 66.9922
R23472 two_stage_opamp_dummy_magic_24_0.VD4.n44 two_stage_opamp_dummy_magic_24_0.VD4.n18 66.9922
R23473 two_stage_opamp_dummy_magic_24_0.VD4.n16 two_stage_opamp_dummy_magic_24_0.VD4.n15 66.9922
R23474 two_stage_opamp_dummy_magic_24_0.VD4.n56 two_stage_opamp_dummy_magic_24_0.VD4.n55 66.0338
R23475 two_stage_opamp_dummy_magic_24_0.VD4.n12 two_stage_opamp_dummy_magic_24_0.VD4.n11 66.0338
R23476 two_stage_opamp_dummy_magic_24_0.VD4.n58 two_stage_opamp_dummy_magic_24_0.VD4.n57 66.0338
R23477 two_stage_opamp_dummy_magic_24_0.VD4.n61 two_stage_opamp_dummy_magic_24_0.VD4.n60 66.0338
R23478 two_stage_opamp_dummy_magic_24_0.VD4.n66 two_stage_opamp_dummy_magic_24_0.VD4.n65 66.0338
R23479 two_stage_opamp_dummy_magic_24_0.VD4.n70 two_stage_opamp_dummy_magic_24_0.VD4.n69 66.0338
R23480 two_stage_opamp_dummy_magic_24_0.VD4.n55 two_stage_opamp_dummy_magic_24_0.VD4.t20 11.2576
R23481 two_stage_opamp_dummy_magic_24_0.VD4.n55 two_stage_opamp_dummy_magic_24_0.VD4.t27 11.2576
R23482 two_stage_opamp_dummy_magic_24_0.VD4.n11 two_stage_opamp_dummy_magic_24_0.VD4.t25 11.2576
R23483 two_stage_opamp_dummy_magic_24_0.VD4.n11 two_stage_opamp_dummy_magic_24_0.VD4.t28 11.2576
R23484 two_stage_opamp_dummy_magic_24_0.VD4.n57 two_stage_opamp_dummy_magic_24_0.VD4.t30 11.2576
R23485 two_stage_opamp_dummy_magic_24_0.VD4.n57 two_stage_opamp_dummy_magic_24_0.VD4.t21 11.2576
R23486 two_stage_opamp_dummy_magic_24_0.VD4.n60 two_stage_opamp_dummy_magic_24_0.VD4.t26 11.2576
R23487 two_stage_opamp_dummy_magic_24_0.VD4.n60 two_stage_opamp_dummy_magic_24_0.VD4.t29 11.2576
R23488 two_stage_opamp_dummy_magic_24_0.VD4.n65 two_stage_opamp_dummy_magic_24_0.VD4.t24 11.2576
R23489 two_stage_opamp_dummy_magic_24_0.VD4.n65 two_stage_opamp_dummy_magic_24_0.VD4.t23 11.2576
R23490 two_stage_opamp_dummy_magic_24_0.VD4.n25 two_stage_opamp_dummy_magic_24_0.VD4.t7 11.2576
R23491 two_stage_opamp_dummy_magic_24_0.VD4.n25 two_stage_opamp_dummy_magic_24_0.VD4.t19 11.2576
R23492 two_stage_opamp_dummy_magic_24_0.VD4.n24 two_stage_opamp_dummy_magic_24_0.VD4.t13 11.2576
R23493 two_stage_opamp_dummy_magic_24_0.VD4.n24 two_stage_opamp_dummy_magic_24_0.VD4.t11 11.2576
R23494 two_stage_opamp_dummy_magic_24_0.VD4.n21 two_stage_opamp_dummy_magic_24_0.VD4.t1 11.2576
R23495 two_stage_opamp_dummy_magic_24_0.VD4.n21 two_stage_opamp_dummy_magic_24_0.VD4.t9 11.2576
R23496 two_stage_opamp_dummy_magic_24_0.VD4.n18 two_stage_opamp_dummy_magic_24_0.VD4.t3 11.2576
R23497 two_stage_opamp_dummy_magic_24_0.VD4.n18 two_stage_opamp_dummy_magic_24_0.VD4.t17 11.2576
R23498 two_stage_opamp_dummy_magic_24_0.VD4.n15 two_stage_opamp_dummy_magic_24_0.VD4.t5 11.2576
R23499 two_stage_opamp_dummy_magic_24_0.VD4.n15 two_stage_opamp_dummy_magic_24_0.VD4.t15 11.2576
R23500 two_stage_opamp_dummy_magic_24_0.VD4.t31 two_stage_opamp_dummy_magic_24_0.VD4.n70 11.2576
R23501 two_stage_opamp_dummy_magic_24_0.VD4.n70 two_stage_opamp_dummy_magic_24_0.VD4.t22 11.2576
R23502 two_stage_opamp_dummy_magic_24_0.VD4.n58 two_stage_opamp_dummy_magic_24_0.VD4.n10 5.91717
R23503 two_stage_opamp_dummy_magic_24_0.VD4.n56 two_stage_opamp_dummy_magic_24_0.VD4.n9 5.91717
R23504 two_stage_opamp_dummy_magic_24_0.VD4.n12 two_stage_opamp_dummy_magic_24_0.VD4.n9 5.29217
R23505 two_stage_opamp_dummy_magic_24_0.VD4.n61 two_stage_opamp_dummy_magic_24_0.VD4.n10 5.29217
R23506 two_stage_opamp_dummy_magic_24_0.VD4.n67 two_stage_opamp_dummy_magic_24_0.VD4.n66 5.29217
R23507 two_stage_opamp_dummy_magic_24_0.VD4.n69 two_stage_opamp_dummy_magic_24_0.VD4.n68 5.29217
R23508 two_stage_opamp_dummy_magic_24_0.VD4.n53 two_stage_opamp_dummy_magic_24_0.VD4.n52 1.5005
R23509 two_stage_opamp_dummy_magic_24_0.VD4.n51 two_stage_opamp_dummy_magic_24_0.VD4.n13 1.5005
R23510 two_stage_opamp_dummy_magic_24_0.VD4.n50 two_stage_opamp_dummy_magic_24_0.VD4.n49 1.5005
R23511 two_stage_opamp_dummy_magic_24_0.VD4.n48 two_stage_opamp_dummy_magic_24_0.VD4.n16 1.5005
R23512 two_stage_opamp_dummy_magic_24_0.VD4.n47 two_stage_opamp_dummy_magic_24_0.VD4.n46 1.5005
R23513 two_stage_opamp_dummy_magic_24_0.VD4.n45 two_stage_opamp_dummy_magic_24_0.VD4.n17 1.5005
R23514 two_stage_opamp_dummy_magic_24_0.VD4.n44 two_stage_opamp_dummy_magic_24_0.VD4.n43 1.5005
R23515 two_stage_opamp_dummy_magic_24_0.VD4.n42 two_stage_opamp_dummy_magic_24_0.VD4.n19 1.5005
R23516 two_stage_opamp_dummy_magic_24_0.VD4.n41 two_stage_opamp_dummy_magic_24_0.VD4.n40 1.5005
R23517 two_stage_opamp_dummy_magic_24_0.VD4.n39 two_stage_opamp_dummy_magic_24_0.VD4.n20 1.5005
R23518 two_stage_opamp_dummy_magic_24_0.VD4.n38 two_stage_opamp_dummy_magic_24_0.VD4.n37 1.5005
R23519 two_stage_opamp_dummy_magic_24_0.VD4.n36 two_stage_opamp_dummy_magic_24_0.VD4.n22 1.5005
R23520 two_stage_opamp_dummy_magic_24_0.VD4.n35 two_stage_opamp_dummy_magic_24_0.VD4.n34 1.5005
R23521 two_stage_opamp_dummy_magic_24_0.VD4.n33 two_stage_opamp_dummy_magic_24_0.VD4.n23 1.5005
R23522 two_stage_opamp_dummy_magic_24_0.VD4.n32 two_stage_opamp_dummy_magic_24_0.VD4.n31 1.5005
R23523 two_stage_opamp_dummy_magic_24_0.VD4.n0 two_stage_opamp_dummy_magic_24_0.VD4.n1 0.740726
R23524 two_stage_opamp_dummy_magic_24_0.VD4.n64 two_stage_opamp_dummy_magic_24_0.VD4.n63 1.5005
R23525 two_stage_opamp_dummy_magic_24_0.VD4.n6 two_stage_opamp_dummy_magic_24_0.VD4.n5 0.740726
R23526 two_stage_opamp_dummy_magic_24_0.VD4.n8 two_stage_opamp_dummy_magic_24_0.VD4.n7 0.740726
R23527 two_stage_opamp_dummy_magic_24_0.VD4.n4 two_stage_opamp_dummy_magic_24_0.VD4.n3 0.740726
R23528 two_stage_opamp_dummy_magic_24_0.VD4.n2 two_stage_opamp_dummy_magic_24_0.VD4.n54 1.5005
R23529 two_stage_opamp_dummy_magic_24_0.VD4.n29 two_stage_opamp_dummy_magic_24_0.VD4.n28 1.03383
R23530 two_stage_opamp_dummy_magic_24_0.VD4.n27 two_stage_opamp_dummy_magic_24_0.VD4.n14 1.03383
R23531 two_stage_opamp_dummy_magic_24_0.VD4.n30 two_stage_opamp_dummy_magic_24_0.VD4.n29 1.02322
R23532 two_stage_opamp_dummy_magic_24_0.VD4.n59 two_stage_opamp_dummy_magic_24_0.VD4.n58 1.02322
R23533 two_stage_opamp_dummy_magic_24_0.VD4.n8 two_stage_opamp_dummy_magic_24_0.VD4.n12 0.958833
R23534 two_stage_opamp_dummy_magic_24_0.VD4.n62 two_stage_opamp_dummy_magic_24_0.VD4.n61 0.958833
R23535 two_stage_opamp_dummy_magic_24_0.VD4.n66 two_stage_opamp_dummy_magic_24_0.VD4.n64 0.958833
R23536 two_stage_opamp_dummy_magic_24_0.VD4.n52 two_stage_opamp_dummy_magic_24_0.VD4.n14 0.958833
R23537 two_stage_opamp_dummy_magic_24_0.VD4.n2 two_stage_opamp_dummy_magic_24_0.VD4.n56 0.958833
R23538 two_stage_opamp_dummy_magic_24_0.VD4.n69 two_stage_opamp_dummy_magic_24_0.VD4.n5 0.958833
R23539 two_stage_opamp_dummy_magic_24_0.VD4.n68 two_stage_opamp_dummy_magic_24_0.VD4.n67 0.6255
R23540 two_stage_opamp_dummy_magic_24_0.VD4.n67 two_stage_opamp_dummy_magic_24_0.VD4.n10 0.6255
R23541 two_stage_opamp_dummy_magic_24_0.VD4.n68 two_stage_opamp_dummy_magic_24_0.VD4.n9 0.6255
R23542 two_stage_opamp_dummy_magic_24_0.VD4.n54 two_stage_opamp_dummy_magic_24_0.VD4.n53 0.443208
R23543 two_stage_opamp_dummy_magic_24_0.VD4.n31 two_stage_opamp_dummy_magic_24_0.VD4.n30 0.427973
R23544 two_stage_opamp_dummy_magic_24_0.VD4.n0 two_stage_opamp_dummy_magic_24_0.VD4.n59 0.427973
R23545 two_stage_opamp_dummy_magic_24_0.VD4.n5 two_stage_opamp_dummy_magic_24_0.VD4.n8 0.0838333
R23546 two_stage_opamp_dummy_magic_24_0.VD4.n30 two_stage_opamp_dummy_magic_24_0.VD4.n26 0.0587394
R23547 two_stage_opamp_dummy_magic_24_0.VD4.n62 two_stage_opamp_dummy_magic_24_0.VD4.n59 0.0587394
R23548 two_stage_opamp_dummy_magic_24_0.VD4.n64 two_stage_opamp_dummy_magic_24_0.VD4.n1 0.0632146
R23549 two_stage_opamp_dummy_magic_24_0.VD4.n62 two_stage_opamp_dummy_magic_24_0.VD4.n1 0.0632146
R23550 two_stage_opamp_dummy_magic_24_0.VD4.n32 two_stage_opamp_dummy_magic_24_0.VD4.n26 0.0421667
R23551 two_stage_opamp_dummy_magic_24_0.VD4.n33 two_stage_opamp_dummy_magic_24_0.VD4.n32 0.0421667
R23552 two_stage_opamp_dummy_magic_24_0.VD4.n34 two_stage_opamp_dummy_magic_24_0.VD4.n33 0.0421667
R23553 two_stage_opamp_dummy_magic_24_0.VD4.n34 two_stage_opamp_dummy_magic_24_0.VD4.n22 0.0421667
R23554 two_stage_opamp_dummy_magic_24_0.VD4.n38 two_stage_opamp_dummy_magic_24_0.VD4.n22 0.0421667
R23555 two_stage_opamp_dummy_magic_24_0.VD4.n39 two_stage_opamp_dummy_magic_24_0.VD4.n38 0.0421667
R23556 two_stage_opamp_dummy_magic_24_0.VD4.n40 two_stage_opamp_dummy_magic_24_0.VD4.n39 0.0421667
R23557 two_stage_opamp_dummy_magic_24_0.VD4.n40 two_stage_opamp_dummy_magic_24_0.VD4.n19 0.0421667
R23558 two_stage_opamp_dummy_magic_24_0.VD4.n44 two_stage_opamp_dummy_magic_24_0.VD4.n19 0.0421667
R23559 two_stage_opamp_dummy_magic_24_0.VD4.n45 two_stage_opamp_dummy_magic_24_0.VD4.n44 0.0421667
R23560 two_stage_opamp_dummy_magic_24_0.VD4.n46 two_stage_opamp_dummy_magic_24_0.VD4.n45 0.0421667
R23561 two_stage_opamp_dummy_magic_24_0.VD4.n46 two_stage_opamp_dummy_magic_24_0.VD4.n16 0.0421667
R23562 two_stage_opamp_dummy_magic_24_0.VD4.n50 two_stage_opamp_dummy_magic_24_0.VD4.n16 0.0421667
R23563 two_stage_opamp_dummy_magic_24_0.VD4.n51 two_stage_opamp_dummy_magic_24_0.VD4.n50 0.0421667
R23564 two_stage_opamp_dummy_magic_24_0.VD4.n52 two_stage_opamp_dummy_magic_24_0.VD4.n51 0.0421667
R23565 two_stage_opamp_dummy_magic_24_0.VD4.n31 two_stage_opamp_dummy_magic_24_0.VD4.n23 0.0421667
R23566 two_stage_opamp_dummy_magic_24_0.VD4.n35 two_stage_opamp_dummy_magic_24_0.VD4.n23 0.0421667
R23567 two_stage_opamp_dummy_magic_24_0.VD4.n36 two_stage_opamp_dummy_magic_24_0.VD4.n35 0.0421667
R23568 two_stage_opamp_dummy_magic_24_0.VD4.n37 two_stage_opamp_dummy_magic_24_0.VD4.n36 0.0421667
R23569 two_stage_opamp_dummy_magic_24_0.VD4.n37 two_stage_opamp_dummy_magic_24_0.VD4.n20 0.0421667
R23570 two_stage_opamp_dummy_magic_24_0.VD4.n41 two_stage_opamp_dummy_magic_24_0.VD4.n20 0.0421667
R23571 two_stage_opamp_dummy_magic_24_0.VD4.n42 two_stage_opamp_dummy_magic_24_0.VD4.n41 0.0421667
R23572 two_stage_opamp_dummy_magic_24_0.VD4.n43 two_stage_opamp_dummy_magic_24_0.VD4.n42 0.0421667
R23573 two_stage_opamp_dummy_magic_24_0.VD4.n43 two_stage_opamp_dummy_magic_24_0.VD4.n17 0.0421667
R23574 two_stage_opamp_dummy_magic_24_0.VD4.n47 two_stage_opamp_dummy_magic_24_0.VD4.n17 0.0421667
R23575 two_stage_opamp_dummy_magic_24_0.VD4.n48 two_stage_opamp_dummy_magic_24_0.VD4.n47 0.0421667
R23576 two_stage_opamp_dummy_magic_24_0.VD4.n49 two_stage_opamp_dummy_magic_24_0.VD4.n48 0.0421667
R23577 two_stage_opamp_dummy_magic_24_0.VD4.n49 two_stage_opamp_dummy_magic_24_0.VD4.n13 0.0421667
R23578 two_stage_opamp_dummy_magic_24_0.VD4.n53 two_stage_opamp_dummy_magic_24_0.VD4.n13 0.0421667
R23579 two_stage_opamp_dummy_magic_24_0.VD4.n4 two_stage_opamp_dummy_magic_24_0.VD4.n54 0.0632146
R23580 two_stage_opamp_dummy_magic_24_0.VD4.n7 two_stage_opamp_dummy_magic_24_0.VD4.n4 0.0842626
R23581 two_stage_opamp_dummy_magic_24_0.VD4.n7 two_stage_opamp_dummy_magic_24_0.VD4.n6 0.0842626
R23582 two_stage_opamp_dummy_magic_24_0.VD4.n63 two_stage_opamp_dummy_magic_24_0.VD4.n6 0.146548
R23583 two_stage_opamp_dummy_magic_24_0.VD4.n8 two_stage_opamp_dummy_magic_24_0.VD4.n3 0.0838333
R23584 two_stage_opamp_dummy_magic_24_0.VD4.n3 two_stage_opamp_dummy_magic_24_0.VD4.n2 0.0838333
R23585 two_stage_opamp_dummy_magic_24_0.VD4.n63 two_stage_opamp_dummy_magic_24_0.VD4.n0 0.0838333
R23586 VOUT+.n19 VOUT+.t2 110.191
R23587 VOUT+.n48 VOUT+.n47 34.9935
R23588 VOUT+.n46 VOUT+.n45 34.9935
R23589 VOUT+.n60 VOUT+.n59 34.9935
R23590 VOUT+.n56 VOUT+.n55 34.9935
R23591 VOUT+.n53 VOUT+.n52 34.9935
R23592 VOUT+.n50 VOUT+.n49 34.9935
R23593 VOUT+.n2 VOUT+.n1 9.73997
R23594 VOUT+.n6 VOUT+.n5 9.73997
R23595 VOUT+.n9 VOUT+.n8 9.73997
R23596 VOUT+.n7 VOUT+.n6 6.64633
R23597 VOUT+.n7 VOUT+.n2 6.64633
R23598 VOUT+.n47 VOUT+.t0 6.56717
R23599 VOUT+.n47 VOUT+.t12 6.56717
R23600 VOUT+.n45 VOUT+.t13 6.56717
R23601 VOUT+.n45 VOUT+.t3 6.56717
R23602 VOUT+.n59 VOUT+.t6 6.56717
R23603 VOUT+.n59 VOUT+.t1 6.56717
R23604 VOUT+.n55 VOUT+.t10 6.56717
R23605 VOUT+.n55 VOUT+.t8 6.56717
R23606 VOUT+.n52 VOUT+.t11 6.56717
R23607 VOUT+.n52 VOUT+.t9 6.56717
R23608 VOUT+.n49 VOUT+.t5 6.56717
R23609 VOUT+.n49 VOUT+.t7 6.56717
R23610 VOUT+.n58 VOUT+.n46 6.3755
R23611 VOUT+.n51 VOUT+.n48 6.3755
R23612 VOUT+.n9 VOUT+.n7 6.02133
R23613 VOUT+.n60 VOUT+.n58 5.813
R23614 VOUT+.n57 VOUT+.n56 5.813
R23615 VOUT+.n54 VOUT+.n53 5.813
R23616 VOUT+.n51 VOUT+.n50 5.813
R23617 VOUT+.n61 VOUT+.n37 5.063
R23618 VOUT+.n64 VOUT+.n44 5.063
R23619 VOUT+.n124 VOUT+.t113 4.8295
R23620 VOUT+.n126 VOUT+.t78 4.8295
R23621 VOUT+.n127 VOUT+.t119 4.8295
R23622 VOUT+.n128 VOUT+.t24 4.8295
R23623 VOUT+.n139 VOUT+.t67 4.8295
R23624 VOUT+.n141 VOUT+.t93 4.8295
R23625 VOUT+.n142 VOUT+.t111 4.8295
R23626 VOUT+.n144 VOUT+.t45 4.8295
R23627 VOUT+.n145 VOUT+.t70 4.8295
R23628 VOUT+.n147 VOUT+.t147 4.8295
R23629 VOUT+.n148 VOUT+.t33 4.8295
R23630 VOUT+.n150 VOUT+.t37 4.8295
R23631 VOUT+.n151 VOUT+.t66 4.8295
R23632 VOUT+.n153 VOUT+.t142 4.8295
R23633 VOUT+.n154 VOUT+.t28 4.8295
R23634 VOUT+.n156 VOUT+.t105 4.8295
R23635 VOUT+.n157 VOUT+.t131 4.8295
R23636 VOUT+.n159 VOUT+.t137 4.8295
R23637 VOUT+.n160 VOUT+.t23 4.8295
R23638 VOUT+.n162 VOUT+.t97 4.8295
R23639 VOUT+.n163 VOUT+.t124 4.8295
R23640 VOUT+.n165 VOUT+.t55 4.8295
R23641 VOUT+.n166 VOUT+.t84 4.8295
R23642 VOUT+.n168 VOUT+.t20 4.8295
R23643 VOUT+.n169 VOUT+.t46 4.8295
R23644 VOUT+.n98 VOUT+.t90 4.8295
R23645 VOUT+.n110 VOUT+.t126 4.8295
R23646 VOUT+.n112 VOUT+.t75 4.8295
R23647 VOUT+.n113 VOUT+.t106 4.8295
R23648 VOUT+.n115 VOUT+.t146 4.8295
R23649 VOUT+.n116 VOUT+.t32 4.8295
R23650 VOUT+.n118 VOUT+.t114 4.8295
R23651 VOUT+.n119 VOUT+.t143 4.8295
R23652 VOUT+.n121 VOUT+.t152 4.8295
R23653 VOUT+.n122 VOUT+.t38 4.8295
R23654 VOUT+.n171 VOUT+.t77 4.8295
R23655 VOUT+.n132 VOUT+.t81 4.8154
R23656 VOUT+.n131 VOUT+.t122 4.8154
R23657 VOUT+.n130 VOUT+.t104 4.8154
R23658 VOUT+.n129 VOUT+.t139 4.8154
R23659 VOUT+.n138 VOUT+.t121 4.806
R23660 VOUT+.n137 VOUT+.t101 4.806
R23661 VOUT+.n136 VOUT+.t138 4.806
R23662 VOUT+.n135 VOUT+.t31 4.806
R23663 VOUT+.n134 VOUT+.t156 4.806
R23664 VOUT+.n133 VOUT+.t47 4.806
R23665 VOUT+.n133 VOUT+.t52 4.806
R23666 VOUT+.n132 VOUT+.t86 4.806
R23667 VOUT+.n131 VOUT+.t127 4.806
R23668 VOUT+.n130 VOUT+.t110 4.806
R23669 VOUT+.n129 VOUT+.t144 4.806
R23670 VOUT+.n109 VOUT+.t154 4.806
R23671 VOUT+.n108 VOUT+.t61 4.806
R23672 VOUT+.n107 VOUT+.t99 4.806
R23673 VOUT+.n106 VOUT+.t133 4.806
R23674 VOUT+.n105 VOUT+.t40 4.806
R23675 VOUT+.n104 VOUT+.t72 4.806
R23676 VOUT+.n103 VOUT+.t116 4.806
R23677 VOUT+.n102 VOUT+.t149 4.806
R23678 VOUT+.n101 VOUT+.t56 4.806
R23679 VOUT+.n100 VOUT+.t92 4.806
R23680 VOUT+.n125 VOUT+.t80 4.5005
R23681 VOUT+.n124 VOUT+.t73 4.5005
R23682 VOUT+.n126 VOUT+.t134 4.5005
R23683 VOUT+.n127 VOUT+.t26 4.5005
R23684 VOUT+.n128 VOUT+.t150 4.5005
R23685 VOUT+.n129 VOUT+.t107 4.5005
R23686 VOUT+.n130 VOUT+.t63 4.5005
R23687 VOUT+.n131 VOUT+.t85 4.5005
R23688 VOUT+.n132 VOUT+.t48 4.5005
R23689 VOUT+.n133 VOUT+.t155 4.5005
R23690 VOUT+.n134 VOUT+.t117 4.5005
R23691 VOUT+.n135 VOUT+.t136 4.5005
R23692 VOUT+.n136 VOUT+.t100 4.5005
R23693 VOUT+.n137 VOUT+.t57 4.5005
R23694 VOUT+.n138 VOUT+.t79 4.5005
R23695 VOUT+.n140 VOUT+.t41 4.5005
R23696 VOUT+.n139 VOUT+.t34 4.5005
R23697 VOUT+.n141 VOUT+.t120 4.5005
R23698 VOUT+.n143 VOUT+.t74 4.5005
R23699 VOUT+.n142 VOUT+.t68 4.5005
R23700 VOUT+.n144 VOUT+.t135 4.5005
R23701 VOUT+.n146 VOUT+.t102 4.5005
R23702 VOUT+.n145 VOUT+.t69 4.5005
R23703 VOUT+.n147 VOUT+.t96 4.5005
R23704 VOUT+.n149 VOUT+.t59 4.5005
R23705 VOUT+.n148 VOUT+.t30 4.5005
R23706 VOUT+.n150 VOUT+.t129 4.5005
R23707 VOUT+.n152 VOUT+.t94 4.5005
R23708 VOUT+.n151 VOUT+.t65 4.5005
R23709 VOUT+.n153 VOUT+.t88 4.5005
R23710 VOUT+.n155 VOUT+.t54 4.5005
R23711 VOUT+.n154 VOUT+.t27 4.5005
R23712 VOUT+.n156 VOUT+.t50 4.5005
R23713 VOUT+.n158 VOUT+.t19 4.5005
R23714 VOUT+.n157 VOUT+.t130 4.5005
R23715 VOUT+.n159 VOUT+.t82 4.5005
R23716 VOUT+.n161 VOUT+.t49 4.5005
R23717 VOUT+.n160 VOUT+.t22 4.5005
R23718 VOUT+.n162 VOUT+.t42 4.5005
R23719 VOUT+.n164 VOUT+.t151 4.5005
R23720 VOUT+.n163 VOUT+.t123 4.5005
R23721 VOUT+.n165 VOUT+.t145 4.5005
R23722 VOUT+.n167 VOUT+.t112 4.5005
R23723 VOUT+.n166 VOUT+.t83 4.5005
R23724 VOUT+.n168 VOUT+.t109 4.5005
R23725 VOUT+.n170 VOUT+.t64 4.5005
R23726 VOUT+.n169 VOUT+.t43 4.5005
R23727 VOUT+.n99 VOUT+.t118 4.5005
R23728 VOUT+.n98 VOUT+.t89 4.5005
R23729 VOUT+.n100 VOUT+.t128 4.5005
R23730 VOUT+.n101 VOUT+.t91 4.5005
R23731 VOUT+.n102 VOUT+.t39 4.5005
R23732 VOUT+.n103 VOUT+.t148 4.5005
R23733 VOUT+.n104 VOUT+.t115 4.5005
R23734 VOUT+.n105 VOUT+.t71 4.5005
R23735 VOUT+.n106 VOUT+.t25 4.5005
R23736 VOUT+.n107 VOUT+.t132 4.5005
R23737 VOUT+.n108 VOUT+.t98 4.5005
R23738 VOUT+.n109 VOUT+.t44 4.5005
R23739 VOUT+.n111 VOUT+.t153 4.5005
R23740 VOUT+.n110 VOUT+.t125 4.5005
R23741 VOUT+.n112 VOUT+.t35 4.5005
R23742 VOUT+.n114 VOUT+.t87 4.5005
R23743 VOUT+.n113 VOUT+.t53 4.5005
R23744 VOUT+.n115 VOUT+.t95 4.5005
R23745 VOUT+.n117 VOUT+.t58 4.5005
R23746 VOUT+.n116 VOUT+.t29 4.5005
R23747 VOUT+.n118 VOUT+.t60 4.5005
R23748 VOUT+.n120 VOUT+.t21 4.5005
R23749 VOUT+.n119 VOUT+.t141 4.5005
R23750 VOUT+.n121 VOUT+.t103 4.5005
R23751 VOUT+.n123 VOUT+.t62 4.5005
R23752 VOUT+.n122 VOUT+.t36 4.5005
R23753 VOUT+.n173 VOUT+.t140 4.5005
R23754 VOUT+.n172 VOUT+.t108 4.5005
R23755 VOUT+.n171 VOUT+.t76 4.5005
R23756 VOUT+.n174 VOUT+.t51 4.5005
R23757 VOUT+.n61 VOUT+.n38 4.5005
R23758 VOUT+.n62 VOUT+.n41 4.5005
R23759 VOUT+.n63 VOUT+.n42 4.5005
R23760 VOUT+.n65 VOUT+.n64 4.5005
R23761 VOUT+.n88 VOUT+.n87 4.5005
R23762 VOUT+.n84 VOUT+.n81 4.5005
R23763 VOUT+.n88 VOUT+.n81 4.5005
R23764 VOUT+.n89 VOUT+.n33 4.5005
R23765 VOUT+.n89 VOUT+.n35 4.5005
R23766 VOUT+.n89 VOUT+.n88 4.5005
R23767 VOUT+.n179 VOUT+.n92 4.5005
R23768 VOUT+.n180 VOUT+.n179 4.5005
R23769 VOUT+.n180 VOUT+.n29 4.5005
R23770 VOUT+.n181 VOUT+.n28 4.5005
R23771 VOUT+.n181 VOUT+.n180 4.5005
R23772 VOUT+.n185 VOUT+.n184 4.5005
R23773 VOUT+.n184 VOUT+.n20 4.5005
R23774 VOUT+.n23 VOUT+.n20 4.5005
R23775 VOUT+.n187 VOUT+.n20 4.5005
R23776 VOUT+.n189 VOUT+.n20 4.5005
R23777 VOUT+.n188 VOUT+.n23 4.5005
R23778 VOUT+.n188 VOUT+.n187 4.5005
R23779 VOUT+.n189 VOUT+.n188 4.5005
R23780 VOUT+.n1 VOUT+.t16 3.42907
R23781 VOUT+.n1 VOUT+.t14 3.42907
R23782 VOUT+.n5 VOUT+.t15 3.42907
R23783 VOUT+.n5 VOUT+.t4 3.42907
R23784 VOUT+.n8 VOUT+.t17 3.42907
R23785 VOUT+.n8 VOUT+.t18 3.42907
R23786 VOUT+.n86 VOUT+.n34 2.26725
R23787 VOUT+.n82 VOUT+.n32 2.24601
R23788 VOUT+.n183 VOUT+.n182 2.24601
R23789 VOUT+.n25 VOUT+.n22 2.24601
R23790 VOUT+.n178 VOUT+.n177 2.24477
R23791 VOUT+.n31 VOUT+.n26 2.24477
R23792 VOUT+.n89 VOUT+.n34 2.24063
R23793 VOUT+.n181 VOUT+.n27 2.24063
R23794 VOUT+.n188 VOUT+.n24 2.24063
R23795 VOUT+.n81 VOUT+.n80 2.24063
R23796 VOUT+.n179 VOUT+.n90 2.24063
R23797 VOUT+.n91 VOUT+.n29 2.24063
R23798 VOUT+.n186 VOUT+.n185 2.24063
R23799 VOUT+.n185 VOUT+.n21 2.24063
R23800 VOUT+.n87 VOUT+.n85 2.23934
R23801 VOUT+.n87 VOUT+.n83 2.23934
R23802 VOUT+.n6 VOUT+.n4 1.62886
R23803 VOUT+.n10 VOUT+.n9 1.52133
R23804 VOUT+.n17 VOUT+.n2 1.52133
R23805 VOUT+.n79 VOUT+.n78 1.5005
R23806 VOUT+.n77 VOUT+.n36 1.5005
R23807 VOUT+.n76 VOUT+.n75 1.5005
R23808 VOUT+.n74 VOUT+.n39 1.5005
R23809 VOUT+.n73 VOUT+.n72 1.5005
R23810 VOUT+.n71 VOUT+.n40 1.5005
R23811 VOUT+.n70 VOUT+.n69 1.5005
R23812 VOUT+.n68 VOUT+.n43 1.5005
R23813 VOUT+.n18 VOUT+.n17 1.5005
R23814 VOUT+.n16 VOUT+.n0 1.5005
R23815 VOUT+.n15 VOUT+.n14 1.5005
R23816 VOUT+.n13 VOUT+.n3 1.5005
R23817 VOUT+.n12 VOUT+.n11 1.5005
R23818 VOUT+.n65 VOUT+.n60 1.313
R23819 VOUT+.n56 VOUT+.n42 1.313
R23820 VOUT+.n53 VOUT+.n41 1.313
R23821 VOUT+.n50 VOUT+.n38 1.313
R23822 VOUT+.n46 VOUT+.n44 1.313
R23823 VOUT+.n48 VOUT+.n37 1.313
R23824 VOUT+.n180 VOUT+.n30 1.1455
R23825 VOUT+.n96 VOUT+.n95 1.13717
R23826 VOUT+.n97 VOUT+.n93 1.13717
R23827 VOUT+.n176 VOUT+.n175 1.13717
R23828 VOUT+.n94 VOUT+.n31 1.13717
R23829 VOUT+.n95 VOUT+.n28 1.13717
R23830 VOUT+.n93 VOUT+.n92 1.13717
R23831 VOUT+.n177 VOUT+.n176 1.13717
R23832 VOUT+.n67 VOUT+.n44 0.715216
R23833 VOUT+.n66 VOUT+.n65 0.65675
R23834 VOUT+.n70 VOUT+.n42 0.65675
R23835 VOUT+.n72 VOUT+.n41 0.65675
R23836 VOUT+.n76 VOUT+.n38 0.65675
R23837 VOUT+.n78 VOUT+.n37 0.65675
R23838 VOUT+.n96 VOUT+.n30 0.585
R23839 VOUT+.n68 VOUT+.n67 0.564601
R23840 VOUT+.n62 VOUT+.n61 0.563
R23841 VOUT+.n63 VOUT+.n62 0.563
R23842 VOUT+.n64 VOUT+.n63 0.563
R23843 VOUT+.n58 VOUT+.n57 0.563
R23844 VOUT+.n57 VOUT+.n54 0.563
R23845 VOUT+.n54 VOUT+.n51 0.563
R23846 VOUT+.n88 VOUT+.n79 0.5005
R23847 VOUT+.n185 VOUT+.n181 0.338
R23848 VOUT+.n125 VOUT+.n124 0.3295
R23849 VOUT+.n130 VOUT+.n129 0.3295
R23850 VOUT+.n131 VOUT+.n130 0.3295
R23851 VOUT+.n132 VOUT+.n131 0.3295
R23852 VOUT+.n133 VOUT+.n132 0.3295
R23853 VOUT+.n134 VOUT+.n133 0.3295
R23854 VOUT+.n135 VOUT+.n134 0.3295
R23855 VOUT+.n136 VOUT+.n135 0.3295
R23856 VOUT+.n137 VOUT+.n136 0.3295
R23857 VOUT+.n138 VOUT+.n137 0.3295
R23858 VOUT+.n140 VOUT+.n138 0.3295
R23859 VOUT+.n140 VOUT+.n139 0.3295
R23860 VOUT+.n143 VOUT+.n141 0.3295
R23861 VOUT+.n143 VOUT+.n142 0.3295
R23862 VOUT+.n146 VOUT+.n144 0.3295
R23863 VOUT+.n146 VOUT+.n145 0.3295
R23864 VOUT+.n149 VOUT+.n147 0.3295
R23865 VOUT+.n149 VOUT+.n148 0.3295
R23866 VOUT+.n152 VOUT+.n150 0.3295
R23867 VOUT+.n152 VOUT+.n151 0.3295
R23868 VOUT+.n155 VOUT+.n153 0.3295
R23869 VOUT+.n155 VOUT+.n154 0.3295
R23870 VOUT+.n158 VOUT+.n156 0.3295
R23871 VOUT+.n158 VOUT+.n157 0.3295
R23872 VOUT+.n161 VOUT+.n159 0.3295
R23873 VOUT+.n161 VOUT+.n160 0.3295
R23874 VOUT+.n164 VOUT+.n162 0.3295
R23875 VOUT+.n164 VOUT+.n163 0.3295
R23876 VOUT+.n167 VOUT+.n165 0.3295
R23877 VOUT+.n167 VOUT+.n166 0.3295
R23878 VOUT+.n170 VOUT+.n168 0.3295
R23879 VOUT+.n170 VOUT+.n169 0.3295
R23880 VOUT+.n99 VOUT+.n98 0.3295
R23881 VOUT+.n101 VOUT+.n100 0.3295
R23882 VOUT+.n102 VOUT+.n101 0.3295
R23883 VOUT+.n103 VOUT+.n102 0.3295
R23884 VOUT+.n104 VOUT+.n103 0.3295
R23885 VOUT+.n105 VOUT+.n104 0.3295
R23886 VOUT+.n106 VOUT+.n105 0.3295
R23887 VOUT+.n107 VOUT+.n106 0.3295
R23888 VOUT+.n108 VOUT+.n107 0.3295
R23889 VOUT+.n109 VOUT+.n108 0.3295
R23890 VOUT+.n111 VOUT+.n109 0.3295
R23891 VOUT+.n111 VOUT+.n110 0.3295
R23892 VOUT+.n114 VOUT+.n112 0.3295
R23893 VOUT+.n114 VOUT+.n113 0.3295
R23894 VOUT+.n117 VOUT+.n115 0.3295
R23895 VOUT+.n117 VOUT+.n116 0.3295
R23896 VOUT+.n120 VOUT+.n118 0.3295
R23897 VOUT+.n120 VOUT+.n119 0.3295
R23898 VOUT+.n123 VOUT+.n121 0.3295
R23899 VOUT+.n123 VOUT+.n122 0.3295
R23900 VOUT+.n173 VOUT+.n172 0.3295
R23901 VOUT+.n172 VOUT+.n171 0.3295
R23902 VOUT+.n179 VOUT+.n89 0.3205
R23903 VOUT+.n12 VOUT+.n4 0.314966
R23904 VOUT+.n174 VOUT+.n173 0.313833
R23905 VOUT+.n136 VOUT+.n126 0.306
R23906 VOUT+.n135 VOUT+.n127 0.306
R23907 VOUT+.n134 VOUT+.n128 0.306
R23908 VOUT+.n140 VOUT+.n125 0.2825
R23909 VOUT+.n143 VOUT+.n140 0.2825
R23910 VOUT+.n146 VOUT+.n143 0.2825
R23911 VOUT+.n149 VOUT+.n146 0.2825
R23912 VOUT+.n152 VOUT+.n149 0.2825
R23913 VOUT+.n155 VOUT+.n152 0.2825
R23914 VOUT+.n158 VOUT+.n155 0.2825
R23915 VOUT+.n161 VOUT+.n158 0.2825
R23916 VOUT+.n164 VOUT+.n161 0.2825
R23917 VOUT+.n167 VOUT+.n164 0.2825
R23918 VOUT+.n170 VOUT+.n167 0.2825
R23919 VOUT+.n111 VOUT+.n99 0.2825
R23920 VOUT+.n114 VOUT+.n111 0.2825
R23921 VOUT+.n117 VOUT+.n114 0.2825
R23922 VOUT+.n120 VOUT+.n117 0.2825
R23923 VOUT+.n123 VOUT+.n120 0.2825
R23924 VOUT+.n172 VOUT+.n123 0.2825
R23925 VOUT+.n172 VOUT+.n170 0.2825
R23926 VOUT+.n19 VOUT+.n18 0.28175
R23927 VOUT+ VOUT+.n19 0.21925
R23928 VOUT+.n175 VOUT+.n174 0.0898
R23929 VOUT+.n10 VOUT+.n4 0.0891864
R23930 VOUT+.n66 VOUT+.n43 0.0577917
R23931 VOUT+.n70 VOUT+.n43 0.0577917
R23932 VOUT+.n71 VOUT+.n70 0.0577917
R23933 VOUT+.n72 VOUT+.n71 0.0577917
R23934 VOUT+.n72 VOUT+.n39 0.0577917
R23935 VOUT+.n76 VOUT+.n39 0.0577917
R23936 VOUT+.n77 VOUT+.n76 0.0577917
R23937 VOUT+.n78 VOUT+.n77 0.0577917
R23938 VOUT+.n69 VOUT+.n68 0.0577917
R23939 VOUT+.n69 VOUT+.n40 0.0577917
R23940 VOUT+.n73 VOUT+.n40 0.0577917
R23941 VOUT+.n74 VOUT+.n73 0.0577917
R23942 VOUT+.n75 VOUT+.n74 0.0577917
R23943 VOUT+.n75 VOUT+.n36 0.0577917
R23944 VOUT+.n79 VOUT+.n36 0.0577917
R23945 VOUT+ VOUT+.n189 0.0577917
R23946 VOUT+.n67 VOUT+.n66 0.054517
R23947 VOUT+.n187 VOUT+.n25 0.047375
R23948 VOUT+.n182 VOUT+.n23 0.047375
R23949 VOUT+.n180 VOUT+.n31 0.0421667
R23950 VOUT+.n88 VOUT+.n82 0.0421667
R23951 VOUT+.n11 VOUT+.n10 0.0421667
R23952 VOUT+.n11 VOUT+.n3 0.0421667
R23953 VOUT+.n15 VOUT+.n3 0.0421667
R23954 VOUT+.n16 VOUT+.n15 0.0421667
R23955 VOUT+.n17 VOUT+.n16 0.0421667
R23956 VOUT+.n13 VOUT+.n12 0.0421667
R23957 VOUT+.n14 VOUT+.n13 0.0421667
R23958 VOUT+.n14 VOUT+.n0 0.0421667
R23959 VOUT+.n18 VOUT+.n0 0.0421667
R23960 VOUT+.n83 VOUT+.n82 0.0243161
R23961 VOUT+.n85 VOUT+.n33 0.0243161
R23962 VOUT+.n85 VOUT+.n84 0.0243161
R23963 VOUT+.n83 VOUT+.n35 0.0243161
R23964 VOUT+.n177 VOUT+.n27 0.0217373
R23965 VOUT+.n84 VOUT+.n34 0.0217373
R23966 VOUT+.n92 VOUT+.n27 0.0217373
R23967 VOUT+.n184 VOUT+.n24 0.0217373
R23968 VOUT+.n182 VOUT+.n24 0.0217373
R23969 VOUT+.n90 VOUT+.n31 0.0217373
R23970 VOUT+.n92 VOUT+.n91 0.0217373
R23971 VOUT+.n80 VOUT+.n33 0.0217373
R23972 VOUT+.n80 VOUT+.n35 0.0217373
R23973 VOUT+.n90 VOUT+.n28 0.0217373
R23974 VOUT+.n91 VOUT+.n28 0.0217373
R23975 VOUT+.n189 VOUT+.n21 0.0217373
R23976 VOUT+.n187 VOUT+.n186 0.0217373
R23977 VOUT+.n186 VOUT+.n23 0.0217373
R23978 VOUT+.n25 VOUT+.n21 0.0217373
R23979 VOUT+.n97 VOUT+.n96 0.0161667
R23980 VOUT+.n175 VOUT+.n97 0.0161667
R23981 VOUT+.n95 VOUT+.n94 0.0161667
R23982 VOUT+.n95 VOUT+.n93 0.0161667
R23983 VOUT+.n176 VOUT+.n93 0.0161667
R23984 VOUT+.n178 VOUT+.n29 0.0134654
R23985 VOUT+.n181 VOUT+.n26 0.0134654
R23986 VOUT+.n179 VOUT+.n178 0.0134654
R23987 VOUT+.n29 VOUT+.n26 0.0134654
R23988 VOUT+.n86 VOUT+.n81 0.0109778
R23989 VOUT+.n89 VOUT+.n32 0.0109778
R23990 VOUT+.n183 VOUT+.n20 0.0109778
R23991 VOUT+.n188 VOUT+.n22 0.0109778
R23992 VOUT+.n87 VOUT+.n86 0.0109778
R23993 VOUT+.n81 VOUT+.n32 0.0109778
R23994 VOUT+.n185 VOUT+.n183 0.0109778
R23995 VOUT+.n22 VOUT+.n20 0.0109778
R23996 VOUT+.n94 VOUT+.n30 0.00872683
R23997 two_stage_opamp_dummy_magic_24_0.cap_res_Y two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 49.2388
R23998 two_stage_opamp_dummy_magic_24_0.cap_res_Y two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 1.45163
R23999 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 0.1603
R24000 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t44 0.1603
R24001 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 0.1603
R24002 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t64 0.1603
R24003 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 0.1603
R24004 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 0.1603
R24005 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t124 0.1603
R24006 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 0.1603
R24007 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 0.1603
R24008 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 0.1603
R24009 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t129 0.1603
R24010 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 0.1603
R24011 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 0.1603
R24012 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 0.1603
R24013 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 0.1603
R24014 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 0.1603
R24015 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t33 0.1603
R24016 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 0.1603
R24017 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 0.1603
R24018 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 0.1603
R24019 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t111 0.1603
R24020 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 0.1603
R24021 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 0.1603
R24022 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 0.1603
R24023 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 0.1603
R24024 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 0.1603
R24025 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t14 0.1603
R24026 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 0.1603
R24027 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 0.1603
R24028 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t11 0.1603
R24029 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t51 0.1603
R24030 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 0.1603
R24031 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t31 0.1603
R24032 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t65 0.1603
R24033 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 0.1603
R24034 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 0.1603
R24035 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 0.1603
R24036 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 0.1603
R24037 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t117 0.1603
R24038 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t24 0.1603
R24039 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t58 0.1603
R24040 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 0.1603
R24041 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t3 0.1603
R24042 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 0.1603
R24043 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t18 0.1603
R24044 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 0.1603
R24045 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 0.1603
R24046 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 0.1603
R24047 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 0.1603
R24048 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 0.1603
R24049 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 0.1603
R24050 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 0.1603
R24051 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 0.1603
R24052 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 0.1603
R24053 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 0.1603
R24054 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 0.159278
R24055 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 0.159278
R24056 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 0.159278
R24057 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 0.159278
R24058 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 0.159278
R24059 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 0.159278
R24060 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 0.159278
R24061 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 0.159278
R24062 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 0.159278
R24063 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 0.159278
R24064 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 0.159278
R24065 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 0.159278
R24066 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 0.159278
R24067 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 0.159278
R24068 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 0.159278
R24069 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 0.159278
R24070 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 0.159278
R24071 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 0.159278
R24072 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t36 0.159278
R24073 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 0.159278
R24074 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t13 0.159278
R24075 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t47 0.159278
R24076 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t30 0.159278
R24077 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t71 0.159278
R24078 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t105 0.159278
R24079 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t1 0.159278
R24080 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 0.159278
R24081 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t19 0.159278
R24082 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 0.137822
R24083 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 0.1368
R24084 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 0.1368
R24085 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 0.1368
R24086 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 0.1368
R24087 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 0.1368
R24088 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 0.1368
R24089 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 0.1368
R24090 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 0.1368
R24091 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 0.1368
R24092 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 0.1368
R24093 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 0.1368
R24094 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 0.1368
R24095 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 0.1368
R24096 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 0.1368
R24097 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 0.1368
R24098 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 0.1368
R24099 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 0.1368
R24100 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 0.1368
R24101 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 0.1368
R24102 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 0.1368
R24103 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 0.1368
R24104 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 0.1368
R24105 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 0.1368
R24106 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 0.1368
R24107 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 0.1368
R24108 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 0.1368
R24109 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 0.1368
R24110 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 0.1368
R24111 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 0.1368
R24112 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 0.1368
R24113 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 0.1368
R24114 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 0.1368
R24115 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 0.1368
R24116 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 0.114322
R24117 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 0.1133
R24118 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 0.1133
R24119 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 0.1133
R24120 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 0.1133
R24121 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 0.1133
R24122 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 0.1133
R24123 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 0.1133
R24124 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 0.1133
R24125 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 0.1133
R24126 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 0.1133
R24127 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 0.1133
R24128 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 0.1133
R24129 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 0.1133
R24130 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 0.1133
R24131 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 0.1133
R24132 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 0.1133
R24133 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 0.1133
R24134 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 0.1133
R24135 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 0.1133
R24136 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 0.00152174
R24137 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 0.00152174
R24138 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 0.00152174
R24139 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 0.00152174
R24140 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 0.00152174
R24141 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 0.00152174
R24142 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 0.00152174
R24143 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 0.00152174
R24144 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 0.00152174
R24145 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 0.00152174
R24146 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 0.00152174
R24147 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 0.00152174
R24148 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 0.00152174
R24149 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 0.00152174
R24150 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 0.00152174
R24151 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 0.00152174
R24152 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 0.00152174
R24153 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 0.00152174
R24154 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 0.00152174
R24155 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 0.00152174
R24156 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 0.00152174
R24157 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 0.00152174
R24158 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 0.00152174
R24159 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 0.00152174
R24160 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 0.00152174
R24161 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 0.00152174
R24162 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 0.00152174
R24163 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 0.00152174
R24164 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t100 0.00152174
R24165 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 0.00152174
R24166 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 0.00152174
R24167 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 0.00152174
R24168 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 0.00152174
R24169 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 0.00152174
R24170 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 0.00152174
R24171 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 0.00152174
R24172 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n36 0.00152174
R24173 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t3 369.534
R24174 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t8 369.534
R24175 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t5 369.534
R24176 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t17 369.534
R24177 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t14 369.534
R24178 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t13 369.534
R24179 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t15 369.534
R24180 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n1 367.397
R24181 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t7 249.034
R24182 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t19 192.8
R24183 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t22 192.8
R24184 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t11 192.8
R24185 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t10 192.8
R24186 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t16 192.8
R24187 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t9 192.8
R24188 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t20 192.8
R24189 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t12 192.8
R24190 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t18 192.8
R24191 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t6 192.8
R24192 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t21 192.8
R24193 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.n11 176.733
R24194 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 176.733
R24195 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R24196 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R24197 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n6 169.602
R24198 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n18 166.727
R24199 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 166.727
R24200 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n9 166.727
R24201 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n0 142.137
R24202 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.n17 56.2338
R24203 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n14 56.2338
R24204 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n13 56.2338
R24205 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 56.2338
R24206 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R24207 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 56.2338
R24208 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n2 56.2338
R24209 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t1 39.4005
R24210 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t0 39.4005
R24211 bgr_11_0.NFET_GATE_10uA.t2 bgr_11_0.NFET_GATE_10uA.n19 24.0005
R24212 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t4 24.0005
R24213 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n16 4.15675
R24214 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n10 2.8755
R24215 two_stage_opamp_dummy_magic_24_0.Vb2.n23 two_stage_opamp_dummy_magic_24_0.Vb2.t15 746.673
R24216 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.t1 721.625
R24217 two_stage_opamp_dummy_magic_24_0.Vb2.n16 two_stage_opamp_dummy_magic_24_0.Vb2.t12 611.739
R24218 two_stage_opamp_dummy_magic_24_0.Vb2.n12 two_stage_opamp_dummy_magic_24_0.Vb2.t27 611.739
R24219 two_stage_opamp_dummy_magic_24_0.Vb2.n7 two_stage_opamp_dummy_magic_24_0.Vb2.t22 611.739
R24220 two_stage_opamp_dummy_magic_24_0.Vb2.n3 two_stage_opamp_dummy_magic_24_0.Vb2.t19 611.739
R24221 two_stage_opamp_dummy_magic_24_0.Vb2.n2 two_stage_opamp_dummy_magic_24_0.Vb2.t28 563.451
R24222 two_stage_opamp_dummy_magic_24_0.Vb2.n16 two_stage_opamp_dummy_magic_24_0.Vb2.t31 421.75
R24223 two_stage_opamp_dummy_magic_24_0.Vb2.n17 two_stage_opamp_dummy_magic_24_0.Vb2.t25 421.75
R24224 two_stage_opamp_dummy_magic_24_0.Vb2.n18 two_stage_opamp_dummy_magic_24_0.Vb2.t21 421.75
R24225 two_stage_opamp_dummy_magic_24_0.Vb2.n19 two_stage_opamp_dummy_magic_24_0.Vb2.t16 421.75
R24226 two_stage_opamp_dummy_magic_24_0.Vb2.n12 two_stage_opamp_dummy_magic_24_0.Vb2.t23 421.75
R24227 two_stage_opamp_dummy_magic_24_0.Vb2.n13 two_stage_opamp_dummy_magic_24_0.Vb2.t29 421.75
R24228 two_stage_opamp_dummy_magic_24_0.Vb2.n14 two_stage_opamp_dummy_magic_24_0.Vb2.t11 421.75
R24229 two_stage_opamp_dummy_magic_24_0.Vb2.n15 two_stage_opamp_dummy_magic_24_0.Vb2.t13 421.75
R24230 two_stage_opamp_dummy_magic_24_0.Vb2.n7 two_stage_opamp_dummy_magic_24_0.Vb2.t18 421.75
R24231 two_stage_opamp_dummy_magic_24_0.Vb2.n8 two_stage_opamp_dummy_magic_24_0.Vb2.t20 421.75
R24232 two_stage_opamp_dummy_magic_24_0.Vb2.n9 two_stage_opamp_dummy_magic_24_0.Vb2.t17 421.75
R24233 two_stage_opamp_dummy_magic_24_0.Vb2.n10 two_stage_opamp_dummy_magic_24_0.Vb2.t14 421.75
R24234 two_stage_opamp_dummy_magic_24_0.Vb2.n3 two_stage_opamp_dummy_magic_24_0.Vb2.t24 421.75
R24235 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.t30 421.75
R24236 two_stage_opamp_dummy_magic_24_0.Vb2.n5 two_stage_opamp_dummy_magic_24_0.Vb2.t26 421.75
R24237 two_stage_opamp_dummy_magic_24_0.Vb2.n6 two_stage_opamp_dummy_magic_24_0.Vb2.t32 421.75
R24238 two_stage_opamp_dummy_magic_24_0.Vb2.n21 two_stage_opamp_dummy_magic_24_0.Vb2.n11 313.776
R24239 two_stage_opamp_dummy_magic_24_0.Vb2.n21 two_stage_opamp_dummy_magic_24_0.Vb2.n20 313.212
R24240 two_stage_opamp_dummy_magic_24_0.Vb2.n17 two_stage_opamp_dummy_magic_24_0.Vb2.n16 167.094
R24241 two_stage_opamp_dummy_magic_24_0.Vb2.n18 two_stage_opamp_dummy_magic_24_0.Vb2.n17 167.094
R24242 two_stage_opamp_dummy_magic_24_0.Vb2.n19 two_stage_opamp_dummy_magic_24_0.Vb2.n18 167.094
R24243 two_stage_opamp_dummy_magic_24_0.Vb2.n13 two_stage_opamp_dummy_magic_24_0.Vb2.n12 167.094
R24244 two_stage_opamp_dummy_magic_24_0.Vb2.n14 two_stage_opamp_dummy_magic_24_0.Vb2.n13 167.094
R24245 two_stage_opamp_dummy_magic_24_0.Vb2.n15 two_stage_opamp_dummy_magic_24_0.Vb2.n14 167.094
R24246 two_stage_opamp_dummy_magic_24_0.Vb2.n8 two_stage_opamp_dummy_magic_24_0.Vb2.n7 167.094
R24247 two_stage_opamp_dummy_magic_24_0.Vb2.n9 two_stage_opamp_dummy_magic_24_0.Vb2.n8 167.094
R24248 two_stage_opamp_dummy_magic_24_0.Vb2.n10 two_stage_opamp_dummy_magic_24_0.Vb2.n9 167.094
R24249 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.n3 167.094
R24250 two_stage_opamp_dummy_magic_24_0.Vb2.n5 two_stage_opamp_dummy_magic_24_0.Vb2.n4 167.094
R24251 two_stage_opamp_dummy_magic_24_0.Vb2.n6 two_stage_opamp_dummy_magic_24_0.Vb2.n5 167.094
R24252 two_stage_opamp_dummy_magic_24_0.Vb2.n26 two_stage_opamp_dummy_magic_24_0.Vb2.n24 140.546
R24253 two_stage_opamp_dummy_magic_24_0.Vb2.n28 two_stage_opamp_dummy_magic_24_0.Vb2.n27 139.297
R24254 two_stage_opamp_dummy_magic_24_0.Vb2.n26 two_stage_opamp_dummy_magic_24_0.Vb2.n25 139.297
R24255 two_stage_opamp_dummy_magic_24_0.Vb2.n30 two_stage_opamp_dummy_magic_24_0.Vb2.n29 139.297
R24256 two_stage_opamp_dummy_magic_24_0.Vb2.n29 two_stage_opamp_dummy_magic_24_0.Vb2.n23 84.7286
R24257 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.n0 67.013
R24258 two_stage_opamp_dummy_magic_24_0.Vb2.n20 two_stage_opamp_dummy_magic_24_0.Vb2.n19 35.3472
R24259 two_stage_opamp_dummy_magic_24_0.Vb2.n20 two_stage_opamp_dummy_magic_24_0.Vb2.n15 35.3472
R24260 two_stage_opamp_dummy_magic_24_0.Vb2.n11 two_stage_opamp_dummy_magic_24_0.Vb2.n10 35.3472
R24261 two_stage_opamp_dummy_magic_24_0.Vb2.n11 two_stage_opamp_dummy_magic_24_0.Vb2.n6 35.3472
R24262 two_stage_opamp_dummy_magic_24_0.Vb2.n27 two_stage_opamp_dummy_magic_24_0.Vb2.t7 24.0005
R24263 two_stage_opamp_dummy_magic_24_0.Vb2.n27 two_stage_opamp_dummy_magic_24_0.Vb2.t5 24.0005
R24264 two_stage_opamp_dummy_magic_24_0.Vb2.n25 two_stage_opamp_dummy_magic_24_0.Vb2.t6 24.0005
R24265 two_stage_opamp_dummy_magic_24_0.Vb2.n25 two_stage_opamp_dummy_magic_24_0.Vb2.t9 24.0005
R24266 two_stage_opamp_dummy_magic_24_0.Vb2.n24 two_stage_opamp_dummy_magic_24_0.Vb2.t8 24.0005
R24267 two_stage_opamp_dummy_magic_24_0.Vb2.n24 two_stage_opamp_dummy_magic_24_0.Vb2.t3 24.0005
R24268 two_stage_opamp_dummy_magic_24_0.Vb2.n30 two_stage_opamp_dummy_magic_24_0.Vb2.t4 24.0005
R24269 two_stage_opamp_dummy_magic_24_0.Vb2.t10 two_stage_opamp_dummy_magic_24_0.Vb2.n30 24.0005
R24270 two_stage_opamp_dummy_magic_24_0.Vb2.n22 two_stage_opamp_dummy_magic_24_0.Vb2.n21 14.2505
R24271 two_stage_opamp_dummy_magic_24_0.Vb2.n0 two_stage_opamp_dummy_magic_24_0.Vb2.t2 11.2576
R24272 two_stage_opamp_dummy_magic_24_0.Vb2.n0 two_stage_opamp_dummy_magic_24_0.Vb2.t0 11.2576
R24273 two_stage_opamp_dummy_magic_24_0.Vb2.n2 two_stage_opamp_dummy_magic_24_0.Vb2.n1 7.35988
R24274 two_stage_opamp_dummy_magic_24_0.Vb2.n28 two_stage_opamp_dummy_magic_24_0.Vb2.n26 5.8755
R24275 two_stage_opamp_dummy_magic_24_0.Vb2.n23 two_stage_opamp_dummy_magic_24_0.Vb2.n22 4.55362
R24276 two_stage_opamp_dummy_magic_24_0.Vb2.n29 two_stage_opamp_dummy_magic_24_0.Vb2.n28 1.2505
R24277 two_stage_opamp_dummy_magic_24_0.Vb2.n22 two_stage_opamp_dummy_magic_24_0.Vb2.n2 1.14112
R24278 two_stage_opamp_dummy_magic_24_0.Y.n74 two_stage_opamp_dummy_magic_24_0.Y.t52 1172.87
R24279 two_stage_opamp_dummy_magic_24_0.Y.n70 two_stage_opamp_dummy_magic_24_0.Y.t44 1172.87
R24280 two_stage_opamp_dummy_magic_24_0.Y.n74 two_stage_opamp_dummy_magic_24_0.Y.t36 996.134
R24281 two_stage_opamp_dummy_magic_24_0.Y.n75 two_stage_opamp_dummy_magic_24_0.Y.t51 996.134
R24282 two_stage_opamp_dummy_magic_24_0.Y.n76 two_stage_opamp_dummy_magic_24_0.Y.t38 996.134
R24283 two_stage_opamp_dummy_magic_24_0.Y.n77 two_stage_opamp_dummy_magic_24_0.Y.t54 996.134
R24284 two_stage_opamp_dummy_magic_24_0.Y.n73 two_stage_opamp_dummy_magic_24_0.Y.t39 996.134
R24285 two_stage_opamp_dummy_magic_24_0.Y.n72 two_stage_opamp_dummy_magic_24_0.Y.t25 996.134
R24286 two_stage_opamp_dummy_magic_24_0.Y.n71 two_stage_opamp_dummy_magic_24_0.Y.t41 996.134
R24287 two_stage_opamp_dummy_magic_24_0.Y.n70 two_stage_opamp_dummy_magic_24_0.Y.t28 996.134
R24288 two_stage_opamp_dummy_magic_24_0.Y.n46 two_stage_opamp_dummy_magic_24_0.Y.t27 690.867
R24289 two_stage_opamp_dummy_magic_24_0.Y.n39 two_stage_opamp_dummy_magic_24_0.Y.t50 690.867
R24290 two_stage_opamp_dummy_magic_24_0.Y.n55 two_stage_opamp_dummy_magic_24_0.Y.t30 530.201
R24291 two_stage_opamp_dummy_magic_24_0.Y.n48 two_stage_opamp_dummy_magic_24_0.Y.t53 530.201
R24292 two_stage_opamp_dummy_magic_24_0.Y.n46 two_stage_opamp_dummy_magic_24_0.Y.t40 514.134
R24293 two_stage_opamp_dummy_magic_24_0.Y.n39 two_stage_opamp_dummy_magic_24_0.Y.t35 514.134
R24294 two_stage_opamp_dummy_magic_24_0.Y.n40 two_stage_opamp_dummy_magic_24_0.Y.t48 514.134
R24295 two_stage_opamp_dummy_magic_24_0.Y.n41 two_stage_opamp_dummy_magic_24_0.Y.t33 514.134
R24296 two_stage_opamp_dummy_magic_24_0.Y.n42 two_stage_opamp_dummy_magic_24_0.Y.t46 514.134
R24297 two_stage_opamp_dummy_magic_24_0.Y.n43 two_stage_opamp_dummy_magic_24_0.Y.t31 514.134
R24298 two_stage_opamp_dummy_magic_24_0.Y.n44 two_stage_opamp_dummy_magic_24_0.Y.t43 514.134
R24299 two_stage_opamp_dummy_magic_24_0.Y.n45 two_stage_opamp_dummy_magic_24_0.Y.t26 514.134
R24300 two_stage_opamp_dummy_magic_24_0.Y.n55 two_stage_opamp_dummy_magic_24_0.Y.t42 353.467
R24301 two_stage_opamp_dummy_magic_24_0.Y.n54 two_stage_opamp_dummy_magic_24_0.Y.t29 353.467
R24302 two_stage_opamp_dummy_magic_24_0.Y.n53 two_stage_opamp_dummy_magic_24_0.Y.t45 353.467
R24303 two_stage_opamp_dummy_magic_24_0.Y.n52 two_stage_opamp_dummy_magic_24_0.Y.t32 353.467
R24304 two_stage_opamp_dummy_magic_24_0.Y.n51 two_stage_opamp_dummy_magic_24_0.Y.t47 353.467
R24305 two_stage_opamp_dummy_magic_24_0.Y.n50 two_stage_opamp_dummy_magic_24_0.Y.t34 353.467
R24306 two_stage_opamp_dummy_magic_24_0.Y.n49 two_stage_opamp_dummy_magic_24_0.Y.t49 353.467
R24307 two_stage_opamp_dummy_magic_24_0.Y.n48 two_stage_opamp_dummy_magic_24_0.Y.t37 353.467
R24308 two_stage_opamp_dummy_magic_24_0.Y.n73 two_stage_opamp_dummy_magic_24_0.Y.n72 176.733
R24309 two_stage_opamp_dummy_magic_24_0.Y.n72 two_stage_opamp_dummy_magic_24_0.Y.n71 176.733
R24310 two_stage_opamp_dummy_magic_24_0.Y.n71 two_stage_opamp_dummy_magic_24_0.Y.n70 176.733
R24311 two_stage_opamp_dummy_magic_24_0.Y.n75 two_stage_opamp_dummy_magic_24_0.Y.n74 176.733
R24312 two_stage_opamp_dummy_magic_24_0.Y.n76 two_stage_opamp_dummy_magic_24_0.Y.n75 176.733
R24313 two_stage_opamp_dummy_magic_24_0.Y.n77 two_stage_opamp_dummy_magic_24_0.Y.n76 176.733
R24314 two_stage_opamp_dummy_magic_24_0.Y.n54 two_stage_opamp_dummy_magic_24_0.Y.n53 176.733
R24315 two_stage_opamp_dummy_magic_24_0.Y.n53 two_stage_opamp_dummy_magic_24_0.Y.n52 176.733
R24316 two_stage_opamp_dummy_magic_24_0.Y.n52 two_stage_opamp_dummy_magic_24_0.Y.n51 176.733
R24317 two_stage_opamp_dummy_magic_24_0.Y.n51 two_stage_opamp_dummy_magic_24_0.Y.n50 176.733
R24318 two_stage_opamp_dummy_magic_24_0.Y.n50 two_stage_opamp_dummy_magic_24_0.Y.n49 176.733
R24319 two_stage_opamp_dummy_magic_24_0.Y.n49 two_stage_opamp_dummy_magic_24_0.Y.n48 176.733
R24320 two_stage_opamp_dummy_magic_24_0.Y.n45 two_stage_opamp_dummy_magic_24_0.Y.n44 176.733
R24321 two_stage_opamp_dummy_magic_24_0.Y.n44 two_stage_opamp_dummy_magic_24_0.Y.n43 176.733
R24322 two_stage_opamp_dummy_magic_24_0.Y.n43 two_stage_opamp_dummy_magic_24_0.Y.n42 176.733
R24323 two_stage_opamp_dummy_magic_24_0.Y.n42 two_stage_opamp_dummy_magic_24_0.Y.n41 176.733
R24324 two_stage_opamp_dummy_magic_24_0.Y.n41 two_stage_opamp_dummy_magic_24_0.Y.n40 176.733
R24325 two_stage_opamp_dummy_magic_24_0.Y.n40 two_stage_opamp_dummy_magic_24_0.Y.n39 176.733
R24326 two_stage_opamp_dummy_magic_24_0.Y.n57 two_stage_opamp_dummy_magic_24_0.Y.n56 165.472
R24327 two_stage_opamp_dummy_magic_24_0.Y.n57 two_stage_opamp_dummy_magic_24_0.Y.n47 165.472
R24328 two_stage_opamp_dummy_magic_24_0.Y.n80 two_stage_opamp_dummy_magic_24_0.Y.n79 152
R24329 two_stage_opamp_dummy_magic_24_0.Y.n81 two_stage_opamp_dummy_magic_24_0.Y.n80 131.571
R24330 two_stage_opamp_dummy_magic_24_0.Y.n80 two_stage_opamp_dummy_magic_24_0.Y.n78 124.517
R24331 two_stage_opamp_dummy_magic_24_0.Y.n147 two_stage_opamp_dummy_magic_24_0.Y.n57 74.3549
R24332 two_stage_opamp_dummy_magic_24_0.Y.n107 two_stage_opamp_dummy_magic_24_0.Y.n106 66.0338
R24333 two_stage_opamp_dummy_magic_24_0.Y.n98 two_stage_opamp_dummy_magic_24_0.Y.n97 66.0338
R24334 two_stage_opamp_dummy_magic_24_0.Y.n96 two_stage_opamp_dummy_magic_24_0.Y.n95 66.0338
R24335 two_stage_opamp_dummy_magic_24_0.Y.n101 two_stage_opamp_dummy_magic_24_0.Y.n100 66.0338
R24336 two_stage_opamp_dummy_magic_24_0.Y.n104 two_stage_opamp_dummy_magic_24_0.Y.n103 66.0338
R24337 two_stage_opamp_dummy_magic_24_0.Y.n110 two_stage_opamp_dummy_magic_24_0.Y.n109 66.0338
R24338 two_stage_opamp_dummy_magic_24_0.Y.n7 two_stage_opamp_dummy_magic_24_0.Y.n6 49.3505
R24339 two_stage_opamp_dummy_magic_24_0.Y.n11 two_stage_opamp_dummy_magic_24_0.Y.n10 49.3505
R24340 two_stage_opamp_dummy_magic_24_0.Y.n20 two_stage_opamp_dummy_magic_24_0.Y.n19 49.3505
R24341 two_stage_opamp_dummy_magic_24_0.Y.n30 two_stage_opamp_dummy_magic_24_0.Y.n29 49.3505
R24342 two_stage_opamp_dummy_magic_24_0.Y.n26 two_stage_opamp_dummy_magic_24_0.Y.n25 49.3505
R24343 two_stage_opamp_dummy_magic_24_0.Y.n23 two_stage_opamp_dummy_magic_24_0.Y.n22 49.3505
R24344 two_stage_opamp_dummy_magic_24_0.Y.n64 two_stage_opamp_dummy_magic_24_0.Y.t10 41.1625
R24345 two_stage_opamp_dummy_magic_24_0.Y.n78 two_stage_opamp_dummy_magic_24_0.Y.n73 40.1672
R24346 two_stage_opamp_dummy_magic_24_0.Y.n78 two_stage_opamp_dummy_magic_24_0.Y.n77 40.1672
R24347 two_stage_opamp_dummy_magic_24_0.Y.n56 two_stage_opamp_dummy_magic_24_0.Y.n54 40.1672
R24348 two_stage_opamp_dummy_magic_24_0.Y.n56 two_stage_opamp_dummy_magic_24_0.Y.n55 40.1672
R24349 two_stage_opamp_dummy_magic_24_0.Y.n47 two_stage_opamp_dummy_magic_24_0.Y.n45 40.1672
R24350 two_stage_opamp_dummy_magic_24_0.Y.n47 two_stage_opamp_dummy_magic_24_0.Y.n46 40.1672
R24351 two_stage_opamp_dummy_magic_24_0.Y.n82 two_stage_opamp_dummy_magic_24_0.Y.n81 16.3217
R24352 two_stage_opamp_dummy_magic_24_0.Y.n6 two_stage_opamp_dummy_magic_24_0.Y.t14 16.0005
R24353 two_stage_opamp_dummy_magic_24_0.Y.n6 two_stage_opamp_dummy_magic_24_0.Y.t12 16.0005
R24354 two_stage_opamp_dummy_magic_24_0.Y.n10 two_stage_opamp_dummy_magic_24_0.Y.t11 16.0005
R24355 two_stage_opamp_dummy_magic_24_0.Y.n10 two_stage_opamp_dummy_magic_24_0.Y.t16 16.0005
R24356 two_stage_opamp_dummy_magic_24_0.Y.n19 two_stage_opamp_dummy_magic_24_0.Y.t20 16.0005
R24357 two_stage_opamp_dummy_magic_24_0.Y.n19 two_stage_opamp_dummy_magic_24_0.Y.t18 16.0005
R24358 two_stage_opamp_dummy_magic_24_0.Y.n29 two_stage_opamp_dummy_magic_24_0.Y.t17 16.0005
R24359 two_stage_opamp_dummy_magic_24_0.Y.n29 two_stage_opamp_dummy_magic_24_0.Y.t19 16.0005
R24360 two_stage_opamp_dummy_magic_24_0.Y.n25 two_stage_opamp_dummy_magic_24_0.Y.t13 16.0005
R24361 two_stage_opamp_dummy_magic_24_0.Y.n25 two_stage_opamp_dummy_magic_24_0.Y.t22 16.0005
R24362 two_stage_opamp_dummy_magic_24_0.Y.n22 two_stage_opamp_dummy_magic_24_0.Y.t15 16.0005
R24363 two_stage_opamp_dummy_magic_24_0.Y.n22 two_stage_opamp_dummy_magic_24_0.Y.t21 16.0005
R24364 two_stage_opamp_dummy_magic_24_0.Y.n79 two_stage_opamp_dummy_magic_24_0.Y.n69 12.8005
R24365 two_stage_opamp_dummy_magic_24_0.Y.n106 two_stage_opamp_dummy_magic_24_0.Y.t2 11.2576
R24366 two_stage_opamp_dummy_magic_24_0.Y.n106 two_stage_opamp_dummy_magic_24_0.Y.t23 11.2576
R24367 two_stage_opamp_dummy_magic_24_0.Y.n97 two_stage_opamp_dummy_magic_24_0.Y.t24 11.2576
R24368 two_stage_opamp_dummy_magic_24_0.Y.n97 two_stage_opamp_dummy_magic_24_0.Y.t8 11.2576
R24369 two_stage_opamp_dummy_magic_24_0.Y.n95 two_stage_opamp_dummy_magic_24_0.Y.t0 11.2576
R24370 two_stage_opamp_dummy_magic_24_0.Y.n95 two_stage_opamp_dummy_magic_24_0.Y.t3 11.2576
R24371 two_stage_opamp_dummy_magic_24_0.Y.n100 two_stage_opamp_dummy_magic_24_0.Y.t5 11.2576
R24372 two_stage_opamp_dummy_magic_24_0.Y.n100 two_stage_opamp_dummy_magic_24_0.Y.t6 11.2576
R24373 two_stage_opamp_dummy_magic_24_0.Y.n103 two_stage_opamp_dummy_magic_24_0.Y.t7 11.2576
R24374 two_stage_opamp_dummy_magic_24_0.Y.n103 two_stage_opamp_dummy_magic_24_0.Y.t9 11.2576
R24375 two_stage_opamp_dummy_magic_24_0.Y.n109 two_stage_opamp_dummy_magic_24_0.Y.t1 11.2576
R24376 two_stage_opamp_dummy_magic_24_0.Y.n109 two_stage_opamp_dummy_magic_24_0.Y.t4 11.2576
R24377 two_stage_opamp_dummy_magic_24_0.Y.n79 two_stage_opamp_dummy_magic_24_0.Y.n67 9.36264
R24378 two_stage_opamp_dummy_magic_24_0.Y.n69 two_stage_opamp_dummy_magic_24_0.Y.n68 9.3005
R24379 two_stage_opamp_dummy_magic_24_0.Y.n99 two_stage_opamp_dummy_magic_24_0.Y.n98 5.91717
R24380 two_stage_opamp_dummy_magic_24_0.Y.n108 two_stage_opamp_dummy_magic_24_0.Y.n107 5.91717
R24381 two_stage_opamp_dummy_magic_24_0.Y.n21 two_stage_opamp_dummy_magic_24_0.Y.n11 5.6255
R24382 two_stage_opamp_dummy_magic_24_0.Y.n24 two_stage_opamp_dummy_magic_24_0.Y.n7 5.6255
R24383 two_stage_opamp_dummy_magic_24_0.Y.n81 two_stage_opamp_dummy_magic_24_0.Y.n69 5.33141
R24384 two_stage_opamp_dummy_magic_24_0.Y.n99 two_stage_opamp_dummy_magic_24_0.Y.n96 5.29217
R24385 two_stage_opamp_dummy_magic_24_0.Y.n102 two_stage_opamp_dummy_magic_24_0.Y.n101 5.29217
R24386 two_stage_opamp_dummy_magic_24_0.Y.n105 two_stage_opamp_dummy_magic_24_0.Y.n104 5.29217
R24387 two_stage_opamp_dummy_magic_24_0.Y.n110 two_stage_opamp_dummy_magic_24_0.Y.n108 5.29217
R24388 two_stage_opamp_dummy_magic_24_0.Y.n112 two_stage_opamp_dummy_magic_24_0.Y.n86 5.1255
R24389 two_stage_opamp_dummy_magic_24_0.Y.n115 two_stage_opamp_dummy_magic_24_0.Y.n94 5.1255
R24390 two_stage_opamp_dummy_magic_24_0.Y.n21 two_stage_opamp_dummy_magic_24_0.Y.n20 5.063
R24391 two_stage_opamp_dummy_magic_24_0.Y.n30 two_stage_opamp_dummy_magic_24_0.Y.n28 5.063
R24392 two_stage_opamp_dummy_magic_24_0.Y.n27 two_stage_opamp_dummy_magic_24_0.Y.n26 5.063
R24393 two_stage_opamp_dummy_magic_24_0.Y.n24 two_stage_opamp_dummy_magic_24_0.Y.n23 5.063
R24394 two_stage_opamp_dummy_magic_24_0.Y.n35 two_stage_opamp_dummy_magic_24_0.Y.n34 5.063
R24395 two_stage_opamp_dummy_magic_24_0.Y.n12 two_stage_opamp_dummy_magic_24_0.Y.n8 5.063
R24396 two_stage_opamp_dummy_magic_24_0.Y.n112 two_stage_opamp_dummy_magic_24_0.Y.n111 4.5005
R24397 two_stage_opamp_dummy_magic_24_0.Y.n113 two_stage_opamp_dummy_magic_24_0.Y.n89 4.5005
R24398 two_stage_opamp_dummy_magic_24_0.Y.n114 two_stage_opamp_dummy_magic_24_0.Y.n92 4.5005
R24399 two_stage_opamp_dummy_magic_24_0.Y.n116 two_stage_opamp_dummy_magic_24_0.Y.n115 4.5005
R24400 two_stage_opamp_dummy_magic_24_0.Y.n141 two_stage_opamp_dummy_magic_24_0.Y.n140 4.5005
R24401 two_stage_opamp_dummy_magic_24_0.Y.n34 two_stage_opamp_dummy_magic_24_0.Y.n5 4.5005
R24402 two_stage_opamp_dummy_magic_24_0.Y.n33 two_stage_opamp_dummy_magic_24_0.Y.n1 4.5005
R24403 two_stage_opamp_dummy_magic_24_0.Y.n32 two_stage_opamp_dummy_magic_24_0.Y.n31 4.5005
R24404 two_stage_opamp_dummy_magic_24_0.Y.n18 two_stage_opamp_dummy_magic_24_0.Y.n8 4.5005
R24405 two_stage_opamp_dummy_magic_24_0.Y.n148 two_stage_opamp_dummy_magic_24_0.Y.n36 4.5005
R24406 two_stage_opamp_dummy_magic_24_0.Y.n147 two_stage_opamp_dummy_magic_24_0.Y.n146 4.5005
R24407 two_stage_opamp_dummy_magic_24_0.Y.n148 two_stage_opamp_dummy_magic_24_0.Y.n147 4.5005
R24408 two_stage_opamp_dummy_magic_24_0.Y.n83 two_stage_opamp_dummy_magic_24_0.Y.n82 4.5005
R24409 two_stage_opamp_dummy_magic_24_0.Y.n61 two_stage_opamp_dummy_magic_24_0.Y.n60 4.5005
R24410 two_stage_opamp_dummy_magic_24_0.Y.n62 two_stage_opamp_dummy_magic_24_0.Y.n59 2.26187
R24411 two_stage_opamp_dummy_magic_24_0.Y.n138 two_stage_opamp_dummy_magic_24_0.Y.n84 2.26187
R24412 two_stage_opamp_dummy_magic_24_0.Y.n139 two_stage_opamp_dummy_magic_24_0.Y.n138 2.26187
R24413 two_stage_opamp_dummy_magic_24_0.Y.n63 two_stage_opamp_dummy_magic_24_0.Y.n62 2.26187
R24414 two_stage_opamp_dummy_magic_24_0.Y.n142 two_stage_opamp_dummy_magic_24_0.Y.n137 2.24063
R24415 two_stage_opamp_dummy_magic_24_0.Y.n143 two_stage_opamp_dummy_magic_24_0.Y.n84 2.24063
R24416 two_stage_opamp_dummy_magic_24_0.Y.n146 two_stage_opamp_dummy_magic_24_0.Y.n145 2.24063
R24417 two_stage_opamp_dummy_magic_24_0.Y.n58 two_stage_opamp_dummy_magic_24_0.Y.n38 2.24063
R24418 two_stage_opamp_dummy_magic_24_0.Y.n66 two_stage_opamp_dummy_magic_24_0.Y.n59 2.24063
R24419 two_stage_opamp_dummy_magic_24_0.Y.n144 two_stage_opamp_dummy_magic_24_0.Y.n37 2.24063
R24420 two_stage_opamp_dummy_magic_24_0.Y.n65 two_stage_opamp_dummy_magic_24_0.Y.n64 2.24063
R24421 two_stage_opamp_dummy_magic_24_0.Y.n83 two_stage_opamp_dummy_magic_24_0.Y.n67 2.22018
R24422 two_stage_opamp_dummy_magic_24_0.Y.n136 two_stage_opamp_dummy_magic_24_0.Y.n135 1.5005
R24423 two_stage_opamp_dummy_magic_24_0.Y.n134 two_stage_opamp_dummy_magic_24_0.Y.n85 1.5005
R24424 two_stage_opamp_dummy_magic_24_0.Y.n133 two_stage_opamp_dummy_magic_24_0.Y.n132 1.5005
R24425 two_stage_opamp_dummy_magic_24_0.Y.n131 two_stage_opamp_dummy_magic_24_0.Y.n87 1.5005
R24426 two_stage_opamp_dummy_magic_24_0.Y.n130 two_stage_opamp_dummy_magic_24_0.Y.n129 1.5005
R24427 two_stage_opamp_dummy_magic_24_0.Y.n128 two_stage_opamp_dummy_magic_24_0.Y.n88 1.5005
R24428 two_stage_opamp_dummy_magic_24_0.Y.n127 two_stage_opamp_dummy_magic_24_0.Y.n126 1.5005
R24429 two_stage_opamp_dummy_magic_24_0.Y.n125 two_stage_opamp_dummy_magic_24_0.Y.n90 1.5005
R24430 two_stage_opamp_dummy_magic_24_0.Y.n124 two_stage_opamp_dummy_magic_24_0.Y.n123 1.5005
R24431 two_stage_opamp_dummy_magic_24_0.Y.n122 two_stage_opamp_dummy_magic_24_0.Y.n91 1.5005
R24432 two_stage_opamp_dummy_magic_24_0.Y.n121 two_stage_opamp_dummy_magic_24_0.Y.n120 1.5005
R24433 two_stage_opamp_dummy_magic_24_0.Y.n119 two_stage_opamp_dummy_magic_24_0.Y.n93 1.5005
R24434 two_stage_opamp_dummy_magic_24_0.Y.n150 two_stage_opamp_dummy_magic_24_0.Y.n149 1.5005
R24435 two_stage_opamp_dummy_magic_24_0.Y.n151 two_stage_opamp_dummy_magic_24_0.Y.n4 1.5005
R24436 two_stage_opamp_dummy_magic_24_0.Y.n153 two_stage_opamp_dummy_magic_24_0.Y.n152 1.5005
R24437 two_stage_opamp_dummy_magic_24_0.Y.n154 two_stage_opamp_dummy_magic_24_0.Y.n2 1.5005
R24438 two_stage_opamp_dummy_magic_24_0.Y.n156 two_stage_opamp_dummy_magic_24_0.Y.n155 1.5005
R24439 two_stage_opamp_dummy_magic_24_0.Y.n3 two_stage_opamp_dummy_magic_24_0.Y.n0 1.5005
R24440 two_stage_opamp_dummy_magic_24_0.Y.n14 two_stage_opamp_dummy_magic_24_0.Y.n9 1.5005
R24441 two_stage_opamp_dummy_magic_24_0.Y.n16 two_stage_opamp_dummy_magic_24_0.Y.n15 1.5005
R24442 two_stage_opamp_dummy_magic_24_0.Y.n144 two_stage_opamp_dummy_magic_24_0.Y.n143 0.891125
R24443 two_stage_opamp_dummy_magic_24_0.Y.n83 two_stage_opamp_dummy_magic_24_0.Y.n66 0.891125
R24444 two_stage_opamp_dummy_magic_24_0.Y.n13 two_stage_opamp_dummy_magic_24_0.Y.n12 0.887091
R24445 two_stage_opamp_dummy_magic_24_0.Y.n18 two_stage_opamp_dummy_magic_24_0.Y.n17 0.828625
R24446 two_stage_opamp_dummy_magic_24_0.Y.n31 two_stage_opamp_dummy_magic_24_0.Y.n9 0.828625
R24447 two_stage_opamp_dummy_magic_24_0.Y.n156 two_stage_opamp_dummy_magic_24_0.Y.n1 0.828625
R24448 two_stage_opamp_dummy_magic_24_0.Y.n152 two_stage_opamp_dummy_magic_24_0.Y.n5 0.828625
R24449 two_stage_opamp_dummy_magic_24_0.Y.n150 two_stage_opamp_dummy_magic_24_0.Y.n35 0.828625
R24450 two_stage_opamp_dummy_magic_24_0.Y.n116 two_stage_opamp_dummy_magic_24_0.Y.n96 0.792167
R24451 two_stage_opamp_dummy_magic_24_0.Y.n101 two_stage_opamp_dummy_magic_24_0.Y.n92 0.792167
R24452 two_stage_opamp_dummy_magic_24_0.Y.n104 two_stage_opamp_dummy_magic_24_0.Y.n89 0.792167
R24453 two_stage_opamp_dummy_magic_24_0.Y.n111 two_stage_opamp_dummy_magic_24_0.Y.n110 0.792167
R24454 two_stage_opamp_dummy_magic_24_0.Y.n98 two_stage_opamp_dummy_magic_24_0.Y.n94 0.792167
R24455 two_stage_opamp_dummy_magic_24_0.Y.n107 two_stage_opamp_dummy_magic_24_0.Y.n86 0.792167
R24456 two_stage_opamp_dummy_magic_24_0.Y.n113 two_stage_opamp_dummy_magic_24_0.Y.n112 0.6255
R24457 two_stage_opamp_dummy_magic_24_0.Y.n114 two_stage_opamp_dummy_magic_24_0.Y.n113 0.6255
R24458 two_stage_opamp_dummy_magic_24_0.Y.n115 two_stage_opamp_dummy_magic_24_0.Y.n114 0.6255
R24459 two_stage_opamp_dummy_magic_24_0.Y.n102 two_stage_opamp_dummy_magic_24_0.Y.n99 0.6255
R24460 two_stage_opamp_dummy_magic_24_0.Y.n105 two_stage_opamp_dummy_magic_24_0.Y.n102 0.6255
R24461 two_stage_opamp_dummy_magic_24_0.Y.n108 two_stage_opamp_dummy_magic_24_0.Y.n105 0.6255
R24462 two_stage_opamp_dummy_magic_24_0.Y.n15 two_stage_opamp_dummy_magic_24_0.Y.n13 0.564601
R24463 two_stage_opamp_dummy_magic_24_0.Y.n34 two_stage_opamp_dummy_magic_24_0.Y.n33 0.563
R24464 two_stage_opamp_dummy_magic_24_0.Y.n33 two_stage_opamp_dummy_magic_24_0.Y.n32 0.563
R24465 two_stage_opamp_dummy_magic_24_0.Y.n32 two_stage_opamp_dummy_magic_24_0.Y.n8 0.563
R24466 two_stage_opamp_dummy_magic_24_0.Y.n28 two_stage_opamp_dummy_magic_24_0.Y.n21 0.563
R24467 two_stage_opamp_dummy_magic_24_0.Y.n28 two_stage_opamp_dummy_magic_24_0.Y.n27 0.563
R24468 two_stage_opamp_dummy_magic_24_0.Y.n27 two_stage_opamp_dummy_magic_24_0.Y.n24 0.563
R24469 two_stage_opamp_dummy_magic_24_0.Y.n118 two_stage_opamp_dummy_magic_24_0.Y.n94 0.533638
R24470 two_stage_opamp_dummy_magic_24_0.Y.n117 two_stage_opamp_dummy_magic_24_0.Y.n116 0.46925
R24471 two_stage_opamp_dummy_magic_24_0.Y.n122 two_stage_opamp_dummy_magic_24_0.Y.n92 0.46925
R24472 two_stage_opamp_dummy_magic_24_0.Y.n127 two_stage_opamp_dummy_magic_24_0.Y.n89 0.46925
R24473 two_stage_opamp_dummy_magic_24_0.Y.n111 two_stage_opamp_dummy_magic_24_0.Y.n87 0.46925
R24474 two_stage_opamp_dummy_magic_24_0.Y.n135 two_stage_opamp_dummy_magic_24_0.Y.n86 0.46925
R24475 two_stage_opamp_dummy_magic_24_0.Y.n146 two_stage_opamp_dummy_magic_24_0.Y.n83 0.46925
R24476 two_stage_opamp_dummy_magic_24_0.Y.n119 two_stage_opamp_dummy_magic_24_0.Y.n118 0.427973
R24477 two_stage_opamp_dummy_magic_24_0.Y.n149 two_stage_opamp_dummy_magic_24_0.Y.n148 0.422375
R24478 two_stage_opamp_dummy_magic_24_0.Y.n137 two_stage_opamp_dummy_magic_24_0.Y.n136 0.401542
R24479 two_stage_opamp_dummy_magic_24_0.Y.n20 two_stage_opamp_dummy_magic_24_0.Y.n18 0.3755
R24480 two_stage_opamp_dummy_magic_24_0.Y.n31 two_stage_opamp_dummy_magic_24_0.Y.n30 0.3755
R24481 two_stage_opamp_dummy_magic_24_0.Y.n26 two_stage_opamp_dummy_magic_24_0.Y.n1 0.3755
R24482 two_stage_opamp_dummy_magic_24_0.Y.n23 two_stage_opamp_dummy_magic_24_0.Y.n5 0.3755
R24483 two_stage_opamp_dummy_magic_24_0.Y.n12 two_stage_opamp_dummy_magic_24_0.Y.n11 0.3755
R24484 two_stage_opamp_dummy_magic_24_0.Y.n35 two_stage_opamp_dummy_magic_24_0.Y.n7 0.3755
R24485 two_stage_opamp_dummy_magic_24_0.Y.n82 two_stage_opamp_dummy_magic_24_0.Y.n68 0.1255
R24486 two_stage_opamp_dummy_magic_24_0.Y.n68 two_stage_opamp_dummy_magic_24_0.Y.n67 0.0626438
R24487 two_stage_opamp_dummy_magic_24_0.Y.n118 two_stage_opamp_dummy_magic_24_0.Y.n117 0.0587394
R24488 two_stage_opamp_dummy_magic_24_0.Y.n17 two_stage_opamp_dummy_magic_24_0.Y.n16 0.0577917
R24489 two_stage_opamp_dummy_magic_24_0.Y.n16 two_stage_opamp_dummy_magic_24_0.Y.n9 0.0577917
R24490 two_stage_opamp_dummy_magic_24_0.Y.n9 two_stage_opamp_dummy_magic_24_0.Y.n0 0.0577917
R24491 two_stage_opamp_dummy_magic_24_0.Y.n156 two_stage_opamp_dummy_magic_24_0.Y.n2 0.0577917
R24492 two_stage_opamp_dummy_magic_24_0.Y.n152 two_stage_opamp_dummy_magic_24_0.Y.n2 0.0577917
R24493 two_stage_opamp_dummy_magic_24_0.Y.n152 two_stage_opamp_dummy_magic_24_0.Y.n151 0.0577917
R24494 two_stage_opamp_dummy_magic_24_0.Y.n151 two_stage_opamp_dummy_magic_24_0.Y.n150 0.0577917
R24495 two_stage_opamp_dummy_magic_24_0.Y.n15 two_stage_opamp_dummy_magic_24_0.Y.n14 0.0577917
R24496 two_stage_opamp_dummy_magic_24_0.Y.n14 two_stage_opamp_dummy_magic_24_0.Y.n3 0.0577917
R24497 two_stage_opamp_dummy_magic_24_0.Y.n155 two_stage_opamp_dummy_magic_24_0.Y.n3 0.0577917
R24498 two_stage_opamp_dummy_magic_24_0.Y.n155 two_stage_opamp_dummy_magic_24_0.Y.n154 0.0577917
R24499 two_stage_opamp_dummy_magic_24_0.Y.n154 two_stage_opamp_dummy_magic_24_0.Y.n153 0.0577917
R24500 two_stage_opamp_dummy_magic_24_0.Y.n153 two_stage_opamp_dummy_magic_24_0.Y.n4 0.0577917
R24501 two_stage_opamp_dummy_magic_24_0.Y.n149 two_stage_opamp_dummy_magic_24_0.Y.n4 0.0577917
R24502 two_stage_opamp_dummy_magic_24_0.Y.n17 two_stage_opamp_dummy_magic_24_0.Y.n13 0.054517
R24503 two_stage_opamp_dummy_magic_24_0.Y.n117 two_stage_opamp_dummy_magic_24_0.Y.n93 0.0421667
R24504 two_stage_opamp_dummy_magic_24_0.Y.n121 two_stage_opamp_dummy_magic_24_0.Y.n93 0.0421667
R24505 two_stage_opamp_dummy_magic_24_0.Y.n122 two_stage_opamp_dummy_magic_24_0.Y.n121 0.0421667
R24506 two_stage_opamp_dummy_magic_24_0.Y.n123 two_stage_opamp_dummy_magic_24_0.Y.n122 0.0421667
R24507 two_stage_opamp_dummy_magic_24_0.Y.n123 two_stage_opamp_dummy_magic_24_0.Y.n90 0.0421667
R24508 two_stage_opamp_dummy_magic_24_0.Y.n127 two_stage_opamp_dummy_magic_24_0.Y.n90 0.0421667
R24509 two_stage_opamp_dummy_magic_24_0.Y.n128 two_stage_opamp_dummy_magic_24_0.Y.n127 0.0421667
R24510 two_stage_opamp_dummy_magic_24_0.Y.n129 two_stage_opamp_dummy_magic_24_0.Y.n128 0.0421667
R24511 two_stage_opamp_dummy_magic_24_0.Y.n129 two_stage_opamp_dummy_magic_24_0.Y.n87 0.0421667
R24512 two_stage_opamp_dummy_magic_24_0.Y.n133 two_stage_opamp_dummy_magic_24_0.Y.n87 0.0421667
R24513 two_stage_opamp_dummy_magic_24_0.Y.n134 two_stage_opamp_dummy_magic_24_0.Y.n133 0.0421667
R24514 two_stage_opamp_dummy_magic_24_0.Y.n135 two_stage_opamp_dummy_magic_24_0.Y.n134 0.0421667
R24515 two_stage_opamp_dummy_magic_24_0.Y.n120 two_stage_opamp_dummy_magic_24_0.Y.n119 0.0421667
R24516 two_stage_opamp_dummy_magic_24_0.Y.n120 two_stage_opamp_dummy_magic_24_0.Y.n91 0.0421667
R24517 two_stage_opamp_dummy_magic_24_0.Y.n124 two_stage_opamp_dummy_magic_24_0.Y.n91 0.0421667
R24518 two_stage_opamp_dummy_magic_24_0.Y.n125 two_stage_opamp_dummy_magic_24_0.Y.n124 0.0421667
R24519 two_stage_opamp_dummy_magic_24_0.Y.n126 two_stage_opamp_dummy_magic_24_0.Y.n125 0.0421667
R24520 two_stage_opamp_dummy_magic_24_0.Y.n126 two_stage_opamp_dummy_magic_24_0.Y.n88 0.0421667
R24521 two_stage_opamp_dummy_magic_24_0.Y.n130 two_stage_opamp_dummy_magic_24_0.Y.n88 0.0421667
R24522 two_stage_opamp_dummy_magic_24_0.Y.n131 two_stage_opamp_dummy_magic_24_0.Y.n130 0.0421667
R24523 two_stage_opamp_dummy_magic_24_0.Y.n132 two_stage_opamp_dummy_magic_24_0.Y.n131 0.0421667
R24524 two_stage_opamp_dummy_magic_24_0.Y.n132 two_stage_opamp_dummy_magic_24_0.Y.n85 0.0421667
R24525 two_stage_opamp_dummy_magic_24_0.Y.n136 two_stage_opamp_dummy_magic_24_0.Y.n85 0.0421667
R24526 two_stage_opamp_dummy_magic_24_0.Y.n146 two_stage_opamp_dummy_magic_24_0.Y.n58 0.0421667
R24527 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.Y.n0 0.0369583
R24528 two_stage_opamp_dummy_magic_24_0.Y.n142 two_stage_opamp_dummy_magic_24_0.Y.n141 0.0217373
R24529 two_stage_opamp_dummy_magic_24_0.Y.n145 two_stage_opamp_dummy_magic_24_0.Y.n144 0.0217373
R24530 two_stage_opamp_dummy_magic_24_0.Y.n147 two_stage_opamp_dummy_magic_24_0.Y.n38 0.0217373
R24531 two_stage_opamp_dummy_magic_24_0.Y.n140 two_stage_opamp_dummy_magic_24_0.Y.n84 0.0217373
R24532 two_stage_opamp_dummy_magic_24_0.Y.n143 two_stage_opamp_dummy_magic_24_0.Y.n142 0.0217373
R24533 two_stage_opamp_dummy_magic_24_0.Y.n145 two_stage_opamp_dummy_magic_24_0.Y.n36 0.0217373
R24534 two_stage_opamp_dummy_magic_24_0.Y.n38 two_stage_opamp_dummy_magic_24_0.Y.n36 0.0217373
R24535 two_stage_opamp_dummy_magic_24_0.Y.n61 two_stage_opamp_dummy_magic_24_0.Y.n59 0.0217373
R24536 two_stage_opamp_dummy_magic_24_0.Y.n62 two_stage_opamp_dummy_magic_24_0.Y.n60 0.0217373
R24537 two_stage_opamp_dummy_magic_24_0.Y.n140 two_stage_opamp_dummy_magic_24_0.Y.n139 0.0217373
R24538 two_stage_opamp_dummy_magic_24_0.Y.n141 two_stage_opamp_dummy_magic_24_0.Y.n138 0.0217373
R24539 two_stage_opamp_dummy_magic_24_0.Y.n139 two_stage_opamp_dummy_magic_24_0.Y.n137 0.0217373
R24540 two_stage_opamp_dummy_magic_24_0.Y.n148 two_stage_opamp_dummy_magic_24_0.Y.n37 0.0217373
R24541 two_stage_opamp_dummy_magic_24_0.Y.n65 two_stage_opamp_dummy_magic_24_0.Y.n60 0.0217373
R24542 two_stage_opamp_dummy_magic_24_0.Y.n58 two_stage_opamp_dummy_magic_24_0.Y.n37 0.0217373
R24543 two_stage_opamp_dummy_magic_24_0.Y.n63 two_stage_opamp_dummy_magic_24_0.Y.n61 0.0217373
R24544 two_stage_opamp_dummy_magic_24_0.Y.n64 two_stage_opamp_dummy_magic_24_0.Y.n63 0.0217373
R24545 two_stage_opamp_dummy_magic_24_0.Y.n66 two_stage_opamp_dummy_magic_24_0.Y.n65 0.0217373
R24546 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.Y.n156 0.0213333
R24547 two_stage_opamp_dummy_magic_24_0.VD2.n15 two_stage_opamp_dummy_magic_24_0.VD2.n14 49.3505
R24548 two_stage_opamp_dummy_magic_24_0.VD2.n18 two_stage_opamp_dummy_magic_24_0.VD2.n17 49.3505
R24549 two_stage_opamp_dummy_magic_24_0.VD2.n4 two_stage_opamp_dummy_magic_24_0.VD2.n3 49.3505
R24550 two_stage_opamp_dummy_magic_24_0.VD2.n7 two_stage_opamp_dummy_magic_24_0.VD2.n6 49.3505
R24551 two_stage_opamp_dummy_magic_24_0.VD2.n39 two_stage_opamp_dummy_magic_24_0.VD2.n38 49.3505
R24552 two_stage_opamp_dummy_magic_24_0.VD2.n32 two_stage_opamp_dummy_magic_24_0.VD2.n31 49.3505
R24553 two_stage_opamp_dummy_magic_24_0.VD2.n12 two_stage_opamp_dummy_magic_24_0.VD2.n11 49.3505
R24554 two_stage_opamp_dummy_magic_24_0.VD2.n25 two_stage_opamp_dummy_magic_24_0.VD2.n24 49.3505
R24555 two_stage_opamp_dummy_magic_24_0.VD2.n9 two_stage_opamp_dummy_magic_24_0.VD2.n8 49.3505
R24556 two_stage_opamp_dummy_magic_24_0.VD2.n43 two_stage_opamp_dummy_magic_24_0.VD2.n42 49.3505
R24557 two_stage_opamp_dummy_magic_24_0.VD2.n28 two_stage_opamp_dummy_magic_24_0.VD2.n27 49.3505
R24558 two_stage_opamp_dummy_magic_24_0.VD2.n14 two_stage_opamp_dummy_magic_24_0.VD2.t9 16.0005
R24559 two_stage_opamp_dummy_magic_24_0.VD2.n14 two_stage_opamp_dummy_magic_24_0.VD2.t4 16.0005
R24560 two_stage_opamp_dummy_magic_24_0.VD2.n17 two_stage_opamp_dummy_magic_24_0.VD2.t0 16.0005
R24561 two_stage_opamp_dummy_magic_24_0.VD2.n17 two_stage_opamp_dummy_magic_24_0.VD2.t8 16.0005
R24562 two_stage_opamp_dummy_magic_24_0.VD2.n3 two_stage_opamp_dummy_magic_24_0.VD2.t3 16.0005
R24563 two_stage_opamp_dummy_magic_24_0.VD2.n3 two_stage_opamp_dummy_magic_24_0.VD2.t5 16.0005
R24564 two_stage_opamp_dummy_magic_24_0.VD2.n6 two_stage_opamp_dummy_magic_24_0.VD2.t1 16.0005
R24565 two_stage_opamp_dummy_magic_24_0.VD2.n6 two_stage_opamp_dummy_magic_24_0.VD2.t10 16.0005
R24566 two_stage_opamp_dummy_magic_24_0.VD2.n38 two_stage_opamp_dummy_magic_24_0.VD2.t21 16.0005
R24567 two_stage_opamp_dummy_magic_24_0.VD2.n38 two_stage_opamp_dummy_magic_24_0.VD2.t6 16.0005
R24568 two_stage_opamp_dummy_magic_24_0.VD2.n31 two_stage_opamp_dummy_magic_24_0.VD2.t13 16.0005
R24569 two_stage_opamp_dummy_magic_24_0.VD2.n31 two_stage_opamp_dummy_magic_24_0.VD2.t19 16.0005
R24570 two_stage_opamp_dummy_magic_24_0.VD2.n11 two_stage_opamp_dummy_magic_24_0.VD2.t16 16.0005
R24571 two_stage_opamp_dummy_magic_24_0.VD2.n11 two_stage_opamp_dummy_magic_24_0.VD2.t11 16.0005
R24572 two_stage_opamp_dummy_magic_24_0.VD2.n24 two_stage_opamp_dummy_magic_24_0.VD2.t14 16.0005
R24573 two_stage_opamp_dummy_magic_24_0.VD2.n24 two_stage_opamp_dummy_magic_24_0.VD2.t17 16.0005
R24574 two_stage_opamp_dummy_magic_24_0.VD2.n8 two_stage_opamp_dummy_magic_24_0.VD2.t12 16.0005
R24575 two_stage_opamp_dummy_magic_24_0.VD2.n8 two_stage_opamp_dummy_magic_24_0.VD2.t18 16.0005
R24576 two_stage_opamp_dummy_magic_24_0.VD2.n42 two_stage_opamp_dummy_magic_24_0.VD2.t2 16.0005
R24577 two_stage_opamp_dummy_magic_24_0.VD2.n42 two_stage_opamp_dummy_magic_24_0.VD2.t7 16.0005
R24578 two_stage_opamp_dummy_magic_24_0.VD2.n27 two_stage_opamp_dummy_magic_24_0.VD2.t15 16.0005
R24579 two_stage_opamp_dummy_magic_24_0.VD2.n27 two_stage_opamp_dummy_magic_24_0.VD2.t20 16.0005
R24580 two_stage_opamp_dummy_magic_24_0.VD2.n23 two_stage_opamp_dummy_magic_24_0.VD2.n13 5.8755
R24581 two_stage_opamp_dummy_magic_24_0.VD2.n36 two_stage_opamp_dummy_magic_24_0.VD2.n35 5.8755
R24582 two_stage_opamp_dummy_magic_24_0.VD2.n21 two_stage_opamp_dummy_magic_24_0.VD2.n20 5.8755
R24583 two_stage_opamp_dummy_magic_24_0.VD2.n33 two_stage_opamp_dummy_magic_24_0.VD2.n2 5.8755
R24584 two_stage_opamp_dummy_magic_24_0.VD2.n30 two_stage_opamp_dummy_magic_24_0.VD2.n9 5.6255
R24585 two_stage_opamp_dummy_magic_24_0.VD2.n26 two_stage_opamp_dummy_magic_24_0.VD2.n12 5.6255
R24586 two_stage_opamp_dummy_magic_24_0.VD2.n40 two_stage_opamp_dummy_magic_24_0.VD2.n7 5.438
R24587 two_stage_opamp_dummy_magic_24_0.VD2.n16 two_stage_opamp_dummy_magic_24_0.VD2.n15 5.438
R24588 two_stage_opamp_dummy_magic_24_0.VD2.n36 two_stage_opamp_dummy_magic_24_0.VD2.n7 5.31821
R24589 two_stage_opamp_dummy_magic_24_0.VD2.n20 two_stage_opamp_dummy_magic_24_0.VD2.n15 5.31821
R24590 two_stage_opamp_dummy_magic_24_0.VD2.n19 two_stage_opamp_dummy_magic_24_0.VD2.n18 5.08383
R24591 two_stage_opamp_dummy_magic_24_0.VD2.n4 two_stage_opamp_dummy_magic_24_0.VD2.n1 5.08383
R24592 two_stage_opamp_dummy_magic_24_0.VD2.n39 two_stage_opamp_dummy_magic_24_0.VD2.n37 5.08383
R24593 two_stage_opamp_dummy_magic_24_0.VD2.n44 two_stage_opamp_dummy_magic_24_0.VD2.n43 5.08383
R24594 two_stage_opamp_dummy_magic_24_0.VD2.n29 two_stage_opamp_dummy_magic_24_0.VD2.n28 5.063
R24595 two_stage_opamp_dummy_magic_24_0.VD2.n26 two_stage_opamp_dummy_magic_24_0.VD2.n25 5.063
R24596 two_stage_opamp_dummy_magic_24_0.VD2.n35 two_stage_opamp_dummy_magic_24_0.VD2.n34 5.063
R24597 two_stage_opamp_dummy_magic_24_0.VD2.n22 two_stage_opamp_dummy_magic_24_0.VD2.n21 5.063
R24598 two_stage_opamp_dummy_magic_24_0.VD2.n32 two_stage_opamp_dummy_magic_24_0.VD2.n30 5.063
R24599 two_stage_opamp_dummy_magic_24_0.VD2.n18 two_stage_opamp_dummy_magic_24_0.VD2.n16 4.8755
R24600 two_stage_opamp_dummy_magic_24_0.VD2.n5 two_stage_opamp_dummy_magic_24_0.VD2.n4 4.8755
R24601 two_stage_opamp_dummy_magic_24_0.VD2.n40 two_stage_opamp_dummy_magic_24_0.VD2.n39 4.8755
R24602 two_stage_opamp_dummy_magic_24_0.VD2.n43 two_stage_opamp_dummy_magic_24_0.VD2.n41 4.8755
R24603 two_stage_opamp_dummy_magic_24_0.VD2 two_stage_opamp_dummy_magic_24_0.VD2.n45 4.60467
R24604 two_stage_opamp_dummy_magic_24_0.VD2.n23 two_stage_opamp_dummy_magic_24_0.VD2.n22 4.5005
R24605 two_stage_opamp_dummy_magic_24_0.VD2.n34 two_stage_opamp_dummy_magic_24_0.VD2.n33 4.5005
R24606 two_stage_opamp_dummy_magic_24_0.VD2.n10 two_stage_opamp_dummy_magic_24_0.VD2.n0 4.5005
R24607 two_stage_opamp_dummy_magic_24_0.VD2 two_stage_opamp_dummy_magic_24_0.VD2.n0 1.27133
R24608 two_stage_opamp_dummy_magic_24_0.VD2.n34 two_stage_opamp_dummy_magic_24_0.VD2.n10 0.563
R24609 two_stage_opamp_dummy_magic_24_0.VD2.n22 two_stage_opamp_dummy_magic_24_0.VD2.n10 0.563
R24610 two_stage_opamp_dummy_magic_24_0.VD2.n29 two_stage_opamp_dummy_magic_24_0.VD2.n26 0.563
R24611 two_stage_opamp_dummy_magic_24_0.VD2.n30 two_stage_opamp_dummy_magic_24_0.VD2.n29 0.563
R24612 two_stage_opamp_dummy_magic_24_0.VD2.n41 two_stage_opamp_dummy_magic_24_0.VD2.n40 0.563
R24613 two_stage_opamp_dummy_magic_24_0.VD2.n41 two_stage_opamp_dummy_magic_24_0.VD2.n5 0.563
R24614 two_stage_opamp_dummy_magic_24_0.VD2.n16 two_stage_opamp_dummy_magic_24_0.VD2.n5 0.563
R24615 two_stage_opamp_dummy_magic_24_0.VD2.n25 two_stage_opamp_dummy_magic_24_0.VD2.n23 0.3755
R24616 two_stage_opamp_dummy_magic_24_0.VD2.n35 two_stage_opamp_dummy_magic_24_0.VD2.n9 0.3755
R24617 two_stage_opamp_dummy_magic_24_0.VD2.n21 two_stage_opamp_dummy_magic_24_0.VD2.n12 0.3755
R24618 two_stage_opamp_dummy_magic_24_0.VD2.n33 two_stage_opamp_dummy_magic_24_0.VD2.n32 0.3755
R24619 two_stage_opamp_dummy_magic_24_0.VD2.n28 two_stage_opamp_dummy_magic_24_0.VD2.n0 0.3755
R24620 two_stage_opamp_dummy_magic_24_0.VD2.n45 two_stage_opamp_dummy_magic_24_0.VD2.n44 0.234875
R24621 two_stage_opamp_dummy_magic_24_0.VD2.n44 two_stage_opamp_dummy_magic_24_0.VD2.n2 0.234875
R24622 two_stage_opamp_dummy_magic_24_0.VD2.n37 two_stage_opamp_dummy_magic_24_0.VD2.n2 0.234875
R24623 two_stage_opamp_dummy_magic_24_0.VD2.n37 two_stage_opamp_dummy_magic_24_0.VD2.n36 0.234875
R24624 two_stage_opamp_dummy_magic_24_0.VD2.n20 two_stage_opamp_dummy_magic_24_0.VD2.n19 0.234875
R24625 two_stage_opamp_dummy_magic_24_0.VD2.n19 two_stage_opamp_dummy_magic_24_0.VD2.n13 0.234875
R24626 two_stage_opamp_dummy_magic_24_0.VD2.n13 two_stage_opamp_dummy_magic_24_0.VD2.n1 0.234875
R24627 two_stage_opamp_dummy_magic_24_0.VD2.n45 two_stage_opamp_dummy_magic_24_0.VD2.n1 0.234875
R24628 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t9 354.854
R24629 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t22 346.8
R24630 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n11 339.522
R24631 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n6 339.522
R24632 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 335.022
R24633 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t24 184.097
R24634 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t7 184.097
R24635 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t20 184.097
R24636 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t11 184.097
R24637 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n10 166.05
R24638 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n7 166.05
R24639 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t0 106.556
R24640 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.n0 53.3384
R24641 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t4 39.4005
R24642 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t5 39.4005
R24643 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t6 39.4005
R24644 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t1 39.4005
R24645 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t3 39.4005
R24646 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t2 39.4005
R24647 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t30 4.8295
R24648 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t15 4.8295
R24649 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t32 4.8295
R24650 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t25 4.8295
R24651 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t28 4.8295
R24652 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t14 4.8295
R24653 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t17 4.8295
R24654 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t8 4.8295
R24655 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t27 4.8295
R24656 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t19 4.5005
R24657 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t26 4.5005
R24658 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t29 4.5005
R24659 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t31 4.5005
R24660 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R24661 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t23 4.5005
R24662 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t10 4.5005
R24663 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t13 4.5005
R24664 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t16 4.5005
R24665 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t21 4.5005
R24666 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t12 4.5005
R24667 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n9 4.5005
R24668 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n2 2.2095
R24669 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n4 2.0005
R24670 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n3 1.813
R24671 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n5 1.813
R24672 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.8935
R24673 bgr_11_0.V_TOP.n0 bgr_11_0.V_TOP.t34 369.534
R24674 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 339.961
R24675 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 339.272
R24676 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 339.272
R24677 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 339.272
R24678 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 339.272
R24679 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 334.772
R24680 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 224.934
R24681 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 224.934
R24682 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 224.934
R24683 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 224.934
R24684 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 224.934
R24685 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 224.934
R24686 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 224.934
R24687 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.n0 224.934
R24688 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 224.934
R24689 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 224.934
R24690 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 224.934
R24691 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 224.934
R24692 bgr_11_0.V_TOP bgr_11_0.V_TOP.t15 214.222
R24693 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 164.113
R24694 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t31 144.601
R24695 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t40 144.601
R24696 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t47 144.601
R24697 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t23 144.601
R24698 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.t21 144.601
R24699 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t33 144.601
R24700 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.t41 144.601
R24701 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t49 144.601
R24702 bgr_11_0.V_TOP.n0 bgr_11_0.V_TOP.t36 144.601
R24703 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t19 144.601
R24704 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t44 144.601
R24705 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t37 144.601
R24706 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t25 144.601
R24707 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t27 144.601
R24708 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t13 108.424
R24709 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t12 95.9779
R24710 bgr_11_0.V_TOP bgr_11_0.V_TOP.n39 69.6227
R24711 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 69.6227
R24712 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n5 69.6227
R24713 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t8 39.4005
R24714 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t1 39.4005
R24715 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t3 39.4005
R24716 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t2 39.4005
R24717 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t7 39.4005
R24718 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t11 39.4005
R24719 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t10 39.4005
R24720 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t6 39.4005
R24721 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t5 39.4005
R24722 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t0 39.4005
R24723 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t4 39.4005
R24724 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t9 39.4005
R24725 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 37.1479
R24726 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n17 26.8996
R24727 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 9.2505
R24728 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.n29 5.188
R24729 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.t26 4.8295
R24730 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t46 4.8295
R24731 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t35 4.8295
R24732 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t18 4.8295
R24733 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t24 4.8295
R24734 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t45 4.8295
R24735 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t48 4.8295
R24736 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t38 4.8295
R24737 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t42 4.8295
R24738 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.t32 4.5005
R24739 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t20 4.5005
R24740 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t39 4.5005
R24741 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t30 4.5005
R24742 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t29 4.5005
R24743 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t17 4.5005
R24744 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t16 4.5005
R24745 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t43 4.5005
R24746 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t22 4.5005
R24747 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t28 4.5005
R24748 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t14 4.5005
R24749 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R24750 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 2.1255
R24751 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 2.1255
R24752 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 2.1255
R24753 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 0.3295
R24754 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R24755 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R24756 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R24757 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.3295
R24758 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R24759 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n7 0.2825
R24760 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R24761 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R24762 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.n13 0.2825
R24763 VOUT-.n190 VOUT-.t17 110.191
R24764 VOUT-.n39 VOUT-.n38 34.9935
R24765 VOUT-.n28 VOUT-.n27 34.9935
R24766 VOUT-.n30 VOUT-.n29 34.9935
R24767 VOUT-.n33 VOUT-.n32 34.9935
R24768 VOUT-.n36 VOUT-.n35 34.9935
R24769 VOUT-.n42 VOUT-.n41 34.9935
R24770 VOUT-.n177 VOUT-.n176 9.73997
R24771 VOUT-.n173 VOUT-.n172 9.73997
R24772 VOUT-.n180 VOUT-.n179 9.73997
R24773 VOUT-.n178 VOUT-.n173 6.64633
R24774 VOUT-.n178 VOUT-.n177 6.64633
R24775 VOUT-.n38 VOUT-.t2 6.56717
R24776 VOUT-.n38 VOUT-.t12 6.56717
R24777 VOUT-.n27 VOUT-.t13 6.56717
R24778 VOUT-.n27 VOUT-.t4 6.56717
R24779 VOUT-.n29 VOUT-.t10 6.56717
R24780 VOUT-.n29 VOUT-.t3 6.56717
R24781 VOUT-.n32 VOUT-.t16 6.56717
R24782 VOUT-.n32 VOUT-.t11 6.56717
R24783 VOUT-.n35 VOUT-.t18 6.56717
R24784 VOUT-.n35 VOUT-.t9 6.56717
R24785 VOUT-.n41 VOUT-.t1 6.56717
R24786 VOUT-.n41 VOUT-.t8 6.56717
R24787 VOUT-.n31 VOUT-.n28 6.3755
R24788 VOUT-.n40 VOUT-.n39 6.3755
R24789 VOUT-.n180 VOUT-.n178 6.02133
R24790 VOUT-.n31 VOUT-.n30 5.813
R24791 VOUT-.n34 VOUT-.n33 5.813
R24792 VOUT-.n37 VOUT-.n36 5.813
R24793 VOUT-.n42 VOUT-.n40 5.813
R24794 VOUT-.n46 VOUT-.n26 5.063
R24795 VOUT-.n43 VOUT-.n19 5.063
R24796 VOUT-.n97 VOUT-.t102 4.8295
R24797 VOUT-.n102 VOUT-.t72 4.8295
R24798 VOUT-.n101 VOUT-.t106 4.8295
R24799 VOUT-.n100 VOUT-.t139 4.8295
R24800 VOUT-.n99 VOUT-.t66 4.8295
R24801 VOUT-.n114 VOUT-.t99 4.8295
R24802 VOUT-.n115 VOUT-.t143 4.8295
R24803 VOUT-.n117 VOUT-.t70 4.8295
R24804 VOUT-.n118 VOUT-.t60 4.8295
R24805 VOUT-.n120 VOUT-.t27 4.8295
R24806 VOUT-.n121 VOUT-.t150 4.8295
R24807 VOUT-.n123 VOUT-.t69 4.8295
R24808 VOUT-.n124 VOUT-.t51 4.8295
R24809 VOUT-.n126 VOUT-.t23 4.8295
R24810 VOUT-.n127 VOUT-.t146 4.8295
R24811 VOUT-.n129 VOUT-.t121 4.8295
R24812 VOUT-.n130 VOUT-.t108 4.8295
R24813 VOUT-.n132 VOUT-.t156 4.8295
R24814 VOUT-.n133 VOUT-.t140 4.8295
R24815 VOUT-.n135 VOUT-.t114 4.8295
R24816 VOUT-.n136 VOUT-.t103 4.8295
R24817 VOUT-.n138 VOUT-.t77 4.8295
R24818 VOUT-.n139 VOUT-.t67 4.8295
R24819 VOUT-.n141 VOUT-.t40 4.8295
R24820 VOUT-.n142 VOUT-.t20 4.8295
R24821 VOUT-.n71 VOUT-.t87 4.8295
R24822 VOUT-.n73 VOUT-.t115 4.8295
R24823 VOUT-.n85 VOUT-.t110 4.8295
R24824 VOUT-.n86 VOUT-.t80 4.8295
R24825 VOUT-.n88 VOUT-.t28 4.8295
R24826 VOUT-.n89 VOUT-.t149 4.8295
R24827 VOUT-.n91 VOUT-.t131 4.8295
R24828 VOUT-.n92 VOUT-.t111 4.8295
R24829 VOUT-.n94 VOUT-.t33 4.8295
R24830 VOUT-.n95 VOUT-.t152 4.8295
R24831 VOUT-.n144 VOUT-.t74 4.8295
R24832 VOUT-.n103 VOUT-.t42 4.8154
R24833 VOUT-.n104 VOUT-.t155 4.8154
R24834 VOUT-.n105 VOUT-.t35 4.8154
R24835 VOUT-.n106 VOUT-.t75 4.8154
R24836 VOUT-.n103 VOUT-.t49 4.806
R24837 VOUT-.n104 VOUT-.t22 4.806
R24838 VOUT-.n105 VOUT-.t43 4.806
R24839 VOUT-.n106 VOUT-.t79 4.806
R24840 VOUT-.n107 VOUT-.t56 4.806
R24841 VOUT-.n107 VOUT-.t62 4.806
R24842 VOUT-.n108 VOUT-.t98 4.806
R24843 VOUT-.n109 VOUT-.t127 4.806
R24844 VOUT-.n110 VOUT-.t30 4.806
R24845 VOUT-.n111 VOUT-.t147 4.806
R24846 VOUT-.n112 VOUT-.t50 4.806
R24847 VOUT-.n74 VOUT-.t128 4.806
R24848 VOUT-.n75 VOUT-.t47 4.806
R24849 VOUT-.n76 VOUT-.t107 4.806
R24850 VOUT-.n77 VOUT-.t138 4.806
R24851 VOUT-.n78 VOUT-.t59 4.806
R24852 VOUT-.n79 VOUT-.t90 4.806
R24853 VOUT-.n80 VOUT-.t117 4.806
R24854 VOUT-.n81 VOUT-.t154 4.806
R24855 VOUT-.n82 VOUT-.t71 4.806
R24856 VOUT-.n83 VOUT-.t105 4.806
R24857 VOUT-.n97 VOUT-.t68 4.5005
R24858 VOUT-.n98 VOUT-.t88 4.5005
R24859 VOUT-.n102 VOUT-.t94 4.5005
R24860 VOUT-.n101 VOUT-.t123 4.5005
R24861 VOUT-.n100 VOUT-.t24 4.5005
R24862 VOUT-.n99 VOUT-.t21 4.5005
R24863 VOUT-.n113 VOUT-.t48 4.5005
R24864 VOUT-.n112 VOUT-.t145 4.5005
R24865 VOUT-.n111 VOUT-.t109 4.5005
R24866 VOUT-.n110 VOUT-.t125 4.5005
R24867 VOUT-.n109 VOUT-.t97 4.5005
R24868 VOUT-.n108 VOUT-.t61 4.5005
R24869 VOUT-.n107 VOUT-.t151 4.5005
R24870 VOUT-.n106 VOUT-.t41 4.5005
R24871 VOUT-.n105 VOUT-.t137 4.5005
R24872 VOUT-.n104 VOUT-.t120 4.5005
R24873 VOUT-.n103 VOUT-.t144 4.5005
R24874 VOUT-.n114 VOUT-.t65 4.5005
R24875 VOUT-.n116 VOUT-.t81 4.5005
R24876 VOUT-.n115 VOUT-.t44 4.5005
R24877 VOUT-.n117 VOUT-.t32 4.5005
R24878 VOUT-.n119 VOUT-.t118 4.5005
R24879 VOUT-.n118 VOUT-.t91 4.5005
R24880 VOUT-.n120 VOUT-.t130 4.5005
R24881 VOUT-.n122 VOUT-.t84 4.5005
R24882 VOUT-.n121 VOUT-.t53 4.5005
R24883 VOUT-.n123 VOUT-.t26 4.5005
R24884 VOUT-.n125 VOUT-.t112 4.5005
R24885 VOUT-.n124 VOUT-.t82 4.5005
R24886 VOUT-.n126 VOUT-.t124 4.5005
R24887 VOUT-.n128 VOUT-.t76 4.5005
R24888 VOUT-.n127 VOUT-.t45 4.5005
R24889 VOUT-.n129 VOUT-.t93 4.5005
R24890 VOUT-.n131 VOUT-.t38 4.5005
R24891 VOUT-.n130 VOUT-.t141 4.5005
R24892 VOUT-.n132 VOUT-.t119 4.5005
R24893 VOUT-.n134 VOUT-.t73 4.5005
R24894 VOUT-.n133 VOUT-.t37 4.5005
R24895 VOUT-.n135 VOUT-.t85 4.5005
R24896 VOUT-.n137 VOUT-.t31 4.5005
R24897 VOUT-.n136 VOUT-.t132 4.5005
R24898 VOUT-.n138 VOUT-.t46 4.5005
R24899 VOUT-.n140 VOUT-.t126 4.5005
R24900 VOUT-.n139 VOUT-.t100 4.5005
R24901 VOUT-.n141 VOUT-.t142 4.5005
R24902 VOUT-.n143 VOUT-.t96 4.5005
R24903 VOUT-.n142 VOUT-.t64 4.5005
R24904 VOUT-.n71 VOUT-.t55 4.5005
R24905 VOUT-.n72 VOUT-.t135 4.5005
R24906 VOUT-.n73 VOUT-.t86 4.5005
R24907 VOUT-.n84 VOUT-.t34 4.5005
R24908 VOUT-.n83 VOUT-.t133 4.5005
R24909 VOUT-.n82 VOUT-.t104 4.5005
R24910 VOUT-.n81 VOUT-.t58 4.5005
R24911 VOUT-.n80 VOUT-.t153 4.5005
R24912 VOUT-.n79 VOUT-.t116 4.5005
R24913 VOUT-.n78 VOUT-.t89 4.5005
R24914 VOUT-.n77 VOUT-.t36 4.5005
R24915 VOUT-.n76 VOUT-.t136 4.5005
R24916 VOUT-.n75 VOUT-.t78 4.5005
R24917 VOUT-.n74 VOUT-.t25 4.5005
R24918 VOUT-.n85 VOUT-.t19 4.5005
R24919 VOUT-.n87 VOUT-.t113 4.5005
R24920 VOUT-.n86 VOUT-.t29 4.5005
R24921 VOUT-.n88 VOUT-.t129 4.5005
R24922 VOUT-.n90 VOUT-.t83 4.5005
R24923 VOUT-.n89 VOUT-.t52 4.5005
R24924 VOUT-.n91 VOUT-.t101 4.5005
R24925 VOUT-.n93 VOUT-.t54 4.5005
R24926 VOUT-.n92 VOUT-.t148 4.5005
R24927 VOUT-.n94 VOUT-.t134 4.5005
R24928 VOUT-.n96 VOUT-.t92 4.5005
R24929 VOUT-.n95 VOUT-.t57 4.5005
R24930 VOUT-.n144 VOUT-.t39 4.5005
R24931 VOUT-.n145 VOUT-.t122 4.5005
R24932 VOUT-.n146 VOUT-.t95 4.5005
R24933 VOUT-.n147 VOUT-.t63 4.5005
R24934 VOUT-.n47 VOUT-.n46 4.5005
R24935 VOUT-.n45 VOUT-.n24 4.5005
R24936 VOUT-.n44 VOUT-.n23 4.5005
R24937 VOUT-.n43 VOUT-.n20 4.5005
R24938 VOUT-.n65 VOUT-.n64 4.5005
R24939 VOUT-.n16 VOUT-.n13 4.5005
R24940 VOUT-.n65 VOUT-.n13 4.5005
R24941 VOUT-.n66 VOUT-.n9 4.5005
R24942 VOUT-.n66 VOUT-.n11 4.5005
R24943 VOUT-.n66 VOUT-.n65 4.5005
R24944 VOUT-.n156 VOUT-.n69 4.5005
R24945 VOUT-.n157 VOUT-.n156 4.5005
R24946 VOUT-.n157 VOUT-.n5 4.5005
R24947 VOUT-.n158 VOUT-.n4 4.5005
R24948 VOUT-.n158 VOUT-.n157 4.5005
R24949 VOUT-.n170 VOUT-.n169 4.5005
R24950 VOUT-.n170 VOUT-.n1 4.5005
R24951 VOUT-.n166 VOUT-.n1 4.5005
R24952 VOUT-.n163 VOUT-.n1 4.5005
R24953 VOUT-.n164 VOUT-.n1 4.5005
R24954 VOUT-.n166 VOUT-.n165 4.5005
R24955 VOUT-.n165 VOUT-.n163 4.5005
R24956 VOUT-.n165 VOUT-.n164 4.5005
R24957 VOUT-.n176 VOUT-.t7 3.42907
R24958 VOUT-.n176 VOUT-.t14 3.42907
R24959 VOUT-.n172 VOUT-.t15 3.42907
R24960 VOUT-.n172 VOUT-.t5 3.42907
R24961 VOUT-.n179 VOUT-.t0 3.42907
R24962 VOUT-.n179 VOUT-.t6 3.42907
R24963 VOUT-.n63 VOUT-.n62 2.24601
R24964 VOUT-.n14 VOUT-.n8 2.24601
R24965 VOUT-.n168 VOUT-.n167 2.24601
R24966 VOUT-.n162 VOUT-.n161 2.24601
R24967 VOUT-.n155 VOUT-.n154 2.24477
R24968 VOUT-.n7 VOUT-.n2 2.24477
R24969 VOUT-.n66 VOUT-.n10 2.24063
R24970 VOUT-.n158 VOUT-.n3 2.24063
R24971 VOUT-.n165 VOUT-.n0 2.24063
R24972 VOUT-.n13 VOUT-.n12 2.24063
R24973 VOUT-.n156 VOUT-.n67 2.24063
R24974 VOUT-.n68 VOUT-.n5 2.24063
R24975 VOUT-.n169 VOUT-.n160 2.24063
R24976 VOUT-.n169 VOUT-.n159 2.24063
R24977 VOUT-.n64 VOUT-.n17 2.23934
R24978 VOUT-.n64 VOUT-.n15 2.23934
R24979 VOUT-.n177 VOUT-.n175 1.62886
R24980 VOUT-.n188 VOUT-.n173 1.52133
R24981 VOUT-.n181 VOUT-.n180 1.52133
R24982 VOUT-.n50 VOUT-.n25 1.5005
R24983 VOUT-.n52 VOUT-.n51 1.5005
R24984 VOUT-.n53 VOUT-.n22 1.5005
R24985 VOUT-.n55 VOUT-.n54 1.5005
R24986 VOUT-.n56 VOUT-.n21 1.5005
R24987 VOUT-.n58 VOUT-.n57 1.5005
R24988 VOUT-.n59 VOUT-.n18 1.5005
R24989 VOUT-.n61 VOUT-.n60 1.5005
R24990 VOUT-.n183 VOUT-.n182 1.5005
R24991 VOUT-.n184 VOUT-.n174 1.5005
R24992 VOUT-.n186 VOUT-.n185 1.5005
R24993 VOUT-.n187 VOUT-.n171 1.5005
R24994 VOUT-.n189 VOUT-.n188 1.5005
R24995 VOUT-.n30 VOUT-.n20 1.313
R24996 VOUT-.n33 VOUT-.n23 1.313
R24997 VOUT-.n36 VOUT-.n24 1.313
R24998 VOUT-.n47 VOUT-.n42 1.313
R24999 VOUT-.n28 VOUT-.n19 1.313
R25000 VOUT-.n39 VOUT-.n26 1.313
R25001 VOUT-.n154 VOUT-.n153 1.1455
R25002 VOUT-.n148 VOUT-.n6 1.13717
R25003 VOUT-.n150 VOUT-.n149 1.13717
R25004 VOUT-.n152 VOUT-.n151 1.13717
R25005 VOUT-.n157 VOUT-.n6 1.13717
R25006 VOUT-.n150 VOUT-.n7 1.13717
R25007 VOUT-.n151 VOUT-.n4 1.13717
R25008 VOUT-.n70 VOUT-.n69 1.13717
R25009 VOUT-.n49 VOUT-.n26 0.715216
R25010 VOUT-.n58 VOUT-.n20 0.65675
R25011 VOUT-.n54 VOUT-.n23 0.65675
R25012 VOUT-.n52 VOUT-.n24 0.65675
R25013 VOUT-.n48 VOUT-.n47 0.65675
R25014 VOUT-.n60 VOUT-.n19 0.65675
R25015 VOUT-.n153 VOUT-.n152 0.585
R25016 VOUT-.n50 VOUT-.n49 0.564601
R25017 VOUT-.n46 VOUT-.n45 0.563
R25018 VOUT-.n45 VOUT-.n44 0.563
R25019 VOUT-.n44 VOUT-.n43 0.563
R25020 VOUT-.n34 VOUT-.n31 0.563
R25021 VOUT-.n37 VOUT-.n34 0.563
R25022 VOUT-.n40 VOUT-.n37 0.563
R25023 VOUT-.n62 VOUT-.n61 0.5005
R25024 VOUT-.n169 VOUT-.n158 0.338
R25025 VOUT-.n98 VOUT-.n97 0.3295
R25026 VOUT-.n113 VOUT-.n99 0.3295
R25027 VOUT-.n113 VOUT-.n112 0.3295
R25028 VOUT-.n112 VOUT-.n111 0.3295
R25029 VOUT-.n111 VOUT-.n110 0.3295
R25030 VOUT-.n110 VOUT-.n109 0.3295
R25031 VOUT-.n109 VOUT-.n108 0.3295
R25032 VOUT-.n108 VOUT-.n107 0.3295
R25033 VOUT-.n107 VOUT-.n106 0.3295
R25034 VOUT-.n106 VOUT-.n105 0.3295
R25035 VOUT-.n105 VOUT-.n104 0.3295
R25036 VOUT-.n104 VOUT-.n103 0.3295
R25037 VOUT-.n116 VOUT-.n114 0.3295
R25038 VOUT-.n116 VOUT-.n115 0.3295
R25039 VOUT-.n119 VOUT-.n117 0.3295
R25040 VOUT-.n119 VOUT-.n118 0.3295
R25041 VOUT-.n122 VOUT-.n120 0.3295
R25042 VOUT-.n122 VOUT-.n121 0.3295
R25043 VOUT-.n125 VOUT-.n123 0.3295
R25044 VOUT-.n125 VOUT-.n124 0.3295
R25045 VOUT-.n128 VOUT-.n126 0.3295
R25046 VOUT-.n128 VOUT-.n127 0.3295
R25047 VOUT-.n131 VOUT-.n129 0.3295
R25048 VOUT-.n131 VOUT-.n130 0.3295
R25049 VOUT-.n134 VOUT-.n132 0.3295
R25050 VOUT-.n134 VOUT-.n133 0.3295
R25051 VOUT-.n137 VOUT-.n135 0.3295
R25052 VOUT-.n137 VOUT-.n136 0.3295
R25053 VOUT-.n140 VOUT-.n138 0.3295
R25054 VOUT-.n140 VOUT-.n139 0.3295
R25055 VOUT-.n143 VOUT-.n141 0.3295
R25056 VOUT-.n143 VOUT-.n142 0.3295
R25057 VOUT-.n72 VOUT-.n71 0.3295
R25058 VOUT-.n84 VOUT-.n73 0.3295
R25059 VOUT-.n84 VOUT-.n83 0.3295
R25060 VOUT-.n83 VOUT-.n82 0.3295
R25061 VOUT-.n82 VOUT-.n81 0.3295
R25062 VOUT-.n81 VOUT-.n80 0.3295
R25063 VOUT-.n80 VOUT-.n79 0.3295
R25064 VOUT-.n79 VOUT-.n78 0.3295
R25065 VOUT-.n78 VOUT-.n77 0.3295
R25066 VOUT-.n77 VOUT-.n76 0.3295
R25067 VOUT-.n76 VOUT-.n75 0.3295
R25068 VOUT-.n75 VOUT-.n74 0.3295
R25069 VOUT-.n87 VOUT-.n85 0.3295
R25070 VOUT-.n87 VOUT-.n86 0.3295
R25071 VOUT-.n90 VOUT-.n88 0.3295
R25072 VOUT-.n90 VOUT-.n89 0.3295
R25073 VOUT-.n93 VOUT-.n91 0.3295
R25074 VOUT-.n93 VOUT-.n92 0.3295
R25075 VOUT-.n96 VOUT-.n94 0.3295
R25076 VOUT-.n96 VOUT-.n95 0.3295
R25077 VOUT-.n145 VOUT-.n144 0.3295
R25078 VOUT-.n146 VOUT-.n145 0.3295
R25079 VOUT-.n156 VOUT-.n66 0.3205
R25080 VOUT-.n183 VOUT-.n175 0.314966
R25081 VOUT-.n147 VOUT-.n146 0.3107
R25082 VOUT-.n108 VOUT-.n102 0.306
R25083 VOUT-.n109 VOUT-.n101 0.306
R25084 VOUT-.n110 VOUT-.n100 0.306
R25085 VOUT-.n113 VOUT-.n98 0.2825
R25086 VOUT-.n116 VOUT-.n113 0.2825
R25087 VOUT-.n119 VOUT-.n116 0.2825
R25088 VOUT-.n122 VOUT-.n119 0.2825
R25089 VOUT-.n125 VOUT-.n122 0.2825
R25090 VOUT-.n128 VOUT-.n125 0.2825
R25091 VOUT-.n131 VOUT-.n128 0.2825
R25092 VOUT-.n134 VOUT-.n131 0.2825
R25093 VOUT-.n137 VOUT-.n134 0.2825
R25094 VOUT-.n140 VOUT-.n137 0.2825
R25095 VOUT-.n143 VOUT-.n140 0.2825
R25096 VOUT-.n84 VOUT-.n72 0.2825
R25097 VOUT-.n87 VOUT-.n84 0.2825
R25098 VOUT-.n90 VOUT-.n87 0.2825
R25099 VOUT-.n93 VOUT-.n90 0.2825
R25100 VOUT-.n96 VOUT-.n93 0.2825
R25101 VOUT-.n145 VOUT-.n96 0.2825
R25102 VOUT-.n145 VOUT-.n143 0.2825
R25103 VOUT-.n190 VOUT-.n189 0.28175
R25104 VOUT- VOUT-.n190 0.172375
R25105 VOUT- VOUT-.n170 0.104667
R25106 VOUT-.n148 VOUT-.n147 0.0898
R25107 VOUT-.n181 VOUT-.n175 0.0891864
R25108 VOUT-.n60 VOUT-.n59 0.0577917
R25109 VOUT-.n59 VOUT-.n58 0.0577917
R25110 VOUT-.n58 VOUT-.n21 0.0577917
R25111 VOUT-.n54 VOUT-.n21 0.0577917
R25112 VOUT-.n54 VOUT-.n53 0.0577917
R25113 VOUT-.n53 VOUT-.n52 0.0577917
R25114 VOUT-.n52 VOUT-.n25 0.0577917
R25115 VOUT-.n48 VOUT-.n25 0.0577917
R25116 VOUT-.n61 VOUT-.n18 0.0577917
R25117 VOUT-.n57 VOUT-.n18 0.0577917
R25118 VOUT-.n57 VOUT-.n56 0.0577917
R25119 VOUT-.n56 VOUT-.n55 0.0577917
R25120 VOUT-.n55 VOUT-.n22 0.0577917
R25121 VOUT-.n51 VOUT-.n22 0.0577917
R25122 VOUT-.n51 VOUT-.n50 0.0577917
R25123 VOUT-.n49 VOUT-.n48 0.054517
R25124 VOUT-.n163 VOUT-.n162 0.047375
R25125 VOUT-.n167 VOUT-.n166 0.047375
R25126 VOUT-.n157 VOUT-.n7 0.0421667
R25127 VOUT-.n65 VOUT-.n14 0.0421667
R25128 VOUT-.n188 VOUT-.n187 0.0421667
R25129 VOUT-.n187 VOUT-.n186 0.0421667
R25130 VOUT-.n186 VOUT-.n174 0.0421667
R25131 VOUT-.n182 VOUT-.n174 0.0421667
R25132 VOUT-.n182 VOUT-.n181 0.0421667
R25133 VOUT-.n189 VOUT-.n171 0.0421667
R25134 VOUT-.n185 VOUT-.n171 0.0421667
R25135 VOUT-.n185 VOUT-.n184 0.0421667
R25136 VOUT-.n184 VOUT-.n183 0.0421667
R25137 VOUT-.n15 VOUT-.n14 0.0243161
R25138 VOUT-.n17 VOUT-.n9 0.0243161
R25139 VOUT-.n17 VOUT-.n16 0.0243161
R25140 VOUT-.n15 VOUT-.n11 0.0243161
R25141 VOUT-.n154 VOUT-.n3 0.0217373
R25142 VOUT-.n62 VOUT-.n10 0.0217373
R25143 VOUT-.n16 VOUT-.n10 0.0217373
R25144 VOUT-.n69 VOUT-.n3 0.0217373
R25145 VOUT-.n170 VOUT-.n0 0.0217373
R25146 VOUT-.n167 VOUT-.n0 0.0217373
R25147 VOUT-.n67 VOUT-.n7 0.0217373
R25148 VOUT-.n69 VOUT-.n68 0.0217373
R25149 VOUT-.n12 VOUT-.n9 0.0217373
R25150 VOUT-.n12 VOUT-.n11 0.0217373
R25151 VOUT-.n67 VOUT-.n4 0.0217373
R25152 VOUT-.n68 VOUT-.n4 0.0217373
R25153 VOUT-.n164 VOUT-.n159 0.0217373
R25154 VOUT-.n163 VOUT-.n160 0.0217373
R25155 VOUT-.n166 VOUT-.n160 0.0217373
R25156 VOUT-.n162 VOUT-.n159 0.0217373
R25157 VOUT-.n149 VOUT-.n148 0.0161667
R25158 VOUT-.n152 VOUT-.n149 0.0161667
R25159 VOUT-.n150 VOUT-.n6 0.0161667
R25160 VOUT-.n151 VOUT-.n150 0.0161667
R25161 VOUT-.n151 VOUT-.n70 0.0161667
R25162 VOUT-.n155 VOUT-.n5 0.0134654
R25163 VOUT-.n158 VOUT-.n2 0.0134654
R25164 VOUT-.n156 VOUT-.n155 0.0134654
R25165 VOUT-.n5 VOUT-.n2 0.0134654
R25166 VOUT-.n63 VOUT-.n13 0.0109778
R25167 VOUT-.n66 VOUT-.n8 0.0109778
R25168 VOUT-.n168 VOUT-.n1 0.0109778
R25169 VOUT-.n165 VOUT-.n161 0.0109778
R25170 VOUT-.n64 VOUT-.n63 0.0109778
R25171 VOUT-.n13 VOUT-.n8 0.0109778
R25172 VOUT-.n169 VOUT-.n168 0.0109778
R25173 VOUT-.n161 VOUT-.n1 0.0109778
R25174 VOUT-.n153 VOUT-.n70 0.00872683
R25175 two_stage_opamp_dummy_magic_24_0.cap_res_X.t0 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 50.689
R25176 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t115 0.1603
R25177 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 0.1603
R25178 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t122 0.1603
R25179 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 two_stage_opamp_dummy_magic_24_0.cap_res_X.t82 0.1603
R25180 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 two_stage_opamp_dummy_magic_24_0.cap_res_X.t101 0.1603
R25181 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 0.1603
R25182 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 0.1603
R25183 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t51 0.1603
R25184 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 0.1603
R25185 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 two_stage_opamp_dummy_magic_24_0.cap_res_X.t91 0.1603
R25186 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 two_stage_opamp_dummy_magic_24_0.cap_res_X.t55 0.1603
R25187 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 0.1603
R25188 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 0.1603
R25189 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 0.1603
R25190 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 two_stage_opamp_dummy_magic_24_0.cap_res_X.t87 0.1603
R25191 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 two_stage_opamp_dummy_magic_24_0.cap_res_X.t7 0.1603
R25192 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 0.1603
R25193 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 0.1603
R25194 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 0.1603
R25195 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 two_stage_opamp_dummy_magic_24_0.cap_res_X.t11 0.1603
R25196 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 0.1603
R25197 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t49 0.1603
R25198 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 0.1603
R25199 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 0.1603
R25200 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 0.1603
R25201 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t54 0.1603
R25202 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 0.1603
R25203 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 two_stage_opamp_dummy_magic_24_0.cap_res_X.t90 0.1603
R25204 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 0.1603
R25205 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 0.1603
R25206 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 0.1603
R25207 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 0.1603
R25208 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 two_stage_opamp_dummy_magic_24_0.cap_res_X.t83 0.1603
R25209 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 0.1603
R25210 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 0.1603
R25211 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 two_stage_opamp_dummy_magic_24_0.cap_res_X.t46 0.1603
R25212 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 0.1603
R25213 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 0.1603
R25214 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 0.1603
R25215 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 two_stage_opamp_dummy_magic_24_0.cap_res_X.t77 0.1603
R25216 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 0.1603
R25217 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 0.1603
R25218 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 two_stage_opamp_dummy_magic_24_0.cap_res_X.t110 0.1603
R25219 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t50 0.1603
R25220 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 0.1603
R25221 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 two_stage_opamp_dummy_magic_24_0.cap_res_X.t98 0.1603
R25222 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 0.1603
R25223 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 two_stage_opamp_dummy_magic_24_0.cap_res_X.t40 0.1603
R25224 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 two_stage_opamp_dummy_magic_24_0.cap_res_X.t3 0.1603
R25225 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 two_stage_opamp_dummy_magic_24_0.cap_res_X.t86 0.1603
R25226 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 0.1603
R25227 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 0.1603
R25228 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 0.1603
R25229 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 0.1603
R25230 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 0.1603
R25231 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 0.159278
R25232 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 two_stage_opamp_dummy_magic_24_0.cap_res_X.t135 0.159278
R25233 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 two_stage_opamp_dummy_magic_24_0.cap_res_X.t114 0.159278
R25234 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 0.159278
R25235 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t95 0.159278
R25236 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t59 0.159278
R25237 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 two_stage_opamp_dummy_magic_24_0.cap_res_X.t30 0.159278
R25238 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 0.159278
R25239 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 0.159278
R25240 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 0.159278
R25241 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 0.159278
R25242 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 0.159278
R25243 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 0.159278
R25244 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 0.159278
R25245 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 0.159278
R25246 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 0.159278
R25247 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 0.159278
R25248 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 0.159278
R25249 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 0.159278
R25250 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 0.159278
R25251 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 0.159278
R25252 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 0.159278
R25253 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 0.159278
R25254 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 0.159278
R25255 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 0.159278
R25256 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 0.159278
R25257 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t10 0.159278
R25258 two_stage_opamp_dummy_magic_24_0.cap_res_X.n36 two_stage_opamp_dummy_magic_24_0.cap_res_X.t127 0.159278
R25259 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 0.137822
R25260 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 0.1368
R25261 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 0.1368
R25262 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 0.1368
R25263 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 0.1368
R25264 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 0.1368
R25265 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 0.1368
R25266 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 0.1368
R25267 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 0.1368
R25268 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 0.1368
R25269 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 0.1368
R25270 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 0.1368
R25271 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 0.1368
R25272 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 0.1368
R25273 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 0.1368
R25274 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 0.1368
R25275 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 0.1368
R25276 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 0.1368
R25277 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 0.1368
R25278 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 0.1368
R25279 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 0.1368
R25280 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 0.1368
R25281 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 0.1368
R25282 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 0.1368
R25283 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 0.1368
R25284 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 0.1368
R25285 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 0.1368
R25286 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 0.1368
R25287 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 0.1368
R25288 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 0.1368
R25289 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 0.1368
R25290 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 0.1368
R25291 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 0.1368
R25292 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 0.1368
R25293 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 0.114322
R25294 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 0.1133
R25295 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 0.1133
R25296 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 0.1133
R25297 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 0.1133
R25298 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 0.1133
R25299 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 0.1133
R25300 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 0.1133
R25301 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 0.1133
R25302 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 0.1133
R25303 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 0.1133
R25304 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 0.1133
R25305 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 0.1133
R25306 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 0.1133
R25307 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 0.1133
R25308 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 0.1133
R25309 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 0.1133
R25310 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 0.1133
R25311 two_stage_opamp_dummy_magic_24_0.cap_res_X.n36 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 0.1133
R25312 two_stage_opamp_dummy_magic_24_0.cap_res_X.n36 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 0.1133
R25313 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 0.00152174
R25314 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 0.00152174
R25315 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 0.00152174
R25316 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 0.00152174
R25317 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 0.00152174
R25318 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 0.00152174
R25319 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 0.00152174
R25320 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 0.00152174
R25321 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 0.00152174
R25322 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 0.00152174
R25323 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 0.00152174
R25324 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 0.00152174
R25325 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 0.00152174
R25326 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 0.00152174
R25327 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 0.00152174
R25328 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 0.00152174
R25329 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 0.00152174
R25330 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 0.00152174
R25331 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 0.00152174
R25332 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 0.00152174
R25333 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 0.00152174
R25334 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 0.00152174
R25335 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 0.00152174
R25336 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 0.00152174
R25337 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 0.00152174
R25338 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 0.00152174
R25339 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 0.00152174
R25340 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 0.00152174
R25341 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 0.00152174
R25342 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 0.00152174
R25343 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 0.00152174
R25344 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 0.00152174
R25345 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 0.00152174
R25346 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 0.00152174
R25347 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 0.00152174
R25348 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 0.00152174
R25349 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 two_stage_opamp_dummy_magic_24_0.cap_res_X.n36 0.00152174
R25350 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t24 731.563
R25351 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n0 621.082
R25352 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n25 617.676
R25353 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t26 369.534
R25354 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t25 369.534
R25355 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t18 369.534
R25356 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t22 369.534
R25357 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t21 369.534
R25358 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t20 369.534
R25359 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 341.397
R25360 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n11 339.272
R25361 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 339.272
R25362 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.n14 334.772
R25363 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t16 249.034
R25364 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t23 249.034
R25365 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t17 192.8
R25366 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t11 192.8
R25367 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t27 192.8
R25368 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t12 192.8
R25369 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t19 192.8
R25370 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t10 192.8
R25371 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t15 192.8
R25372 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t14 192.8
R25373 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t13 192.8
R25374 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t28 192.8
R25375 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R25376 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R25377 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.n22 176.733
R25378 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R25379 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n7 168.633
R25380 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n3 166.821
R25381 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t1 137.48
R25382 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.t6 101.165
R25383 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.n6 56.2338
R25384 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.n5 56.2338
R25385 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n2 56.2338
R25386 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R25387 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n21 56.2338
R25388 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 56.2338
R25389 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R25390 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R25391 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t0 39.4005
R25392 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R25393 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t3 39.4005
R25394 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t2 39.4005
R25395 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.t9 39.4005
R25396 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R25397 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n17 28.438
R25398 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n15 10.4693
R25399 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.n13 4.5005
R25400 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n4 4.438
R25401 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n18 2.5005
R25402 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n10 2.1255
R25403 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 2.1255
R25404 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 1.688
R25405 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t15 610.534
R25406 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t13 610.534
R25407 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t24 433.8
R25408 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t21 433.8
R25409 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t30 433.8
R25410 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t18 433.8
R25411 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t27 433.8
R25412 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t17 433.8
R25413 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t26 433.8
R25414 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t16 433.8
R25415 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t19 433.8
R25416 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t14 433.8
R25417 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t23 433.8
R25418 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t12 433.8
R25419 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t22 433.8
R25420 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t31 433.8
R25421 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t20 433.8
R25422 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t29 433.8
R25423 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t28 433.8
R25424 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t25 433.8
R25425 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 287.264
R25426 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 287.264
R25427 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 287.264
R25428 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 287.264
R25429 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 176.733
R25430 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 176.733
R25431 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 176.733
R25432 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 176.733
R25433 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 176.733
R25434 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 176.733
R25435 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 176.733
R25436 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 176.733
R25437 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 176.733
R25438 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 176.733
R25439 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 176.733
R25440 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 176.733
R25441 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 176.733
R25442 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 176.733
R25443 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 176.733
R25444 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 161.504
R25445 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n35 161.425
R25446 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 63.7586
R25447 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 63.7578
R25448 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 63.7578
R25449 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 52.5725
R25450 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 52.5725
R25451 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 52.01
R25452 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 52.01
R25453 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 50.3975
R25454 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 50.3975
R25455 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_24_0.V_tail_gate 46.7517
R25456 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 45.5227
R25457 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 45.5227
R25458 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n34 45.5227
R25459 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 45.5227
R25460 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t4 39.4005
R25461 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t1 39.4005
R25462 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t6 39.4005
R25463 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t2 39.4005
R25464 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t7 39.4005
R25465 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t3 39.4005
R25466 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t8 39.4005
R25467 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t5 39.4005
R25468 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 17.0067
R25469 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t0 16.0005
R25470 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t10 16.0005
R25471 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t11 16.0005
R25472 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t9 16.0005
R25473 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 0.170949
R25474 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 6.6358
R25475 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 0.563
R25476 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 0.170106
R25477 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 0.237927
R25478 two_stage_opamp_dummy_magic_24_0.VD3.n37 two_stage_opamp_dummy_magic_24_0.VD3.t0 672.293
R25479 two_stage_opamp_dummy_magic_24_0.VD3.n47 two_stage_opamp_dummy_magic_24_0.VD3.t3 672.293
R25480 two_stage_opamp_dummy_magic_24_0.VD3.t1 two_stage_opamp_dummy_magic_24_0.VD3.n45 213.131
R25481 two_stage_opamp_dummy_magic_24_0.VD3.n46 two_stage_opamp_dummy_magic_24_0.VD3.t4 213.131
R25482 two_stage_opamp_dummy_magic_24_0.VD3.t14 two_stage_opamp_dummy_magic_24_0.VD3.t1 146.155
R25483 two_stage_opamp_dummy_magic_24_0.VD3.t20 two_stage_opamp_dummy_magic_24_0.VD3.t14 146.155
R25484 two_stage_opamp_dummy_magic_24_0.VD3.t16 two_stage_opamp_dummy_magic_24_0.VD3.t20 146.155
R25485 two_stage_opamp_dummy_magic_24_0.VD3.t22 two_stage_opamp_dummy_magic_24_0.VD3.t16 146.155
R25486 two_stage_opamp_dummy_magic_24_0.VD3.t24 two_stage_opamp_dummy_magic_24_0.VD3.t22 146.155
R25487 two_stage_opamp_dummy_magic_24_0.VD3.t6 two_stage_opamp_dummy_magic_24_0.VD3.t24 146.155
R25488 two_stage_opamp_dummy_magic_24_0.VD3.t10 two_stage_opamp_dummy_magic_24_0.VD3.t6 146.155
R25489 two_stage_opamp_dummy_magic_24_0.VD3.t8 two_stage_opamp_dummy_magic_24_0.VD3.t10 146.155
R25490 two_stage_opamp_dummy_magic_24_0.VD3.t12 two_stage_opamp_dummy_magic_24_0.VD3.t8 146.155
R25491 two_stage_opamp_dummy_magic_24_0.VD3.t18 two_stage_opamp_dummy_magic_24_0.VD3.t12 146.155
R25492 two_stage_opamp_dummy_magic_24_0.VD3.t4 two_stage_opamp_dummy_magic_24_0.VD3.t18 146.155
R25493 two_stage_opamp_dummy_magic_24_0.VD3.n45 two_stage_opamp_dummy_magic_24_0.VD3.t2 76.2576
R25494 two_stage_opamp_dummy_magic_24_0.VD3.n46 two_stage_opamp_dummy_magic_24_0.VD3.t5 76.2576
R25495 two_stage_opamp_dummy_magic_24_0.VD3.n39 two_stage_opamp_dummy_magic_24_0.VD3.n38 66.9922
R25496 two_stage_opamp_dummy_magic_24_0.VD3.n51 two_stage_opamp_dummy_magic_24_0.VD3.n40 66.9922
R25497 two_stage_opamp_dummy_magic_24_0.VD3.n50 two_stage_opamp_dummy_magic_24_0.VD3.n41 66.9922
R25498 two_stage_opamp_dummy_magic_24_0.VD3.n49 two_stage_opamp_dummy_magic_24_0.VD3.n42 66.9922
R25499 two_stage_opamp_dummy_magic_24_0.VD3.n44 two_stage_opamp_dummy_magic_24_0.VD3.n43 66.9922
R25500 two_stage_opamp_dummy_magic_24_0.VD3.n36 two_stage_opamp_dummy_magic_24_0.VD3.n35 66.0338
R25501 two_stage_opamp_dummy_magic_24_0.VD3.n33 two_stage_opamp_dummy_magic_24_0.VD3.n32 66.0338
R25502 two_stage_opamp_dummy_magic_24_0.VD3.n31 two_stage_opamp_dummy_magic_24_0.VD3.n30 66.0338
R25503 two_stage_opamp_dummy_magic_24_0.VD3.n5 two_stage_opamp_dummy_magic_24_0.VD3.n29 66.0338
R25504 two_stage_opamp_dummy_magic_24_0.VD3.n55 two_stage_opamp_dummy_magic_24_0.VD3.n54 66.0338
R25505 two_stage_opamp_dummy_magic_24_0.VD3.n59 two_stage_opamp_dummy_magic_24_0.VD3.n58 66.0338
R25506 two_stage_opamp_dummy_magic_24_0.VD3.n35 two_stage_opamp_dummy_magic_24_0.VD3.t27 11.2576
R25507 two_stage_opamp_dummy_magic_24_0.VD3.n35 two_stage_opamp_dummy_magic_24_0.VD3.t30 11.2576
R25508 two_stage_opamp_dummy_magic_24_0.VD3.n32 two_stage_opamp_dummy_magic_24_0.VD3.t28 11.2576
R25509 two_stage_opamp_dummy_magic_24_0.VD3.n32 two_stage_opamp_dummy_magic_24_0.VD3.t31 11.2576
R25510 two_stage_opamp_dummy_magic_24_0.VD3.n30 two_stage_opamp_dummy_magic_24_0.VD3.t33 11.2576
R25511 two_stage_opamp_dummy_magic_24_0.VD3.n30 two_stage_opamp_dummy_magic_24_0.VD3.t35 11.2576
R25512 two_stage_opamp_dummy_magic_24_0.VD3.n38 two_stage_opamp_dummy_magic_24_0.VD3.t15 11.2576
R25513 two_stage_opamp_dummy_magic_24_0.VD3.n38 two_stage_opamp_dummy_magic_24_0.VD3.t21 11.2576
R25514 two_stage_opamp_dummy_magic_24_0.VD3.n40 two_stage_opamp_dummy_magic_24_0.VD3.t17 11.2576
R25515 two_stage_opamp_dummy_magic_24_0.VD3.n40 two_stage_opamp_dummy_magic_24_0.VD3.t23 11.2576
R25516 two_stage_opamp_dummy_magic_24_0.VD3.n41 two_stage_opamp_dummy_magic_24_0.VD3.t25 11.2576
R25517 two_stage_opamp_dummy_magic_24_0.VD3.n41 two_stage_opamp_dummy_magic_24_0.VD3.t7 11.2576
R25518 two_stage_opamp_dummy_magic_24_0.VD3.n42 two_stage_opamp_dummy_magic_24_0.VD3.t11 11.2576
R25519 two_stage_opamp_dummy_magic_24_0.VD3.n42 two_stage_opamp_dummy_magic_24_0.VD3.t9 11.2576
R25520 two_stage_opamp_dummy_magic_24_0.VD3.n43 two_stage_opamp_dummy_magic_24_0.VD3.t13 11.2576
R25521 two_stage_opamp_dummy_magic_24_0.VD3.n43 two_stage_opamp_dummy_magic_24_0.VD3.t19 11.2576
R25522 two_stage_opamp_dummy_magic_24_0.VD3.n29 two_stage_opamp_dummy_magic_24_0.VD3.t34 11.2576
R25523 two_stage_opamp_dummy_magic_24_0.VD3.n29 two_stage_opamp_dummy_magic_24_0.VD3.t26 11.2576
R25524 two_stage_opamp_dummy_magic_24_0.VD3.n54 two_stage_opamp_dummy_magic_24_0.VD3.t29 11.2576
R25525 two_stage_opamp_dummy_magic_24_0.VD3.n54 two_stage_opamp_dummy_magic_24_0.VD3.t32 11.2576
R25526 two_stage_opamp_dummy_magic_24_0.VD3.n59 two_stage_opamp_dummy_magic_24_0.VD3.t36 11.2576
R25527 two_stage_opamp_dummy_magic_24_0.VD3.t37 two_stage_opamp_dummy_magic_24_0.VD3.n59 11.2576
R25528 two_stage_opamp_dummy_magic_24_0.VD3.n56 two_stage_opamp_dummy_magic_24_0.VD3.n5 5.91717
R25529 two_stage_opamp_dummy_magic_24_0.VD3.n36 two_stage_opamp_dummy_magic_24_0.VD3.n34 5.91717
R25530 two_stage_opamp_dummy_magic_24_0.VD3.n34 two_stage_opamp_dummy_magic_24_0.VD3.n33 5.29217
R25531 two_stage_opamp_dummy_magic_24_0.VD3.n31 two_stage_opamp_dummy_magic_24_0.VD3.n28 5.29217
R25532 two_stage_opamp_dummy_magic_24_0.VD3.n56 two_stage_opamp_dummy_magic_24_0.VD3.n55 5.29217
R25533 two_stage_opamp_dummy_magic_24_0.VD3.n58 two_stage_opamp_dummy_magic_24_0.VD3.n57 5.29217
R25534 two_stage_opamp_dummy_magic_24_0.VD3.n7 two_stage_opamp_dummy_magic_24_0.VD3.n6 0.740726
R25535 two_stage_opamp_dummy_magic_24_0.VD3.n9 two_stage_opamp_dummy_magic_24_0.VD3.n8 0.740726
R25536 two_stage_opamp_dummy_magic_24_0.VD3.n0 two_stage_opamp_dummy_magic_24_0.VD3.n8 0.0215479
R25537 two_stage_opamp_dummy_magic_24_0.VD3.n4 two_stage_opamp_dummy_magic_24_0.VD3.n2 0.740726
R25538 two_stage_opamp_dummy_magic_24_0.VD3.n3 two_stage_opamp_dummy_magic_24_0.VD3.n1 1.5005
R25539 two_stage_opamp_dummy_magic_24_0.VD3.n23 two_stage_opamp_dummy_magic_24_0.VD3.n21 0.740726
R25540 two_stage_opamp_dummy_magic_24_0.VD3.n19 two_stage_opamp_dummy_magic_24_0.VD3.n22 0.740726
R25541 two_stage_opamp_dummy_magic_24_0.VD3.n20 two_stage_opamp_dummy_magic_24_0.VD3.n17 0.740726
R25542 two_stage_opamp_dummy_magic_24_0.VD3.n50 two_stage_opamp_dummy_magic_24_0.VD3.n20 0.0215479
R25543 two_stage_opamp_dummy_magic_24_0.VD3.n15 two_stage_opamp_dummy_magic_24_0.VD3.n18 0.740726
R25544 two_stage_opamp_dummy_magic_24_0.VD3.n16 two_stage_opamp_dummy_magic_24_0.VD3.n13 0.740726
R25545 two_stage_opamp_dummy_magic_24_0.VD3.n10 two_stage_opamp_dummy_magic_24_0.VD3.n14 0.740726
R25546 two_stage_opamp_dummy_magic_24_0.VD3.n14 two_stage_opamp_dummy_magic_24_0.VD3.n39 0.0215479
R25547 two_stage_opamp_dummy_magic_24_0.VD3.n12 two_stage_opamp_dummy_magic_24_0.VD3.n11 0.740726
R25548 two_stage_opamp_dummy_magic_24_0.VD3.n53 two_stage_opamp_dummy_magic_24_0.VD3.n52 1.5005
R25549 two_stage_opamp_dummy_magic_24_0.VD3.n27 two_stage_opamp_dummy_magic_24_0.VD3.n26 0.740726
R25550 two_stage_opamp_dummy_magic_24_0.VD3.n24 two_stage_opamp_dummy_magic_24_0.VD3.n25 0.0749176
R25551 two_stage_opamp_dummy_magic_24_0.VD3.n45 two_stage_opamp_dummy_magic_24_0.VD3.n37 1.03383
R25552 two_stage_opamp_dummy_magic_24_0.VD3.n47 two_stage_opamp_dummy_magic_24_0.VD3.n46 1.03383
R25553 two_stage_opamp_dummy_magic_24_0.VD3.n25 two_stage_opamp_dummy_magic_24_0.VD3.n36 1.04479
R25554 two_stage_opamp_dummy_magic_24_0.VD3.n48 two_stage_opamp_dummy_magic_24_0.VD3.n47 1.02322
R25555 two_stage_opamp_dummy_magic_24_0.VD3.n33 two_stage_opamp_dummy_magic_24_0.VD3.n24 0.958833
R25556 two_stage_opamp_dummy_magic_24_0.VD3.n26 two_stage_opamp_dummy_magic_24_0.VD3.n31 0.958833
R25557 two_stage_opamp_dummy_magic_24_0.VD3.n52 two_stage_opamp_dummy_magic_24_0.VD3.n37 0.958833
R25558 two_stage_opamp_dummy_magic_24_0.VD3.n55 two_stage_opamp_dummy_magic_24_0.VD3.n0 0.958833
R25559 two_stage_opamp_dummy_magic_24_0.VD3.n7 two_stage_opamp_dummy_magic_24_0.VD3.n5 0.979881
R25560 two_stage_opamp_dummy_magic_24_0.VD3.n58 two_stage_opamp_dummy_magic_24_0.VD3.n1 0.958833
R25561 two_stage_opamp_dummy_magic_24_0.VD3.n57 two_stage_opamp_dummy_magic_24_0.VD3.n56 0.6255
R25562 two_stage_opamp_dummy_magic_24_0.VD3.n34 two_stage_opamp_dummy_magic_24_0.VD3.n28 0.6255
R25563 two_stage_opamp_dummy_magic_24_0.VD3.n57 two_stage_opamp_dummy_magic_24_0.VD3.n28 0.6255
R25564 two_stage_opamp_dummy_magic_24_0.VD3.n6 two_stage_opamp_dummy_magic_24_0.VD3.n53 0.443208
R25565 two_stage_opamp_dummy_magic_24_0.VD3.n27 two_stage_opamp_dummy_magic_24_0.VD3.n25 0.37999
R25566 two_stage_opamp_dummy_magic_24_0.VD3.n21 two_stage_opamp_dummy_magic_24_0.VD3.n48 0.427973
R25567 two_stage_opamp_dummy_magic_24_0.VD3.n26 two_stage_opamp_dummy_magic_24_0.VD3.n24 0.0838333
R25568 two_stage_opamp_dummy_magic_24_0.VD3.n48 two_stage_opamp_dummy_magic_24_0.VD3.n44 0.0587394
R25569 two_stage_opamp_dummy_magic_24_0.VD3.n52 two_stage_opamp_dummy_magic_24_0.VD3.n12 0.0632146
R25570 two_stage_opamp_dummy_magic_24_0.VD3.n12 two_stage_opamp_dummy_magic_24_0.VD3.n39 0.0632146
R25571 two_stage_opamp_dummy_magic_24_0.VD3.n16 two_stage_opamp_dummy_magic_24_0.VD3.n14 0.0842626
R25572 two_stage_opamp_dummy_magic_24_0.VD3.n16 two_stage_opamp_dummy_magic_24_0.VD3.n51 0.0215479
R25573 two_stage_opamp_dummy_magic_24_0.VD3.n51 two_stage_opamp_dummy_magic_24_0.VD3.n18 0.0632146
R25574 two_stage_opamp_dummy_magic_24_0.VD3.n50 two_stage_opamp_dummy_magic_24_0.VD3.n18 0.0632146
R25575 two_stage_opamp_dummy_magic_24_0.VD3.n20 two_stage_opamp_dummy_magic_24_0.VD3.n22 0.0842626
R25576 two_stage_opamp_dummy_magic_24_0.VD3.n49 two_stage_opamp_dummy_magic_24_0.VD3.n22 0.0215479
R25577 two_stage_opamp_dummy_magic_24_0.VD3.n49 two_stage_opamp_dummy_magic_24_0.VD3.n23 0.0632146
R25578 two_stage_opamp_dummy_magic_24_0.VD3.n23 two_stage_opamp_dummy_magic_24_0.VD3.n44 0.0632146
R25579 two_stage_opamp_dummy_magic_24_0.VD3.n2 two_stage_opamp_dummy_magic_24_0.VD3.n1 0.0632146
R25580 two_stage_opamp_dummy_magic_24_0.VD3.n2 two_stage_opamp_dummy_magic_24_0.VD3.n0 0.0632146
R25581 two_stage_opamp_dummy_magic_24_0.VD3.n8 two_stage_opamp_dummy_magic_24_0.VD3.n7 0.0842626
R25582 two_stage_opamp_dummy_magic_24_0.VD3.n3 two_stage_opamp_dummy_magic_24_0.VD3.n27 0.146548
R25583 two_stage_opamp_dummy_magic_24_0.VD3.n19 two_stage_opamp_dummy_magic_24_0.VD3.n21 0.0838333
R25584 two_stage_opamp_dummy_magic_24_0.VD3.n17 two_stage_opamp_dummy_magic_24_0.VD3.n19 0.0838333
R25585 two_stage_opamp_dummy_magic_24_0.VD3.n15 two_stage_opamp_dummy_magic_24_0.VD3.n17 0.0838333
R25586 two_stage_opamp_dummy_magic_24_0.VD3.n13 two_stage_opamp_dummy_magic_24_0.VD3.n15 0.0838333
R25587 two_stage_opamp_dummy_magic_24_0.VD3.n10 two_stage_opamp_dummy_magic_24_0.VD3.n13 0.0838333
R25588 two_stage_opamp_dummy_magic_24_0.VD3.n11 two_stage_opamp_dummy_magic_24_0.VD3.n10 0.0838333
R25589 two_stage_opamp_dummy_magic_24_0.VD3.n53 two_stage_opamp_dummy_magic_24_0.VD3.n11 0.0838333
R25590 two_stage_opamp_dummy_magic_24_0.VD3.n9 two_stage_opamp_dummy_magic_24_0.VD3.n6 0.0838333
R25591 two_stage_opamp_dummy_magic_24_0.VD3.n9 two_stage_opamp_dummy_magic_24_0.VD3.n4 0.0838333
R25592 two_stage_opamp_dummy_magic_24_0.VD3.n4 two_stage_opamp_dummy_magic_24_0.VD3.n3 0.0838333
R25593 a_13430_3858.t0 a_13430_3858.t1 294.339
R25594 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t11 119.722
R25595 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 107.121
R25596 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 97.4332
R25597 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 57.7974
R25598 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 24.288
R25599 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 24.288
R25600 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 24.288
R25601 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 24.288
R25602 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 24.288
R25603 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t14 24.0005
R25604 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t7 24.0005
R25605 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t12 24.0005
R25606 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t13 24.0005
R25607 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 17.6657
R25608 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t8 8.0005
R25609 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t5 8.0005
R25610 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t1 8.0005
R25611 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t4 8.0005
R25612 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t9 8.0005
R25613 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t3 8.0005
R25614 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t0 8.0005
R25615 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t2 8.0005
R25616 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t10 8.0005
R25617 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t6 8.0005
R25618 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 5.7505
R25619 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 5.7505
R25620 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 5.7505
R25621 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 5.65675
R25622 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 5.188
R25623 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 5.188
R25624 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 5.188
R25625 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 5.188
R25626 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 5.188
R25627 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 5.188
R25628 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 5.188
R25629 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 0.563
R25630 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 0.563
R25631 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 0.563
R25632 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 0.563
R25633 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 0.563
R25634 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t0 119.722
R25635 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 107.121
R25636 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 97.4332
R25637 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 57.7974
R25638 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 24.288
R25639 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 24.288
R25640 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 24.288
R25641 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 24.288
R25642 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 24.288
R25643 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t1 24.0005
R25644 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t13 24.0005
R25645 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t12 24.0005
R25646 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t14 24.0005
R25647 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 17.6657
R25648 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t10 8.0005
R25649 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t6 8.0005
R25650 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t11 8.0005
R25651 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t5 8.0005
R25652 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t9 8.0005
R25653 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t4 8.0005
R25654 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t8 8.0005
R25655 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t3 8.0005
R25656 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t7 8.0005
R25657 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t2 8.0005
R25658 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 5.7505
R25659 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 5.7505
R25660 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 5.7505
R25661 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 5.65675
R25662 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 5.188
R25663 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 5.188
R25664 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 5.188
R25665 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 5.188
R25666 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 5.188
R25667 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 5.188
R25668 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 5.188
R25669 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 0.563
R25670 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 0.563
R25671 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 0.563
R25672 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 0.563
R25673 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 0.563
R25674 bgr_11_0.cap_res1.t20 bgr_11_0.cap_res1.t13 121.245
R25675 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t17 0.1603
R25676 bgr_11_0.cap_res1.t16 bgr_11_0.cap_res1.t19 0.1603
R25677 bgr_11_0.cap_res1.t8 bgr_11_0.cap_res1.t15 0.1603
R25678 bgr_11_0.cap_res1.t1 bgr_11_0.cap_res1.t7 0.1603
R25679 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.t14 0.1603
R25680 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t10 0.159278
R25681 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t3 0.159278
R25682 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t11 0.159278
R25683 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t18 0.159278
R25684 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t9 0.1368
R25685 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t5 0.1368
R25686 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t16 0.1368
R25687 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t12 0.1368
R25688 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t8 0.1368
R25689 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t4 0.1368
R25690 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t1 0.1368
R25691 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t0 0.1368
R25692 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t6 0.1368
R25693 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t2 0.1368
R25694 bgr_11_0.cap_res1.t10 bgr_11_0.cap_res1.n0 0.00152174
R25695 bgr_11_0.cap_res1.t3 bgr_11_0.cap_res1.n1 0.00152174
R25696 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.n2 0.00152174
R25697 bgr_11_0.cap_res1.t18 bgr_11_0.cap_res1.n3 0.00152174
R25698 bgr_11_0.cap_res1.t13 bgr_11_0.cap_res1.n4 0.00152174
R25699 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 194.296
R25700 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R25701 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R25702 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R25703 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R25704 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R25705 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R25706 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R25707 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R25708 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R25709 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R25710 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R25711 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R25712 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R25713 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R25714 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R25715 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R25716 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R25717 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R25718 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R25719 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R25720 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R25721 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R25722 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R25723 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R25724 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R25725 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R25726 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R25727 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R25728 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R25729 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R25730 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R25731 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R25732 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R25733 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R25734 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R25735 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R25736 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 65.0299
R25737 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R25738 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R25739 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R25740 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R25741 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R25742 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R25743 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R25744 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R25745 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R25746 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R25747 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R25748 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R25749 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R25750 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R25751 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R25752 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R25753 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25754 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25755 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R25756 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25757 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25758 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25759 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R25760 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25761 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25762 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25763 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25764 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R25765 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R25766 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25767 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25768 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25769 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R25770 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R25771 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25772 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25773 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R25774 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R25775 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R25776 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R25777 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R25778 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R25779 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R25780 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25781 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25782 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25783 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R25784 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25785 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25786 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25787 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R25788 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25789 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25790 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25791 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25792 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25793 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25794 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25795 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25796 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25797 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25798 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25799 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25800 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R25801 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R25802 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R25803 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R25804 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R25805 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R25806 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R25807 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R25808 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R25809 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R25810 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R25811 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R25812 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R25813 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R25814 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R25815 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R25816 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R25817 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R25818 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R25819 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R25820 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R25821 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R25822 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R25823 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R25824 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R25825 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R25826 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R25827 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R25828 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R25829 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R25830 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R25831 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R25832 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R25833 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R25834 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R25835 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R25836 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R25837 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R25838 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R25839 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R25840 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R25841 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R25842 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R25843 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R25844 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R25845 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R25846 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R25847 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R25848 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R25849 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R25850 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R25851 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R25852 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R25853 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R25854 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R25855 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R25856 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R25857 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R25858 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R25859 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R25860 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R25861 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R25862 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R25863 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R25864 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R25865 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R25866 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R25867 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R25868 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R25869 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R25870 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R25871 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R25872 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R25873 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R25874 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R25875 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R25876 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R25877 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R25878 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R25879 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R25880 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R25881 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R25882 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R25883 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R25884 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R25885 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R25886 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R25887 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R25888 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R25889 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R25890 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R25891 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R25892 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R25893 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R25894 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R25895 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R25896 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R25897 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R25898 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R25899 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R25900 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R25901 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R25902 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R25903 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R25904 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R25905 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R25906 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R25907 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R25908 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R25909 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R25910 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R25911 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R25912 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R25913 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R25914 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R25915 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25916 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25917 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25918 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R25919 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R25920 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R25921 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R25922 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R25923 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R25924 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R25925 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R25926 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R25927 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R25928 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R25929 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R25930 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R25931 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R25932 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R25933 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R25934 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R25935 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R25936 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R25937 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R25938 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R25939 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R25940 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R25941 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R25942 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R25943 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R25944 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R25945 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R25946 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R25947 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R25948 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R25949 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R25950 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R25951 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R25952 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R25953 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R25954 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R25955 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R25956 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R25957 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R25958 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R25959 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R25960 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R25961 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R25962 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R25963 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R25964 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R25965 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R25966 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R25967 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R25968 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R25969 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R25970 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R25971 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R25972 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R25973 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 two_stage_opamp_dummy_magic_24_0.V_err_gate.t6 479.322
R25974 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 two_stage_opamp_dummy_magic_24_0.V_err_gate.t8 479.322
R25975 two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 two_stage_opamp_dummy_magic_24_0.V_err_gate.t9 479.322
R25976 two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 two_stage_opamp_dummy_magic_24_0.V_err_gate.t7 479.322
R25977 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 178.625
R25978 two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 177.987
R25979 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 170.452
R25980 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 165.8
R25981 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 165.8
R25982 two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 two_stage_opamp_dummy_magic_24_0.V_err_gate.t4 24.0005
R25983 two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 two_stage_opamp_dummy_magic_24_0.V_err_gate.t5 24.0005
R25984 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 two_stage_opamp_dummy_magic_24_0.V_err_gate.t2 15.7605
R25985 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 two_stage_opamp_dummy_magic_24_0.V_err_gate.t1 15.7605
R25986 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 two_stage_opamp_dummy_magic_24_0.V_err_gate.t0 15.7605
R25987 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 two_stage_opamp_dummy_magic_24_0.V_err_gate.t3 15.7605
R25988 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 1.76612
R25989 two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 0.641125
R25990 two_stage_opamp_dummy_magic_24_0.Vb2_2.n2 two_stage_opamp_dummy_magic_24_0.Vb2_2.t3 661.375
R25991 two_stage_opamp_dummy_magic_24_0.Vb2_2.n4 two_stage_opamp_dummy_magic_24_0.Vb2_2.t0 661.375
R25992 two_stage_opamp_dummy_magic_24_0.Vb2_2.t4 two_stage_opamp_dummy_magic_24_0.Vb2_2.n0 213.131
R25993 two_stage_opamp_dummy_magic_24_0.Vb2_2.n3 two_stage_opamp_dummy_magic_24_0.Vb2_2.t1 213.131
R25994 two_stage_opamp_dummy_magic_24_0.Vb2_2.n6 two_stage_opamp_dummy_magic_24_0.Vb2_2.n1 154.983
R25995 two_stage_opamp_dummy_magic_24_0.Vb2_2.t6 two_stage_opamp_dummy_magic_24_0.Vb2_2.t4 146.155
R25996 two_stage_opamp_dummy_magic_24_0.Vb2_2.t1 two_stage_opamp_dummy_magic_24_0.Vb2_2.t6 146.155
R25997 two_stage_opamp_dummy_magic_24_0.Vb2_2.t5 two_stage_opamp_dummy_magic_24_0.Vb2_2.n0 76.2576
R25998 two_stage_opamp_dummy_magic_24_0.Vb2_2.n3 two_stage_opamp_dummy_magic_24_0.Vb2_2.t2 76.2576
R25999 two_stage_opamp_dummy_magic_24_0.Vb2_2.n7 two_stage_opamp_dummy_magic_24_0.Vb2_2.n6 66.4421
R26000 two_stage_opamp_dummy_magic_24_0.Vb2_2.n1 two_stage_opamp_dummy_magic_24_0.Vb2_2.t9 21.8894
R26001 two_stage_opamp_dummy_magic_24_0.Vb2_2.n1 two_stage_opamp_dummy_magic_24_0.Vb2_2.t8 21.8894
R26002 two_stage_opamp_dummy_magic_24_0.Vb2_2.t5 two_stage_opamp_dummy_magic_24_0.Vb2_2.n7 11.2576
R26003 two_stage_opamp_dummy_magic_24_0.Vb2_2.n7 two_stage_opamp_dummy_magic_24_0.Vb2_2.t7 11.2576
R26004 two_stage_opamp_dummy_magic_24_0.Vb2_2.n5 two_stage_opamp_dummy_magic_24_0.Vb2_2.n4 5.1255
R26005 two_stage_opamp_dummy_magic_24_0.Vb2_2.n6 two_stage_opamp_dummy_magic_24_0.Vb2_2.n5 4.92067
R26006 two_stage_opamp_dummy_magic_24_0.Vb2_2.n5 two_stage_opamp_dummy_magic_24_0.Vb2_2.n2 4.7505
R26007 two_stage_opamp_dummy_magic_24_0.Vb2_2.n4 two_stage_opamp_dummy_magic_24_0.Vb2_2.n3 1.888
R26008 two_stage_opamp_dummy_magic_24_0.Vb2_2.n2 two_stage_opamp_dummy_magic_24_0.Vb2_2.n0 1.888
R26009 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.n15 325.473
R26010 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 325.473
R26011 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 325.473
R26012 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t15 310.488
R26013 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t17 310.488
R26014 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t16 310.488
R26015 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.t9 184.097
R26016 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t11 184.097
R26017 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t1 184.097
R26018 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 167.094
R26019 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R26020 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R26021 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 152
R26022 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 152
R26023 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 152
R26024 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t14 120.501
R26025 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t3 120.501
R26026 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t13 120.501
R26027 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t5 120.501
R26028 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t18 120.501
R26029 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t7 120.501
R26030 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.t0 106.933
R26031 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 40.7027
R26032 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R26033 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R26034 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t12 39.4005
R26035 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t6 39.4005
R26036 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t2 39.4005
R26037 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t8 39.4005
R26038 bgr_11_0.V_mir1.t10 bgr_11_0.V_mir1.n16 39.4005
R26039 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.t4 39.4005
R26040 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.n4 15.9255
R26041 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n11 15.9255
R26042 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 9.3005
R26043 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.n10 4.5005
R26044 two_stage_opamp_dummy_magic_24_0.V_source.n63 two_stage_opamp_dummy_magic_24_0.V_source.t38 66.9963
R26045 two_stage_opamp_dummy_magic_24_0.V_source.n28 two_stage_opamp_dummy_magic_24_0.V_source.n27 49.3505
R26046 two_stage_opamp_dummy_magic_24_0.V_source.n25 two_stage_opamp_dummy_magic_24_0.V_source.n24 49.3505
R26047 two_stage_opamp_dummy_magic_24_0.V_source.n10 two_stage_opamp_dummy_magic_24_0.V_source.n9 49.3505
R26048 two_stage_opamp_dummy_magic_24_0.V_source.n37 two_stage_opamp_dummy_magic_24_0.V_source.n36 49.3505
R26049 two_stage_opamp_dummy_magic_24_0.V_source.n33 two_stage_opamp_dummy_magic_24_0.V_source.n32 49.3505
R26050 two_stage_opamp_dummy_magic_24_0.V_source.n31 two_stage_opamp_dummy_magic_24_0.V_source.n30 49.3505
R26051 two_stage_opamp_dummy_magic_24_0.V_source.n22 two_stage_opamp_dummy_magic_24_0.V_source.n21 49.3505
R26052 two_stage_opamp_dummy_magic_24_0.V_source.n20 two_stage_opamp_dummy_magic_24_0.V_source.n19 49.3505
R26053 two_stage_opamp_dummy_magic_24_0.V_source.n16 two_stage_opamp_dummy_magic_24_0.V_source.n15 49.3505
R26054 two_stage_opamp_dummy_magic_24_0.V_source.n12 two_stage_opamp_dummy_magic_24_0.V_source.n11 49.3505
R26055 two_stage_opamp_dummy_magic_24_0.V_source.n62 two_stage_opamp_dummy_magic_24_0.V_source.n61 32.3838
R26056 two_stage_opamp_dummy_magic_24_0.V_source.n66 two_stage_opamp_dummy_magic_24_0.V_source.n65 32.3838
R26057 two_stage_opamp_dummy_magic_24_0.V_source.n69 two_stage_opamp_dummy_magic_24_0.V_source.n68 32.3838
R26058 two_stage_opamp_dummy_magic_24_0.V_source.n56 two_stage_opamp_dummy_magic_24_0.V_source.n55 32.3838
R26059 two_stage_opamp_dummy_magic_24_0.V_source.n53 two_stage_opamp_dummy_magic_24_0.V_source.n52 32.3838
R26060 two_stage_opamp_dummy_magic_24_0.V_source.n49 two_stage_opamp_dummy_magic_24_0.V_source.n48 32.3838
R26061 two_stage_opamp_dummy_magic_24_0.V_source.n47 two_stage_opamp_dummy_magic_24_0.V_source.n46 32.3838
R26062 two_stage_opamp_dummy_magic_24_0.V_source.n43 two_stage_opamp_dummy_magic_24_0.V_source.n42 32.3838
R26063 two_stage_opamp_dummy_magic_24_0.V_source.n41 two_stage_opamp_dummy_magic_24_0.V_source.n40 32.3838
R26064 two_stage_opamp_dummy_magic_24_0.V_source.n59 two_stage_opamp_dummy_magic_24_0.V_source.n58 32.3838
R26065 two_stage_opamp_dummy_magic_24_0.V_source.n27 two_stage_opamp_dummy_magic_24_0.V_source.t36 16.0005
R26066 two_stage_opamp_dummy_magic_24_0.V_source.n27 two_stage_opamp_dummy_magic_24_0.V_source.t6 16.0005
R26067 two_stage_opamp_dummy_magic_24_0.V_source.n24 two_stage_opamp_dummy_magic_24_0.V_source.t7 16.0005
R26068 two_stage_opamp_dummy_magic_24_0.V_source.n24 two_stage_opamp_dummy_magic_24_0.V_source.t1 16.0005
R26069 two_stage_opamp_dummy_magic_24_0.V_source.n9 two_stage_opamp_dummy_magic_24_0.V_source.t29 16.0005
R26070 two_stage_opamp_dummy_magic_24_0.V_source.n9 two_stage_opamp_dummy_magic_24_0.V_source.t27 16.0005
R26071 two_stage_opamp_dummy_magic_24_0.V_source.n36 two_stage_opamp_dummy_magic_24_0.V_source.t28 16.0005
R26072 two_stage_opamp_dummy_magic_24_0.V_source.n36 two_stage_opamp_dummy_magic_24_0.V_source.t4 16.0005
R26073 two_stage_opamp_dummy_magic_24_0.V_source.n32 two_stage_opamp_dummy_magic_24_0.V_source.t35 16.0005
R26074 two_stage_opamp_dummy_magic_24_0.V_source.n32 two_stage_opamp_dummy_magic_24_0.V_source.t39 16.0005
R26075 two_stage_opamp_dummy_magic_24_0.V_source.n30 two_stage_opamp_dummy_magic_24_0.V_source.t32 16.0005
R26076 two_stage_opamp_dummy_magic_24_0.V_source.n30 two_stage_opamp_dummy_magic_24_0.V_source.t3 16.0005
R26077 two_stage_opamp_dummy_magic_24_0.V_source.n21 two_stage_opamp_dummy_magic_24_0.V_source.t31 16.0005
R26078 two_stage_opamp_dummy_magic_24_0.V_source.n21 two_stage_opamp_dummy_magic_24_0.V_source.t0 16.0005
R26079 two_stage_opamp_dummy_magic_24_0.V_source.n19 two_stage_opamp_dummy_magic_24_0.V_source.t26 16.0005
R26080 two_stage_opamp_dummy_magic_24_0.V_source.n19 two_stage_opamp_dummy_magic_24_0.V_source.t40 16.0005
R26081 two_stage_opamp_dummy_magic_24_0.V_source.n15 two_stage_opamp_dummy_magic_24_0.V_source.t2 16.0005
R26082 two_stage_opamp_dummy_magic_24_0.V_source.n15 two_stage_opamp_dummy_magic_24_0.V_source.t34 16.0005
R26083 two_stage_opamp_dummy_magic_24_0.V_source.n11 two_stage_opamp_dummy_magic_24_0.V_source.t5 16.0005
R26084 two_stage_opamp_dummy_magic_24_0.V_source.n11 two_stage_opamp_dummy_magic_24_0.V_source.t30 16.0005
R26085 two_stage_opamp_dummy_magic_24_0.V_source.n61 two_stage_opamp_dummy_magic_24_0.V_source.t18 9.6005
R26086 two_stage_opamp_dummy_magic_24_0.V_source.n61 two_stage_opamp_dummy_magic_24_0.V_source.t8 9.6005
R26087 two_stage_opamp_dummy_magic_24_0.V_source.n65 two_stage_opamp_dummy_magic_24_0.V_source.t24 9.6005
R26088 two_stage_opamp_dummy_magic_24_0.V_source.n65 two_stage_opamp_dummy_magic_24_0.V_source.t10 9.6005
R26089 two_stage_opamp_dummy_magic_24_0.V_source.n68 two_stage_opamp_dummy_magic_24_0.V_source.t37 9.6005
R26090 two_stage_opamp_dummy_magic_24_0.V_source.n68 two_stage_opamp_dummy_magic_24_0.V_source.t33 9.6005
R26091 two_stage_opamp_dummy_magic_24_0.V_source.n55 two_stage_opamp_dummy_magic_24_0.V_source.t15 9.6005
R26092 two_stage_opamp_dummy_magic_24_0.V_source.n55 two_stage_opamp_dummy_magic_24_0.V_source.t23 9.6005
R26093 two_stage_opamp_dummy_magic_24_0.V_source.n52 two_stage_opamp_dummy_magic_24_0.V_source.t14 9.6005
R26094 two_stage_opamp_dummy_magic_24_0.V_source.n52 two_stage_opamp_dummy_magic_24_0.V_source.t11 9.6005
R26095 two_stage_opamp_dummy_magic_24_0.V_source.n48 two_stage_opamp_dummy_magic_24_0.V_source.t19 9.6005
R26096 two_stage_opamp_dummy_magic_24_0.V_source.n48 two_stage_opamp_dummy_magic_24_0.V_source.t22 9.6005
R26097 two_stage_opamp_dummy_magic_24_0.V_source.n46 two_stage_opamp_dummy_magic_24_0.V_source.t9 9.6005
R26098 two_stage_opamp_dummy_magic_24_0.V_source.n46 two_stage_opamp_dummy_magic_24_0.V_source.t17 9.6005
R26099 two_stage_opamp_dummy_magic_24_0.V_source.n42 two_stage_opamp_dummy_magic_24_0.V_source.t12 9.6005
R26100 two_stage_opamp_dummy_magic_24_0.V_source.n42 two_stage_opamp_dummy_magic_24_0.V_source.t20 9.6005
R26101 two_stage_opamp_dummy_magic_24_0.V_source.n40 two_stage_opamp_dummy_magic_24_0.V_source.t13 9.6005
R26102 two_stage_opamp_dummy_magic_24_0.V_source.n40 two_stage_opamp_dummy_magic_24_0.V_source.t21 9.6005
R26103 two_stage_opamp_dummy_magic_24_0.V_source.n58 two_stage_opamp_dummy_magic_24_0.V_source.t16 9.6005
R26104 two_stage_opamp_dummy_magic_24_0.V_source.n58 two_stage_opamp_dummy_magic_24_0.V_source.t25 9.6005
R26105 two_stage_opamp_dummy_magic_24_0.V_source.n47 two_stage_opamp_dummy_magic_24_0.V_source.n45 5.89633
R26106 two_stage_opamp_dummy_magic_24_0.V_source.n69 two_stage_opamp_dummy_magic_24_0.V_source.n67 5.89633
R26107 two_stage_opamp_dummy_magic_24_0.V_source.n70 two_stage_opamp_dummy_magic_24_0.V_source.n69 5.85187
R26108 two_stage_opamp_dummy_magic_24_0.V_source.n31 two_stage_opamp_dummy_magic_24_0.V_source.n7 5.51092
R26109 two_stage_opamp_dummy_magic_24_0.V_source.n13 two_stage_opamp_dummy_magic_24_0.V_source.n10 5.51092
R26110 two_stage_opamp_dummy_magic_24_0.V_source.n34 two_stage_opamp_dummy_magic_24_0.V_source.n31 5.45883
R26111 two_stage_opamp_dummy_magic_24_0.V_source.n10 two_stage_opamp_dummy_magic_24_0.V_source.n8 5.45883
R26112 two_stage_opamp_dummy_magic_24_0.V_source.n67 two_stage_opamp_dummy_magic_24_0.V_source.n66 5.33383
R26113 two_stage_opamp_dummy_magic_24_0.V_source.n54 two_stage_opamp_dummy_magic_24_0.V_source.n53 5.33383
R26114 two_stage_opamp_dummy_magic_24_0.V_source.n49 two_stage_opamp_dummy_magic_24_0.V_source.n5 5.33383
R26115 two_stage_opamp_dummy_magic_24_0.V_source.n45 two_stage_opamp_dummy_magic_24_0.V_source.n43 5.33383
R26116 two_stage_opamp_dummy_magic_24_0.V_source.n44 two_stage_opamp_dummy_magic_24_0.V_source.n41 5.33383
R26117 two_stage_opamp_dummy_magic_24_0.V_source.n57 two_stage_opamp_dummy_magic_24_0.V_source.n56 5.33383
R26118 two_stage_opamp_dummy_magic_24_0.V_source.n60 two_stage_opamp_dummy_magic_24_0.V_source.n59 5.33383
R26119 two_stage_opamp_dummy_magic_24_0.V_source.n53 two_stage_opamp_dummy_magic_24_0.V_source.n51 5.188
R26120 two_stage_opamp_dummy_magic_24_0.V_source.n50 two_stage_opamp_dummy_magic_24_0.V_source.n49 5.188
R26121 two_stage_opamp_dummy_magic_24_0.V_source.n56 two_stage_opamp_dummy_magic_24_0.V_source.n4 5.188
R26122 two_stage_opamp_dummy_magic_24_0.V_source.n33 two_stage_opamp_dummy_magic_24_0.V_source.n7 5.16717
R26123 two_stage_opamp_dummy_magic_24_0.V_source.n38 two_stage_opamp_dummy_magic_24_0.V_source.n37 5.16717
R26124 two_stage_opamp_dummy_magic_24_0.V_source.n16 two_stage_opamp_dummy_magic_24_0.V_source.n14 5.16717
R26125 two_stage_opamp_dummy_magic_24_0.V_source.n13 two_stage_opamp_dummy_magic_24_0.V_source.n12 5.16717
R26126 two_stage_opamp_dummy_magic_24_0.V_source.n34 two_stage_opamp_dummy_magic_24_0.V_source.n33 4.89633
R26127 two_stage_opamp_dummy_magic_24_0.V_source.n29 two_stage_opamp_dummy_magic_24_0.V_source.n28 4.89633
R26128 two_stage_opamp_dummy_magic_24_0.V_source.n37 two_stage_opamp_dummy_magic_24_0.V_source.n35 4.89633
R26129 two_stage_opamp_dummy_magic_24_0.V_source.n23 two_stage_opamp_dummy_magic_24_0.V_source.n22 4.89633
R26130 two_stage_opamp_dummy_magic_24_0.V_source.n20 two_stage_opamp_dummy_magic_24_0.V_source.n18 4.89633
R26131 two_stage_opamp_dummy_magic_24_0.V_source.n17 two_stage_opamp_dummy_magic_24_0.V_source.n16 4.89633
R26132 two_stage_opamp_dummy_magic_24_0.V_source.n12 two_stage_opamp_dummy_magic_24_0.V_source.n8 4.89633
R26133 two_stage_opamp_dummy_magic_24_0.V_source.n26 two_stage_opamp_dummy_magic_24_0.V_source.n25 4.89633
R26134 two_stage_opamp_dummy_magic_24_0.V_source.n64 two_stage_opamp_dummy_magic_24_0.V_source.n63 4.5005
R26135 two_stage_opamp_dummy_magic_24_0.V_source.n26 two_stage_opamp_dummy_magic_24_0.V_source.n23 3.6255
R26136 two_stage_opamp_dummy_magic_24_0.V_source.n39 two_stage_opamp_dummy_magic_24_0.V_source.n6 2.2076
R26137 two_stage_opamp_dummy_magic_24_0.V_source.n6 two_stage_opamp_dummy_magic_24_0.V_source.n0 2.16822
R26138 two_stage_opamp_dummy_magic_24_0.V_source.n2 two_stage_opamp_dummy_magic_24_0.V_source.n39 2.16822
R26139 two_stage_opamp_dummy_magic_24_0.V_source.n50 two_stage_opamp_dummy_magic_24_0.V_source.n3 2.02255
R26140 two_stage_opamp_dummy_magic_24_0.V_source.n1 two_stage_opamp_dummy_magic_24_0.V_source.n70 1.36007
R26141 two_stage_opamp_dummy_magic_24_0.V_source.n63 two_stage_opamp_dummy_magic_24_0.V_source.n62 0.833833
R26142 two_stage_opamp_dummy_magic_24_0.V_source.n70 two_stage_opamp_dummy_magic_24_0.V_source.n4 0.66477
R26143 two_stage_opamp_dummy_magic_24_0.V_source.n62 two_stage_opamp_dummy_magic_24_0.V_source.n1 0.6255
R26144 two_stage_opamp_dummy_magic_24_0.V_source.n66 two_stage_opamp_dummy_magic_24_0.V_source.n1 0.6255
R26145 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n41 0.6255
R26146 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n43 0.6255
R26147 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n47 0.6255
R26148 two_stage_opamp_dummy_magic_24_0.V_source.n59 two_stage_opamp_dummy_magic_24_0.V_source.n1 0.6255
R26149 two_stage_opamp_dummy_magic_24_0.V_source.n0 two_stage_opamp_dummy_magic_24_0.V_source.n20 0.604667
R26150 two_stage_opamp_dummy_magic_24_0.V_source.n22 two_stage_opamp_dummy_magic_24_0.V_source.n0 0.604667
R26151 two_stage_opamp_dummy_magic_24_0.V_source.n25 two_stage_opamp_dummy_magic_24_0.V_source.n2 0.604667
R26152 two_stage_opamp_dummy_magic_24_0.V_source.n28 two_stage_opamp_dummy_magic_24_0.V_source.n2 0.604667
R26153 two_stage_opamp_dummy_magic_24_0.V_source.n35 two_stage_opamp_dummy_magic_24_0.V_source.n34 0.563
R26154 two_stage_opamp_dummy_magic_24_0.V_source.n29 two_stage_opamp_dummy_magic_24_0.V_source.n26 0.563
R26155 two_stage_opamp_dummy_magic_24_0.V_source.n35 two_stage_opamp_dummy_magic_24_0.V_source.n29 0.563
R26156 two_stage_opamp_dummy_magic_24_0.V_source.n17 two_stage_opamp_dummy_magic_24_0.V_source.n8 0.563
R26157 two_stage_opamp_dummy_magic_24_0.V_source.n18 two_stage_opamp_dummy_magic_24_0.V_source.n17 0.563
R26158 two_stage_opamp_dummy_magic_24_0.V_source.n23 two_stage_opamp_dummy_magic_24_0.V_source.n18 0.563
R26159 two_stage_opamp_dummy_magic_24_0.V_source.n45 two_stage_opamp_dummy_magic_24_0.V_source.n44 0.563
R26160 two_stage_opamp_dummy_magic_24_0.V_source.n44 two_stage_opamp_dummy_magic_24_0.V_source.n5 0.563
R26161 two_stage_opamp_dummy_magic_24_0.V_source.n54 two_stage_opamp_dummy_magic_24_0.V_source.n5 0.563
R26162 two_stage_opamp_dummy_magic_24_0.V_source.n57 two_stage_opamp_dummy_magic_24_0.V_source.n54 0.563
R26163 two_stage_opamp_dummy_magic_24_0.V_source.n60 two_stage_opamp_dummy_magic_24_0.V_source.n57 0.563
R26164 two_stage_opamp_dummy_magic_24_0.V_source.n67 two_stage_opamp_dummy_magic_24_0.V_source.n64 0.563
R26165 two_stage_opamp_dummy_magic_24_0.V_source.n64 two_stage_opamp_dummy_magic_24_0.V_source.n60 0.563
R26166 two_stage_opamp_dummy_magic_24_0.V_source.n14 two_stage_opamp_dummy_magic_24_0.V_source.n6 0.510302
R26167 two_stage_opamp_dummy_magic_24_0.V_source.n39 two_stage_opamp_dummy_magic_24_0.V_source.n38 0.510302
R26168 two_stage_opamp_dummy_magic_24_0.V_source.n14 two_stage_opamp_dummy_magic_24_0.V_source.n13 0.34425
R26169 two_stage_opamp_dummy_magic_24_0.V_source.n38 two_stage_opamp_dummy_magic_24_0.V_source.n7 0.34425
R26170 two_stage_opamp_dummy_magic_24_0.V_source.n51 two_stage_opamp_dummy_magic_24_0.V_source.n4 0.34425
R26171 two_stage_opamp_dummy_magic_24_0.V_source.n51 two_stage_opamp_dummy_magic_24_0.V_source.n50 0.34425
R26172 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n2 0.190404
R26173 two_stage_opamp_dummy_magic_24_0.V_source two_stage_opamp_dummy_magic_24_0.V_source.n1 0.120692
R26174 two_stage_opamp_dummy_magic_24_0.V_source two_stage_opamp_dummy_magic_24_0.V_source.n0 0.0702115
R26175 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t5 573.044
R26176 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t3 433.8
R26177 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n0 185.237
R26178 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n1 163.978
R26179 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n2 33.0088
R26180 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t0 15.7605
R26181 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t1 15.7605
R26182 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t4 9.6005
R26183 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n3 9.6005
R26184 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t8 651.343
R26185 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t9 647.968
R26186 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t7 540.458
R26187 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 173.591
R26188 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 169.216
R26189 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 169.216
R26190 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t6 125.111
R26191 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 70.8755
R26192 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t3 13.1338
R26193 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t5 13.1338
R26194 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t0 13.1338
R26195 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t1 13.1338
R26196 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t4 13.1338
R26197 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t2 13.1338
R26198 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 10.0317
R26199 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 4.3755
R26200 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 3.688
R26201 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 1.53175
R26202 a_4380_346.t0 a_4380_346.t1 169.905
R26203 two_stage_opamp_dummy_magic_24_0.X.n51 two_stage_opamp_dummy_magic_24_0.X.t36 1172.87
R26204 two_stage_opamp_dummy_magic_24_0.X.n47 two_stage_opamp_dummy_magic_24_0.X.t30 1172.87
R26205 two_stage_opamp_dummy_magic_24_0.X.n51 two_stage_opamp_dummy_magic_24_0.X.t52 996.134
R26206 two_stage_opamp_dummy_magic_24_0.X.n52 two_stage_opamp_dummy_magic_24_0.X.t40 996.134
R26207 two_stage_opamp_dummy_magic_24_0.X.n53 two_stage_opamp_dummy_magic_24_0.X.t33 996.134
R26208 two_stage_opamp_dummy_magic_24_0.X.n54 two_stage_opamp_dummy_magic_24_0.X.t50 996.134
R26209 two_stage_opamp_dummy_magic_24_0.X.n50 two_stage_opamp_dummy_magic_24_0.X.t34 996.134
R26210 two_stage_opamp_dummy_magic_24_0.X.n49 two_stage_opamp_dummy_magic_24_0.X.t51 996.134
R26211 two_stage_opamp_dummy_magic_24_0.X.n48 two_stage_opamp_dummy_magic_24_0.X.t37 996.134
R26212 two_stage_opamp_dummy_magic_24_0.X.n47 two_stage_opamp_dummy_magic_24_0.X.t53 996.134
R26213 two_stage_opamp_dummy_magic_24_0.X.n18 two_stage_opamp_dummy_magic_24_0.X.t43 690.867
R26214 two_stage_opamp_dummy_magic_24_0.X.n17 two_stage_opamp_dummy_magic_24_0.X.t35 690.867
R26215 two_stage_opamp_dummy_magic_24_0.X.n27 two_stage_opamp_dummy_magic_24_0.X.t46 530.201
R26216 two_stage_opamp_dummy_magic_24_0.X.n26 two_stage_opamp_dummy_magic_24_0.X.t38 530.201
R26217 two_stage_opamp_dummy_magic_24_0.X.n24 two_stage_opamp_dummy_magic_24_0.X.t45 514.134
R26218 two_stage_opamp_dummy_magic_24_0.X.n23 two_stage_opamp_dummy_magic_24_0.X.t26 514.134
R26219 two_stage_opamp_dummy_magic_24_0.X.n22 two_stage_opamp_dummy_magic_24_0.X.t42 514.134
R26220 two_stage_opamp_dummy_magic_24_0.X.n21 two_stage_opamp_dummy_magic_24_0.X.t54 514.134
R26221 two_stage_opamp_dummy_magic_24_0.X.n20 two_stage_opamp_dummy_magic_24_0.X.t39 514.134
R26222 two_stage_opamp_dummy_magic_24_0.X.n19 two_stage_opamp_dummy_magic_24_0.X.t47 514.134
R26223 two_stage_opamp_dummy_magic_24_0.X.n18 two_stage_opamp_dummy_magic_24_0.X.t27 514.134
R26224 two_stage_opamp_dummy_magic_24_0.X.n17 two_stage_opamp_dummy_magic_24_0.X.t29 514.134
R26225 two_stage_opamp_dummy_magic_24_0.X.n27 two_stage_opamp_dummy_magic_24_0.X.t31 353.467
R26226 two_stage_opamp_dummy_magic_24_0.X.n28 two_stage_opamp_dummy_magic_24_0.X.t49 353.467
R26227 two_stage_opamp_dummy_magic_24_0.X.n29 two_stage_opamp_dummy_magic_24_0.X.t41 353.467
R26228 two_stage_opamp_dummy_magic_24_0.X.n30 two_stage_opamp_dummy_magic_24_0.X.t25 353.467
R26229 two_stage_opamp_dummy_magic_24_0.X.n31 two_stage_opamp_dummy_magic_24_0.X.t44 353.467
R26230 two_stage_opamp_dummy_magic_24_0.X.n32 two_stage_opamp_dummy_magic_24_0.X.t28 353.467
R26231 two_stage_opamp_dummy_magic_24_0.X.n33 two_stage_opamp_dummy_magic_24_0.X.t48 353.467
R26232 two_stage_opamp_dummy_magic_24_0.X.n26 two_stage_opamp_dummy_magic_24_0.X.t32 353.467
R26233 two_stage_opamp_dummy_magic_24_0.X.n50 two_stage_opamp_dummy_magic_24_0.X.n49 176.733
R26234 two_stage_opamp_dummy_magic_24_0.X.n49 two_stage_opamp_dummy_magic_24_0.X.n48 176.733
R26235 two_stage_opamp_dummy_magic_24_0.X.n48 two_stage_opamp_dummy_magic_24_0.X.n47 176.733
R26236 two_stage_opamp_dummy_magic_24_0.X.n52 two_stage_opamp_dummy_magic_24_0.X.n51 176.733
R26237 two_stage_opamp_dummy_magic_24_0.X.n53 two_stage_opamp_dummy_magic_24_0.X.n52 176.733
R26238 two_stage_opamp_dummy_magic_24_0.X.n54 two_stage_opamp_dummy_magic_24_0.X.n53 176.733
R26239 two_stage_opamp_dummy_magic_24_0.X.n28 two_stage_opamp_dummy_magic_24_0.X.n27 176.733
R26240 two_stage_opamp_dummy_magic_24_0.X.n29 two_stage_opamp_dummy_magic_24_0.X.n28 176.733
R26241 two_stage_opamp_dummy_magic_24_0.X.n30 two_stage_opamp_dummy_magic_24_0.X.n29 176.733
R26242 two_stage_opamp_dummy_magic_24_0.X.n31 two_stage_opamp_dummy_magic_24_0.X.n30 176.733
R26243 two_stage_opamp_dummy_magic_24_0.X.n32 two_stage_opamp_dummy_magic_24_0.X.n31 176.733
R26244 two_stage_opamp_dummy_magic_24_0.X.n33 two_stage_opamp_dummy_magic_24_0.X.n32 176.733
R26245 two_stage_opamp_dummy_magic_24_0.X.n19 two_stage_opamp_dummy_magic_24_0.X.n18 176.733
R26246 two_stage_opamp_dummy_magic_24_0.X.n20 two_stage_opamp_dummy_magic_24_0.X.n19 176.733
R26247 two_stage_opamp_dummy_magic_24_0.X.n21 two_stage_opamp_dummy_magic_24_0.X.n20 176.733
R26248 two_stage_opamp_dummy_magic_24_0.X.n22 two_stage_opamp_dummy_magic_24_0.X.n21 176.733
R26249 two_stage_opamp_dummy_magic_24_0.X.n23 two_stage_opamp_dummy_magic_24_0.X.n22 176.733
R26250 two_stage_opamp_dummy_magic_24_0.X.n24 two_stage_opamp_dummy_magic_24_0.X.n23 176.733
R26251 two_stage_opamp_dummy_magic_24_0.X.n35 two_stage_opamp_dummy_magic_24_0.X.n34 165.472
R26252 two_stage_opamp_dummy_magic_24_0.X.n35 two_stage_opamp_dummy_magic_24_0.X.n25 165.472
R26253 two_stage_opamp_dummy_magic_24_0.X.n57 two_stage_opamp_dummy_magic_24_0.X.n56 152
R26254 two_stage_opamp_dummy_magic_24_0.X.n58 two_stage_opamp_dummy_magic_24_0.X.n57 131.571
R26255 two_stage_opamp_dummy_magic_24_0.X.n57 two_stage_opamp_dummy_magic_24_0.X.n55 124.517
R26256 two_stage_opamp_dummy_magic_24_0.X.n125 two_stage_opamp_dummy_magic_24_0.X.n35 74.3539
R26257 two_stage_opamp_dummy_magic_24_0.X.n79 two_stage_opamp_dummy_magic_24_0.X.n78 66.0338
R26258 two_stage_opamp_dummy_magic_24_0.X.n77 two_stage_opamp_dummy_magic_24_0.X.n76 66.0338
R26259 two_stage_opamp_dummy_magic_24_0.X.n89 two_stage_opamp_dummy_magic_24_0.X.n88 66.0338
R26260 two_stage_opamp_dummy_magic_24_0.X.n85 two_stage_opamp_dummy_magic_24_0.X.n84 66.0338
R26261 two_stage_opamp_dummy_magic_24_0.X.n82 two_stage_opamp_dummy_magic_24_0.X.n81 66.0338
R26262 two_stage_opamp_dummy_magic_24_0.X.n75 two_stage_opamp_dummy_magic_24_0.X.n74 66.0338
R26263 two_stage_opamp_dummy_magic_24_0.X.n6 two_stage_opamp_dummy_magic_24_0.X.n5 49.3505
R26264 two_stage_opamp_dummy_magic_24_0.X.n10 two_stage_opamp_dummy_magic_24_0.X.n9 49.3505
R26265 two_stage_opamp_dummy_magic_24_0.X.n134 two_stage_opamp_dummy_magic_24_0.X.n133 49.3505
R26266 two_stage_opamp_dummy_magic_24_0.X.n140 two_stage_opamp_dummy_magic_24_0.X.n139 49.3505
R26267 two_stage_opamp_dummy_magic_24_0.X.n143 two_stage_opamp_dummy_magic_24_0.X.n142 49.3505
R26268 two_stage_opamp_dummy_magic_24_0.X.n147 two_stage_opamp_dummy_magic_24_0.X.n146 49.3505
R26269 two_stage_opamp_dummy_magic_24_0.X.n41 two_stage_opamp_dummy_magic_24_0.X.t0 41.054
R26270 two_stage_opamp_dummy_magic_24_0.X.n55 two_stage_opamp_dummy_magic_24_0.X.n50 40.1672
R26271 two_stage_opamp_dummy_magic_24_0.X.n55 two_stage_opamp_dummy_magic_24_0.X.n54 40.1672
R26272 two_stage_opamp_dummy_magic_24_0.X.n34 two_stage_opamp_dummy_magic_24_0.X.n26 40.1672
R26273 two_stage_opamp_dummy_magic_24_0.X.n34 two_stage_opamp_dummy_magic_24_0.X.n33 40.1672
R26274 two_stage_opamp_dummy_magic_24_0.X.n25 two_stage_opamp_dummy_magic_24_0.X.n17 40.1672
R26275 two_stage_opamp_dummy_magic_24_0.X.n25 two_stage_opamp_dummy_magic_24_0.X.n24 40.1672
R26276 two_stage_opamp_dummy_magic_24_0.X.n59 two_stage_opamp_dummy_magic_24_0.X.n58 16.3217
R26277 two_stage_opamp_dummy_magic_24_0.X.n5 two_stage_opamp_dummy_magic_24_0.X.t23 16.0005
R26278 two_stage_opamp_dummy_magic_24_0.X.n5 two_stage_opamp_dummy_magic_24_0.X.t13 16.0005
R26279 two_stage_opamp_dummy_magic_24_0.X.n9 two_stage_opamp_dummy_magic_24_0.X.t14 16.0005
R26280 two_stage_opamp_dummy_magic_24_0.X.n9 two_stage_opamp_dummy_magic_24_0.X.t22 16.0005
R26281 two_stage_opamp_dummy_magic_24_0.X.n133 two_stage_opamp_dummy_magic_24_0.X.t16 16.0005
R26282 two_stage_opamp_dummy_magic_24_0.X.n133 two_stage_opamp_dummy_magic_24_0.X.t24 16.0005
R26283 two_stage_opamp_dummy_magic_24_0.X.n139 two_stage_opamp_dummy_magic_24_0.X.t18 16.0005
R26284 two_stage_opamp_dummy_magic_24_0.X.n139 two_stage_opamp_dummy_magic_24_0.X.t21 16.0005
R26285 two_stage_opamp_dummy_magic_24_0.X.n142 two_stage_opamp_dummy_magic_24_0.X.t15 16.0005
R26286 two_stage_opamp_dummy_magic_24_0.X.n142 two_stage_opamp_dummy_magic_24_0.X.t19 16.0005
R26287 two_stage_opamp_dummy_magic_24_0.X.n146 two_stage_opamp_dummy_magic_24_0.X.t17 16.0005
R26288 two_stage_opamp_dummy_magic_24_0.X.n146 two_stage_opamp_dummy_magic_24_0.X.t20 16.0005
R26289 two_stage_opamp_dummy_magic_24_0.X.n56 two_stage_opamp_dummy_magic_24_0.X.n46 12.8005
R26290 two_stage_opamp_dummy_magic_24_0.X.n78 two_stage_opamp_dummy_magic_24_0.X.t9 11.2576
R26291 two_stage_opamp_dummy_magic_24_0.X.n78 two_stage_opamp_dummy_magic_24_0.X.t2 11.2576
R26292 two_stage_opamp_dummy_magic_24_0.X.n76 two_stage_opamp_dummy_magic_24_0.X.t1 11.2576
R26293 two_stage_opamp_dummy_magic_24_0.X.n76 two_stage_opamp_dummy_magic_24_0.X.t7 11.2576
R26294 two_stage_opamp_dummy_magic_24_0.X.n88 two_stage_opamp_dummy_magic_24_0.X.t10 11.2576
R26295 two_stage_opamp_dummy_magic_24_0.X.n88 two_stage_opamp_dummy_magic_24_0.X.t8 11.2576
R26296 two_stage_opamp_dummy_magic_24_0.X.n84 two_stage_opamp_dummy_magic_24_0.X.t11 11.2576
R26297 two_stage_opamp_dummy_magic_24_0.X.n84 two_stage_opamp_dummy_magic_24_0.X.t12 11.2576
R26298 two_stage_opamp_dummy_magic_24_0.X.n81 two_stage_opamp_dummy_magic_24_0.X.t3 11.2576
R26299 two_stage_opamp_dummy_magic_24_0.X.n81 two_stage_opamp_dummy_magic_24_0.X.t5 11.2576
R26300 two_stage_opamp_dummy_magic_24_0.X.n74 two_stage_opamp_dummy_magic_24_0.X.t4 11.2576
R26301 two_stage_opamp_dummy_magic_24_0.X.n74 two_stage_opamp_dummy_magic_24_0.X.t6 11.2576
R26302 two_stage_opamp_dummy_magic_24_0.X.n56 two_stage_opamp_dummy_magic_24_0.X.n44 9.36264
R26303 two_stage_opamp_dummy_magic_24_0.X.n46 two_stage_opamp_dummy_magic_24_0.X.n45 9.3005
R26304 two_stage_opamp_dummy_magic_24_0.X.n87 two_stage_opamp_dummy_magic_24_0.X.n77 5.91717
R26305 two_stage_opamp_dummy_magic_24_0.X.n80 two_stage_opamp_dummy_magic_24_0.X.n79 5.91717
R26306 two_stage_opamp_dummy_magic_24_0.X.n10 two_stage_opamp_dummy_magic_24_0.X.n8 5.6255
R26307 two_stage_opamp_dummy_magic_24_0.X.n145 two_stage_opamp_dummy_magic_24_0.X.n6 5.6255
R26308 two_stage_opamp_dummy_magic_24_0.X.n58 two_stage_opamp_dummy_magic_24_0.X.n46 5.33141
R26309 two_stage_opamp_dummy_magic_24_0.X.n89 two_stage_opamp_dummy_magic_24_0.X.n87 5.29217
R26310 two_stage_opamp_dummy_magic_24_0.X.n86 two_stage_opamp_dummy_magic_24_0.X.n85 5.29217
R26311 two_stage_opamp_dummy_magic_24_0.X.n83 two_stage_opamp_dummy_magic_24_0.X.n82 5.29217
R26312 two_stage_opamp_dummy_magic_24_0.X.n80 two_stage_opamp_dummy_magic_24_0.X.n75 5.29217
R26313 two_stage_opamp_dummy_magic_24_0.X.n94 two_stage_opamp_dummy_magic_24_0.X.n73 5.1255
R26314 two_stage_opamp_dummy_magic_24_0.X.n91 two_stage_opamp_dummy_magic_24_0.X.n65 5.1255
R26315 two_stage_opamp_dummy_magic_24_0.X.n134 two_stage_opamp_dummy_magic_24_0.X.n8 5.063
R26316 two_stage_opamp_dummy_magic_24_0.X.n141 two_stage_opamp_dummy_magic_24_0.X.n140 5.063
R26317 two_stage_opamp_dummy_magic_24_0.X.n144 two_stage_opamp_dummy_magic_24_0.X.n143 5.063
R26318 two_stage_opamp_dummy_magic_24_0.X.n147 two_stage_opamp_dummy_magic_24_0.X.n145 5.063
R26319 two_stage_opamp_dummy_magic_24_0.X.n150 two_stage_opamp_dummy_magic_24_0.X.n149 5.063
R26320 two_stage_opamp_dummy_magic_24_0.X.n136 two_stage_opamp_dummy_magic_24_0.X.n11 5.063
R26321 two_stage_opamp_dummy_magic_24_0.X.n95 two_stage_opamp_dummy_magic_24_0.X.n94 4.5005
R26322 two_stage_opamp_dummy_magic_24_0.X.n93 two_stage_opamp_dummy_magic_24_0.X.n71 4.5005
R26323 two_stage_opamp_dummy_magic_24_0.X.n92 two_stage_opamp_dummy_magic_24_0.X.n68 4.5005
R26324 two_stage_opamp_dummy_magic_24_0.X.n91 two_stage_opamp_dummy_magic_24_0.X.n90 4.5005
R26325 two_stage_opamp_dummy_magic_24_0.X.n119 two_stage_opamp_dummy_magic_24_0.X.n118 4.5005
R26326 two_stage_opamp_dummy_magic_24_0.X.n149 two_stage_opamp_dummy_magic_24_0.X.n148 4.5005
R26327 two_stage_opamp_dummy_magic_24_0.X.n7 two_stage_opamp_dummy_magic_24_0.X.n3 4.5005
R26328 two_stage_opamp_dummy_magic_24_0.X.n138 two_stage_opamp_dummy_magic_24_0.X.n137 4.5005
R26329 two_stage_opamp_dummy_magic_24_0.X.n136 two_stage_opamp_dummy_magic_24_0.X.n135 4.5005
R26330 two_stage_opamp_dummy_magic_24_0.X.n124 two_stage_opamp_dummy_magic_24_0.X.n61 4.5005
R26331 two_stage_opamp_dummy_magic_24_0.X.n126 two_stage_opamp_dummy_magic_24_0.X.n125 4.5005
R26332 two_stage_opamp_dummy_magic_24_0.X.n125 two_stage_opamp_dummy_magic_24_0.X.n124 4.5005
R26333 two_stage_opamp_dummy_magic_24_0.X.n60 two_stage_opamp_dummy_magic_24_0.X.n59 4.5005
R26334 two_stage_opamp_dummy_magic_24_0.X.n38 two_stage_opamp_dummy_magic_24_0.X.n37 4.5005
R26335 two_stage_opamp_dummy_magic_24_0.X.n120 two_stage_opamp_dummy_magic_24_0.X.n63 2.26187
R26336 two_stage_opamp_dummy_magic_24_0.X.n40 two_stage_opamp_dummy_magic_24_0.X.n39 2.26187
R26337 two_stage_opamp_dummy_magic_24_0.X.n39 two_stage_opamp_dummy_magic_24_0.X.n36 2.26187
R26338 two_stage_opamp_dummy_magic_24_0.X.n117 two_stage_opamp_dummy_magic_24_0.X.n63 2.26187
R26339 two_stage_opamp_dummy_magic_24_0.X.n121 two_stage_opamp_dummy_magic_24_0.X.n62 2.24063
R26340 two_stage_opamp_dummy_magic_24_0.X.n126 two_stage_opamp_dummy_magic_24_0.X.n15 2.24063
R26341 two_stage_opamp_dummy_magic_24_0.X.n16 two_stage_opamp_dummy_magic_24_0.X.n14 2.24063
R26342 two_stage_opamp_dummy_magic_24_0.X.n117 two_stage_opamp_dummy_magic_24_0.X.n116 2.24063
R26343 two_stage_opamp_dummy_magic_24_0.X.n123 two_stage_opamp_dummy_magic_24_0.X.n122 2.24063
R26344 two_stage_opamp_dummy_magic_24_0.X.n41 two_stage_opamp_dummy_magic_24_0.X.n40 2.24063
R26345 two_stage_opamp_dummy_magic_24_0.X.n43 two_stage_opamp_dummy_magic_24_0.X.n42 2.24063
R26346 two_stage_opamp_dummy_magic_24_0.X.n60 two_stage_opamp_dummy_magic_24_0.X.n44 2.22018
R26347 two_stage_opamp_dummy_magic_24_0.X.n98 two_stage_opamp_dummy_magic_24_0.X.n72 1.5005
R26348 two_stage_opamp_dummy_magic_24_0.X.n100 two_stage_opamp_dummy_magic_24_0.X.n99 1.5005
R26349 two_stage_opamp_dummy_magic_24_0.X.n101 two_stage_opamp_dummy_magic_24_0.X.n70 1.5005
R26350 two_stage_opamp_dummy_magic_24_0.X.n103 two_stage_opamp_dummy_magic_24_0.X.n102 1.5005
R26351 two_stage_opamp_dummy_magic_24_0.X.n104 two_stage_opamp_dummy_magic_24_0.X.n69 1.5005
R26352 two_stage_opamp_dummy_magic_24_0.X.n106 two_stage_opamp_dummy_magic_24_0.X.n105 1.5005
R26353 two_stage_opamp_dummy_magic_24_0.X.n107 two_stage_opamp_dummy_magic_24_0.X.n67 1.5005
R26354 two_stage_opamp_dummy_magic_24_0.X.n109 two_stage_opamp_dummy_magic_24_0.X.n108 1.5005
R26355 two_stage_opamp_dummy_magic_24_0.X.n110 two_stage_opamp_dummy_magic_24_0.X.n66 1.5005
R26356 two_stage_opamp_dummy_magic_24_0.X.n112 two_stage_opamp_dummy_magic_24_0.X.n111 1.5005
R26357 two_stage_opamp_dummy_magic_24_0.X.n113 two_stage_opamp_dummy_magic_24_0.X.n64 1.5005
R26358 two_stage_opamp_dummy_magic_24_0.X.n115 two_stage_opamp_dummy_magic_24_0.X.n114 1.5005
R26359 two_stage_opamp_dummy_magic_24_0.X.n153 two_stage_opamp_dummy_magic_24_0.X.n152 1.5005
R26360 two_stage_opamp_dummy_magic_24_0.X.n154 two_stage_opamp_dummy_magic_24_0.X.n1 1.5005
R26361 two_stage_opamp_dummy_magic_24_0.X.n156 two_stage_opamp_dummy_magic_24_0.X.n155 1.5005
R26362 two_stage_opamp_dummy_magic_24_0.X.n2 two_stage_opamp_dummy_magic_24_0.X.n0 1.5005
R26363 two_stage_opamp_dummy_magic_24_0.X.n130 two_stage_opamp_dummy_magic_24_0.X.n13 1.5005
R26364 two_stage_opamp_dummy_magic_24_0.X.n132 two_stage_opamp_dummy_magic_24_0.X.n131 1.5005
R26365 two_stage_opamp_dummy_magic_24_0.X.n129 two_stage_opamp_dummy_magic_24_0.X.n12 1.5005
R26366 two_stage_opamp_dummy_magic_24_0.X.n128 two_stage_opamp_dummy_magic_24_0.X.n127 1.5005
R26367 two_stage_opamp_dummy_magic_24_0.X.n122 two_stage_opamp_dummy_magic_24_0.X.n121 0.891125
R26368 two_stage_opamp_dummy_magic_24_0.X.n60 two_stage_opamp_dummy_magic_24_0.X.n43 0.891125
R26369 two_stage_opamp_dummy_magic_24_0.X.n151 two_stage_opamp_dummy_magic_24_0.X.n150 0.887091
R26370 two_stage_opamp_dummy_magic_24_0.X.n135 two_stage_opamp_dummy_magic_24_0.X.n132 0.828625
R26371 two_stage_opamp_dummy_magic_24_0.X.n138 two_stage_opamp_dummy_magic_24_0.X.n2 0.828625
R26372 two_stage_opamp_dummy_magic_24_0.X.n154 two_stage_opamp_dummy_magic_24_0.X.n3 0.828625
R26373 two_stage_opamp_dummy_magic_24_0.X.n148 two_stage_opamp_dummy_magic_24_0.X.n4 0.828625
R26374 two_stage_opamp_dummy_magic_24_0.X.n127 two_stage_opamp_dummy_magic_24_0.X.n11 0.828625
R26375 two_stage_opamp_dummy_magic_24_0.X.n90 two_stage_opamp_dummy_magic_24_0.X.n89 0.792167
R26376 two_stage_opamp_dummy_magic_24_0.X.n85 two_stage_opamp_dummy_magic_24_0.X.n68 0.792167
R26377 two_stage_opamp_dummy_magic_24_0.X.n82 two_stage_opamp_dummy_magic_24_0.X.n71 0.792167
R26378 two_stage_opamp_dummy_magic_24_0.X.n95 two_stage_opamp_dummy_magic_24_0.X.n75 0.792167
R26379 two_stage_opamp_dummy_magic_24_0.X.n77 two_stage_opamp_dummy_magic_24_0.X.n65 0.792167
R26380 two_stage_opamp_dummy_magic_24_0.X.n79 two_stage_opamp_dummy_magic_24_0.X.n73 0.792167
R26381 two_stage_opamp_dummy_magic_24_0.X.n94 two_stage_opamp_dummy_magic_24_0.X.n93 0.6255
R26382 two_stage_opamp_dummy_magic_24_0.X.n93 two_stage_opamp_dummy_magic_24_0.X.n92 0.6255
R26383 two_stage_opamp_dummy_magic_24_0.X.n92 two_stage_opamp_dummy_magic_24_0.X.n91 0.6255
R26384 two_stage_opamp_dummy_magic_24_0.X.n87 two_stage_opamp_dummy_magic_24_0.X.n86 0.6255
R26385 two_stage_opamp_dummy_magic_24_0.X.n86 two_stage_opamp_dummy_magic_24_0.X.n83 0.6255
R26386 two_stage_opamp_dummy_magic_24_0.X.n83 two_stage_opamp_dummy_magic_24_0.X.n80 0.6255
R26387 two_stage_opamp_dummy_magic_24_0.X.n152 two_stage_opamp_dummy_magic_24_0.X.n151 0.564601
R26388 two_stage_opamp_dummy_magic_24_0.X.n149 two_stage_opamp_dummy_magic_24_0.X.n7 0.563
R26389 two_stage_opamp_dummy_magic_24_0.X.n137 two_stage_opamp_dummy_magic_24_0.X.n7 0.563
R26390 two_stage_opamp_dummy_magic_24_0.X.n137 two_stage_opamp_dummy_magic_24_0.X.n136 0.563
R26391 two_stage_opamp_dummy_magic_24_0.X.n141 two_stage_opamp_dummy_magic_24_0.X.n8 0.563
R26392 two_stage_opamp_dummy_magic_24_0.X.n144 two_stage_opamp_dummy_magic_24_0.X.n141 0.563
R26393 two_stage_opamp_dummy_magic_24_0.X.n145 two_stage_opamp_dummy_magic_24_0.X.n144 0.563
R26394 two_stage_opamp_dummy_magic_24_0.X.n97 two_stage_opamp_dummy_magic_24_0.X.n73 0.533638
R26395 two_stage_opamp_dummy_magic_24_0.X.n90 two_stage_opamp_dummy_magic_24_0.X.n66 0.46925
R26396 two_stage_opamp_dummy_magic_24_0.X.n106 two_stage_opamp_dummy_magic_24_0.X.n68 0.46925
R26397 two_stage_opamp_dummy_magic_24_0.X.n101 two_stage_opamp_dummy_magic_24_0.X.n71 0.46925
R26398 two_stage_opamp_dummy_magic_24_0.X.n96 two_stage_opamp_dummy_magic_24_0.X.n95 0.46925
R26399 two_stage_opamp_dummy_magic_24_0.X.n114 two_stage_opamp_dummy_magic_24_0.X.n65 0.46925
R26400 two_stage_opamp_dummy_magic_24_0.X.n124 two_stage_opamp_dummy_magic_24_0.X.n60 0.46925
R26401 two_stage_opamp_dummy_magic_24_0.X.n98 two_stage_opamp_dummy_magic_24_0.X.n97 0.427973
R26402 two_stage_opamp_dummy_magic_24_0.X.n128 two_stage_opamp_dummy_magic_24_0.X.n126 0.422375
R26403 two_stage_opamp_dummy_magic_24_0.X.n116 two_stage_opamp_dummy_magic_24_0.X.n115 0.401542
R26404 two_stage_opamp_dummy_magic_24_0.X.n135 two_stage_opamp_dummy_magic_24_0.X.n134 0.3755
R26405 two_stage_opamp_dummy_magic_24_0.X.n140 two_stage_opamp_dummy_magic_24_0.X.n138 0.3755
R26406 two_stage_opamp_dummy_magic_24_0.X.n143 two_stage_opamp_dummy_magic_24_0.X.n3 0.3755
R26407 two_stage_opamp_dummy_magic_24_0.X.n148 two_stage_opamp_dummy_magic_24_0.X.n147 0.3755
R26408 two_stage_opamp_dummy_magic_24_0.X.n11 two_stage_opamp_dummy_magic_24_0.X.n10 0.3755
R26409 two_stage_opamp_dummy_magic_24_0.X.n150 two_stage_opamp_dummy_magic_24_0.X.n6 0.3755
R26410 two_stage_opamp_dummy_magic_24_0.X.n59 two_stage_opamp_dummy_magic_24_0.X.n45 0.1255
R26411 two_stage_opamp_dummy_magic_24_0.X.n45 two_stage_opamp_dummy_magic_24_0.X.n44 0.0626438
R26412 two_stage_opamp_dummy_magic_24_0.X.n97 two_stage_opamp_dummy_magic_24_0.X.n96 0.0587394
R26413 two_stage_opamp_dummy_magic_24_0.X.n127 two_stage_opamp_dummy_magic_24_0.X.n12 0.0577917
R26414 two_stage_opamp_dummy_magic_24_0.X.n132 two_stage_opamp_dummy_magic_24_0.X.n12 0.0577917
R26415 two_stage_opamp_dummy_magic_24_0.X.n132 two_stage_opamp_dummy_magic_24_0.X.n13 0.0577917
R26416 two_stage_opamp_dummy_magic_24_0.X.n13 two_stage_opamp_dummy_magic_24_0.X.n2 0.0577917
R26417 two_stage_opamp_dummy_magic_24_0.X.n155 two_stage_opamp_dummy_magic_24_0.X.n2 0.0577917
R26418 two_stage_opamp_dummy_magic_24_0.X.n155 two_stage_opamp_dummy_magic_24_0.X.n154 0.0577917
R26419 two_stage_opamp_dummy_magic_24_0.X.n154 two_stage_opamp_dummy_magic_24_0.X.n153 0.0577917
R26420 two_stage_opamp_dummy_magic_24_0.X.n153 two_stage_opamp_dummy_magic_24_0.X.n4 0.0577917
R26421 two_stage_opamp_dummy_magic_24_0.X.n129 two_stage_opamp_dummy_magic_24_0.X.n128 0.0577917
R26422 two_stage_opamp_dummy_magic_24_0.X.n131 two_stage_opamp_dummy_magic_24_0.X.n129 0.0577917
R26423 two_stage_opamp_dummy_magic_24_0.X.n131 two_stage_opamp_dummy_magic_24_0.X.n130 0.0577917
R26424 two_stage_opamp_dummy_magic_24_0.X.n130 two_stage_opamp_dummy_magic_24_0.X.n0 0.0577917
R26425 two_stage_opamp_dummy_magic_24_0.X.n156 two_stage_opamp_dummy_magic_24_0.X.n1 0.0577917
R26426 two_stage_opamp_dummy_magic_24_0.X.n152 two_stage_opamp_dummy_magic_24_0.X.n1 0.0577917
R26427 two_stage_opamp_dummy_magic_24_0.X.n151 two_stage_opamp_dummy_magic_24_0.X.n4 0.054517
R26428 two_stage_opamp_dummy_magic_24_0.X.n114 two_stage_opamp_dummy_magic_24_0.X.n113 0.0421667
R26429 two_stage_opamp_dummy_magic_24_0.X.n113 two_stage_opamp_dummy_magic_24_0.X.n112 0.0421667
R26430 two_stage_opamp_dummy_magic_24_0.X.n112 two_stage_opamp_dummy_magic_24_0.X.n66 0.0421667
R26431 two_stage_opamp_dummy_magic_24_0.X.n108 two_stage_opamp_dummy_magic_24_0.X.n66 0.0421667
R26432 two_stage_opamp_dummy_magic_24_0.X.n108 two_stage_opamp_dummy_magic_24_0.X.n107 0.0421667
R26433 two_stage_opamp_dummy_magic_24_0.X.n107 two_stage_opamp_dummy_magic_24_0.X.n106 0.0421667
R26434 two_stage_opamp_dummy_magic_24_0.X.n106 two_stage_opamp_dummy_magic_24_0.X.n69 0.0421667
R26435 two_stage_opamp_dummy_magic_24_0.X.n102 two_stage_opamp_dummy_magic_24_0.X.n69 0.0421667
R26436 two_stage_opamp_dummy_magic_24_0.X.n102 two_stage_opamp_dummy_magic_24_0.X.n101 0.0421667
R26437 two_stage_opamp_dummy_magic_24_0.X.n101 two_stage_opamp_dummy_magic_24_0.X.n100 0.0421667
R26438 two_stage_opamp_dummy_magic_24_0.X.n100 two_stage_opamp_dummy_magic_24_0.X.n72 0.0421667
R26439 two_stage_opamp_dummy_magic_24_0.X.n96 two_stage_opamp_dummy_magic_24_0.X.n72 0.0421667
R26440 two_stage_opamp_dummy_magic_24_0.X.n115 two_stage_opamp_dummy_magic_24_0.X.n64 0.0421667
R26441 two_stage_opamp_dummy_magic_24_0.X.n111 two_stage_opamp_dummy_magic_24_0.X.n64 0.0421667
R26442 two_stage_opamp_dummy_magic_24_0.X.n111 two_stage_opamp_dummy_magic_24_0.X.n110 0.0421667
R26443 two_stage_opamp_dummy_magic_24_0.X.n110 two_stage_opamp_dummy_magic_24_0.X.n109 0.0421667
R26444 two_stage_opamp_dummy_magic_24_0.X.n109 two_stage_opamp_dummy_magic_24_0.X.n67 0.0421667
R26445 two_stage_opamp_dummy_magic_24_0.X.n105 two_stage_opamp_dummy_magic_24_0.X.n67 0.0421667
R26446 two_stage_opamp_dummy_magic_24_0.X.n105 two_stage_opamp_dummy_magic_24_0.X.n104 0.0421667
R26447 two_stage_opamp_dummy_magic_24_0.X.n104 two_stage_opamp_dummy_magic_24_0.X.n103 0.0421667
R26448 two_stage_opamp_dummy_magic_24_0.X.n103 two_stage_opamp_dummy_magic_24_0.X.n70 0.0421667
R26449 two_stage_opamp_dummy_magic_24_0.X.n99 two_stage_opamp_dummy_magic_24_0.X.n70 0.0421667
R26450 two_stage_opamp_dummy_magic_24_0.X.n99 two_stage_opamp_dummy_magic_24_0.X.n98 0.0421667
R26451 two_stage_opamp_dummy_magic_24_0.X.n126 two_stage_opamp_dummy_magic_24_0.X.n14 0.0421667
R26452 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.X.n156 0.0369583
R26453 two_stage_opamp_dummy_magic_24_0.X.n116 two_stage_opamp_dummy_magic_24_0.X.n62 0.0217373
R26454 two_stage_opamp_dummy_magic_24_0.X.n120 two_stage_opamp_dummy_magic_24_0.X.n119 0.0217373
R26455 two_stage_opamp_dummy_magic_24_0.X.n122 two_stage_opamp_dummy_magic_24_0.X.n15 0.0217373
R26456 two_stage_opamp_dummy_magic_24_0.X.n125 two_stage_opamp_dummy_magic_24_0.X.n16 0.0217373
R26457 two_stage_opamp_dummy_magic_24_0.X.n118 two_stage_opamp_dummy_magic_24_0.X.n62 0.0217373
R26458 two_stage_opamp_dummy_magic_24_0.X.n121 two_stage_opamp_dummy_magic_24_0.X.n120 0.0217373
R26459 two_stage_opamp_dummy_magic_24_0.X.n43 two_stage_opamp_dummy_magic_24_0.X.n36 0.0217373
R26460 two_stage_opamp_dummy_magic_24_0.X.n61 two_stage_opamp_dummy_magic_24_0.X.n15 0.0217373
R26461 two_stage_opamp_dummy_magic_24_0.X.n61 two_stage_opamp_dummy_magic_24_0.X.n16 0.0217373
R26462 two_stage_opamp_dummy_magic_24_0.X.n39 two_stage_opamp_dummy_magic_24_0.X.n37 0.0217373
R26463 two_stage_opamp_dummy_magic_24_0.X.n38 two_stage_opamp_dummy_magic_24_0.X.n36 0.0217373
R26464 two_stage_opamp_dummy_magic_24_0.X.n118 two_stage_opamp_dummy_magic_24_0.X.n63 0.0217373
R26465 two_stage_opamp_dummy_magic_24_0.X.n119 two_stage_opamp_dummy_magic_24_0.X.n117 0.0217373
R26466 two_stage_opamp_dummy_magic_24_0.X.n40 two_stage_opamp_dummy_magic_24_0.X.n38 0.0217373
R26467 two_stage_opamp_dummy_magic_24_0.X.n124 two_stage_opamp_dummy_magic_24_0.X.n123 0.0217373
R26468 two_stage_opamp_dummy_magic_24_0.X.n123 two_stage_opamp_dummy_magic_24_0.X.n14 0.0217373
R26469 two_stage_opamp_dummy_magic_24_0.X.n42 two_stage_opamp_dummy_magic_24_0.X.n37 0.0217373
R26470 two_stage_opamp_dummy_magic_24_0.X.n42 two_stage_opamp_dummy_magic_24_0.X.n41 0.0217373
R26471 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.X.n0 0.0213333
R26472 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 344.837
R26473 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 344.274
R26474 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 292.5
R26475 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t16 121.724
R26476 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 118.861
R26477 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 118.861
R26478 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 118.861
R26479 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 118.861
R26480 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 118.861
R26481 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 75.063
R26482 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 52.3363
R26483 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 52.1563
R26484 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t15 39.4005
R26485 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t12 39.4005
R26486 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t10 39.4005
R26487 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t13 39.4005
R26488 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t11 39.4005
R26489 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t14 39.4005
R26490 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t6 19.7005
R26491 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t5 19.7005
R26492 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t8 19.7005
R26493 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t1 19.7005
R26494 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t9 19.7005
R26495 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t3 19.7005
R26496 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t0 19.7005
R26497 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t4 19.7005
R26498 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t2 19.7005
R26499 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t7 19.7005
R26500 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 5.938
R26501 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 5.60467
R26502 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 5.54217
R26503 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 5.54217
R26504 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 5.04217
R26505 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 5.04217
R26506 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 5.04217
R26507 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 5.04217
R26508 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 4.97967
R26509 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 4.97967
R26510 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 4.97967
R26511 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 0.563
R26512 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 0.563
R26513 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 0.563
R26514 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 0.563
R26515 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 0.563
R26516 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t7 355.293
R26517 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t8 346.8
R26518 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n10 339.522
R26519 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n6 339.522
R26520 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n5 335.022
R26521 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t19 184.097
R26522 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t27 184.097
R26523 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t14 184.097
R26524 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t26 184.097
R26525 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n11 166.05
R26526 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n8 166.05
R26527 bgr_11_0.1st_Vout_2.t4 bgr_11_0.1st_Vout_2.n12 106.556
R26528 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n0 51.9009
R26529 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t1 39.4005
R26530 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t3 39.4005
R26531 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t6 39.4005
R26532 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t2 39.4005
R26533 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t0 39.4005
R26534 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t5 39.4005
R26535 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t32 4.8295
R26536 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t12 4.8295
R26537 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t13 4.8295
R26538 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t18 4.8295
R26539 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t30 4.8295
R26540 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t11 4.8295
R26541 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t22 4.8295
R26542 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t28 4.8295
R26543 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t9 4.8295
R26544 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t25 4.5005
R26545 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t20 4.5005
R26546 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t31 4.5005
R26547 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t24 4.5005
R26548 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t23 4.5005
R26549 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t17 4.5005
R26550 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t16 4.5005
R26551 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t10 4.5005
R26552 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t29 4.5005
R26553 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t21 4.5005
R26554 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t15 4.5005
R26555 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n4 4.5005
R26556 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n2 2.2095
R26557 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n3 2.0005
R26558 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n9 1.813
R26559 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n7 1.3755
R26560 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n1 0.8935
R26561 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 1057.5
R26562 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 1057.5
R26563 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t6 525.38
R26564 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t8 525.38
R26565 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t9 525.38
R26566 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t3 525.38
R26567 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t5 281.168
R26568 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t2 281.168
R26569 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t4 281.168
R26570 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t7 281.168
R26571 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 244.214
R26572 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 244.214
R26573 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t1 119.004
R26574 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 119.004
R26575 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 21.1255
R26576 VIN-.n0 VIN-.t9 1097.62
R26577 VIN- VIN-.n9 433.019
R26578 VIN-.n9 VIN-.t1 273.134
R26579 VIN-.n0 VIN-.t0 273.134
R26580 VIN-.n1 VIN-.t5 273.134
R26581 VIN-.n2 VIN-.t10 273.134
R26582 VIN-.n3 VIN-.t3 273.134
R26583 VIN-.n4 VIN-.t7 273.134
R26584 VIN-.n5 VIN-.t4 273.134
R26585 VIN-.n6 VIN-.t8 273.134
R26586 VIN-.n7 VIN-.t2 273.134
R26587 VIN-.n8 VIN-.t6 273.134
R26588 VIN-.n9 VIN-.n8 176.733
R26589 VIN-.n8 VIN-.n7 176.733
R26590 VIN-.n7 VIN-.n6 176.733
R26591 VIN-.n6 VIN-.n5 176.733
R26592 VIN-.n5 VIN-.n4 176.733
R26593 VIN-.n4 VIN-.n3 176.733
R26594 VIN-.n3 VIN-.n2 176.733
R26595 VIN-.n2 VIN-.n1 176.733
R26596 VIN-.n1 VIN-.n0 176.733
R26597 two_stage_opamp_dummy_magic_24_0.VD1.n15 two_stage_opamp_dummy_magic_24_0.VD1.n14 49.3505
R26598 two_stage_opamp_dummy_magic_24_0.VD1.n18 two_stage_opamp_dummy_magic_24_0.VD1.n17 49.3505
R26599 two_stage_opamp_dummy_magic_24_0.VD1.n4 two_stage_opamp_dummy_magic_24_0.VD1.n3 49.3505
R26600 two_stage_opamp_dummy_magic_24_0.VD1.n43 two_stage_opamp_dummy_magic_24_0.VD1.n42 49.3505
R26601 two_stage_opamp_dummy_magic_24_0.VD1.n39 two_stage_opamp_dummy_magic_24_0.VD1.n38 49.3505
R26602 two_stage_opamp_dummy_magic_24_0.VD1.n9 two_stage_opamp_dummy_magic_24_0.VD1.n8 49.3505
R26603 two_stage_opamp_dummy_magic_24_0.VD1.n12 two_stage_opamp_dummy_magic_24_0.VD1.n11 49.3505
R26604 two_stage_opamp_dummy_magic_24_0.VD1.n25 two_stage_opamp_dummy_magic_24_0.VD1.n24 49.3505
R26605 two_stage_opamp_dummy_magic_24_0.VD1.n28 two_stage_opamp_dummy_magic_24_0.VD1.n27 49.3505
R26606 two_stage_opamp_dummy_magic_24_0.VD1.n32 two_stage_opamp_dummy_magic_24_0.VD1.n31 49.3505
R26607 two_stage_opamp_dummy_magic_24_0.VD1.n7 two_stage_opamp_dummy_magic_24_0.VD1.n6 49.3505
R26608 two_stage_opamp_dummy_magic_24_0.VD1.n14 two_stage_opamp_dummy_magic_24_0.VD1.t11 16.0005
R26609 two_stage_opamp_dummy_magic_24_0.VD1.n14 two_stage_opamp_dummy_magic_24_0.VD1.t8 16.0005
R26610 two_stage_opamp_dummy_magic_24_0.VD1.n17 two_stage_opamp_dummy_magic_24_0.VD1.t3 16.0005
R26611 two_stage_opamp_dummy_magic_24_0.VD1.n17 two_stage_opamp_dummy_magic_24_0.VD1.t7 16.0005
R26612 two_stage_opamp_dummy_magic_24_0.VD1.n3 two_stage_opamp_dummy_magic_24_0.VD1.t1 16.0005
R26613 two_stage_opamp_dummy_magic_24_0.VD1.n3 two_stage_opamp_dummy_magic_24_0.VD1.t5 16.0005
R26614 two_stage_opamp_dummy_magic_24_0.VD1.n42 two_stage_opamp_dummy_magic_24_0.VD1.t2 16.0005
R26615 two_stage_opamp_dummy_magic_24_0.VD1.n42 two_stage_opamp_dummy_magic_24_0.VD1.t6 16.0005
R26616 two_stage_opamp_dummy_magic_24_0.VD1.n38 two_stage_opamp_dummy_magic_24_0.VD1.t0 16.0005
R26617 two_stage_opamp_dummy_magic_24_0.VD1.n38 two_stage_opamp_dummy_magic_24_0.VD1.t4 16.0005
R26618 two_stage_opamp_dummy_magic_24_0.VD1.n8 two_stage_opamp_dummy_magic_24_0.VD1.t12 16.0005
R26619 two_stage_opamp_dummy_magic_24_0.VD1.n8 two_stage_opamp_dummy_magic_24_0.VD1.t17 16.0005
R26620 two_stage_opamp_dummy_magic_24_0.VD1.n11 two_stage_opamp_dummy_magic_24_0.VD1.t16 16.0005
R26621 two_stage_opamp_dummy_magic_24_0.VD1.n11 two_stage_opamp_dummy_magic_24_0.VD1.t21 16.0005
R26622 two_stage_opamp_dummy_magic_24_0.VD1.n24 two_stage_opamp_dummy_magic_24_0.VD1.t15 16.0005
R26623 two_stage_opamp_dummy_magic_24_0.VD1.n24 two_stage_opamp_dummy_magic_24_0.VD1.t19 16.0005
R26624 two_stage_opamp_dummy_magic_24_0.VD1.n27 two_stage_opamp_dummy_magic_24_0.VD1.t13 16.0005
R26625 two_stage_opamp_dummy_magic_24_0.VD1.n27 two_stage_opamp_dummy_magic_24_0.VD1.t20 16.0005
R26626 two_stage_opamp_dummy_magic_24_0.VD1.n31 two_stage_opamp_dummy_magic_24_0.VD1.t14 16.0005
R26627 two_stage_opamp_dummy_magic_24_0.VD1.n31 two_stage_opamp_dummy_magic_24_0.VD1.t18 16.0005
R26628 two_stage_opamp_dummy_magic_24_0.VD1.n6 two_stage_opamp_dummy_magic_24_0.VD1.t9 16.0005
R26629 two_stage_opamp_dummy_magic_24_0.VD1.n6 two_stage_opamp_dummy_magic_24_0.VD1.t10 16.0005
R26630 two_stage_opamp_dummy_magic_24_0.VD1.n23 two_stage_opamp_dummy_magic_24_0.VD1.n13 5.8755
R26631 two_stage_opamp_dummy_magic_24_0.VD1.n33 two_stage_opamp_dummy_magic_24_0.VD1.n2 5.8755
R26632 two_stage_opamp_dummy_magic_24_0.VD1.n21 two_stage_opamp_dummy_magic_24_0.VD1.n20 5.8755
R26633 two_stage_opamp_dummy_magic_24_0.VD1.n36 two_stage_opamp_dummy_magic_24_0.VD1.n35 5.8755
R26634 two_stage_opamp_dummy_magic_24_0.VD1.n26 two_stage_opamp_dummy_magic_24_0.VD1.n12 5.6255
R26635 two_stage_opamp_dummy_magic_24_0.VD1.n30 two_stage_opamp_dummy_magic_24_0.VD1.n9 5.6255
R26636 two_stage_opamp_dummy_magic_24_0.VD1.n16 two_stage_opamp_dummy_magic_24_0.VD1.n15 5.438
R26637 two_stage_opamp_dummy_magic_24_0.VD1.n40 two_stage_opamp_dummy_magic_24_0.VD1.n7 5.438
R26638 two_stage_opamp_dummy_magic_24_0.VD1.n36 two_stage_opamp_dummy_magic_24_0.VD1.n7 5.31821
R26639 two_stage_opamp_dummy_magic_24_0.VD1.n20 two_stage_opamp_dummy_magic_24_0.VD1.n15 5.31821
R26640 two_stage_opamp_dummy_magic_24_0.VD1.n19 two_stage_opamp_dummy_magic_24_0.VD1.n18 5.08383
R26641 two_stage_opamp_dummy_magic_24_0.VD1.n4 two_stage_opamp_dummy_magic_24_0.VD1.n1 5.08383
R26642 two_stage_opamp_dummy_magic_24_0.VD1.n44 two_stage_opamp_dummy_magic_24_0.VD1.n43 5.08383
R26643 two_stage_opamp_dummy_magic_24_0.VD1.n39 two_stage_opamp_dummy_magic_24_0.VD1.n37 5.08383
R26644 two_stage_opamp_dummy_magic_24_0.VD1.n26 two_stage_opamp_dummy_magic_24_0.VD1.n25 5.063
R26645 two_stage_opamp_dummy_magic_24_0.VD1.n29 two_stage_opamp_dummy_magic_24_0.VD1.n28 5.063
R26646 two_stage_opamp_dummy_magic_24_0.VD1.n32 two_stage_opamp_dummy_magic_24_0.VD1.n30 5.063
R26647 two_stage_opamp_dummy_magic_24_0.VD1.n35 two_stage_opamp_dummy_magic_24_0.VD1.n34 5.063
R26648 two_stage_opamp_dummy_magic_24_0.VD1.n22 two_stage_opamp_dummy_magic_24_0.VD1.n21 5.063
R26649 two_stage_opamp_dummy_magic_24_0.VD1.n18 two_stage_opamp_dummy_magic_24_0.VD1.n16 4.8755
R26650 two_stage_opamp_dummy_magic_24_0.VD1.n5 two_stage_opamp_dummy_magic_24_0.VD1.n4 4.8755
R26651 two_stage_opamp_dummy_magic_24_0.VD1.n43 two_stage_opamp_dummy_magic_24_0.VD1.n41 4.8755
R26652 two_stage_opamp_dummy_magic_24_0.VD1.n40 two_stage_opamp_dummy_magic_24_0.VD1.n39 4.8755
R26653 two_stage_opamp_dummy_magic_24_0.VD1 two_stage_opamp_dummy_magic_24_0.VD1.n45 4.60467
R26654 two_stage_opamp_dummy_magic_24_0.VD1.n34 two_stage_opamp_dummy_magic_24_0.VD1.n33 4.5005
R26655 two_stage_opamp_dummy_magic_24_0.VD1.n10 two_stage_opamp_dummy_magic_24_0.VD1.n0 4.5005
R26656 two_stage_opamp_dummy_magic_24_0.VD1.n23 two_stage_opamp_dummy_magic_24_0.VD1.n22 4.5005
R26657 two_stage_opamp_dummy_magic_24_0.VD1 two_stage_opamp_dummy_magic_24_0.VD1.n0 1.27133
R26658 two_stage_opamp_dummy_magic_24_0.VD1.n34 two_stage_opamp_dummy_magic_24_0.VD1.n10 0.563
R26659 two_stage_opamp_dummy_magic_24_0.VD1.n22 two_stage_opamp_dummy_magic_24_0.VD1.n10 0.563
R26660 two_stage_opamp_dummy_magic_24_0.VD1.n29 two_stage_opamp_dummy_magic_24_0.VD1.n26 0.563
R26661 two_stage_opamp_dummy_magic_24_0.VD1.n30 two_stage_opamp_dummy_magic_24_0.VD1.n29 0.563
R26662 two_stage_opamp_dummy_magic_24_0.VD1.n16 two_stage_opamp_dummy_magic_24_0.VD1.n5 0.563
R26663 two_stage_opamp_dummy_magic_24_0.VD1.n41 two_stage_opamp_dummy_magic_24_0.VD1.n5 0.563
R26664 two_stage_opamp_dummy_magic_24_0.VD1.n41 two_stage_opamp_dummy_magic_24_0.VD1.n40 0.563
R26665 two_stage_opamp_dummy_magic_24_0.VD1.n25 two_stage_opamp_dummy_magic_24_0.VD1.n23 0.3755
R26666 two_stage_opamp_dummy_magic_24_0.VD1.n28 two_stage_opamp_dummy_magic_24_0.VD1.n0 0.3755
R26667 two_stage_opamp_dummy_magic_24_0.VD1.n33 two_stage_opamp_dummy_magic_24_0.VD1.n32 0.3755
R26668 two_stage_opamp_dummy_magic_24_0.VD1.n21 two_stage_opamp_dummy_magic_24_0.VD1.n12 0.3755
R26669 two_stage_opamp_dummy_magic_24_0.VD1.n35 two_stage_opamp_dummy_magic_24_0.VD1.n9 0.3755
R26670 two_stage_opamp_dummy_magic_24_0.VD1.n37 two_stage_opamp_dummy_magic_24_0.VD1.n36 0.234875
R26671 two_stage_opamp_dummy_magic_24_0.VD1.n37 two_stage_opamp_dummy_magic_24_0.VD1.n2 0.234875
R26672 two_stage_opamp_dummy_magic_24_0.VD1.n44 two_stage_opamp_dummy_magic_24_0.VD1.n2 0.234875
R26673 two_stage_opamp_dummy_magic_24_0.VD1.n45 two_stage_opamp_dummy_magic_24_0.VD1.n44 0.234875
R26674 two_stage_opamp_dummy_magic_24_0.VD1.n45 two_stage_opamp_dummy_magic_24_0.VD1.n1 0.234875
R26675 two_stage_opamp_dummy_magic_24_0.VD1.n13 two_stage_opamp_dummy_magic_24_0.VD1.n1 0.234875
R26676 two_stage_opamp_dummy_magic_24_0.VD1.n19 two_stage_opamp_dummy_magic_24_0.VD1.n13 0.234875
R26677 two_stage_opamp_dummy_magic_24_0.VD1.n20 two_stage_opamp_dummy_magic_24_0.VD1.n19 0.234875
R26678 two_stage_opamp_dummy_magic_24_0.V_tot.n2 two_stage_opamp_dummy_magic_24_0.V_tot.t4 648.28
R26679 two_stage_opamp_dummy_magic_24_0.V_tot.n1 two_stage_opamp_dummy_magic_24_0.V_tot.t5 648.28
R26680 two_stage_opamp_dummy_magic_24_0.V_tot.n0 two_stage_opamp_dummy_magic_24_0.V_tot.t1 117.591
R26681 two_stage_opamp_dummy_magic_24_0.V_tot.t0 two_stage_opamp_dummy_magic_24_0.V_tot.n3 117.591
R26682 two_stage_opamp_dummy_magic_24_0.V_tot.n3 two_stage_opamp_dummy_magic_24_0.V_tot.t3 108.424
R26683 two_stage_opamp_dummy_magic_24_0.V_tot.n0 two_stage_opamp_dummy_magic_24_0.V_tot.t2 108.424
R26684 two_stage_opamp_dummy_magic_24_0.V_tot.n1 two_stage_opamp_dummy_magic_24_0.V_tot.n0 38.5809
R26685 two_stage_opamp_dummy_magic_24_0.V_tot.n3 two_stage_opamp_dummy_magic_24_0.V_tot.n2 38.5809
R26686 two_stage_opamp_dummy_magic_24_0.V_tot.n2 two_stage_opamp_dummy_magic_24_0.V_tot.n1 1.563
R26687 two_stage_opamp_dummy_magic_24_0.V_err_mir_p two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n0 187.315
R26688 two_stage_opamp_dummy_magic_24_0.V_err_mir_p two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n1 177.755
R26689 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t3 15.7605
R26690 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t1 15.7605
R26691 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t2 15.7605
R26692 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t0 15.7605
R26693 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R26694 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R26695 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 175.56
R26696 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 168.936
R26697 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 166.925
R26698 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t1 130.001
R26699 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t0 81.7074
R26700 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.3864
R26701 bgr_11_0.START_UP bgr_11_0.START_UP.n5 14.938
R26702 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t2 13.1338
R26703 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t4 13.1338
R26704 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t3 13.1338
R26705 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t5 13.1338
R26706 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R26707 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 two_stage_opamp_dummy_magic_24_0.err_amp_out.t4 989.788
R26708 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 179.913
R26709 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 39.3422
R26710 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 two_stage_opamp_dummy_magic_24_0.err_amp_out.t1 15.7605
R26711 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 two_stage_opamp_dummy_magic_24_0.err_amp_out.t0 15.7605
R26712 two_stage_opamp_dummy_magic_24_0.err_amp_out.t2 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 9.6005
R26713 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 two_stage_opamp_dummy_magic_24_0.err_amp_out.t3 9.6005
R26714 bgr_11_0.cap_res2.t0 bgr_11_0.cap_res2.t15 121.245
R26715 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.t4 0.1603
R26716 bgr_11_0.cap_res2.t14 bgr_11_0.cap_res2.t9 0.1603
R26717 bgr_11_0.cap_res2.t8 bgr_11_0.cap_res2.t3 0.1603
R26718 bgr_11_0.cap_res2.t2 bgr_11_0.cap_res2.t16 0.1603
R26719 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.t1 0.1603
R26720 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t11 0.159278
R26721 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t7 0.159278
R26722 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t13 0.159278
R26723 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t19 0.159278
R26724 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t20 0.1368
R26725 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t10 0.1368
R26726 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t5 0.1368
R26727 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t14 0.1368
R26728 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t18 0.1368
R26729 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t8 0.1368
R26730 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t12 0.1368
R26731 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t2 0.1368
R26732 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t17 0.1368
R26733 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t6 0.1368
R26734 bgr_11_0.cap_res2.t11 bgr_11_0.cap_res2.n0 0.00152174
R26735 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.n1 0.00152174
R26736 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.n2 0.00152174
R26737 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.n3 0.00152174
R26738 bgr_11_0.cap_res2.t15 bgr_11_0.cap_res2.n4 0.00152174
R26739 VIN+.n0 VIN+.t3 1097.62
R26740 VIN+ VIN+.n9 433.019
R26741 VIN+.n9 VIN+.t9 273.134
R26742 VIN+.n0 VIN+.t0 273.134
R26743 VIN+.n8 VIN+.t5 273.134
R26744 VIN+.n7 VIN+.t8 273.134
R26745 VIN+.n6 VIN+.t4 273.134
R26746 VIN+.n5 VIN+.t7 273.134
R26747 VIN+.n4 VIN+.t1 273.134
R26748 VIN+.n3 VIN+.t10 273.134
R26749 VIN+.n2 VIN+.t2 273.134
R26750 VIN+.n1 VIN+.t6 273.134
R26751 VIN+.n1 VIN+.n0 176.733
R26752 VIN+.n2 VIN+.n1 176.733
R26753 VIN+.n3 VIN+.n2 176.733
R26754 VIN+.n4 VIN+.n3 176.733
R26755 VIN+.n5 VIN+.n4 176.733
R26756 VIN+.n6 VIN+.n5 176.733
R26757 VIN+.n7 VIN+.n6 176.733
R26758 VIN+.n8 VIN+.n7 176.733
R26759 VIN+.n9 VIN+.n8 176.733
R26760 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 528.612
R26761 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.n1 168.435
R26762 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 168.435
R26763 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t0 156.141
R26764 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t1 115.74
R26765 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.n0 22.5317
R26766 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 17.4224
R26767 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t2 13.1338
R26768 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t5 13.1338
R26769 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.t4 13.1338
R26770 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.t3 13.1338
R26771 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n2 1.1255
R26772 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.n15 325.473
R26773 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.n8 325.473
R26774 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.n3 325.473
R26775 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t17 310.488
R26776 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t18 310.488
R26777 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t13 310.488
R26778 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.t11 184.097
R26779 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.t9 184.097
R26780 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.t7 184.097
R26781 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.n12 167.094
R26782 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.n5 167.094
R26783 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.n0 167.094
R26784 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.n7 152
R26785 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.n2 152
R26786 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n14 152
R26787 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t14 120.501
R26788 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.t3 120.501
R26789 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t16 120.501
R26790 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.t5 120.501
R26791 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t15 120.501
R26792 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.t1 120.501
R26793 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.t0 106.933
R26794 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.n13 40.7027
R26795 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.n6 40.7027
R26796 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.n1 40.7027
R26797 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.t6 39.4005
R26798 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.t10 39.4005
R26799 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.t2 39.4005
R26800 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.t8 39.4005
R26801 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.t4 39.4005
R26802 bgr_11_0.V_mir2.t12 bgr_11_0.V_mir2.n16 39.4005
R26803 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n4 15.9255
R26804 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n11 15.9255
R26805 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.n9 9.3005
R26806 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n10 4.5005
R26807 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.t8 539.803
R26808 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n5 351.522
R26809 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n2 173.029
R26810 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n3 168.654
R26811 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t0 118.442
R26812 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n11 83.5719
R26813 bgr_11_0.Vin-.n1 bgr_11_0.Vin-.n0 83.5719
R26814 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n1 73.8495
R26815 bgr_11_0.Vin-.t7 bgr_11_0.Vin-.n10 65.0341
R26816 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.t2 39.4005
R26817 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.t1 39.4005
R26818 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 28.1567
R26819 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n1 26.074
R26820 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 16.188
R26821 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t4 13.1338
R26822 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t5 13.1338
R26823 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.t6 13.1338
R26824 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.t3 13.1338
R26825 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 11.8755
R26826 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n4 3.8755
R26827 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n10 1.56483
R26828 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 1.5505
R26829 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n0 0.885803
R26830 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 0.77514
R26831 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R26832 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 0.711459
R26833 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n15 0.576566
R26834 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 0.531499
R26835 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t7 0.290206
R26836 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n9 0.00817857
R26837 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t2 99.353
R26838 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t1 9.6005
R26839 bgr_11_0.V_p_1.t0 bgr_11_0.V_p_1.n0 9.6005
R26840 a_11300_28850.t0 a_11300_28850.t1 178.133
R26841 a_4100_3858.t0 a_4100_3858.t1 294.339
R26842 a_13390_346.t0 a_13390_346.t1 169.905
R26843 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t5 661.375
R26844 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t2 661.375
R26845 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n6 213.131
R26846 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t6 213.131
R26847 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t3 146.155
R26848 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t0 146.155
R26849 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t4 76.2576
R26850 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n7 76.2576
R26851 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n1 72.4424
R26852 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n2 66.4532
R26853 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t1 11.2576
R26854 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t7 11.2576
R26855 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t10 11.2576
R26856 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t9 11.2576
R26857 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n4 5.1255
R26858 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n3 4.9096
R26859 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n0 4.7505
R26860 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n5 1.888
R26861 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n0 1.888
R26862 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 345.264
R26863 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 344.7
R26864 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 292.5
R26865 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t4 121.849
R26866 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 118.861
R26867 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 118.861
R26868 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 118.861
R26869 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 118.861
R26870 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 118.861
R26871 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 75.063
R26872 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 52.763
R26873 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 51.7297
R26874 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t0 39.4005
R26875 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t6 39.4005
R26876 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t3 39.4005
R26877 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t2 39.4005
R26878 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t5 39.4005
R26879 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t1 39.4005
R26880 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t15 19.7005
R26881 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t11 19.7005
R26882 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t16 19.7005
R26883 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t10 19.7005
R26884 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t14 19.7005
R26885 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t9 19.7005
R26886 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t13 19.7005
R26887 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t8 19.7005
R26888 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t12 19.7005
R26889 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t7 19.7005
R26890 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 5.938
R26891 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 5.60467
R26892 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 5.54217
R26893 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 5.54217
R26894 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 5.04217
R26895 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 5.04217
R26896 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 5.04217
R26897 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 5.04217
R26898 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 4.97967
R26899 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 4.97967
R26900 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 4.97967
R26901 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 0.563
R26902 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 0.563
R26903 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 0.563
R26904 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 0.563
R26905 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 0.563
R26906 a_5700_30308.t0 a_5700_30308.t1 178.133
R26907 a_5820_29044.t0 a_5820_29044.t1 178.133
R26908 a_13550_3858.t0 a_13550_3858.t1 169.905
R26909 two_stage_opamp_dummy_magic_24_0.V_p_mir.n1 two_stage_opamp_dummy_magic_24_0.V_p_mir.n0 89.9957
R26910 two_stage_opamp_dummy_magic_24_0.V_p_mir.n0 two_stage_opamp_dummy_magic_24_0.V_p_mir.t0 16.0005
R26911 two_stage_opamp_dummy_magic_24_0.V_p_mir.n0 two_stage_opamp_dummy_magic_24_0.V_p_mir.t3 16.0005
R26912 two_stage_opamp_dummy_magic_24_0.V_p_mir.n1 two_stage_opamp_dummy_magic_24_0.V_p_mir.t1 9.6005
R26913 two_stage_opamp_dummy_magic_24_0.V_p_mir.t2 two_stage_opamp_dummy_magic_24_0.V_p_mir.n1 9.6005
R26914 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 200.749
R26915 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t1 9.6005
R26916 bgr_11_0.V_p_2.t0 bgr_11_0.V_p_2.n0 9.6005
R26917 a_6350_30458.t0 a_6350_30458.t1 178.133
R26918 a_6470_28850.t0 a_6470_28850.t1 178.133
R26919 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 two_stage_opamp_dummy_magic_24_0.Vb1_2.t0 65.3505
R26920 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 49.3505
R26921 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 49.3505
R26922 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 two_stage_opamp_dummy_magic_24_0.Vb1_2.t2 16.0005
R26923 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 two_stage_opamp_dummy_magic_24_0.Vb1_2.t4 16.0005
R26924 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 two_stage_opamp_dummy_magic_24_0.Vb1_2.t1 16.0005
R26925 two_stage_opamp_dummy_magic_24_0.Vb1_2.t3 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 16.0005
R26926 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 6.3755
R26927 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 6.1255
R26928 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 5.688
R26929 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 5.438
R26930 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 5.1255
R26931 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 4.8755
R26932 a_12070_30308.t0 a_12070_30308.t1 178.133
R26933 a_11950_29100.t0 a_11950_29100.t1 178.133
R26934 two_stage_opamp_dummy_magic_24_0.V_err_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_p.n0 365.07
R26935 two_stage_opamp_dummy_magic_24_0.V_err_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_p.t1 15.7605
R26936 two_stage_opamp_dummy_magic_24_0.V_err_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_p.t3 15.7605
R26937 two_stage_opamp_dummy_magic_24_0.V_err_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_p.t0 15.7605
R26938 two_stage_opamp_dummy_magic_24_0.V_err_p.t2 two_stage_opamp_dummy_magic_24_0.V_err_p.n1 15.7605
R26939 a_11420_30458.t0 a_11420_30458.t1 178.133
R26940 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t3 536.909
R26941 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 371.678
R26942 bgr_11_0.V_CUR_REF_REG.t1 bgr_11_0.V_CUR_REF_REG.n1 151.849
R26943 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t0 39.4005
R26944 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R26945 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R26946 a_4220_3858.t0 a_4220_3858.t1 169.905
C0 bgr_11_0.START_UP_NFET1 VDDA 0.378868f
C1 bgr_11_0.PFET_GATE_10uA VDDA 8.25933f
C2 VDDA VOUT+ 15.1488f
C3 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.019707f
C4 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.V_TOP 0.581096f
C5 two_stage_opamp_dummy_magic_24_0.V_source VDDA 0.010606f
C6 VDDA VOUT- 15.152599f
C7 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_mir_p 0.429395f
C8 two_stage_opamp_dummy_magic_24_0.cap_res_Y VDDA 7.74732f
C9 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_gate 0.80454f
C10 two_stage_opamp_dummy_magic_24_0.X VDDA 6.31959f
C11 two_stage_opamp_dummy_magic_24_0.Y VDDA 5.6772f
C12 two_stage_opamp_dummy_magic_24_0.VD1 two_stage_opamp_dummy_magic_24_0.V_source 5.04286f
C13 bgr_11_0.1st_Vout_1 VDDA 1.384f
C14 two_stage_opamp_dummy_magic_24_0.VD2 two_stage_opamp_dummy_magic_24_0.V_source 5.0406f
C15 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.START_UP 1.36559f
C16 VOUT+ VOUT- 0.305434f
C17 two_stage_opamp_dummy_magic_24_0.cap_res_Y VOUT+ 51.283f
C18 two_stage_opamp_dummy_magic_24_0.V_tail_gate VDDA 8.50828f
C19 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.VD1 6.05003f
C20 two_stage_opamp_dummy_magic_24_0.Y VOUT+ 4.16524f
C21 bgr_11_0.Vin+ VDDA 1.43659f
C22 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.VD2 6.19572f
C23 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.576305f
C24 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_mir_p 0.047303f
C25 two_stage_opamp_dummy_magic_24_0.cap_res_Y VOUT- 0.028842f
C26 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.VD1 0.017519f
C27 two_stage_opamp_dummy_magic_24_0.V_tail_gate VOUT+ 2.21052f
C28 two_stage_opamp_dummy_magic_24_0.VD2 VIN+ 0.532981f
C29 two_stage_opamp_dummy_magic_24_0.X VOUT- 4.1657f
C30 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.VD2 0.018539f
C31 two_stage_opamp_dummy_magic_24_0.V_source VIN+ 0.525732f
C32 bgr_11_0.PFET_GATE_10uA bgr_11_0.Vin+ 0.294564f
C33 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.cap_res_Y 0.08087f
C34 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_source 3.97214f
C35 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.X 0.063916f
C36 two_stage_opamp_dummy_magic_24_0.VD1 VIN- 0.532981f
C37 bgr_11_0.V_TOP VDDA 14.430401f
C38 two_stage_opamp_dummy_magic_24_0.V_tail_gate VOUT- 2.21048f
C39 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.cap_res_Y 5.64371f
C40 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C41 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.X 0.033547f
C42 two_stage_opamp_dummy_magic_24_0.V_source VIN- 0.526626f
C43 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.Y 0.033068f
C44 two_stage_opamp_dummy_magic_24_0.V_err_gate VDDA 2.96245f
C45 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.211226f
C46 two_stage_opamp_dummy_magic_24_0.V_tail_gate VIN+ 0.063737f
C47 bgr_11_0.Vin+ bgr_11_0.1st_Vout_1 0.172624f
C48 bgr_11_0.START_UP VDDA 1.50797f
C49 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C50 VIN+ VIN- 0.075694f
C51 two_stage_opamp_dummy_magic_24_0.V_tail_gate VIN- 0.060623f
C52 two_stage_opamp_dummy_magic_24_0.V_err_mir_p VDDA 0.671298f
C53 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref VDDA 2.76164f
C54 bgr_11_0.V_TOP bgr_11_0.1st_Vout_1 2.44008f
C55 two_stage_opamp_dummy_magic_24_0.V_err_gate VOUT- 0.033453f
C56 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.X 0.201432f
C57 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.Y 0.019251f
C58 two_stage_opamp_dummy_magic_24_0.V_err_gate bgr_11_0.1st_Vout_1 0.040807f
C59 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_24_0.V_err_amp_ref 1.65222f
C60 bgr_11_0.Vin+ bgr_11_0.V_TOP 1.10602f
C61 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref VOUT+ 0.032828f
C62 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.169248f
C63 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.895203f
C64 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.040465f
C65 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.cap_res_Y 0.222453f
C66 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.X 0.010979f
C67 bgr_11_0.Vin+ bgr_11_0.START_UP 0.407102f
C68 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.V_err_mir_p 0.026615f
C69 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.Y 0.218439f
C70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.055802f
C71 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_24_0.V_err_gate 0.08574f
C72 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.138416f
C73 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.Vin+ 3.11453f
C74 bgr_11_0.V_TOP bgr_11_0.START_UP 0.746692f
C75 VIN- GNDA 1.81825f
C76 VIN+ GNDA 1.8149f
C77 VOUT- GNDA 22.797924f
C78 VOUT+ GNDA 22.816366f
C79 VDDA GNDA 0.482204p
C80 two_stage_opamp_dummy_magic_24_0.V_source GNDA 16.871408f
C81 two_stage_opamp_dummy_magic_24_0.VD1 GNDA 2.618378f
C82 two_stage_opamp_dummy_magic_24_0.VD2 GNDA 2.234519f
C83 two_stage_opamp_dummy_magic_24_0.V_err_mir_p GNDA 0.099889f
C84 two_stage_opamp_dummy_magic_24_0.cap_res_Y GNDA 37.32978f
C85 two_stage_opamp_dummy_magic_24_0.X GNDA 10.345821f
C86 two_stage_opamp_dummy_magic_24_0.Y GNDA 9.788177f
C87 two_stage_opamp_dummy_magic_24_0.V_tail_gate GNDA 29.262648f
C88 bgr_11_0.1st_Vout_1 GNDA 7.197568f
C89 bgr_11_0.START_UP GNDA 6.096303f
C90 bgr_11_0.START_UP_NFET1 GNDA 4.52649f
C91 two_stage_opamp_dummy_magic_24_0.V_err_gate GNDA 11.29427f
C92 bgr_11_0.V_TOP GNDA 9.923664f
C93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.6726f
C94 bgr_11_0.Vin+ GNDA 4.730191f
C95 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref GNDA 8.255939f
C96 bgr_11_0.PFET_GATE_10uA GNDA 7.532079f
C97 bgr_11_0.V_CUR_REF_REG.n0 GNDA 0.065451f
C98 bgr_11_0.V_CUR_REF_REG.t3 GNDA 0.045935f
C99 bgr_11_0.V_CUR_REF_REG.n1 GNDA 2.00566f
C100 bgr_11_0.V_CUR_REF_REG.t1 GNDA 0.264844f
C101 two_stage_opamp_dummy_magic_24_0.Vb1_2.t1 GNDA 0.047649f
C102 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 GNDA 0.318351f
C103 two_stage_opamp_dummy_magic_24_0.Vb1_2.t0 GNDA 0.161927f
C104 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 GNDA 0.491746f
C105 two_stage_opamp_dummy_magic_24_0.Vb1_2.t2 GNDA 0.047649f
C106 two_stage_opamp_dummy_magic_24_0.Vb1_2.t4 GNDA 0.047649f
C107 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 GNDA 0.103679f
C108 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 GNDA 0.407675f
C109 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 GNDA 0.297965f
C110 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 GNDA 0.42438f
C111 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 GNDA 0.103679f
C112 two_stage_opamp_dummy_magic_24_0.Vb1_2.t3 GNDA 0.047649f
C113 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t5 GNDA 0.020037f
C114 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t1 GNDA 0.020037f
C115 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 GNDA 0.050247f
C116 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t3 GNDA 0.020037f
C117 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t2 GNDA 0.020037f
C118 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 GNDA 0.049983f
C119 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 GNDA 0.444327f
C120 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t0 GNDA 0.020037f
C121 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t6 GNDA 0.020037f
C122 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 GNDA 0.040074f
C123 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 GNDA 0.07461f
C124 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t4 GNDA 0.252398f
C125 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 GNDA 0.063297f
C126 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 GNDA 0.111959f
C127 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t15 GNDA 0.040074f
C128 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t11 GNDA 0.040074f
C129 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 GNDA 0.081935f
C130 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 GNDA 0.275217f
C131 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t16 GNDA 0.040074f
C132 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t10 GNDA 0.040074f
C133 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 GNDA 0.081935f
C134 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 GNDA 0.265036f
C135 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 GNDA 0.107622f
C136 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 GNDA 0.063297f
C137 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t14 GNDA 0.040074f
C138 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t9 GNDA 0.040074f
C139 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 GNDA 0.081935f
C140 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 GNDA 0.265036f
C141 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 GNDA 0.065611f
C142 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t13 GNDA 0.040074f
C143 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t8 GNDA 0.040074f
C144 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 GNDA 0.081935f
C145 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 GNDA 0.265036f
C146 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 GNDA 0.111959f
C147 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t12 GNDA 0.040074f
C148 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t7 GNDA 0.040074f
C149 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 GNDA 0.081935f
C150 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 GNDA 0.270272f
C151 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 GNDA 0.147536f
C152 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 GNDA 2.3493f
C153 bgr_11_0.V_CMFB_S3 GNDA 2.19655f
C154 bgr_11_0.Vin-.n0 GNDA 0.077003f
C155 bgr_11_0.Vin-.n1 GNDA 0.349039f
C156 bgr_11_0.Vin-.t6 GNDA 0.02992f
C157 bgr_11_0.Vin-.t3 GNDA 0.02992f
C158 bgr_11_0.Vin-.n2 GNDA 0.104161f
C159 bgr_11_0.Vin-.t4 GNDA 0.02992f
C160 bgr_11_0.Vin-.t5 GNDA 0.02992f
C161 bgr_11_0.Vin-.n3 GNDA 0.099464f
C162 bgr_11_0.Vin-.n4 GNDA 0.426698f
C163 bgr_11_0.Vin-.n5 GNDA 0.030561f
C164 bgr_11_0.Vin-.n6 GNDA 0.411767f
C165 bgr_11_0.Vin-.t8 GNDA 0.048458f
C166 bgr_11_0.Vin-.n7 GNDA 0.589708f
C167 bgr_11_0.Vin-.t0 GNDA 0.12816f
C168 bgr_11_0.Vin-.n8 GNDA 0.693577f
C169 bgr_11_0.Vin-.n9 GNDA 1.17523f
C170 bgr_11_0.Vin-.n10 GNDA 0.520358f
C171 bgr_11_0.Vin-.t7 GNDA 0.28885f
C172 bgr_11_0.Vin-.n11 GNDA 0.077145f
C173 bgr_11_0.Vin-.n12 GNDA 0.132035f
C174 bgr_11_0.Vin-.n13 GNDA 0.077868f
C175 bgr_11_0.Vin-.n14 GNDA 0.639268f
C176 bgr_11_0.Vin-.n15 GNDA 0.395484f
C177 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.095541f
C178 bgr_11_0.Vin+.t0 GNDA 0.123845f
C179 bgr_11_0.Vin+.t1 GNDA 0.173539f
C180 bgr_11_0.Vin+.n0 GNDA 2.15533f
C181 bgr_11_0.Vin+.t2 GNDA 0.038796f
C182 bgr_11_0.Vin+.t5 GNDA 0.038796f
C183 bgr_11_0.Vin+.n1 GNDA 0.128171f
C184 bgr_11_0.Vin+.n2 GNDA 1.45471f
C185 bgr_11_0.Vin+.t4 GNDA 0.038796f
C186 bgr_11_0.Vin+.t3 GNDA 0.038796f
C187 bgr_11_0.Vin+.n3 GNDA 0.128171f
C188 bgr_11_0.Vin+.n4 GNDA 1.04273f
C189 bgr_11_0.Vin+.t6 GNDA 0.061838f
C190 bgr_11_0.cap_res2.t4 GNDA 0.358376f
C191 bgr_11_0.cap_res2.t10 GNDA 0.359675f
C192 bgr_11_0.cap_res2.t20 GNDA 0.340442f
C193 bgr_11_0.cap_res2.t9 GNDA 0.358376f
C194 bgr_11_0.cap_res2.t14 GNDA 0.359675f
C195 bgr_11_0.cap_res2.t5 GNDA 0.340442f
C196 bgr_11_0.cap_res2.t3 GNDA 0.358376f
C197 bgr_11_0.cap_res2.t8 GNDA 0.359675f
C198 bgr_11_0.cap_res2.t18 GNDA 0.340442f
C199 bgr_11_0.cap_res2.t16 GNDA 0.358376f
C200 bgr_11_0.cap_res2.t2 GNDA 0.359675f
C201 bgr_11_0.cap_res2.t12 GNDA 0.340442f
C202 bgr_11_0.cap_res2.t1 GNDA 0.358376f
C203 bgr_11_0.cap_res2.t6 GNDA 0.359675f
C204 bgr_11_0.cap_res2.t17 GNDA 0.340442f
C205 bgr_11_0.cap_res2.n0 GNDA 0.24022f
C206 bgr_11_0.cap_res2.t11 GNDA 0.1913f
C207 bgr_11_0.cap_res2.n1 GNDA 0.260644f
C208 bgr_11_0.cap_res2.t7 GNDA 0.1913f
C209 bgr_11_0.cap_res2.n2 GNDA 0.260644f
C210 bgr_11_0.cap_res2.t13 GNDA 0.1913f
C211 bgr_11_0.cap_res2.n3 GNDA 0.260644f
C212 bgr_11_0.cap_res2.t19 GNDA 0.1913f
C213 bgr_11_0.cap_res2.n4 GNDA 0.260644f
C214 bgr_11_0.cap_res2.t15 GNDA 0.373116f
C215 bgr_11_0.cap_res2.t0 GNDA 0.086426f
C216 bgr_11_0.START_UP.t0 GNDA 1.81996f
C217 bgr_11_0.START_UP.t1 GNDA 0.047842f
C218 bgr_11_0.START_UP.n0 GNDA 1.21481f
C219 bgr_11_0.START_UP.t2 GNDA 0.045656f
C220 bgr_11_0.START_UP.t4 GNDA 0.045656f
C221 bgr_11_0.START_UP.n1 GNDA 0.165632f
C222 bgr_11_0.START_UP.t3 GNDA 0.045656f
C223 bgr_11_0.START_UP.t5 GNDA 0.045656f
C224 bgr_11_0.START_UP.n2 GNDA 0.152372f
C225 bgr_11_0.START_UP.n3 GNDA 0.789149f
C226 bgr_11_0.START_UP.t6 GNDA 0.017156f
C227 bgr_11_0.START_UP.t7 GNDA 0.017156f
C228 bgr_11_0.START_UP.n4 GNDA 0.048434f
C229 bgr_11_0.START_UP.n5 GNDA 0.475003f
C230 two_stage_opamp_dummy_magic_24_0.V_tot.t3 GNDA 0.101695f
C231 two_stage_opamp_dummy_magic_24_0.V_tot.t1 GNDA 0.10833f
C232 two_stage_opamp_dummy_magic_24_0.V_tot.t2 GNDA 0.101695f
C233 two_stage_opamp_dummy_magic_24_0.V_tot.n0 GNDA 0.544778f
C234 two_stage_opamp_dummy_magic_24_0.V_tot.t5 GNDA 0.030796f
C235 two_stage_opamp_dummy_magic_24_0.V_tot.n1 GNDA 0.514402f
C236 two_stage_opamp_dummy_magic_24_0.V_tot.t4 GNDA 0.030796f
C237 two_stage_opamp_dummy_magic_24_0.V_tot.n2 GNDA 0.514402f
C238 two_stage_opamp_dummy_magic_24_0.V_tot.n3 GNDA 0.544778f
C239 two_stage_opamp_dummy_magic_24_0.V_tot.t0 GNDA 0.10833f
C240 two_stage_opamp_dummy_magic_24_0.VD1.n0 GNDA 0.224083f
C241 two_stage_opamp_dummy_magic_24_0.VD1.n1 GNDA 0.076567f
C242 two_stage_opamp_dummy_magic_24_0.VD1.n2 GNDA 0.102761f
C243 two_stage_opamp_dummy_magic_24_0.VD1.t1 GNDA 0.051027f
C244 two_stage_opamp_dummy_magic_24_0.VD1.t5 GNDA 0.051027f
C245 two_stage_opamp_dummy_magic_24_0.VD1.n3 GNDA 0.111028f
C246 two_stage_opamp_dummy_magic_24_0.VD1.n4 GNDA 0.427784f
C247 two_stage_opamp_dummy_magic_24_0.VD1.n5 GNDA 0.108519f
C248 two_stage_opamp_dummy_magic_24_0.VD1.t9 GNDA 0.051027f
C249 two_stage_opamp_dummy_magic_24_0.VD1.t10 GNDA 0.051027f
C250 two_stage_opamp_dummy_magic_24_0.VD1.n6 GNDA 0.111028f
C251 two_stage_opamp_dummy_magic_24_0.VD1.n7 GNDA 0.439712f
C252 two_stage_opamp_dummy_magic_24_0.VD1.t12 GNDA 0.051027f
C253 two_stage_opamp_dummy_magic_24_0.VD1.t17 GNDA 0.051027f
C254 two_stage_opamp_dummy_magic_24_0.VD1.n8 GNDA 0.111028f
C255 two_stage_opamp_dummy_magic_24_0.VD1.n9 GNDA 0.354798f
C256 two_stage_opamp_dummy_magic_24_0.VD1.n10 GNDA 0.102053f
C257 two_stage_opamp_dummy_magic_24_0.VD1.t16 GNDA 0.051027f
C258 two_stage_opamp_dummy_magic_24_0.VD1.t21 GNDA 0.051027f
C259 two_stage_opamp_dummy_magic_24_0.VD1.n11 GNDA 0.111028f
C260 two_stage_opamp_dummy_magic_24_0.VD1.n12 GNDA 0.354798f
C261 two_stage_opamp_dummy_magic_24_0.VD1.n13 GNDA 0.102761f
C262 two_stage_opamp_dummy_magic_24_0.VD1.t11 GNDA 0.051027f
C263 two_stage_opamp_dummy_magic_24_0.VD1.t8 GNDA 0.051027f
C264 two_stage_opamp_dummy_magic_24_0.VD1.n14 GNDA 0.111028f
C265 two_stage_opamp_dummy_magic_24_0.VD1.n15 GNDA 0.439711f
C266 two_stage_opamp_dummy_magic_24_0.VD1.n16 GNDA 0.184463f
C267 two_stage_opamp_dummy_magic_24_0.VD1.t3 GNDA 0.051027f
C268 two_stage_opamp_dummy_magic_24_0.VD1.t7 GNDA 0.051027f
C269 two_stage_opamp_dummy_magic_24_0.VD1.n17 GNDA 0.111028f
C270 two_stage_opamp_dummy_magic_24_0.VD1.n18 GNDA 0.427784f
C271 two_stage_opamp_dummy_magic_24_0.VD1.n19 GNDA 0.076567f
C272 two_stage_opamp_dummy_magic_24_0.VD1.n20 GNDA 0.171401f
C273 two_stage_opamp_dummy_magic_24_0.VD1.n21 GNDA 0.390374f
C274 two_stage_opamp_dummy_magic_24_0.VD1.n22 GNDA 0.171601f
C275 two_stage_opamp_dummy_magic_24_0.VD1.n23 GNDA 0.381681f
C276 two_stage_opamp_dummy_magic_24_0.VD1.t15 GNDA 0.051027f
C277 two_stage_opamp_dummy_magic_24_0.VD1.t19 GNDA 0.051027f
C278 two_stage_opamp_dummy_magic_24_0.VD1.n24 GNDA 0.111028f
C279 two_stage_opamp_dummy_magic_24_0.VD1.n25 GNDA 0.345781f
C280 two_stage_opamp_dummy_magic_24_0.VD1.n26 GNDA 0.195132f
C281 two_stage_opamp_dummy_magic_24_0.VD1.t13 GNDA 0.051027f
C282 two_stage_opamp_dummy_magic_24_0.VD1.t20 GNDA 0.051027f
C283 two_stage_opamp_dummy_magic_24_0.VD1.n27 GNDA 0.111028f
C284 two_stage_opamp_dummy_magic_24_0.VD1.n28 GNDA 0.345781f
C285 two_stage_opamp_dummy_magic_24_0.VD1.n29 GNDA 0.113981f
C286 two_stage_opamp_dummy_magic_24_0.VD1.n30 GNDA 0.195132f
C287 two_stage_opamp_dummy_magic_24_0.VD1.t14 GNDA 0.051027f
C288 two_stage_opamp_dummy_magic_24_0.VD1.t18 GNDA 0.051027f
C289 two_stage_opamp_dummy_magic_24_0.VD1.n31 GNDA 0.111028f
C290 two_stage_opamp_dummy_magic_24_0.VD1.n32 GNDA 0.345781f
C291 two_stage_opamp_dummy_magic_24_0.VD1.n33 GNDA 0.381681f
C292 two_stage_opamp_dummy_magic_24_0.VD1.n34 GNDA 0.171601f
C293 two_stage_opamp_dummy_magic_24_0.VD1.n35 GNDA 0.390374f
C294 two_stage_opamp_dummy_magic_24_0.VD1.n36 GNDA 0.171401f
C295 two_stage_opamp_dummy_magic_24_0.VD1.n37 GNDA 0.076567f
C296 two_stage_opamp_dummy_magic_24_0.VD1.t0 GNDA 0.051027f
C297 two_stage_opamp_dummy_magic_24_0.VD1.t4 GNDA 0.051027f
C298 two_stage_opamp_dummy_magic_24_0.VD1.n38 GNDA 0.111028f
C299 two_stage_opamp_dummy_magic_24_0.VD1.n39 GNDA 0.427784f
C300 two_stage_opamp_dummy_magic_24_0.VD1.n40 GNDA 0.184463f
C301 two_stage_opamp_dummy_magic_24_0.VD1.n41 GNDA 0.108519f
C302 two_stage_opamp_dummy_magic_24_0.VD1.t2 GNDA 0.051027f
C303 two_stage_opamp_dummy_magic_24_0.VD1.t6 GNDA 0.051027f
C304 two_stage_opamp_dummy_magic_24_0.VD1.n42 GNDA 0.111028f
C305 two_stage_opamp_dummy_magic_24_0.VD1.n43 GNDA 0.427784f
C306 two_stage_opamp_dummy_magic_24_0.VD1.n44 GNDA 0.076567f
C307 two_stage_opamp_dummy_magic_24_0.VD1.n45 GNDA 0.059261f
C308 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t1 GNDA 0.294683f
C309 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t4 GNDA 0.711146f
C310 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t7 GNDA 0.711146f
C311 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t3 GNDA 0.844019f
C312 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 GNDA 0.445804f
C313 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t9 GNDA 0.844019f
C314 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 GNDA 0.551177f
C315 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 GNDA 1.59801f
C316 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t5 GNDA 0.711146f
C317 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t8 GNDA 0.844019f
C318 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t2 GNDA 0.711146f
C319 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t6 GNDA 0.844019f
C320 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 GNDA 0.445804f
C321 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 GNDA 0.551177f
C322 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 GNDA 1.59801f
C323 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t0 GNDA 0.294683f
C324 bgr_11_0.1st_Vout_2.n0 GNDA 1.42188f
C325 bgr_11_0.1st_Vout_2.n1 GNDA 0.433567f
C326 bgr_11_0.1st_Vout_2.n2 GNDA 0.97351f
C327 bgr_11_0.1st_Vout_2.n3 GNDA 0.150653f
C328 bgr_11_0.1st_Vout_2.n4 GNDA 0.097613f
C329 bgr_11_0.1st_Vout_2.n5 GNDA 0.017136f
C330 bgr_11_0.1st_Vout_2.t7 GNDA 0.01702f
C331 bgr_11_0.1st_Vout_2.n6 GNDA 0.017877f
C332 bgr_11_0.1st_Vout_2.n7 GNDA 0.136013f
C333 bgr_11_0.1st_Vout_2.t26 GNDA 0.010803f
C334 bgr_11_0.1st_Vout_2.t14 GNDA 0.010803f
C335 bgr_11_0.1st_Vout_2.n8 GNDA 0.024033f
C336 bgr_11_0.1st_Vout_2.t29 GNDA 0.283668f
C337 bgr_11_0.1st_Vout_2.t32 GNDA 0.288499f
C338 bgr_11_0.1st_Vout_2.t25 GNDA 0.283668f
C339 bgr_11_0.1st_Vout_2.t20 GNDA 0.283668f
C340 bgr_11_0.1st_Vout_2.t12 GNDA 0.288499f
C341 bgr_11_0.1st_Vout_2.t13 GNDA 0.288499f
C342 bgr_11_0.1st_Vout_2.t31 GNDA 0.283668f
C343 bgr_11_0.1st_Vout_2.t24 GNDA 0.283668f
C344 bgr_11_0.1st_Vout_2.t18 GNDA 0.288499f
C345 bgr_11_0.1st_Vout_2.t30 GNDA 0.288499f
C346 bgr_11_0.1st_Vout_2.t23 GNDA 0.283668f
C347 bgr_11_0.1st_Vout_2.t17 GNDA 0.283668f
C348 bgr_11_0.1st_Vout_2.t11 GNDA 0.288499f
C349 bgr_11_0.1st_Vout_2.t22 GNDA 0.288499f
C350 bgr_11_0.1st_Vout_2.t16 GNDA 0.283668f
C351 bgr_11_0.1st_Vout_2.t10 GNDA 0.283668f
C352 bgr_11_0.1st_Vout_2.t28 GNDA 0.288499f
C353 bgr_11_0.1st_Vout_2.t9 GNDA 0.288499f
C354 bgr_11_0.1st_Vout_2.t15 GNDA 0.283668f
C355 bgr_11_0.1st_Vout_2.t21 GNDA 0.283668f
C356 bgr_11_0.1st_Vout_2.t8 GNDA 0.018531f
C357 bgr_11_0.1st_Vout_2.n9 GNDA 0.547784f
C358 bgr_11_0.1st_Vout_2.n10 GNDA 0.017877f
C359 bgr_11_0.1st_Vout_2.t27 GNDA 0.010803f
C360 bgr_11_0.1st_Vout_2.t19 GNDA 0.010803f
C361 bgr_11_0.1st_Vout_2.n11 GNDA 0.024033f
C362 bgr_11_0.1st_Vout_2.n12 GNDA 0.103502f
C363 bgr_11_0.1st_Vout_2.t4 GNDA 0.096368f
C364 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t11 GNDA 0.020261f
C365 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t14 GNDA 0.020261f
C366 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 GNDA 0.050788f
C367 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t10 GNDA 0.020261f
C368 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t13 GNDA 0.020261f
C369 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 GNDA 0.05052f
C370 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 GNDA 0.449015f
C371 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t15 GNDA 0.020261f
C372 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t12 GNDA 0.020261f
C373 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 GNDA 0.040522f
C374 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 GNDA 0.075475f
C375 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t16 GNDA 0.255451f
C376 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 GNDA 0.064004f
C377 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 GNDA 0.113211f
C378 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t6 GNDA 0.040522f
C379 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t5 GNDA 0.040522f
C380 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 GNDA 0.082851f
C381 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 GNDA 0.278294f
C382 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t8 GNDA 0.040522f
C383 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t1 GNDA 0.040522f
C384 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 GNDA 0.082851f
C385 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 GNDA 0.267999f
C386 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 GNDA 0.108825f
C387 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 GNDA 0.064004f
C388 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t9 GNDA 0.040522f
C389 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t3 GNDA 0.040522f
C390 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 GNDA 0.082851f
C391 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 GNDA 0.267999f
C392 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 GNDA 0.066344f
C393 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t0 GNDA 0.040522f
C394 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t4 GNDA 0.040522f
C395 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 GNDA 0.082851f
C396 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 GNDA 0.267999f
C397 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 GNDA 0.113211f
C398 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t2 GNDA 0.040522f
C399 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t7 GNDA 0.040522f
C400 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 GNDA 0.082851f
C401 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 GNDA 0.273294f
C402 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 GNDA 0.149186f
C403 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 GNDA 2.38141f
C404 bgr_11_0.V_CMFB_S1 GNDA 2.2214f
C405 two_stage_opamp_dummy_magic_24_0.X.n0 GNDA 0.068212f
C406 two_stage_opamp_dummy_magic_24_0.X.n1 GNDA 0.100044f
C407 two_stage_opamp_dummy_magic_24_0.X.n2 GNDA 0.180382f
C408 two_stage_opamp_dummy_magic_24_0.X.n3 GNDA 0.105665f
C409 two_stage_opamp_dummy_magic_24_0.X.n4 GNDA 0.213297f
C410 two_stage_opamp_dummy_magic_24_0.X.t23 GNDA 0.022737f
C411 two_stage_opamp_dummy_magic_24_0.X.t13 GNDA 0.022737f
C412 two_stage_opamp_dummy_magic_24_0.X.n5 GNDA 0.049474f
C413 two_stage_opamp_dummy_magic_24_0.X.n6 GNDA 0.158096f
C414 two_stage_opamp_dummy_magic_24_0.X.n7 GNDA 0.045474f
C415 two_stage_opamp_dummy_magic_24_0.X.n8 GNDA 0.08695f
C416 two_stage_opamp_dummy_magic_24_0.X.t14 GNDA 0.022737f
C417 two_stage_opamp_dummy_magic_24_0.X.t22 GNDA 0.022737f
C418 two_stage_opamp_dummy_magic_24_0.X.n9 GNDA 0.049474f
C419 two_stage_opamp_dummy_magic_24_0.X.n10 GNDA 0.158096f
C420 two_stage_opamp_dummy_magic_24_0.X.n11 GNDA 0.109539f
C421 two_stage_opamp_dummy_magic_24_0.X.n12 GNDA 0.100044f
C422 two_stage_opamp_dummy_magic_24_0.X.n13 GNDA 0.100044f
C423 two_stage_opamp_dummy_magic_24_0.X.n14 GNDA 0.072759f
C424 two_stage_opamp_dummy_magic_24_0.X.t29 GNDA 0.048885f
C425 two_stage_opamp_dummy_magic_24_0.X.t35 GNDA 0.055574f
C426 two_stage_opamp_dummy_magic_24_0.X.n17 GNDA 0.045322f
C427 two_stage_opamp_dummy_magic_24_0.X.t45 GNDA 0.048885f
C428 two_stage_opamp_dummy_magic_24_0.X.t26 GNDA 0.048885f
C429 two_stage_opamp_dummy_magic_24_0.X.t42 GNDA 0.048885f
C430 two_stage_opamp_dummy_magic_24_0.X.t54 GNDA 0.048885f
C431 two_stage_opamp_dummy_magic_24_0.X.t39 GNDA 0.048885f
C432 two_stage_opamp_dummy_magic_24_0.X.t47 GNDA 0.048885f
C433 two_stage_opamp_dummy_magic_24_0.X.t27 GNDA 0.048885f
C434 two_stage_opamp_dummy_magic_24_0.X.t43 GNDA 0.055574f
C435 two_stage_opamp_dummy_magic_24_0.X.n18 GNDA 0.050154f
C436 two_stage_opamp_dummy_magic_24_0.X.n19 GNDA 0.030695f
C437 two_stage_opamp_dummy_magic_24_0.X.n20 GNDA 0.030695f
C438 two_stage_opamp_dummy_magic_24_0.X.n21 GNDA 0.030695f
C439 two_stage_opamp_dummy_magic_24_0.X.n22 GNDA 0.030695f
C440 two_stage_opamp_dummy_magic_24_0.X.n23 GNDA 0.030695f
C441 two_stage_opamp_dummy_magic_24_0.X.n24 GNDA 0.025864f
C442 two_stage_opamp_dummy_magic_24_0.X.n25 GNDA 0.012559f
C443 two_stage_opamp_dummy_magic_24_0.X.t32 GNDA 0.031832f
C444 two_stage_opamp_dummy_magic_24_0.X.t38 GNDA 0.038653f
C445 two_stage_opamp_dummy_magic_24_0.X.n26 GNDA 0.033822f
C446 two_stage_opamp_dummy_magic_24_0.X.t48 GNDA 0.031832f
C447 two_stage_opamp_dummy_magic_24_0.X.t28 GNDA 0.031832f
C448 two_stage_opamp_dummy_magic_24_0.X.t44 GNDA 0.031832f
C449 two_stage_opamp_dummy_magic_24_0.X.t25 GNDA 0.031832f
C450 two_stage_opamp_dummy_magic_24_0.X.t41 GNDA 0.031832f
C451 two_stage_opamp_dummy_magic_24_0.X.t49 GNDA 0.031832f
C452 two_stage_opamp_dummy_magic_24_0.X.t31 GNDA 0.031832f
C453 two_stage_opamp_dummy_magic_24_0.X.t46 GNDA 0.038653f
C454 two_stage_opamp_dummy_magic_24_0.X.n27 GNDA 0.038653f
C455 two_stage_opamp_dummy_magic_24_0.X.n28 GNDA 0.025011f
C456 two_stage_opamp_dummy_magic_24_0.X.n29 GNDA 0.025011f
C457 two_stage_opamp_dummy_magic_24_0.X.n30 GNDA 0.025011f
C458 two_stage_opamp_dummy_magic_24_0.X.n31 GNDA 0.025011f
C459 two_stage_opamp_dummy_magic_24_0.X.n32 GNDA 0.025011f
C460 two_stage_opamp_dummy_magic_24_0.X.n33 GNDA 0.020179f
C461 two_stage_opamp_dummy_magic_24_0.X.n34 GNDA 0.012559f
C462 two_stage_opamp_dummy_magic_24_0.X.n35 GNDA 0.073548f
C463 two_stage_opamp_dummy_magic_24_0.X.n37 GNDA 0.072759f
C464 two_stage_opamp_dummy_magic_24_0.X.t0 GNDA 0.629399f
C465 two_stage_opamp_dummy_magic_24_0.X.n38 GNDA 0.072759f
C466 two_stage_opamp_dummy_magic_24_0.X.n39 GNDA 0.072759f
C467 two_stage_opamp_dummy_magic_24_0.X.n40 GNDA 0.072076f
C468 two_stage_opamp_dummy_magic_24_0.X.n41 GNDA 0.702092f
C469 two_stage_opamp_dummy_magic_24_0.X.n43 GNDA 0.813992f
C470 two_stage_opamp_dummy_magic_24_0.X.n44 GNDA 0.024092f
C471 two_stage_opamp_dummy_magic_24_0.X.n45 GNDA 0.024253f
C472 two_stage_opamp_dummy_magic_24_0.X.n46 GNDA 0.024253f
C473 two_stage_opamp_dummy_magic_24_0.X.t34 GNDA 0.100044f
C474 two_stage_opamp_dummy_magic_24_0.X.t51 GNDA 0.100044f
C475 two_stage_opamp_dummy_magic_24_0.X.t37 GNDA 0.100044f
C476 two_stage_opamp_dummy_magic_24_0.X.t53 GNDA 0.100044f
C477 two_stage_opamp_dummy_magic_24_0.X.t30 GNDA 0.106553f
C478 two_stage_opamp_dummy_magic_24_0.X.n47 GNDA 0.084439f
C479 two_stage_opamp_dummy_magic_24_0.X.n48 GNDA 0.047748f
C480 two_stage_opamp_dummy_magic_24_0.X.n49 GNDA 0.047748f
C481 two_stage_opamp_dummy_magic_24_0.X.n50 GNDA 0.042916f
C482 two_stage_opamp_dummy_magic_24_0.X.t50 GNDA 0.100044f
C483 two_stage_opamp_dummy_magic_24_0.X.t33 GNDA 0.100044f
C484 two_stage_opamp_dummy_magic_24_0.X.t40 GNDA 0.100044f
C485 two_stage_opamp_dummy_magic_24_0.X.t52 GNDA 0.100044f
C486 two_stage_opamp_dummy_magic_24_0.X.t36 GNDA 0.106553f
C487 two_stage_opamp_dummy_magic_24_0.X.n51 GNDA 0.084439f
C488 two_stage_opamp_dummy_magic_24_0.X.n52 GNDA 0.047748f
C489 two_stage_opamp_dummy_magic_24_0.X.n53 GNDA 0.047748f
C490 two_stage_opamp_dummy_magic_24_0.X.n54 GNDA 0.042916f
C491 two_stage_opamp_dummy_magic_24_0.X.n55 GNDA 0.010305f
C492 two_stage_opamp_dummy_magic_24_0.X.n56 GNDA 0.024414f
C493 two_stage_opamp_dummy_magic_24_0.X.n57 GNDA 0.057469f
C494 two_stage_opamp_dummy_magic_24_0.X.n58 GNDA 0.032778f
C495 two_stage_opamp_dummy_magic_24_0.X.n59 GNDA 0.037198f
C496 two_stage_opamp_dummy_magic_24_0.X.n60 GNDA 1.18688f
C497 two_stage_opamp_dummy_magic_24_0.X.n61 GNDA 0.072759f
C498 two_stage_opamp_dummy_magic_24_0.X.n63 GNDA 0.072759f
C499 two_stage_opamp_dummy_magic_24_0.X.n64 GNDA 0.072759f
C500 two_stage_opamp_dummy_magic_24_0.X.n65 GNDA 0.098208f
C501 two_stage_opamp_dummy_magic_24_0.X.n66 GNDA 0.118233f
C502 two_stage_opamp_dummy_magic_24_0.X.n67 GNDA 0.072759f
C503 two_stage_opamp_dummy_magic_24_0.X.n68 GNDA 0.093771f
C504 two_stage_opamp_dummy_magic_24_0.X.n69 GNDA 0.072759f
C505 two_stage_opamp_dummy_magic_24_0.X.n70 GNDA 0.072759f
C506 two_stage_opamp_dummy_magic_24_0.X.n71 GNDA 0.093771f
C507 two_stage_opamp_dummy_magic_24_0.X.n72 GNDA 0.072759f
C508 two_stage_opamp_dummy_magic_24_0.X.n73 GNDA 0.119891f
C509 two_stage_opamp_dummy_magic_24_0.X.t4 GNDA 0.053054f
C510 two_stage_opamp_dummy_magic_24_0.X.t6 GNDA 0.053054f
C511 two_stage_opamp_dummy_magic_24_0.X.n74 GNDA 0.108526f
C512 two_stage_opamp_dummy_magic_24_0.X.n75 GNDA 0.290397f
C513 two_stage_opamp_dummy_magic_24_0.X.t1 GNDA 0.053054f
C514 two_stage_opamp_dummy_magic_24_0.X.t7 GNDA 0.053054f
C515 two_stage_opamp_dummy_magic_24_0.X.n76 GNDA 0.108526f
C516 two_stage_opamp_dummy_magic_24_0.X.n77 GNDA 0.295195f
C517 two_stage_opamp_dummy_magic_24_0.X.t9 GNDA 0.053054f
C518 two_stage_opamp_dummy_magic_24_0.X.t2 GNDA 0.053054f
C519 two_stage_opamp_dummy_magic_24_0.X.n78 GNDA 0.108526f
C520 two_stage_opamp_dummy_magic_24_0.X.n79 GNDA 0.295195f
C521 two_stage_opamp_dummy_magic_24_0.X.n80 GNDA 0.098167f
C522 two_stage_opamp_dummy_magic_24_0.X.t3 GNDA 0.053054f
C523 two_stage_opamp_dummy_magic_24_0.X.t5 GNDA 0.053054f
C524 two_stage_opamp_dummy_magic_24_0.X.n81 GNDA 0.108526f
C525 two_stage_opamp_dummy_magic_24_0.X.n82 GNDA 0.290397f
C526 two_stage_opamp_dummy_magic_24_0.X.n83 GNDA 0.057546f
C527 two_stage_opamp_dummy_magic_24_0.X.t11 GNDA 0.053054f
C528 two_stage_opamp_dummy_magic_24_0.X.t12 GNDA 0.053054f
C529 two_stage_opamp_dummy_magic_24_0.X.n84 GNDA 0.108526f
C530 two_stage_opamp_dummy_magic_24_0.X.n85 GNDA 0.290397f
C531 two_stage_opamp_dummy_magic_24_0.X.n86 GNDA 0.057546f
C532 two_stage_opamp_dummy_magic_24_0.X.n87 GNDA 0.098167f
C533 two_stage_opamp_dummy_magic_24_0.X.t10 GNDA 0.053054f
C534 two_stage_opamp_dummy_magic_24_0.X.t8 GNDA 0.053054f
C535 two_stage_opamp_dummy_magic_24_0.X.n88 GNDA 0.108526f
C536 two_stage_opamp_dummy_magic_24_0.X.n89 GNDA 0.290397f
C537 two_stage_opamp_dummy_magic_24_0.X.n90 GNDA 0.093771f
C538 two_stage_opamp_dummy_magic_24_0.X.n91 GNDA 0.080449f
C539 two_stage_opamp_dummy_magic_24_0.X.n92 GNDA 0.048506f
C540 two_stage_opamp_dummy_magic_24_0.X.n93 GNDA 0.048506f
C541 two_stage_opamp_dummy_magic_24_0.X.n94 GNDA 0.080449f
C542 two_stage_opamp_dummy_magic_24_0.X.n95 GNDA 0.093771f
C543 two_stage_opamp_dummy_magic_24_0.X.n96 GNDA 0.165892f
C544 two_stage_opamp_dummy_magic_24_0.X.n97 GNDA 0.245724f
C545 two_stage_opamp_dummy_magic_24_0.X.n98 GNDA 0.312481f
C546 two_stage_opamp_dummy_magic_24_0.X.n99 GNDA 0.072759f
C547 two_stage_opamp_dummy_magic_24_0.X.n100 GNDA 0.072759f
C548 two_stage_opamp_dummy_magic_24_0.X.n101 GNDA 0.118233f
C549 two_stage_opamp_dummy_magic_24_0.X.n102 GNDA 0.072759f
C550 two_stage_opamp_dummy_magic_24_0.X.n103 GNDA 0.072759f
C551 two_stage_opamp_dummy_magic_24_0.X.n104 GNDA 0.072759f
C552 two_stage_opamp_dummy_magic_24_0.X.n105 GNDA 0.072759f
C553 two_stage_opamp_dummy_magic_24_0.X.n106 GNDA 0.118233f
C554 two_stage_opamp_dummy_magic_24_0.X.n107 GNDA 0.072759f
C555 two_stage_opamp_dummy_magic_24_0.X.n108 GNDA 0.072759f
C556 two_stage_opamp_dummy_magic_24_0.X.n109 GNDA 0.072759f
C557 two_stage_opamp_dummy_magic_24_0.X.n110 GNDA 0.072759f
C558 two_stage_opamp_dummy_magic_24_0.X.n111 GNDA 0.072759f
C559 two_stage_opamp_dummy_magic_24_0.X.n112 GNDA 0.072759f
C560 two_stage_opamp_dummy_magic_24_0.X.n113 GNDA 0.072759f
C561 two_stage_opamp_dummy_magic_24_0.X.n114 GNDA 0.118233f
C562 two_stage_opamp_dummy_magic_24_0.X.n115 GNDA 0.386532f
C563 two_stage_opamp_dummy_magic_24_0.X.n116 GNDA 0.386532f
C564 two_stage_opamp_dummy_magic_24_0.X.n117 GNDA 0.072076f
C565 two_stage_opamp_dummy_magic_24_0.X.n118 GNDA 0.072759f
C566 two_stage_opamp_dummy_magic_24_0.X.n119 GNDA 0.072759f
C567 two_stage_opamp_dummy_magic_24_0.X.n121 GNDA 0.813992f
C568 two_stage_opamp_dummy_magic_24_0.X.n122 GNDA 0.813992f
C569 two_stage_opamp_dummy_magic_24_0.X.n124 GNDA 0.445649f
C570 two_stage_opamp_dummy_magic_24_0.X.n125 GNDA 1.83665f
C571 two_stage_opamp_dummy_magic_24_0.X.n126 GNDA 0.404722f
C572 two_stage_opamp_dummy_magic_24_0.X.n127 GNDA 0.16674f
C573 two_stage_opamp_dummy_magic_24_0.X.n128 GNDA 0.418365f
C574 two_stage_opamp_dummy_magic_24_0.X.n129 GNDA 0.100044f
C575 two_stage_opamp_dummy_magic_24_0.X.n130 GNDA 0.100044f
C576 two_stage_opamp_dummy_magic_24_0.X.n131 GNDA 0.100044f
C577 two_stage_opamp_dummy_magic_24_0.X.n132 GNDA 0.180382f
C578 two_stage_opamp_dummy_magic_24_0.X.t16 GNDA 0.022737f
C579 two_stage_opamp_dummy_magic_24_0.X.t24 GNDA 0.022737f
C580 two_stage_opamp_dummy_magic_24_0.X.n133 GNDA 0.049474f
C581 two_stage_opamp_dummy_magic_24_0.X.n134 GNDA 0.154078f
C582 two_stage_opamp_dummy_magic_24_0.X.n135 GNDA 0.105665f
C583 two_stage_opamp_dummy_magic_24_0.X.n136 GNDA 0.076464f
C584 two_stage_opamp_dummy_magic_24_0.X.n137 GNDA 0.045474f
C585 two_stage_opamp_dummy_magic_24_0.X.n138 GNDA 0.105665f
C586 two_stage_opamp_dummy_magic_24_0.X.t18 GNDA 0.022737f
C587 two_stage_opamp_dummy_magic_24_0.X.t21 GNDA 0.022737f
C588 two_stage_opamp_dummy_magic_24_0.X.n139 GNDA 0.049474f
C589 two_stage_opamp_dummy_magic_24_0.X.n140 GNDA 0.154078f
C590 two_stage_opamp_dummy_magic_24_0.X.n141 GNDA 0.050789f
C591 two_stage_opamp_dummy_magic_24_0.X.t15 GNDA 0.022737f
C592 two_stage_opamp_dummy_magic_24_0.X.t19 GNDA 0.022737f
C593 two_stage_opamp_dummy_magic_24_0.X.n142 GNDA 0.049474f
C594 two_stage_opamp_dummy_magic_24_0.X.n143 GNDA 0.154078f
C595 two_stage_opamp_dummy_magic_24_0.X.n144 GNDA 0.050789f
C596 two_stage_opamp_dummy_magic_24_0.X.n145 GNDA 0.08695f
C597 two_stage_opamp_dummy_magic_24_0.X.t17 GNDA 0.022737f
C598 two_stage_opamp_dummy_magic_24_0.X.t20 GNDA 0.022737f
C599 two_stage_opamp_dummy_magic_24_0.X.n146 GNDA 0.049474f
C600 two_stage_opamp_dummy_magic_24_0.X.n147 GNDA 0.154078f
C601 two_stage_opamp_dummy_magic_24_0.X.n148 GNDA 0.105665f
C602 two_stage_opamp_dummy_magic_24_0.X.n149 GNDA 0.076464f
C603 two_stage_opamp_dummy_magic_24_0.X.n150 GNDA 0.123394f
C604 two_stage_opamp_dummy_magic_24_0.X.n151 GNDA 0.263643f
C605 two_stage_opamp_dummy_magic_24_0.X.n152 GNDA 0.342902f
C606 two_stage_opamp_dummy_magic_24_0.X.n153 GNDA 0.100044f
C607 two_stage_opamp_dummy_magic_24_0.X.n154 GNDA 0.180382f
C608 two_stage_opamp_dummy_magic_24_0.X.n155 GNDA 0.100044f
C609 two_stage_opamp_dummy_magic_24_0.X.n156 GNDA 0.081854f
C610 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t8 GNDA 0.070681f
C611 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t9 GNDA 0.069492f
C612 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 GNDA 0.503602f
C613 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t6 GNDA 0.318882f
C614 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t7 GNDA 0.100545f
C615 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 GNDA 1.73362f
C616 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t4 GNDA 0.061551f
C617 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t2 GNDA 0.061551f
C618 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 GNDA 0.216779f
C619 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t0 GNDA 0.061551f
C620 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t1 GNDA 0.061551f
C621 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 GNDA 0.206258f
C622 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 GNDA 0.963909f
C623 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t3 GNDA 0.061551f
C624 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t5 GNDA 0.061551f
C625 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 GNDA 0.206258f
C626 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 GNDA 0.689269f
C627 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 GNDA 2.33472f
C628 two_stage_opamp_dummy_magic_24_0.V_source.n0 GNDA 0.406711f
C629 two_stage_opamp_dummy_magic_24_0.V_source.n1 GNDA 0.659723f
C630 two_stage_opamp_dummy_magic_24_0.V_source.n2 GNDA 0.878055f
C631 two_stage_opamp_dummy_magic_24_0.V_source.n3 GNDA 0.962374f
C632 two_stage_opamp_dummy_magic_24_0.V_source.n4 GNDA 0.121245f
C633 two_stage_opamp_dummy_magic_24_0.V_source.n5 GNDA 0.057482f
C634 two_stage_opamp_dummy_magic_24_0.V_source.n6 GNDA 0.270618f
C635 two_stage_opamp_dummy_magic_24_0.V_source.n7 GNDA 0.12763f
C636 two_stage_opamp_dummy_magic_24_0.V_source.n8 GNDA 0.085972f
C637 two_stage_opamp_dummy_magic_24_0.V_source.t29 GNDA 0.023646f
C638 two_stage_opamp_dummy_magic_24_0.V_source.t27 GNDA 0.023646f
C639 two_stage_opamp_dummy_magic_24_0.V_source.n9 GNDA 0.051451f
C640 two_stage_opamp_dummy_magic_24_0.V_source.n10 GNDA 0.215937f
C641 two_stage_opamp_dummy_magic_24_0.V_source.t5 GNDA 0.023646f
C642 two_stage_opamp_dummy_magic_24_0.V_source.t30 GNDA 0.023646f
C643 two_stage_opamp_dummy_magic_24_0.V_source.n11 GNDA 0.051451f
C644 two_stage_opamp_dummy_magic_24_0.V_source.n12 GNDA 0.208467f
C645 two_stage_opamp_dummy_magic_24_0.V_source.n13 GNDA 0.12763f
C646 two_stage_opamp_dummy_magic_24_0.V_source.n14 GNDA 0.099142f
C647 two_stage_opamp_dummy_magic_24_0.V_source.t2 GNDA 0.023646f
C648 two_stage_opamp_dummy_magic_24_0.V_source.t34 GNDA 0.023646f
C649 two_stage_opamp_dummy_magic_24_0.V_source.n15 GNDA 0.051451f
C650 two_stage_opamp_dummy_magic_24_0.V_source.n16 GNDA 0.208467f
C651 two_stage_opamp_dummy_magic_24_0.V_source.n17 GNDA 0.050539f
C652 two_stage_opamp_dummy_magic_24_0.V_source.n18 GNDA 0.050539f
C653 two_stage_opamp_dummy_magic_24_0.V_source.t26 GNDA 0.023646f
C654 two_stage_opamp_dummy_magic_24_0.V_source.t40 GNDA 0.023646f
C655 two_stage_opamp_dummy_magic_24_0.V_source.n19 GNDA 0.051451f
C656 two_stage_opamp_dummy_magic_24_0.V_source.n20 GNDA 0.156146f
C657 two_stage_opamp_dummy_magic_24_0.V_source.t31 GNDA 0.023646f
C658 two_stage_opamp_dummy_magic_24_0.V_source.t0 GNDA 0.023646f
C659 two_stage_opamp_dummy_magic_24_0.V_source.n21 GNDA 0.051451f
C660 two_stage_opamp_dummy_magic_24_0.V_source.n22 GNDA 0.156146f
C661 two_stage_opamp_dummy_magic_24_0.V_source.n23 GNDA 0.127782f
C662 two_stage_opamp_dummy_magic_24_0.V_source.t7 GNDA 0.023646f
C663 two_stage_opamp_dummy_magic_24_0.V_source.t1 GNDA 0.023646f
C664 two_stage_opamp_dummy_magic_24_0.V_source.n24 GNDA 0.051451f
C665 two_stage_opamp_dummy_magic_24_0.V_source.n25 GNDA 0.156146f
C666 two_stage_opamp_dummy_magic_24_0.V_source.n26 GNDA 0.127782f
C667 two_stage_opamp_dummy_magic_24_0.V_source.t36 GNDA 0.023646f
C668 two_stage_opamp_dummy_magic_24_0.V_source.t6 GNDA 0.023646f
C669 two_stage_opamp_dummy_magic_24_0.V_source.n27 GNDA 0.051451f
C670 two_stage_opamp_dummy_magic_24_0.V_source.n28 GNDA 0.156146f
C671 two_stage_opamp_dummy_magic_24_0.V_source.n29 GNDA 0.050539f
C672 two_stage_opamp_dummy_magic_24_0.V_source.t32 GNDA 0.023646f
C673 two_stage_opamp_dummy_magic_24_0.V_source.t3 GNDA 0.023646f
C674 two_stage_opamp_dummy_magic_24_0.V_source.n30 GNDA 0.051451f
C675 two_stage_opamp_dummy_magic_24_0.V_source.n31 GNDA 0.215937f
C676 two_stage_opamp_dummy_magic_24_0.V_source.t35 GNDA 0.023646f
C677 two_stage_opamp_dummy_magic_24_0.V_source.t39 GNDA 0.023646f
C678 two_stage_opamp_dummy_magic_24_0.V_source.n32 GNDA 0.051451f
C679 two_stage_opamp_dummy_magic_24_0.V_source.n33 GNDA 0.208467f
C680 two_stage_opamp_dummy_magic_24_0.V_source.n34 GNDA 0.085972f
C681 two_stage_opamp_dummy_magic_24_0.V_source.n35 GNDA 0.050539f
C682 two_stage_opamp_dummy_magic_24_0.V_source.t28 GNDA 0.023646f
C683 two_stage_opamp_dummy_magic_24_0.V_source.t4 GNDA 0.023646f
C684 two_stage_opamp_dummy_magic_24_0.V_source.n36 GNDA 0.051451f
C685 two_stage_opamp_dummy_magic_24_0.V_source.n37 GNDA 0.208467f
C686 two_stage_opamp_dummy_magic_24_0.V_source.n38 GNDA 0.099142f
C687 two_stage_opamp_dummy_magic_24_0.V_source.n39 GNDA 0.270618f
C688 two_stage_opamp_dummy_magic_24_0.V_source.t13 GNDA 0.03941f
C689 two_stage_opamp_dummy_magic_24_0.V_source.t21 GNDA 0.03941f
C690 two_stage_opamp_dummy_magic_24_0.V_source.n40 GNDA 0.084253f
C691 two_stage_opamp_dummy_magic_24_0.V_source.n41 GNDA 0.24606f
C692 two_stage_opamp_dummy_magic_24_0.V_source.t12 GNDA 0.03941f
C693 two_stage_opamp_dummy_magic_24_0.V_source.t20 GNDA 0.03941f
C694 two_stage_opamp_dummy_magic_24_0.V_source.n42 GNDA 0.084253f
C695 two_stage_opamp_dummy_magic_24_0.V_source.n43 GNDA 0.24606f
C696 two_stage_opamp_dummy_magic_24_0.V_source.n44 GNDA 0.057482f
C697 two_stage_opamp_dummy_magic_24_0.V_source.n45 GNDA 0.099497f
C698 two_stage_opamp_dummy_magic_24_0.V_source.t9 GNDA 0.03941f
C699 two_stage_opamp_dummy_magic_24_0.V_source.t17 GNDA 0.03941f
C700 two_stage_opamp_dummy_magic_24_0.V_source.n46 GNDA 0.084253f
C701 two_stage_opamp_dummy_magic_24_0.V_source.n47 GNDA 0.250491f
C702 two_stage_opamp_dummy_magic_24_0.V_source.t19 GNDA 0.03941f
C703 two_stage_opamp_dummy_magic_24_0.V_source.t22 GNDA 0.03941f
C704 two_stage_opamp_dummy_magic_24_0.V_source.n48 GNDA 0.084253f
C705 two_stage_opamp_dummy_magic_24_0.V_source.n49 GNDA 0.299211f
C706 two_stage_opamp_dummy_magic_24_0.V_source.n50 GNDA 0.216431f
C707 two_stage_opamp_dummy_magic_24_0.V_source.n51 GNDA 0.076902f
C708 two_stage_opamp_dummy_magic_24_0.V_source.t14 GNDA 0.03941f
C709 two_stage_opamp_dummy_magic_24_0.V_source.t11 GNDA 0.03941f
C710 two_stage_opamp_dummy_magic_24_0.V_source.n52 GNDA 0.084253f
C711 two_stage_opamp_dummy_magic_24_0.V_source.n53 GNDA 0.299211f
C712 two_stage_opamp_dummy_magic_24_0.V_source.n54 GNDA 0.057482f
C713 two_stage_opamp_dummy_magic_24_0.V_source.t15 GNDA 0.03941f
C714 two_stage_opamp_dummy_magic_24_0.V_source.t23 GNDA 0.03941f
C715 two_stage_opamp_dummy_magic_24_0.V_source.n55 GNDA 0.084253f
C716 two_stage_opamp_dummy_magic_24_0.V_source.n56 GNDA 0.299211f
C717 two_stage_opamp_dummy_magic_24_0.V_source.n57 GNDA 0.057482f
C718 two_stage_opamp_dummy_magic_24_0.V_source.t16 GNDA 0.03941f
C719 two_stage_opamp_dummy_magic_24_0.V_source.t25 GNDA 0.03941f
C720 two_stage_opamp_dummy_magic_24_0.V_source.n58 GNDA 0.084253f
C721 two_stage_opamp_dummy_magic_24_0.V_source.n59 GNDA 0.24606f
C722 two_stage_opamp_dummy_magic_24_0.V_source.n60 GNDA 0.057482f
C723 two_stage_opamp_dummy_magic_24_0.V_source.t18 GNDA 0.03941f
C724 two_stage_opamp_dummy_magic_24_0.V_source.t8 GNDA 0.03941f
C725 two_stage_opamp_dummy_magic_24_0.V_source.n61 GNDA 0.084253f
C726 two_stage_opamp_dummy_magic_24_0.V_source.n62 GNDA 0.191036f
C727 two_stage_opamp_dummy_magic_24_0.V_source.t38 GNDA 0.085443f
C728 two_stage_opamp_dummy_magic_24_0.V_source.n63 GNDA 0.353377f
C729 two_stage_opamp_dummy_magic_24_0.V_source.n64 GNDA 0.047292f
C730 two_stage_opamp_dummy_magic_24_0.V_source.t24 GNDA 0.03941f
C731 two_stage_opamp_dummy_magic_24_0.V_source.t10 GNDA 0.03941f
C732 two_stage_opamp_dummy_magic_24_0.V_source.n65 GNDA 0.084253f
C733 two_stage_opamp_dummy_magic_24_0.V_source.n66 GNDA 0.24606f
C734 two_stage_opamp_dummy_magic_24_0.V_source.n67 GNDA 0.099497f
C735 two_stage_opamp_dummy_magic_24_0.V_source.t37 GNDA 0.03941f
C736 two_stage_opamp_dummy_magic_24_0.V_source.t33 GNDA 0.03941f
C737 two_stage_opamp_dummy_magic_24_0.V_source.n68 GNDA 0.084253f
C738 two_stage_opamp_dummy_magic_24_0.V_source.n69 GNDA 0.314894f
C739 two_stage_opamp_dummy_magic_24_0.V_source.n70 GNDA 0.207322f
C740 two_stage_opamp_dummy_magic_24_0.V_err_gate.t4 GNDA 0.020119f
C741 two_stage_opamp_dummy_magic_24_0.V_err_gate.t5 GNDA 0.020119f
C742 two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 GNDA 0.248145f
C743 two_stage_opamp_dummy_magic_24_0.V_err_gate.t0 GNDA 0.050298f
C744 two_stage_opamp_dummy_magic_24_0.V_err_gate.t3 GNDA 0.050298f
C745 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 GNDA 0.154097f
C746 two_stage_opamp_dummy_magic_24_0.V_err_gate.t8 GNDA 0.056165f
C747 two_stage_opamp_dummy_magic_24_0.V_err_gate.t6 GNDA 0.056165f
C748 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 GNDA 0.084365f
C749 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 GNDA 0.311368f
C750 two_stage_opamp_dummy_magic_24_0.V_err_gate.t2 GNDA 0.050298f
C751 two_stage_opamp_dummy_magic_24_0.V_err_gate.t1 GNDA 0.050298f
C752 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 GNDA 0.153429f
C753 two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 GNDA 0.23824f
C754 two_stage_opamp_dummy_magic_24_0.V_err_gate.t7 GNDA 0.056165f
C755 two_stage_opamp_dummy_magic_24_0.V_err_gate.t9 GNDA 0.056165f
C756 two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 GNDA 0.084365f
C757 bgr_11_0.cap_res1.t5 GNDA 0.331712f
C758 bgr_11_0.cap_res1.t17 GNDA 0.349187f
C759 bgr_11_0.cap_res1.t9 GNDA 0.350452f
C760 bgr_11_0.cap_res1.t12 GNDA 0.331712f
C761 bgr_11_0.cap_res1.t19 GNDA 0.349187f
C762 bgr_11_0.cap_res1.t16 GNDA 0.350452f
C763 bgr_11_0.cap_res1.t4 GNDA 0.331712f
C764 bgr_11_0.cap_res1.t15 GNDA 0.349187f
C765 bgr_11_0.cap_res1.t8 GNDA 0.350452f
C766 bgr_11_0.cap_res1.t0 GNDA 0.331712f
C767 bgr_11_0.cap_res1.t7 GNDA 0.349187f
C768 bgr_11_0.cap_res1.t1 GNDA 0.350452f
C769 bgr_11_0.cap_res1.t2 GNDA 0.331712f
C770 bgr_11_0.cap_res1.t14 GNDA 0.349187f
C771 bgr_11_0.cap_res1.t6 GNDA 0.350452f
C772 bgr_11_0.cap_res1.n0 GNDA 0.23406f
C773 bgr_11_0.cap_res1.t10 GNDA 0.186395f
C774 bgr_11_0.cap_res1.n1 GNDA 0.253961f
C775 bgr_11_0.cap_res1.t3 GNDA 0.186395f
C776 bgr_11_0.cap_res1.n2 GNDA 0.253961f
C777 bgr_11_0.cap_res1.t11 GNDA 0.186395f
C778 bgr_11_0.cap_res1.n3 GNDA 0.253961f
C779 bgr_11_0.cap_res1.t18 GNDA 0.186395f
C780 bgr_11_0.cap_res1.n4 GNDA 0.253961f
C781 bgr_11_0.cap_res1.t13 GNDA 0.363549f
C782 bgr_11_0.cap_res1.t20 GNDA 0.08421f
C783 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t1 GNDA 0.023655f
C784 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t13 GNDA 0.023655f
C785 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 GNDA 0.074393f
C786 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t12 GNDA 0.023655f
C787 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t14 GNDA 0.023655f
C788 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 GNDA 0.050743f
C789 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 GNDA 3.78749f
C790 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t0 GNDA 0.289539f
C791 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 GNDA 0.082281f
C792 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 GNDA 0.141574f
C793 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t10 GNDA 0.070966f
C794 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t6 GNDA 0.070966f
C795 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 GNDA 0.151783f
C796 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 GNDA 0.474777f
C797 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t11 GNDA 0.070966f
C798 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t5 GNDA 0.070966f
C799 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 GNDA 0.151783f
C800 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 GNDA 0.461918f
C801 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 GNDA 0.141574f
C802 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 GNDA 0.082281f
C803 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t9 GNDA 0.070966f
C804 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t4 GNDA 0.070966f
C805 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 GNDA 0.151783f
C806 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 GNDA 0.461918f
C807 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 GNDA 0.082281f
C808 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t8 GNDA 0.070966f
C809 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t3 GNDA 0.070966f
C810 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 GNDA 0.151783f
C811 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 GNDA 0.461918f
C812 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 GNDA 0.141574f
C813 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t7 GNDA 0.070966f
C814 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t2 GNDA 0.070966f
C815 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 GNDA 0.151783f
C816 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 GNDA 0.468348f
C817 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 GNDA 0.165918f
C818 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 GNDA 2.34089f
C819 bgr_11_0.V_CMFB_S4 GNDA 6.72738f
C820 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t14 GNDA 0.022867f
C821 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t7 GNDA 0.022867f
C822 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 GNDA 0.071913f
C823 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t12 GNDA 0.022867f
C824 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t13 GNDA 0.022867f
C825 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 GNDA 0.049052f
C826 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 GNDA 3.66124f
C827 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t11 GNDA 0.279888f
C828 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 GNDA 0.079538f
C829 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 GNDA 0.136855f
C830 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t8 GNDA 0.068601f
C831 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t5 GNDA 0.068601f
C832 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 GNDA 0.146724f
C833 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 GNDA 0.458951f
C834 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t1 GNDA 0.068601f
C835 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t4 GNDA 0.068601f
C836 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 GNDA 0.146724f
C837 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 GNDA 0.446521f
C838 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 GNDA 0.136855f
C839 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 GNDA 0.079538f
C840 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t9 GNDA 0.068601f
C841 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t3 GNDA 0.068601f
C842 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 GNDA 0.146724f
C843 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 GNDA 0.446521f
C844 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 GNDA 0.079538f
C845 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t0 GNDA 0.068601f
C846 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t2 GNDA 0.068601f
C847 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 GNDA 0.146724f
C848 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 GNDA 0.446521f
C849 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 GNDA 0.136855f
C850 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t10 GNDA 0.068601f
C851 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t6 GNDA 0.068601f
C852 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 GNDA 0.146724f
C853 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 GNDA 0.452736f
C854 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 GNDA 0.160387f
C855 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 GNDA 2.26286f
C856 bgr_11_0.V_CMFB_S2 GNDA 6.50314f
C857 two_stage_opamp_dummy_magic_24_0.VD3.n0 GNDA 0.141913f
C858 two_stage_opamp_dummy_magic_24_0.VD3.n1 GNDA 0.141913f
C859 two_stage_opamp_dummy_magic_24_0.VD3.n2 GNDA 0.09179f
C860 two_stage_opamp_dummy_magic_24_0.VD3.n3 GNDA 0.158068f
C861 two_stage_opamp_dummy_magic_24_0.VD3.n4 GNDA 0.138157f
C862 two_stage_opamp_dummy_magic_24_0.VD3.n5 GNDA 0.291251f
C863 two_stage_opamp_dummy_magic_24_0.VD3.n6 GNDA 0.470599f
C864 two_stage_opamp_dummy_magic_24_0.VD3.n7 GNDA 0.185256f
C865 two_stage_opamp_dummy_magic_24_0.VD3.n8 GNDA 0.069079f
C866 two_stage_opamp_dummy_magic_24_0.VD3.n9 GNDA 0.138157f
C867 two_stage_opamp_dummy_magic_24_0.VD3.n10 GNDA 0.138157f
C868 two_stage_opamp_dummy_magic_24_0.VD3.n11 GNDA 0.138157f
C869 two_stage_opamp_dummy_magic_24_0.VD3.n12 GNDA 0.09179f
C870 two_stage_opamp_dummy_magic_24_0.VD3.n13 GNDA 0.138157f
C871 two_stage_opamp_dummy_magic_24_0.VD3.n14 GNDA 0.069079f
C872 two_stage_opamp_dummy_magic_24_0.VD3.n15 GNDA 0.138157f
C873 two_stage_opamp_dummy_magic_24_0.VD3.n16 GNDA 0.069079f
C874 two_stage_opamp_dummy_magic_24_0.VD3.n17 GNDA 0.138157f
C875 two_stage_opamp_dummy_magic_24_0.VD3.n18 GNDA 0.09179f
C876 two_stage_opamp_dummy_magic_24_0.VD3.n19 GNDA 0.138157f
C877 two_stage_opamp_dummy_magic_24_0.VD3.n20 GNDA 0.069079f
C878 two_stage_opamp_dummy_magic_24_0.VD3.n21 GNDA 0.365754f
C879 two_stage_opamp_dummy_magic_24_0.VD3.n22 GNDA 0.069079f
C880 two_stage_opamp_dummy_magic_24_0.VD3.n23 GNDA 0.09179f
C881 two_stage_opamp_dummy_magic_24_0.VD3.n24 GNDA 0.233055f
C882 two_stage_opamp_dummy_magic_24_0.VD3.n25 GNDA 0.296931f
C883 two_stage_opamp_dummy_magic_24_0.VD3.n26 GNDA 0.187808f
C884 two_stage_opamp_dummy_magic_24_0.VD3.n27 GNDA 0.43114f
C885 two_stage_opamp_dummy_magic_24_0.VD3.t36 GNDA 0.05037f
C886 two_stage_opamp_dummy_magic_24_0.VD3.n28 GNDA 0.054635f
C887 two_stage_opamp_dummy_magic_24_0.VD3.t34 GNDA 0.05037f
C888 two_stage_opamp_dummy_magic_24_0.VD3.t26 GNDA 0.05037f
C889 two_stage_opamp_dummy_magic_24_0.VD3.n29 GNDA 0.103037f
C890 two_stage_opamp_dummy_magic_24_0.VD3.t33 GNDA 0.05037f
C891 two_stage_opamp_dummy_magic_24_0.VD3.t35 GNDA 0.05037f
C892 two_stage_opamp_dummy_magic_24_0.VD3.n30 GNDA 0.103037f
C893 two_stage_opamp_dummy_magic_24_0.VD3.n31 GNDA 0.284144f
C894 two_stage_opamp_dummy_magic_24_0.VD3.t28 GNDA 0.05037f
C895 two_stage_opamp_dummy_magic_24_0.VD3.t31 GNDA 0.05037f
C896 two_stage_opamp_dummy_magic_24_0.VD3.n32 GNDA 0.103037f
C897 two_stage_opamp_dummy_magic_24_0.VD3.n33 GNDA 0.284144f
C898 two_stage_opamp_dummy_magic_24_0.VD3.n34 GNDA 0.093202f
C899 two_stage_opamp_dummy_magic_24_0.VD3.t27 GNDA 0.05037f
C900 two_stage_opamp_dummy_magic_24_0.VD3.t30 GNDA 0.05037f
C901 two_stage_opamp_dummy_magic_24_0.VD3.n35 GNDA 0.103037f
C902 two_stage_opamp_dummy_magic_24_0.VD3.n36 GNDA 0.304985f
C903 two_stage_opamp_dummy_magic_24_0.VD3.t0 GNDA 0.088322f
C904 two_stage_opamp_dummy_magic_24_0.VD3.n37 GNDA 0.201305f
C905 two_stage_opamp_dummy_magic_24_0.VD3.t15 GNDA 0.05037f
C906 two_stage_opamp_dummy_magic_24_0.VD3.t21 GNDA 0.05037f
C907 two_stage_opamp_dummy_magic_24_0.VD3.n38 GNDA 0.106864f
C908 two_stage_opamp_dummy_magic_24_0.VD3.n39 GNDA 0.405627f
C909 two_stage_opamp_dummy_magic_24_0.VD3.t17 GNDA 0.05037f
C910 two_stage_opamp_dummy_magic_24_0.VD3.t23 GNDA 0.05037f
C911 two_stage_opamp_dummy_magic_24_0.VD3.n40 GNDA 0.106864f
C912 two_stage_opamp_dummy_magic_24_0.VD3.t25 GNDA 0.05037f
C913 two_stage_opamp_dummy_magic_24_0.VD3.t7 GNDA 0.05037f
C914 two_stage_opamp_dummy_magic_24_0.VD3.n41 GNDA 0.106864f
C915 two_stage_opamp_dummy_magic_24_0.VD3.t11 GNDA 0.05037f
C916 two_stage_opamp_dummy_magic_24_0.VD3.t9 GNDA 0.05037f
C917 two_stage_opamp_dummy_magic_24_0.VD3.n42 GNDA 0.106864f
C918 two_stage_opamp_dummy_magic_24_0.VD3.t13 GNDA 0.05037f
C919 two_stage_opamp_dummy_magic_24_0.VD3.t19 GNDA 0.05037f
C920 two_stage_opamp_dummy_magic_24_0.VD3.n43 GNDA 0.106864f
C921 two_stage_opamp_dummy_magic_24_0.VD3.n44 GNDA 0.450875f
C922 two_stage_opamp_dummy_magic_24_0.VD3.t3 GNDA 0.088322f
C923 two_stage_opamp_dummy_magic_24_0.VD3.t5 GNDA 0.179173f
C924 two_stage_opamp_dummy_magic_24_0.VD3.t2 GNDA 0.179173f
C925 two_stage_opamp_dummy_magic_24_0.VD3.n45 GNDA 0.519765f
C926 two_stage_opamp_dummy_magic_24_0.VD3.t1 GNDA 0.429348f
C927 two_stage_opamp_dummy_magic_24_0.VD3.t14 GNDA 0.336759f
C928 two_stage_opamp_dummy_magic_24_0.VD3.t20 GNDA 0.336759f
C929 two_stage_opamp_dummy_magic_24_0.VD3.t16 GNDA 0.336759f
C930 two_stage_opamp_dummy_magic_24_0.VD3.t22 GNDA 0.336759f
C931 two_stage_opamp_dummy_magic_24_0.VD3.t24 GNDA 0.336759f
C932 two_stage_opamp_dummy_magic_24_0.VD3.t6 GNDA 0.336759f
C933 two_stage_opamp_dummy_magic_24_0.VD3.t10 GNDA 0.336759f
C934 two_stage_opamp_dummy_magic_24_0.VD3.t8 GNDA 0.336759f
C935 two_stage_opamp_dummy_magic_24_0.VD3.t12 GNDA 0.336759f
C936 two_stage_opamp_dummy_magic_24_0.VD3.t18 GNDA 0.336759f
C937 two_stage_opamp_dummy_magic_24_0.VD3.t4 GNDA 0.429348f
C938 two_stage_opamp_dummy_magic_24_0.VD3.n46 GNDA 0.519765f
C939 two_stage_opamp_dummy_magic_24_0.VD3.n47 GNDA 0.212445f
C940 two_stage_opamp_dummy_magic_24_0.VD3.n48 GNDA 0.249218f
C941 two_stage_opamp_dummy_magic_24_0.VD3.n49 GNDA 0.405627f
C942 two_stage_opamp_dummy_magic_24_0.VD3.n50 GNDA 0.405627f
C943 two_stage_opamp_dummy_magic_24_0.VD3.n51 GNDA 0.405627f
C944 two_stage_opamp_dummy_magic_24_0.VD3.n52 GNDA 0.141913f
C945 two_stage_opamp_dummy_magic_24_0.VD3.n53 GNDA 0.40152f
C946 two_stage_opamp_dummy_magic_24_0.VD3.t29 GNDA 0.05037f
C947 two_stage_opamp_dummy_magic_24_0.VD3.t32 GNDA 0.05037f
C948 two_stage_opamp_dummy_magic_24_0.VD3.n54 GNDA 0.103037f
C949 two_stage_opamp_dummy_magic_24_0.VD3.n55 GNDA 0.284144f
C950 two_stage_opamp_dummy_magic_24_0.VD3.n56 GNDA 0.093202f
C951 two_stage_opamp_dummy_magic_24_0.VD3.n57 GNDA 0.054635f
C952 two_stage_opamp_dummy_magic_24_0.VD3.n58 GNDA 0.284144f
C953 two_stage_opamp_dummy_magic_24_0.VD3.n59 GNDA 0.103037f
C954 two_stage_opamp_dummy_magic_24_0.VD3.t37 GNDA 0.05037f
C955 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 GNDA 8.08f
C956 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 GNDA 0.995855f
C957 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 GNDA 0.21811f
C958 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 GNDA 8.5645f
C959 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 GNDA 12.484099f
C960 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 GNDA 0.018875f
C961 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 GNDA 0.018875f
C962 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 GNDA 0.217564f
C963 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 GNDA 0.108068f
C964 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 GNDA 0.018875f
C965 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 GNDA 0.034273f
C966 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 GNDA 0.108068f
C967 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 GNDA 0.018875f
C968 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 GNDA 0.218122f
C969 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t0 GNDA 0.014156f
C970 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t10 GNDA 0.014156f
C971 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 GNDA 0.033385f
C972 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t11 GNDA 0.014156f
C973 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t9 GNDA 0.014156f
C974 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 GNDA 0.033385f
C975 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t14 GNDA 0.025127f
C976 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t23 GNDA 0.025127f
C977 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t12 GNDA 0.025127f
C978 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t22 GNDA 0.025127f
C979 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t31 GNDA 0.025127f
C980 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t20 GNDA 0.025127f
C981 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t29 GNDA 0.025127f
C982 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t13 GNDA 0.029328f
C983 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 GNDA 0.027651f
C984 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 GNDA 0.017341f
C985 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 GNDA 0.017341f
C986 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 GNDA 0.017341f
C987 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 GNDA 0.017341f
C988 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 GNDA 0.017341f
C989 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 GNDA 0.016228f
C990 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t25 GNDA 0.025127f
C991 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t28 GNDA 0.025127f
C992 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t19 GNDA 0.025127f
C993 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t16 GNDA 0.025127f
C994 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t26 GNDA 0.025127f
C995 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t17 GNDA 0.025127f
C996 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t27 GNDA 0.025127f
C997 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t18 GNDA 0.025127f
C998 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t30 GNDA 0.025127f
C999 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t21 GNDA 0.025127f
C1000 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t24 GNDA 0.025127f
C1001 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t15 GNDA 0.029328f
C1002 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 GNDA 0.027651f
C1003 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 GNDA 0.017341f
C1004 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 GNDA 0.017341f
C1005 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 GNDA 0.017341f
C1006 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 GNDA 0.017341f
C1007 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 GNDA 0.017341f
C1008 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 GNDA 0.017341f
C1009 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 GNDA 0.017341f
C1010 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 GNDA 0.016228f
C1011 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 GNDA 0.014466f
C1012 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 GNDA 0.016228f
C1013 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n34 GNDA 0.016228f
C1014 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n35 GNDA 0.014446f
C1015 bgr_11_0.PFET_GATE_10uA.t23 GNDA 0.0233f
C1016 bgr_11_0.PFET_GATE_10uA.t16 GNDA 0.0233f
C1017 bgr_11_0.PFET_GATE_10uA.n0 GNDA 0.089931f
C1018 bgr_11_0.PFET_GATE_10uA.t28 GNDA 0.020075f
C1019 bgr_11_0.PFET_GATE_10uA.t20 GNDA 0.029676f
C1020 bgr_11_0.PFET_GATE_10uA.n1 GNDA 0.032699f
C1021 bgr_11_0.PFET_GATE_10uA.t13 GNDA 0.020075f
C1022 bgr_11_0.PFET_GATE_10uA.t21 GNDA 0.029676f
C1023 bgr_11_0.PFET_GATE_10uA.n2 GNDA 0.032699f
C1024 bgr_11_0.PFET_GATE_10uA.n3 GNDA 0.032212f
C1025 bgr_11_0.PFET_GATE_10uA.n4 GNDA 0.671121f
C1026 bgr_11_0.PFET_GATE_10uA.t11 GNDA 0.020075f
C1027 bgr_11_0.PFET_GATE_10uA.t25 GNDA 0.029676f
C1028 bgr_11_0.PFET_GATE_10uA.n5 GNDA 0.032699f
C1029 bgr_11_0.PFET_GATE_10uA.t17 GNDA 0.020075f
C1030 bgr_11_0.PFET_GATE_10uA.t26 GNDA 0.029676f
C1031 bgr_11_0.PFET_GATE_10uA.n6 GNDA 0.032699f
C1032 bgr_11_0.PFET_GATE_10uA.n7 GNDA 0.034608f
C1033 bgr_11_0.PFET_GATE_10uA.t6 GNDA 0.304658f
C1034 bgr_11_0.PFET_GATE_10uA.t9 GNDA 0.020589f
C1035 bgr_11_0.PFET_GATE_10uA.t4 GNDA 0.020589f
C1036 bgr_11_0.PFET_GATE_10uA.n8 GNDA 0.052625f
C1037 bgr_11_0.PFET_GATE_10uA.t3 GNDA 0.020589f
C1038 bgr_11_0.PFET_GATE_10uA.t2 GNDA 0.020589f
C1039 bgr_11_0.PFET_GATE_10uA.n9 GNDA 0.051265f
C1040 bgr_11_0.PFET_GATE_10uA.n10 GNDA 0.501438f
C1041 bgr_11_0.PFET_GATE_10uA.t0 GNDA 0.020589f
C1042 bgr_11_0.PFET_GATE_10uA.t8 GNDA 0.020589f
C1043 bgr_11_0.PFET_GATE_10uA.n11 GNDA 0.051265f
C1044 bgr_11_0.PFET_GATE_10uA.n12 GNDA 0.284342f
C1045 bgr_11_0.PFET_GATE_10uA.n13 GNDA 0.61157f
C1046 bgr_11_0.PFET_GATE_10uA.t5 GNDA 0.020589f
C1047 bgr_11_0.PFET_GATE_10uA.t7 GNDA 0.020589f
C1048 bgr_11_0.PFET_GATE_10uA.n14 GNDA 0.049657f
C1049 bgr_11_0.PFET_GATE_10uA.n15 GNDA 0.310845f
C1050 bgr_11_0.PFET_GATE_10uA.t1 GNDA 0.44755f
C1051 bgr_11_0.PFET_GATE_10uA.t24 GNDA 0.066286f
C1052 bgr_11_0.PFET_GATE_10uA.n16 GNDA 1.83377f
C1053 bgr_11_0.PFET_GATE_10uA.n17 GNDA 0.788794f
C1054 bgr_11_0.PFET_GATE_10uA.n18 GNDA 0.796613f
C1055 bgr_11_0.PFET_GATE_10uA.t10 GNDA 0.020075f
C1056 bgr_11_0.PFET_GATE_10uA.t15 GNDA 0.020075f
C1057 bgr_11_0.PFET_GATE_10uA.t14 GNDA 0.020075f
C1058 bgr_11_0.PFET_GATE_10uA.t22 GNDA 0.029676f
C1059 bgr_11_0.PFET_GATE_10uA.n19 GNDA 0.036725f
C1060 bgr_11_0.PFET_GATE_10uA.n20 GNDA 0.026252f
C1061 bgr_11_0.PFET_GATE_10uA.n21 GNDA 0.020461f
C1062 bgr_11_0.PFET_GATE_10uA.t19 GNDA 0.020075f
C1063 bgr_11_0.PFET_GATE_10uA.t12 GNDA 0.020075f
C1064 bgr_11_0.PFET_GATE_10uA.t27 GNDA 0.020075f
C1065 bgr_11_0.PFET_GATE_10uA.t18 GNDA 0.029676f
C1066 bgr_11_0.PFET_GATE_10uA.n22 GNDA 0.036725f
C1067 bgr_11_0.PFET_GATE_10uA.n23 GNDA 0.026252f
C1068 bgr_11_0.PFET_GATE_10uA.n24 GNDA 0.020461f
C1069 bgr_11_0.PFET_GATE_10uA.n25 GNDA 0.066415f
C1070 two_stage_opamp_dummy_magic_24_0.cap_res_X.t91 GNDA 0.43829f
C1071 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 GNDA 0.439878f
C1072 two_stage_opamp_dummy_magic_24_0.cap_res_X.t55 GNDA 0.43829f
C1073 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 GNDA 0.441726f
C1074 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 GNDA 0.48044f
C1075 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 GNDA 0.43829f
C1076 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 GNDA 0.439878f
C1077 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 GNDA 0.43829f
C1078 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 GNDA 0.439878f
C1079 two_stage_opamp_dummy_magic_24_0.cap_res_X.t87 GNDA 0.43829f
C1080 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 GNDA 0.439878f
C1081 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 GNDA 0.43829f
C1082 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 GNDA 0.439878f
C1083 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 GNDA 0.43829f
C1084 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 GNDA 0.439878f
C1085 two_stage_opamp_dummy_magic_24_0.cap_res_X.t7 GNDA 0.43829f
C1086 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 GNDA 0.439878f
C1087 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 GNDA 0.43829f
C1088 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 GNDA 0.439878f
C1089 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 GNDA 0.43829f
C1090 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 GNDA 0.439878f
C1091 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 GNDA 0.43829f
C1092 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 GNDA 0.439878f
C1093 two_stage_opamp_dummy_magic_24_0.cap_res_X.t11 GNDA 0.43829f
C1094 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 GNDA 0.439878f
C1095 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 GNDA 0.43829f
C1096 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 GNDA 0.439878f
C1097 two_stage_opamp_dummy_magic_24_0.cap_res_X.t49 GNDA 0.43829f
C1098 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 GNDA 0.439878f
C1099 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 GNDA 0.43829f
C1100 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 GNDA 0.439878f
C1101 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 GNDA 0.43829f
C1102 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 GNDA 0.439878f
C1103 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 GNDA 0.43829f
C1104 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 GNDA 0.439878f
C1105 two_stage_opamp_dummy_magic_24_0.cap_res_X.t54 GNDA 0.43829f
C1106 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 GNDA 0.439878f
C1107 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 GNDA 0.43829f
C1108 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 GNDA 0.439878f
C1109 two_stage_opamp_dummy_magic_24_0.cap_res_X.t90 GNDA 0.43829f
C1110 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 GNDA 0.439878f
C1111 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 GNDA 0.43829f
C1112 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 GNDA 0.439878f
C1113 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 GNDA 0.43829f
C1114 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 GNDA 0.439878f
C1115 two_stage_opamp_dummy_magic_24_0.cap_res_X.t83 GNDA 0.43829f
C1116 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 GNDA 0.439878f
C1117 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 GNDA 0.43829f
C1118 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 GNDA 0.439878f
C1119 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 GNDA 0.43829f
C1120 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 GNDA 0.439878f
C1121 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 GNDA 0.43829f
C1122 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 GNDA 0.439878f
C1123 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 GNDA 0.43829f
C1124 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 GNDA 0.439878f
C1125 two_stage_opamp_dummy_magic_24_0.cap_res_X.t46 GNDA 0.43829f
C1126 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 GNDA 0.439878f
C1127 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 GNDA 0.43829f
C1128 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 GNDA 0.439878f
C1129 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 GNDA 0.43829f
C1130 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 GNDA 0.439878f
C1131 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 GNDA 0.43829f
C1132 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 GNDA 0.439878f
C1133 two_stage_opamp_dummy_magic_24_0.cap_res_X.t77 GNDA 0.43829f
C1134 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 GNDA 0.439878f
C1135 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 GNDA 0.43829f
C1136 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 GNDA 0.439878f
C1137 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 GNDA 0.43829f
C1138 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 GNDA 0.459779f
C1139 two_stage_opamp_dummy_magic_24_0.cap_res_X.t110 GNDA 0.43829f
C1140 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 GNDA 0.235414f
C1141 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 GNDA 0.251952f
C1142 two_stage_opamp_dummy_magic_24_0.cap_res_X.t50 GNDA 0.43829f
C1143 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 GNDA 0.235414f
C1144 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 GNDA 0.249919f
C1145 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 GNDA 0.43829f
C1146 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 GNDA 0.235414f
C1147 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 GNDA 0.249919f
C1148 two_stage_opamp_dummy_magic_24_0.cap_res_X.t98 GNDA 0.43829f
C1149 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 GNDA 0.235414f
C1150 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 GNDA 0.249919f
C1151 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 GNDA 0.43829f
C1152 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 GNDA 0.235414f
C1153 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 GNDA 0.249919f
C1154 two_stage_opamp_dummy_magic_24_0.cap_res_X.t40 GNDA 0.43829f
C1155 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 GNDA 0.235414f
C1156 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 GNDA 0.249919f
C1157 two_stage_opamp_dummy_magic_24_0.cap_res_X.t3 GNDA 0.43829f
C1158 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 GNDA 0.235414f
C1159 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 GNDA 0.249919f
C1160 two_stage_opamp_dummy_magic_24_0.cap_res_X.t86 GNDA 0.43829f
C1161 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 GNDA 0.235414f
C1162 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 GNDA 0.249919f
C1163 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 GNDA 0.43829f
C1164 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 GNDA 0.235414f
C1165 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 GNDA 0.249919f
C1166 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 GNDA 0.43829f
C1167 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 GNDA 0.439878f
C1168 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 GNDA 0.211892f
C1169 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 GNDA 0.27331f
C1170 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 GNDA 0.233957f
C1171 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 GNDA 0.296831f
C1172 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 GNDA 0.233957f
C1173 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 GNDA 0.318765f
C1174 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 GNDA 0.233957f
C1175 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 GNDA 0.318765f
C1176 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 GNDA 0.233957f
C1177 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 GNDA 0.318765f
C1178 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 GNDA 0.233957f
C1179 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 GNDA 0.318765f
C1180 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 GNDA 0.233957f
C1181 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 GNDA 0.318765f
C1182 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 GNDA 0.233957f
C1183 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 GNDA 0.318765f
C1184 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 GNDA 0.233957f
C1185 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 GNDA 0.318765f
C1186 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 GNDA 0.233957f
C1187 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 GNDA 0.318765f
C1188 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 GNDA 0.233957f
C1189 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 GNDA 0.318765f
C1190 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 GNDA 0.233957f
C1191 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 GNDA 0.318765f
C1192 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 GNDA 0.233957f
C1193 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 GNDA 0.318765f
C1194 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 GNDA 0.233957f
C1195 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 GNDA 0.318765f
C1196 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 GNDA 0.233957f
C1197 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 GNDA 0.318765f
C1198 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 GNDA 0.233957f
C1199 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 GNDA 0.318765f
C1200 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 GNDA 0.233957f
C1201 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 GNDA 0.318765f
C1202 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 GNDA 0.233957f
C1203 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 GNDA 0.296831f
C1204 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 GNDA 0.436833f
C1205 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 GNDA 0.211892f
C1206 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 GNDA 0.274898f
C1207 two_stage_opamp_dummy_magic_24_0.cap_res_X.t10 GNDA 0.436833f
C1208 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 GNDA 0.211892f
C1209 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 GNDA 0.274898f
C1210 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 GNDA 0.436833f
C1211 two_stage_opamp_dummy_magic_24_0.cap_res_X.t115 GNDA 0.43829f
C1212 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 GNDA 0.235414f
C1213 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 GNDA 0.251376f
C1214 two_stage_opamp_dummy_magic_24_0.cap_res_X.t135 GNDA 0.436833f
C1215 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 GNDA 0.43829f
C1216 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 GNDA 0.235414f
C1217 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 GNDA 0.274898f
C1218 two_stage_opamp_dummy_magic_24_0.cap_res_X.t114 GNDA 0.436833f
C1219 two_stage_opamp_dummy_magic_24_0.cap_res_X.t122 GNDA 0.43829f
C1220 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 GNDA 0.235414f
C1221 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 GNDA 0.274898f
C1222 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 GNDA 0.436833f
C1223 two_stage_opamp_dummy_magic_24_0.cap_res_X.t82 GNDA 0.43829f
C1224 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 GNDA 0.235414f
C1225 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 GNDA 0.274898f
C1226 two_stage_opamp_dummy_magic_24_0.cap_res_X.t95 GNDA 0.436833f
C1227 two_stage_opamp_dummy_magic_24_0.cap_res_X.t101 GNDA 0.43829f
C1228 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 GNDA 0.235414f
C1229 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 GNDA 0.274898f
C1230 two_stage_opamp_dummy_magic_24_0.cap_res_X.t59 GNDA 0.436833f
C1231 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 GNDA 0.43829f
C1232 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 GNDA 0.461812f
C1233 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 GNDA 0.235414f
C1234 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 GNDA 0.274898f
C1235 two_stage_opamp_dummy_magic_24_0.cap_res_X.t30 GNDA 0.436833f
C1236 two_stage_opamp_dummy_magic_24_0.cap_res_X.t51 GNDA 0.43829f
C1237 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 GNDA 0.461812f
C1238 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 GNDA 0.235414f
C1239 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 GNDA 0.274898f
C1240 two_stage_opamp_dummy_magic_24_0.cap_res_X.t127 GNDA 0.436833f
C1241 two_stage_opamp_dummy_magic_24_0.cap_res_X.n36 GNDA 0.274898f
C1242 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 GNDA 0.235414f
C1243 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 GNDA 0.461812f
C1244 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 GNDA 1.07126f
C1245 two_stage_opamp_dummy_magic_24_0.cap_res_X.t0 GNDA 0.384111f
C1246 VOUT-.n1 GNDA 0.078254f
C1247 VOUT-.n4 GNDA 0.05869f
C1248 VOUT-.n5 GNDA 0.097817f
C1249 VOUT-.n6 GNDA 0.05869f
C1250 VOUT-.n7 GNDA 0.05869f
C1251 VOUT-.n9 GNDA 0.03991f
C1252 VOUT-.n11 GNDA 0.03991f
C1253 VOUT-.n13 GNDA 0.078254f
C1254 VOUT-.n14 GNDA 0.03991f
C1255 VOUT-.n16 GNDA 0.03991f
C1256 VOUT-.n18 GNDA 0.051647f
C1257 VOUT-.n19 GNDA 0.074515f
C1258 VOUT-.n20 GNDA 0.072515f
C1259 VOUT-.n21 GNDA 0.051647f
C1260 VOUT-.n22 GNDA 0.051647f
C1261 VOUT-.n23 GNDA 0.072515f
C1262 VOUT-.n24 GNDA 0.072515f
C1263 VOUT-.n25 GNDA 0.051647f
C1264 VOUT-.n26 GNDA 0.082684f
C1265 VOUT-.t13 GNDA 0.046952f
C1266 VOUT-.t4 GNDA 0.046952f
C1267 VOUT-.n27 GNDA 0.096205f
C1268 VOUT-.n28 GNDA 0.248334f
C1269 VOUT-.t10 GNDA 0.046952f
C1270 VOUT-.t3 GNDA 0.046952f
C1271 VOUT-.n29 GNDA 0.096205f
C1272 VOUT-.n30 GNDA 0.245831f
C1273 VOUT-.n31 GNDA 0.059705f
C1274 VOUT-.t16 GNDA 0.046952f
C1275 VOUT-.t11 GNDA 0.046952f
C1276 VOUT-.n32 GNDA 0.096205f
C1277 VOUT-.n33 GNDA 0.245831f
C1278 VOUT-.n34 GNDA 0.033843f
C1279 VOUT-.t18 GNDA 0.046952f
C1280 VOUT-.t9 GNDA 0.046952f
C1281 VOUT-.n35 GNDA 0.096205f
C1282 VOUT-.n36 GNDA 0.245831f
C1283 VOUT-.n37 GNDA 0.033843f
C1284 VOUT-.t2 GNDA 0.046952f
C1285 VOUT-.t12 GNDA 0.046952f
C1286 VOUT-.n38 GNDA 0.096205f
C1287 VOUT-.n39 GNDA 0.248334f
C1288 VOUT-.n40 GNDA 0.059705f
C1289 VOUT-.t1 GNDA 0.046952f
C1290 VOUT-.t8 GNDA 0.046952f
C1291 VOUT-.n41 GNDA 0.096205f
C1292 VOUT-.n42 GNDA 0.245831f
C1293 VOUT-.n43 GNDA 0.039475f
C1294 VOUT-.n44 GNDA 0.023476f
C1295 VOUT-.n45 GNDA 0.023476f
C1296 VOUT-.n46 GNDA 0.039475f
C1297 VOUT-.n47 GNDA 0.072515f
C1298 VOUT-.n48 GNDA 0.101507f
C1299 VOUT-.n49 GNDA 0.126482f
C1300 VOUT-.n50 GNDA 0.177023f
C1301 VOUT-.n51 GNDA 0.051647f
C1302 VOUT-.n52 GNDA 0.084514f
C1303 VOUT-.n53 GNDA 0.051647f
C1304 VOUT-.n54 GNDA 0.084514f
C1305 VOUT-.n55 GNDA 0.051647f
C1306 VOUT-.n56 GNDA 0.051647f
C1307 VOUT-.n57 GNDA 0.051647f
C1308 VOUT-.n58 GNDA 0.084514f
C1309 VOUT-.n59 GNDA 0.051647f
C1310 VOUT-.n60 GNDA 0.077471f
C1311 VOUT-.n61 GNDA 0.251195f
C1312 VOUT-.n62 GNDA 0.244152f
C1313 VOUT-.n64 GNDA 0.078254f
C1314 VOUT-.n65 GNDA 0.037562f
C1315 VOUT-.n66 GNDA 0.665158f
C1316 VOUT-.n69 GNDA 0.05869f
C1317 VOUT-.n70 GNDA 0.05869f
C1318 VOUT-.t87 GNDA 0.318347f
C1319 VOUT-.t55 GNDA 0.313015f
C1320 VOUT-.n71 GNDA 0.209867f
C1321 VOUT-.t135 GNDA 0.313015f
C1322 VOUT-.n72 GNDA 0.136944f
C1323 VOUT-.t115 GNDA 0.318347f
C1324 VOUT-.t86 GNDA 0.313015f
C1325 VOUT-.n73 GNDA 0.209867f
C1326 VOUT-.t34 GNDA 0.313015f
C1327 VOUT-.t105 GNDA 0.317679f
C1328 VOUT-.t71 GNDA 0.317679f
C1329 VOUT-.t154 GNDA 0.317679f
C1330 VOUT-.t117 GNDA 0.317679f
C1331 VOUT-.t90 GNDA 0.317679f
C1332 VOUT-.t59 GNDA 0.317679f
C1333 VOUT-.t138 GNDA 0.317679f
C1334 VOUT-.t107 GNDA 0.317679f
C1335 VOUT-.t47 GNDA 0.317679f
C1336 VOUT-.t128 GNDA 0.317679f
C1337 VOUT-.t25 GNDA 0.313015f
C1338 VOUT-.n74 GNDA 0.210534f
C1339 VOUT-.t78 GNDA 0.313015f
C1340 VOUT-.n75 GNDA 0.269225f
C1341 VOUT-.t136 GNDA 0.313015f
C1342 VOUT-.n76 GNDA 0.269225f
C1343 VOUT-.t36 GNDA 0.313015f
C1344 VOUT-.n77 GNDA 0.269225f
C1345 VOUT-.t89 GNDA 0.313015f
C1346 VOUT-.n78 GNDA 0.269225f
C1347 VOUT-.t116 GNDA 0.313015f
C1348 VOUT-.n79 GNDA 0.269225f
C1349 VOUT-.t153 GNDA 0.313015f
C1350 VOUT-.n80 GNDA 0.269225f
C1351 VOUT-.t58 GNDA 0.313015f
C1352 VOUT-.n81 GNDA 0.269225f
C1353 VOUT-.t104 GNDA 0.313015f
C1354 VOUT-.n82 GNDA 0.269225f
C1355 VOUT-.t133 GNDA 0.313015f
C1356 VOUT-.n83 GNDA 0.269225f
C1357 VOUT-.n84 GNDA 0.254325f
C1358 VOUT-.t110 GNDA 0.318347f
C1359 VOUT-.t19 GNDA 0.313015f
C1360 VOUT-.n85 GNDA 0.209867f
C1361 VOUT-.t113 GNDA 0.313015f
C1362 VOUT-.t80 GNDA 0.318347f
C1363 VOUT-.t29 GNDA 0.313015f
C1364 VOUT-.n86 GNDA 0.209867f
C1365 VOUT-.n87 GNDA 0.254325f
C1366 VOUT-.t28 GNDA 0.318347f
C1367 VOUT-.t129 GNDA 0.313015f
C1368 VOUT-.n88 GNDA 0.209867f
C1369 VOUT-.t83 GNDA 0.313015f
C1370 VOUT-.t149 GNDA 0.318347f
C1371 VOUT-.t52 GNDA 0.313015f
C1372 VOUT-.n89 GNDA 0.209867f
C1373 VOUT-.n90 GNDA 0.254325f
C1374 VOUT-.t131 GNDA 0.318347f
C1375 VOUT-.t101 GNDA 0.313015f
C1376 VOUT-.n91 GNDA 0.209867f
C1377 VOUT-.t54 GNDA 0.313015f
C1378 VOUT-.t111 GNDA 0.318347f
C1379 VOUT-.t148 GNDA 0.313015f
C1380 VOUT-.n92 GNDA 0.209867f
C1381 VOUT-.n93 GNDA 0.254325f
C1382 VOUT-.t33 GNDA 0.318347f
C1383 VOUT-.t134 GNDA 0.313015f
C1384 VOUT-.n94 GNDA 0.209867f
C1385 VOUT-.t92 GNDA 0.313015f
C1386 VOUT-.t152 GNDA 0.318347f
C1387 VOUT-.t57 GNDA 0.313015f
C1388 VOUT-.n95 GNDA 0.209867f
C1389 VOUT-.n96 GNDA 0.254325f
C1390 VOUT-.t102 GNDA 0.318347f
C1391 VOUT-.t68 GNDA 0.313015f
C1392 VOUT-.n97 GNDA 0.209867f
C1393 VOUT-.t88 GNDA 0.313015f
C1394 VOUT-.n98 GNDA 0.136944f
C1395 VOUT-.t66 GNDA 0.318347f
C1396 VOUT-.t21 GNDA 0.313015f
C1397 VOUT-.n99 GNDA 0.209867f
C1398 VOUT-.t48 GNDA 0.313015f
C1399 VOUT-.t50 GNDA 0.317679f
C1400 VOUT-.t147 GNDA 0.317679f
C1401 VOUT-.t139 GNDA 0.318347f
C1402 VOUT-.t24 GNDA 0.313015f
C1403 VOUT-.n100 GNDA 0.204976f
C1404 VOUT-.t30 GNDA 0.317679f
C1405 VOUT-.t106 GNDA 0.318347f
C1406 VOUT-.t123 GNDA 0.313015f
C1407 VOUT-.n101 GNDA 0.204976f
C1408 VOUT-.t127 GNDA 0.317679f
C1409 VOUT-.t72 GNDA 0.318347f
C1410 VOUT-.t94 GNDA 0.313015f
C1411 VOUT-.n102 GNDA 0.204976f
C1412 VOUT-.t98 GNDA 0.317679f
C1413 VOUT-.t56 GNDA 0.317679f
C1414 VOUT-.t62 GNDA 0.317679f
C1415 VOUT-.t75 GNDA 0.317941f
C1416 VOUT-.t79 GNDA 0.317679f
C1417 VOUT-.t35 GNDA 0.317941f
C1418 VOUT-.t43 GNDA 0.317679f
C1419 VOUT-.t155 GNDA 0.317941f
C1420 VOUT-.t22 GNDA 0.317679f
C1421 VOUT-.t42 GNDA 0.317941f
C1422 VOUT-.t49 GNDA 0.317679f
C1423 VOUT-.t144 GNDA 0.313015f
C1424 VOUT-.n103 GNDA 0.346465f
C1425 VOUT-.t120 GNDA 0.313015f
C1426 VOUT-.n104 GNDA 0.405156f
C1427 VOUT-.t137 GNDA 0.313015f
C1428 VOUT-.n105 GNDA 0.405156f
C1429 VOUT-.t41 GNDA 0.313015f
C1430 VOUT-.n106 GNDA 0.405156f
C1431 VOUT-.t151 GNDA 0.313015f
C1432 VOUT-.n107 GNDA 0.401505f
C1433 VOUT-.t61 GNDA 0.313015f
C1434 VOUT-.n108 GNDA 0.332806f
C1435 VOUT-.t97 GNDA 0.313015f
C1436 VOUT-.n109 GNDA 0.332806f
C1437 VOUT-.t125 GNDA 0.313015f
C1438 VOUT-.n110 GNDA 0.332806f
C1439 VOUT-.t109 GNDA 0.313015f
C1440 VOUT-.n111 GNDA 0.269225f
C1441 VOUT-.t145 GNDA 0.313015f
C1442 VOUT-.n112 GNDA 0.269225f
C1443 VOUT-.n113 GNDA 0.254325f
C1444 VOUT-.t99 GNDA 0.318347f
C1445 VOUT-.t65 GNDA 0.313015f
C1446 VOUT-.n114 GNDA 0.209867f
C1447 VOUT-.t81 GNDA 0.313015f
C1448 VOUT-.t143 GNDA 0.318347f
C1449 VOUT-.t44 GNDA 0.313015f
C1450 VOUT-.n115 GNDA 0.209867f
C1451 VOUT-.n116 GNDA 0.254325f
C1452 VOUT-.t70 GNDA 0.318347f
C1453 VOUT-.t32 GNDA 0.313015f
C1454 VOUT-.n117 GNDA 0.209867f
C1455 VOUT-.t118 GNDA 0.313015f
C1456 VOUT-.t60 GNDA 0.318347f
C1457 VOUT-.t91 GNDA 0.313015f
C1458 VOUT-.n118 GNDA 0.209867f
C1459 VOUT-.n119 GNDA 0.254325f
C1460 VOUT-.t27 GNDA 0.318347f
C1461 VOUT-.t130 GNDA 0.313015f
C1462 VOUT-.n120 GNDA 0.209867f
C1463 VOUT-.t84 GNDA 0.313015f
C1464 VOUT-.t150 GNDA 0.318347f
C1465 VOUT-.t53 GNDA 0.313015f
C1466 VOUT-.n121 GNDA 0.209867f
C1467 VOUT-.n122 GNDA 0.254325f
C1468 VOUT-.t69 GNDA 0.318347f
C1469 VOUT-.t26 GNDA 0.313015f
C1470 VOUT-.n123 GNDA 0.209867f
C1471 VOUT-.t112 GNDA 0.313015f
C1472 VOUT-.t51 GNDA 0.318347f
C1473 VOUT-.t82 GNDA 0.313015f
C1474 VOUT-.n124 GNDA 0.209867f
C1475 VOUT-.n125 GNDA 0.254325f
C1476 VOUT-.t23 GNDA 0.318347f
C1477 VOUT-.t124 GNDA 0.313015f
C1478 VOUT-.n126 GNDA 0.209867f
C1479 VOUT-.t76 GNDA 0.313015f
C1480 VOUT-.t146 GNDA 0.318347f
C1481 VOUT-.t45 GNDA 0.313015f
C1482 VOUT-.n127 GNDA 0.209867f
C1483 VOUT-.n128 GNDA 0.254325f
C1484 VOUT-.t121 GNDA 0.318347f
C1485 VOUT-.t93 GNDA 0.313015f
C1486 VOUT-.n129 GNDA 0.209867f
C1487 VOUT-.t38 GNDA 0.313015f
C1488 VOUT-.t108 GNDA 0.318347f
C1489 VOUT-.t141 GNDA 0.313015f
C1490 VOUT-.n130 GNDA 0.209867f
C1491 VOUT-.n131 GNDA 0.254325f
C1492 VOUT-.t156 GNDA 0.318347f
C1493 VOUT-.t119 GNDA 0.313015f
C1494 VOUT-.n132 GNDA 0.209867f
C1495 VOUT-.t73 GNDA 0.313015f
C1496 VOUT-.t140 GNDA 0.318347f
C1497 VOUT-.t37 GNDA 0.313015f
C1498 VOUT-.n133 GNDA 0.209867f
C1499 VOUT-.n134 GNDA 0.254325f
C1500 VOUT-.t114 GNDA 0.318347f
C1501 VOUT-.t85 GNDA 0.313015f
C1502 VOUT-.n135 GNDA 0.209867f
C1503 VOUT-.t31 GNDA 0.313015f
C1504 VOUT-.t103 GNDA 0.318347f
C1505 VOUT-.t132 GNDA 0.313015f
C1506 VOUT-.n136 GNDA 0.209867f
C1507 VOUT-.n137 GNDA 0.254325f
C1508 VOUT-.t77 GNDA 0.318347f
C1509 VOUT-.t46 GNDA 0.313015f
C1510 VOUT-.n138 GNDA 0.209867f
C1511 VOUT-.t126 GNDA 0.313015f
C1512 VOUT-.t67 GNDA 0.318347f
C1513 VOUT-.t100 GNDA 0.313015f
C1514 VOUT-.n139 GNDA 0.209867f
C1515 VOUT-.n140 GNDA 0.254325f
C1516 VOUT-.t40 GNDA 0.318347f
C1517 VOUT-.t142 GNDA 0.313015f
C1518 VOUT-.n141 GNDA 0.209867f
C1519 VOUT-.t96 GNDA 0.313015f
C1520 VOUT-.t20 GNDA 0.318347f
C1521 VOUT-.t64 GNDA 0.313015f
C1522 VOUT-.n142 GNDA 0.209867f
C1523 VOUT-.n143 GNDA 0.254325f
C1524 VOUT-.t74 GNDA 0.318347f
C1525 VOUT-.t39 GNDA 0.313015f
C1526 VOUT-.n144 GNDA 0.209867f
C1527 VOUT-.t122 GNDA 0.313015f
C1528 VOUT-.n145 GNDA 0.254325f
C1529 VOUT-.t95 GNDA 0.313015f
C1530 VOUT-.n146 GNDA 0.133506f
C1531 VOUT-.t63 GNDA 0.313015f
C1532 VOUT-.n147 GNDA 0.262654f
C1533 VOUT-.n148 GNDA 0.196613f
C1534 VOUT-.n149 GNDA 0.05869f
C1535 VOUT-.n150 GNDA 0.05869f
C1536 VOUT-.n151 GNDA 0.05869f
C1537 VOUT-.n152 GNDA 0.172148f
C1538 VOUT-.n153 GNDA 0.06218f
C1539 VOUT-.n154 GNDA 0.059123f
C1540 VOUT-.n156 GNDA 0.674939f
C1541 VOUT-.n157 GNDA 0.05869f
C1542 VOUT-.n158 GNDA 0.709175f
C1543 VOUT-.n162 GNDA 0.03991f
C1544 VOUT-.n163 GNDA 0.03991f
C1545 VOUT-.n164 GNDA 0.037562f
C1546 VOUT-.n165 GNDA 0.078254f
C1547 VOUT-.n166 GNDA 0.03991f
C1548 VOUT-.n167 GNDA 0.03991f
C1549 VOUT-.n169 GNDA 0.699394f
C1550 VOUT-.n170 GNDA 0.065733f
C1551 VOUT-.n171 GNDA 0.037562f
C1552 VOUT-.t15 GNDA 0.054778f
C1553 VOUT-.t5 GNDA 0.054778f
C1554 VOUT-.n172 GNDA 0.117696f
C1555 VOUT-.n173 GNDA 0.283057f
C1556 VOUT-.n174 GNDA 0.037562f
C1557 VOUT-.n175 GNDA 0.242565f
C1558 VOUT-.t7 GNDA 0.054778f
C1559 VOUT-.t14 GNDA 0.054778f
C1560 VOUT-.n176 GNDA 0.117696f
C1561 VOUT-.n177 GNDA 0.292945f
C1562 VOUT-.n178 GNDA 0.167445f
C1563 VOUT-.t0 GNDA 0.054778f
C1564 VOUT-.t6 GNDA 0.054778f
C1565 VOUT-.n179 GNDA 0.117696f
C1566 VOUT-.n180 GNDA 0.278295f
C1567 VOUT-.n181 GNDA 0.127717f
C1568 VOUT-.n182 GNDA 0.037562f
C1569 VOUT-.n183 GNDA 0.193823f
C1570 VOUT-.n184 GNDA 0.037562f
C1571 VOUT-.n185 GNDA 0.037562f
C1572 VOUT-.n186 GNDA 0.037562f
C1573 VOUT-.n187 GNDA 0.037562f
C1574 VOUT-.n188 GNDA 0.080406f
C1575 VOUT-.n189 GNDA 0.145552f
C1576 VOUT-.t17 GNDA 0.089346f
C1577 VOUT-.n190 GNDA 0.289403f
C1578 bgr_11_0.V_TOP.t31 GNDA 0.101858f
C1579 bgr_11_0.V_TOP.t40 GNDA 0.101858f
C1580 bgr_11_0.V_TOP.t47 GNDA 0.101858f
C1581 bgr_11_0.V_TOP.t23 GNDA 0.101858f
C1582 bgr_11_0.V_TOP.t21 GNDA 0.101858f
C1583 bgr_11_0.V_TOP.t33 GNDA 0.101858f
C1584 bgr_11_0.V_TOP.t41 GNDA 0.101858f
C1585 bgr_11_0.V_TOP.t49 GNDA 0.101858f
C1586 bgr_11_0.V_TOP.t27 GNDA 0.101858f
C1587 bgr_11_0.V_TOP.t25 GNDA 0.101858f
C1588 bgr_11_0.V_TOP.t37 GNDA 0.101858f
C1589 bgr_11_0.V_TOP.t44 GNDA 0.101858f
C1590 bgr_11_0.V_TOP.t19 GNDA 0.101858f
C1591 bgr_11_0.V_TOP.t36 GNDA 0.101858f
C1592 bgr_11_0.V_TOP.t34 GNDA 0.133153f
C1593 bgr_11_0.V_TOP.n0 GNDA 0.074443f
C1594 bgr_11_0.V_TOP.n1 GNDA 0.054324f
C1595 bgr_11_0.V_TOP.n2 GNDA 0.054324f
C1596 bgr_11_0.V_TOP.n3 GNDA 0.054324f
C1597 bgr_11_0.V_TOP.n4 GNDA 0.054324f
C1598 bgr_11_0.V_TOP.n5 GNDA 0.050658f
C1599 bgr_11_0.V_TOP.t12 GNDA 0.132092f
C1600 bgr_11_0.V_TOP.t22 GNDA 0.38803f
C1601 bgr_11_0.V_TOP.t26 GNDA 0.394639f
C1602 bgr_11_0.V_TOP.t32 GNDA 0.38803f
C1603 bgr_11_0.V_TOP.n6 GNDA 0.260161f
C1604 bgr_11_0.V_TOP.t20 GNDA 0.38803f
C1605 bgr_11_0.V_TOP.t46 GNDA 0.394639f
C1606 bgr_11_0.V_TOP.n7 GNDA 0.332917f
C1607 bgr_11_0.V_TOP.t35 GNDA 0.394639f
C1608 bgr_11_0.V_TOP.t39 GNDA 0.38803f
C1609 bgr_11_0.V_TOP.n8 GNDA 0.260161f
C1610 bgr_11_0.V_TOP.t30 GNDA 0.38803f
C1611 bgr_11_0.V_TOP.t18 GNDA 0.394639f
C1612 bgr_11_0.V_TOP.n9 GNDA 0.405673f
C1613 bgr_11_0.V_TOP.t24 GNDA 0.394639f
C1614 bgr_11_0.V_TOP.t29 GNDA 0.38803f
C1615 bgr_11_0.V_TOP.n10 GNDA 0.260161f
C1616 bgr_11_0.V_TOP.t17 GNDA 0.38803f
C1617 bgr_11_0.V_TOP.t45 GNDA 0.394639f
C1618 bgr_11_0.V_TOP.n11 GNDA 0.405673f
C1619 bgr_11_0.V_TOP.t48 GNDA 0.394639f
C1620 bgr_11_0.V_TOP.t16 GNDA 0.38803f
C1621 bgr_11_0.V_TOP.n12 GNDA 0.260161f
C1622 bgr_11_0.V_TOP.t43 GNDA 0.38803f
C1623 bgr_11_0.V_TOP.t38 GNDA 0.394639f
C1624 bgr_11_0.V_TOP.n13 GNDA 0.405673f
C1625 bgr_11_0.V_TOP.t42 GNDA 0.394639f
C1626 bgr_11_0.V_TOP.t14 GNDA 0.38803f
C1627 bgr_11_0.V_TOP.n14 GNDA 0.332917f
C1628 bgr_11_0.V_TOP.t28 GNDA 0.38803f
C1629 bgr_11_0.V_TOP.n15 GNDA 0.169763f
C1630 bgr_11_0.V_TOP.n16 GNDA 0.58097f
C1631 bgr_11_0.V_TOP.t13 GNDA 0.109158f
C1632 bgr_11_0.V_TOP.n17 GNDA 0.757626f
C1633 bgr_11_0.V_TOP.n18 GNDA 0.024154f
C1634 bgr_11_0.V_TOP.n19 GNDA 0.428712f
C1635 bgr_11_0.V_TOP.n20 GNDA 0.023396f
C1636 bgr_11_0.V_TOP.n21 GNDA 0.024317f
C1637 bgr_11_0.V_TOP.n22 GNDA 0.024154f
C1638 bgr_11_0.V_TOP.n23 GNDA 0.233507f
C1639 bgr_11_0.V_TOP.n24 GNDA 0.155412f
C1640 bgr_11_0.V_TOP.n25 GNDA 0.077606f
C1641 bgr_11_0.V_TOP.n26 GNDA 0.024154f
C1642 bgr_11_0.V_TOP.n27 GNDA 0.133969f
C1643 bgr_11_0.V_TOP.n28 GNDA 0.024154f
C1644 bgr_11_0.V_TOP.n29 GNDA 0.132695f
C1645 bgr_11_0.V_TOP.n30 GNDA 0.335602f
C1646 bgr_11_0.V_TOP.n31 GNDA 0.021099f
C1647 bgr_11_0.V_TOP.n32 GNDA 0.050658f
C1648 bgr_11_0.V_TOP.n33 GNDA 0.054324f
C1649 bgr_11_0.V_TOP.n34 GNDA 0.054324f
C1650 bgr_11_0.V_TOP.n35 GNDA 0.054324f
C1651 bgr_11_0.V_TOP.n36 GNDA 0.054324f
C1652 bgr_11_0.V_TOP.n37 GNDA 0.054324f
C1653 bgr_11_0.V_TOP.n38 GNDA 0.054324f
C1654 bgr_11_0.V_TOP.n39 GNDA 0.050658f
C1655 bgr_11_0.V_TOP.t15 GNDA 0.117376f
C1656 bgr_11_0.1st_Vout_1.n0 GNDA 1.44728f
C1657 bgr_11_0.1st_Vout_1.n1 GNDA 0.436509f
C1658 bgr_11_0.1st_Vout_1.n2 GNDA 0.980114f
C1659 bgr_11_0.1st_Vout_1.n3 GNDA 0.098275f
C1660 bgr_11_0.1st_Vout_1.n4 GNDA 0.151675f
C1661 bgr_11_0.1st_Vout_1.t30 GNDA 0.290456f
C1662 bgr_11_0.1st_Vout_1.t19 GNDA 0.285592f
C1663 bgr_11_0.1st_Vout_1.t15 GNDA 0.290456f
C1664 bgr_11_0.1st_Vout_1.t26 GNDA 0.285592f
C1665 bgr_11_0.1st_Vout_1.t32 GNDA 0.290456f
C1666 bgr_11_0.1st_Vout_1.t29 GNDA 0.285592f
C1667 bgr_11_0.1st_Vout_1.t25 GNDA 0.290456f
C1668 bgr_11_0.1st_Vout_1.t31 GNDA 0.285592f
C1669 bgr_11_0.1st_Vout_1.t28 GNDA 0.290456f
C1670 bgr_11_0.1st_Vout_1.t18 GNDA 0.285592f
C1671 bgr_11_0.1st_Vout_1.t14 GNDA 0.290456f
C1672 bgr_11_0.1st_Vout_1.t23 GNDA 0.285592f
C1673 bgr_11_0.1st_Vout_1.t17 GNDA 0.290456f
C1674 bgr_11_0.1st_Vout_1.t10 GNDA 0.285592f
C1675 bgr_11_0.1st_Vout_1.t8 GNDA 0.290456f
C1676 bgr_11_0.1st_Vout_1.t13 GNDA 0.285592f
C1677 bgr_11_0.1st_Vout_1.t27 GNDA 0.290456f
C1678 bgr_11_0.1st_Vout_1.t16 GNDA 0.285592f
C1679 bgr_11_0.1st_Vout_1.t21 GNDA 0.285592f
C1680 bgr_11_0.1st_Vout_1.t12 GNDA 0.285592f
C1681 bgr_11_0.1st_Vout_1.t22 GNDA 0.018657f
C1682 bgr_11_0.1st_Vout_1.n5 GNDA 0.568592f
C1683 bgr_11_0.1st_Vout_1.n6 GNDA 0.017998f
C1684 bgr_11_0.1st_Vout_1.t11 GNDA 0.010877f
C1685 bgr_11_0.1st_Vout_1.t20 GNDA 0.010877f
C1686 bgr_11_0.1st_Vout_1.n7 GNDA 0.024196f
C1687 bgr_11_0.1st_Vout_1.t0 GNDA 0.097022f
C1688 bgr_11_0.1st_Vout_1.n8 GNDA 0.017252f
C1689 bgr_11_0.1st_Vout_1.n9 GNDA 0.104204f
C1690 bgr_11_0.1st_Vout_1.t7 GNDA 0.010877f
C1691 bgr_11_0.1st_Vout_1.t24 GNDA 0.010877f
C1692 bgr_11_0.1st_Vout_1.n10 GNDA 0.024196f
C1693 bgr_11_0.1st_Vout_1.n11 GNDA 0.017998f
C1694 bgr_11_0.1st_Vout_1.t9 GNDA 0.017072f
C1695 two_stage_opamp_dummy_magic_24_0.VD2.n0 GNDA 0.226102f
C1696 two_stage_opamp_dummy_magic_24_0.VD2.n1 GNDA 0.077257f
C1697 two_stage_opamp_dummy_magic_24_0.VD2.n2 GNDA 0.103687f
C1698 two_stage_opamp_dummy_magic_24_0.VD2.t3 GNDA 0.051486f
C1699 two_stage_opamp_dummy_magic_24_0.VD2.t5 GNDA 0.051486f
C1700 two_stage_opamp_dummy_magic_24_0.VD2.n3 GNDA 0.112028f
C1701 two_stage_opamp_dummy_magic_24_0.VD2.n4 GNDA 0.431638f
C1702 two_stage_opamp_dummy_magic_24_0.VD2.n5 GNDA 0.109497f
C1703 two_stage_opamp_dummy_magic_24_0.VD2.t1 GNDA 0.051486f
C1704 two_stage_opamp_dummy_magic_24_0.VD2.t10 GNDA 0.051486f
C1705 two_stage_opamp_dummy_magic_24_0.VD2.n6 GNDA 0.112028f
C1706 two_stage_opamp_dummy_magic_24_0.VD2.n7 GNDA 0.443673f
C1707 two_stage_opamp_dummy_magic_24_0.VD2.t12 GNDA 0.051486f
C1708 two_stage_opamp_dummy_magic_24_0.VD2.t18 GNDA 0.051486f
C1709 two_stage_opamp_dummy_magic_24_0.VD2.n8 GNDA 0.112028f
C1710 two_stage_opamp_dummy_magic_24_0.VD2.n9 GNDA 0.357994f
C1711 two_stage_opamp_dummy_magic_24_0.VD2.n10 GNDA 0.102973f
C1712 two_stage_opamp_dummy_magic_24_0.VD2.t16 GNDA 0.051486f
C1713 two_stage_opamp_dummy_magic_24_0.VD2.t11 GNDA 0.051486f
C1714 two_stage_opamp_dummy_magic_24_0.VD2.n11 GNDA 0.112028f
C1715 two_stage_opamp_dummy_magic_24_0.VD2.n12 GNDA 0.357994f
C1716 two_stage_opamp_dummy_magic_24_0.VD2.n13 GNDA 0.103687f
C1717 two_stage_opamp_dummy_magic_24_0.VD2.t9 GNDA 0.051486f
C1718 two_stage_opamp_dummy_magic_24_0.VD2.t4 GNDA 0.051486f
C1719 two_stage_opamp_dummy_magic_24_0.VD2.n14 GNDA 0.112028f
C1720 two_stage_opamp_dummy_magic_24_0.VD2.n15 GNDA 0.443673f
C1721 two_stage_opamp_dummy_magic_24_0.VD2.n16 GNDA 0.186124f
C1722 two_stage_opamp_dummy_magic_24_0.VD2.t0 GNDA 0.051486f
C1723 two_stage_opamp_dummy_magic_24_0.VD2.t8 GNDA 0.051486f
C1724 two_stage_opamp_dummy_magic_24_0.VD2.n17 GNDA 0.112028f
C1725 two_stage_opamp_dummy_magic_24_0.VD2.n18 GNDA 0.431638f
C1726 two_stage_opamp_dummy_magic_24_0.VD2.n19 GNDA 0.077257f
C1727 two_stage_opamp_dummy_magic_24_0.VD2.n20 GNDA 0.172945f
C1728 two_stage_opamp_dummy_magic_24_0.VD2.n21 GNDA 0.393891f
C1729 two_stage_opamp_dummy_magic_24_0.VD2.n22 GNDA 0.173147f
C1730 two_stage_opamp_dummy_magic_24_0.VD2.n23 GNDA 0.385119f
C1731 two_stage_opamp_dummy_magic_24_0.VD2.t14 GNDA 0.051486f
C1732 two_stage_opamp_dummy_magic_24_0.VD2.t17 GNDA 0.051486f
C1733 two_stage_opamp_dummy_magic_24_0.VD2.n24 GNDA 0.112028f
C1734 two_stage_opamp_dummy_magic_24_0.VD2.n25 GNDA 0.348896f
C1735 two_stage_opamp_dummy_magic_24_0.VD2.n26 GNDA 0.19689f
C1736 two_stage_opamp_dummy_magic_24_0.VD2.t15 GNDA 0.051486f
C1737 two_stage_opamp_dummy_magic_24_0.VD2.t20 GNDA 0.051486f
C1738 two_stage_opamp_dummy_magic_24_0.VD2.n27 GNDA 0.112028f
C1739 two_stage_opamp_dummy_magic_24_0.VD2.n28 GNDA 0.348896f
C1740 two_stage_opamp_dummy_magic_24_0.VD2.n29 GNDA 0.115007f
C1741 two_stage_opamp_dummy_magic_24_0.VD2.n30 GNDA 0.19689f
C1742 two_stage_opamp_dummy_magic_24_0.VD2.t13 GNDA 0.051486f
C1743 two_stage_opamp_dummy_magic_24_0.VD2.t19 GNDA 0.051486f
C1744 two_stage_opamp_dummy_magic_24_0.VD2.n31 GNDA 0.112028f
C1745 two_stage_opamp_dummy_magic_24_0.VD2.n32 GNDA 0.348896f
C1746 two_stage_opamp_dummy_magic_24_0.VD2.n33 GNDA 0.385119f
C1747 two_stage_opamp_dummy_magic_24_0.VD2.n34 GNDA 0.173147f
C1748 two_stage_opamp_dummy_magic_24_0.VD2.n35 GNDA 0.393891f
C1749 two_stage_opamp_dummy_magic_24_0.VD2.n36 GNDA 0.172945f
C1750 two_stage_opamp_dummy_magic_24_0.VD2.n37 GNDA 0.077257f
C1751 two_stage_opamp_dummy_magic_24_0.VD2.t21 GNDA 0.051486f
C1752 two_stage_opamp_dummy_magic_24_0.VD2.t6 GNDA 0.051486f
C1753 two_stage_opamp_dummy_magic_24_0.VD2.n38 GNDA 0.112028f
C1754 two_stage_opamp_dummy_magic_24_0.VD2.n39 GNDA 0.431638f
C1755 two_stage_opamp_dummy_magic_24_0.VD2.n40 GNDA 0.186124f
C1756 two_stage_opamp_dummy_magic_24_0.VD2.n41 GNDA 0.109497f
C1757 two_stage_opamp_dummy_magic_24_0.VD2.t2 GNDA 0.051486f
C1758 two_stage_opamp_dummy_magic_24_0.VD2.t7 GNDA 0.051486f
C1759 two_stage_opamp_dummy_magic_24_0.VD2.n42 GNDA 0.112028f
C1760 two_stage_opamp_dummy_magic_24_0.VD2.n43 GNDA 0.431638f
C1761 two_stage_opamp_dummy_magic_24_0.VD2.n44 GNDA 0.077257f
C1762 two_stage_opamp_dummy_magic_24_0.VD2.n45 GNDA 0.059795f
C1763 two_stage_opamp_dummy_magic_24_0.Y.n0 GNDA 0.080325f
C1764 two_stage_opamp_dummy_magic_24_0.Y.n1 GNDA 0.103691f
C1765 two_stage_opamp_dummy_magic_24_0.Y.n2 GNDA 0.098175f
C1766 two_stage_opamp_dummy_magic_24_0.Y.n3 GNDA 0.098175f
C1767 two_stage_opamp_dummy_magic_24_0.Y.n4 GNDA 0.098175f
C1768 two_stage_opamp_dummy_magic_24_0.Y.n5 GNDA 0.103691f
C1769 two_stage_opamp_dummy_magic_24_0.Y.t14 GNDA 0.022313f
C1770 two_stage_opamp_dummy_magic_24_0.Y.t12 GNDA 0.022313f
C1771 two_stage_opamp_dummy_magic_24_0.Y.n6 GNDA 0.048549f
C1772 two_stage_opamp_dummy_magic_24_0.Y.n7 GNDA 0.155143f
C1773 two_stage_opamp_dummy_magic_24_0.Y.n8 GNDA 0.075036f
C1774 two_stage_opamp_dummy_magic_24_0.Y.n9 GNDA 0.177012f
C1775 two_stage_opamp_dummy_magic_24_0.Y.t11 GNDA 0.022313f
C1776 two_stage_opamp_dummy_magic_24_0.Y.t16 GNDA 0.022313f
C1777 two_stage_opamp_dummy_magic_24_0.Y.n10 GNDA 0.048549f
C1778 two_stage_opamp_dummy_magic_24_0.Y.n11 GNDA 0.155143f
C1779 two_stage_opamp_dummy_magic_24_0.Y.n12 GNDA 0.121089f
C1780 two_stage_opamp_dummy_magic_24_0.Y.n13 GNDA 0.258718f
C1781 two_stage_opamp_dummy_magic_24_0.Y.n14 GNDA 0.098175f
C1782 two_stage_opamp_dummy_magic_24_0.Y.n15 GNDA 0.336497f
C1783 two_stage_opamp_dummy_magic_24_0.Y.n16 GNDA 0.098175f
C1784 two_stage_opamp_dummy_magic_24_0.Y.n17 GNDA 0.209313f
C1785 two_stage_opamp_dummy_magic_24_0.Y.n18 GNDA 0.103691f
C1786 two_stage_opamp_dummy_magic_24_0.Y.t20 GNDA 0.022313f
C1787 two_stage_opamp_dummy_magic_24_0.Y.t18 GNDA 0.022313f
C1788 two_stage_opamp_dummy_magic_24_0.Y.n19 GNDA 0.048549f
C1789 two_stage_opamp_dummy_magic_24_0.Y.n20 GNDA 0.1512f
C1790 two_stage_opamp_dummy_magic_24_0.Y.n21 GNDA 0.085325f
C1791 two_stage_opamp_dummy_magic_24_0.Y.t15 GNDA 0.022313f
C1792 two_stage_opamp_dummy_magic_24_0.Y.t21 GNDA 0.022313f
C1793 two_stage_opamp_dummy_magic_24_0.Y.n22 GNDA 0.048549f
C1794 two_stage_opamp_dummy_magic_24_0.Y.n23 GNDA 0.1512f
C1795 two_stage_opamp_dummy_magic_24_0.Y.n24 GNDA 0.085325f
C1796 two_stage_opamp_dummy_magic_24_0.Y.t13 GNDA 0.022313f
C1797 two_stage_opamp_dummy_magic_24_0.Y.t22 GNDA 0.022313f
C1798 two_stage_opamp_dummy_magic_24_0.Y.n25 GNDA 0.048549f
C1799 two_stage_opamp_dummy_magic_24_0.Y.n26 GNDA 0.1512f
C1800 two_stage_opamp_dummy_magic_24_0.Y.n27 GNDA 0.04984f
C1801 two_stage_opamp_dummy_magic_24_0.Y.n28 GNDA 0.04984f
C1802 two_stage_opamp_dummy_magic_24_0.Y.t17 GNDA 0.022313f
C1803 two_stage_opamp_dummy_magic_24_0.Y.t19 GNDA 0.022313f
C1804 two_stage_opamp_dummy_magic_24_0.Y.n29 GNDA 0.048549f
C1805 two_stage_opamp_dummy_magic_24_0.Y.n30 GNDA 0.1512f
C1806 two_stage_opamp_dummy_magic_24_0.Y.n31 GNDA 0.103691f
C1807 two_stage_opamp_dummy_magic_24_0.Y.n32 GNDA 0.044625f
C1808 two_stage_opamp_dummy_magic_24_0.Y.n33 GNDA 0.044625f
C1809 two_stage_opamp_dummy_magic_24_0.Y.n34 GNDA 0.075036f
C1810 two_stage_opamp_dummy_magic_24_0.Y.n35 GNDA 0.107492f
C1811 two_stage_opamp_dummy_magic_24_0.Y.n36 GNDA 0.0714f
C1812 two_stage_opamp_dummy_magic_24_0.Y.t26 GNDA 0.047972f
C1813 two_stage_opamp_dummy_magic_24_0.Y.t43 GNDA 0.047972f
C1814 two_stage_opamp_dummy_magic_24_0.Y.t31 GNDA 0.047972f
C1815 two_stage_opamp_dummy_magic_24_0.Y.t46 GNDA 0.047972f
C1816 two_stage_opamp_dummy_magic_24_0.Y.t33 GNDA 0.047972f
C1817 two_stage_opamp_dummy_magic_24_0.Y.t48 GNDA 0.047972f
C1818 two_stage_opamp_dummy_magic_24_0.Y.t35 GNDA 0.047972f
C1819 two_stage_opamp_dummy_magic_24_0.Y.t50 GNDA 0.054536f
C1820 two_stage_opamp_dummy_magic_24_0.Y.n39 GNDA 0.049217f
C1821 two_stage_opamp_dummy_magic_24_0.Y.n40 GNDA 0.030122f
C1822 two_stage_opamp_dummy_magic_24_0.Y.n41 GNDA 0.030122f
C1823 two_stage_opamp_dummy_magic_24_0.Y.n42 GNDA 0.030122f
C1824 two_stage_opamp_dummy_magic_24_0.Y.n43 GNDA 0.030122f
C1825 two_stage_opamp_dummy_magic_24_0.Y.n44 GNDA 0.030122f
C1826 two_stage_opamp_dummy_magic_24_0.Y.n45 GNDA 0.02538f
C1827 two_stage_opamp_dummy_magic_24_0.Y.t40 GNDA 0.047972f
C1828 two_stage_opamp_dummy_magic_24_0.Y.t27 GNDA 0.054536f
C1829 two_stage_opamp_dummy_magic_24_0.Y.n46 GNDA 0.044476f
C1830 two_stage_opamp_dummy_magic_24_0.Y.n47 GNDA 0.012324f
C1831 two_stage_opamp_dummy_magic_24_0.Y.t29 GNDA 0.031237f
C1832 two_stage_opamp_dummy_magic_24_0.Y.t45 GNDA 0.031237f
C1833 two_stage_opamp_dummy_magic_24_0.Y.t32 GNDA 0.031237f
C1834 two_stage_opamp_dummy_magic_24_0.Y.t47 GNDA 0.031237f
C1835 two_stage_opamp_dummy_magic_24_0.Y.t34 GNDA 0.031237f
C1836 two_stage_opamp_dummy_magic_24_0.Y.t49 GNDA 0.031237f
C1837 two_stage_opamp_dummy_magic_24_0.Y.t37 GNDA 0.031237f
C1838 two_stage_opamp_dummy_magic_24_0.Y.t53 GNDA 0.037931f
C1839 two_stage_opamp_dummy_magic_24_0.Y.n48 GNDA 0.037931f
C1840 two_stage_opamp_dummy_magic_24_0.Y.n49 GNDA 0.024544f
C1841 two_stage_opamp_dummy_magic_24_0.Y.n50 GNDA 0.024544f
C1842 two_stage_opamp_dummy_magic_24_0.Y.n51 GNDA 0.024544f
C1843 two_stage_opamp_dummy_magic_24_0.Y.n52 GNDA 0.024544f
C1844 two_stage_opamp_dummy_magic_24_0.Y.n53 GNDA 0.024544f
C1845 two_stage_opamp_dummy_magic_24_0.Y.n54 GNDA 0.019802f
C1846 two_stage_opamp_dummy_magic_24_0.Y.t42 GNDA 0.031237f
C1847 two_stage_opamp_dummy_magic_24_0.Y.t30 GNDA 0.037931f
C1848 two_stage_opamp_dummy_magic_24_0.Y.n55 GNDA 0.03319f
C1849 two_stage_opamp_dummy_magic_24_0.Y.n56 GNDA 0.012324f
C1850 two_stage_opamp_dummy_magic_24_0.Y.n57 GNDA 0.07218f
C1851 two_stage_opamp_dummy_magic_24_0.Y.n58 GNDA 0.0714f
C1852 two_stage_opamp_dummy_magic_24_0.Y.n59 GNDA 0.070729f
C1853 two_stage_opamp_dummy_magic_24_0.Y.n60 GNDA 0.0714f
C1854 two_stage_opamp_dummy_magic_24_0.Y.t10 GNDA 0.618914f
C1855 two_stage_opamp_dummy_magic_24_0.Y.n61 GNDA 0.0714f
C1856 two_stage_opamp_dummy_magic_24_0.Y.n62 GNDA 0.0714f
C1857 two_stage_opamp_dummy_magic_24_0.Y.n64 GNDA 0.647244f
C1858 two_stage_opamp_dummy_magic_24_0.Y.n66 GNDA 0.798786f
C1859 two_stage_opamp_dummy_magic_24_0.Y.n67 GNDA 0.023642f
C1860 two_stage_opamp_dummy_magic_24_0.Y.n68 GNDA 0.0238f
C1861 two_stage_opamp_dummy_magic_24_0.Y.n69 GNDA 0.0238f
C1862 two_stage_opamp_dummy_magic_24_0.Y.t39 GNDA 0.098175f
C1863 two_stage_opamp_dummy_magic_24_0.Y.t25 GNDA 0.098175f
C1864 two_stage_opamp_dummy_magic_24_0.Y.t41 GNDA 0.098175f
C1865 two_stage_opamp_dummy_magic_24_0.Y.t28 GNDA 0.098175f
C1866 two_stage_opamp_dummy_magic_24_0.Y.t44 GNDA 0.104563f
C1867 two_stage_opamp_dummy_magic_24_0.Y.n70 GNDA 0.082862f
C1868 two_stage_opamp_dummy_magic_24_0.Y.n71 GNDA 0.046856f
C1869 two_stage_opamp_dummy_magic_24_0.Y.n72 GNDA 0.046856f
C1870 two_stage_opamp_dummy_magic_24_0.Y.n73 GNDA 0.042115f
C1871 two_stage_opamp_dummy_magic_24_0.Y.t54 GNDA 0.098175f
C1872 two_stage_opamp_dummy_magic_24_0.Y.t38 GNDA 0.098175f
C1873 two_stage_opamp_dummy_magic_24_0.Y.t51 GNDA 0.098175f
C1874 two_stage_opamp_dummy_magic_24_0.Y.t36 GNDA 0.098175f
C1875 two_stage_opamp_dummy_magic_24_0.Y.t52 GNDA 0.104563f
C1876 two_stage_opamp_dummy_magic_24_0.Y.n74 GNDA 0.082862f
C1877 two_stage_opamp_dummy_magic_24_0.Y.n75 GNDA 0.046856f
C1878 two_stage_opamp_dummy_magic_24_0.Y.n76 GNDA 0.046856f
C1879 two_stage_opamp_dummy_magic_24_0.Y.n77 GNDA 0.042115f
C1880 two_stage_opamp_dummy_magic_24_0.Y.n78 GNDA 0.010113f
C1881 two_stage_opamp_dummy_magic_24_0.Y.n79 GNDA 0.023958f
C1882 two_stage_opamp_dummy_magic_24_0.Y.n80 GNDA 0.056395f
C1883 two_stage_opamp_dummy_magic_24_0.Y.n81 GNDA 0.032165f
C1884 two_stage_opamp_dummy_magic_24_0.Y.n82 GNDA 0.036504f
C1885 two_stage_opamp_dummy_magic_24_0.Y.n83 GNDA 1.16471f
C1886 two_stage_opamp_dummy_magic_24_0.Y.n84 GNDA 0.070729f
C1887 two_stage_opamp_dummy_magic_24_0.Y.n85 GNDA 0.0714f
C1888 two_stage_opamp_dummy_magic_24_0.Y.n86 GNDA 0.096373f
C1889 two_stage_opamp_dummy_magic_24_0.Y.n87 GNDA 0.116025f
C1890 two_stage_opamp_dummy_magic_24_0.Y.n88 GNDA 0.0714f
C1891 two_stage_opamp_dummy_magic_24_0.Y.n89 GNDA 0.092019f
C1892 two_stage_opamp_dummy_magic_24_0.Y.n90 GNDA 0.0714f
C1893 two_stage_opamp_dummy_magic_24_0.Y.n91 GNDA 0.0714f
C1894 two_stage_opamp_dummy_magic_24_0.Y.n92 GNDA 0.092019f
C1895 two_stage_opamp_dummy_magic_24_0.Y.n93 GNDA 0.0714f
C1896 two_stage_opamp_dummy_magic_24_0.Y.n94 GNDA 0.117651f
C1897 two_stage_opamp_dummy_magic_24_0.Y.t0 GNDA 0.052062f
C1898 two_stage_opamp_dummy_magic_24_0.Y.t3 GNDA 0.052062f
C1899 two_stage_opamp_dummy_magic_24_0.Y.n95 GNDA 0.106499f
C1900 two_stage_opamp_dummy_magic_24_0.Y.n96 GNDA 0.284972f
C1901 two_stage_opamp_dummy_magic_24_0.Y.t24 GNDA 0.052062f
C1902 two_stage_opamp_dummy_magic_24_0.Y.t8 GNDA 0.052062f
C1903 two_stage_opamp_dummy_magic_24_0.Y.n97 GNDA 0.106499f
C1904 two_stage_opamp_dummy_magic_24_0.Y.n98 GNDA 0.289681f
C1905 two_stage_opamp_dummy_magic_24_0.Y.n99 GNDA 0.096333f
C1906 two_stage_opamp_dummy_magic_24_0.Y.t5 GNDA 0.052062f
C1907 two_stage_opamp_dummy_magic_24_0.Y.t6 GNDA 0.052062f
C1908 two_stage_opamp_dummy_magic_24_0.Y.n100 GNDA 0.106499f
C1909 two_stage_opamp_dummy_magic_24_0.Y.n101 GNDA 0.284972f
C1910 two_stage_opamp_dummy_magic_24_0.Y.n102 GNDA 0.056471f
C1911 two_stage_opamp_dummy_magic_24_0.Y.t7 GNDA 0.052062f
C1912 two_stage_opamp_dummy_magic_24_0.Y.t9 GNDA 0.052062f
C1913 two_stage_opamp_dummy_magic_24_0.Y.n103 GNDA 0.106499f
C1914 two_stage_opamp_dummy_magic_24_0.Y.n104 GNDA 0.284972f
C1915 two_stage_opamp_dummy_magic_24_0.Y.n105 GNDA 0.056471f
C1916 two_stage_opamp_dummy_magic_24_0.Y.t2 GNDA 0.052062f
C1917 two_stage_opamp_dummy_magic_24_0.Y.t23 GNDA 0.052062f
C1918 two_stage_opamp_dummy_magic_24_0.Y.n106 GNDA 0.106499f
C1919 two_stage_opamp_dummy_magic_24_0.Y.n107 GNDA 0.289681f
C1920 two_stage_opamp_dummy_magic_24_0.Y.n108 GNDA 0.096333f
C1921 two_stage_opamp_dummy_magic_24_0.Y.t1 GNDA 0.052062f
C1922 two_stage_opamp_dummy_magic_24_0.Y.t4 GNDA 0.052062f
C1923 two_stage_opamp_dummy_magic_24_0.Y.n109 GNDA 0.106499f
C1924 two_stage_opamp_dummy_magic_24_0.Y.n110 GNDA 0.284972f
C1925 two_stage_opamp_dummy_magic_24_0.Y.n111 GNDA 0.092019f
C1926 two_stage_opamp_dummy_magic_24_0.Y.n112 GNDA 0.078946f
C1927 two_stage_opamp_dummy_magic_24_0.Y.n113 GNDA 0.0476f
C1928 two_stage_opamp_dummy_magic_24_0.Y.n114 GNDA 0.0476f
C1929 two_stage_opamp_dummy_magic_24_0.Y.n115 GNDA 0.078946f
C1930 two_stage_opamp_dummy_magic_24_0.Y.n116 GNDA 0.092019f
C1931 two_stage_opamp_dummy_magic_24_0.Y.n117 GNDA 0.162793f
C1932 two_stage_opamp_dummy_magic_24_0.Y.n118 GNDA 0.241134f
C1933 two_stage_opamp_dummy_magic_24_0.Y.n119 GNDA 0.306644f
C1934 two_stage_opamp_dummy_magic_24_0.Y.n120 GNDA 0.0714f
C1935 two_stage_opamp_dummy_magic_24_0.Y.n121 GNDA 0.0714f
C1936 two_stage_opamp_dummy_magic_24_0.Y.n122 GNDA 0.116025f
C1937 two_stage_opamp_dummy_magic_24_0.Y.n123 GNDA 0.0714f
C1938 two_stage_opamp_dummy_magic_24_0.Y.n124 GNDA 0.0714f
C1939 two_stage_opamp_dummy_magic_24_0.Y.n125 GNDA 0.0714f
C1940 two_stage_opamp_dummy_magic_24_0.Y.n126 GNDA 0.0714f
C1941 two_stage_opamp_dummy_magic_24_0.Y.n127 GNDA 0.116025f
C1942 two_stage_opamp_dummy_magic_24_0.Y.n128 GNDA 0.0714f
C1943 two_stage_opamp_dummy_magic_24_0.Y.n129 GNDA 0.0714f
C1944 two_stage_opamp_dummy_magic_24_0.Y.n130 GNDA 0.0714f
C1945 two_stage_opamp_dummy_magic_24_0.Y.n131 GNDA 0.0714f
C1946 two_stage_opamp_dummy_magic_24_0.Y.n132 GNDA 0.0714f
C1947 two_stage_opamp_dummy_magic_24_0.Y.n133 GNDA 0.0714f
C1948 two_stage_opamp_dummy_magic_24_0.Y.n134 GNDA 0.0714f
C1949 two_stage_opamp_dummy_magic_24_0.Y.n135 GNDA 0.116025f
C1950 two_stage_opamp_dummy_magic_24_0.Y.n136 GNDA 0.379312f
C1951 two_stage_opamp_dummy_magic_24_0.Y.n137 GNDA 0.379312f
C1952 two_stage_opamp_dummy_magic_24_0.Y.n138 GNDA 0.0714f
C1953 two_stage_opamp_dummy_magic_24_0.Y.n140 GNDA 0.0714f
C1954 two_stage_opamp_dummy_magic_24_0.Y.n141 GNDA 0.0714f
C1955 two_stage_opamp_dummy_magic_24_0.Y.n143 GNDA 0.798786f
C1956 two_stage_opamp_dummy_magic_24_0.Y.n144 GNDA 0.798786f
C1957 two_stage_opamp_dummy_magic_24_0.Y.n146 GNDA 0.437324f
C1958 two_stage_opamp_dummy_magic_24_0.Y.n147 GNDA 1.80233f
C1959 two_stage_opamp_dummy_magic_24_0.Y.n148 GNDA 0.397162f
C1960 two_stage_opamp_dummy_magic_24_0.Y.n149 GNDA 0.410549f
C1961 two_stage_opamp_dummy_magic_24_0.Y.n150 GNDA 0.163625f
C1962 two_stage_opamp_dummy_magic_24_0.Y.n151 GNDA 0.098175f
C1963 two_stage_opamp_dummy_magic_24_0.Y.n152 GNDA 0.177012f
C1964 two_stage_opamp_dummy_magic_24_0.Y.n153 GNDA 0.098175f
C1965 two_stage_opamp_dummy_magic_24_0.Y.n154 GNDA 0.098175f
C1966 two_stage_opamp_dummy_magic_24_0.Y.n155 GNDA 0.098175f
C1967 two_stage_opamp_dummy_magic_24_0.Y.n156 GNDA 0.145775f
C1968 two_stage_opamp_dummy_magic_24_0.Vb2.t4 GNDA 0.019226f
C1969 two_stage_opamp_dummy_magic_24_0.Vb2.t2 GNDA 0.06729f
C1970 two_stage_opamp_dummy_magic_24_0.Vb2.t0 GNDA 0.06729f
C1971 two_stage_opamp_dummy_magic_24_0.Vb2.n0 GNDA 0.142896f
C1972 two_stage_opamp_dummy_magic_24_0.Vb2.t1 GNDA 0.125612f
C1973 two_stage_opamp_dummy_magic_24_0.Vb2.n1 GNDA 0.581662f
C1974 two_stage_opamp_dummy_magic_24_0.Vb2.t28 GNDA 0.075436f
C1975 two_stage_opamp_dummy_magic_24_0.Vb2.n2 GNDA 0.2896f
C1976 two_stage_opamp_dummy_magic_24_0.Vb2.t32 GNDA 0.095168f
C1977 two_stage_opamp_dummy_magic_24_0.Vb2.t26 GNDA 0.095168f
C1978 two_stage_opamp_dummy_magic_24_0.Vb2.t30 GNDA 0.095168f
C1979 two_stage_opamp_dummy_magic_24_0.Vb2.t24 GNDA 0.095168f
C1980 two_stage_opamp_dummy_magic_24_0.Vb2.t19 GNDA 0.109823f
C1981 two_stage_opamp_dummy_magic_24_0.Vb2.n3 GNDA 0.089164f
C1982 two_stage_opamp_dummy_magic_24_0.Vb2.n4 GNDA 0.054793f
C1983 two_stage_opamp_dummy_magic_24_0.Vb2.n5 GNDA 0.054793f
C1984 two_stage_opamp_dummy_magic_24_0.Vb2.n6 GNDA 0.048043f
C1985 two_stage_opamp_dummy_magic_24_0.Vb2.t14 GNDA 0.095168f
C1986 two_stage_opamp_dummy_magic_24_0.Vb2.t17 GNDA 0.095168f
C1987 two_stage_opamp_dummy_magic_24_0.Vb2.t20 GNDA 0.095168f
C1988 two_stage_opamp_dummy_magic_24_0.Vb2.t18 GNDA 0.095168f
C1989 two_stage_opamp_dummy_magic_24_0.Vb2.t22 GNDA 0.109823f
C1990 two_stage_opamp_dummy_magic_24_0.Vb2.n7 GNDA 0.089164f
C1991 two_stage_opamp_dummy_magic_24_0.Vb2.n8 GNDA 0.054793f
C1992 two_stage_opamp_dummy_magic_24_0.Vb2.n9 GNDA 0.054793f
C1993 two_stage_opamp_dummy_magic_24_0.Vb2.n10 GNDA 0.048043f
C1994 two_stage_opamp_dummy_magic_24_0.Vb2.n11 GNDA 0.035607f
C1995 two_stage_opamp_dummy_magic_24_0.Vb2.t13 GNDA 0.095168f
C1996 two_stage_opamp_dummy_magic_24_0.Vb2.t11 GNDA 0.095168f
C1997 two_stage_opamp_dummy_magic_24_0.Vb2.t29 GNDA 0.095168f
C1998 two_stage_opamp_dummy_magic_24_0.Vb2.t23 GNDA 0.095168f
C1999 two_stage_opamp_dummy_magic_24_0.Vb2.t27 GNDA 0.109823f
C2000 two_stage_opamp_dummy_magic_24_0.Vb2.n12 GNDA 0.089164f
C2001 two_stage_opamp_dummy_magic_24_0.Vb2.n13 GNDA 0.054793f
C2002 two_stage_opamp_dummy_magic_24_0.Vb2.n14 GNDA 0.054793f
C2003 two_stage_opamp_dummy_magic_24_0.Vb2.n15 GNDA 0.048043f
C2004 two_stage_opamp_dummy_magic_24_0.Vb2.t16 GNDA 0.095168f
C2005 two_stage_opamp_dummy_magic_24_0.Vb2.t21 GNDA 0.095168f
C2006 two_stage_opamp_dummy_magic_24_0.Vb2.t25 GNDA 0.095168f
C2007 two_stage_opamp_dummy_magic_24_0.Vb2.t31 GNDA 0.095168f
C2008 two_stage_opamp_dummy_magic_24_0.Vb2.t12 GNDA 0.109823f
C2009 two_stage_opamp_dummy_magic_24_0.Vb2.n16 GNDA 0.089164f
C2010 two_stage_opamp_dummy_magic_24_0.Vb2.n17 GNDA 0.054793f
C2011 two_stage_opamp_dummy_magic_24_0.Vb2.n18 GNDA 0.054793f
C2012 two_stage_opamp_dummy_magic_24_0.Vb2.n19 GNDA 0.048043f
C2013 two_stage_opamp_dummy_magic_24_0.Vb2.n20 GNDA 0.035084f
C2014 two_stage_opamp_dummy_magic_24_0.Vb2.n21 GNDA 0.794556f
C2015 two_stage_opamp_dummy_magic_24_0.Vb2.n22 GNDA 0.386457f
C2016 two_stage_opamp_dummy_magic_24_0.Vb2.t15 GNDA 0.123675f
C2017 two_stage_opamp_dummy_magic_24_0.Vb2.n23 GNDA 2.28086f
C2018 two_stage_opamp_dummy_magic_24_0.Vb2.t8 GNDA 0.019226f
C2019 two_stage_opamp_dummy_magic_24_0.Vb2.t3 GNDA 0.019226f
C2020 two_stage_opamp_dummy_magic_24_0.Vb2.n24 GNDA 0.064461f
C2021 two_stage_opamp_dummy_magic_24_0.Vb2.t6 GNDA 0.019226f
C2022 two_stage_opamp_dummy_magic_24_0.Vb2.t9 GNDA 0.019226f
C2023 two_stage_opamp_dummy_magic_24_0.Vb2.n25 GNDA 0.062693f
C2024 two_stage_opamp_dummy_magic_24_0.Vb2.n26 GNDA 0.572663f
C2025 two_stage_opamp_dummy_magic_24_0.Vb2.t7 GNDA 0.019226f
C2026 two_stage_opamp_dummy_magic_24_0.Vb2.t5 GNDA 0.019226f
C2027 two_stage_opamp_dummy_magic_24_0.Vb2.n27 GNDA 0.062693f
C2028 two_stage_opamp_dummy_magic_24_0.Vb2.n28 GNDA 0.375654f
C2029 two_stage_opamp_dummy_magic_24_0.Vb2.n29 GNDA 2.49016f
C2030 two_stage_opamp_dummy_magic_24_0.Vb2.n30 GNDA 0.062693f
C2031 two_stage_opamp_dummy_magic_24_0.Vb2.t10 GNDA 0.019226f
C2032 bgr_11_0.NFET_GATE_10uA.n0 GNDA 1.04726f
C2033 bgr_11_0.NFET_GATE_10uA.t1 GNDA 0.011025f
C2034 bgr_11_0.NFET_GATE_10uA.t0 GNDA 0.011025f
C2035 bgr_11_0.NFET_GATE_10uA.n1 GNDA 0.061322f
C2036 bgr_11_0.NFET_GATE_10uA.t21 GNDA 0.010749f
C2037 bgr_11_0.NFET_GATE_10uA.t15 GNDA 0.01589f
C2038 bgr_11_0.NFET_GATE_10uA.n2 GNDA 0.017509f
C2039 bgr_11_0.NFET_GATE_10uA.t12 GNDA 0.010749f
C2040 bgr_11_0.NFET_GATE_10uA.t18 GNDA 0.010749f
C2041 bgr_11_0.NFET_GATE_10uA.t6 GNDA 0.010749f
C2042 bgr_11_0.NFET_GATE_10uA.t13 GNDA 0.01589f
C2043 bgr_11_0.NFET_GATE_10uA.n3 GNDA 0.019665f
C2044 bgr_11_0.NFET_GATE_10uA.n4 GNDA 0.014057f
C2045 bgr_11_0.NFET_GATE_10uA.n5 GNDA 0.011901f
C2046 bgr_11_0.NFET_GATE_10uA.n6 GNDA 0.019415f
C2047 bgr_11_0.NFET_GATE_10uA.t20 GNDA 0.010749f
C2048 bgr_11_0.NFET_GATE_10uA.t14 GNDA 0.01589f
C2049 bgr_11_0.NFET_GATE_10uA.n7 GNDA 0.017509f
C2050 bgr_11_0.NFET_GATE_10uA.t9 GNDA 0.010749f
C2051 bgr_11_0.NFET_GATE_10uA.t17 GNDA 0.01589f
C2052 bgr_11_0.NFET_GATE_10uA.n8 GNDA 0.017509f
C2053 bgr_11_0.NFET_GATE_10uA.n9 GNDA 0.017128f
C2054 bgr_11_0.NFET_GATE_10uA.n10 GNDA 0.316054f
C2055 bgr_11_0.NFET_GATE_10uA.t16 GNDA 0.010749f
C2056 bgr_11_0.NFET_GATE_10uA.t10 GNDA 0.010749f
C2057 bgr_11_0.NFET_GATE_10uA.t11 GNDA 0.010749f
C2058 bgr_11_0.NFET_GATE_10uA.t5 GNDA 0.01589f
C2059 bgr_11_0.NFET_GATE_10uA.n11 GNDA 0.019665f
C2060 bgr_11_0.NFET_GATE_10uA.n12 GNDA 0.014057f
C2061 bgr_11_0.NFET_GATE_10uA.n13 GNDA 0.011901f
C2062 bgr_11_0.NFET_GATE_10uA.t22 GNDA 0.010749f
C2063 bgr_11_0.NFET_GATE_10uA.t8 GNDA 0.01589f
C2064 bgr_11_0.NFET_GATE_10uA.n14 GNDA 0.017509f
C2065 bgr_11_0.NFET_GATE_10uA.n15 GNDA 0.017128f
C2066 bgr_11_0.NFET_GATE_10uA.n16 GNDA 0.196104f
C2067 bgr_11_0.NFET_GATE_10uA.t19 GNDA 0.010749f
C2068 bgr_11_0.NFET_GATE_10uA.t3 GNDA 0.01589f
C2069 bgr_11_0.NFET_GATE_10uA.n17 GNDA 0.017509f
C2070 bgr_11_0.NFET_GATE_10uA.t7 GNDA 0.01269f
C2071 bgr_11_0.NFET_GATE_10uA.n18 GNDA 0.023781f
C2072 bgr_11_0.NFET_GATE_10uA.t4 GNDA 0.011025f
C2073 bgr_11_0.NFET_GATE_10uA.n19 GNDA 0.03676f
C2074 bgr_11_0.NFET_GATE_10uA.t2 GNDA 0.011025f
C2075 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t13 GNDA 0.436158f
C2076 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t18 GNDA 0.437612f
C2077 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 GNDA 0.23505f
C2078 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 GNDA 0.250988f
C2079 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t47 GNDA 0.436158f
C2080 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 GNDA 0.437612f
C2081 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 GNDA 0.23505f
C2082 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 GNDA 0.274473f
C2083 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t30 GNDA 0.436158f
C2084 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 GNDA 0.437612f
C2085 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 GNDA 0.23505f
C2086 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 GNDA 0.274473f
C2087 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t71 GNDA 0.436158f
C2088 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 GNDA 0.437612f
C2089 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 GNDA 0.23505f
C2090 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 GNDA 0.274473f
C2091 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t105 GNDA 0.436158f
C2092 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 GNDA 0.437612f
C2093 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 GNDA 0.23505f
C2094 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 GNDA 0.274473f
C2095 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t1 GNDA 0.436158f
C2096 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 GNDA 0.437612f
C2097 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 GNDA 0.461098f
C2098 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 GNDA 0.23505f
C2099 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 GNDA 0.274473f
C2100 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 GNDA 0.436158f
C2101 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 GNDA 0.437612f
C2102 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 GNDA 0.461098f
C2103 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 GNDA 0.23505f
C2104 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 GNDA 0.274473f
C2105 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 GNDA 0.437612f
C2106 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 GNDA 0.439198f
C2107 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t44 GNDA 0.437612f
C2108 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 GNDA 0.441043f
C2109 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 GNDA 0.479698f
C2110 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t64 GNDA 0.437612f
C2111 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 GNDA 0.439198f
C2112 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 GNDA 0.437612f
C2113 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 GNDA 0.439198f
C2114 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 GNDA 0.437612f
C2115 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 GNDA 0.439198f
C2116 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 GNDA 0.437612f
C2117 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 GNDA 0.439198f
C2118 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 GNDA 0.437612f
C2119 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 GNDA 0.439198f
C2120 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t124 GNDA 0.437612f
C2121 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 GNDA 0.439198f
C2122 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 GNDA 0.437612f
C2123 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 GNDA 0.439198f
C2124 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 GNDA 0.437612f
C2125 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 GNDA 0.439198f
C2126 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 GNDA 0.437612f
C2127 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 GNDA 0.439198f
C2128 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t129 GNDA 0.437612f
C2129 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 GNDA 0.439198f
C2130 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 GNDA 0.437612f
C2131 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 GNDA 0.439198f
C2132 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 GNDA 0.437612f
C2133 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 GNDA 0.439198f
C2134 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 GNDA 0.437612f
C2135 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 GNDA 0.439198f
C2136 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 GNDA 0.437612f
C2137 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 GNDA 0.439198f
C2138 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 GNDA 0.437612f
C2139 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 GNDA 0.439198f
C2140 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t33 GNDA 0.437612f
C2141 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 GNDA 0.439198f
C2142 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 GNDA 0.437612f
C2143 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 GNDA 0.439198f
C2144 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 GNDA 0.437612f
C2145 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 GNDA 0.439198f
C2146 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 GNDA 0.437612f
C2147 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 GNDA 0.439198f
C2148 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t111 GNDA 0.437612f
C2149 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 GNDA 0.439198f
C2150 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 GNDA 0.437612f
C2151 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 GNDA 0.439198f
C2152 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 GNDA 0.437612f
C2153 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 GNDA 0.439198f
C2154 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 GNDA 0.437612f
C2155 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 GNDA 0.439198f
C2156 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 GNDA 0.437612f
C2157 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 GNDA 0.439198f
C2158 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 GNDA 0.437612f
C2159 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 GNDA 0.439198f
C2160 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t14 GNDA 0.437612f
C2161 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 GNDA 0.439198f
C2162 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t11 GNDA 0.437612f
C2163 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 GNDA 0.439198f
C2164 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 GNDA 0.437612f
C2165 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 GNDA 0.439198f
C2166 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 GNDA 0.437612f
C2167 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 GNDA 0.439198f
C2168 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t51 GNDA 0.437612f
C2169 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 GNDA 0.439198f
C2170 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t65 GNDA 0.437612f
C2171 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 GNDA 0.459069f
C2172 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 GNDA 0.437612f
C2173 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 GNDA 0.23505f
C2174 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 GNDA 0.251562f
C2175 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 GNDA 0.437612f
C2176 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 GNDA 0.23505f
C2177 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 GNDA 0.249533f
C2178 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 GNDA 0.437612f
C2179 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 GNDA 0.23505f
C2180 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 GNDA 0.249533f
C2181 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 GNDA 0.437612f
C2182 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 GNDA 0.23505f
C2183 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 GNDA 0.249533f
C2184 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t117 GNDA 0.437612f
C2185 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 GNDA 0.23505f
C2186 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 GNDA 0.249533f
C2187 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t24 GNDA 0.437612f
C2188 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 GNDA 0.23505f
C2189 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 GNDA 0.249533f
C2190 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t58 GNDA 0.437612f
C2191 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 GNDA 0.23505f
C2192 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 GNDA 0.249533f
C2193 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 GNDA 0.437612f
C2194 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 GNDA 0.23505f
C2195 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 GNDA 0.249533f
C2196 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t3 GNDA 0.437612f
C2197 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 GNDA 0.23505f
C2198 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 GNDA 0.249533f
C2199 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t31 GNDA 0.437612f
C2200 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 GNDA 0.439198f
C2201 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 GNDA 0.437612f
C2202 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 GNDA 0.439198f
C2203 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 GNDA 0.211565f
C2204 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 GNDA 0.272887f
C2205 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 GNDA 0.233596f
C2206 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 GNDA 0.296373f
C2207 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 GNDA 0.233596f
C2208 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 GNDA 0.318272f
C2209 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 GNDA 0.233596f
C2210 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 GNDA 0.318272f
C2211 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 GNDA 0.233596f
C2212 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 GNDA 0.318272f
C2213 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 GNDA 0.233596f
C2214 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 GNDA 0.318272f
C2215 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 GNDA 0.233596f
C2216 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 GNDA 0.318272f
C2217 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 GNDA 0.233596f
C2218 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 GNDA 0.318272f
C2219 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 GNDA 0.233596f
C2220 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 GNDA 0.318272f
C2221 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 GNDA 0.233596f
C2222 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 GNDA 0.318272f
C2223 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 GNDA 0.233596f
C2224 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 GNDA 0.318272f
C2225 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 GNDA 0.233596f
C2226 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 GNDA 0.318272f
C2227 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 GNDA 0.233596f
C2228 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 GNDA 0.318272f
C2229 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 GNDA 0.233596f
C2230 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 GNDA 0.318272f
C2231 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 GNDA 0.233596f
C2232 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 GNDA 0.318272f
C2233 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 GNDA 0.233596f
C2234 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 GNDA 0.318272f
C2235 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 GNDA 0.233596f
C2236 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 GNDA 0.318272f
C2237 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 GNDA 0.233596f
C2238 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 GNDA 0.296373f
C2239 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t36 GNDA 0.436158f
C2240 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 GNDA 0.211565f
C2241 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 GNDA 0.274473f
C2242 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 GNDA 0.436158f
C2243 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t100 GNDA 0.211565f
C2244 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 GNDA 0.274473f
C2245 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t19 GNDA 0.436158f
C2246 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n36 GNDA 0.274473f
C2247 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 GNDA 0.23505f
C2248 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 GNDA 0.461098f
C2249 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 GNDA 0.623087f
C2250 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 GNDA 0.37036f
C2251 VOUT+.n0 GNDA 0.037514f
C2252 VOUT+.t16 GNDA 0.054708f
C2253 VOUT+.t14 GNDA 0.054708f
C2254 VOUT+.n1 GNDA 0.117546f
C2255 VOUT+.n2 GNDA 0.282696f
C2256 VOUT+.n3 GNDA 0.037514f
C2257 VOUT+.n4 GNDA 0.242255f
C2258 VOUT+.t15 GNDA 0.054708f
C2259 VOUT+.t4 GNDA 0.054708f
C2260 VOUT+.n5 GNDA 0.117546f
C2261 VOUT+.n6 GNDA 0.29257f
C2262 VOUT+.n7 GNDA 0.167231f
C2263 VOUT+.t17 GNDA 0.054708f
C2264 VOUT+.t18 GNDA 0.054708f
C2265 VOUT+.n8 GNDA 0.117546f
C2266 VOUT+.n9 GNDA 0.277939f
C2267 VOUT+.n10 GNDA 0.127554f
C2268 VOUT+.n11 GNDA 0.037514f
C2269 VOUT+.n12 GNDA 0.193575f
C2270 VOUT+.n13 GNDA 0.037514f
C2271 VOUT+.n14 GNDA 0.037514f
C2272 VOUT+.n15 GNDA 0.037514f
C2273 VOUT+.n16 GNDA 0.037514f
C2274 VOUT+.n17 GNDA 0.080303f
C2275 VOUT+.n18 GNDA 0.145366f
C2276 VOUT+.t2 GNDA 0.089232f
C2277 VOUT+.n19 GNDA 0.310134f
C2278 VOUT+.n20 GNDA 0.078154f
C2279 VOUT+.n23 GNDA 0.039859f
C2280 VOUT+.n25 GNDA 0.039859f
C2281 VOUT+.n28 GNDA 0.058615f
C2282 VOUT+.n29 GNDA 0.097692f
C2283 VOUT+.n30 GNDA 0.062101f
C2284 VOUT+.n31 GNDA 0.058615f
C2285 VOUT+.n33 GNDA 0.039859f
C2286 VOUT+.n34 GNDA 0.037162f
C2287 VOUT+.n35 GNDA 0.039859f
C2288 VOUT+.n36 GNDA 0.051582f
C2289 VOUT+.n37 GNDA 0.07442f
C2290 VOUT+.n38 GNDA 0.072423f
C2291 VOUT+.n39 GNDA 0.051582f
C2292 VOUT+.n40 GNDA 0.051582f
C2293 VOUT+.n41 GNDA 0.072423f
C2294 VOUT+.n42 GNDA 0.072423f
C2295 VOUT+.n43 GNDA 0.051582f
C2296 VOUT+.n44 GNDA 0.082578f
C2297 VOUT+.t13 GNDA 0.046892f
C2298 VOUT+.t3 GNDA 0.046892f
C2299 VOUT+.n45 GNDA 0.096082f
C2300 VOUT+.n46 GNDA 0.248017f
C2301 VOUT+.t0 GNDA 0.046892f
C2302 VOUT+.t12 GNDA 0.046892f
C2303 VOUT+.n47 GNDA 0.096082f
C2304 VOUT+.n48 GNDA 0.248017f
C2305 VOUT+.t5 GNDA 0.046892f
C2306 VOUT+.t7 GNDA 0.046892f
C2307 VOUT+.n49 GNDA 0.096082f
C2308 VOUT+.n50 GNDA 0.245517f
C2309 VOUT+.n51 GNDA 0.059628f
C2310 VOUT+.t11 GNDA 0.046892f
C2311 VOUT+.t9 GNDA 0.046892f
C2312 VOUT+.n52 GNDA 0.096082f
C2313 VOUT+.n53 GNDA 0.245517f
C2314 VOUT+.n54 GNDA 0.033799f
C2315 VOUT+.t10 GNDA 0.046892f
C2316 VOUT+.t8 GNDA 0.046892f
C2317 VOUT+.n55 GNDA 0.096082f
C2318 VOUT+.n56 GNDA 0.245517f
C2319 VOUT+.n57 GNDA 0.033799f
C2320 VOUT+.n58 GNDA 0.059628f
C2321 VOUT+.t6 GNDA 0.046892f
C2322 VOUT+.t1 GNDA 0.046892f
C2323 VOUT+.n59 GNDA 0.096082f
C2324 VOUT+.n60 GNDA 0.245517f
C2325 VOUT+.n61 GNDA 0.039424f
C2326 VOUT+.n62 GNDA 0.023446f
C2327 VOUT+.n63 GNDA 0.023446f
C2328 VOUT+.n64 GNDA 0.039424f
C2329 VOUT+.n65 GNDA 0.072423f
C2330 VOUT+.n66 GNDA 0.101377f
C2331 VOUT+.n67 GNDA 0.12632f
C2332 VOUT+.n68 GNDA 0.176797f
C2333 VOUT+.n69 GNDA 0.051582f
C2334 VOUT+.n70 GNDA 0.084406f
C2335 VOUT+.n71 GNDA 0.051582f
C2336 VOUT+.n72 GNDA 0.084406f
C2337 VOUT+.n73 GNDA 0.051582f
C2338 VOUT+.n74 GNDA 0.051582f
C2339 VOUT+.n75 GNDA 0.051582f
C2340 VOUT+.n76 GNDA 0.084406f
C2341 VOUT+.n77 GNDA 0.051582f
C2342 VOUT+.n78 GNDA 0.077372f
C2343 VOUT+.n79 GNDA 0.250874f
C2344 VOUT+.n81 GNDA 0.078154f
C2345 VOUT+.n82 GNDA 0.039859f
C2346 VOUT+.n84 GNDA 0.039859f
C2347 VOUT+.n87 GNDA 0.078154f
C2348 VOUT+.n88 GNDA 0.24384f
C2349 VOUT+.n89 GNDA 0.664308f
C2350 VOUT+.n92 GNDA 0.058615f
C2351 VOUT+.n93 GNDA 0.058615f
C2352 VOUT+.n94 GNDA 0.058615f
C2353 VOUT+.n95 GNDA 0.058615f
C2354 VOUT+.n96 GNDA 0.171928f
C2355 VOUT+.n97 GNDA 0.058615f
C2356 VOUT+.t118 GNDA 0.312615f
C2357 VOUT+.t90 GNDA 0.31794f
C2358 VOUT+.t89 GNDA 0.312615f
C2359 VOUT+.n98 GNDA 0.209598f
C2360 VOUT+.n99 GNDA 0.136769f
C2361 VOUT+.t154 GNDA 0.317273f
C2362 VOUT+.t61 GNDA 0.317273f
C2363 VOUT+.t99 GNDA 0.317273f
C2364 VOUT+.t133 GNDA 0.317273f
C2365 VOUT+.t40 GNDA 0.317273f
C2366 VOUT+.t72 GNDA 0.317273f
C2367 VOUT+.t116 GNDA 0.317273f
C2368 VOUT+.t149 GNDA 0.317273f
C2369 VOUT+.t56 GNDA 0.317273f
C2370 VOUT+.t92 GNDA 0.317273f
C2371 VOUT+.t128 GNDA 0.312615f
C2372 VOUT+.n100 GNDA 0.210265f
C2373 VOUT+.t91 GNDA 0.312615f
C2374 VOUT+.n101 GNDA 0.268881f
C2375 VOUT+.t39 GNDA 0.312615f
C2376 VOUT+.n102 GNDA 0.268881f
C2377 VOUT+.t148 GNDA 0.312615f
C2378 VOUT+.n103 GNDA 0.268881f
C2379 VOUT+.t115 GNDA 0.312615f
C2380 VOUT+.n104 GNDA 0.268881f
C2381 VOUT+.t71 GNDA 0.312615f
C2382 VOUT+.n105 GNDA 0.268881f
C2383 VOUT+.t25 GNDA 0.312615f
C2384 VOUT+.n106 GNDA 0.268881f
C2385 VOUT+.t132 GNDA 0.312615f
C2386 VOUT+.n107 GNDA 0.268881f
C2387 VOUT+.t98 GNDA 0.312615f
C2388 VOUT+.n108 GNDA 0.268881f
C2389 VOUT+.t44 GNDA 0.312615f
C2390 VOUT+.n109 GNDA 0.268881f
C2391 VOUT+.t153 GNDA 0.312615f
C2392 VOUT+.t126 GNDA 0.31794f
C2393 VOUT+.t125 GNDA 0.312615f
C2394 VOUT+.n110 GNDA 0.209598f
C2395 VOUT+.n111 GNDA 0.254f
C2396 VOUT+.t75 GNDA 0.31794f
C2397 VOUT+.t35 GNDA 0.312615f
C2398 VOUT+.n112 GNDA 0.209598f
C2399 VOUT+.t87 GNDA 0.312615f
C2400 VOUT+.t106 GNDA 0.31794f
C2401 VOUT+.t53 GNDA 0.312615f
C2402 VOUT+.n113 GNDA 0.209598f
C2403 VOUT+.n114 GNDA 0.254f
C2404 VOUT+.t146 GNDA 0.31794f
C2405 VOUT+.t95 GNDA 0.312615f
C2406 VOUT+.n115 GNDA 0.209598f
C2407 VOUT+.t58 GNDA 0.312615f
C2408 VOUT+.t32 GNDA 0.31794f
C2409 VOUT+.t29 GNDA 0.312615f
C2410 VOUT+.n116 GNDA 0.209598f
C2411 VOUT+.n117 GNDA 0.254f
C2412 VOUT+.t114 GNDA 0.31794f
C2413 VOUT+.t60 GNDA 0.312615f
C2414 VOUT+.n118 GNDA 0.209598f
C2415 VOUT+.t21 GNDA 0.312615f
C2416 VOUT+.t143 GNDA 0.31794f
C2417 VOUT+.t141 GNDA 0.312615f
C2418 VOUT+.n119 GNDA 0.209598f
C2419 VOUT+.n120 GNDA 0.254f
C2420 VOUT+.t152 GNDA 0.31794f
C2421 VOUT+.t103 GNDA 0.312615f
C2422 VOUT+.n121 GNDA 0.209598f
C2423 VOUT+.t62 GNDA 0.312615f
C2424 VOUT+.t38 GNDA 0.31794f
C2425 VOUT+.t36 GNDA 0.312615f
C2426 VOUT+.n122 GNDA 0.209598f
C2427 VOUT+.n123 GNDA 0.254f
C2428 VOUT+.t80 GNDA 0.312615f
C2429 VOUT+.t113 GNDA 0.31794f
C2430 VOUT+.t73 GNDA 0.312615f
C2431 VOUT+.n124 GNDA 0.209598f
C2432 VOUT+.n125 GNDA 0.136769f
C2433 VOUT+.t121 GNDA 0.317273f
C2434 VOUT+.t101 GNDA 0.317273f
C2435 VOUT+.t78 GNDA 0.31794f
C2436 VOUT+.t134 GNDA 0.312615f
C2437 VOUT+.n126 GNDA 0.204714f
C2438 VOUT+.t138 GNDA 0.317273f
C2439 VOUT+.t119 GNDA 0.31794f
C2440 VOUT+.t26 GNDA 0.312615f
C2441 VOUT+.n127 GNDA 0.204714f
C2442 VOUT+.t31 GNDA 0.317273f
C2443 VOUT+.t24 GNDA 0.31794f
C2444 VOUT+.t150 GNDA 0.312615f
C2445 VOUT+.n128 GNDA 0.204714f
C2446 VOUT+.t156 GNDA 0.317273f
C2447 VOUT+.t47 GNDA 0.317273f
C2448 VOUT+.t52 GNDA 0.317273f
C2449 VOUT+.t81 GNDA 0.317535f
C2450 VOUT+.t86 GNDA 0.317273f
C2451 VOUT+.t122 GNDA 0.317535f
C2452 VOUT+.t127 GNDA 0.317273f
C2453 VOUT+.t104 GNDA 0.317535f
C2454 VOUT+.t110 GNDA 0.317273f
C2455 VOUT+.t139 GNDA 0.317535f
C2456 VOUT+.t144 GNDA 0.317273f
C2457 VOUT+.t107 GNDA 0.312615f
C2458 VOUT+.n129 GNDA 0.346022f
C2459 VOUT+.t63 GNDA 0.312615f
C2460 VOUT+.n130 GNDA 0.404638f
C2461 VOUT+.t85 GNDA 0.312615f
C2462 VOUT+.n131 GNDA 0.404638f
C2463 VOUT+.t48 GNDA 0.312615f
C2464 VOUT+.n132 GNDA 0.404638f
C2465 VOUT+.t155 GNDA 0.312615f
C2466 VOUT+.n133 GNDA 0.400992f
C2467 VOUT+.t117 GNDA 0.312615f
C2468 VOUT+.n134 GNDA 0.332381f
C2469 VOUT+.t136 GNDA 0.312615f
C2470 VOUT+.n135 GNDA 0.332381f
C2471 VOUT+.t100 GNDA 0.312615f
C2472 VOUT+.n136 GNDA 0.332381f
C2473 VOUT+.t57 GNDA 0.312615f
C2474 VOUT+.n137 GNDA 0.268881f
C2475 VOUT+.t79 GNDA 0.312615f
C2476 VOUT+.n138 GNDA 0.268881f
C2477 VOUT+.t41 GNDA 0.312615f
C2478 VOUT+.t67 GNDA 0.31794f
C2479 VOUT+.t34 GNDA 0.312615f
C2480 VOUT+.n139 GNDA 0.209598f
C2481 VOUT+.n140 GNDA 0.254f
C2482 VOUT+.t93 GNDA 0.31794f
C2483 VOUT+.t120 GNDA 0.312615f
C2484 VOUT+.n141 GNDA 0.209598f
C2485 VOUT+.t74 GNDA 0.312615f
C2486 VOUT+.t111 GNDA 0.31794f
C2487 VOUT+.t68 GNDA 0.312615f
C2488 VOUT+.n142 GNDA 0.209598f
C2489 VOUT+.n143 GNDA 0.254f
C2490 VOUT+.t45 GNDA 0.31794f
C2491 VOUT+.t135 GNDA 0.312615f
C2492 VOUT+.n144 GNDA 0.209598f
C2493 VOUT+.t102 GNDA 0.312615f
C2494 VOUT+.t70 GNDA 0.31794f
C2495 VOUT+.t69 GNDA 0.312615f
C2496 VOUT+.n145 GNDA 0.209598f
C2497 VOUT+.n146 GNDA 0.254f
C2498 VOUT+.t147 GNDA 0.31794f
C2499 VOUT+.t96 GNDA 0.312615f
C2500 VOUT+.n147 GNDA 0.209598f
C2501 VOUT+.t59 GNDA 0.312615f
C2502 VOUT+.t33 GNDA 0.31794f
C2503 VOUT+.t30 GNDA 0.312615f
C2504 VOUT+.n148 GNDA 0.209598f
C2505 VOUT+.n149 GNDA 0.254f
C2506 VOUT+.t37 GNDA 0.31794f
C2507 VOUT+.t129 GNDA 0.312615f
C2508 VOUT+.n150 GNDA 0.209598f
C2509 VOUT+.t94 GNDA 0.312615f
C2510 VOUT+.t66 GNDA 0.31794f
C2511 VOUT+.t65 GNDA 0.312615f
C2512 VOUT+.n151 GNDA 0.209598f
C2513 VOUT+.n152 GNDA 0.254f
C2514 VOUT+.t142 GNDA 0.31794f
C2515 VOUT+.t88 GNDA 0.312615f
C2516 VOUT+.n153 GNDA 0.209598f
C2517 VOUT+.t54 GNDA 0.312615f
C2518 VOUT+.t28 GNDA 0.31794f
C2519 VOUT+.t27 GNDA 0.312615f
C2520 VOUT+.n154 GNDA 0.209598f
C2521 VOUT+.n155 GNDA 0.254f
C2522 VOUT+.t105 GNDA 0.31794f
C2523 VOUT+.t50 GNDA 0.312615f
C2524 VOUT+.n156 GNDA 0.209598f
C2525 VOUT+.t19 GNDA 0.312615f
C2526 VOUT+.t131 GNDA 0.31794f
C2527 VOUT+.t130 GNDA 0.312615f
C2528 VOUT+.n157 GNDA 0.209598f
C2529 VOUT+.n158 GNDA 0.254f
C2530 VOUT+.t137 GNDA 0.31794f
C2531 VOUT+.t82 GNDA 0.312615f
C2532 VOUT+.n159 GNDA 0.209598f
C2533 VOUT+.t49 GNDA 0.312615f
C2534 VOUT+.t23 GNDA 0.31794f
C2535 VOUT+.t22 GNDA 0.312615f
C2536 VOUT+.n160 GNDA 0.209598f
C2537 VOUT+.n161 GNDA 0.254f
C2538 VOUT+.t97 GNDA 0.31794f
C2539 VOUT+.t42 GNDA 0.312615f
C2540 VOUT+.n162 GNDA 0.209598f
C2541 VOUT+.t151 GNDA 0.312615f
C2542 VOUT+.t124 GNDA 0.31794f
C2543 VOUT+.t123 GNDA 0.312615f
C2544 VOUT+.n163 GNDA 0.209598f
C2545 VOUT+.n164 GNDA 0.254f
C2546 VOUT+.t55 GNDA 0.31794f
C2547 VOUT+.t145 GNDA 0.312615f
C2548 VOUT+.n165 GNDA 0.209598f
C2549 VOUT+.t112 GNDA 0.312615f
C2550 VOUT+.t84 GNDA 0.31794f
C2551 VOUT+.t83 GNDA 0.312615f
C2552 VOUT+.n166 GNDA 0.209598f
C2553 VOUT+.n167 GNDA 0.254f
C2554 VOUT+.t20 GNDA 0.31794f
C2555 VOUT+.t109 GNDA 0.312615f
C2556 VOUT+.n168 GNDA 0.209598f
C2557 VOUT+.t64 GNDA 0.312615f
C2558 VOUT+.t46 GNDA 0.31794f
C2559 VOUT+.t43 GNDA 0.312615f
C2560 VOUT+.n169 GNDA 0.209598f
C2561 VOUT+.n170 GNDA 0.254f
C2562 VOUT+.t77 GNDA 0.31794f
C2563 VOUT+.t76 GNDA 0.312615f
C2564 VOUT+.n171 GNDA 0.209598f
C2565 VOUT+.t108 GNDA 0.312615f
C2566 VOUT+.n172 GNDA 0.254f
C2567 VOUT+.t140 GNDA 0.312615f
C2568 VOUT+.n173 GNDA 0.133838f
C2569 VOUT+.t51 GNDA 0.312615f
C2570 VOUT+.n174 GNDA 0.257908f
C2571 VOUT+.n175 GNDA 0.196362f
C2572 VOUT+.n176 GNDA 0.058615f
C2573 VOUT+.n177 GNDA 0.058615f
C2574 VOUT+.n179 GNDA 0.674077f
C2575 VOUT+.n180 GNDA 0.059048f
C2576 VOUT+.n181 GNDA 0.708269f
C2577 VOUT+.n182 GNDA 0.039859f
C2578 VOUT+.n184 GNDA 0.037514f
C2579 VOUT+.n185 GNDA 0.6985f
C2580 VOUT+.n187 GNDA 0.039859f
C2581 VOUT+.n188 GNDA 0.078154f
C2582 VOUT+.n189 GNDA 0.044548f
C2583 two_stage_opamp_dummy_magic_24_0.VD4.n0 GNDA 0.365754f
C2584 two_stage_opamp_dummy_magic_24_0.VD4.n1 GNDA 0.09179f
C2585 two_stage_opamp_dummy_magic_24_0.VD4.n2 GNDA 0.118729f
C2586 two_stage_opamp_dummy_magic_24_0.VD4.n3 GNDA 0.138157f
C2587 two_stage_opamp_dummy_magic_24_0.VD4.n4 GNDA 0.114974f
C2588 two_stage_opamp_dummy_magic_24_0.VD4.n5 GNDA 0.187808f
C2589 two_stage_opamp_dummy_magic_24_0.VD4.n6 GNDA 0.187325f
C2590 two_stage_opamp_dummy_magic_24_0.VD4.n7 GNDA 0.138157f
C2591 two_stage_opamp_dummy_magic_24_0.VD4.n8 GNDA 0.187808f
C2592 two_stage_opamp_dummy_magic_24_0.VD4.t22 GNDA 0.05037f
C2593 two_stage_opamp_dummy_magic_24_0.VD4.n9 GNDA 0.093202f
C2594 two_stage_opamp_dummy_magic_24_0.VD4.n10 GNDA 0.093202f
C2595 two_stage_opamp_dummy_magic_24_0.VD4.t25 GNDA 0.05037f
C2596 two_stage_opamp_dummy_magic_24_0.VD4.t28 GNDA 0.05037f
C2597 two_stage_opamp_dummy_magic_24_0.VD4.n11 GNDA 0.103037f
C2598 two_stage_opamp_dummy_magic_24_0.VD4.n12 GNDA 0.284144f
C2599 two_stage_opamp_dummy_magic_24_0.VD4.n13 GNDA 0.069079f
C2600 two_stage_opamp_dummy_magic_24_0.VD4.t32 GNDA 0.088322f
C2601 two_stage_opamp_dummy_magic_24_0.VD4.n14 GNDA 0.201305f
C2602 two_stage_opamp_dummy_magic_24_0.VD4.t5 GNDA 0.05037f
C2603 two_stage_opamp_dummy_magic_24_0.VD4.t15 GNDA 0.05037f
C2604 two_stage_opamp_dummy_magic_24_0.VD4.n15 GNDA 0.106864f
C2605 two_stage_opamp_dummy_magic_24_0.VD4.n16 GNDA 0.382443f
C2606 two_stage_opamp_dummy_magic_24_0.VD4.n17 GNDA 0.069079f
C2607 two_stage_opamp_dummy_magic_24_0.VD4.t3 GNDA 0.05037f
C2608 two_stage_opamp_dummy_magic_24_0.VD4.t17 GNDA 0.05037f
C2609 two_stage_opamp_dummy_magic_24_0.VD4.n18 GNDA 0.106864f
C2610 two_stage_opamp_dummy_magic_24_0.VD4.n19 GNDA 0.069079f
C2611 two_stage_opamp_dummy_magic_24_0.VD4.n20 GNDA 0.069079f
C2612 two_stage_opamp_dummy_magic_24_0.VD4.t1 GNDA 0.05037f
C2613 two_stage_opamp_dummy_magic_24_0.VD4.t9 GNDA 0.05037f
C2614 two_stage_opamp_dummy_magic_24_0.VD4.n21 GNDA 0.106864f
C2615 two_stage_opamp_dummy_magic_24_0.VD4.n22 GNDA 0.069079f
C2616 two_stage_opamp_dummy_magic_24_0.VD4.n23 GNDA 0.069079f
C2617 two_stage_opamp_dummy_magic_24_0.VD4.t13 GNDA 0.05037f
C2618 two_stage_opamp_dummy_magic_24_0.VD4.t11 GNDA 0.05037f
C2619 two_stage_opamp_dummy_magic_24_0.VD4.n24 GNDA 0.106864f
C2620 two_stage_opamp_dummy_magic_24_0.VD4.t7 GNDA 0.05037f
C2621 two_stage_opamp_dummy_magic_24_0.VD4.t19 GNDA 0.05037f
C2622 two_stage_opamp_dummy_magic_24_0.VD4.n25 GNDA 0.106864f
C2623 two_stage_opamp_dummy_magic_24_0.VD4.n26 GNDA 0.427691f
C2624 two_stage_opamp_dummy_magic_24_0.VD4.t35 GNDA 0.088322f
C2625 two_stage_opamp_dummy_magic_24_0.VD4.t34 GNDA 0.179173f
C2626 two_stage_opamp_dummy_magic_24_0.VD4.n27 GNDA 0.519765f
C2627 two_stage_opamp_dummy_magic_24_0.VD4.t33 GNDA 0.429348f
C2628 two_stage_opamp_dummy_magic_24_0.VD4.t14 GNDA 0.336759f
C2629 two_stage_opamp_dummy_magic_24_0.VD4.t4 GNDA 0.336759f
C2630 two_stage_opamp_dummy_magic_24_0.VD4.t16 GNDA 0.336759f
C2631 two_stage_opamp_dummy_magic_24_0.VD4.t2 GNDA 0.336759f
C2632 two_stage_opamp_dummy_magic_24_0.VD4.t8 GNDA 0.336759f
C2633 two_stage_opamp_dummy_magic_24_0.VD4.t0 GNDA 0.336759f
C2634 two_stage_opamp_dummy_magic_24_0.VD4.t10 GNDA 0.336759f
C2635 two_stage_opamp_dummy_magic_24_0.VD4.t12 GNDA 0.336759f
C2636 two_stage_opamp_dummy_magic_24_0.VD4.t18 GNDA 0.336759f
C2637 two_stage_opamp_dummy_magic_24_0.VD4.t6 GNDA 0.336759f
C2638 two_stage_opamp_dummy_magic_24_0.VD4.t36 GNDA 0.429348f
C2639 two_stage_opamp_dummy_magic_24_0.VD4.t37 GNDA 0.179173f
C2640 two_stage_opamp_dummy_magic_24_0.VD4.n28 GNDA 0.519765f
C2641 two_stage_opamp_dummy_magic_24_0.VD4.n29 GNDA 0.212445f
C2642 two_stage_opamp_dummy_magic_24_0.VD4.n30 GNDA 0.249218f
C2643 two_stage_opamp_dummy_magic_24_0.VD4.n31 GNDA 0.296675f
C2644 two_stage_opamp_dummy_magic_24_0.VD4.n32 GNDA 0.069079f
C2645 two_stage_opamp_dummy_magic_24_0.VD4.n33 GNDA 0.069079f
C2646 two_stage_opamp_dummy_magic_24_0.VD4.n34 GNDA 0.382443f
C2647 two_stage_opamp_dummy_magic_24_0.VD4.n35 GNDA 0.069079f
C2648 two_stage_opamp_dummy_magic_24_0.VD4.n36 GNDA 0.069079f
C2649 two_stage_opamp_dummy_magic_24_0.VD4.n37 GNDA 0.069079f
C2650 two_stage_opamp_dummy_magic_24_0.VD4.n38 GNDA 0.069079f
C2651 two_stage_opamp_dummy_magic_24_0.VD4.n39 GNDA 0.382443f
C2652 two_stage_opamp_dummy_magic_24_0.VD4.n40 GNDA 0.069079f
C2653 two_stage_opamp_dummy_magic_24_0.VD4.n41 GNDA 0.069079f
C2654 two_stage_opamp_dummy_magic_24_0.VD4.n42 GNDA 0.069079f
C2655 two_stage_opamp_dummy_magic_24_0.VD4.n43 GNDA 0.069079f
C2656 two_stage_opamp_dummy_magic_24_0.VD4.n44 GNDA 0.382443f
C2657 two_stage_opamp_dummy_magic_24_0.VD4.n45 GNDA 0.069079f
C2658 two_stage_opamp_dummy_magic_24_0.VD4.n46 GNDA 0.069079f
C2659 two_stage_opamp_dummy_magic_24_0.VD4.n47 GNDA 0.069079f
C2660 two_stage_opamp_dummy_magic_24_0.VD4.n48 GNDA 0.069079f
C2661 two_stage_opamp_dummy_magic_24_0.VD4.n49 GNDA 0.069079f
C2662 two_stage_opamp_dummy_magic_24_0.VD4.n50 GNDA 0.069079f
C2663 two_stage_opamp_dummy_magic_24_0.VD4.n51 GNDA 0.069079f
C2664 two_stage_opamp_dummy_magic_24_0.VD4.n52 GNDA 0.118729f
C2665 two_stage_opamp_dummy_magic_24_0.VD4.n53 GNDA 0.40152f
C2666 two_stage_opamp_dummy_magic_24_0.VD4.n54 GNDA 0.424704f
C2667 two_stage_opamp_dummy_magic_24_0.VD4.t20 GNDA 0.05037f
C2668 two_stage_opamp_dummy_magic_24_0.VD4.t27 GNDA 0.05037f
C2669 two_stage_opamp_dummy_magic_24_0.VD4.n55 GNDA 0.103037f
C2670 two_stage_opamp_dummy_magic_24_0.VD4.n56 GNDA 0.288699f
C2671 two_stage_opamp_dummy_magic_24_0.VD4.t30 GNDA 0.05037f
C2672 two_stage_opamp_dummy_magic_24_0.VD4.t21 GNDA 0.05037f
C2673 two_stage_opamp_dummy_magic_24_0.VD4.n57 GNDA 0.103037f
C2674 two_stage_opamp_dummy_magic_24_0.VD4.n58 GNDA 0.299839f
C2675 two_stage_opamp_dummy_magic_24_0.VD4.n59 GNDA 0.249218f
C2676 two_stage_opamp_dummy_magic_24_0.VD4.t26 GNDA 0.05037f
C2677 two_stage_opamp_dummy_magic_24_0.VD4.t29 GNDA 0.05037f
C2678 two_stage_opamp_dummy_magic_24_0.VD4.n60 GNDA 0.103037f
C2679 two_stage_opamp_dummy_magic_24_0.VD4.n61 GNDA 0.284144f
C2680 two_stage_opamp_dummy_magic_24_0.VD4.n62 GNDA 0.187161f
C2681 two_stage_opamp_dummy_magic_24_0.VD4.n63 GNDA 0.158068f
C2682 two_stage_opamp_dummy_magic_24_0.VD4.n64 GNDA 0.141913f
C2683 two_stage_opamp_dummy_magic_24_0.VD4.t24 GNDA 0.05037f
C2684 two_stage_opamp_dummy_magic_24_0.VD4.t23 GNDA 0.05037f
C2685 two_stage_opamp_dummy_magic_24_0.VD4.n65 GNDA 0.103037f
C2686 two_stage_opamp_dummy_magic_24_0.VD4.n66 GNDA 0.284144f
C2687 two_stage_opamp_dummy_magic_24_0.VD4.n67 GNDA 0.054635f
C2688 two_stage_opamp_dummy_magic_24_0.VD4.n68 GNDA 0.054635f
C2689 two_stage_opamp_dummy_magic_24_0.VD4.n69 GNDA 0.284144f
C2690 two_stage_opamp_dummy_magic_24_0.VD4.n70 GNDA 0.103037f
C2691 two_stage_opamp_dummy_magic_24_0.VD4.t31 GNDA 0.05037f
C2692 two_stage_opamp_dummy_magic_24_0.Vb3.t6 GNDA 0.011238f
C2693 two_stage_opamp_dummy_magic_24_0.Vb3.t3 GNDA 0.011238f
C2694 two_stage_opamp_dummy_magic_24_0.Vb3.n0 GNDA 0.036199f
C2695 two_stage_opamp_dummy_magic_24_0.Vb3.t0 GNDA 0.011238f
C2696 two_stage_opamp_dummy_magic_24_0.Vb3.t5 GNDA 0.011238f
C2697 two_stage_opamp_dummy_magic_24_0.Vb3.n1 GNDA 0.036199f
C2698 two_stage_opamp_dummy_magic_24_0.Vb3.n2 GNDA 0.199565f
C2699 two_stage_opamp_dummy_magic_24_0.Vb3.t1 GNDA 0.011238f
C2700 two_stage_opamp_dummy_magic_24_0.Vb3.t7 GNDA 0.011238f
C2701 two_stage_opamp_dummy_magic_24_0.Vb3.n3 GNDA 0.033944f
C2702 two_stage_opamp_dummy_magic_24_0.Vb3.n4 GNDA 0.639061f
C2703 two_stage_opamp_dummy_magic_24_0.Vb3.t2 GNDA 0.039333f
C2704 two_stage_opamp_dummy_magic_24_0.Vb3.t4 GNDA 0.039333f
C2705 two_stage_opamp_dummy_magic_24_0.Vb3.n5 GNDA 0.108511f
C2706 two_stage_opamp_dummy_magic_24_0.Vb3.t11 GNDA 0.055629f
C2707 two_stage_opamp_dummy_magic_24_0.Vb3.t9 GNDA 0.055629f
C2708 two_stage_opamp_dummy_magic_24_0.Vb3.t27 GNDA 0.055629f
C2709 two_stage_opamp_dummy_magic_24_0.Vb3.t22 GNDA 0.055629f
C2710 two_stage_opamp_dummy_magic_24_0.Vb3.t17 GNDA 0.064195f
C2711 two_stage_opamp_dummy_magic_24_0.Vb3.n6 GNDA 0.05212f
C2712 two_stage_opamp_dummy_magic_24_0.Vb3.n7 GNDA 0.032029f
C2713 two_stage_opamp_dummy_magic_24_0.Vb3.n8 GNDA 0.032029f
C2714 two_stage_opamp_dummy_magic_24_0.Vb3.n9 GNDA 0.028083f
C2715 two_stage_opamp_dummy_magic_24_0.Vb3.t13 GNDA 0.055629f
C2716 two_stage_opamp_dummy_magic_24_0.Vb3.t19 GNDA 0.055629f
C2717 two_stage_opamp_dummy_magic_24_0.Vb3.t24 GNDA 0.055629f
C2718 two_stage_opamp_dummy_magic_24_0.Vb3.t28 GNDA 0.055629f
C2719 two_stage_opamp_dummy_magic_24_0.Vb3.t26 GNDA 0.064195f
C2720 two_stage_opamp_dummy_magic_24_0.Vb3.n10 GNDA 0.05212f
C2721 two_stage_opamp_dummy_magic_24_0.Vb3.n11 GNDA 0.032029f
C2722 two_stage_opamp_dummy_magic_24_0.Vb3.n12 GNDA 0.032029f
C2723 two_stage_opamp_dummy_magic_24_0.Vb3.n13 GNDA 0.028083f
C2724 two_stage_opamp_dummy_magic_24_0.Vb3.n14 GNDA 0.028342f
C2725 two_stage_opamp_dummy_magic_24_0.Vb3.t21 GNDA 0.055629f
C2726 two_stage_opamp_dummy_magic_24_0.Vb3.t23 GNDA 0.055629f
C2727 two_stage_opamp_dummy_magic_24_0.Vb3.t18 GNDA 0.055629f
C2728 two_stage_opamp_dummy_magic_24_0.Vb3.t12 GNDA 0.055629f
C2729 two_stage_opamp_dummy_magic_24_0.Vb3.t10 GNDA 0.064195f
C2730 two_stage_opamp_dummy_magic_24_0.Vb3.n15 GNDA 0.05212f
C2731 two_stage_opamp_dummy_magic_24_0.Vb3.n16 GNDA 0.032029f
C2732 two_stage_opamp_dummy_magic_24_0.Vb3.n17 GNDA 0.032029f
C2733 two_stage_opamp_dummy_magic_24_0.Vb3.n18 GNDA 0.028083f
C2734 two_stage_opamp_dummy_magic_24_0.Vb3.t25 GNDA 0.055629f
C2735 two_stage_opamp_dummy_magic_24_0.Vb3.t8 GNDA 0.055629f
C2736 two_stage_opamp_dummy_magic_24_0.Vb3.t14 GNDA 0.055629f
C2737 two_stage_opamp_dummy_magic_24_0.Vb3.t20 GNDA 0.055629f
C2738 two_stage_opamp_dummy_magic_24_0.Vb3.t16 GNDA 0.064195f
C2739 two_stage_opamp_dummy_magic_24_0.Vb3.n19 GNDA 0.05212f
C2740 two_stage_opamp_dummy_magic_24_0.Vb3.n20 GNDA 0.032029f
C2741 two_stage_opamp_dummy_magic_24_0.Vb3.n21 GNDA 0.032029f
C2742 two_stage_opamp_dummy_magic_24_0.Vb3.n22 GNDA 0.028083f
C2743 two_stage_opamp_dummy_magic_24_0.Vb3.n23 GNDA 0.028889f
C2744 two_stage_opamp_dummy_magic_24_0.Vb3.n24 GNDA 0.966028f
C2745 two_stage_opamp_dummy_magic_24_0.Vb3.t15 GNDA 0.072669f
C2746 two_stage_opamp_dummy_magic_24_0.Vb3.n25 GNDA 0.272086f
C2747 two_stage_opamp_dummy_magic_24_0.Vb3.n26 GNDA 1.13609f
C2748 bgr_11_0.VB3_CUR_BIAS GNDA 1.77244f
C2749 two_stage_opamp_dummy_magic_24_0.Vb1.t28 GNDA 0.045649f
C2750 two_stage_opamp_dummy_magic_24_0.Vb1.t34 GNDA 0.04781f
C2751 two_stage_opamp_dummy_magic_24_0.Vb1.t189 GNDA 0.04781f
C2752 two_stage_opamp_dummy_magic_24_0.Vb1.t129 GNDA 0.04781f
C2753 two_stage_opamp_dummy_magic_24_0.Vb1.t181 GNDA 0.04781f
C2754 two_stage_opamp_dummy_magic_24_0.Vb1.t121 GNDA 0.04781f
C2755 two_stage_opamp_dummy_magic_24_0.Vb1.t59 GNDA 0.04781f
C2756 two_stage_opamp_dummy_magic_24_0.Vb1.t110 GNDA 0.04781f
C2757 two_stage_opamp_dummy_magic_24_0.Vb1.t51 GNDA 0.04781f
C2758 two_stage_opamp_dummy_magic_24_0.Vb1.t205 GNDA 0.04781f
C2759 two_stage_opamp_dummy_magic_24_0.Vb1.t45 GNDA 0.04781f
C2760 two_stage_opamp_dummy_magic_24_0.Vb1.t197 GNDA 0.04781f
C2761 two_stage_opamp_dummy_magic_24_0.Vb1.t136 GNDA 0.04781f
C2762 two_stage_opamp_dummy_magic_24_0.Vb1.t75 GNDA 0.04781f
C2763 two_stage_opamp_dummy_magic_24_0.Vb1.t130 GNDA 0.04781f
C2764 two_stage_opamp_dummy_magic_24_0.Vb1.t76 GNDA 0.04781f
C2765 two_stage_opamp_dummy_magic_24_0.Vb1.t14 GNDA 0.04781f
C2766 two_stage_opamp_dummy_magic_24_0.Vb1.t69 GNDA 0.04781f
C2767 two_stage_opamp_dummy_magic_24_0.Vb1.t9 GNDA 0.04781f
C2768 two_stage_opamp_dummy_magic_24_0.Vb1.t162 GNDA 0.04781f
C2769 two_stage_opamp_dummy_magic_24_0.Vb1.t214 GNDA 0.04781f
C2770 two_stage_opamp_dummy_magic_24_0.Vb1.t150 GNDA 0.04781f
C2771 two_stage_opamp_dummy_magic_24_0.Vb1.t91 GNDA 0.04781f
C2772 two_stage_opamp_dummy_magic_24_0.Vb1.t152 GNDA 0.037912f
C2773 two_stage_opamp_dummy_magic_24_0.Vb1.t210 GNDA 0.039946f
C2774 two_stage_opamp_dummy_magic_24_0.Vb1.t174 GNDA 0.039946f
C2775 two_stage_opamp_dummy_magic_24_0.Vb1.t16 GNDA 0.038049f
C2776 two_stage_opamp_dummy_magic_24_0.Vb1.t161 GNDA 0.037912f
C2777 two_stage_opamp_dummy_magic_24_0.Vb1.t5 GNDA 0.039946f
C2778 two_stage_opamp_dummy_magic_24_0.Vb1.t62 GNDA 0.039946f
C2779 two_stage_opamp_dummy_magic_24_0.Vb1.t25 GNDA 0.038049f
C2780 two_stage_opamp_dummy_magic_24_0.Vb1.t100 GNDA 0.037912f
C2781 two_stage_opamp_dummy_magic_24_0.Vb1.t160 GNDA 0.039946f
C2782 two_stage_opamp_dummy_magic_24_0.Vb1.t125 GNDA 0.039946f
C2783 two_stage_opamp_dummy_magic_24_0.Vb1.t177 GNDA 0.038049f
C2784 two_stage_opamp_dummy_magic_24_0.Vb1.t98 GNDA 0.037912f
C2785 two_stage_opamp_dummy_magic_24_0.Vb1.t157 GNDA 0.039946f
C2786 two_stage_opamp_dummy_magic_24_0.Vb1.t216 GNDA 0.039946f
C2787 two_stage_opamp_dummy_magic_24_0.Vb1.t179 GNDA 0.038049f
C2788 two_stage_opamp_dummy_magic_24_0.Vb1.t39 GNDA 0.037912f
C2789 two_stage_opamp_dummy_magic_24_0.Vb1.t97 GNDA 0.039946f
C2790 two_stage_opamp_dummy_magic_24_0.Vb1.t65 GNDA 0.039946f
C2791 two_stage_opamp_dummy_magic_24_0.Vb1.t116 GNDA 0.038049f
C2792 two_stage_opamp_dummy_magic_24_0.Vb1.t37 GNDA 0.037912f
C2793 two_stage_opamp_dummy_magic_24_0.Vb1.t94 GNDA 0.039946f
C2794 two_stage_opamp_dummy_magic_24_0.Vb1.t153 GNDA 0.039946f
C2795 two_stage_opamp_dummy_magic_24_0.Vb1.t118 GNDA 0.038049f
C2796 two_stage_opamp_dummy_magic_24_0.Vb1.t192 GNDA 0.037912f
C2797 two_stage_opamp_dummy_magic_24_0.Vb1.t35 GNDA 0.039946f
C2798 two_stage_opamp_dummy_magic_24_0.Vb1.t3 GNDA 0.039946f
C2799 two_stage_opamp_dummy_magic_24_0.Vb1.t56 GNDA 0.038049f
C2800 two_stage_opamp_dummy_magic_24_0.Vb1.t90 GNDA 0.037912f
C2801 two_stage_opamp_dummy_magic_24_0.Vb1.t147 GNDA 0.039946f
C2802 two_stage_opamp_dummy_magic_24_0.Vb1.t207 GNDA 0.039946f
C2803 two_stage_opamp_dummy_magic_24_0.Vb1.t171 GNDA 0.038049f
C2804 two_stage_opamp_dummy_magic_24_0.Vb1.t29 GNDA 0.037912f
C2805 two_stage_opamp_dummy_magic_24_0.Vb1.t89 GNDA 0.039946f
C2806 two_stage_opamp_dummy_magic_24_0.Vb1.t54 GNDA 0.039946f
C2807 two_stage_opamp_dummy_magic_24_0.Vb1.t108 GNDA 0.038049f
C2808 two_stage_opamp_dummy_magic_24_0.Vb1.t27 GNDA 0.037912f
C2809 two_stage_opamp_dummy_magic_24_0.Vb1.t86 GNDA 0.039946f
C2810 two_stage_opamp_dummy_magic_24_0.Vb1.t145 GNDA 0.039946f
C2811 two_stage_opamp_dummy_magic_24_0.Vb1.t109 GNDA 0.038049f
C2812 two_stage_opamp_dummy_magic_24_0.Vb1.t184 GNDA 0.037912f
C2813 two_stage_opamp_dummy_magic_24_0.Vb1.t26 GNDA 0.039946f
C2814 two_stage_opamp_dummy_magic_24_0.Vb1.t208 GNDA 0.039946f
C2815 two_stage_opamp_dummy_magic_24_0.Vb1.t49 GNDA 0.038049f
C2816 two_stage_opamp_dummy_magic_24_0.Vb1.t183 GNDA 0.037912f
C2817 two_stage_opamp_dummy_magic_24_0.Vb1.t24 GNDA 0.039946f
C2818 two_stage_opamp_dummy_magic_24_0.Vb1.t84 GNDA 0.039946f
C2819 two_stage_opamp_dummy_magic_24_0.Vb1.t50 GNDA 0.038049f
C2820 two_stage_opamp_dummy_magic_24_0.Vb1.t124 GNDA 0.037912f
C2821 two_stage_opamp_dummy_magic_24_0.Vb1.t182 GNDA 0.039946f
C2822 two_stage_opamp_dummy_magic_24_0.Vb1.t146 GNDA 0.039946f
C2823 two_stage_opamp_dummy_magic_24_0.Vb1.t204 GNDA 0.038049f
C2824 two_stage_opamp_dummy_magic_24_0.Vb1.t21 GNDA 0.037912f
C2825 two_stage_opamp_dummy_magic_24_0.Vb1.t80 GNDA 0.039946f
C2826 two_stage_opamp_dummy_magic_24_0.Vb1.t138 GNDA 0.039946f
C2827 two_stage_opamp_dummy_magic_24_0.Vb1.t104 GNDA 0.038049f
C2828 two_stage_opamp_dummy_magic_24_0.Vb1.t175 GNDA 0.037912f
C2829 two_stage_opamp_dummy_magic_24_0.Vb1.t19 GNDA 0.039946f
C2830 two_stage_opamp_dummy_magic_24_0.Vb1.t203 GNDA 0.039946f
C2831 two_stage_opamp_dummy_magic_24_0.Vb1.t41 GNDA 0.038049f
C2832 two_stage_opamp_dummy_magic_24_0.Vb1.t173 GNDA 0.037912f
C2833 two_stage_opamp_dummy_magic_24_0.Vb1.t17 GNDA 0.039946f
C2834 two_stage_opamp_dummy_magic_24_0.Vb1.t77 GNDA 0.039946f
C2835 two_stage_opamp_dummy_magic_24_0.Vb1.t43 GNDA 0.038049f
C2836 two_stage_opamp_dummy_magic_24_0.Vb1.t114 GNDA 0.037912f
C2837 two_stage_opamp_dummy_magic_24_0.Vb1.t172 GNDA 0.039946f
C2838 two_stage_opamp_dummy_magic_24_0.Vb1.t142 GNDA 0.039946f
C2839 two_stage_opamp_dummy_magic_24_0.Vb1.t194 GNDA 0.038049f
C2840 two_stage_opamp_dummy_magic_24_0.Vb1.t113 GNDA 0.037912f
C2841 two_stage_opamp_dummy_magic_24_0.Vb1.t169 GNDA 0.039946f
C2842 two_stage_opamp_dummy_magic_24_0.Vb1.t15 GNDA 0.039946f
C2843 two_stage_opamp_dummy_magic_24_0.Vb1.t195 GNDA 0.038049f
C2844 two_stage_opamp_dummy_magic_24_0.Vb1.t52 GNDA 0.037912f
C2845 two_stage_opamp_dummy_magic_24_0.Vb1.t111 GNDA 0.039946f
C2846 two_stage_opamp_dummy_magic_24_0.Vb1.t79 GNDA 0.039946f
C2847 two_stage_opamp_dummy_magic_24_0.Vb1.t135 GNDA 0.038049f
C2848 two_stage_opamp_dummy_magic_24_0.Vb1.t168 GNDA 0.037912f
C2849 two_stage_opamp_dummy_magic_24_0.Vb1.t13 GNDA 0.039946f
C2850 two_stage_opamp_dummy_magic_24_0.Vb1.t71 GNDA 0.039946f
C2851 two_stage_opamp_dummy_magic_24_0.Vb1.t33 GNDA 0.038049f
C2852 two_stage_opamp_dummy_magic_24_0.Vb1.t107 GNDA 0.037912f
C2853 two_stage_opamp_dummy_magic_24_0.Vb1.t167 GNDA 0.039946f
C2854 two_stage_opamp_dummy_magic_24_0.Vb1.t133 GNDA 0.039946f
C2855 two_stage_opamp_dummy_magic_24_0.Vb1.t186 GNDA 0.038049f
C2856 two_stage_opamp_dummy_magic_24_0.Vb1.t106 GNDA 0.037912f
C2857 two_stage_opamp_dummy_magic_24_0.Vb1.t166 GNDA 0.039946f
C2858 two_stage_opamp_dummy_magic_24_0.Vb1.t10 GNDA 0.039946f
C2859 two_stage_opamp_dummy_magic_24_0.Vb1.t188 GNDA 0.038049f
C2860 two_stage_opamp_dummy_magic_24_0.Vb1.t48 GNDA 0.037912f
C2861 two_stage_opamp_dummy_magic_24_0.Vb1.t105 GNDA 0.039946f
C2862 two_stage_opamp_dummy_magic_24_0.Vb1.t73 GNDA 0.039946f
C2863 two_stage_opamp_dummy_magic_24_0.Vb1.t126 GNDA 0.038049f
C2864 two_stage_opamp_dummy_magic_24_0.Vb1.t47 GNDA 0.037912f
C2865 two_stage_opamp_dummy_magic_24_0.Vb1.t103 GNDA 0.039946f
C2866 two_stage_opamp_dummy_magic_24_0.Vb1.t163 GNDA 0.039946f
C2867 two_stage_opamp_dummy_magic_24_0.Vb1.t128 GNDA 0.038049f
C2868 two_stage_opamp_dummy_magic_24_0.Vb1.t202 GNDA 0.037912f
C2869 two_stage_opamp_dummy_magic_24_0.Vb1.t46 GNDA 0.039946f
C2870 two_stage_opamp_dummy_magic_24_0.Vb1.t11 GNDA 0.039946f
C2871 two_stage_opamp_dummy_magic_24_0.Vb1.t66 GNDA 0.038049f
C2872 two_stage_opamp_dummy_magic_24_0.Vb1.t200 GNDA 0.037912f
C2873 two_stage_opamp_dummy_magic_24_0.Vb1.t42 GNDA 0.039946f
C2874 two_stage_opamp_dummy_magic_24_0.Vb1.t99 GNDA 0.039946f
C2875 two_stage_opamp_dummy_magic_24_0.Vb1.t67 GNDA 0.038049f
C2876 two_stage_opamp_dummy_magic_24_0.Vb1.t140 GNDA 0.037912f
C2877 two_stage_opamp_dummy_magic_24_0.Vb1.t198 GNDA 0.039946f
C2878 two_stage_opamp_dummy_magic_24_0.Vb1.t164 GNDA 0.039946f
C2879 two_stage_opamp_dummy_magic_24_0.Vb1.t6 GNDA 0.038049f
C2880 two_stage_opamp_dummy_magic_24_0.Vb1.t38 GNDA 0.037912f
C2881 two_stage_opamp_dummy_magic_24_0.Vb1.t95 GNDA 0.039946f
C2882 two_stage_opamp_dummy_magic_24_0.Vb1.t154 GNDA 0.039946f
C2883 two_stage_opamp_dummy_magic_24_0.Vb1.t119 GNDA 0.038049f
C2884 two_stage_opamp_dummy_magic_24_0.Vb1.t193 GNDA 0.037912f
C2885 two_stage_opamp_dummy_magic_24_0.Vb1.t36 GNDA 0.039946f
C2886 two_stage_opamp_dummy_magic_24_0.Vb1.t4 GNDA 0.039946f
C2887 two_stage_opamp_dummy_magic_24_0.Vb1.t57 GNDA 0.038049f
C2888 two_stage_opamp_dummy_magic_24_0.Vb1.t201 GNDA 0.037912f
C2889 two_stage_opamp_dummy_magic_24_0.Vb1.t44 GNDA 0.039946f
C2890 two_stage_opamp_dummy_magic_24_0.Vb1.t101 GNDA 0.039946f
C2891 two_stage_opamp_dummy_magic_24_0.Vb1.t68 GNDA 0.038049f
C2892 two_stage_opamp_dummy_magic_24_0.Vb1.t141 GNDA 0.037912f
C2893 two_stage_opamp_dummy_magic_24_0.Vb1.t199 GNDA 0.039946f
C2894 two_stage_opamp_dummy_magic_24_0.Vb1.t165 GNDA 0.039946f
C2895 two_stage_opamp_dummy_magic_24_0.Vb1.t7 GNDA 0.038049f
C2896 two_stage_opamp_dummy_magic_24_0.Vb1.t139 GNDA 0.037912f
C2897 two_stage_opamp_dummy_magic_24_0.Vb1.t196 GNDA 0.039946f
C2898 two_stage_opamp_dummy_magic_24_0.Vb1.t40 GNDA 0.039946f
C2899 two_stage_opamp_dummy_magic_24_0.Vb1.t8 GNDA 0.038049f
C2900 two_stage_opamp_dummy_magic_24_0.Vb1.t78 GNDA 0.037912f
C2901 two_stage_opamp_dummy_magic_24_0.Vb1.t137 GNDA 0.039946f
C2902 two_stage_opamp_dummy_magic_24_0.Vb1.t102 GNDA 0.039946f
C2903 two_stage_opamp_dummy_magic_24_0.Vb1.t159 GNDA 0.038049f
C2904 two_stage_opamp_dummy_magic_24_0.Vb1.t191 GNDA 0.037912f
C2905 two_stage_opamp_dummy_magic_24_0.Vb1.t32 GNDA 0.039946f
C2906 two_stage_opamp_dummy_magic_24_0.Vb1.t92 GNDA 0.039946f
C2907 two_stage_opamp_dummy_magic_24_0.Vb1.t60 GNDA 0.038049f
C2908 two_stage_opamp_dummy_magic_24_0.Vb1.t134 GNDA 0.037912f
C2909 two_stage_opamp_dummy_magic_24_0.Vb1.t190 GNDA 0.039946f
C2910 two_stage_opamp_dummy_magic_24_0.Vb1.t158 GNDA 0.039946f
C2911 two_stage_opamp_dummy_magic_24_0.Vb1.t209 GNDA 0.038049f
C2912 two_stage_opamp_dummy_magic_24_0.Vb1.t132 GNDA 0.037912f
C2913 two_stage_opamp_dummy_magic_24_0.Vb1.t187 GNDA 0.039946f
C2914 two_stage_opamp_dummy_magic_24_0.Vb1.t30 GNDA 0.039946f
C2915 two_stage_opamp_dummy_magic_24_0.Vb1.t213 GNDA 0.038049f
C2916 two_stage_opamp_dummy_magic_24_0.Vb1.t74 GNDA 0.037912f
C2917 two_stage_opamp_dummy_magic_24_0.Vb1.t131 GNDA 0.039946f
C2918 two_stage_opamp_dummy_magic_24_0.Vb1.t96 GNDA 0.039946f
C2919 two_stage_opamp_dummy_magic_24_0.Vb1.t148 GNDA 0.038049f
C2920 two_stage_opamp_dummy_magic_24_0.Vb1.t72 GNDA 0.037912f
C2921 two_stage_opamp_dummy_magic_24_0.Vb1.t127 GNDA 0.039946f
C2922 two_stage_opamp_dummy_magic_24_0.Vb1.t185 GNDA 0.039946f
C2923 two_stage_opamp_dummy_magic_24_0.Vb1.t149 GNDA 0.038049f
C2924 two_stage_opamp_dummy_magic_24_0.Vb1.t12 GNDA 0.037912f
C2925 two_stage_opamp_dummy_magic_24_0.Vb1.t70 GNDA 0.039946f
C2926 two_stage_opamp_dummy_magic_24_0.Vb1.t31 GNDA 0.039946f
C2927 two_stage_opamp_dummy_magic_24_0.Vb1.t87 GNDA 0.038049f
C2928 two_stage_opamp_dummy_magic_24_0.Vb1.t123 GNDA 0.037912f
C2929 two_stage_opamp_dummy_magic_24_0.Vb1.t180 GNDA 0.039946f
C2930 two_stage_opamp_dummy_magic_24_0.Vb1.t22 GNDA 0.039946f
C2931 two_stage_opamp_dummy_magic_24_0.Vb1.t206 GNDA 0.038049f
C2932 two_stage_opamp_dummy_magic_24_0.Vb1.t64 GNDA 0.037912f
C2933 two_stage_opamp_dummy_magic_24_0.Vb1.t122 GNDA 0.039946f
C2934 two_stage_opamp_dummy_magic_24_0.Vb1.t85 GNDA 0.039946f
C2935 two_stage_opamp_dummy_magic_24_0.Vb1.t143 GNDA 0.038049f
C2936 two_stage_opamp_dummy_magic_24_0.Vb1.t63 GNDA 0.037912f
C2937 two_stage_opamp_dummy_magic_24_0.Vb1.t120 GNDA 0.039946f
C2938 two_stage_opamp_dummy_magic_24_0.Vb1.t176 GNDA 0.039946f
C2939 two_stage_opamp_dummy_magic_24_0.Vb1.t144 GNDA 0.038049f
C2940 two_stage_opamp_dummy_magic_24_0.Vb1.t2 GNDA 0.037912f
C2941 two_stage_opamp_dummy_magic_24_0.Vb1.t61 GNDA 0.039946f
C2942 two_stage_opamp_dummy_magic_24_0.Vb1.t23 GNDA 0.039946f
C2943 two_stage_opamp_dummy_magic_24_0.Vb1.t82 GNDA 0.038049f
C2944 two_stage_opamp_dummy_magic_24_0.Vb1.t156 GNDA 0.037912f
C2945 two_stage_opamp_dummy_magic_24_0.Vb1.t215 GNDA 0.039946f
C2946 two_stage_opamp_dummy_magic_24_0.Vb1.t178 GNDA 0.039946f
C2947 two_stage_opamp_dummy_magic_24_0.Vb1.t18 GNDA 0.038049f
C2948 two_stage_opamp_dummy_magic_24_0.Vb1.t155 GNDA 0.037912f
C2949 two_stage_opamp_dummy_magic_24_0.Vb1.t211 GNDA 0.039946f
C2950 two_stage_opamp_dummy_magic_24_0.Vb1.t53 GNDA 0.039946f
C2951 two_stage_opamp_dummy_magic_24_0.Vb1.t20 GNDA 0.038049f
C2952 two_stage_opamp_dummy_magic_24_0.Vb1.t93 GNDA 0.037912f
C2953 two_stage_opamp_dummy_magic_24_0.Vb1.t151 GNDA 0.039946f
C2954 two_stage_opamp_dummy_magic_24_0.Vb1.t117 GNDA 0.039946f
C2955 two_stage_opamp_dummy_magic_24_0.Vb1.t170 GNDA 0.038049f
C2956 two_stage_opamp_dummy_magic_24_0.Vb1.n1 GNDA -0.109581f
C2957 two_stage_opamp_dummy_magic_24_0.Vb1.t217 GNDA 0.147492f
C2958 two_stage_opamp_dummy_magic_24_0.Vb1.t58 GNDA 0.039946f
C2959 two_stage_opamp_dummy_magic_24_0.Vb1.t115 GNDA 0.039946f
C2960 two_stage_opamp_dummy_magic_24_0.Vb1.t83 GNDA 0.038049f
C2961 two_stage_opamp_dummy_magic_24_0.Vb1.t88 GNDA 0.045901f
C2962 two_stage_opamp_dummy_magic_24_0.Vb1.t81 GNDA 0.038049f
C2963 two_stage_opamp_dummy_magic_24_0.Vb1.t112 GNDA 0.039946f
C2964 two_stage_opamp_dummy_magic_24_0.Vb1.t55 GNDA 0.039946f
C2965 two_stage_opamp_dummy_magic_24_0.Vb1.t212 GNDA 0.060601f
C2966 two_stage_opamp_dummy_magic_24_0.Vb1.n2 GNDA 0.037338f
C2967 two_stage_opamp_dummy_magic_24_0.Vb1.t241 GNDA 0.031784f
C2968 two_stage_opamp_dummy_magic_24_0.Vb1.n16 GNDA 0.017627f
C2969 two_stage_opamp_dummy_magic_24_0.Vb1.n36 GNDA 0.082195f
C2970 bgr_11_0.VB1_CUR_BIAS GNDA 0.056727f
C2971 VDDA.n15 GNDA 0.498447f
C2972 VDDA.n16 GNDA 0.45208f
C2973 VDDA.n17 GNDA 1.62285f
C2974 VDDA.n44 GNDA 0.012171f
C2975 VDDA.n48 GNDA 0.011737f
C2976 VDDA.n52 GNDA 0.010867f
C2977 VDDA.n56 GNDA 0.012171f
C2978 VDDA.n60 GNDA 0.011737f
C2979 VDDA.n64 GNDA 0.010867f
C2980 VDDA.n68 GNDA 0.012171f
C2981 VDDA.n72 GNDA 0.011737f
C2982 VDDA.n76 GNDA 0.010867f
C2983 VDDA.n80 GNDA 0.012171f
C2984 VDDA.n84 GNDA 0.011737f
C2985 VDDA.n91 GNDA 0.033905f
C2986 VDDA.n92 GNDA 0.012171f
C2987 VDDA.n98 GNDA 0.010867f
C2988 VDDA.n99 GNDA 0.010867f
C2989 VDDA.n100 GNDA 0.011737f
C2990 VDDA.n106 GNDA 0.012171f
C2991 VDDA.n107 GNDA 0.011737f
C2992 VDDA.n108 GNDA 0.010867f
C2993 VDDA.n114 GNDA 0.011737f
C2994 VDDA.n115 GNDA 0.012171f
C2995 VDDA.n116 GNDA 0.012171f
C2996 VDDA.n122 GNDA 0.010867f
C2997 VDDA.n123 GNDA 0.010867f
C2998 VDDA.n124 GNDA 0.011737f
C2999 VDDA.n130 GNDA 0.012171f
C3000 VDDA.n131 GNDA 0.011737f
C3001 VDDA.n132 GNDA 0.010867f
C3002 VDDA.n138 GNDA 0.011737f
C3003 VDDA.n139 GNDA 0.012171f
C3004 VDDA.n140 GNDA 0.012171f
C3005 VDDA.n146 GNDA 0.010867f
C3006 VDDA.n147 GNDA 0.010867f
C3007 VDDA.n148 GNDA 0.011737f
C3008 VDDA.n154 GNDA 0.012171f
C3009 VDDA.n155 GNDA 0.011737f
C3010 VDDA.n156 GNDA 0.010867f
C3011 VDDA.n162 GNDA 0.011737f
C3012 VDDA.n163 GNDA 0.012171f
C3013 VDDA.n164 GNDA 0.012171f
C3014 VDDA.n170 GNDA 0.010867f
C3015 VDDA.n171 GNDA 0.010867f
C3016 VDDA.n172 GNDA 0.011737f
C3017 VDDA.n178 GNDA 0.012171f
C3018 VDDA.n179 GNDA 0.011737f
C3019 VDDA.n180 GNDA 0.14168f
C3020 VDDA.n181 GNDA 0.011737f
C3021 VDDA.t195 GNDA 0.080998f
C3022 VDDA.t102 GNDA 0.081291f
C3023 VDDA.t185 GNDA 0.076944f
C3024 VDDA.t105 GNDA 0.080998f
C3025 VDDA.t167 GNDA 0.081291f
C3026 VDDA.t213 GNDA 0.076944f
C3027 VDDA.t66 GNDA 0.080998f
C3028 VDDA.t106 GNDA 0.081291f
C3029 VDDA.t57 GNDA 0.076944f
C3030 VDDA.t9 GNDA 0.080998f
C3031 VDDA.t112 GNDA 0.081291f
C3032 VDDA.t229 GNDA 0.076944f
C3033 VDDA.t110 GNDA 0.080998f
C3034 VDDA.t190 GNDA 0.081291f
C3035 VDDA.t58 GNDA 0.076944f
C3036 VDDA.n232 GNDA 0.054293f
C3037 VDDA.t118 GNDA 0.043236f
C3038 VDDA.n233 GNDA 0.058909f
C3039 VDDA.t107 GNDA 0.043236f
C3040 VDDA.n234 GNDA 0.058909f
C3041 VDDA.t228 GNDA 0.043236f
C3042 VDDA.n235 GNDA 0.058909f
C3043 VDDA.t214 GNDA 0.043236f
C3044 VDDA.n236 GNDA 0.058909f
C3045 VDDA.t73 GNDA 0.17947f
C3046 VDDA.n237 GNDA 0.29228f
C3047 VDDA.n351 GNDA 0.016551f
C3048 VDDA.n354 GNDA 2.8168f
C3049 VDDA.n381 GNDA 0.012171f
C3050 VDDA.n385 GNDA 0.011737f
C3051 VDDA.n389 GNDA 0.010867f
C3052 VDDA.n393 GNDA 0.012171f
C3053 VDDA.n397 GNDA 0.011737f
C3054 VDDA.n401 GNDA 0.010867f
C3055 VDDA.n405 GNDA 0.012171f
C3056 VDDA.n409 GNDA 0.011737f
C3057 VDDA.n413 GNDA 0.010867f
C3058 VDDA.n417 GNDA 0.012171f
C3059 VDDA.n421 GNDA 0.011737f
C3060 VDDA.n428 GNDA 0.033905f
C3061 VDDA.n429 GNDA 0.012171f
C3062 VDDA.n435 GNDA 0.010867f
C3063 VDDA.n436 GNDA 0.010867f
C3064 VDDA.n437 GNDA 0.011737f
C3065 VDDA.n443 GNDA 0.012171f
C3066 VDDA.n444 GNDA 0.011737f
C3067 VDDA.n445 GNDA 0.010867f
C3068 VDDA.n451 GNDA 0.011737f
C3069 VDDA.n452 GNDA 0.012171f
C3070 VDDA.n453 GNDA 0.012171f
C3071 VDDA.n459 GNDA 0.010867f
C3072 VDDA.n460 GNDA 0.010867f
C3073 VDDA.n461 GNDA 0.011737f
C3074 VDDA.n467 GNDA 0.012171f
C3075 VDDA.n468 GNDA 0.011737f
C3076 VDDA.n469 GNDA 0.010867f
C3077 VDDA.n475 GNDA 0.011737f
C3078 VDDA.n476 GNDA 0.012171f
C3079 VDDA.n477 GNDA 0.012171f
C3080 VDDA.n483 GNDA 0.010867f
C3081 VDDA.n484 GNDA 0.010867f
C3082 VDDA.n485 GNDA 0.011737f
C3083 VDDA.n491 GNDA 0.012171f
C3084 VDDA.n492 GNDA 0.011737f
C3085 VDDA.n493 GNDA 0.010867f
C3086 VDDA.n499 GNDA 0.011737f
C3087 VDDA.n500 GNDA 0.012171f
C3088 VDDA.n501 GNDA 0.012171f
C3089 VDDA.n507 GNDA 0.010867f
C3090 VDDA.n508 GNDA 0.010867f
C3091 VDDA.n509 GNDA 0.011737f
C3092 VDDA.n515 GNDA 0.012171f
C3093 VDDA.n516 GNDA 0.011737f
C3094 VDDA.n517 GNDA 0.14168f
C3095 VDDA.n518 GNDA 0.011737f
C3096 VDDA.n521 GNDA 1.62285f
C3097 VDDA.n548 GNDA 0.012171f
C3098 VDDA.n552 GNDA 0.011737f
C3099 VDDA.n556 GNDA 0.010867f
C3100 VDDA.n560 GNDA 0.012171f
C3101 VDDA.n564 GNDA 0.011737f
C3102 VDDA.n568 GNDA 0.010867f
C3103 VDDA.n572 GNDA 0.012171f
C3104 VDDA.n576 GNDA 0.011737f
C3105 VDDA.n580 GNDA 0.010867f
C3106 VDDA.n584 GNDA 0.012171f
C3107 VDDA.n588 GNDA 0.011737f
C3108 VDDA.n595 GNDA 0.033905f
C3109 VDDA.n596 GNDA 0.012171f
C3110 VDDA.n602 GNDA 0.010867f
C3111 VDDA.n603 GNDA 0.010867f
C3112 VDDA.n604 GNDA 0.011737f
C3113 VDDA.n610 GNDA 0.012171f
C3114 VDDA.n611 GNDA 0.011737f
C3115 VDDA.n612 GNDA 0.010867f
C3116 VDDA.n618 GNDA 0.011737f
C3117 VDDA.n619 GNDA 0.012171f
C3118 VDDA.n620 GNDA 0.012171f
C3119 VDDA.n626 GNDA 0.010867f
C3120 VDDA.n627 GNDA 0.010867f
C3121 VDDA.n628 GNDA 0.011737f
C3122 VDDA.n634 GNDA 0.012171f
C3123 VDDA.n635 GNDA 0.011737f
C3124 VDDA.n636 GNDA 0.010867f
C3125 VDDA.n642 GNDA 0.011737f
C3126 VDDA.n643 GNDA 0.012171f
C3127 VDDA.n644 GNDA 0.012171f
C3128 VDDA.n650 GNDA 0.010867f
C3129 VDDA.n651 GNDA 0.010867f
C3130 VDDA.n652 GNDA 0.011737f
C3131 VDDA.n658 GNDA 0.012171f
C3132 VDDA.n659 GNDA 0.011737f
C3133 VDDA.n660 GNDA 0.010867f
C3134 VDDA.n666 GNDA 0.011737f
C3135 VDDA.n667 GNDA 0.012171f
C3136 VDDA.n668 GNDA 0.012171f
C3137 VDDA.n674 GNDA 0.010867f
C3138 VDDA.n675 GNDA 0.010867f
C3139 VDDA.n676 GNDA 0.011737f
C3140 VDDA.n682 GNDA 0.012171f
C3141 VDDA.n683 GNDA 0.011737f
C3142 VDDA.n684 GNDA 0.011737f
C3143 VDDA.t463 GNDA 0.058946f
C3144 VDDA.t551 GNDA 0.057959f
C3145 VDDA.n687 GNDA 0.03886f
C3146 VDDA.t952 GNDA 0.057959f
C3147 VDDA.n688 GNDA 0.025357f
C3148 VDDA.t801 GNDA 0.057959f
C3149 VDDA.n689 GNDA 0.025357f
C3150 VDDA.t887 GNDA 0.057959f
C3151 VDDA.n690 GNDA 0.025357f
C3152 VDDA.t735 GNDA 0.057959f
C3153 VDDA.n691 GNDA 0.025357f
C3154 VDDA.t590 GNDA 0.057959f
C3155 VDDA.n692 GNDA 0.025357f
C3156 VDDA.t674 GNDA 0.057959f
C3157 VDDA.n693 GNDA 0.025357f
C3158 VDDA.t526 GNDA 0.057959f
C3159 VDDA.t578 GNDA 0.058946f
C3160 VDDA.t727 GNDA 0.057959f
C3161 VDDA.n694 GNDA 0.03886f
C3162 VDDA.t877 GNDA 0.057959f
C3163 VDDA.n695 GNDA 0.025357f
C3164 VDDA.t792 GNDA 0.057959f
C3165 VDDA.n696 GNDA 0.025357f
C3166 VDDA.t715 GNDA 0.057959f
C3167 VDDA.n697 GNDA 0.025357f
C3168 VDDA.t866 GNDA 0.057959f
C3169 VDDA.n698 GNDA 0.025357f
C3170 VDDA.t782 GNDA 0.057959f
C3171 VDDA.n699 GNDA 0.025357f
C3172 VDDA.t928 GNDA 0.057959f
C3173 VDDA.n700 GNDA 0.025357f
C3174 VDDA.n701 GNDA 0.036224f
C3175 VDDA.t855 GNDA 0.058946f
C3176 VDDA.t943 GNDA 0.057959f
C3177 VDDA.n702 GNDA 0.03886f
C3178 VDDA.t796 GNDA 0.057959f
C3179 VDDA.n703 GNDA 0.025357f
C3180 VDDA.t643 GNDA 0.057959f
C3181 VDDA.n704 GNDA 0.025357f
C3182 VDDA.t728 GNDA 0.057959f
C3183 VDDA.n705 GNDA 0.025357f
C3184 VDDA.t580 GNDA 0.057959f
C3185 VDDA.n706 GNDA 0.025357f
C3186 VDDA.t434 GNDA 0.057959f
C3187 VDDA.n707 GNDA 0.025357f
C3188 VDDA.t516 GNDA 0.057959f
C3189 VDDA.n708 GNDA 0.025357f
C3190 VDDA.t919 GNDA 0.057959f
C3191 VDDA.t423 GNDA 0.058946f
C3192 VDDA.t571 GNDA 0.057959f
C3193 VDDA.n709 GNDA 0.03886f
C3194 VDDA.t719 GNDA 0.057959f
C3195 VDDA.n710 GNDA 0.025357f
C3196 VDDA.t633 GNDA 0.057959f
C3197 VDDA.n711 GNDA 0.025357f
C3198 VDDA.t560 GNDA 0.057959f
C3199 VDDA.n712 GNDA 0.025357f
C3200 VDDA.t708 GNDA 0.057959f
C3201 VDDA.n713 GNDA 0.025357f
C3202 VDDA.t623 GNDA 0.057959f
C3203 VDDA.n714 GNDA 0.025357f
C3204 VDDA.t772 GNDA 0.057959f
C3205 VDDA.n715 GNDA 0.025357f
C3206 VDDA.n716 GNDA 0.047092f
C3207 VDDA.t446 GNDA 0.058946f
C3208 VDDA.t529 GNDA 0.057959f
C3209 VDDA.n717 GNDA 0.03886f
C3210 VDDA.t931 GNDA 0.057959f
C3211 VDDA.n718 GNDA 0.025357f
C3212 VDDA.t784 GNDA 0.057959f
C3213 VDDA.n719 GNDA 0.025357f
C3214 VDDA.t867 GNDA 0.057959f
C3215 VDDA.n720 GNDA 0.025357f
C3216 VDDA.t718 GNDA 0.057959f
C3217 VDDA.n721 GNDA 0.025357f
C3218 VDDA.t569 GNDA 0.057959f
C3219 VDDA.n722 GNDA 0.025357f
C3220 VDDA.t652 GNDA 0.057959f
C3221 VDDA.n723 GNDA 0.025357f
C3222 VDDA.t505 GNDA 0.057959f
C3223 VDDA.t559 GNDA 0.058946f
C3224 VDDA.t707 GNDA 0.057959f
C3225 VDDA.n724 GNDA 0.03886f
C3226 VDDA.t857 GNDA 0.057959f
C3227 VDDA.n725 GNDA 0.025357f
C3228 VDDA.t770 GNDA 0.057959f
C3229 VDDA.n726 GNDA 0.025357f
C3230 VDDA.t695 GNDA 0.057959f
C3231 VDDA.n727 GNDA 0.025357f
C3232 VDDA.t845 GNDA 0.057959f
C3233 VDDA.n728 GNDA 0.025357f
C3234 VDDA.t758 GNDA 0.057959f
C3235 VDDA.n729 GNDA 0.025357f
C3236 VDDA.t906 GNDA 0.057959f
C3237 VDDA.n730 GNDA 0.025357f
C3238 VDDA.n731 GNDA 0.047092f
C3239 VDDA.t835 GNDA 0.058946f
C3240 VDDA.t920 GNDA 0.057959f
C3241 VDDA.n732 GNDA 0.03886f
C3242 VDDA.t775 GNDA 0.057959f
C3243 VDDA.n733 GNDA 0.025357f
C3244 VDDA.t626 GNDA 0.057959f
C3245 VDDA.n734 GNDA 0.025357f
C3246 VDDA.t709 GNDA 0.057959f
C3247 VDDA.n735 GNDA 0.025357f
C3248 VDDA.t563 GNDA 0.057959f
C3249 VDDA.n736 GNDA 0.025357f
C3250 VDDA.t963 GNDA 0.057959f
C3251 VDDA.n737 GNDA 0.025357f
C3252 VDDA.t496 GNDA 0.057959f
C3253 VDDA.n738 GNDA 0.025357f
C3254 VDDA.t899 GNDA 0.057959f
C3255 VDDA.t954 GNDA 0.058946f
C3256 VDDA.t553 GNDA 0.057959f
C3257 VDDA.n739 GNDA 0.03886f
C3258 VDDA.t698 GNDA 0.057959f
C3259 VDDA.n740 GNDA 0.025357f
C3260 VDDA.t614 GNDA 0.057959f
C3261 VDDA.n741 GNDA 0.025357f
C3262 VDDA.t541 GNDA 0.057959f
C3263 VDDA.n742 GNDA 0.025357f
C3264 VDDA.t688 GNDA 0.057959f
C3265 VDDA.n743 GNDA 0.025357f
C3266 VDDA.t603 GNDA 0.057959f
C3267 VDDA.n744 GNDA 0.025357f
C3268 VDDA.t750 GNDA 0.057959f
C3269 VDDA.n745 GNDA 0.025357f
C3270 VDDA.n746 GNDA 0.047092f
C3271 VDDA.t679 GNDA 0.058946f
C3272 VDDA.t764 GNDA 0.057959f
C3273 VDDA.n747 GNDA 0.03886f
C3274 VDDA.t619 GNDA 0.057959f
C3275 VDDA.n748 GNDA 0.025357f
C3276 VDDA.t471 GNDA 0.057959f
C3277 VDDA.n749 GNDA 0.025357f
C3278 VDDA.t555 GNDA 0.057959f
C3279 VDDA.n750 GNDA 0.025357f
C3280 VDDA.t958 GNDA 0.057959f
C3281 VDDA.n751 GNDA 0.025357f
C3282 VDDA.t807 GNDA 0.057959f
C3283 VDDA.n752 GNDA 0.025357f
C3284 VDDA.t892 GNDA 0.057959f
C3285 VDDA.n753 GNDA 0.025357f
C3286 VDDA.t743 GNDA 0.057959f
C3287 VDDA.t798 GNDA 0.058946f
C3288 VDDA.t946 GNDA 0.057959f
C3289 VDDA.n754 GNDA 0.03886f
C3290 VDDA.t546 GNDA 0.057959f
C3291 VDDA.n755 GNDA 0.025357f
C3292 VDDA.t459 GNDA 0.057959f
C3293 VDDA.n756 GNDA 0.025357f
C3294 VDDA.t933 GNDA 0.057959f
C3295 VDDA.n757 GNDA 0.025357f
C3296 VDDA.t534 GNDA 0.057959f
C3297 VDDA.n758 GNDA 0.025357f
C3298 VDDA.t448 GNDA 0.057959f
C3299 VDDA.n759 GNDA 0.025357f
C3300 VDDA.t596 GNDA 0.057959f
C3301 VDDA.n760 GNDA 0.025357f
C3302 VDDA.n761 GNDA 0.047092f
C3303 VDDA.t814 GNDA 0.058946f
C3304 VDDA.t901 GNDA 0.057959f
C3305 VDDA.n762 GNDA 0.03886f
C3306 VDDA.t752 GNDA 0.057959f
C3307 VDDA.n763 GNDA 0.025357f
C3308 VDDA.t605 GNDA 0.057959f
C3309 VDDA.n764 GNDA 0.025357f
C3310 VDDA.t690 GNDA 0.057959f
C3311 VDDA.n765 GNDA 0.025357f
C3312 VDDA.t544 GNDA 0.057959f
C3313 VDDA.n766 GNDA 0.025357f
C3314 VDDA.t947 GNDA 0.057959f
C3315 VDDA.n767 GNDA 0.025357f
C3316 VDDA.t481 GNDA 0.057959f
C3317 VDDA.n768 GNDA 0.025357f
C3318 VDDA.t881 GNDA 0.057959f
C3319 VDDA.t932 GNDA 0.058946f
C3320 VDDA.t533 GNDA 0.057959f
C3321 VDDA.n769 GNDA 0.03886f
C3322 VDDA.t680 GNDA 0.057959f
C3323 VDDA.n770 GNDA 0.025357f
C3324 VDDA.t594 GNDA 0.057959f
C3325 VDDA.n771 GNDA 0.025357f
C3326 VDDA.t517 GNDA 0.057959f
C3327 VDDA.n772 GNDA 0.025357f
C3328 VDDA.t666 GNDA 0.057959f
C3329 VDDA.n773 GNDA 0.025357f
C3330 VDDA.t583 GNDA 0.057959f
C3331 VDDA.n774 GNDA 0.025357f
C3332 VDDA.t730 GNDA 0.057959f
C3333 VDDA.n775 GNDA 0.025357f
C3334 VDDA.n776 GNDA 0.047092f
C3335 VDDA.t656 GNDA 0.058946f
C3336 VDDA.t744 GNDA 0.057959f
C3337 VDDA.n777 GNDA 0.03886f
C3338 VDDA.t598 GNDA 0.057959f
C3339 VDDA.n778 GNDA 0.025357f
C3340 VDDA.t450 GNDA 0.057959f
C3341 VDDA.n779 GNDA 0.025357f
C3342 VDDA.t535 GNDA 0.057959f
C3343 VDDA.n780 GNDA 0.025357f
C3344 VDDA.t936 GNDA 0.057959f
C3345 VDDA.n781 GNDA 0.025357f
C3346 VDDA.t787 GNDA 0.057959f
C3347 VDDA.n782 GNDA 0.025357f
C3348 VDDA.t872 GNDA 0.057959f
C3349 VDDA.n783 GNDA 0.025357f
C3350 VDDA.t722 GNDA 0.057959f
C3351 VDDA.t776 GNDA 0.058946f
C3352 VDDA.t923 GNDA 0.057959f
C3353 VDDA.n784 GNDA 0.03886f
C3354 VDDA.t520 GNDA 0.057959f
C3355 VDDA.n785 GNDA 0.025357f
C3356 VDDA.t439 GNDA 0.057959f
C3357 VDDA.n786 GNDA 0.025357f
C3358 VDDA.t909 GNDA 0.057959f
C3359 VDDA.n787 GNDA 0.025357f
C3360 VDDA.t509 GNDA 0.057959f
C3361 VDDA.n788 GNDA 0.025357f
C3362 VDDA.t427 GNDA 0.057959f
C3363 VDDA.n789 GNDA 0.025357f
C3364 VDDA.t573 GNDA 0.057959f
C3365 VDDA.n790 GNDA 0.025357f
C3366 VDDA.n791 GNDA 0.047092f
C3367 VDDA.t522 GNDA 0.058946f
C3368 VDDA.t610 GNDA 0.057959f
C3369 VDDA.n792 GNDA 0.03886f
C3370 VDDA.t464 GNDA 0.057959f
C3371 VDDA.n793 GNDA 0.025357f
C3372 VDDA.t863 GNDA 0.057959f
C3373 VDDA.n794 GNDA 0.025357f
C3374 VDDA.t950 GNDA 0.057959f
C3375 VDDA.n795 GNDA 0.025357f
C3376 VDDA.t802 GNDA 0.057959f
C3377 VDDA.n796 GNDA 0.025357f
C3378 VDDA.t649 GNDA 0.057959f
C3379 VDDA.n797 GNDA 0.025357f
C3380 VDDA.t733 GNDA 0.057959f
C3381 VDDA.n798 GNDA 0.025357f
C3382 VDDA.t587 GNDA 0.057959f
C3383 VDDA.t639 GNDA 0.058946f
C3384 VDDA.t790 GNDA 0.057959f
C3385 VDDA.n799 GNDA 0.03886f
C3386 VDDA.t940 GNDA 0.057959f
C3387 VDDA.n800 GNDA 0.025357f
C3388 VDDA.t850 GNDA 0.057959f
C3389 VDDA.n801 GNDA 0.025357f
C3390 VDDA.t780 GNDA 0.057959f
C3391 VDDA.n802 GNDA 0.025357f
C3392 VDDA.t926 GNDA 0.057959f
C3393 VDDA.n803 GNDA 0.025357f
C3394 VDDA.t838 GNDA 0.057959f
C3395 VDDA.n804 GNDA 0.025357f
C3396 VDDA.t443 GNDA 0.057959f
C3397 VDDA.n805 GNDA 0.025357f
C3398 VDDA.n806 GNDA 0.047092f
C3399 VDDA.t659 GNDA 0.058946f
C3400 VDDA.t746 GNDA 0.057959f
C3401 VDDA.n807 GNDA 0.03886f
C3402 VDDA.t599 GNDA 0.057959f
C3403 VDDA.n808 GNDA 0.025357f
C3404 VDDA.t452 GNDA 0.057959f
C3405 VDDA.n809 GNDA 0.025357f
C3406 VDDA.t537 GNDA 0.057959f
C3407 VDDA.n810 GNDA 0.025357f
C3408 VDDA.t937 GNDA 0.057959f
C3409 VDDA.n811 GNDA 0.025357f
C3410 VDDA.t791 GNDA 0.057959f
C3411 VDDA.n812 GNDA 0.025357f
C3412 VDDA.t874 GNDA 0.057959f
C3413 VDDA.n813 GNDA 0.025357f
C3414 VDDA.t723 GNDA 0.057959f
C3415 VDDA.t777 GNDA 0.058946f
C3416 VDDA.t925 GNDA 0.057959f
C3417 VDDA.n814 GNDA 0.03886f
C3418 VDDA.t524 GNDA 0.057959f
C3419 VDDA.n815 GNDA 0.025357f
C3420 VDDA.t440 GNDA 0.057959f
C3421 VDDA.n816 GNDA 0.025357f
C3422 VDDA.t914 GNDA 0.057959f
C3423 VDDA.n817 GNDA 0.025357f
C3424 VDDA.t510 GNDA 0.057959f
C3425 VDDA.n818 GNDA 0.025357f
C3426 VDDA.t431 GNDA 0.057959f
C3427 VDDA.n819 GNDA 0.025357f
C3428 VDDA.t577 GNDA 0.057959f
C3429 VDDA.n820 GNDA 0.025357f
C3430 VDDA.n821 GNDA 0.047092f
C3431 VDDA.t503 GNDA 0.058946f
C3432 VDDA.t591 GNDA 0.057959f
C3433 VDDA.n822 GNDA 0.03886f
C3434 VDDA.t445 GNDA 0.057959f
C3435 VDDA.n823 GNDA 0.025357f
C3436 VDDA.t842 GNDA 0.057959f
C3437 VDDA.n824 GNDA 0.025357f
C3438 VDDA.t929 GNDA 0.057959f
C3439 VDDA.n825 GNDA 0.025357f
C3440 VDDA.t783 GNDA 0.057959f
C3441 VDDA.n826 GNDA 0.025357f
C3442 VDDA.t632 GNDA 0.057959f
C3443 VDDA.n827 GNDA 0.025357f
C3444 VDDA.t716 GNDA 0.057959f
C3445 VDDA.n828 GNDA 0.025357f
C3446 VDDA.t568 GNDA 0.057959f
C3447 VDDA.t621 GNDA 0.058946f
C3448 VDDA.t769 GNDA 0.057959f
C3449 VDDA.n829 GNDA 0.03886f
C3450 VDDA.t917 GNDA 0.057959f
C3451 VDDA.n830 GNDA 0.025357f
C3452 VDDA.t830 GNDA 0.057959f
C3453 VDDA.n831 GNDA 0.025357f
C3454 VDDA.t757 GNDA 0.057959f
C3455 VDDA.n832 GNDA 0.025357f
C3456 VDDA.t905 GNDA 0.057959f
C3457 VDDA.n833 GNDA 0.025357f
C3458 VDDA.t821 GNDA 0.057959f
C3459 VDDA.n834 GNDA 0.025357f
C3460 VDDA.t422 GNDA 0.057959f
C3461 VDDA.n835 GNDA 0.025357f
C3462 VDDA.n836 GNDA 0.047092f
C3463 VDDA.t896 GNDA 0.058946f
C3464 VDDA.t436 GNDA 0.057959f
C3465 VDDA.n837 GNDA 0.03886f
C3466 VDDA.t834 GNDA 0.057959f
C3467 VDDA.n838 GNDA 0.025357f
C3468 VDDA.t684 GNDA 0.057959f
C3469 VDDA.n839 GNDA 0.025357f
C3470 VDDA.t773 GNDA 0.057959f
C3471 VDDA.n840 GNDA 0.025357f
C3472 VDDA.t624 GNDA 0.057959f
C3473 VDDA.n841 GNDA 0.025357f
C3474 VDDA.t476 GNDA 0.057959f
C3475 VDDA.n842 GNDA 0.025357f
C3476 VDDA.t561 GNDA 0.057959f
C3477 VDDA.n843 GNDA 0.025357f
C3478 VDDA.t962 GNDA 0.057959f
C3479 VDDA.t466 GNDA 0.058946f
C3480 VDDA.t613 GNDA 0.057959f
C3481 VDDA.n844 GNDA 0.03886f
C3482 VDDA.t761 GNDA 0.057959f
C3483 VDDA.n845 GNDA 0.025357f
C3484 VDDA.t670 GNDA 0.057959f
C3485 VDDA.n846 GNDA 0.025357f
C3486 VDDA.t602 GNDA 0.057959f
C3487 VDDA.n847 GNDA 0.025357f
C3488 VDDA.t749 GNDA 0.057959f
C3489 VDDA.n848 GNDA 0.025357f
C3490 VDDA.t663 GNDA 0.057959f
C3491 VDDA.n849 GNDA 0.025357f
C3492 VDDA.t813 GNDA 0.057959f
C3493 VDDA.n850 GNDA 0.025357f
C3494 VDDA.n851 GNDA 0.047092f
C3495 VDDA.t738 GNDA 0.058946f
C3496 VDDA.t825 GNDA 0.057959f
C3497 VDDA.n852 GNDA 0.03886f
C3498 VDDA.t677 GNDA 0.057959f
C3499 VDDA.n853 GNDA 0.025357f
C3500 VDDA.t530 GNDA 0.057959f
C3501 VDDA.n854 GNDA 0.025357f
C3502 VDDA.t616 GNDA 0.057959f
C3503 VDDA.n855 GNDA 0.025357f
C3504 VDDA.t468 GNDA 0.057959f
C3505 VDDA.n856 GNDA 0.025357f
C3506 VDDA.t869 GNDA 0.057959f
C3507 VDDA.n857 GNDA 0.025357f
C3508 VDDA.t956 GNDA 0.057959f
C3509 VDDA.n858 GNDA 0.025357f
C3510 VDDA.t806 GNDA 0.057959f
C3511 VDDA.t858 GNDA 0.058946f
C3512 VDDA.t458 GNDA 0.057959f
C3513 VDDA.n859 GNDA 0.03886f
C3514 VDDA.t606 GNDA 0.057959f
C3515 VDDA.n860 GNDA 0.025357f
C3516 VDDA.t514 GNDA 0.057959f
C3517 VDDA.n861 GNDA 0.025357f
C3518 VDDA.t449 GNDA 0.057959f
C3519 VDDA.n862 GNDA 0.025357f
C3520 VDDA.t595 GNDA 0.057959f
C3521 VDDA.n863 GNDA 0.025357f
C3522 VDDA.t506 GNDA 0.057959f
C3523 VDDA.n864 GNDA 0.025357f
C3524 VDDA.t655 GNDA 0.057959f
C3525 VDDA.n865 GNDA 0.025357f
C3526 VDDA.n866 GNDA 0.047092f
C3527 VDDA.t879 GNDA 0.058946f
C3528 VDDA.t965 GNDA 0.057959f
C3529 VDDA.n867 GNDA 0.03886f
C3530 VDDA.t815 GNDA 0.057959f
C3531 VDDA.n868 GNDA 0.025357f
C3532 VDDA.t664 GNDA 0.057959f
C3533 VDDA.n869 GNDA 0.025357f
C3534 VDDA.t751 GNDA 0.057959f
C3535 VDDA.n870 GNDA 0.025357f
C3536 VDDA.t604 GNDA 0.057959f
C3537 VDDA.n871 GNDA 0.025357f
C3538 VDDA.t457 GNDA 0.057959f
C3539 VDDA.n872 GNDA 0.025357f
C3540 VDDA.t542 GNDA 0.057959f
C3541 VDDA.n873 GNDA 0.025357f
C3542 VDDA.t944 GNDA 0.057959f
C3543 VDDA.t447 GNDA 0.058946f
C3544 VDDA.t593 GNDA 0.057959f
C3545 VDDA.n874 GNDA 0.03886f
C3546 VDDA.t740 GNDA 0.057959f
C3547 VDDA.n875 GNDA 0.025357f
C3548 VDDA.t653 GNDA 0.057959f
C3549 VDDA.n876 GNDA 0.025357f
C3550 VDDA.t581 GNDA 0.057959f
C3551 VDDA.n877 GNDA 0.025357f
C3552 VDDA.t729 GNDA 0.057959f
C3553 VDDA.n878 GNDA 0.025357f
C3554 VDDA.t645 GNDA 0.057959f
C3555 VDDA.n879 GNDA 0.025357f
C3556 VDDA.t797 GNDA 0.057959f
C3557 VDDA.n880 GNDA 0.025357f
C3558 VDDA.n881 GNDA 0.047092f
C3559 VDDA.t720 GNDA 0.058946f
C3560 VDDA.t809 GNDA 0.057959f
C3561 VDDA.n882 GNDA 0.03886f
C3562 VDDA.t657 GNDA 0.057959f
C3563 VDDA.n883 GNDA 0.025357f
C3564 VDDA.t507 GNDA 0.057959f
C3565 VDDA.n884 GNDA 0.025357f
C3566 VDDA.t597 GNDA 0.057959f
C3567 VDDA.n885 GNDA 0.025357f
C3568 VDDA.t451 GNDA 0.057959f
C3569 VDDA.n886 GNDA 0.025357f
C3570 VDDA.t847 GNDA 0.057959f
C3571 VDDA.n887 GNDA 0.025357f
C3572 VDDA.t934 GNDA 0.057959f
C3573 VDDA.n888 GNDA 0.025357f
C3574 VDDA.t786 GNDA 0.057959f
C3575 VDDA.t836 GNDA 0.058946f
C3576 VDDA.t438 GNDA 0.057959f
C3577 VDDA.n889 GNDA 0.03886f
C3578 VDDA.t585 GNDA 0.057959f
C3579 VDDA.n890 GNDA 0.025357f
C3580 VDDA.t497 GNDA 0.057959f
C3581 VDDA.n891 GNDA 0.025357f
C3582 VDDA.t426 GNDA 0.057959f
C3583 VDDA.n892 GNDA 0.025357f
C3584 VDDA.t572 GNDA 0.057959f
C3585 VDDA.n893 GNDA 0.025357f
C3586 VDDA.t488 GNDA 0.057959f
C3587 VDDA.n894 GNDA 0.025357f
C3588 VDDA.t636 GNDA 0.057959f
C3589 VDDA.n895 GNDA 0.025357f
C3590 VDDA.n896 GNDA 0.047092f
C3591 VDDA.t565 GNDA 0.058946f
C3592 VDDA.t647 GNDA 0.057959f
C3593 VDDA.n897 GNDA 0.03886f
C3594 VDDA.t500 GNDA 0.057959f
C3595 VDDA.n898 GNDA 0.025357f
C3596 VDDA.t902 GNDA 0.057959f
C3597 VDDA.n899 GNDA 0.025357f
C3598 VDDA.t441 GNDA 0.057959f
C3599 VDDA.n900 GNDA 0.025357f
C3600 VDDA.t839 GNDA 0.057959f
C3601 VDDA.n901 GNDA 0.025357f
C3602 VDDA.t691 GNDA 0.057959f
C3603 VDDA.n902 GNDA 0.025357f
C3604 VDDA.t778 GNDA 0.057959f
C3605 VDDA.n903 GNDA 0.025357f
C3606 VDDA.t630 GNDA 0.057959f
C3607 VDDA.t681 GNDA 0.058946f
C3608 VDDA.t828 GNDA 0.057959f
C3609 VDDA.n904 GNDA 0.03886f
C3610 VDDA.t432 GNDA 0.057959f
C3611 VDDA.n905 GNDA 0.025357f
C3612 VDDA.t893 GNDA 0.057959f
C3613 VDDA.n906 GNDA 0.025357f
C3614 VDDA.t818 GNDA 0.057959f
C3615 VDDA.n907 GNDA 0.025357f
C3616 VDDA.t968 GNDA 0.057959f
C3617 VDDA.n908 GNDA 0.025357f
C3618 VDDA.t883 GNDA 0.057959f
C3619 VDDA.n909 GNDA 0.025357f
C3620 VDDA.t482 GNDA 0.057959f
C3621 VDDA.n910 GNDA 0.025357f
C3622 VDDA.n911 GNDA 0.047092f
C3623 VDDA.t699 GNDA 0.058946f
C3624 VDDA.t788 GNDA 0.057959f
C3625 VDDA.n912 GNDA 0.03886f
C3626 VDDA.t638 GNDA 0.057959f
C3627 VDDA.n913 GNDA 0.025357f
C3628 VDDA.t491 GNDA 0.057959f
C3629 VDDA.n914 GNDA 0.025357f
C3630 VDDA.t575 GNDA 0.057959f
C3631 VDDA.n915 GNDA 0.025357f
C3632 VDDA.t429 GNDA 0.057959f
C3633 VDDA.n916 GNDA 0.025357f
C3634 VDDA.t829 GNDA 0.057959f
C3635 VDDA.n917 GNDA 0.025357f
C3636 VDDA.t912 GNDA 0.057959f
C3637 VDDA.n918 GNDA 0.025357f
C3638 VDDA.t765 GNDA 0.057959f
C3639 VDDA.t816 GNDA 0.058946f
C3640 VDDA.t967 GNDA 0.057959f
C3641 VDDA.n919 GNDA 0.03886f
C3642 VDDA.t566 GNDA 0.057959f
C3643 VDDA.n920 GNDA 0.025357f
C3644 VDDA.t479 GNDA 0.057959f
C3645 VDDA.n921 GNDA 0.025357f
C3646 VDDA.t959 GNDA 0.057959f
C3647 VDDA.n922 GNDA 0.025357f
C3648 VDDA.t556 GNDA 0.057959f
C3649 VDDA.n923 GNDA 0.025357f
C3650 VDDA.t472 GNDA 0.057959f
C3651 VDDA.n924 GNDA 0.025357f
C3652 VDDA.t620 GNDA 0.057959f
C3653 VDDA.n925 GNDA 0.025357f
C3654 VDDA.n926 GNDA 0.047092f
C3655 VDDA.t547 GNDA 0.058946f
C3656 VDDA.t631 GNDA 0.057959f
C3657 VDDA.n927 GNDA 0.03886f
C3658 VDDA.t484 GNDA 0.057959f
C3659 VDDA.n928 GNDA 0.025357f
C3660 VDDA.t885 GNDA 0.057959f
C3661 VDDA.n929 GNDA 0.025357f
C3662 VDDA.t421 GNDA 0.057959f
C3663 VDDA.n930 GNDA 0.025357f
C3664 VDDA.t820 GNDA 0.057959f
C3665 VDDA.n931 GNDA 0.025357f
C3666 VDDA.t668 GNDA 0.057959f
C3667 VDDA.n932 GNDA 0.025357f
C3668 VDDA.t756 GNDA 0.057959f
C3669 VDDA.n933 GNDA 0.025357f
C3670 VDDA.t609 GNDA 0.057959f
C3671 VDDA.t658 GNDA 0.058946f
C3672 VDDA.t810 GNDA 0.057959f
C3673 VDDA.n934 GNDA 0.03886f
C3674 VDDA.t960 GNDA 0.057959f
C3675 VDDA.n935 GNDA 0.025357f
C3676 VDDA.t871 GNDA 0.057959f
C3677 VDDA.n936 GNDA 0.025357f
C3678 VDDA.t799 GNDA 0.057959f
C3679 VDDA.n937 GNDA 0.025357f
C3680 VDDA.t949 GNDA 0.057959f
C3681 VDDA.n938 GNDA 0.025357f
C3682 VDDA.t861 GNDA 0.057959f
C3683 VDDA.n939 GNDA 0.025357f
C3684 VDDA.t461 GNDA 0.057959f
C3685 VDDA.n940 GNDA 0.025357f
C3686 VDDA.n941 GNDA 0.047092f
C3687 VDDA.t938 GNDA 0.058946f
C3688 VDDA.t474 GNDA 0.057959f
C3689 VDDA.n942 GNDA 0.03886f
C3690 VDDA.t875 GNDA 0.057959f
C3691 VDDA.n943 GNDA 0.025357f
C3692 VDDA.t724 GNDA 0.057959f
C3693 VDDA.n944 GNDA 0.025357f
C3694 VDDA.t811 GNDA 0.057959f
C3695 VDDA.n945 GNDA 0.025357f
C3696 VDDA.t661 GNDA 0.057959f
C3697 VDDA.n946 GNDA 0.025357f
C3698 VDDA.t512 GNDA 0.057959f
C3699 VDDA.n947 GNDA 0.025357f
C3700 VDDA.t601 GNDA 0.057959f
C3701 VDDA.n948 GNDA 0.025357f
C3702 VDDA.t455 GNDA 0.057959f
C3703 VDDA.t502 GNDA 0.058946f
C3704 VDDA.t651 GNDA 0.057959f
C3705 VDDA.n949 GNDA 0.03886f
C3706 VDDA.t804 GNDA 0.057959f
C3707 VDDA.n950 GNDA 0.025357f
C3708 VDDA.t714 GNDA 0.057959f
C3709 VDDA.n951 GNDA 0.025357f
C3710 VDDA.t641 GNDA 0.057959f
C3711 VDDA.n952 GNDA 0.025357f
C3712 VDDA.t793 GNDA 0.057959f
C3713 VDDA.n953 GNDA 0.025357f
C3714 VDDA.t704 GNDA 0.057959f
C3715 VDDA.n954 GNDA 0.025357f
C3716 VDDA.t853 GNDA 0.057959f
C3717 VDDA.n955 GNDA 0.025357f
C3718 VDDA.n956 GNDA 0.047092f
C3719 VDDA.t523 GNDA 0.058946f
C3720 VDDA.t611 GNDA 0.057959f
C3721 VDDA.n957 GNDA 0.03886f
C3722 VDDA.t465 GNDA 0.057959f
C3723 VDDA.n958 GNDA 0.025357f
C3724 VDDA.t864 GNDA 0.057959f
C3725 VDDA.n959 GNDA 0.025357f
C3726 VDDA.t951 GNDA 0.057959f
C3727 VDDA.n960 GNDA 0.025357f
C3728 VDDA.t803 GNDA 0.057959f
C3729 VDDA.n961 GNDA 0.025357f
C3730 VDDA.t650 GNDA 0.057959f
C3731 VDDA.n962 GNDA 0.025357f
C3732 VDDA.t736 GNDA 0.057959f
C3733 VDDA.n963 GNDA 0.025357f
C3734 VDDA.t588 GNDA 0.057959f
C3735 VDDA.t640 GNDA 0.058946f
C3736 VDDA.t794 GNDA 0.057959f
C3737 VDDA.n964 GNDA 0.03886f
C3738 VDDA.t941 GNDA 0.057959f
C3739 VDDA.n965 GNDA 0.025357f
C3740 VDDA.t851 GNDA 0.057959f
C3741 VDDA.n966 GNDA 0.025357f
C3742 VDDA.t781 GNDA 0.057959f
C3743 VDDA.n967 GNDA 0.025357f
C3744 VDDA.t927 GNDA 0.057959f
C3745 VDDA.n968 GNDA 0.025357f
C3746 VDDA.t841 GNDA 0.057959f
C3747 VDDA.n969 GNDA 0.025357f
C3748 VDDA.t444 GNDA 0.057959f
C3749 VDDA.n970 GNDA 0.025357f
C3750 VDDA.n971 GNDA 0.047092f
C3751 VDDA.t916 GNDA 0.058946f
C3752 VDDA.t456 GNDA 0.057959f
C3753 VDDA.n972 GNDA 0.03886f
C3754 VDDA.t856 GNDA 0.057959f
C3755 VDDA.n973 GNDA 0.025357f
C3756 VDDA.t706 GNDA 0.057959f
C3757 VDDA.n974 GNDA 0.025357f
C3758 VDDA.t795 GNDA 0.057959f
C3759 VDDA.n975 GNDA 0.025357f
C3760 VDDA.t644 GNDA 0.057959f
C3761 VDDA.n976 GNDA 0.025357f
C3762 VDDA.t494 GNDA 0.057959f
C3763 VDDA.n977 GNDA 0.025357f
C3764 VDDA.t582 GNDA 0.057959f
C3765 VDDA.n978 GNDA 0.025357f
C3766 VDDA.t435 GNDA 0.057959f
C3767 VDDA.t485 GNDA 0.058946f
C3768 VDDA.t634 GNDA 0.057959f
C3769 VDDA.n979 GNDA 0.03886f
C3770 VDDA.t785 GNDA 0.057959f
C3771 VDDA.n980 GNDA 0.025357f
C3772 VDDA.t694 GNDA 0.057959f
C3773 VDDA.n981 GNDA 0.025357f
C3774 VDDA.t622 GNDA 0.057959f
C3775 VDDA.n982 GNDA 0.025357f
C3776 VDDA.t771 GNDA 0.057959f
C3777 VDDA.n983 GNDA 0.025357f
C3778 VDDA.t683 GNDA 0.057959f
C3779 VDDA.n984 GNDA 0.025357f
C3780 VDDA.t832 GNDA 0.057959f
C3781 VDDA.n985 GNDA 0.025357f
C3782 VDDA.n986 GNDA 0.047092f
C3783 VDDA.t760 GNDA 0.058946f
C3784 VDDA.t846 GNDA 0.057959f
C3785 VDDA.n987 GNDA 0.03886f
C3786 VDDA.t697 GNDA 0.057959f
C3787 VDDA.n988 GNDA 0.025357f
C3788 VDDA.t552 GNDA 0.057959f
C3789 VDDA.n989 GNDA 0.025357f
C3790 VDDA.t635 GNDA 0.057959f
C3791 VDDA.n990 GNDA 0.025357f
C3792 VDDA.t487 GNDA 0.057959f
C3793 VDDA.n991 GNDA 0.025357f
C3794 VDDA.t888 GNDA 0.057959f
C3795 VDDA.n992 GNDA 0.025357f
C3796 VDDA.t424 GNDA 0.057959f
C3797 VDDA.n993 GNDA 0.025357f
C3798 VDDA.t824 GNDA 0.057959f
C3799 VDDA.t878 GNDA 0.058946f
C3800 VDDA.t477 GNDA 0.057959f
C3801 VDDA.n994 GNDA 0.03886f
C3802 VDDA.t627 GNDA 0.057959f
C3803 VDDA.n995 GNDA 0.025357f
C3804 VDDA.t540 GNDA 0.057959f
C3805 VDDA.n996 GNDA 0.025357f
C3806 VDDA.t467 GNDA 0.057959f
C3807 VDDA.n997 GNDA 0.025357f
C3808 VDDA.t615 GNDA 0.057959f
C3809 VDDA.n998 GNDA 0.025357f
C3810 VDDA.t528 GNDA 0.057959f
C3811 VDDA.n999 GNDA 0.025357f
C3812 VDDA.t675 GNDA 0.057959f
C3813 VDDA.n1000 GNDA 0.025357f
C3814 VDDA.n1001 GNDA 0.047092f
C3815 VDDA.t628 GNDA 0.058946f
C3816 VDDA.t711 GNDA 0.057959f
C3817 VDDA.n1002 GNDA 0.03886f
C3818 VDDA.t564 GNDA 0.057959f
C3819 VDDA.n1003 GNDA 0.025357f
C3820 VDDA.t966 GNDA 0.057959f
C3821 VDDA.n1004 GNDA 0.025357f
C3822 VDDA.t499 GNDA 0.057959f
C3823 VDDA.n1005 GNDA 0.025357f
C3824 VDDA.t900 GNDA 0.057959f
C3825 VDDA.n1006 GNDA 0.025357f
C3826 VDDA.t753 GNDA 0.057959f
C3827 VDDA.n1007 GNDA 0.025357f
C3828 VDDA.t837 GNDA 0.057959f
C3829 VDDA.n1008 GNDA 0.025357f
C3830 VDDA.t689 GNDA 0.057959f
C3831 VDDA.t741 GNDA 0.058946f
C3832 VDDA.t891 GNDA 0.057959f
C3833 VDDA.n1009 GNDA 0.03886f
C3834 VDDA.t492 GNDA 0.057959f
C3835 VDDA.n1010 GNDA 0.025357f
C3836 VDDA.t955 GNDA 0.057959f
C3837 VDDA.n1011 GNDA 0.025357f
C3838 VDDA.t882 GNDA 0.057959f
C3839 VDDA.n1012 GNDA 0.025357f
C3840 VDDA.t480 GNDA 0.057959f
C3841 VDDA.n1013 GNDA 0.025357f
C3842 VDDA.t945 GNDA 0.057959f
C3843 VDDA.n1014 GNDA 0.025357f
C3844 VDDA.t545 GNDA 0.057959f
C3845 VDDA.n1015 GNDA 0.025357f
C3846 VDDA.n1016 GNDA 0.047092f
C3847 VDDA.t763 GNDA 0.058946f
C3848 VDDA.t848 GNDA 0.057959f
C3849 VDDA.n1017 GNDA 0.03886f
C3850 VDDA.t700 GNDA 0.057959f
C3851 VDDA.n1018 GNDA 0.025357f
C3852 VDDA.t554 GNDA 0.057959f
C3853 VDDA.n1019 GNDA 0.025357f
C3854 VDDA.t637 GNDA 0.057959f
C3855 VDDA.n1020 GNDA 0.025357f
C3856 VDDA.t489 GNDA 0.057959f
C3857 VDDA.n1021 GNDA 0.025357f
C3858 VDDA.t890 GNDA 0.057959f
C3859 VDDA.n1022 GNDA 0.025357f
C3860 VDDA.t428 GNDA 0.057959f
C3861 VDDA.n1023 GNDA 0.025357f
C3862 VDDA.t826 GNDA 0.057959f
C3863 VDDA.t880 GNDA 0.058946f
C3864 VDDA.t478 GNDA 0.057959f
C3865 VDDA.n1024 GNDA 0.03886f
C3866 VDDA.t629 GNDA 0.057959f
C3867 VDDA.n1025 GNDA 0.025357f
C3868 VDDA.t543 GNDA 0.057959f
C3869 VDDA.n1026 GNDA 0.025357f
C3870 VDDA.t469 GNDA 0.057959f
C3871 VDDA.n1027 GNDA 0.025357f
C3872 VDDA.t617 GNDA 0.057959f
C3873 VDDA.n1028 GNDA 0.025357f
C3874 VDDA.t532 GNDA 0.057959f
C3875 VDDA.n1029 GNDA 0.025357f
C3876 VDDA.t678 GNDA 0.057959f
C3877 VDDA.n1030 GNDA 0.025357f
C3878 VDDA.n1031 GNDA 0.047092f
C3879 VDDA.t608 GNDA 0.058946f
C3880 VDDA.t692 GNDA 0.057959f
C3881 VDDA.n1032 GNDA 0.03886f
C3882 VDDA.t548 GNDA 0.057959f
C3883 VDDA.n1033 GNDA 0.025357f
C3884 VDDA.t948 GNDA 0.057959f
C3885 VDDA.n1034 GNDA 0.025357f
C3886 VDDA.t483 GNDA 0.057959f
C3887 VDDA.n1035 GNDA 0.025357f
C3888 VDDA.t884 GNDA 0.057959f
C3889 VDDA.n1036 GNDA 0.025357f
C3890 VDDA.t732 GNDA 0.057959f
C3891 VDDA.n1037 GNDA 0.025357f
C3892 VDDA.t819 GNDA 0.057959f
C3893 VDDA.n1038 GNDA 0.025357f
C3894 VDDA.t667 GNDA 0.057959f
C3895 VDDA.t721 GNDA 0.058946f
C3896 VDDA.t870 GNDA 0.057959f
C3897 VDDA.n1039 GNDA 0.03886f
C3898 VDDA.t473 GNDA 0.057959f
C3899 VDDA.n1040 GNDA 0.025357f
C3900 VDDA.t935 GNDA 0.057959f
C3901 VDDA.n1041 GNDA 0.025357f
C3902 VDDA.t859 GNDA 0.057959f
C3903 VDDA.n1042 GNDA 0.025357f
C3904 VDDA.t460 GNDA 0.057959f
C3905 VDDA.n1043 GNDA 0.025357f
C3906 VDDA.t922 GNDA 0.057959f
C3907 VDDA.n1044 GNDA 0.025357f
C3908 VDDA.t519 GNDA 0.057959f
C3909 VDDA.n1045 GNDA 0.025357f
C3910 VDDA.n1046 GNDA 0.047092f
C3911 VDDA.t453 GNDA 0.058946f
C3912 VDDA.t536 GNDA 0.057959f
C3913 VDDA.n1047 GNDA 0.03886f
C3914 VDDA.t939 GNDA 0.057959f
C3915 VDDA.n1048 GNDA 0.025357f
C3916 VDDA.t789 GNDA 0.057959f
C3917 VDDA.n1049 GNDA 0.025357f
C3918 VDDA.t873 GNDA 0.057959f
C3919 VDDA.n1050 GNDA 0.025357f
C3920 VDDA.t725 GNDA 0.057959f
C3921 VDDA.n1051 GNDA 0.025357f
C3922 VDDA.t576 GNDA 0.057959f
C3923 VDDA.n1052 GNDA 0.025357f
C3924 VDDA.t660 GNDA 0.057959f
C3925 VDDA.n1053 GNDA 0.025357f
C3926 VDDA.t511 GNDA 0.057959f
C3927 VDDA.t567 GNDA 0.058946f
C3928 VDDA.t712 GNDA 0.057959f
C3929 VDDA.n1054 GNDA 0.03886f
C3930 VDDA.t865 GNDA 0.057959f
C3931 VDDA.n1055 GNDA 0.025357f
C3932 VDDA.t779 GNDA 0.057959f
C3933 VDDA.n1056 GNDA 0.025357f
C3934 VDDA.t703 GNDA 0.057959f
C3935 VDDA.n1057 GNDA 0.025357f
C3936 VDDA.t852 GNDA 0.057959f
C3937 VDDA.n1058 GNDA 0.025357f
C3938 VDDA.t767 GNDA 0.057959f
C3939 VDDA.n1059 GNDA 0.025357f
C3940 VDDA.t913 GNDA 0.057959f
C3941 VDDA.n1060 GNDA 0.025357f
C3942 VDDA.n1061 GNDA 0.047092f
C3943 VDDA.t586 GNDA 0.058946f
C3944 VDDA.t669 GNDA 0.057959f
C3945 VDDA.n1062 GNDA 0.03886f
C3946 VDDA.t521 GNDA 0.057959f
C3947 VDDA.n1063 GNDA 0.025357f
C3948 VDDA.t924 GNDA 0.057959f
C3949 VDDA.n1064 GNDA 0.025357f
C3950 VDDA.t462 GNDA 0.057959f
C3951 VDDA.n1065 GNDA 0.025357f
C3952 VDDA.t862 GNDA 0.057959f
C3953 VDDA.n1066 GNDA 0.025357f
C3954 VDDA.t713 GNDA 0.057959f
C3955 VDDA.n1067 GNDA 0.025357f
C3956 VDDA.t800 GNDA 0.057959f
C3957 VDDA.n1068 GNDA 0.025357f
C3958 VDDA.t648 GNDA 0.057959f
C3959 VDDA.t701 GNDA 0.058946f
C3960 VDDA.t849 GNDA 0.057959f
C3961 VDDA.n1069 GNDA 0.03886f
C3962 VDDA.t454 GNDA 0.057959f
C3963 VDDA.n1070 GNDA 0.025357f
C3964 VDDA.t910 GNDA 0.057959f
C3965 VDDA.n1071 GNDA 0.025357f
C3966 VDDA.t840 GNDA 0.057959f
C3967 VDDA.n1072 GNDA 0.025357f
C3968 VDDA.t442 GNDA 0.057959f
C3969 VDDA.n1073 GNDA 0.025357f
C3970 VDDA.t903 GNDA 0.057959f
C3971 VDDA.n1074 GNDA 0.025357f
C3972 VDDA.t501 GNDA 0.057959f
C3973 VDDA.n1075 GNDA 0.025357f
C3974 VDDA.n1076 GNDA 0.047092f
C3975 VDDA.t433 GNDA 0.058946f
C3976 VDDA.t513 GNDA 0.057959f
C3977 VDDA.n1077 GNDA 0.03886f
C3978 VDDA.t915 GNDA 0.057959f
C3979 VDDA.n1078 GNDA 0.025357f
C3980 VDDA.t768 GNDA 0.057959f
C3981 VDDA.n1079 GNDA 0.025357f
C3982 VDDA.t854 GNDA 0.057959f
C3983 VDDA.n1080 GNDA 0.025357f
C3984 VDDA.t705 GNDA 0.057959f
C3985 VDDA.n1081 GNDA 0.025357f
C3986 VDDA.t558 GNDA 0.057959f
C3987 VDDA.n1082 GNDA 0.025357f
C3988 VDDA.t642 GNDA 0.057959f
C3989 VDDA.n1083 GNDA 0.025357f
C3990 VDDA.t493 GNDA 0.057959f
C3991 VDDA.t549 GNDA 0.058946f
C3992 VDDA.t693 GNDA 0.057959f
C3993 VDDA.n1084 GNDA 0.03886f
C3994 VDDA.t843 GNDA 0.057959f
C3995 VDDA.n1085 GNDA 0.025357f
C3996 VDDA.t755 GNDA 0.057959f
C3997 VDDA.n1086 GNDA 0.025357f
C3998 VDDA.t682 GNDA 0.057959f
C3999 VDDA.n1087 GNDA 0.025357f
C4000 VDDA.t831 GNDA 0.057959f
C4001 VDDA.n1088 GNDA 0.025357f
C4002 VDDA.t745 GNDA 0.057959f
C4003 VDDA.n1089 GNDA 0.025357f
C4004 VDDA.t895 GNDA 0.057959f
C4005 VDDA.n1090 GNDA 0.025357f
C4006 VDDA.n1091 GNDA 0.047092f
C4007 VDDA.t822 GNDA 0.058946f
C4008 VDDA.t907 GNDA 0.057959f
C4009 VDDA.n1092 GNDA 0.03886f
C4010 VDDA.t759 GNDA 0.057959f
C4011 VDDA.n1093 GNDA 0.025357f
C4012 VDDA.t612 GNDA 0.057959f
C4013 VDDA.n1094 GNDA 0.025357f
C4014 VDDA.t696 GNDA 0.057959f
C4015 VDDA.n1095 GNDA 0.025357f
C4016 VDDA.t550 GNDA 0.057959f
C4017 VDDA.n1096 GNDA 0.025357f
C4018 VDDA.t953 GNDA 0.057959f
C4019 VDDA.n1097 GNDA 0.025357f
C4020 VDDA.t486 GNDA 0.057959f
C4021 VDDA.n1098 GNDA 0.025357f
C4022 VDDA.t886 GNDA 0.057959f
C4023 VDDA.t942 GNDA 0.058946f
C4024 VDDA.t539 GNDA 0.057959f
C4025 VDDA.n1099 GNDA 0.03886f
C4026 VDDA.t687 GNDA 0.057959f
C4027 VDDA.n1100 GNDA 0.025357f
C4028 VDDA.t600 GNDA 0.057959f
C4029 VDDA.n1101 GNDA 0.025357f
C4030 VDDA.t527 GNDA 0.057959f
C4031 VDDA.n1102 GNDA 0.025357f
C4032 VDDA.t672 GNDA 0.057959f
C4033 VDDA.n1103 GNDA 0.025357f
C4034 VDDA.t589 GNDA 0.057959f
C4035 VDDA.n1104 GNDA 0.025357f
C4036 VDDA.t737 GNDA 0.057959f
C4037 VDDA.n1105 GNDA 0.025357f
C4038 VDDA.n1106 GNDA 0.047092f
C4039 VDDA.t961 GNDA 0.058946f
C4040 VDDA.t495 GNDA 0.057959f
C4041 VDDA.n1107 GNDA 0.03886f
C4042 VDDA.t897 GNDA 0.057959f
C4043 VDDA.n1108 GNDA 0.025357f
C4044 VDDA.t747 GNDA 0.057959f
C4045 VDDA.n1109 GNDA 0.025357f
C4046 VDDA.t833 GNDA 0.057959f
C4047 VDDA.n1110 GNDA 0.025357f
C4048 VDDA.t685 GNDA 0.057959f
C4049 VDDA.n1111 GNDA 0.025357f
C4050 VDDA.t538 GNDA 0.057959f
C4051 VDDA.n1112 GNDA 0.025357f
C4052 VDDA.t625 GNDA 0.057959f
C4053 VDDA.n1113 GNDA 0.025357f
C4054 VDDA.t475 GNDA 0.057959f
C4055 VDDA.t525 GNDA 0.058946f
C4056 VDDA.t671 GNDA 0.057959f
C4057 VDDA.n1114 GNDA 0.03886f
C4058 VDDA.t823 GNDA 0.057959f
C4059 VDDA.n1115 GNDA 0.025357f
C4060 VDDA.t734 GNDA 0.057959f
C4061 VDDA.n1116 GNDA 0.025357f
C4062 VDDA.t662 GNDA 0.057959f
C4063 VDDA.n1117 GNDA 0.025357f
C4064 VDDA.t812 GNDA 0.057959f
C4065 VDDA.n1118 GNDA 0.025357f
C4066 VDDA.t726 GNDA 0.057959f
C4067 VDDA.n1119 GNDA 0.025357f
C4068 VDDA.t876 GNDA 0.057959f
C4069 VDDA.n1120 GNDA 0.025357f
C4070 VDDA.n1121 GNDA 0.047092f
C4071 VDDA.t805 GNDA 0.058946f
C4072 VDDA.t889 GNDA 0.057959f
C4073 VDDA.n1122 GNDA 0.03886f
C4074 VDDA.t739 GNDA 0.057959f
C4075 VDDA.n1123 GNDA 0.025357f
C4076 VDDA.t592 GNDA 0.057959f
C4077 VDDA.n1124 GNDA 0.025357f
C4078 VDDA.t676 GNDA 0.057959f
C4079 VDDA.n1125 GNDA 0.025357f
C4080 VDDA.t531 GNDA 0.057959f
C4081 VDDA.n1126 GNDA 0.025357f
C4082 VDDA.t930 GNDA 0.057959f
C4083 VDDA.n1127 GNDA 0.025357f
C4084 VDDA.t470 GNDA 0.057959f
C4085 VDDA.n1128 GNDA 0.025357f
C4086 VDDA.t868 GNDA 0.057959f
C4087 VDDA.t918 GNDA 0.058946f
C4088 VDDA.t515 GNDA 0.057959f
C4089 VDDA.n1129 GNDA 0.03886f
C4090 VDDA.t665 GNDA 0.057959f
C4091 VDDA.n1130 GNDA 0.025357f
C4092 VDDA.t579 GNDA 0.057959f
C4093 VDDA.n1131 GNDA 0.025357f
C4094 VDDA.t504 GNDA 0.057959f
C4095 VDDA.n1132 GNDA 0.025357f
C4096 VDDA.t654 GNDA 0.057959f
C4097 VDDA.n1133 GNDA 0.025357f
C4098 VDDA.t570 GNDA 0.057959f
C4099 VDDA.n1134 GNDA 0.025357f
C4100 VDDA.t717 GNDA 0.057959f
C4101 VDDA.n1135 GNDA 0.025357f
C4102 VDDA.n1136 GNDA 0.047092f
C4103 VDDA.t646 GNDA 0.058946f
C4104 VDDA.t731 GNDA 0.057959f
C4105 VDDA.n1137 GNDA 0.03886f
C4106 VDDA.t584 GNDA 0.057959f
C4107 VDDA.n1138 GNDA 0.025357f
C4108 VDDA.t437 GNDA 0.057959f
C4109 VDDA.n1139 GNDA 0.025357f
C4110 VDDA.t518 GNDA 0.057959f
C4111 VDDA.n1140 GNDA 0.025357f
C4112 VDDA.t921 GNDA 0.057959f
C4113 VDDA.n1141 GNDA 0.025357f
C4114 VDDA.t774 GNDA 0.057959f
C4115 VDDA.n1142 GNDA 0.025357f
C4116 VDDA.t860 GNDA 0.057959f
C4117 VDDA.n1143 GNDA 0.025357f
C4118 VDDA.t710 GNDA 0.057959f
C4119 VDDA.t762 GNDA 0.058946f
C4120 VDDA.t908 GNDA 0.057959f
C4121 VDDA.n1144 GNDA 0.03886f
C4122 VDDA.t508 GNDA 0.057959f
C4123 VDDA.n1145 GNDA 0.025357f
C4124 VDDA.t425 GNDA 0.057959f
C4125 VDDA.n1146 GNDA 0.025357f
C4126 VDDA.t898 GNDA 0.057959f
C4127 VDDA.n1147 GNDA 0.025357f
C4128 VDDA.t498 GNDA 0.057959f
C4129 VDDA.n1148 GNDA 0.025357f
C4130 VDDA.t964 GNDA 0.057959f
C4131 VDDA.n1149 GNDA 0.025357f
C4132 VDDA.t562 GNDA 0.057959f
C4133 VDDA.n1150 GNDA 0.025357f
C4134 VDDA.n1151 GNDA 0.047092f
C4135 VDDA.t490 GNDA 0.058946f
C4136 VDDA.t574 GNDA 0.057959f
C4137 VDDA.n1152 GNDA 0.03886f
C4138 VDDA.t430 GNDA 0.057959f
C4139 VDDA.n1153 GNDA 0.025357f
C4140 VDDA.t827 GNDA 0.057959f
C4141 VDDA.n1154 GNDA 0.025357f
C4142 VDDA.t911 GNDA 0.057959f
C4143 VDDA.n1155 GNDA 0.025357f
C4144 VDDA.t766 GNDA 0.057959f
C4145 VDDA.n1156 GNDA 0.025357f
C4146 VDDA.t618 GNDA 0.057959f
C4147 VDDA.n1157 GNDA 0.025357f
C4148 VDDA.t702 GNDA 0.057959f
C4149 VDDA.n1158 GNDA 0.025357f
C4150 VDDA.t557 GNDA 0.057959f
C4151 VDDA.n1159 GNDA 0.036224f
C4152 VDDA.t957 GNDA 0.057959f
C4153 VDDA.n1160 GNDA 0.025357f
C4154 VDDA.t808 GNDA 0.057959f
C4155 VDDA.n1161 GNDA 0.025357f
C4156 VDDA.t894 GNDA 0.057959f
C4157 VDDA.n1162 GNDA 0.025357f
C4158 VDDA.t742 GNDA 0.057959f
C4159 VDDA.n1163 GNDA 0.025357f
C4160 VDDA.t817 GNDA 0.057959f
C4161 VDDA.n1164 GNDA 0.025357f
C4162 VDDA.t904 GNDA 0.057959f
C4163 VDDA.n1165 GNDA 0.025357f
C4164 VDDA.t754 GNDA 0.057959f
C4165 VDDA.n1166 GNDA 0.025357f
C4166 VDDA.t607 GNDA 0.057959f
C4167 VDDA.n1167 GNDA 0.020771f
C4168 VDDA.n1193 GNDA 0.010867f
C4169 VDDA.n1195 GNDA 0.012171f
C4170 VDDA.n1197 GNDA 0.011737f
C4171 VDDA.n1199 GNDA 0.010867f
C4172 VDDA.n1201 GNDA 0.012171f
C4173 VDDA.n1203 GNDA 0.011737f
C4174 VDDA.n1205 GNDA 0.010867f
C4175 VDDA.n1207 GNDA 0.012171f
C4176 VDDA.n1209 GNDA 0.011737f
C4177 VDDA.n1211 GNDA 0.010867f
C4178 VDDA.n1213 GNDA 0.033905f
C4179 VDDA.n1221 GNDA 0.012171f
C4180 VDDA.n1222 GNDA 0.011737f
C4181 VDDA.n1223 GNDA 0.010867f
C4182 VDDA.n1231 GNDA 0.011737f
C4183 VDDA.n1232 GNDA 0.012171f
C4184 VDDA.n1233 GNDA 0.012171f
C4185 VDDA.n1241 GNDA 0.010867f
C4186 VDDA.n1242 GNDA 0.010867f
C4187 VDDA.n1243 GNDA 0.011737f
C4188 VDDA.n1251 GNDA 0.012171f
C4189 VDDA.n1252 GNDA 0.011737f
C4190 VDDA.n1253 GNDA 0.010867f
C4191 VDDA.n1261 GNDA 0.011737f
C4192 VDDA.n1262 GNDA 0.012171f
C4193 VDDA.n1263 GNDA 0.012171f
C4194 VDDA.n1271 GNDA 0.010867f
C4195 VDDA.n1272 GNDA 0.010867f
C4196 VDDA.n1273 GNDA 0.011737f
C4197 VDDA.n1281 GNDA 0.012171f
C4198 VDDA.n1282 GNDA 0.011737f
C4199 VDDA.n1283 GNDA 0.010867f
C4200 VDDA.n1291 GNDA 0.011737f
C4201 VDDA.n1292 GNDA 0.012171f
C4202 VDDA.n1293 GNDA 0.012171f
C4203 VDDA.n1301 GNDA 0.010867f
C4204 VDDA.n1302 GNDA 0.010867f
C4205 VDDA.n1303 GNDA 0.011737f
C4206 VDDA.n1311 GNDA 0.012171f
C4207 VDDA.n1312 GNDA 0.011737f
C4208 VDDA.n1313 GNDA 0.010867f
C4209 VDDA.n1321 GNDA 0.011737f
C4210 VDDA.n1322 GNDA 0.012171f
C4211 VDDA.n1323 GNDA 0.012171f
C4212 VDDA.n1327 GNDA 1.09639f
C4213 VDDA.n1330 GNDA 0.290123f
C4214 VDDA.n1331 GNDA 0.011737f
C4215 VDDA.n1335 GNDA 0.010867f
C4216 VDDA.n1339 GNDA 0.012171f
C4217 VDDA.n1343 GNDA 0.011737f
C4218 VDDA.n1347 GNDA 0.010867f
C4219 VDDA.n1351 GNDA 0.012171f
C4220 VDDA.n1355 GNDA 0.011737f
C4221 VDDA.n1359 GNDA 0.010867f
C4222 VDDA.n1363 GNDA 0.012171f
C4223 VDDA.n1367 GNDA 0.011737f
C4224 VDDA.n1371 GNDA 0.010867f
C4225 VDDA.n1375 GNDA 0.033905f
C4226 VDDA.n1386 GNDA 0.012171f
C4227 VDDA.n1387 GNDA 0.011737f
C4228 VDDA.n1388 GNDA 0.010867f
C4229 VDDA.n1396 GNDA 0.011737f
C4230 VDDA.n1397 GNDA 0.012171f
C4231 VDDA.n1398 GNDA 0.012171f
C4232 VDDA.n1406 GNDA 0.010867f
C4233 VDDA.n1407 GNDA 0.010867f
C4234 VDDA.n1408 GNDA 0.011737f
C4235 VDDA.n1416 GNDA 0.012171f
C4236 VDDA.n1417 GNDA 0.011737f
C4237 VDDA.n1418 GNDA 0.010867f
C4238 VDDA.n1426 GNDA 0.011737f
C4239 VDDA.n1427 GNDA 0.012171f
C4240 VDDA.n1428 GNDA 0.012171f
C4241 VDDA.n1436 GNDA 0.010867f
C4242 VDDA.n1437 GNDA 0.010867f
C4243 VDDA.n1438 GNDA 0.011737f
C4244 VDDA.n1446 GNDA 0.012171f
C4245 VDDA.n1447 GNDA 0.011737f
C4246 VDDA.n1448 GNDA 0.010867f
C4247 VDDA.n1456 GNDA 0.011737f
C4248 VDDA.n1457 GNDA 0.012171f
C4249 VDDA.n1458 GNDA 0.012171f
C4250 VDDA.n1466 GNDA 0.010867f
C4251 VDDA.n1467 GNDA 0.010867f
C4252 VDDA.n1468 GNDA 0.011737f
C4253 VDDA.n1476 GNDA 0.012171f
C4254 VDDA.n1477 GNDA 0.011737f
C4255 VDDA.n1478 GNDA 0.010867f
C4256 VDDA.n1486 GNDA 0.011737f
C4257 VDDA.n1487 GNDA 0.012171f
C4258 VDDA.n1488 GNDA 0.012171f
C4259 VDDA.n1495 GNDA 0.26128f
C4260 VDDA.n1496 GNDA 0.227568f
C4261 VDDA.n1497 GNDA 0.14168f
C4262 VDDA.n1498 GNDA 0.26128f
C4263 VDDA.n1501 GNDA 2.43427f
C4264 VDDA.n1528 GNDA 0.012171f
C4265 VDDA.n1532 GNDA 0.011737f
C4266 VDDA.n1536 GNDA 0.010867f
C4267 VDDA.n1540 GNDA 0.012171f
C4268 VDDA.n1544 GNDA 0.011737f
C4269 VDDA.n1548 GNDA 0.010867f
C4270 VDDA.n1552 GNDA 0.012171f
C4271 VDDA.n1556 GNDA 0.011737f
C4272 VDDA.n1560 GNDA 0.010867f
C4273 VDDA.n1564 GNDA 0.012171f
C4274 VDDA.n1568 GNDA 0.011737f
C4275 VDDA.n1575 GNDA 0.033905f
C4276 VDDA.n1576 GNDA 0.012171f
C4277 VDDA.n1582 GNDA 0.010867f
C4278 VDDA.n1583 GNDA 0.010867f
C4279 VDDA.n1584 GNDA 0.011737f
C4280 VDDA.n1590 GNDA 0.012171f
C4281 VDDA.n1591 GNDA 0.011737f
C4282 VDDA.n1592 GNDA 0.010867f
C4283 VDDA.n1598 GNDA 0.011737f
C4284 VDDA.n1599 GNDA 0.012171f
C4285 VDDA.n1600 GNDA 0.012171f
C4286 VDDA.n1606 GNDA 0.010867f
C4287 VDDA.n1607 GNDA 0.010867f
C4288 VDDA.n1608 GNDA 0.011737f
C4289 VDDA.n1614 GNDA 0.012171f
C4290 VDDA.n1615 GNDA 0.011737f
C4291 VDDA.n1616 GNDA 0.010867f
C4292 VDDA.n1622 GNDA 0.011737f
C4293 VDDA.n1623 GNDA 0.012171f
C4294 VDDA.n1624 GNDA 0.012171f
C4295 VDDA.n1630 GNDA 0.010867f
C4296 VDDA.n1631 GNDA 0.010867f
C4297 VDDA.n1632 GNDA 0.011737f
C4298 VDDA.n1638 GNDA 0.012171f
C4299 VDDA.n1639 GNDA 0.011737f
C4300 VDDA.n1640 GNDA 0.010867f
C4301 VDDA.n1646 GNDA 0.011737f
C4302 VDDA.n1647 GNDA 0.012171f
C4303 VDDA.n1648 GNDA 0.012171f
C4304 VDDA.n1654 GNDA 0.010867f
C4305 VDDA.n1655 GNDA 0.010867f
C4306 VDDA.n1656 GNDA 0.011737f
C4307 VDDA.n1662 GNDA 0.012171f
C4308 VDDA.n1663 GNDA 0.011737f
C4309 VDDA.n1664 GNDA 0.26128f
C4310 VDDA.n1667 GNDA 2.43427f
C4311 VDDA.n1693 GNDA 0.010867f
C4312 VDDA.n1697 GNDA 0.012171f
C4313 VDDA.n1701 GNDA 0.011737f
C4314 VDDA.n1705 GNDA 0.010867f
C4315 VDDA.n1709 GNDA 0.012171f
C4316 VDDA.n1713 GNDA 0.011737f
C4317 VDDA.n1717 GNDA 0.010867f
C4318 VDDA.n1721 GNDA 0.012171f
C4319 VDDA.n1725 GNDA 0.011737f
C4320 VDDA.n1729 GNDA 0.010867f
C4321 VDDA.n1733 GNDA 0.033905f
C4322 VDDA.n1741 GNDA 0.012171f
C4323 VDDA.n1742 GNDA 0.011737f
C4324 VDDA.n1743 GNDA 0.010867f
C4325 VDDA.n1749 GNDA 0.011737f
C4326 VDDA.n1750 GNDA 0.012171f
C4327 VDDA.n1751 GNDA 0.012171f
C4328 VDDA.n1757 GNDA 0.010867f
C4329 VDDA.n1758 GNDA 0.010867f
C4330 VDDA.n1759 GNDA 0.011737f
C4331 VDDA.n1765 GNDA 0.012171f
C4332 VDDA.n1766 GNDA 0.011737f
C4333 VDDA.n1767 GNDA 0.010867f
C4334 VDDA.n1773 GNDA 0.011737f
C4335 VDDA.n1774 GNDA 0.012171f
C4336 VDDA.n1775 GNDA 0.012171f
C4337 VDDA.n1781 GNDA 0.010867f
C4338 VDDA.n1782 GNDA 0.010867f
C4339 VDDA.n1783 GNDA 0.011737f
C4340 VDDA.n1789 GNDA 0.012171f
C4341 VDDA.n1790 GNDA 0.011737f
C4342 VDDA.n1791 GNDA 0.010867f
C4343 VDDA.n1797 GNDA 0.011737f
C4344 VDDA.n1798 GNDA 0.012171f
C4345 VDDA.n1799 GNDA 0.012171f
C4346 VDDA.n1805 GNDA 0.010867f
C4347 VDDA.n1806 GNDA 0.010867f
C4348 VDDA.n1807 GNDA 0.011737f
C4349 VDDA.n1813 GNDA 0.012171f
C4350 VDDA.n1814 GNDA 0.011737f
C4351 VDDA.n1815 GNDA 0.010867f
C4352 VDDA.n1821 GNDA 0.011737f
C4353 VDDA.n1822 GNDA 0.012171f
C4354 VDDA.n1823 GNDA 0.012171f
C4355 VDDA.n1947 GNDA 0.014166f
C4356 VDDA.n1948 GNDA 0.061035f
C4357 VDDA.t261 GNDA 0.020728f
C4358 VDDA.n1961 GNDA 0.02539f
C4359 VDDA.t317 GNDA 0.017582f
C4360 VDDA.t163 GNDA 0.011157f
C4361 VDDA.t164 GNDA 0.011157f
C4362 VDDA.t354 GNDA 0.017969f
C4363 VDDA.n1962 GNDA 0.026592f
C4364 VDDA.n1964 GNDA 0.115084f
C4365 VDDA.n1965 GNDA 0.014166f
C4366 VDDA.n1966 GNDA 0.014166f
C4367 VDDA.n1967 GNDA 0.014166f
C4368 VDDA.n1968 GNDA 0.014166f
C4369 VDDA.n1969 GNDA 0.014166f
C4370 VDDA.n1970 GNDA 0.014166f
C4371 VDDA.n1971 GNDA 0.014166f
C4372 VDDA.n1972 GNDA 0.061035f
C4373 VDDA.n1973 GNDA 0.061035f
C4374 VDDA.n1974 GNDA 0.061035f
C4375 VDDA.n1975 GNDA 0.061035f
C4376 VDDA.n1976 GNDA 0.061035f
C4377 VDDA.n1977 GNDA 0.061035f
C4378 VDDA.n1978 GNDA 0.061035f
C4379 VDDA.n1979 GNDA 0.065661f
C4380 VDDA.n1989 GNDA 0.040644f
C4381 VDDA.t262 GNDA 0.043107f
C4382 VDDA.t61 GNDA 0.044339f
C4383 VDDA.t10 GNDA 0.044339f
C4384 VDDA.t116 GNDA 0.044339f
C4385 VDDA.t215 GNDA 0.044339f
C4386 VDDA.t211 GNDA 0.044339f
C4387 VDDA.t108 GNDA 0.044339f
C4388 VDDA.t100 GNDA 0.044339f
C4389 VDDA.t98 GNDA 0.044339f
C4390 VDDA.t183 GNDA 0.044339f
C4391 VDDA.t59 GNDA 0.044339f
C4392 VDDA.t193 GNDA 0.044339f
C4393 VDDA.t64 GNDA 0.044339f
C4394 VDDA.t103 GNDA 0.044339f
C4395 VDDA.t113 GNDA 0.044339f
C4396 VDDA.t188 GNDA 0.044339f
C4397 VDDA.t165 GNDA 0.044339f
C4398 VDDA.t348 GNDA 0.043107f
C4399 VDDA.n2002 GNDA 0.040644f
C4400 VDDA.t347 GNDA 0.020728f
C4401 VDDA.n2006 GNDA 0.065661f
C4402 VDDA.n2007 GNDA 0.057547f
C4403 VDDA.n2021 GNDA 0.025647f
C4404 VDDA.t308 GNDA 0.0213f
C4405 VDDA.t78 GNDA 0.019126f
C4406 VDDA.t344 GNDA 0.0213f
C4407 VDDA.n2027 GNDA 0.025647f
C4408 VDDA.n2031 GNDA 0.039491f
C4409 VDDA.n2033 GNDA 0.042211f
C4410 VDDA.n2034 GNDA 0.033089f
C4411 VDDA.n2148 GNDA 0.016551f
C4412 VDDA.n2151 GNDA 7.557839f
C4413 VDDA.n2177 GNDA 0.02525f
C4414 VDDA.t268 GNDA 0.017581f
C4415 VDDA.t76 GNDA 0.011157f
C4416 VDDA.t84 GNDA 0.011157f
C4417 VDDA.t351 GNDA 0.017581f
C4418 VDDA.n2178 GNDA 0.02525f
C4419 VDDA.n2181 GNDA 0.053652f
C4420 VDDA.n2185 GNDA 0.015083f
C4421 VDDA.t293 GNDA 0.015895f
C4422 VDDA.t88 GNDA 0.011157f
C4423 VDDA.t376 GNDA 0.011157f
C4424 VDDA.t45 GNDA 0.011157f
C4425 VDDA.t30 GNDA 0.011157f
C4426 VDDA.t256 GNDA 0.015895f
C4427 VDDA.n2186 GNDA 0.015083f
C4428 VDDA.n2194 GNDA 0.02525f
C4429 VDDA.t329 GNDA 0.017581f
C4430 VDDA.t51 GNDA 0.011157f
C4431 VDDA.t374 GNDA 0.011157f
C4432 VDDA.t43 GNDA 0.011157f
C4433 VDDA.t86 GNDA 0.011157f
C4434 VDDA.t80 GNDA 0.011157f
C4435 VDDA.t82 GNDA 0.011157f
C4436 VDDA.t47 GNDA 0.011157f
C4437 VDDA.t32 GNDA 0.011157f
C4438 VDDA.t363 GNDA 0.017581f
C4439 VDDA.n2195 GNDA 0.02525f
C4440 VDDA.n2200 GNDA 0.015086f
C4441 VDDA.t299 GNDA 0.015895f
C4442 VDDA.t122 GNDA 0.011157f
C4443 VDDA.t14 GNDA 0.011157f
C4444 VDDA.t49 GNDA 0.011157f
C4445 VDDA.t124 GNDA 0.011157f
C4446 VDDA.t332 GNDA 0.015895f
C4447 VDDA.n2201 GNDA 0.015086f
C4448 VDDA.n2203 GNDA 0.051064f
C4449 VDDA.n2204 GNDA 0.032227f
C4450 VDDA.n2205 GNDA 0.039901f
C4451 VDDA.n2206 GNDA 0.035988f
C4452 VDDA.n2207 GNDA 0.028323f
C4453 VDDA.n2208 GNDA 0.032235f
C4454 VDDA.n2209 GNDA 0.032235f
C4455 VDDA.n2210 GNDA 0.032235f
C4456 VDDA.n2211 GNDA 0.028323f
C4457 VDDA.n2212 GNDA 0.035988f
C4458 VDDA.n2213 GNDA 0.039901f
C4459 VDDA.n2214 GNDA 0.032226f
C4460 VDDA.n2215 GNDA 0.032226f
C4461 VDDA.n2216 GNDA 0.039901f
C4462 VDDA.n2217 GNDA 0.034775f
C4463 VDDA.n2218 GNDA 0.01937f
C4464 VDDA.n2219 GNDA 0.02022f
C4465 VDDA.n2333 GNDA 0.016551f
C4466 VDDA.n2336 GNDA 7.10576f
C4467 VDDA.n2362 GNDA 0.035547f
C4468 VDDA.n2365 GNDA 0.035547f
C4469 VDDA.n2367 GNDA 0.035547f
C4470 VDDA.n2369 GNDA 0.035547f
C4471 VDDA.n2371 GNDA 0.035547f
C4472 VDDA.n2373 GNDA 0.035547f
C4473 VDDA.n2375 GNDA 0.035547f
C4474 VDDA.n2377 GNDA 0.035547f
C4475 VDDA.n2379 GNDA 0.035547f
C4476 VDDA.n2381 GNDA 0.035547f
C4477 VDDA.n2385 GNDA 0.035547f
C4478 VDDA.n2387 GNDA 0.035547f
C4479 VDDA.n2389 GNDA 0.035547f
C4480 VDDA.n2391 GNDA 0.035547f
C4481 VDDA.n2393 GNDA 0.035547f
C4482 VDDA.n2395 GNDA 0.035547f
C4483 VDDA.n2397 GNDA 0.035547f
C4484 VDDA.n2399 GNDA 0.057235f
C4485 VDDA.n2403 GNDA 0.017861f
C4486 VDDA.t284 GNDA 0.015037f
C4487 VDDA.t404 GNDA 0.012171f
C4488 VDDA.t153 GNDA 0.012171f
C4489 VDDA.t136 GNDA 0.012171f
C4490 VDDA.t128 GNDA 0.012171f
C4491 VDDA.t41 GNDA 0.012171f
C4492 VDDA.t139 GNDA 0.012171f
C4493 VDDA.t202 GNDA 0.012171f
C4494 VDDA.t141 GNDA 0.012171f
C4495 VDDA.t91 GNDA 0.012171f
C4496 VDDA.t410 GNDA 0.012171f
C4497 VDDA.t38 GNDA 0.012171f
C4498 VDDA.t402 GNDA 0.012171f
C4499 VDDA.t16 GNDA 0.012171f
C4500 VDDA.t169 GNDA 0.012171f
C4501 VDDA.t93 GNDA 0.012171f
C4502 VDDA.t126 GNDA 0.012171f
C4503 VDDA.t412 GNDA 0.012171f
C4504 VDDA.t387 GNDA 0.012171f
C4505 VDDA.t305 GNDA 0.018213f
C4506 VDDA.n2404 GNDA 0.014685f
C4507 VDDA.n2407 GNDA 0.046275f
C4508 VDDA.n2408 GNDA 0.046275f
C4509 VDDA.n2410 GNDA 0.026435f
C4510 VDDA.t290 GNDA 0.018566f
C4511 VDDA.t415 GNDA 0.012171f
C4512 VDDA.t224 GNDA 0.012171f
C4513 VDDA.t222 GNDA 0.012171f
C4514 VDDA.t394 GNDA 0.012171f
C4515 VDDA.t19 GNDA 0.012171f
C4516 VDDA.t366 GNDA 0.012171f
C4517 VDDA.t419 GNDA 0.012171f
C4518 VDDA.t71 GNDA 0.012171f
C4519 VDDA.t149 GNDA 0.012171f
C4520 VDDA.t130 GNDA 0.012171f
C4521 VDDA.t147 GNDA 0.012171f
C4522 VDDA.t368 GNDA 0.012171f
C4523 VDDA.t417 GNDA 0.012171f
C4524 VDDA.t69 GNDA 0.012171f
C4525 VDDA.t385 GNDA 0.012171f
C4526 VDDA.t226 GNDA 0.012171f
C4527 VDDA.t151 GNDA 0.012171f
C4528 VDDA.t237 GNDA 0.012171f
C4529 VDDA.t250 GNDA 0.018213f
C4530 VDDA.n2411 GNDA 0.014685f
C4531 VDDA.n2414 GNDA 0.142184f
C4532 VDDA.n2415 GNDA 0.073548f
C4533 VDDA.n2529 GNDA 0.016551f
C4534 VDDA.n2532 GNDA 2.19085f
C4535 VDDA.t686 GNDA 0.16012f
C4536 VDDA.t844 GNDA 0.163012f
C4537 VDDA.t748 GNDA 0.170732f
C4538 VDDA.n2557 GNDA 0.143492f
C4539 VDDA.t673 GNDA 0.170665f
C4540 VDDA.n2558 GNDA 0.071512f
C4541 VDDA.n2559 GNDA 0.12884f
C4542 VDDA.n2560 GNDA 0.131316f
C4543 VDDA.n2674 GNDA 0.016551f
C4544 VDDA.n2677 GNDA 1.43738f
C4545 VDDA.n2678 GNDA 1.57648f
C4546 VDDA.n2681 GNDA 0.26128f
C4547 VDDA.n2682 GNDA 0.146011f
C4548 VDDA.n2683 GNDA 0.010683f
C4549 VDDA.n2684 GNDA 0.012674f
C4550 VDDA.n2685 GNDA 0.0342f
C4551 VDDA.t361 GNDA 0.01804f
C4552 VDDA.n2686 GNDA 0.012674f
C4553 VDDA.n2687 GNDA 0.038083f
C4554 VDDA.n2688 GNDA 0.024789f
C4555 VDDA.n2689 GNDA 0.052332f
C4556 VDDA.t360 GNDA 0.043228f
C4557 VDDA.t231 GNDA 0.033906f
C4558 VDDA.t235 GNDA 0.033906f
C4559 VDDA.t207 GNDA 0.033906f
C4560 VDDA.t161 GNDA 0.033906f
C4561 VDDA.t55 GNDA 0.033906f
C4562 VDDA.t145 GNDA 0.033906f
C4563 VDDA.t134 GNDA 0.033906f
C4564 VDDA.t233 GNDA 0.033906f
C4565 VDDA.t389 GNDA 0.033906f
C4566 VDDA.t36 GNDA 0.033906f
C4567 VDDA.t314 GNDA 0.043793f
C4568 VDDA.t315 GNDA 0.01804f
C4569 VDDA.n2690 GNDA 0.054592f
C4570 VDDA.n2691 GNDA 0.024789f
C4571 VDDA.n2692 GNDA 0.012674f
C4572 VDDA.n2693 GNDA 0.038083f
C4573 VDDA.n2694 GNDA 0.012674f
C4574 VDDA.n2695 GNDA 0.0342f
C4575 VDDA.n2697 GNDA 0.043807f
C4576 VDDA.n2698 GNDA 0.039053f
C4577 VDDA.n2699 GNDA 0.014947f
C4578 VDDA.n2700 GNDA 0.014436f
C4579 VDDA.n2701 GNDA 0.055527f
C4580 VDDA.n2702 GNDA 0.014436f
C4581 VDDA.n2703 GNDA 0.028526f
C4582 VDDA.n2704 GNDA 0.014436f
C4583 VDDA.n2705 GNDA 0.028526f
C4584 VDDA.n2706 GNDA 0.014436f
C4585 VDDA.n2707 GNDA 0.028526f
C4586 VDDA.n2708 GNDA 0.014436f
C4587 VDDA.n2709 GNDA 0.043911f
C4588 VDDA.n2710 GNDA 0.022132f
C4589 VDDA.t312 GNDA 0.010339f
C4590 VDDA.n2711 GNDA 0.031762f
C4591 VDDA.t311 GNDA 0.025757f
C4592 VDDA.t373 GNDA 0.019126f
C4593 VDDA.t168 GNDA 0.019126f
C4594 VDDA.t155 GNDA 0.019126f
C4595 VDDA.t90 GNDA 0.019126f
C4596 VDDA.t177 GNDA 0.019126f
C4597 VDDA.t396 GNDA 0.019126f
C4598 VDDA.t0 GNDA 0.019126f
C4599 VDDA.t63 GNDA 0.019126f
C4600 VDDA.t230 GNDA 0.019126f
C4601 VDDA.t40 GNDA 0.019126f
C4602 VDDA.t253 GNDA 0.025757f
C4603 VDDA.t254 GNDA 0.010339f
C4604 VDDA.n2712 GNDA 0.031762f
C4605 VDDA.n2713 GNDA 0.016903f
C4606 VDDA.n2714 GNDA 0.025074f
C4607 VDDA.n2715 GNDA 0.040618f
C4608 VDDA.n2716 GNDA 0.025902f
C4609 VDDA.n2717 GNDA 0.05314f
C4610 VDDA.t336 GNDA 0.030596f
C4611 VDDA.n2718 GNDA 0.025902f
C4612 VDDA.n2719 GNDA 0.05314f
C4613 VDDA.n2720 GNDA 0.025902f
C4614 VDDA.n2721 GNDA 0.05314f
C4615 VDDA.n2722 GNDA 0.025902f
C4616 VDDA.n2723 GNDA 0.05314f
C4617 VDDA.n2724 GNDA 0.025902f
C4618 VDDA.n2725 GNDA 0.056256f
C4619 VDDA.t334 GNDA 0.010548f
C4620 VDDA.n2726 GNDA 0.024087f
C4621 VDDA.n2727 GNDA 0.102346f
C4622 VDDA.t335 GNDA 0.066286f
C4623 VDDA.t120 GNDA 0.051004f
C4624 VDDA.t217 GNDA 0.050681f
C4625 VDDA.t95 GNDA 0.050312f
C4626 VDDA.t381 GNDA 0.051004f
C4627 VDDA.t219 GNDA 0.051004f
C4628 VDDA.t398 GNDA 0.051004f
C4629 VDDA.t191 GNDA 0.051004f
C4630 VDDA.t67 GNDA 0.051004f
C4631 VDDA.t186 GNDA 0.051004f
C4632 VDDA.t74 GNDA 0.051004f
C4633 VDDA.t274 GNDA 0.066286f
C4634 VDDA.t275 GNDA 0.030596f
C4635 VDDA.n2728 GNDA 0.102346f
C4636 VDDA.t273 GNDA 0.010548f
C4637 VDDA.n2729 GNDA 0.023718f
C4638 VDDA.n2731 GNDA 0.012491f
C4639 VDDA.n2732 GNDA 0.016152f
C4640 VDDA.n2733 GNDA 0.010867f
C4641 VDDA.t296 GNDA 0.025737f
C4642 VDDA.n2742 GNDA 0.010867f
C4643 VDDA.t221 GNDA 0.023111f
C4644 VDDA.t383 GNDA 0.023111f
C4645 VDDA.t157 GNDA 0.023111f
C4646 VDDA.t97 GNDA 0.023111f
C4647 VDDA.t302 GNDA 0.025737f
C4648 VDDA.n2753 GNDA 0.03099f
C4649 VDDA.n2757 GNDA 0.012491f
C4650 VDDA.n2758 GNDA 0.02151f
C4651 VDDA.n2769 GNDA 0.010867f
C4652 VDDA.n2772 GNDA 0.010867f
C4653 VDDA.n2775 GNDA 0.028364f
C4654 VDDA.t357 GNDA 0.025737f
C4655 VDDA.t18 GNDA 0.023111f
C4656 VDDA.t196 GNDA 0.023111f
C4657 VDDA.t400 GNDA 0.023111f
C4658 VDDA.t414 GNDA 0.023111f
C4659 VDDA.t326 GNDA 0.025737f
C4660 VDDA.n2782 GNDA 0.03099f
C4661 VDDA.n2786 GNDA 0.016293f
C4662 VDDA.n2787 GNDA 0.016084f
C4663 VDDA.n2788 GNDA 0.037065f
C4664 VDDA.n2789 GNDA 0.0548f
C4665 VDDA.n2790 GNDA 0.036388f
C4666 VDDA.n2791 GNDA 0.01274f
C4667 VDDA.t278 GNDA 0.023111f
C4668 VDDA.n2792 GNDA 0.018969f
C4669 VDDA.n2793 GNDA 0.0577f
C4670 VDDA.t277 GNDA 0.043228f
C4671 VDDA.t28 GNDA 0.033906f
C4672 VDDA.t320 GNDA 0.043228f
C4673 VDDA.t321 GNDA 0.01804f
C4674 VDDA.n2794 GNDA 0.0577f
C4675 VDDA.n2795 GNDA 0.018832f
C4676 VDDA.n2798 GNDA 0.023522f
C4677 VDDA.n2799 GNDA 0.01443f
C4678 VDDA.n2800 GNDA 0.028344f
C4679 VDDA.t280 GNDA 0.025234f
C4680 VDDA.t241 GNDA 0.019126f
C4681 VDDA.t265 GNDA 0.025234f
C4682 VDDA.n2801 GNDA 0.028344f
C4683 VDDA.n2802 GNDA 0.014293f
C4684 VDDA.n2804 GNDA 0.019742f
C4685 VDDA.n2805 GNDA 0.069063f
C4686 VDDA.n2806 GNDA 0.014947f
C4687 VDDA.n2807 GNDA 0.014436f
C4688 VDDA.n2808 GNDA 0.055527f
C4689 VDDA.n2809 GNDA 0.014436f
C4690 VDDA.n2810 GNDA 0.028526f
C4691 VDDA.n2811 GNDA 0.014436f
C4692 VDDA.n2812 GNDA 0.028526f
C4693 VDDA.n2813 GNDA 0.014436f
C4694 VDDA.n2814 GNDA 0.028526f
C4695 VDDA.n2815 GNDA 0.014436f
C4696 VDDA.n2816 GNDA 0.043911f
C4697 VDDA.n2817 GNDA 0.022132f
C4698 VDDA.t339 GNDA 0.010339f
C4699 VDDA.n2818 GNDA 0.031762f
C4700 VDDA.t338 GNDA 0.025757f
C4701 VDDA.t25 GNDA 0.019126f
C4702 VDDA.t180 GNDA 0.019126f
C4703 VDDA.t175 GNDA 0.019126f
C4704 VDDA.t181 GNDA 0.019126f
C4705 VDDA.t22 GNDA 0.019126f
C4706 VDDA.t198 GNDA 0.019126f
C4707 VDDA.t3 GNDA 0.019126f
C4708 VDDA.t206 GNDA 0.019126f
C4709 VDDA.t7 GNDA 0.019126f
C4710 VDDA.t200 GNDA 0.019126f
C4711 VDDA.t287 GNDA 0.025757f
C4712 VDDA.t288 GNDA 0.010339f
C4713 VDDA.n2819 GNDA 0.031762f
C4714 VDDA.n2820 GNDA 0.016903f
C4715 VDDA.n2821 GNDA 0.025074f
C4716 VDDA.n2822 GNDA 0.040618f
C4717 VDDA.n2823 GNDA 0.025902f
C4718 VDDA.n2824 GNDA 0.05314f
C4719 VDDA.t260 GNDA 0.030596f
C4720 VDDA.n2825 GNDA 0.025902f
C4721 VDDA.n2826 GNDA 0.05314f
C4722 VDDA.n2827 GNDA 0.025902f
C4723 VDDA.n2828 GNDA 0.05314f
C4724 VDDA.n2829 GNDA 0.025902f
C4725 VDDA.n2830 GNDA 0.05314f
C4726 VDDA.n2831 GNDA 0.025902f
C4727 VDDA.n2832 GNDA 0.056256f
C4728 VDDA.t258 GNDA 0.010548f
C4729 VDDA.n2833 GNDA 0.024087f
C4730 VDDA.n2834 GNDA 0.102346f
C4731 VDDA.t259 GNDA 0.066286f
C4732 VDDA.t1 GNDA 0.051004f
C4733 VDDA.t204 GNDA 0.051004f
C4734 VDDA.t172 GNDA 0.051004f
C4735 VDDA.t243 GNDA 0.051004f
C4736 VDDA.t247 GNDA 0.051004f
C4737 VDDA.t239 GNDA 0.051004f
C4738 VDDA.t245 GNDA 0.051004f
C4739 VDDA.t5 GNDA 0.051004f
C4740 VDDA.t178 GNDA 0.051004f
C4741 VDDA.t23 GNDA 0.051004f
C4742 VDDA.t323 GNDA 0.066286f
C4743 VDDA.t324 GNDA 0.030596f
C4744 VDDA.n2835 GNDA 0.102346f
C4745 VDDA.t322 GNDA 0.010548f
C4746 VDDA.n2836 GNDA 0.023718f
C4747 VDDA.n2837 GNDA 0.010803f
C4748 VDDA.n2838 GNDA 0.038442f
C4749 VDDA.n2839 GNDA 0.0548f
C4750 VDDA.n2840 GNDA 0.010683f
C4751 VDDA.n2841 GNDA 0.012674f
C4752 VDDA.n2842 GNDA 0.0342f
C4753 VDDA.t272 GNDA 0.01804f
C4754 VDDA.n2843 GNDA 0.012674f
C4755 VDDA.n2844 GNDA 0.038083f
C4756 VDDA.n2845 GNDA 0.024789f
C4757 VDDA.n2846 GNDA 0.054592f
C4758 VDDA.t271 GNDA 0.043793f
C4759 VDDA.t34 GNDA 0.033906f
C4760 VDDA.t406 GNDA 0.033906f
C4761 VDDA.t26 GNDA 0.033906f
C4762 VDDA.t132 GNDA 0.033906f
C4763 VDDA.t209 GNDA 0.033906f
C4764 VDDA.t408 GNDA 0.033906f
C4765 VDDA.t391 GNDA 0.033906f
C4766 VDDA.t159 GNDA 0.033906f
C4767 VDDA.t53 GNDA 0.033906f
C4768 VDDA.t143 GNDA 0.033906f
C4769 VDDA.t341 GNDA 0.043228f
C4770 VDDA.t342 GNDA 0.01804f
C4771 VDDA.n2847 GNDA 0.052332f
C4772 VDDA.n2848 GNDA 0.024789f
C4773 VDDA.n2849 GNDA 0.012674f
C4774 VDDA.n2850 GNDA 0.038083f
C4775 VDDA.n2851 GNDA 0.012674f
C4776 VDDA.n2852 GNDA 0.0342f
C4777 VDDA.n2854 GNDA 0.043807f
C4778 VDDA.n2855 GNDA 0.039057f
C4779 VDDA.n2856 GNDA 0.146014f
C4780 VDDA.n2857 GNDA 0.26128f
C4781 VDDA.n2860 GNDA 1.65763f
C4782 VDDA.n2887 GNDA 0.012171f
C4783 VDDA.n2891 GNDA 0.011737f
C4784 VDDA.n2895 GNDA 0.010867f
C4785 VDDA.n2899 GNDA 0.012171f
C4786 VDDA.n2903 GNDA 0.011737f
C4787 VDDA.n2907 GNDA 0.010867f
C4788 VDDA.n2911 GNDA 0.012171f
C4789 VDDA.n2915 GNDA 0.011737f
C4790 VDDA.n2919 GNDA 0.010867f
C4791 VDDA.n2923 GNDA 0.012171f
C4792 VDDA.n2927 GNDA 0.011737f
C4793 VDDA.n2934 GNDA 0.033905f
C4794 VDDA.n2935 GNDA 0.012171f
C4795 VDDA.n2941 GNDA 0.010867f
C4796 VDDA.n2942 GNDA 0.010867f
C4797 VDDA.n2943 GNDA 0.011737f
C4798 VDDA.n2949 GNDA 0.012171f
C4799 VDDA.n2950 GNDA 0.011737f
C4800 VDDA.n2951 GNDA 0.010867f
C4801 VDDA.n2957 GNDA 0.011737f
C4802 VDDA.n2958 GNDA 0.012171f
C4803 VDDA.n2959 GNDA 0.012171f
C4804 VDDA.n2965 GNDA 0.010867f
C4805 VDDA.n2966 GNDA 0.010867f
C4806 VDDA.n2967 GNDA 0.011737f
C4807 VDDA.n2973 GNDA 0.012171f
C4808 VDDA.n2974 GNDA 0.011737f
C4809 VDDA.n2975 GNDA 0.010867f
C4810 VDDA.n2981 GNDA 0.011737f
C4811 VDDA.n2982 GNDA 0.012171f
C4812 VDDA.n2983 GNDA 0.012171f
C4813 VDDA.n2989 GNDA 0.010867f
C4814 VDDA.n2990 GNDA 0.010867f
C4815 VDDA.n2991 GNDA 0.011737f
C4816 VDDA.n2997 GNDA 0.012171f
C4817 VDDA.n2998 GNDA 0.011737f
C4818 VDDA.n2999 GNDA 0.010867f
C4819 VDDA.n3005 GNDA 0.011737f
C4820 VDDA.n3006 GNDA 0.012171f
C4821 VDDA.n3007 GNDA 0.012171f
C4822 VDDA.n3013 GNDA 0.010867f
C4823 VDDA.n3014 GNDA 0.010867f
C4824 VDDA.n3015 GNDA 0.011737f
C4825 VDDA.n3021 GNDA 0.012171f
C4826 VDDA.n3022 GNDA 0.011737f
C4827 VDDA.n3023 GNDA 0.26128f
C4828 VDDA.n3026 GNDA 2.43427f
C4829 VDDA.n3052 GNDA 0.010867f
C4830 VDDA.n3056 GNDA 0.012171f
C4831 VDDA.n3060 GNDA 0.011737f
C4832 VDDA.n3064 GNDA 0.010867f
C4833 VDDA.n3068 GNDA 0.012171f
C4834 VDDA.n3072 GNDA 0.011737f
C4835 VDDA.n3076 GNDA 0.010867f
C4836 VDDA.n3080 GNDA 0.012171f
C4837 VDDA.n3084 GNDA 0.011737f
C4838 VDDA.n3088 GNDA 0.010867f
C4839 VDDA.n3092 GNDA 0.033905f
C4840 VDDA.n3100 GNDA 0.012171f
C4841 VDDA.n3101 GNDA 0.011737f
C4842 VDDA.n3102 GNDA 0.010867f
C4843 VDDA.n3108 GNDA 0.011737f
C4844 VDDA.n3109 GNDA 0.012171f
C4845 VDDA.n3110 GNDA 0.012171f
C4846 VDDA.n3116 GNDA 0.010867f
C4847 VDDA.n3117 GNDA 0.010867f
C4848 VDDA.n3118 GNDA 0.011737f
C4849 VDDA.n3124 GNDA 0.012171f
C4850 VDDA.n3125 GNDA 0.011737f
C4851 VDDA.n3126 GNDA 0.010867f
C4852 VDDA.n3132 GNDA 0.011737f
C4853 VDDA.n3133 GNDA 0.012171f
C4854 VDDA.n3134 GNDA 0.012171f
C4855 VDDA.n3140 GNDA 0.010867f
C4856 VDDA.n3141 GNDA 0.010867f
C4857 VDDA.n3142 GNDA 0.011737f
C4858 VDDA.n3148 GNDA 0.012171f
C4859 VDDA.n3149 GNDA 0.011737f
C4860 VDDA.n3150 GNDA 0.010867f
C4861 VDDA.n3156 GNDA 0.011737f
C4862 VDDA.n3157 GNDA 0.012171f
C4863 VDDA.n3158 GNDA 0.012171f
C4864 VDDA.n3164 GNDA 0.010867f
C4865 VDDA.n3165 GNDA 0.010867f
C4866 VDDA.n3166 GNDA 0.011737f
C4867 VDDA.n3172 GNDA 0.012171f
C4868 VDDA.n3173 GNDA 0.011737f
C4869 VDDA.n3174 GNDA 0.010867f
C4870 VDDA.n3180 GNDA 0.011737f
C4871 VDDA.n3181 GNDA 0.012171f
C4872 VDDA.n3182 GNDA 0.012171f
C4873 VDDA.n3186 GNDA 2.43427f
C4874 VDDA.n3189 GNDA 0.26128f
C4875 VDDA.n3190 GNDA 0.14168f
C4876 VDDA.n3191 GNDA 0.011737f
C4877 VDDA.n3195 GNDA 0.010867f
C4878 VDDA.n3199 GNDA 0.012171f
C4879 VDDA.n3203 GNDA 0.011737f
C4880 VDDA.n3207 GNDA 0.010867f
C4881 VDDA.n3211 GNDA 0.012171f
C4882 VDDA.n3215 GNDA 0.011737f
C4883 VDDA.n3219 GNDA 0.010867f
C4884 VDDA.n3223 GNDA 0.012171f
C4885 VDDA.n3227 GNDA 0.011737f
C4886 VDDA.n3231 GNDA 0.010867f
C4887 VDDA.n3235 GNDA 0.033905f
C4888 VDDA.n3246 GNDA 0.012171f
C4889 VDDA.n3247 GNDA 0.011737f
C4890 VDDA.n3248 GNDA 0.010867f
C4891 VDDA.n3256 GNDA 0.011737f
C4892 VDDA.n3257 GNDA 0.012171f
C4893 VDDA.n3258 GNDA 0.012171f
C4894 VDDA.n3266 GNDA 0.010867f
C4895 VDDA.n3267 GNDA 0.010867f
C4896 VDDA.n3268 GNDA 0.011737f
C4897 VDDA.n3276 GNDA 0.012171f
C4898 VDDA.n3277 GNDA 0.011737f
C4899 VDDA.n3278 GNDA 0.010867f
C4900 VDDA.n3286 GNDA 0.011737f
C4901 VDDA.n3287 GNDA 0.012171f
C4902 VDDA.n3288 GNDA 0.012171f
C4903 VDDA.n3296 GNDA 0.010867f
C4904 VDDA.n3297 GNDA 0.010867f
C4905 VDDA.n3298 GNDA 0.011737f
C4906 VDDA.n3306 GNDA 0.012171f
C4907 VDDA.n3307 GNDA 0.011737f
C4908 VDDA.n3308 GNDA 0.010867f
C4909 VDDA.n3316 GNDA 0.011737f
C4910 VDDA.n3317 GNDA 0.012171f
C4911 VDDA.n3318 GNDA 0.012171f
C4912 VDDA.n3326 GNDA 0.010867f
C4913 VDDA.n3327 GNDA 0.010867f
C4914 VDDA.n3328 GNDA 0.011737f
C4915 VDDA.n3336 GNDA 0.012171f
C4916 VDDA.n3337 GNDA 0.011737f
C4917 VDDA.n3338 GNDA 0.010867f
C4918 VDDA.n3346 GNDA 0.011737f
C4919 VDDA.n3347 GNDA 0.012171f
C4920 VDDA.n3348 GNDA 0.012171f
C4921 VDDA.n3355 GNDA 0.26128f
C4922 VDDA.n3356 GNDA 0.227567f
C4923 VDDA.n3357 GNDA 0.290119f
C4924 VDDA.n3360 GNDA 5.42495f
C4925 VDDA.n3361 GNDA 0.440488f
C4926 VDDA.n3362 GNDA 0.486855f
C4927 VDDA.n3363 GNDA 0.440488f
C4928 VDDA.n3364 GNDA 0.486855f
C4929 VDDA.n3365 GNDA 0.440488f
C4930 VDDA.n3366 GNDA 0.486855f
C4931 VDDA.n3367 GNDA 0.440488f
C4932 VDDA.n3368 GNDA 0.486855f
C4933 VDDA.n3369 GNDA 0.440488f
C4934 VDDA.n3370 GNDA 0.486855f
C4935 VDDA.n3371 GNDA 0.440488f
C4936 VDDA.n3372 GNDA 0.486855f
C4937 VDDA.n3373 GNDA 0.440488f
C4938 VDDA.n3374 GNDA 0.486855f
C4939 VDDA.n3375 GNDA 0.440488f
C4940 VDDA.n3376 GNDA 0.440488f
C4941 VDDA.n3378 GNDA 0.440488f
C4942 VDDA.n3381 GNDA 0.486855f
C4943 VDDA.n3384 GNDA 0.440488f
C4944 VDDA.n3387 GNDA 0.486855f
C4945 VDDA.n3390 GNDA 0.440488f
C4946 VDDA.n3393 GNDA 0.486855f
C4947 VDDA.n3396 GNDA 0.440488f
C4948 VDDA.n3399 GNDA 0.486855f
C4949 VDDA.n3402 GNDA 0.440488f
C4950 VDDA.n3405 GNDA 0.486855f
C4951 VDDA.n3408 GNDA 0.440488f
C4952 VDDA.n3411 GNDA 0.486855f
C4953 VDDA.n3414 GNDA 0.440488f
C4954 VDDA.n3417 GNDA 0.486855f
C4955 VDDA.n3420 GNDA 0.440488f
C4956 VDDA.n3423 GNDA 0.463671f
C4957 VDDA.n3424 GNDA 0.45208f
C4958 VDDA.n3425 GNDA 0.498447f
C4959 VDDA.n3426 GNDA 0.440488f
C4960 VDDA.n3427 GNDA 0.463671f
C4961 VDDA.n3428 GNDA 0.45208f
C4962 VDDA.n3429 GNDA 0.498447f
C4963 VDDA.n3430 GNDA 0.440488f
C4964 VDDA.n3431 GNDA 0.463671f
C4965 VDDA.n3432 GNDA 0.45208f
C4966 VDDA.n3433 GNDA 0.498447f
C4967 VDDA.n3434 GNDA 0.440488f
C4968 VDDA.n3435 GNDA 0.463671f
C4969 VDDA.n3436 GNDA 0.45208f
C4970 VDDA.n3437 GNDA 0.440488f
C4971 VDDA.n3440 GNDA 0.463671f
C4972 VDDA.n3442 GNDA 0.45208f
C4973 VDDA.n3444 GNDA 0.498447f
C4974 VDDA.n3446 GNDA 0.440488f
C4975 VDDA.n3448 GNDA 0.463671f
C4976 VDDA.n3450 GNDA 0.45208f
C4977 VDDA.n3452 GNDA 0.498447f
C4978 VDDA.n3454 GNDA 0.440488f
C4979 VDDA.n3456 GNDA 0.463671f
C4980 VDDA.n3458 GNDA 0.45208f
C4981 VDDA.n3460 GNDA 0.498447f
C4982 VDDA.n3462 GNDA 0.440488f
C4983 VDDA.n3464 GNDA 0.463671f
C4984 VDDA.n3465 GNDA 0.486855f
C4985 VDDA.n3466 GNDA 4.83377f
C4986 VDDA.n3467 GNDA 1.51852f
.ends

