magic
tech sky130A
timestamp 1740540882
<< poly >>
rect -130 960 -90 975
rect 2180 945 2220 955
rect 2180 930 2190 945
rect 2090 925 2190 930
rect 2210 925 2220 945
rect 2090 915 2220 925
rect 3090 680 3130 690
rect 3090 660 3100 680
rect 3120 660 3130 680
rect 3090 650 3130 660
rect 3850 680 3890 690
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 3850 650 3890 660
rect 4070 490 4110 500
rect 4070 470 4080 490
rect 4100 470 4110 490
rect 4070 460 4110 470
rect -130 260 -90 270
rect -130 240 -120 260
rect -100 240 -90 260
rect -130 230 -90 240
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
rect 6010 -310 6050 -300
rect 6010 -330 6020 -310
rect 6040 -330 6050 -310
rect 6010 -340 6050 -330
rect 4965 -600 4985 -585
<< polycont >>
rect 2190 925 2210 945
rect 3100 660 3120 680
rect 3860 660 3880 680
rect 4080 470 4100 490
rect -120 240 -100 260
rect 2085 65 2105 85
rect 6020 -330 6040 -310
<< locali >>
rect 2775 2815 2825 2830
rect 2775 2795 2790 2815
rect 2810 2795 2825 2815
rect 2775 2780 2825 2795
rect 4820 2540 4860 2550
rect 4820 2520 4830 2540
rect 4850 2520 4860 2540
rect 4820 2510 4860 2520
rect 2775 2220 2825 2235
rect 2775 2200 2790 2220
rect 2810 2200 2825 2220
rect 2775 2185 2825 2200
rect 2380 1220 2430 1230
rect 2380 1210 2390 1220
rect 2355 1190 2390 1210
rect 2420 1190 2430 1220
rect 2380 1180 2430 1190
rect 2040 1155 2080 1165
rect 2040 1135 2050 1155
rect 2070 1135 2080 1155
rect 2040 1125 2080 1135
rect 2040 1105 2060 1125
rect 2735 1015 2785 1030
rect 2735 995 2750 1015
rect 2770 995 2785 1015
rect 2735 980 2785 995
rect 2180 945 2220 955
rect 2180 925 2190 945
rect 2210 925 2220 945
rect 2180 915 2220 925
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 925 2340 945
rect 2300 915 2340 925
rect 3090 680 3130 690
rect 3090 660 3100 680
rect 3120 660 3130 680
rect 3850 680 3890 690
rect 3090 650 3130 660
rect 3155 645 3195 665
rect 3850 660 3860 680
rect 3880 660 3890 680
rect 3850 650 3890 660
rect -190 625 -140 635
rect -190 595 -180 625
rect -150 620 -140 625
rect 2460 625 2510 640
rect 2460 620 2475 625
rect -150 600 -130 620
rect 2370 600 2400 620
rect 2420 605 2475 620
rect 2495 605 2510 625
rect 3155 625 3165 645
rect 3185 625 3195 645
rect 3155 615 3195 625
rect 2420 600 2510 605
rect -150 595 -140 600
rect -190 585 -140 595
rect 2460 590 2510 600
rect 4450 595 4490 605
rect 4450 575 4460 595
rect 4480 575 4490 595
rect 4450 565 4490 575
rect 2040 550 2220 560
rect 2040 540 2190 550
rect 2040 505 2060 540
rect 2180 530 2190 540
rect 2210 530 2220 550
rect 2180 520 2220 530
rect 4070 490 4110 500
rect 4070 470 4080 490
rect 4100 470 4110 490
rect 4070 460 4110 470
rect 2305 275 2345 285
rect -130 260 -90 270
rect -130 240 -120 260
rect -100 240 -90 260
rect 2305 255 2315 275
rect 2335 255 2345 275
rect 2305 245 2345 255
rect -130 230 -90 240
rect 2735 165 2785 180
rect 2735 145 2750 165
rect 2770 145 2785 165
rect 2735 130 2785 145
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
rect 2380 30 2430 40
rect 2355 10 2390 30
rect 2380 0 2390 10
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 2380 -125 2430 -115
rect 2380 -155 2390 -125
rect 2420 -135 2430 -125
rect 7550 -135 7570 30
rect 2420 -155 2460 -135
rect 2480 -155 2510 -135
rect 2530 -155 2560 -135
rect 2580 -155 2610 -135
rect 2630 -155 2660 -135
rect 2680 -155 2710 -135
rect 2730 -155 2760 -135
rect 2780 -155 2810 -135
rect 2830 -155 2860 -135
rect 2880 -155 2910 -135
rect 2930 -155 2960 -135
rect 2980 -155 3010 -135
rect 3030 -155 3060 -135
rect 3080 -155 3110 -135
rect 3130 -155 3160 -135
rect 3180 -155 3210 -135
rect 3230 -155 3260 -135
rect 3280 -155 3310 -135
rect 3330 -155 3360 -135
rect 3380 -155 3410 -135
rect 3430 -155 3460 -135
rect 3480 -155 3510 -135
rect 3530 -155 3560 -135
rect 3580 -155 3610 -135
rect 3630 -155 3660 -135
rect 3680 -155 3710 -135
rect 3730 -155 3760 -135
rect 3780 -155 3810 -135
rect 3830 -155 3860 -135
rect 3880 -155 3910 -135
rect 3930 -155 3960 -135
rect 3980 -155 4010 -135
rect 4030 -155 4060 -135
rect 4080 -155 4110 -135
rect 4130 -155 4160 -135
rect 4180 -155 4210 -135
rect 4230 -155 4260 -135
rect 4280 -155 4310 -135
rect 4330 -155 4360 -135
rect 4380 -155 4410 -135
rect 4430 -155 4460 -135
rect 4480 -155 4510 -135
rect 4530 -155 4560 -135
rect 4580 -155 4610 -135
rect 4630 -155 4660 -135
rect 4680 -155 4710 -135
rect 4730 -155 4760 -135
rect 4780 -155 4810 -135
rect 4830 -155 4860 -135
rect 4880 -155 4910 -135
rect 4930 -155 4945 -135
rect 6180 -155 6210 -135
rect 6230 -155 6260 -135
rect 6280 -155 6310 -135
rect 6330 -155 6360 -135
rect 6380 -155 6410 -135
rect 6430 -155 6460 -135
rect 6480 -155 6510 -135
rect 6530 -155 6560 -135
rect 6580 -155 6610 -135
rect 6630 -155 6660 -135
rect 6680 -155 6710 -135
rect 6730 -155 6760 -135
rect 6780 -155 6810 -135
rect 6830 -155 6860 -135
rect 6880 -155 6910 -135
rect 6930 -155 6960 -135
rect 6980 -155 7010 -135
rect 7030 -155 7060 -135
rect 7080 -155 7110 -135
rect 7130 -155 7160 -135
rect 7180 -155 7210 -135
rect 7230 -155 7260 -135
rect 7280 -155 7310 -135
rect 7330 -155 7360 -135
rect 7380 -155 7410 -135
rect 7430 -155 7460 -135
rect 7480 -155 7510 -135
rect 7530 -155 7570 -135
rect 2380 -165 2430 -155
rect 6010 -310 6050 -300
rect 6010 -330 6020 -310
rect 6040 -330 6050 -310
rect 6010 -340 6050 -330
rect -330 -585 -290 -575
rect -330 -605 -320 -585
rect -300 -605 -290 -585
rect -330 -615 -290 -605
rect -330 -775 -280 -765
rect -330 -805 -320 -775
rect -290 -805 -280 -775
rect -330 -815 -280 -805
<< viali >>
rect 2790 2795 2810 2815
rect 4830 2520 4850 2540
rect 2790 2200 2810 2220
rect 2390 1190 2420 1220
rect 2050 1135 2070 1155
rect 2750 995 2770 1015
rect 2190 925 2210 945
rect 2310 925 2330 945
rect 3100 660 3120 680
rect 3860 660 3880 680
rect -180 595 -150 625
rect 2350 600 2370 620
rect 2400 600 2420 620
rect 2475 605 2495 625
rect 3165 625 3185 645
rect 4460 575 4480 595
rect 2190 530 2210 550
rect 3065 520 3085 540
rect 4080 470 4100 490
rect -120 240 -100 260
rect 2315 255 2335 275
rect 2750 145 2770 165
rect 2085 65 2105 85
rect 2390 0 2420 30
rect 2390 -155 2420 -125
rect 2460 -155 2480 -135
rect 2510 -155 2530 -135
rect 2560 -155 2580 -135
rect 2610 -155 2630 -135
rect 2660 -155 2680 -135
rect 2710 -155 2730 -135
rect 2760 -155 2780 -135
rect 2810 -155 2830 -135
rect 2860 -155 2880 -135
rect 2910 -155 2930 -135
rect 2960 -155 2980 -135
rect 3010 -155 3030 -135
rect 3060 -155 3080 -135
rect 3110 -155 3130 -135
rect 3160 -155 3180 -135
rect 3210 -155 3230 -135
rect 3260 -155 3280 -135
rect 3310 -155 3330 -135
rect 3360 -155 3380 -135
rect 3410 -155 3430 -135
rect 3460 -155 3480 -135
rect 3510 -155 3530 -135
rect 3560 -155 3580 -135
rect 3610 -155 3630 -135
rect 3660 -155 3680 -135
rect 3710 -155 3730 -135
rect 3760 -155 3780 -135
rect 3810 -155 3830 -135
rect 3860 -155 3880 -135
rect 3910 -155 3930 -135
rect 3960 -155 3980 -135
rect 4010 -155 4030 -135
rect 4060 -155 4080 -135
rect 4110 -155 4130 -135
rect 4160 -155 4180 -135
rect 4210 -155 4230 -135
rect 4260 -155 4280 -135
rect 4310 -155 4330 -135
rect 4360 -155 4380 -135
rect 4410 -155 4430 -135
rect 4460 -155 4480 -135
rect 4510 -155 4530 -135
rect 4560 -155 4580 -135
rect 4610 -155 4630 -135
rect 4660 -155 4680 -135
rect 4710 -155 4730 -135
rect 4760 -155 4780 -135
rect 4810 -155 4830 -135
rect 4860 -155 4880 -135
rect 4910 -155 4930 -135
rect 6160 -155 6180 -135
rect 6210 -155 6230 -135
rect 6260 -155 6280 -135
rect 6310 -155 6330 -135
rect 6360 -155 6380 -135
rect 6410 -155 6430 -135
rect 6460 -155 6480 -135
rect 6510 -155 6530 -135
rect 6560 -155 6580 -135
rect 6610 -155 6630 -135
rect 6660 -155 6680 -135
rect 6710 -155 6730 -135
rect 6760 -155 6780 -135
rect 6810 -155 6830 -135
rect 6860 -155 6880 -135
rect 6910 -155 6930 -135
rect 6960 -155 6980 -135
rect 7010 -155 7030 -135
rect 7060 -155 7080 -135
rect 7110 -155 7130 -135
rect 7160 -155 7180 -135
rect 7210 -155 7230 -135
rect 7260 -155 7280 -135
rect 7310 -155 7330 -135
rect 7360 -155 7380 -135
rect 7410 -155 7430 -135
rect 7460 -155 7480 -135
rect 7510 -155 7530 -135
rect 6020 -330 6040 -310
rect -320 -605 -300 -585
rect -320 -805 -290 -775
<< metal1 >>
rect 2775 2820 2825 2830
rect 2775 2790 2785 2820
rect 2815 2790 2825 2820
rect 2775 2780 2825 2790
rect 2635 2595 2675 2600
rect 2635 2565 2640 2595
rect 2670 2580 2675 2595
rect 2670 2565 3005 2580
rect 2635 2560 2675 2565
rect 4820 2540 4860 2550
rect 5975 2545 6015 2550
rect 5975 2540 5980 2545
rect 4820 2520 4830 2540
rect 4850 2525 5980 2540
rect 4850 2520 4860 2525
rect 2580 2510 2620 2515
rect 4820 2510 4860 2520
rect 5975 2515 5980 2525
rect 6010 2515 6015 2545
rect 5975 2510 6015 2515
rect 2580 2480 2585 2510
rect 2615 2500 2620 2510
rect 2615 2485 3005 2500
rect 2615 2480 2620 2485
rect 2580 2475 2620 2480
rect 2775 2225 2825 2235
rect 2775 2195 2785 2225
rect 2815 2195 2825 2225
rect 2775 2185 2825 2195
rect 2690 1390 2730 1395
rect 2690 1360 2695 1390
rect 2725 1380 2730 1390
rect 5975 1385 6015 1390
rect 5975 1380 5980 1385
rect 2725 1365 5980 1380
rect 2725 1360 2730 1365
rect 2690 1355 2730 1360
rect 5975 1355 5980 1365
rect 6010 1355 6015 1385
rect 5975 1350 6015 1355
rect 2580 1335 2620 1340
rect 2580 1305 2585 1335
rect 2615 1325 2620 1335
rect 5450 1330 5490 1335
rect 5450 1325 5455 1330
rect 2615 1310 5455 1325
rect 2615 1305 2620 1310
rect 2580 1300 2620 1305
rect 5450 1300 5455 1310
rect 5485 1300 5490 1330
rect 5450 1295 5490 1300
rect 2540 1280 2580 1285
rect 2540 1250 2545 1280
rect 2575 1275 2580 1280
rect 2575 1260 2805 1275
rect 2575 1250 2580 1260
rect 2540 1245 2580 1250
rect 2380 1220 2430 1230
rect 2355 1190 2390 1220
rect 2420 1190 2430 1220
rect 2355 1180 2430 1190
rect 2040 1155 2080 1165
rect 2040 1135 2050 1155
rect 2070 1150 2080 1155
rect 2580 1160 2620 1165
rect 2580 1150 2585 1160
rect 2070 1135 2585 1150
rect 2040 1125 2080 1135
rect 2580 1130 2585 1135
rect 2615 1130 2620 1160
rect 2580 1125 2620 1130
rect 2180 1095 2220 1100
rect 2180 1065 2185 1095
rect 2215 1085 2220 1095
rect 2535 1095 2575 1100
rect 2535 1085 2540 1095
rect 2215 1070 2540 1085
rect 2215 1065 2220 1070
rect 2180 1060 2220 1065
rect 2535 1065 2540 1070
rect 2570 1065 2575 1095
rect 2535 1060 2575 1065
rect 2735 1020 2785 1030
rect 2735 990 2745 1020
rect 2775 990 2785 1020
rect 2735 980 2785 990
rect 2180 950 2220 955
rect 2180 920 2185 950
rect 2215 920 2220 950
rect 2180 915 2220 920
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 940 2340 945
rect 2535 950 2575 955
rect 2535 940 2540 950
rect 2330 925 2540 940
rect 2300 915 2340 925
rect 2535 920 2540 925
rect 2570 920 2575 950
rect 2535 915 2575 920
rect 2580 695 2620 700
rect 2580 665 2585 695
rect 2615 685 2620 695
rect 2690 695 2730 700
rect 2690 685 2695 695
rect 2615 670 2695 685
rect 2615 665 2620 670
rect 2580 660 2620 665
rect 2690 665 2695 670
rect 2725 675 2730 695
rect 3090 680 3130 690
rect 3090 675 3100 680
rect 2725 665 3100 675
rect 2690 660 3100 665
rect 3120 660 3130 680
rect 2635 650 2675 655
rect 3090 650 3130 660
rect 3850 685 3890 690
rect 3850 655 3855 685
rect 3885 655 3890 685
rect -190 630 -140 635
rect 2460 630 2510 640
rect -190 625 -115 630
rect -190 595 -180 625
rect -150 595 -115 625
rect 2355 620 2470 630
rect 2370 600 2400 620
rect 2420 600 2470 620
rect 2500 600 2510 630
rect 2635 620 2640 650
rect 2670 635 2675 650
rect 3155 645 3195 655
rect 3850 650 3890 655
rect 3155 635 3165 645
rect 2670 625 3165 635
rect 3185 625 3195 645
rect 2670 620 3195 625
rect 2635 615 2675 620
rect 3155 615 3195 620
rect 3850 615 3890 620
rect -190 590 -115 595
rect 2355 590 2510 600
rect 2535 610 2575 615
rect -190 585 -140 590
rect 2535 580 2540 610
rect 2570 600 2575 610
rect 3850 600 3855 615
rect 2570 585 3855 600
rect 3885 585 3890 615
rect 2570 580 2575 585
rect 3850 580 3890 585
rect 4450 595 4490 605
rect 2535 575 2575 580
rect 4450 575 4460 595
rect 4480 590 4490 595
rect 5450 595 5490 600
rect 5450 590 5455 595
rect 4480 575 5455 590
rect 4450 565 4490 575
rect 5450 565 5455 575
rect 5485 565 5490 595
rect 5450 560 5490 565
rect 2180 550 2220 560
rect 2180 530 2190 550
rect 2210 535 2220 550
rect 3055 540 3095 550
rect 3055 535 3065 540
rect 2210 530 3065 535
rect 2180 520 3065 530
rect 3085 520 3095 540
rect 3055 510 3095 520
rect 2535 495 2575 500
rect 2535 465 2540 495
rect 2570 490 2575 495
rect 4070 490 4110 500
rect 2570 475 4080 490
rect 2570 465 2575 475
rect 2535 460 2575 465
rect 4070 470 4080 475
rect 4100 470 4110 490
rect 4070 460 4110 470
rect 2305 275 2345 285
rect -335 265 -295 270
rect -335 235 -330 265
rect -300 260 -295 265
rect -130 260 -90 270
rect -300 245 -120 260
rect -300 235 -295 245
rect -335 230 -295 235
rect -130 240 -120 245
rect -100 240 -90 260
rect 2305 255 2315 275
rect 2335 270 2345 275
rect 2535 280 2575 285
rect 2535 270 2540 280
rect 2335 255 2540 270
rect 2305 245 2345 255
rect 2535 250 2540 255
rect 2570 250 2575 280
rect 2535 245 2575 250
rect -130 230 -90 240
rect 2735 170 2785 180
rect 2735 140 2745 170
rect 2775 140 2785 170
rect 2735 130 2785 140
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 70 2740 85
rect 2105 65 2115 70
rect 2075 55 2115 65
rect 2355 30 2430 40
rect 2355 0 2390 30
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 6010 -5 6065 0
rect 5450 -10 5490 -5
rect 5450 -40 5455 -10
rect 5485 -15 5490 -10
rect 6010 -15 6015 -5
rect 5485 -30 6015 -15
rect 5485 -40 5490 -30
rect 6010 -35 6015 -30
rect 6045 -15 6065 -5
rect 6045 -30 6610 -15
rect 6045 -35 6065 -30
rect 6010 -40 6065 -35
rect 5450 -45 5490 -40
rect 2380 -125 2430 -115
rect 2380 -155 2390 -125
rect 2420 -135 4945 -125
rect 6180 -135 7570 -125
rect 2420 -155 2460 -135
rect 2480 -155 2510 -135
rect 2530 -155 2560 -135
rect 2580 -155 2610 -135
rect 2630 -155 2660 -135
rect 2680 -155 2710 -135
rect 2730 -155 2760 -135
rect 2780 -155 2810 -135
rect 2830 -155 2860 -135
rect 2880 -155 2910 -135
rect 2930 -155 2960 -135
rect 2980 -155 3010 -135
rect 3030 -155 3060 -135
rect 3080 -155 3110 -135
rect 3130 -155 3160 -135
rect 3180 -155 3210 -135
rect 3230 -155 3260 -135
rect 3280 -155 3310 -135
rect 3330 -155 3360 -135
rect 3380 -155 3410 -135
rect 3430 -155 3460 -135
rect 3480 -155 3510 -135
rect 3530 -155 3560 -135
rect 3580 -155 3610 -135
rect 3630 -155 3660 -135
rect 3680 -155 3710 -135
rect 3730 -155 3760 -135
rect 3780 -155 3810 -135
rect 3830 -155 3860 -135
rect 3880 -155 3910 -135
rect 3930 -155 3960 -135
rect 3980 -155 4010 -135
rect 4030 -155 4060 -135
rect 4080 -155 4110 -135
rect 4130 -155 4160 -135
rect 4180 -155 4210 -135
rect 4230 -155 4260 -135
rect 4280 -155 4310 -135
rect 4330 -155 4360 -135
rect 4380 -155 4410 -135
rect 4430 -155 4460 -135
rect 4480 -155 4510 -135
rect 4530 -155 4560 -135
rect 4580 -155 4610 -135
rect 4630 -155 4660 -135
rect 4680 -155 4710 -135
rect 4730 -155 4760 -135
rect 4780 -155 4810 -135
rect 4830 -155 4860 -135
rect 4880 -155 4910 -135
rect 4930 -155 4945 -135
rect 6180 -155 6210 -135
rect 6230 -155 6260 -135
rect 6280 -155 6310 -135
rect 6330 -155 6360 -135
rect 6380 -155 6410 -135
rect 6430 -155 6460 -135
rect 6480 -155 6510 -135
rect 6530 -155 6560 -135
rect 6580 -155 6610 -135
rect 6630 -155 6660 -135
rect 6680 -155 6710 -135
rect 6730 -155 6760 -135
rect 6780 -155 6810 -135
rect 6830 -155 6860 -135
rect 6880 -155 6910 -135
rect 6930 -155 6960 -135
rect 6980 -155 7010 -135
rect 7030 -155 7060 -135
rect 7080 -155 7110 -135
rect 7130 -155 7160 -135
rect 7180 -155 7210 -135
rect 7230 -155 7260 -135
rect 7280 -155 7310 -135
rect 7330 -155 7360 -135
rect 7380 -155 7410 -135
rect 7430 -155 7460 -135
rect 7480 -155 7510 -135
rect 7530 -155 7570 -135
rect 2380 -165 4945 -155
rect 6180 -165 7570 -155
rect 6010 -305 6050 -300
rect 6010 -335 6015 -305
rect 6045 -335 6050 -305
rect 6010 -340 6050 -335
rect -330 -580 -290 -575
rect -330 -610 -325 -580
rect -295 -610 -290 -580
rect -330 -615 -290 -610
rect -330 -775 -280 -765
rect -330 -805 -320 -775
rect -290 -805 -280 -775
rect -330 -815 -280 -805
<< via1 >>
rect 2785 2815 2815 2820
rect 2785 2795 2790 2815
rect 2790 2795 2810 2815
rect 2810 2795 2815 2815
rect 2785 2790 2815 2795
rect 2640 2565 2670 2595
rect 5980 2515 6010 2545
rect 2585 2480 2615 2510
rect 2785 2220 2815 2225
rect 2785 2200 2790 2220
rect 2790 2200 2810 2220
rect 2810 2200 2815 2220
rect 2785 2195 2815 2200
rect 2695 1360 2725 1390
rect 5980 1355 6010 1385
rect 2585 1305 2615 1335
rect 5455 1300 5485 1330
rect 2545 1250 2575 1280
rect 2390 1190 2420 1220
rect 2585 1130 2615 1160
rect 2185 1065 2215 1095
rect 2540 1065 2570 1095
rect 2745 1015 2775 1020
rect 2745 995 2750 1015
rect 2750 995 2770 1015
rect 2770 995 2775 1015
rect 2745 990 2775 995
rect 2185 945 2215 950
rect 2185 925 2190 945
rect 2190 925 2210 945
rect 2210 925 2215 945
rect 2185 920 2215 925
rect 2540 920 2570 950
rect 2585 665 2615 695
rect 2695 665 2725 695
rect 3855 680 3885 685
rect 3855 660 3860 680
rect 3860 660 3880 680
rect 3880 660 3885 680
rect 3855 655 3885 660
rect -180 595 -150 625
rect 2470 625 2500 630
rect 2470 605 2475 625
rect 2475 605 2495 625
rect 2495 605 2500 625
rect 2470 600 2500 605
rect 2640 620 2670 650
rect 2540 580 2570 610
rect 3855 585 3885 615
rect 5455 565 5485 595
rect 2540 465 2570 495
rect -330 235 -300 265
rect 2540 250 2570 280
rect 2745 165 2775 170
rect 2745 145 2750 165
rect 2750 145 2770 165
rect 2770 145 2775 165
rect 2745 140 2775 145
rect 2390 0 2420 30
rect 5455 -40 5485 -10
rect 6015 -35 6045 -5
rect 2390 -155 2420 -125
rect 6015 -310 6045 -305
rect 6015 -330 6020 -310
rect 6020 -330 6040 -310
rect 6040 -330 6045 -310
rect 6015 -335 6045 -330
rect -325 -585 -295 -580
rect -325 -605 -320 -585
rect -320 -605 -300 -585
rect -300 -605 -295 -585
rect -325 -610 -295 -605
rect -320 -805 -290 -775
<< metal2 >>
rect 2775 2820 2825 2830
rect 2775 2790 2785 2820
rect 2815 2790 2825 2820
rect 2775 2780 2825 2790
rect 2635 2595 2675 2600
rect 2635 2565 2640 2595
rect 2670 2565 2675 2595
rect 2635 2560 2675 2565
rect 2580 2510 2620 2515
rect 2580 2480 2585 2510
rect 2615 2480 2620 2510
rect 2580 2475 2620 2480
rect 2590 1340 2605 2475
rect 2580 1335 2620 1340
rect 2580 1305 2585 1335
rect 2615 1305 2620 1335
rect 2580 1300 2620 1305
rect 2540 1280 2580 1285
rect 2540 1250 2545 1280
rect 2575 1250 2580 1280
rect 2540 1245 2580 1250
rect 2380 1220 2430 1230
rect 2380 1190 2390 1220
rect 2420 1190 2430 1220
rect 2380 1180 2430 1190
rect 2550 1100 2565 1245
rect 2580 1160 2620 1165
rect 2580 1130 2585 1160
rect 2615 1130 2620 1160
rect 2580 1125 2620 1130
rect 2180 1095 2220 1100
rect 2180 1065 2185 1095
rect 2215 1065 2220 1095
rect 2180 1060 2220 1065
rect 2535 1095 2575 1100
rect 2535 1065 2540 1095
rect 2570 1065 2575 1095
rect 2535 1060 2575 1065
rect 2195 955 2210 1060
rect 2180 950 2220 955
rect 2180 920 2185 950
rect 2215 920 2220 950
rect 2180 915 2220 920
rect 2535 950 2575 955
rect 2535 920 2540 950
rect 2570 920 2575 950
rect 2535 915 2575 920
rect -190 625 -140 635
rect -190 595 -180 625
rect -150 595 -140 625
rect -190 585 -140 595
rect 2460 630 2510 640
rect 2460 600 2470 630
rect 2500 600 2510 630
rect 2550 615 2565 915
rect 2590 700 2605 1125
rect 2580 695 2620 700
rect 2580 665 2585 695
rect 2615 665 2620 695
rect 2580 660 2620 665
rect 2650 655 2665 2560
rect 5975 2545 6015 2550
rect 5975 2515 5980 2545
rect 6010 2515 6015 2545
rect 5975 2510 6015 2515
rect 2775 2225 2825 2235
rect 2775 2195 2785 2225
rect 2815 2195 2825 2225
rect 2775 2185 2825 2195
rect 2690 1390 2730 1395
rect 5985 1390 6000 2510
rect 2690 1360 2695 1390
rect 2725 1360 2730 1390
rect 2690 1355 2730 1360
rect 5975 1385 6015 1390
rect 5975 1355 5980 1385
rect 6010 1355 6015 1385
rect 2705 700 2720 1355
rect 5975 1350 6015 1355
rect 5450 1330 5490 1335
rect 5450 1300 5455 1330
rect 5485 1300 5490 1330
rect 5450 1295 5490 1300
rect 2735 1020 2785 1030
rect 2735 990 2745 1020
rect 2775 990 2785 1020
rect 2735 980 2785 990
rect 2690 695 2730 700
rect 2690 665 2695 695
rect 2725 665 2730 695
rect 2690 660 2730 665
rect 3850 685 3890 690
rect 3850 655 3855 685
rect 3885 655 3890 685
rect 2635 650 2675 655
rect 3850 650 3890 655
rect 2635 620 2640 650
rect 2670 620 2675 650
rect 3860 620 3875 650
rect 2635 615 2675 620
rect 3850 615 3890 620
rect 2460 590 2510 600
rect 2535 610 2575 615
rect 2535 580 2540 610
rect 2570 580 2575 610
rect 3850 585 3855 615
rect 3885 585 3890 615
rect 5465 600 5480 1295
rect 3850 580 3890 585
rect 5450 595 5490 600
rect 2535 575 2575 580
rect 5450 565 5455 595
rect 5485 565 5490 595
rect 5450 560 5490 565
rect 2535 495 2575 500
rect 2535 465 2540 495
rect 2570 465 2575 495
rect 2535 460 2575 465
rect 2550 285 2565 460
rect 2535 280 2575 285
rect -335 265 -295 270
rect -335 235 -330 265
rect -300 235 -295 265
rect 2535 250 2540 280
rect 2570 250 2575 280
rect 2535 245 2575 250
rect -335 230 -295 235
rect -320 -575 -305 230
rect 2735 170 2785 180
rect 2735 140 2745 170
rect 2775 140 2785 170
rect 2735 130 2785 140
rect 2380 30 2430 40
rect 2380 0 2390 30
rect 2420 0 2430 30
rect 2380 -10 2430 0
rect 5465 -5 5480 560
rect 6010 -5 6065 0
rect 5450 -10 5490 -5
rect 5450 -40 5455 -10
rect 5485 -40 5490 -10
rect 6010 -35 6015 -5
rect 6045 -35 6065 -5
rect 6010 -40 6065 -35
rect 5450 -45 5490 -40
rect 2380 -125 2430 -115
rect 2380 -155 2390 -125
rect 2420 -155 2430 -125
rect 2380 -165 2430 -155
rect 6020 -300 6035 -40
rect 6010 -305 6050 -300
rect 6010 -335 6015 -305
rect 6045 -335 6050 -305
rect 6010 -340 6050 -335
rect -330 -580 -290 -575
rect -330 -610 -325 -580
rect -295 -610 -290 -580
rect -330 -615 -290 -610
rect -330 -775 -280 -765
rect -330 -805 -320 -775
rect -290 -805 -280 -775
rect -330 -815 -280 -805
<< via2 >>
rect 2785 2790 2815 2820
rect 2390 1190 2420 1220
rect -180 595 -150 625
rect 2470 600 2500 630
rect 2785 2195 2815 2225
rect 2745 990 2775 1020
rect 2745 140 2775 170
rect 2390 0 2420 30
rect 2390 -155 2420 -125
rect -320 -805 -290 -775
<< metal3 >>
rect 2380 2825 2825 2830
rect 2380 2785 2385 2825
rect 2425 2820 2825 2825
rect 2425 2790 2785 2820
rect 2815 2790 2825 2820
rect 2425 2785 2825 2790
rect 2380 2780 2825 2785
rect 2460 2230 2825 2235
rect 2460 2190 2465 2230
rect 2505 2225 2825 2230
rect 2505 2195 2785 2225
rect 2815 2195 2825 2225
rect 2505 2190 2825 2195
rect 2460 2185 2825 2190
rect 2380 1225 2430 1230
rect 2380 1185 2385 1225
rect 2425 1185 2430 1225
rect 2380 1180 2430 1185
rect 2460 1025 2785 1030
rect 2460 985 2465 1025
rect 2505 1020 2785 1025
rect 2505 990 2745 1020
rect 2775 990 2785 1020
rect 2505 985 2785 990
rect 2460 980 2785 985
rect 2460 635 2510 640
rect -430 630 -140 635
rect -430 590 -425 630
rect -385 625 -140 630
rect -385 595 -180 625
rect -150 595 -140 625
rect -385 590 -140 595
rect 2460 595 2465 635
rect 2505 595 2510 635
rect 2460 590 2510 595
rect -430 585 -140 590
rect 2380 175 2785 180
rect 2380 135 2385 175
rect 2425 170 2785 175
rect 2425 140 2745 170
rect 2775 140 2785 170
rect 2425 135 2785 140
rect 2380 130 2785 135
rect 2380 35 2430 40
rect 2380 -5 2385 35
rect 2425 -5 2430 35
rect 2380 -10 2430 -5
rect 2380 -120 2430 -115
rect 2380 -160 2385 -120
rect 2425 -160 2430 -120
rect 2380 -165 2430 -160
rect -430 -770 -280 -765
rect -430 -810 -425 -770
rect -385 -775 -280 -770
rect -385 -805 -320 -775
rect -290 -805 -280 -775
rect -385 -810 -280 -805
rect -430 -815 -280 -810
<< via3 >>
rect 2385 2785 2425 2825
rect 2465 2190 2505 2230
rect 2385 1220 2425 1225
rect 2385 1190 2390 1220
rect 2390 1190 2420 1220
rect 2420 1190 2425 1220
rect 2385 1185 2425 1190
rect 2465 985 2505 1025
rect -425 590 -385 630
rect 2465 630 2505 635
rect 2465 600 2470 630
rect 2470 600 2500 630
rect 2500 600 2505 630
rect 2465 595 2505 600
rect 2385 135 2425 175
rect 2385 30 2425 35
rect 2385 0 2390 30
rect 2390 0 2420 30
rect 2420 0 2425 30
rect 2385 -5 2425 0
rect 2385 -125 2425 -120
rect 2385 -155 2390 -125
rect 2390 -155 2420 -125
rect 2420 -155 2425 -125
rect 2385 -160 2425 -155
rect -425 -810 -385 -770
<< metal4 >>
rect 2380 2825 2430 2830
rect 2380 2785 2385 2825
rect 2425 2785 2430 2825
rect 2380 1225 2430 2785
rect 2380 1185 2385 1225
rect 2425 1185 2430 1225
rect -430 630 -380 635
rect -430 590 -425 630
rect -385 590 -380 630
rect -430 -770 -380 590
rect 2380 175 2430 1185
rect 2460 2230 2510 2235
rect 2460 2190 2465 2230
rect 2505 2190 2510 2230
rect 2460 1025 2510 2190
rect 2460 985 2465 1025
rect 2505 985 2510 1025
rect 2460 635 2510 985
rect 2460 595 2465 635
rect 2505 595 2510 635
rect 2460 590 2510 595
rect -280 105 -230 155
rect 2380 135 2385 175
rect 2425 135 2430 175
rect 2380 35 2430 135
rect 2380 -5 2385 35
rect 2425 -5 2430 35
rect 2380 -120 2430 -5
rect 2380 -160 2385 -120
rect 2425 -160 2430 -120
rect 2380 -165 2430 -160
rect -430 -810 -425 -770
rect -385 -810 -380 -770
rect -430 -815 -380 -810
use charge_pump_cell_6  charge_pump_cell_6_0
timestamp 1740156359
transform 1 0 -6370 0 1 -1565
box 9105 1615 11630 2860
use loop_filter_2  loop_filter_2_0
timestamp 1740116583
transform 1 0 4930 0 -1 290
box 1135 -5975 9720 330
use opamp_cell_4  opamp_cell_4_0
timestamp 1740145811
transform 1 0 -425 0 -1 4625
box 3110 897 6365 3205
use pfd_8  pfd_8_0
timestamp 1739770731
transform 1 0 -930 0 1 4655
box 650 -4655 3290 -3435
use VCO_FD_magic  VCO_FD_magic_0
timestamp 1740284885
transform -1 0 6180 0 -1 -65
box 0 60 6470 1150
<< labels >>
flabel metal1 -140 610 -140 610 7 FreeSans 400 0 -200 0 VDDA
port 2 w
flabel metal4 -280 130 -280 130 7 FreeSans 400 0 -200 0 GNDA
port 3 w
flabel poly -130 250 -130 250 7 FreeSans 400 0 -200 0 F_VCO
flabel poly -130 965 -130 965 7 FreeSans 400 0 -200 0 F_REF
port 4 w
flabel poly 4975 -585 4975 -585 1 FreeSans 400 0 0 200 V_OSC
port 1 n
flabel metal1 3095 530 3095 530 3 FreeSans 400 0 200 0 I_IN
port 5 e
flabel metal2 5480 730 5480 730 3 FreeSans 400 0 200 0 V_CONT
<< end >>
