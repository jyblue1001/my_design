magic
tech sky130A
timestamp 1738158477
<< nwell >>
rect -170 190 255 430
rect 470 190 835 430
<< pwell >>
rect 470 -5 835 105
<< nmos >>
rect 0 0 15 100
rect 700 0 715 100
<< pmos >>
rect 0 210 15 410
rect 700 210 715 410
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 650 85 700 100
rect 650 15 665 85
rect 685 15 700 85
rect 650 0 700 15
rect 715 85 765 100
rect 715 15 730 85
rect 750 15 765 85
rect 715 0 765 15
<< pdiff >>
rect -50 395 0 410
rect -50 225 -35 395
rect -15 225 0 395
rect -50 210 0 225
rect 15 395 65 410
rect 15 225 30 395
rect 50 225 65 395
rect 15 210 65 225
rect 650 395 700 410
rect 650 225 665 395
rect 685 225 700 395
rect 650 210 700 225
rect 715 395 765 410
rect 715 225 730 395
rect 750 225 765 395
rect 715 210 765 225
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 665 15 685 85
rect 730 15 750 85
<< pdiffc >>
rect -35 225 -15 395
rect 30 225 50 395
rect 665 225 685 395
rect 730 225 750 395
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
rect 475 85 525 100
rect 475 15 490 85
rect 510 15 525 85
rect 475 0 525 15
<< nsubdiff >>
rect -100 395 -50 410
rect -100 225 -85 395
rect -65 225 -50 395
rect -100 210 -50 225
rect 535 395 585 410
rect 535 225 550 395
rect 570 225 585 395
rect 535 210 585 225
<< psubdiffcont >>
rect -85 15 -65 85
rect 490 15 510 85
<< nsubdiffcont >>
rect -85 225 -65 395
rect 550 225 570 395
<< poly >>
rect 700 430 720 450
rect 0 410 15 425
rect 700 410 715 430
rect 0 165 15 210
rect 700 195 715 210
rect -185 150 15 165
rect 0 100 15 150
rect 700 100 715 115
rect 0 -15 15 0
rect 700 -20 715 0
rect 700 -40 720 -20
<< locali >>
rect -175 430 -85 450
rect -65 430 -40 450
rect -20 430 5 450
rect 25 430 50 450
rect 70 430 95 450
rect 115 430 140 450
rect 160 430 185 450
rect 205 430 230 450
rect 250 430 275 450
rect 295 430 320 450
rect 340 430 365 450
rect 385 430 410 450
rect 430 430 490 450
rect 510 430 545 450
rect 565 430 590 450
rect 610 430 635 450
rect 655 430 700 450
rect 720 430 770 450
rect 790 430 815 450
rect 835 430 860 450
rect -85 405 -65 430
rect -40 405 -20 430
rect -95 395 -5 405
rect -95 225 -85 395
rect -65 225 -35 395
rect -15 225 -5 395
rect -95 215 -5 225
rect 20 395 65 405
rect 20 225 30 395
rect 50 225 65 395
rect 20 215 65 225
rect 30 165 50 215
rect 30 145 145 165
rect 30 95 50 145
rect 490 95 510 430
rect 540 395 580 405
rect 540 225 550 395
rect 570 225 580 395
rect 540 215 580 225
rect 655 395 695 405
rect 655 225 665 395
rect 685 225 695 395
rect 655 215 695 225
rect 720 395 760 405
rect 720 225 730 395
rect 750 225 760 395
rect 720 215 760 225
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 20 85 60 95
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 480 85 520 95
rect 480 15 490 85
rect 510 15 520 85
rect 480 5 520 15
rect -85 -20 -65 5
rect -40 -20 -20 5
rect 550 -20 570 215
rect 665 195 685 215
rect 615 175 685 195
rect 665 95 685 175
rect 730 135 750 215
rect 730 115 880 135
rect 730 95 750 115
rect 655 85 695 95
rect 655 15 665 85
rect 685 15 695 85
rect 655 5 695 15
rect 720 85 760 95
rect 720 15 730 85
rect 750 15 760 85
rect 720 5 760 15
rect -180 -40 -85 -20
rect -65 -40 -40 -20
rect -20 -40 5 -20
rect 25 -40 50 -20
rect 70 -40 95 -20
rect 115 -40 140 -20
rect 160 -40 185 -20
rect 205 -40 230 -20
rect 250 -40 275 -20
rect 295 -40 320 -20
rect 340 -40 365 -20
rect 385 -40 410 -20
rect 430 -40 455 -20
rect 475 -40 500 -20
rect 520 -40 550 -20
rect 570 -40 635 -20
rect 655 -40 700 -20
rect 720 -40 770 -20
rect 790 -40 815 -20
rect 835 -40 860 -20
<< viali >>
rect -85 430 -65 450
rect -40 430 -20 450
rect 5 430 25 450
rect 50 430 70 450
rect 95 430 115 450
rect 140 430 160 450
rect 185 430 205 450
rect 230 430 250 450
rect 275 430 295 450
rect 320 430 340 450
rect 365 430 385 450
rect 410 430 430 450
rect 490 430 510 450
rect 545 430 565 450
rect 590 430 610 450
rect 635 430 655 450
rect 700 430 720 450
rect 770 430 790 450
rect 815 430 835 450
rect 860 430 880 450
rect -85 -40 -65 -20
rect -40 -40 -20 -20
rect 5 -40 25 -20
rect 50 -40 70 -20
rect 95 -40 115 -20
rect 140 -40 160 -20
rect 185 -40 205 -20
rect 230 -40 250 -20
rect 275 -40 295 -20
rect 320 -40 340 -20
rect 365 -40 385 -20
rect 410 -40 430 -20
rect 455 -40 475 -20
rect 500 -40 520 -20
rect 550 -40 570 -20
rect 635 -40 655 -20
rect 700 -40 720 -20
rect 770 -40 790 -20
rect 815 -40 835 -20
rect 860 -40 880 -20
<< metal1 >>
rect -175 450 885 465
rect -175 430 -85 450
rect -65 430 -40 450
rect -20 430 5 450
rect 25 430 50 450
rect 70 430 95 450
rect 115 430 140 450
rect 160 430 185 450
rect 205 430 230 450
rect 250 430 275 450
rect 295 430 320 450
rect 340 430 365 450
rect 385 430 410 450
rect 430 430 490 450
rect 510 430 545 450
rect 565 430 590 450
rect 610 430 635 450
rect 655 430 700 450
rect 720 430 770 450
rect 790 430 815 450
rect 835 430 860 450
rect 880 430 885 450
rect -175 415 885 430
rect -180 -20 885 -5
rect -180 -40 -85 -20
rect -65 -40 -40 -20
rect -20 -40 5 -20
rect 25 -40 50 -20
rect 70 -40 95 -20
rect 115 -40 140 -20
rect 160 -40 185 -20
rect 205 -40 230 -20
rect 250 -40 275 -20
rect 295 -40 320 -20
rect 340 -40 365 -20
rect 385 -40 410 -20
rect 430 -40 455 -20
rect 475 -40 500 -20
rect 520 -40 550 -20
rect 570 -40 635 -20
rect 655 -40 700 -20
rect 720 -40 770 -20
rect 790 -40 815 -20
rect 835 -40 860 -20
rect 880 -40 885 -20
rect -180 -55 885 -40
<< labels >>
flabel locali 145 155 145 155 3 FreeSans 400 0 80 0 B
flabel poly -185 155 -185 155 7 FreeSans 400 0 -80 0 A
flabel metal1 -175 440 -175 440 7 FreeSans 400 0 -80 0 VDDA
flabel metal1 -180 -30 -180 -30 7 FreeSans 400 0 -80 0 GNDA
flabel locali 880 125 880 125 3 FreeSans 400 0 80 0 D
flabel locali 615 185 615 185 7 FreeSans 400 0 -80 0 C
<< end >>
