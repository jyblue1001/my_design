** sch_path: /foss/designs/my_design/projects/pll/pfd/magic/tb_phase_frequency_detector_magic.sch
**.subckt tb_phase_frequency_detector_magic
V1 F_REF GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
V2 F_VCO GND pulse(0 1.8 13ns 1ns 1ns 24ns 50ns)
VDD VDDA GND 1.8
x1 F_REF F_VCO VDDA QA QB GND phase_frequency_detector_magic
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /foss/designs/my_design/projects/pll/pfd/magic/phase_frequency_detector_magic.spice

.option wnflag=1
.option method=gear trtol=1

.control

  save all
  tran 1ns 1us
  remzerovec
  write tb_phase_frequency_detector_magic.raw
  set appendwrite

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
