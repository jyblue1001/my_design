* PEX produced on Tue Aug  5 02:13:48 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_16.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_16 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 two_stage_opamp_dummy_magic_23_0.Vb3.t6 GNDA.t461 GNDA.t463 GNDA.t462 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X1 VOUT+.t16 two_stage_opamp_dummy_magic_23_0.Y.t25 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X2 GNDA.t586 bgr_11_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_23_0.Vb3.t7 GNDA.t585 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X3 VDDA.t424 GNDA.t507 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 VDDA.t425 GNDA.t508 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VDDA.t426 GNDA.t502 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VDDA.t427 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VDDA.t428 GNDA.t503 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VOUT-.t19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VDDA.t429 GNDA.t544 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_23_0.VD1.t10 two_stage_opamp_dummy_magic_23_0.Vb1.t12 two_stage_opamp_dummy_magic_23_0.X.t4 GNDA.t244 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X11 two_stage_opamp_dummy_magic_23_0.X.t14 two_stage_opamp_dummy_magic_23_0.Vb2.t11 two_stage_opamp_dummy_magic_23_0.VD3.t31 two_stage_opamp_dummy_magic_23_0.VD3.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X12 VOUT-.t14 VDDA.t390 VDDA.t392 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X13 GNDA.t292 a_5820_23644.t1 GNDA.t41 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X14 VOUT+.t19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 GNDA.t460 GNDA.t458 VDDA.t102 GNDA.t459 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X16 VDDA.t430 GNDA.t545 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDDA.t431 GNDA.t546 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 w_6100_17280.t27 bgr_11_0.V_mir1.t13 bgr_11_0.1st_Vout_1.t4 w_6100_17280.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X19 bgr_11_0.1st_Vout_1.t7 bgr_11_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VDDA.t432 GNDA.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 GNDA.t457 GNDA.t454 GNDA.t456 GNDA.t455 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X22 VDDA.t433 GNDA.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 VDDA.t79 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t1 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X24 two_stage_opamp_dummy_magic_23_0.VD2.t10 two_stage_opamp_dummy_magic_23_0.Vb1.t13 two_stage_opamp_dummy_magic_23_0.Y.t9 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X25 GNDA.t277 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_23_0.V_source.t39 GNDA.t276 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X26 VDDA.t434 GNDA.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 bgr_11_0.1st_Vout_1.t8 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 GNDA.t453 GNDA.t451 two_stage_opamp_dummy_magic_23_0.Vb2.t8 GNDA.t452 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X29 two_stage_opamp_dummy_magic_23_0.VD1.t9 two_stage_opamp_dummy_magic_23_0.Vb1.t14 two_stage_opamp_dummy_magic_23_0.X.t6 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X30 VOUT-.t20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 two_stage_opamp_dummy_magic_23_0.VD4.t15 two_stage_opamp_dummy_magic_23_0.Vb3.t8 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X32 VDDA.t435 GNDA.t359 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_23_0.X.t25 GNDA.t328 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X34 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.t3 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X35 VOUT-.t21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VDDA.t436 GNDA.t360 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VDDA.t437 GNDA.t361 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 GNDA.t166 a_6470_23450.t0 GNDA.t165 sky130_fd_pr__res_xhigh_po_0p35 l=6
X39 VDDA.t438 GNDA.t469 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VOUT+.t20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VDDA.t439 GNDA.t470 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT-.t22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VDDA.t440 GNDA.t471 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT-.t23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 GNDA.t233 bgr_11_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t2 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X46 w_6100_17280.t47 w_6100_17280.t45 VDDA.t53 w_6100_17280.t46 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X47 two_stage_opamp_dummy_magic_23_0.err_amp_out.t8 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_23_0.V_err_p.t12 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X48 VDDA.t182 two_stage_opamp_dummy_magic_23_0.Y.t26 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t13 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X49 VOUT+.t21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VOUT+.t22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 two_stage_opamp_dummy_magic_23_0.Vb2.t7 GNDA.t448 GNDA.t450 GNDA.t449 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X52 VDDA.t441 GNDA.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VDDA.t442 GNDA.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 VOUT+.t23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VDDA.t378 VDDA.t379 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 VDDA.t31 two_stage_opamp_dummy_magic_23_0.V_err_gate.t14 two_stage_opamp_dummy_magic_23_0.V_err_p.t6 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X57 VDDA.t443 GNDA.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VDDA.t444 GNDA.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 GNDA.t325 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t17 two_stage_opamp_dummy_magic_23_0.err_amp_out.t9 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X60 VOUT-.t24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VDDA.t84 two_stage_opamp_dummy_magic_23_0.V_err_gate.t15 a_7460_6300.t10 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X62 GNDA.t314 two_stage_opamp_dummy_magic_23_0.Y.t27 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t10 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X63 VOUT-.t25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 two_stage_opamp_dummy_magic_23_0.V_source.t6 VIN-.t0 two_stage_opamp_dummy_magic_23_0.VD1.t13 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X65 VDDA.t445 GNDA.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VDDA.t446 GNDA.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VDDA.t389 VDDA.t386 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X68 w_6100_17280.t61 bgr_11_0.1st_Vout_1.t9 VDDA.t80 w_6100_17280.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X69 VDDA.t385 VDDA.t383 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t11 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X70 two_stage_opamp_dummy_magic_23_0.err_amp_out.t7 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_23_0.V_err_p.t13 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X71 VDDA.t376 VDDA.t377 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT+.t24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VOUT-.t26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 VDDA.t447 GNDA.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VDDA.t448 GNDA.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VDDA.t449 GNDA.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VOUT-.t27 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 VOUT-.t28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VDDA.t142 two_stage_opamp_dummy_magic_23_0.Vb3.t9 two_stage_opamp_dummy_magic_23_0.VD3.t9 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X80 two_stage_opamp_dummy_magic_23_0.V_err_p.t8 two_stage_opamp_dummy_magic_23_0.V_err_gate.t16 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X81 VDDA.t450 GNDA.t541 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VOUT-.t29 two_stage_opamp_dummy_magic_23_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VDDA.t140 two_stage_opamp_dummy_magic_23_0.Vb3.t10 two_stage_opamp_dummy_magic_23_0.VD4.t14 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X84 VOUT+.t15 two_stage_opamp_dummy_magic_23_0.Y.t28 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X85 VDDA.t374 VDDA.t375 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT-.t30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 two_stage_opamp_dummy_magic_23_0.VD1.t15 VIN-.t1 two_stage_opamp_dummy_magic_23_0.V_source.t9 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X88 VOUT-.t31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VOUT+.t25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 VOUT-.t32 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 two_stage_opamp_dummy_magic_23_0.V_err_gate.t4 bgr_11_0.NFET_GATE_10uA.t7 GNDA.t235 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X92 two_stage_opamp_dummy_magic_23_0.Y.t3 two_stage_opamp_dummy_magic_23_0.Vb2.t12 two_stage_opamp_dummy_magic_23_0.VD4.t37 two_stage_opamp_dummy_magic_23_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X93 VDDA.t382 VDDA.t380 two_stage_opamp_dummy_magic_23_0.err_amp_out.t11 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X94 VDDA.t451 GNDA.t542 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 VOUT+.t26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT-.t33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT+.t27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 VDDA.t452 GNDA.t543 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VDDA.t453 GNDA.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 VDDA.t454 GNDA.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t13 two_stage_opamp_dummy_magic_23_0.X.t26 VDDA.t87 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X102 w_6100_17280.t25 bgr_11_0.V_mir1.t8 bgr_11_0.V_mir1.t9 w_6100_17280.t24 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X103 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_23_0.Y.t29 GNDA.t240 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X104 two_stage_opamp_dummy_magic_23_0.VD2.t21 VIN+.t0 two_stage_opamp_dummy_magic_23_0.V_source.t21 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X105 VDDA.t455 GNDA.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 VDDA.t456 GNDA.t538 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT-.t34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VDDA.t373 VDDA.t371 two_stage_opamp_dummy_magic_23_0.V_err_gate.t12 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X109 VDDA.t342 VDDA.t343 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 VOUT-.t35 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT+.t28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 w_6100_17280.t59 bgr_11_0.1st_Vout_1.t10 VDDA.t54 w_6100_17280.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X113 w_7200_15600.t31 VDDA.t457 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t3 w_7200_15600.t30 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X114 GNDA.t164 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_23_0.V_source.t38 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X115 VOUT-.t36 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VOUT-.t37 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VOUT+.t29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 GNDA.t447 GNDA.t445 two_stage_opamp_dummy_magic_23_0.Vb1.t9 GNDA.t446 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X119 VDDA.t458 GNDA.t539 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VDDA.t397 w_7200_15600.t43 w_7200_15600.t45 w_7200_15600.t44 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X121 two_stage_opamp_dummy_magic_23_0.VD1.t8 two_stage_opamp_dummy_magic_23_0.Vb1.t15 two_stage_opamp_dummy_magic_23_0.X.t5 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X122 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_23_0.X.t27 GNDA.t331 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X123 VOUT-.t38 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_23_0.X.t28 GNDA.t301 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X125 VDDA.t459 GNDA.t535 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VDDA.t460 GNDA.t536 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VDDA.t461 GNDA.t537 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VDDA.t462 GNDA.t533 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VDDA.t364 VDDA.t365 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VOUT+.t30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 a_12070_24908.t1 bgr_11_0.V_CUR_REF_REG.t0 GNDA.t289 sky130_fd_pr__res_xhigh_po_0p35 l=4
X132 VDDA.t138 two_stage_opamp_dummy_magic_23_0.Vb3.t11 two_stage_opamp_dummy_magic_23_0.VD4.t13 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X133 VOUT+.t31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VOUT-.t39 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 VDDA.t463 GNDA.t534 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 VOUT+.t32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 VOUT+.t33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VDDA.t464 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VDDA.t465 GNDA.t529 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VDDA.t370 VDDA.t369 w_6100_17280.t77 w_6100_17280.t76 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X141 VDDA.t466 GNDA.t530 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 two_stage_opamp_dummy_magic_23_0.X.t13 two_stage_opamp_dummy_magic_23_0.Vb1.t16 two_stage_opamp_dummy_magic_23_0.VD1.t7 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X143 VDDA.t368 VDDA.t366 VOUT-.t13 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X144 GNDA.t98 a_6520_18930# bgr_11_0.V_p_2.t0 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X145 VDDA.t363 VDDA.t361 bgr_11_0.NFET_GATE_10uA.t4 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X146 VDDA.t467 GNDA.t531 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 w_6100_17280.t23 bgr_11_0.V_mir1.t10 bgr_11_0.V_mir1.t11 w_6100_17280.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X148 VDDA.t468 GNDA.t527 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 VOUT+.t35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t1 w_7200_15600.t40 w_7200_15600.t42 w_7200_15600.t41 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X153 VDDA.t75 two_stage_opamp_dummy_magic_23_0.V_err_gate.t17 a_7460_6300.t9 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X154 GNDA.t53 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t15 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t16 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X155 VDDA.t469 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VDDA.t470 GNDA.t528 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VOUT-.t40 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X159 VDDA.t471 GNDA.t524 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VOUT-.t41 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT+.t36 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 w_6100_17280.t75 VDDA.t359 VDDA.t360 w_6100_17280.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X163 GNDA.t532 VDDA.t356 VDDA.t358 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X164 two_stage_opamp_dummy_magic_23_0.Y.t0 two_stage_opamp_dummy_magic_23_0.Vb1.t17 two_stage_opamp_dummy_magic_23_0.VD2.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X165 two_stage_opamp_dummy_magic_23_0.V_source.t37 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t14 GNDA.t555 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X166 two_stage_opamp_dummy_magic_23_0.V_source.t36 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t15 GNDA.t311 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X167 VDDA.t136 two_stage_opamp_dummy_magic_23_0.Vb3.t12 two_stage_opamp_dummy_magic_23_0.VD4.t12 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X168 VOUT-.t42 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT-.t43 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT+.t37 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VDDA.t472 GNDA.t525 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t5 VDDA.t353 VDDA.t355 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X173 VDDA.t473 GNDA.t526 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 VOUT+.t38 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VDDA.t474 GNDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 bgr_11_0.START_UP.t5 VDDA.t475 w_7200_15600.t29 w_7200_15600.t28 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X177 VOUT+.t39 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 two_stage_opamp_dummy_magic_23_0.X.t20 two_stage_opamp_dummy_magic_23_0.VD3.t35 two_stage_opamp_dummy_magic_23_0.VD3.t37 two_stage_opamp_dummy_magic_23_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X179 VDDA.t476 GNDA.t307 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VOUT+.t40 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT+.t41 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT-.t44 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 VOUT+.t42 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 VDDA.t477 GNDA.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 VDDA.t478 GNDA.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VDDA.t479 GNDA.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 a_5700_24908.t1 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t6 GNDA.t41 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X188 two_stage_opamp_dummy_magic_23_0.VD3.t29 two_stage_opamp_dummy_magic_23_0.Vb2.t13 two_stage_opamp_dummy_magic_23_0.X.t1 two_stage_opamp_dummy_magic_23_0.VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X189 VOUT+.t14 two_stage_opamp_dummy_magic_23_0.Y.t30 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X190 VOUT-.t45 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_11_0.Vin+.t5 VDDA.t480 w_7200_15600.t27 w_7200_15600.t26 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X192 w_6100_17280.t49 bgr_11_0.V_mir2.t13 VDDA.t57 w_6100_17280.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X193 VDDA.t481 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 VOUT-.t46 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT+.t43 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VDDA.t482 GNDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_11_0.V_mir1.t12 bgr_11_0.Vin-.t8 VDDA.t28 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X198 VDDA.t483 GNDA.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 two_stage_opamp_dummy_magic_23_0.VD2.t14 VIN+.t1 two_stage_opamp_dummy_magic_23_0.V_source.t11 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X200 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_23_0.X.t29 VDDA.t73 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X201 VDDA.t348 VDDA.t349 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_23_0.Y.t31 GNDA.t241 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X203 two_stage_opamp_dummy_magic_23_0.VD2.t18 VIN+.t2 two_stage_opamp_dummy_magic_23_0.V_source.t19 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X204 two_stage_opamp_dummy_magic_23_0.V_p_mir.t0 VIN+.t3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t0 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X205 VOUT+.t44 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT+.t45 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VDDA.t484 GNDA.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VDDA.t352 VDDA.t350 two_stage_opamp_dummy_magic_23_0.VD4.t17 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X209 a_7460_6300.t17 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_23_0.V_err_gate.t5 VDDA.t421 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X210 VDDA.t485 GNDA.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 VOUT-.t47 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VDDA.t486 GNDA.t145 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT+.t46 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VDDA.t347 VDDA.t344 VDDA.t346 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X215 GNDA.t63 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_23_0.V_source.t35 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X216 VDDA.t487 GNDA.t146 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 a_6350_25058.t1 bgr_11_0.Vin+.t1 GNDA.t165 sky130_fd_pr__res_xhigh_po_0p35 l=6
X218 a_8260_1600.t3 two_stage_opamp_dummy_magic_23_0.Vb1.t4 two_stage_opamp_dummy_magic_23_0.Vb1.t5 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X219 VDDA.t488 GNDA.t147 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_23_0.X.t30 GNDA.t304 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X221 VOUT-.t48 two_stage_opamp_dummy_magic_23_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT+.t47 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT-.t49 two_stage_opamp_dummy_magic_23_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 two_stage_opamp_dummy_magic_23_0.VD3.t11 VDDA.t339 VDDA.t341 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X225 VDDA.t489 GNDA.t185 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VDDA.t490 GNDA.t186 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT-.t50 two_stage_opamp_dummy_magic_23_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VDDA.t491 GNDA.t187 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 bgr_11_0.V_mir2.t11 bgr_11_0.V_mir2.t10 w_6100_17280.t31 w_6100_17280.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X230 w_7200_15600.t25 VDDA.t492 bgr_11_0.Vin-.t7 w_7200_15600.t24 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X231 VDDA.t169 two_stage_opamp_dummy_magic_23_0.Y.t32 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t12 GNDA.t587 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X232 VOUT-.t51 two_stage_opamp_dummy_magic_23_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VDDA.t493 GNDA.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT-.t52 two_stage_opamp_dummy_magic_23_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VOUT-.t53 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VOUT-.t54 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VDDA.t494 GNDA.t248 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 VDDA.t78 two_stage_opamp_dummy_magic_23_0.X.t31 VOUT-.t7 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X239 GNDA.t237 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_23_0.Vb3.t3 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X240 VDDA.t303 VDDA.t304 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VDDA.t495 GNDA.t168 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 GNDA.t316 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t14 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X243 VOUT-.t55 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT+.t48 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT+.t49 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VOUT+.t50 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 VOUT+.t51 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 VDDA.t418 two_stage_opamp_dummy_magic_23_0.V_err_gate.t18 two_stage_opamp_dummy_magic_23_0.V_err_p.t21 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X249 two_stage_opamp_dummy_magic_23_0.Y.t7 two_stage_opamp_dummy_magic_23_0.Vb1.t18 two_stage_opamp_dummy_magic_23_0.VD2.t8 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X250 VDDA.t496 GNDA.t169 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VDDA.t497 GNDA.t170 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 two_stage_opamp_dummy_magic_23_0.Y.t8 two_stage_opamp_dummy_magic_23_0.Vb1.t19 two_stage_opamp_dummy_magic_23_0.VD2.t7 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X253 VDDA.t498 GNDA.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VOUT+.t52 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 two_stage_opamp_dummy_magic_23_0.V_source.t34 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t17 GNDA.t320 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X256 two_stage_opamp_dummy_magic_23_0.VD3.t27 two_stage_opamp_dummy_magic_23_0.Vb2.t14 two_stage_opamp_dummy_magic_23_0.X.t2 two_stage_opamp_dummy_magic_23_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X257 GNDA.t444 GNDA.t442 VOUT+.t6 GNDA.t443 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X258 GNDA.t366 GNDA.t365 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X259 VDDA.t499 GNDA.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 VOUT-.t56 two_stage_opamp_dummy_magic_23_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 two_stage_opamp_dummy_magic_23_0.VD3.t8 two_stage_opamp_dummy_magic_23_0.Vb3.t13 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X262 VDDA.t500 GNDA.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 VDDA.t338 VDDA.t336 bgr_11_0.V_CMFB_S3.t5 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X264 two_stage_opamp_dummy_magic_23_0.VD4.t11 two_stage_opamp_dummy_magic_23_0.Vb3.t14 VDDA.t132 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X265 VDDA.t501 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VDDA.t502 GNDA.t209 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 bgr_11_0.V_CMFB_S3.t4 VDDA.t333 VDDA.t335 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X268 VOUT-.t57 two_stage_opamp_dummy_magic_23_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 w_7200_15600.t23 VDDA.t503 bgr_11_0.Vin+.t4 w_7200_15600.t22 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X270 VOUT-.t58 two_stage_opamp_dummy_magic_23_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 VDDA.t504 GNDA.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X273 w_6100_17280.t21 bgr_11_0.V_mir1.t14 bgr_11_0.1st_Vout_1.t5 w_6100_17280.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X274 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_23_0.Y.t33 VDDA.t174 GNDA.t588 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X275 VDDA.t505 GNDA.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 VDDA.t506 GNDA.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VOUT+.t53 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VDDA.t507 GNDA.t494 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 bgr_11_0.V_p_2.t2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t10 bgr_11_0.V_mir2.t12 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X280 VOUT+.t54 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 bgr_11_0.cap_res1.t0 VDDA.t52 GNDA.t229 sky130_fd_pr__res_high_po_0p35 l=2.05
X282 VOUT+.t55 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VOUT+.t56 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t11 two_stage_opamp_dummy_magic_23_0.X.t32 VDDA.t8 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X285 VDDA.t508 GNDA.t495 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 a_7460_6300.t8 two_stage_opamp_dummy_magic_23_0.V_err_gate.t19 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X287 a_7460_6300.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t20 VDDA.t82 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X288 two_stage_opamp_dummy_magic_23_0.VD2.t13 VIN+.t4 two_stage_opamp_dummy_magic_23_0.V_source.t10 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X289 VDDA.t509 GNDA.t496 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 a_7460_6300.t16 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_23_0.V_err_gate.t9 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X291 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_23_0.Y.t34 GNDA.t238 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X292 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_23_0.X.t33 VDDA.t9 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X293 VOUT+.t57 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 GNDA.t259 bgr_11_0.NFET_GATE_10uA.t9 two_stage_opamp_dummy_magic_23_0.Vb2.t6 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X295 VDDA.t332 VDDA.t330 GNDA.t540 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X296 VDDA.t510 GNDA.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 VDDA.t511 GNDA.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VDDA.t512 GNDA.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 two_stage_opamp_dummy_magic_23_0.Vb2.t5 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t261 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X300 VDDA.t513 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT-.t59 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 VDDA.t514 GNDA.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 bgr_11_0.Vin+.t3 VDDA.t515 w_7200_15600.t21 w_7200_15600.t20 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X304 a_8260_1600.t2 two_stage_opamp_dummy_magic_23_0.Vb1.t6 two_stage_opamp_dummy_magic_23_0.Vb1.t7 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X305 VOUT+.t58 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 VDDA.t32 bgr_11_0.V_mir2.t14 w_6100_17280.t33 w_6100_17280.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 w_6100_17280.t57 bgr_11_0.1st_Vout_1.t12 VDDA.t51 w_6100_17280.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X308 VOUT-.t4 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t2 GNDA.t219 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X309 VOUT-.t60 two_stage_opamp_dummy_magic_23_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VDDA.t329 VDDA.t327 VDDA.t329 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X311 VDDA.t516 GNDA.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VDDA.t326 VDDA.t324 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t10 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X313 VDDA.t517 GNDA.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VOUT+.t59 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VDDA.t518 GNDA.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 w_6100_17280.t19 bgr_11_0.V_mir1.t15 bgr_11_0.1st_Vout_1.t2 w_6100_17280.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X317 VDDA.t519 GNDA.t547 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VDDA.t101 GNDA.t439 GNDA.t441 GNDA.t440 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X319 bgr_11_0.1st_Vout_1.t13 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT+.t60 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VOUT-.t61 two_stage_opamp_dummy_magic_23_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT+.t61 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VDDA.t520 GNDA.t548 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 VDDA.t521 GNDA.t549 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VDDA.t522 GNDA.t182 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 two_stage_opamp_dummy_magic_23_0.Vb3.t1 two_stage_opamp_dummy_magic_23_0.Vb2.t15 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X327 VDDA.t39 two_stage_opamp_dummy_magic_23_0.X.t34 VOUT-.t1 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X328 a_4200_4468.t1 two_stage_opamp_dummy_magic_23_0.V_tot.t0 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X329 VOUT+.t62 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 bgr_11_0.NFET_GATE_10uA.t1 bgr_11_0.NFET_GATE_10uA.t0 GNDA.t251 GNDA.t250 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X331 two_stage_opamp_dummy_magic_23_0.VD4.t10 two_stage_opamp_dummy_magic_23_0.Vb3.t15 VDDA.t130 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X332 GNDA.t31 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t18 two_stage_opamp_dummy_magic_23_0.err_amp_out.t0 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X333 bgr_11_0.V_CMFB_S1.t5 VDDA.t321 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X334 VDDA.t523 GNDA.t183 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 VDDA.t70 two_stage_opamp_dummy_magic_23_0.V_err_gate.t21 a_7460_6300.t6 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X336 two_stage_opamp_dummy_magic_23_0.Y.t12 two_stage_opamp_dummy_magic_23_0.Vb1.t20 two_stage_opamp_dummy_magic_23_0.VD2.t6 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X337 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_11_0.Vin+.t0 GNDA.t257 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X339 VOUT-.t0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t3 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X340 VOUT+.t63 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VDDA.t524 GNDA.t184 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 two_stage_opamp_dummy_magic_23_0.VD3.t25 two_stage_opamp_dummy_magic_23_0.Vb2.t16 two_stage_opamp_dummy_magic_23_0.X.t18 two_stage_opamp_dummy_magic_23_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X343 two_stage_opamp_dummy_magic_23_0.V_source.t33 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t18 GNDA.t584 GNDA.t583 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X344 VDDA.t525 GNDA.t490 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 two_stage_opamp_dummy_magic_23_0.X.t19 two_stage_opamp_dummy_magic_23_0.Vb2.t17 two_stage_opamp_dummy_magic_23_0.VD3.t23 two_stage_opamp_dummy_magic_23_0.VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X346 VOUT+.t5 GNDA.t436 GNDA.t438 GNDA.t437 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X347 VDDA.t526 GNDA.t491 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT-.t62 two_stage_opamp_dummy_magic_23_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VDDA.t527 GNDA.t492 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VOUT-.t63 two_stage_opamp_dummy_magic_23_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VOUT+.t13 two_stage_opamp_dummy_magic_23_0.Y.t35 VDDA.t172 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X352 VOUT+.t64 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 VOUT-.t64 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 bgr_11_0.V_mir2.t9 bgr_11_0.V_mir2.t8 w_6100_17280.t29 w_6100_17280.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X355 two_stage_opamp_dummy_magic_23_0.VD4.t35 two_stage_opamp_dummy_magic_23_0.Vb2.t18 two_stage_opamp_dummy_magic_23_0.Y.t15 two_stage_opamp_dummy_magic_23_0.VD4.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X356 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_23_0.Y.t36 VDDA.t170 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X357 VDDA.t528 GNDA.t487 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 VOUT+.t65 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT+.t66 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 a_11420_25058.t1 bgr_11_0.Vin-.t2 GNDA.t249 sky130_fd_pr__res_xhigh_po_0p35 l=6
X361 VDDA.t301 VDDA.t302 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 VOUT+.t67 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VDDA.t529 GNDA.t488 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VDDA.t530 GNDA.t489 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_23_0.X.t35 VDDA.t40 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X366 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 two_stage_opamp_dummy_magic_23_0.V_err_p.t0 two_stage_opamp_dummy_magic_23_0.V_err_gate.t22 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X368 two_stage_opamp_dummy_magic_23_0.VD2.t0 VIN+.t5 two_stage_opamp_dummy_magic_23_0.V_source.t0 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X369 VDDA.t531 GNDA.t483 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 a_7460_6300.t18 two_stage_opamp_dummy_magic_23_0.V_tot.t4 two_stage_opamp_dummy_magic_23_0.V_err_gate.t10 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X371 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_23_0.Y.t37 GNDA.t221 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X372 VOUT+.t1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t4 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X373 GNDA.t318 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_23_0.V_source.t32 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X374 VDDA.t299 VDDA.t300 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VOUT+.t68 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VOUT-.t65 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VDDA.t128 two_stage_opamp_dummy_magic_23_0.Vb3.t16 two_stage_opamp_dummy_magic_23_0.VD3.t7 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X378 VOUT-.t66 two_stage_opamp_dummy_magic_23_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 VDDA.t532 GNDA.t484 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 two_stage_opamp_dummy_magic_23_0.Vb2.t4 bgr_11_0.NFET_GATE_10uA.t11 GNDA.t577 GNDA.t576 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X381 VOUT-.t67 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VDDA.t533 GNDA.t485 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VOUT-.t68 two_stage_opamp_dummy_magic_23_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 VDDA.t534 GNDA.t480 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VDDA.t320 VDDA.t319 w_6100_17280.t73 w_6100_17280.t72 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X386 VDDA.t535 GNDA.t481 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t167 two_stage_opamp_dummy_magic_23_0.Y.t38 VOUT+.t12 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X388 VOUT-.t69 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VDDA.t536 GNDA.t482 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VDDA.t537 GNDA.t477 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 VDDA.t317 VDDA.t318 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VOUT+.t69 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 VDDA.t538 GNDA.t478 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t8 VDDA.t314 VDDA.t316 VDDA.t315 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X395 VOUT+.t70 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t1 bgr_11_0.NFET_GATE_10uA.t12 GNDA.t579 GNDA.t578 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X397 VDDA.t42 two_stage_opamp_dummy_magic_23_0.X.t36 VOUT-.t2 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X398 VDDA.t539 GNDA.t479 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 two_stage_opamp_dummy_magic_23_0.Y.t10 two_stage_opamp_dummy_magic_23_0.VD4.t3 two_stage_opamp_dummy_magic_23_0.VD4.t5 two_stage_opamp_dummy_magic_23_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X400 VDDA.t44 two_stage_opamp_dummy_magic_23_0.X.t37 VOUT-.t3 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X401 VDDA.t540 GNDA.t474 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VDDA.t541 GNDA.t475 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 VDDA.t297 VDDA.t298 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 GNDA.t256 a_11950_23700.t1 GNDA.t255 sky130_fd_pr__res_xhigh_po_0p35 l=4
X405 two_stage_opamp_dummy_magic_23_0.X.t17 two_stage_opamp_dummy_magic_23_0.Vb2.t19 two_stage_opamp_dummy_magic_23_0.VD3.t21 two_stage_opamp_dummy_magic_23_0.VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X406 VOUT-.t70 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VOUT+.t71 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 two_stage_opamp_dummy_magic_23_0.Y.t13 two_stage_opamp_dummy_magic_23_0.Vb1.t21 two_stage_opamp_dummy_magic_23_0.VD2.t5 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X409 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t0 a_4600_1446.t1 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X410 VDDA.t542 GNDA.t476 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VDDA.t126 two_stage_opamp_dummy_magic_23_0.Vb3.t17 two_stage_opamp_dummy_magic_23_0.VD3.t6 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X412 a_4080_4468.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t3 GNDA.t288 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X413 VDDA.t543 GNDA.t472 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VDDA.t313 VDDA.t311 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t9 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X415 VOUT-.t5 a_13130_1456.t1 GNDA.t274 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X416 VDDA.t544 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VOUT-.t71 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 two_stage_opamp_dummy_magic_23_0.V_source.t31 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t20 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X419 VDDA.t545 GNDA.t473 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VDDA.t546 GNDA.t160 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+.t72 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VOUT-.t72 two_stage_opamp_dummy_magic_23_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t8 VDDA.t308 VDDA.t310 VDDA.t309 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X424 GNDA.t366 GNDA.t432 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X425 GNDA.t348 two_stage_opamp_dummy_magic_23_0.X.t38 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t6 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X426 VOUT-.t73 two_stage_opamp_dummy_magic_23_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VDDA.t547 GNDA.t161 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VOUT+.t73 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 bgr_11_0.START_UP.t4 VDDA.t548 w_7200_15600.t19 w_7200_15600.t18 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X430 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VDDA.t549 GNDA.t279 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VOUT+.t74 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VDDA.t550 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VDDA.t551 GNDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT+.t75 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 VDDA.t552 GNDA.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VDDA.t419 bgr_11_0.V_mir2.t15 w_6100_17280.t81 w_6100_17280.t80 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X438 VOUT+.t18 VDDA.t305 VDDA.t307 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X439 two_stage_opamp_dummy_magic_23_0.cap_res_X.t0 two_stage_opamp_dummy_magic_23_0.X.t3 GNDA.t43 sky130_fd_pr__res_high_po_1p41 l=1.41
X440 VOUT+.t76 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_23_0.Y.t39 VDDA.t165 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X442 two_stage_opamp_dummy_magic_23_0.VD1.t16 VIN-.t2 two_stage_opamp_dummy_magic_23_0.V_source.t13 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X443 GNDA.t435 GNDA.t433 two_stage_opamp_dummy_magic_23_0.V_source.t20 GNDA.t434 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X444 GNDA.t431 GNDA.t428 GNDA.t430 GNDA.t429 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X445 GNDA.t427 GNDA.t425 VDDA.t100 GNDA.t426 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X446 VDDA.t553 GNDA.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 two_stage_opamp_dummy_magic_23_0.V_err_p.t11 two_stage_opamp_dummy_magic_23_0.V_tot.t5 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t2 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X448 VDDA.t554 GNDA.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 bgr_11_0.1st_Vout_1.t17 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 VDDA.t555 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 VOUT+.t77 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 two_stage_opamp_dummy_magic_23_0.err_amp_out.t1 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t19 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X453 VDDA.t556 GNDA.t158 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VOUT-.t74 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 GNDA.t337 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t5 VOUT-.t9 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X456 VOUT-.t75 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 two_stage_opamp_dummy_magic_23_0.VD2.t20 GNDA.t423 GNDA.t424 GNDA.t418 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X458 VOUT-.t76 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 VOUT+.t78 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 a_7460_6300.t5 two_stage_opamp_dummy_magic_23_0.V_err_gate.t23 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X461 VDDA.t557 GNDA.t159 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VDDA.t558 GNDA.t521 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 a_7460_6300.t15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_23_0.V_err_gate.t6 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X464 VDDA.t559 GNDA.t522 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 bgr_11_0.V_mir1.t1 bgr_11_0.V_mir1.t0 w_6100_17280.t17 w_6100_17280.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X466 GNDA.t422 GNDA.t421 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t3 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X467 two_stage_opamp_dummy_magic_23_0.VD1.t17 VIN-.t3 two_stage_opamp_dummy_magic_23_0.V_source.t16 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X468 GNDA.t366 GNDA.t420 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X469 two_stage_opamp_dummy_magic_23_0.V_err_p.t17 two_stage_opamp_dummy_magic_23_0.V_tot.t6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t3 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X470 VDDA.t393 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t1 w_7200_15600.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X471 VOUT+.t79 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT-.t77 two_stage_opamp_dummy_magic_23_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VOUT+.t80 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VOUT-.t78 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VDDA.t560 GNDA.t523 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 w_7200_15600.t39 w_7200_15600.t37 VDDA.t35 w_7200_15600.t38 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X477 VDDA.t561 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VDDA.t562 GNDA.t519 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VDDA.t563 GNDA.t520 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VDDA.t564 GNDA.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 two_stage_opamp_dummy_magic_23_0.Y.t21 two_stage_opamp_dummy_magic_23_0.Vb2.t20 two_stage_opamp_dummy_magic_23_0.VD4.t33 two_stage_opamp_dummy_magic_23_0.VD4.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X482 VOUT+.t81 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VDDA.t164 two_stage_opamp_dummy_magic_23_0.Y.t40 VOUT+.t11 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X484 VOUT+.t82 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VDDA.t565 GNDA.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 VDDA.t566 GNDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_23_0.Vb3.t4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X488 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 a_4200_4468.t0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t0 GNDA.t42 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X490 VDDA.t567 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 VOUT-.t79 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 two_stage_opamp_dummy_magic_23_0.X.t12 two_stage_opamp_dummy_magic_23_0.Vb1.t22 two_stage_opamp_dummy_magic_23_0.VD1.t6 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X493 VDDA.t568 GNDA.t180 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VOUT-.t80 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VDDA.t124 two_stage_opamp_dummy_magic_23_0.Vb3.t18 two_stage_opamp_dummy_magic_23_0.VD4.t9 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X496 VDDA.t98 two_stage_opamp_dummy_magic_23_0.X.t39 VOUT-.t10 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X497 VDDA.t295 VDDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 VDDA.t569 GNDA.t181 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VOUT-.t81 two_stage_opamp_dummy_magic_23_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 VOUT-.t82 two_stage_opamp_dummy_magic_23_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 bgr_11_0.NFET_GATE_10uA.t3 VDDA.t292 VDDA.t294 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X502 VOUT-.t83 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 VOUT-.t84 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 VDDA.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t24 a_7460_6300.t4 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X505 VDDA.t570 GNDA.t516 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 VDDA.t571 GNDA.t517 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 VOUT-.t85 two_stage_opamp_dummy_magic_23_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT+.t83 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 two_stage_opamp_dummy_magic_23_0.X.t21 two_stage_opamp_dummy_magic_23_0.Vb2.t21 two_stage_opamp_dummy_magic_23_0.VD3.t19 two_stage_opamp_dummy_magic_23_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X510 VDDA.t572 GNDA.t518 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT+.t84 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 w_7200_15600.t17 VDDA.t573 bgr_11_0.Vin+.t2 w_7200_15600.t16 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X513 two_stage_opamp_dummy_magic_23_0.Y.t24 GNDA.t417 GNDA.t419 GNDA.t418 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X514 two_stage_opamp_dummy_magic_23_0.V_p_mir.t3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t21 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X515 two_stage_opamp_dummy_magic_23_0.V_source.t30 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t22 GNDA.t591 GNDA.t590 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X516 VDDA.t574 GNDA.t514 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VOUT+.t85 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 GNDA.t366 GNDA.t367 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X519 two_stage_opamp_dummy_magic_23_0.X.t11 two_stage_opamp_dummy_magic_23_0.Vb1.t23 two_stage_opamp_dummy_magic_23_0.VD1.t5 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X520 VDDA.t575 GNDA.t515 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VDDA.t576 GNDA.t511 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VOUT-.t86 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VOUT-.t87 two_stage_opamp_dummy_magic_23_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 bgr_11_0.START_UP.t1 bgr_11_0.START_UP.t0 bgr_11_0.START_UP_NFET1.t0 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X525 VDDA.t285 VDDA.t284 w_6100_17280.t71 w_6100_17280.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X526 GNDA.t191 two_stage_opamp_dummy_magic_23_0.X.t40 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t5 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X527 GNDA.t282 a_11300_23450.t1 GNDA.t281 sky130_fd_pr__res_xhigh_po_0p35 l=6
X528 two_stage_opamp_dummy_magic_23_0.Y.t22 two_stage_opamp_dummy_magic_23_0.Vb2.t22 two_stage_opamp_dummy_magic_23_0.VD4.t31 two_stage_opamp_dummy_magic_23_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X529 VOUT-.t88 two_stage_opamp_dummy_magic_23_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT+.t86 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VDDA.t577 GNDA.t512 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VDDA.t578 GNDA.t513 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VOUT-.t89 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VDDA.t579 GNDA.t509 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 VDDA.t580 GNDA.t510 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 two_stage_opamp_dummy_magic_23_0.VD1.t18 VIN-.t4 two_stage_opamp_dummy_magic_23_0.V_source.t17 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X537 VDDA.t282 VDDA.t283 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_23_0.Y.t41 VDDA.t162 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X539 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t4 VDDA.t581 w_7200_15600.t15 w_7200_15600.t14 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X540 two_stage_opamp_dummy_magic_23_0.V_err_p.t16 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_23_0.err_amp_out.t6 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X541 VOUT-.t90 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VOUT+.t87 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VDDA.t582 GNDA.t504 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VDDA.t583 GNDA.t505 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VOUT+.t88 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VDDA.t280 VDDA.t281 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT-.t91 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 VDDA.t584 GNDA.t506 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 two_stage_opamp_dummy_magic_23_0.VD3.t5 two_stage_opamp_dummy_magic_23_0.Vb3.t19 VDDA.t122 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X550 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t11 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X551 VOUT+.t89 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 VDDA.t93 bgr_11_0.V_mir2.t16 w_6100_17280.t65 w_6100_17280.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X553 two_stage_opamp_dummy_magic_23_0.V_err_p.t10 two_stage_opamp_dummy_magic_23_0.V_err_gate.t25 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X554 VDDA.t3 bgr_11_0.1st_Vout_1.t19 w_6100_17280.t55 w_6100_17280.t54 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X555 VDDA.t585 GNDA.t499 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VDDA.t586 GNDA.t500 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 VDDA.t587 GNDA.t501 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 a_7460_6300.t12 two_stage_opamp_dummy_magic_23_0.V_tot.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t2 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X559 two_stage_opamp_dummy_magic_23_0.VD1.t12 VIN-.t5 two_stage_opamp_dummy_magic_23_0.V_source.t5 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X560 VDDA.t588 GNDA.t225 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 VDDA.t291 VDDA.t289 two_stage_opamp_dummy_magic_23_0.Vb1.t11 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X562 two_stage_opamp_dummy_magic_23_0.V_err_p.t14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_23_0.err_amp_out.t5 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X563 VOUT-.t92 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 VOUT+.t90 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 bgr_11_0.1st_Vout_1.t1 bgr_11_0.V_mir1.t16 w_6100_17280.t15 w_6100_17280.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X566 VOUT+.t91 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 VOUT-.t93 two_stage_opamp_dummy_magic_23_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 VOUT-.t94 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VDDA.t589 GNDA.t226 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VDDA.t120 two_stage_opamp_dummy_magic_23_0.Vb3.t20 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t7 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X571 VDDA.t590 GNDA.t227 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 VDDA.t161 two_stage_opamp_dummy_magic_23_0.Y.t42 VOUT+.t10 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X573 VDDA.t288 VDDA.t286 two_stage_opamp_dummy_magic_23_0.V_err_p.t19 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X574 two_stage_opamp_dummy_magic_23_0.X.t22 two_stage_opamp_dummy_magic_23_0.Vb2.t23 two_stage_opamp_dummy_magic_23_0.VD3.t17 two_stage_opamp_dummy_magic_23_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X575 VDDA.t279 VDDA.t277 VOUT+.t17 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X576 VOUT+.t92 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 w_7200_15600.t11 VDDA.t591 bgr_11_0.START_UP.t3 w_7200_15600.t10 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X578 GNDA.t416 GNDA.t415 two_stage_opamp_dummy_magic_23_0.VD1.t20 GNDA.t408 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X579 VDDA.t592 GNDA.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 two_stage_opamp_dummy_magic_23_0.VD4.t29 two_stage_opamp_dummy_magic_23_0.Vb2.t24 two_stage_opamp_dummy_magic_23_0.Y.t5 two_stage_opamp_dummy_magic_23_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X581 VOUT-.t95 two_stage_opamp_dummy_magic_23_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 VDDA.t593 GNDA.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 VOUT+.t93 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 VOUT+.t94 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 bgr_11_0.Vin-.t6 VDDA.t594 w_7200_15600.t13 w_7200_15600.t12 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X586 VOUT+.t95 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 VDDA.t595 GNDA.t242 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 VDDA.t596 GNDA.t243 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 GNDA.t414 GNDA.t412 two_stage_opamp_dummy_magic_23_0.Vb3.t5 GNDA.t413 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X590 two_stage_opamp_dummy_magic_23_0.VD3.t34 two_stage_opamp_dummy_magic_23_0.VD3.t32 two_stage_opamp_dummy_magic_23_0.X.t15 two_stage_opamp_dummy_magic_23_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X591 two_stage_opamp_dummy_magic_23_0.X.t10 two_stage_opamp_dummy_magic_23_0.Vb1.t24 two_stage_opamp_dummy_magic_23_0.VD1.t4 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X592 VDDA.t597 GNDA.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 VOUT+.t96 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 w_6100_17280.t44 w_6100_17280.t42 VDDA.t412 w_6100_17280.t43 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X595 VOUT+.t97 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 VOUT+.t0 a_4600_1446.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X597 VOUT+.t98 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 two_stage_opamp_dummy_magic_23_0.VD3.t4 two_stage_opamp_dummy_magic_23_0.Vb3.t21 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X599 VDDA.t37 two_stage_opamp_dummy_magic_23_0.X.t41 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t8 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X600 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t1 a_13130_1456.t0 GNDA.t228 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X601 GNDA.t411 GNDA.t410 two_stage_opamp_dummy_magic_23_0.VD2.t19 GNDA.t402 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X602 VDDA.t598 GNDA.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VDDA.t599 GNDA.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VOUT+.t99 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 VDDA.t600 GNDA.t175 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 two_stage_opamp_dummy_magic_23_0.V_source.t29 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t23 GNDA.t554 GNDA.t553 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X607 two_stage_opamp_dummy_magic_23_0.X.t9 two_stage_opamp_dummy_magic_23_0.Vb1.t25 two_stage_opamp_dummy_magic_23_0.VD1.t3 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X608 VOUT+.t100 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 bgr_11_0.V_mir2.t7 bgr_11_0.V_mir2.t6 w_6100_17280.t63 w_6100_17280.t62 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X610 two_stage_opamp_dummy_magic_23_0.V_source.t2 two_stage_opamp_dummy_magic_23_0.Vb1.t26 a_8260_1600.t4 GNDA.t278 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X611 VOUT-.t96 two_stage_opamp_dummy_magic_23_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VDDA.t601 GNDA.t176 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VDDA.t276 VDDA.t274 bgr_11_0.V_CMFB_S3.t3 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X614 GNDA.t497 two_stage_opamp_dummy_magic_23_0.X.t42 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t4 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X615 VDDA.t602 GNDA.t177 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 bgr_11_0.V_CMFB_S3.t2 VDDA.t271 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X617 VOUT-.t97 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 VDDA.t603 GNDA.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 VOUT-.t98 two_stage_opamp_dummy_magic_23_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VOUT-.t99 two_stage_opamp_dummy_magic_23_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 bgr_11_0.1st_Vout_1.t20 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VOUT+.t101 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 VOUT+.t102 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 VDDA.t604 GNDA.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VDDA.t605 GNDA.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 VDDA.t606 GNDA.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 a_5700_24908.t0 a_5820_23644.t0 GNDA.t41 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X628 GNDA.t409 GNDA.t407 two_stage_opamp_dummy_magic_23_0.X.t24 GNDA.t408 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X629 VOUT+.t103 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 VOUT+.t104 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VOUT+.t105 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 bgr_11_0.1st_Vout_1.t0 bgr_11_0.V_mir1.t17 w_6100_17280.t13 w_6100_17280.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X633 VDDA.t607 GNDA.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 VDDA.t608 GNDA.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 VDDA.t609 GNDA.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 two_stage_opamp_dummy_magic_23_0.V_err_p.t18 VDDA.t268 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X638 two_stage_opamp_dummy_magic_23_0.V_err_p.t9 two_stage_opamp_dummy_magic_23_0.V_err_gate.t26 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X639 two_stage_opamp_dummy_magic_23_0.err_amp_out.t2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t20 GNDA.t119 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X640 GNDA.t406 GNDA.t404 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t3 GNDA.t405 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X641 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_23_0.Y.t43 GNDA.t267 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X642 GNDA.t403 GNDA.t401 two_stage_opamp_dummy_magic_23_0.Y.t23 GNDA.t402 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X643 VOUT-.t100 two_stage_opamp_dummy_magic_23_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 two_stage_opamp_dummy_magic_23_0.VD4.t16 VDDA.t265 VDDA.t267 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X645 two_stage_opamp_dummy_magic_23_0.VD1.t19 GNDA.t399 GNDA.t400 GNDA.t394 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X646 VOUT-.t101 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 VOUT-.t102 two_stage_opamp_dummy_magic_23_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 VOUT+.t106 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 GNDA.t366 GNDA.t398 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X650 GNDA.t65 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t3 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X651 two_stage_opamp_dummy_magic_23_0.VD4.t27 two_stage_opamp_dummy_magic_23_0.Vb2.t25 two_stage_opamp_dummy_magic_23_0.Y.t6 two_stage_opamp_dummy_magic_23_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X652 two_stage_opamp_dummy_magic_23_0.V_err_p.t2 two_stage_opamp_dummy_magic_23_0.V_tot.t8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X653 VOUT+.t107 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 VDDA.t610 GNDA.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 VDDA.t611 GNDA.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 a_6350_25058.t0 a_6470_23450.t1 GNDA.t165 sky130_fd_pr__res_xhigh_po_0p35 l=6
X657 VOUT+.t108 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VDDA.t264 VDDA.t262 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t7 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X660 a_4080_4468.t1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t14 GNDA.t589 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X661 VDDA.t612 GNDA.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 VDDA.t613 GNDA.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t6 VDDA.t259 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X664 two_stage_opamp_dummy_magic_23_0.VD3.t3 two_stage_opamp_dummy_magic_23_0.Vb3.t22 VDDA.t116 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X665 a_13450_4368.t1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t0 GNDA.t151 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X666 VDDA.t614 GNDA.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 VDDA.t29 bgr_11_0.1st_Vout_1.t23 w_6100_17280.t53 w_6100_17280.t52 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X668 VDDA.t158 two_stage_opamp_dummy_magic_23_0.Y.t44 VOUT+.t9 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X669 VDDA.t257 VDDA.t258 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 VOUT+.t109 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 two_stage_opamp_dummy_magic_23_0.err_amp_out.t4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_23_0.V_err_p.t15 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X672 VDDA.t615 GNDA.t204 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_23_0.VD3.t15 two_stage_opamp_dummy_magic_23_0.Vb2.t26 two_stage_opamp_dummy_magic_23_0.X.t0 two_stage_opamp_dummy_magic_23_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X675 VDDA.t616 GNDA.t205 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 VDDA.t617 GNDA.t206 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 GNDA.t67 bgr_11_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_23_0.V_err_gate.t3 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X678 bgr_11_0.V_CMFB_S1.t4 VDDA.t254 VDDA.t256 VDDA.t255 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X679 GNDA.t231 two_stage_opamp_dummy_magic_23_0.Y.t45 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t4 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X680 VDDA.t407 two_stage_opamp_dummy_magic_23_0.X.t43 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t7 GNDA.t498 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X681 bgr_11_0.cap_res2.t20 VDDA.t423 GNDA.t594 sky130_fd_pr__res_high_po_0p35 l=2.05
X682 VDDA.t253 VDDA.t251 bgr_11_0.V_CMFB_S1.t3 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X683 two_stage_opamp_dummy_magic_23_0.V_source.t3 VIN+.t6 two_stage_opamp_dummy_magic_23_0.VD2.t11 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X684 VOUT-.t103 two_stage_opamp_dummy_magic_23_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VOUT+.t110 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 VDDA.t411 bgr_11_0.1st_Vout_1.t25 w_6100_17280.t51 w_6100_17280.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X687 VDDA.t250 VDDA.t248 bgr_11_0.V_CMFB_S1.t2 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X688 VDDA.t618 GNDA.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 two_stage_opamp_dummy_magic_23_0.V_err_gate.t13 two_stage_opamp_dummy_magic_23_0.V_tot.t9 a_7460_6300.t19 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X690 VOUT-.t104 two_stage_opamp_dummy_magic_23_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 VOUT-.t105 two_stage_opamp_dummy_magic_23_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 VDDA.t619 GNDA.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 GNDA.t366 GNDA.t397 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X694 two_stage_opamp_dummy_magic_23_0.VD4.t25 two_stage_opamp_dummy_magic_23_0.Vb2.t27 two_stage_opamp_dummy_magic_23_0.Y.t2 two_stage_opamp_dummy_magic_23_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X695 two_stage_opamp_dummy_magic_23_0.V_source.t28 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t24 GNDA.t124 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X696 GNDA.t366 GNDA.t396 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X697 two_stage_opamp_dummy_magic_23_0.X.t23 GNDA.t393 GNDA.t395 GNDA.t394 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X698 two_stage_opamp_dummy_magic_23_0.Vb1.t1 two_stage_opamp_dummy_magic_23_0.Vb1.t0 a_8260_1600.t1 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X699 GNDA.t346 two_stage_opamp_dummy_magic_23_0.X.t44 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t3 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X700 VOUT+.t111 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 GNDA.t347 two_stage_opamp_dummy_magic_23_0.X.t45 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t2 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X702 VDDA.t620 GNDA.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 VDDA.t621 GNDA.t356 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 VDDA.t622 GNDA.t357 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 VDDA.t239 VDDA.t240 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 VDDA.t623 GNDA.t358 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 VOUT-.t106 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT+.t112 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 two_stage_opamp_dummy_magic_23_0.Vb3.t0 bgr_11_0.NFET_GATE_10uA.t15 GNDA.t14 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X710 VDDA.t624 GNDA.t354 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 VDDA.t625 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 VDDA.t626 GNDA.t355 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 VDDA.t247 VDDA.t244 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X714 bgr_11_0.V_mir1.t7 bgr_11_0.V_mir1.t6 w_6100_17280.t11 w_6100_17280.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X715 VDDA.t114 two_stage_opamp_dummy_magic_23_0.Vb3.t23 two_stage_opamp_dummy_magic_23_0.VD3.t2 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X716 VOUT-.t17 two_stage_opamp_dummy_magic_23_0.X.t46 VDDA.t404 VDDA.t403 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X717 VDDA.t627 GNDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 VOUT-.t107 two_stage_opamp_dummy_magic_23_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 VDDA.t416 w_6100_17280.t39 w_6100_17280.t41 w_6100_17280.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X720 a_7460_6300.t3 two_stage_opamp_dummy_magic_23_0.V_err_gate.t27 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X721 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t9 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X722 VDDA.t628 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 VDDA.t629 GNDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VOUT-.t108 two_stage_opamp_dummy_magic_23_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VDDA.t630 GNDA.t351 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 two_stage_opamp_dummy_magic_23_0.VD2.t4 two_stage_opamp_dummy_magic_23_0.Vb1.t27 two_stage_opamp_dummy_magic_23_0.Y.t11 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X727 GNDA.t263 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_23_0.V_source.t27 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X728 GNDA.t272 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_23_0.V_source.t26 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X729 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t2 bgr_11_0.NFET_GATE_10uA.t16 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X730 VDDA.t631 GNDA.t352 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 GNDA.t153 bgr_11_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t1 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X732 VDDA.t243 VDDA.t241 VDDA.t243 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X733 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 VDDA.t632 GNDA.t353 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 VDDA.t633 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 VOUT+.t113 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VDDA.t634 GNDA.t467 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 a_12070_24908.t0 a_11950_23700.t0 GNDA.t156 sky130_fd_pr__res_xhigh_po_0p35 l=4
X739 two_stage_opamp_dummy_magic_23_0.VD3.t13 two_stage_opamp_dummy_magic_23_0.Vb2.t28 two_stage_opamp_dummy_magic_23_0.X.t16 two_stage_opamp_dummy_magic_23_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X740 VOUT-.t109 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 VOUT+.t114 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 VOUT+.t115 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 w_6100_17280.t1 bgr_11_0.V_mir2.t17 VDDA.t0 w_6100_17280.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X744 VDDA.t635 GNDA.t468 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VDDA.t636 GNDA.t286 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 two_stage_opamp_dummy_magic_23_0.Vb2.t3 bgr_11_0.NFET_GATE_10uA.t18 GNDA.t155 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X748 bgr_11_0.V_mir1.t5 bgr_11_0.V_mir1.t4 w_6100_17280.t9 w_6100_17280.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X749 w_7200_15600.t9 VDDA.t637 bgr_11_0.START_UP.t2 w_7200_15600.t8 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X750 VDDA.t112 two_stage_opamp_dummy_magic_23_0.Vb3.t24 two_stage_opamp_dummy_magic_23_0.VD3.t1 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X751 VDDA.t638 GNDA.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VOUT-.t110 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 GNDA.t215 bgr_11_0.NFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_23_0.Vb2.t2 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X754 VDDA.t639 GNDA.t349 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VOUT-.t111 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 two_stage_opamp_dummy_magic_23_0.Vb2.t0 two_stage_opamp_dummy_magic_23_0.Vb2_2.t0 two_stage_opamp_dummy_magic_23_0.Vb2_2.t2 two_stage_opamp_dummy_magic_23_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X757 VOUT-.t112 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VOUT+.t3 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t6 GNDA.t291 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X759 VDDA.t640 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VDDA.t641 GNDA.t350 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 VOUT-.t113 two_stage_opamp_dummy_magic_23_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 VOUT-.t114 two_stage_opamp_dummy_magic_23_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 VDDA.t71 w_6100_17280.t36 w_6100_17280.t38 w_6100_17280.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X764 two_stage_opamp_dummy_magic_23_0.V_source.t18 VIN+.t7 two_stage_opamp_dummy_magic_23_0.VD2.t17 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X765 VDDA.t405 two_stage_opamp_dummy_magic_23_0.X.t47 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t6 GNDA.t493 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X766 VOUT-.t115 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 two_stage_opamp_dummy_magic_23_0.V_err_gate.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t10 a_7460_6300.t0 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X768 GNDA.t265 two_stage_opamp_dummy_magic_23_0.Y.t46 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t3 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X769 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t2 GNDA.t391 GNDA.t392 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X770 VOUT+.t116 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 VOUT+.t117 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 two_stage_opamp_dummy_magic_23_0.V_err_gate.t7 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t16 a_7460_6300.t14 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X773 VDDA.t642 GNDA.t464 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 VDDA.t643 GNDA.t465 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 VOUT+.t118 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t5 VDDA.t236 VDDA.t238 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X777 bgr_11_0.1st_Vout_1.t28 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 VDDA.t644 GNDA.t466 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 two_stage_opamp_dummy_magic_23_0.V_source.t25 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t27 GNDA.t593 GNDA.t592 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X780 VDDA.t645 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 VDDA.t646 GNDA.t293 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 two_stage_opamp_dummy_magic_23_0.Vb1.t3 two_stage_opamp_dummy_magic_23_0.Vb1.t2 a_8260_1600.t0 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X783 VDDA.t647 GNDA.t294 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 GNDA.t239 VDDA.t233 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X785 VOUT+.t119 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 VOUT-.t116 two_stage_opamp_dummy_magic_23_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 VDDA.t232 VDDA.t230 two_stage_opamp_dummy_magic_23_0.Vb2_2.t6 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X788 VOUT-.t117 two_stage_opamp_dummy_magic_23_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X789 VDDA.t648 GNDA.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 VDDA.t649 GNDA.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 bgr_11_0.1st_Vout_1.t29 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X792 VDDA.t650 GNDA.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 VOUT-.t118 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X794 VDDA.t651 GNDA.t561 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X795 VDDA.t652 GNDA.t562 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 VDDA.t653 GNDA.t563 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X797 VDDA.t61 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t6 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X798 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_23_0.Y.t47 VDDA.t153 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X799 VOUT-.t119 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X800 w_6100_17280.t3 bgr_11_0.V_mir2.t4 bgr_11_0.V_mir2.t5 w_6100_17280.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X801 VDDA.t654 GNDA.t573 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X802 VDDA.t655 GNDA.t574 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X803 VOUT-.t120 two_stage_opamp_dummy_magic_23_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X804 VOUT-.t8 two_stage_opamp_dummy_magic_23_0.X.t48 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X805 VOUT+.t120 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X806 VOUT+.t121 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X807 VOUT+.t122 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X808 VDDA.t110 two_stage_opamp_dummy_magic_23_0.Vb3.t25 two_stage_opamp_dummy_magic_23_0.VD4.t8 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X809 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t7 GNDA.t552 GNDA.t551 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X810 VDDA.t656 GNDA.t575 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X811 VOUT+.t123 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 two_stage_opamp_dummy_magic_23_0.Y.t14 two_stage_opamp_dummy_magic_23_0.Vb2.t29 two_stage_opamp_dummy_magic_23_0.VD4.t23 two_stage_opamp_dummy_magic_23_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X813 two_stage_opamp_dummy_magic_23_0.V_err_p.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t28 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X814 two_stage_opamp_dummy_magic_23_0.VD2.t3 two_stage_opamp_dummy_magic_23_0.Vb1.t28 two_stage_opamp_dummy_magic_23_0.Y.t17 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X815 VOUT-.t121 two_stage_opamp_dummy_magic_23_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X816 VDDA.t657 GNDA.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X817 VDDA.t658 GNDA.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X818 VDDA.t659 GNDA.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X819 VDDA.t660 GNDA.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X820 GNDA.t269 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_23_0.V_source.t24 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X821 VOUT-.t122 two_stage_opamp_dummy_magic_23_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X822 bgr_11_0.Vin-.t0 bgr_11_0.START_UP.t7 VDDA.t395 w_7200_15600.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X823 VOUT-.t123 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X824 VOUT+.t124 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X825 VDDA.t661 GNDA.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X826 VDDA.t662 GNDA.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X827 VDDA.t229 VDDA.t227 two_stage_opamp_dummy_magic_23_0.VD3.t10 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X828 a_13570_4368.t1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t0 GNDA.t230 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X829 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t5 VDDA.t663 w_7200_15600.t7 w_7200_15600.t6 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X830 VDDA.t217 VDDA.t218 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X831 VDDA.t664 GNDA.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X832 VOUT-.t124 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X833 VOUT-.t125 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X834 VDDA.t665 GNDA.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X835 VOUT-.t126 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X836 w_6100_17280.t69 VDDA.t222 VDDA.t223 w_6100_17280.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X837 VOUT+.t125 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X838 VDDA.t154 two_stage_opamp_dummy_magic_23_0.Y.t48 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t6 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X839 VDDA.t666 GNDA.t343 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X840 VOUT-.t127 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X841 VDDA.t667 GNDA.t344 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X842 VDDA.t668 GNDA.t345 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X843 VDDA.t215 VDDA.t216 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X844 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t224 VDDA.t226 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X845 GNDA.t298 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t7 VOUT-.t6 GNDA.t297 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X846 VOUT+.t126 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X847 VOUT+.t127 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X848 VOUT+.t128 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X849 VDDA.t669 GNDA.t148 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X850 VOUT+.t129 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X851 VOUT-.t128 two_stage_opamp_dummy_magic_23_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X852 VDDA.t221 VDDA.t219 bgr_11_0.V_CUR_REF_REG.t1 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X853 VDDA.t91 two_stage_opamp_dummy_magic_23_0.X.t49 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t5 GNDA.t335 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X854 VOUT+.t130 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X855 VDDA.t20 two_stage_opamp_dummy_magic_23_0.V_err_gate.t29 two_stage_opamp_dummy_magic_23_0.V_err_p.t4 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X856 two_stage_opamp_dummy_magic_23_0.V_source.t7 VIN+.t8 two_stage_opamp_dummy_magic_23_0.VD2.t12 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X857 VDDA.t670 GNDA.t149 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X858 VDDA.t671 GNDA.t150 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X859 VDDA.t18 two_stage_opamp_dummy_magic_23_0.V_err_gate.t30 two_stage_opamp_dummy_magic_23_0.V_err_p.t3 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X860 VDDA.t408 two_stage_opamp_dummy_magic_23_0.X.t50 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t4 GNDA.t550 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X861 VOUT-.t129 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X862 two_stage_opamp_dummy_magic_23_0.Y.t4 two_stage_opamp_dummy_magic_23_0.Vb2.t30 two_stage_opamp_dummy_magic_23_0.VD4.t21 two_stage_opamp_dummy_magic_23_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X863 two_stage_opamp_dummy_magic_23_0.V_err_gate.t8 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t17 a_7460_6300.t13 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X864 w_7200_15600.t36 w_7200_15600.t34 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t0 w_7200_15600.t35 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X865 GNDA.t327 two_stage_opamp_dummy_magic_23_0.Y.t49 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t2 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X866 VOUT-.t130 two_stage_opamp_dummy_magic_23_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X867 VDDA.t672 GNDA.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X868 VOUT-.t131 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X869 VOUT+.t131 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X870 two_stage_opamp_dummy_magic_23_0.Vb1.t8 GNDA.t388 GNDA.t390 GNDA.t389 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X871 VOUT-.t132 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X872 VDDA.t673 GNDA.t189 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X873 VDDA.t674 GNDA.t190 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X874 VDDA.t675 GNDA.t558 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X875 VOUT+.t132 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X876 GNDA.t96 a_6520_18930# VDDA.t27 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X877 GNDA.t387 GNDA.t385 VOUT-.t12 GNDA.t386 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X878 VOUT-.t133 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X879 bgr_11_0.1st_Vout_1.t3 bgr_11_0.V_mir1.t18 w_6100_17280.t7 w_6100_17280.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X880 VDDA.t676 GNDA.t559 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X881 VOUT-.t134 two_stage_opamp_dummy_magic_23_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X882 VOUT-.t135 two_stage_opamp_dummy_magic_23_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X883 VDDA.t677 GNDA.t560 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X884 two_stage_opamp_dummy_magic_23_0.Vb2_2.t9 two_stage_opamp_dummy_magic_23_0.Vb2.t31 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X885 VOUT+.t133 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X886 two_stage_opamp_dummy_magic_23_0.VD3.t0 two_stage_opamp_dummy_magic_23_0.Vb3.t26 VDDA.t108 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X887 VDDA.t213 VDDA.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X888 VDDA.t678 GNDA.t570 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X889 VOUT+.t134 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X890 VOUT+.t135 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X891 GNDA.t322 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t8 VOUT+.t4 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X892 VOUT+.t136 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X893 VOUT+.t137 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X894 VOUT-.t136 two_stage_opamp_dummy_magic_23_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X895 VDDA.t679 GNDA.t571 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X896 VOUT-.t18 two_stage_opamp_dummy_magic_23_0.X.t51 VDDA.t410 VDDA.t409 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X897 VDDA.t680 GNDA.t572 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X898 VDDA.t681 GNDA.t341 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X899 VDDA.t26 a_6520_18930# GNDA.t94 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X900 a_13450_4368.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t1 GNDA.t47 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X901 two_stage_opamp_dummy_magic_23_0.err_amp_out.t10 GNDA.t382 GNDA.t384 GNDA.t383 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X902 w_7200_15600.t3 VDDA.t682 bgr_11_0.Vin-.t5 w_7200_15600.t2 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X903 VOUT-.t137 two_stage_opamp_dummy_magic_23_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X904 a_7460_6300.t2 two_stage_opamp_dummy_magic_23_0.V_err_gate.t31 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X905 two_stage_opamp_dummy_magic_23_0.VD2.t2 two_stage_opamp_dummy_magic_23_0.Vb1.t29 two_stage_opamp_dummy_magic_23_0.Y.t18 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X906 GNDA.t366 GNDA.t368 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X907 VOUT-.t138 two_stage_opamp_dummy_magic_23_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X908 VDDA.t683 GNDA.t342 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X909 two_stage_opamp_dummy_magic_23_0.Vb1.t10 VDDA.t210 VDDA.t212 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X910 GNDA.t174 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t29 two_stage_opamp_dummy_magic_23_0.V_source.t23 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X911 VDDA.t684 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X912 VDDA.t685 GNDA.t556 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X913 VOUT-.t139 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X914 VOUT-.t140 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X915 VOUT-.t141 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X916 w_6100_17280.t79 bgr_11_0.V_mir2.t2 bgr_11_0.V_mir2.t3 w_6100_17280.t78 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X917 VDDA.t209 VDDA.t207 GNDA.t126 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X918 w_6100_17280.t5 bgr_11_0.V_mir1.t2 bgr_11_0.V_mir1.t3 w_6100_17280.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X919 VDDA.t686 GNDA.t557 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X920 VDDA.t687 GNDA.t567 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X921 GNDA.t224 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t9 VOUT+.t2 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X922 bgr_11_0.1st_Vout_1.t30 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X923 VDDA.t688 GNDA.t568 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X924 VOUT+.t138 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X925 VDDA.t689 GNDA.t569 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X926 VDDA.t690 GNDA.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X927 VOUT-.t142 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X928 VOUT+.t139 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X929 VDDA.t151 two_stage_opamp_dummy_magic_23_0.Y.t50 VOUT+.t8 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X930 two_stage_opamp_dummy_magic_23_0.Vb2_2.t8 two_stage_opamp_dummy_magic_23_0.Vb2.t9 two_stage_opamp_dummy_magic_23_0.Vb2.t10 two_stage_opamp_dummy_magic_23_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X931 VDDA.t149 two_stage_opamp_dummy_magic_23_0.Y.t51 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t5 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X932 two_stage_opamp_dummy_magic_23_0.V_source.t8 VIN-.t6 two_stage_opamp_dummy_magic_23_0.VD1.t14 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X933 VOUT+.t140 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X934 VDDA.t691 GNDA.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X935 VDDA.t692 GNDA.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X936 two_stage_opamp_dummy_magic_23_0.Vb3.t2 bgr_11_0.NFET_GATE_10uA.t20 GNDA.t217 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X937 GNDA.t211 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_23_0.err_amp_out.t3 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X938 VOUT-.t143 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X939 VDDA.t99 GNDA.t379 GNDA.t381 GNDA.t380 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X940 VOUT-.t144 two_stage_opamp_dummy_magic_23_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X941 VDDA.t63 two_stage_opamp_dummy_magic_23_0.V_err_gate.t32 a_7460_6300.t1 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X942 two_stage_opamp_dummy_magic_23_0.V_source.t15 VIN+.t9 two_stage_opamp_dummy_magic_23_0.VD2.t16 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X943 VOUT-.t145 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X944 VOUT+.t141 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X945 VDDA.t693 GNDA.t201 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X946 two_stage_opamp_dummy_magic_23_0.V_err_gate.t1 two_stage_opamp_dummy_magic_23_0.V_tot.t11 a_7460_6300.t11 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X947 VDDA.t694 GNDA.t202 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X948 GNDA.t299 two_stage_opamp_dummy_magic_23_0.Y.t52 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t1 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X949 two_stage_opamp_dummy_magic_23_0.V_source.t4 VIN-.t7 two_stage_opamp_dummy_magic_23_0.VD1.t11 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X950 VDDA.t188 VDDA.t189 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X951 GNDA.t366 GNDA.t378 bgr_11_0.Vin-.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X952 VDDA.t695 GNDA.t203 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X953 VOUT+.t142 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X954 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X955 VOUT+.t143 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X956 VOUT+.t144 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X957 bgr_11_0.Vin-.t4 VDDA.t696 w_7200_15600.t5 w_7200_15600.t4 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X958 bgr_11_0.V_CMFB_S3.t1 VDDA.t204 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X959 VDDA.t697 GNDA.t339 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X960 VDDA.t698 GNDA.t340 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X961 VDDA.t699 GNDA.t252 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X962 VDDA.t203 VDDA.t201 bgr_11_0.V_CMFB_S3.t0 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X963 VDDA.t700 GNDA.t253 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X964 VDDA.t701 GNDA.t254 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X965 w_6100_17280.t67 VDDA.t190 VDDA.t191 w_6100_17280.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X966 VOUT+.t145 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X967 VOUT+.t7 two_stage_opamp_dummy_magic_23_0.Y.t53 VDDA.t147 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X968 VOUT+.t146 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X969 VOUT+.t147 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 VOUT+.t148 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X971 a_11420_25058.t0 a_11300_23450.t0 GNDA.t198 sky130_fd_pr__res_xhigh_po_0p35 l=6
X972 VDDA.t702 GNDA.t564 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X973 VDDA.t703 GNDA.t565 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X974 VOUT-.t11 GNDA.t375 GNDA.t377 GNDA.t376 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X975 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_23_0.Y.t16 GNDA.t285 sky130_fd_pr__res_high_po_1p41 l=1.41
X976 VDDA.t704 GNDA.t566 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X977 two_stage_opamp_dummy_magic_23_0.VD4.t7 two_stage_opamp_dummy_magic_23_0.Vb3.t27 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X978 two_stage_opamp_dummy_magic_23_0.VD1.t2 two_stage_opamp_dummy_magic_23_0.Vb1.t30 two_stage_opamp_dummy_magic_23_0.X.t8 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X979 VOUT-.t15 two_stage_opamp_dummy_magic_23_0.X.t52 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X980 VOUT+.t149 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X981 VOUT-.t146 two_stage_opamp_dummy_magic_23_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X982 two_stage_opamp_dummy_magic_23_0.VD4.t19 two_stage_opamp_dummy_magic_23_0.Vb2.t32 two_stage_opamp_dummy_magic_23_0.Y.t1 two_stage_opamp_dummy_magic_23_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X983 VOUT-.t16 two_stage_opamp_dummy_magic_23_0.X.t53 VDDA.t402 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X984 VOUT-.t147 two_stage_opamp_dummy_magic_23_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X985 VOUT-.t148 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X986 VDDA.t705 GNDA.t580 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X987 VOUT-.t149 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X988 VDDA.t706 GNDA.t581 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X989 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t0 bgr_11_0.NFET_GATE_10uA.t21 GNDA.t195 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X990 VOUT-.t150 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X991 VDDA.t707 GNDA.t582 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X992 two_stage_opamp_dummy_magic_23_0.VD2.t1 two_stage_opamp_dummy_magic_23_0.Vb1.t31 two_stage_opamp_dummy_magic_23_0.Y.t19 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X993 GNDA.t309 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_23_0.V_p_mir.t2 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X994 a_13570_4368.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t2 GNDA.t200 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X995 VOUT+.t150 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X996 GNDA.t197 bgr_11_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_23_0.Vb2.t1 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X997 w_6100_17280.t83 bgr_11_0.V_mir2.t18 VDDA.t422 w_6100_17280.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X998 two_stage_opamp_dummy_magic_23_0.VD1.t1 two_stage_opamp_dummy_magic_23_0.Vb1.t32 two_stage_opamp_dummy_magic_23_0.X.t7 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X999 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t14 GNDA.t372 GNDA.t374 GNDA.t373 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X1000 GNDA.t338 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t31 two_stage_opamp_dummy_magic_23_0.V_source.t22 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1001 VDDA.t708 GNDA.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1002 VOUT-.t151 two_stage_opamp_dummy_magic_23_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1003 VDDA.t709 GNDA.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1004 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t1 two_stage_opamp_dummy_magic_23_0.X.t54 GNDA.t486 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1005 VDDA.t710 GNDA.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1006 VOUT+.t151 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1007 VDDA.t711 GNDA.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1008 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t4 VDDA.t198 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1009 VDDA.t712 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1010 VDDA.t713 GNDA.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1011 VDDA.t25 a_6520_18930# GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X1012 two_stage_opamp_dummy_magic_23_0.V_source.t14 two_stage_opamp_dummy_magic_23_0.err_amp_out.t12 GNDA.t284 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1013 two_stage_opamp_dummy_magic_23_0.VD4.t6 two_stage_opamp_dummy_magic_23_0.Vb3.t28 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1014 VDDA.t145 two_stage_opamp_dummy_magic_23_0.Y.t54 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t4 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1015 two_stage_opamp_dummy_magic_23_0.V_source.t40 VIN-.t8 two_stage_opamp_dummy_magic_23_0.VD1.t21 GNDA.t244 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1016 VOUT-.t152 two_stage_opamp_dummy_magic_23_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1017 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t12 two_stage_opamp_dummy_magic_23_0.V_err_p.t1 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1018 VOUT-.t153 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1019 VDDA.t714 GNDA.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1020 two_stage_opamp_dummy_magic_23_0.VD4.t2 two_stage_opamp_dummy_magic_23_0.VD4.t0 two_stage_opamp_dummy_magic_23_0.Y.t20 two_stage_opamp_dummy_magic_23_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X1021 VDDA.t715 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1022 VOUT-.t154 two_stage_opamp_dummy_magic_23_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1023 VDDA.t716 GNDA.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1024 GNDA.t371 GNDA.t369 bgr_11_0.NFET_GATE_10uA.t2 GNDA.t370 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X1025 GNDA.t364 GNDA.t362 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t4 GNDA.t363 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1026 w_7200_15600.t1 VDDA.t717 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t2 w_7200_15600.t0 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1027 VDDA.t197 VDDA.t195 bgr_11_0.V_CMFB_S1.t1 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1028 VOUT+.t152 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1029 VOUT+.t153 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1030 VOUT+.t154 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1031 bgr_11_0.V_CMFB_S1.t0 VDDA.t192 VDDA.t194 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X1032 VDDA.t22 two_stage_opamp_dummy_magic_23_0.V_err_gate.t33 two_stage_opamp_dummy_magic_23_0.V_err_p.t5 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1033 VOUT+.t155 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1034 two_stage_opamp_dummy_magic_23_0.V_err_gate.t11 VDDA.t185 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X1035 two_stage_opamp_dummy_magic_23_0.V_source.t12 VIN+.t10 two_stage_opamp_dummy_magic_23_0.VD2.t15 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1036 VDDA.t718 GNDA.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1037 VDDA.t719 GNDA.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1038 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t1 VIN-.t9 two_stage_opamp_dummy_magic_23_0.V_p_mir.t1 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1039 two_stage_opamp_dummy_magic_23_0.V_source.t1 VIN-.t10 two_stage_opamp_dummy_magic_23_0.VD1.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1040 bgr_11_0.1st_Vout_1.t32 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1041 VDDA.t720 GNDA.t332 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 VDDA.t721 GNDA.t333 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1043 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t6 two_stage_opamp_dummy_magic_23_0.V_tot.t13 two_stage_opamp_dummy_magic_23_0.V_err_p.t20 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1044 VOUT-.t155 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1045 VDDA.t722 GNDA.t334 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1046 VOUT+.t156 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1047 VDDA.t723 bgr_11_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1048 w_6100_17280.t35 bgr_11_0.V_mir2.t0 bgr_11_0.V_mir2.t1 w_6100_17280.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1049 VOUT-.t156 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 GNDA.n2000 GNDA.n1820 331711
R1 GNDA.n2125 GNDA.n2124 162800
R2 GNDA.n1999 GNDA.n530 162800
R3 GNDA.n2126 GNDA.n2125 150171
R4 GNDA.n2002 GNDA.n530 150171
R5 GNDA.n1820 GNDA.n1819 112519
R6 GNDA.n2124 GNDA.n2123 111525
R7 GNDA.n1999 GNDA.n1998 111525
R8 GNDA.n1820 GNDA.n1814 86240
R9 GNDA.n2129 GNDA.n506 68514.3
R10 GNDA.n2000 GNDA.t249 63894.4
R11 GNDA.n2129 GNDA.n2128 41014.3
R12 GNDA.n1816 GNDA.n1815 18211.5
R13 GNDA.n2005 GNDA.n530 14938
R14 GNDA.n2125 GNDA.n510 14922.8
R15 GNDA.n2004 GNDA.n518 13700
R16 GNDA.n518 GNDA.n517 13700
R17 GNDA.n532 GNDA.n508 13528.5
R18 GNDA.n1819 GNDA.n507 13213.9
R19 GNDA.n507 GNDA.n506 13034.3
R20 GNDA.n2128 GNDA.n2127 12177.8
R21 GNDA.n2127 GNDA.n2126 11518.4
R22 GNDA.n533 GNDA.n531 11440
R23 GNDA.n2002 GNDA.n2001 11267.1
R24 GNDA.n1817 GNDA.n1816 9910.09
R25 GNDA.n2001 GNDA.n2000 9881.97
R26 GNDA.n1818 GNDA.n1817 9724.16
R27 GNDA.n2001 GNDA.n534 9222.08
R28 GNDA.n1815 GNDA.n1814 8404
R29 GNDA.n2003 GNDA.n531 7648.94
R30 GNDA.n531 GNDA.n509 7630.38
R31 GNDA.n533 GNDA.n508 7385.71
R32 GNDA.n2127 GNDA.n508 6364.29
R33 GNDA.n534 GNDA.n532 5234.66
R34 GNDA.t229 GNDA.t47 5225.11
R35 GNDA.n1818 GNDA.n1814 4106.67
R36 GNDA.n1817 GNDA.n507 4031.21
R37 GNDA.n1815 GNDA.n324 3974.19
R38 GNDA.n2129 GNDA.t288 3568.35
R39 GNDA.n517 GNDA.n509 3498
R40 GNDA.n2004 GNDA.n2003 3463.37
R41 GNDA.n2128 GNDA.n507 2977.78
R42 GNDA.n532 GNDA.n507 2954.29
R43 GNDA.n534 GNDA.n533 2928.92
R44 GNDA.n517 GNDA.n510 2520.94
R45 GNDA.n2005 GNDA.n2004 2481.49
R46 GNDA.t97 GNDA.n2129 2451.21
R47 GNDA.n2000 GNDA.n507 2416.39
R48 GNDA.n2035 GNDA.n518 1800
R49 GNDA.t408 GNDA.n2005 1441.38
R50 GNDA.t418 GNDA.n510 1426.21
R51 GNDA.n2364 GNDA.n2363 1214.72
R52 GNDA.n2363 GNDA.n2362 1214.72
R53 GNDA.n2362 GNDA.n117 1214.72
R54 GNDA.n2356 GNDA.n117 1214.72
R55 GNDA.n2356 GNDA.n55 1214.72
R56 GNDA.n129 GNDA.n56 1214.72
R57 GNDA.n2349 GNDA.n129 1214.72
R58 GNDA.n2349 GNDA.n2348 1214.72
R59 GNDA.n2348 GNDA.n2347 1214.72
R60 GNDA.n2347 GNDA.n57 1214.72
R61 GNDA.n2052 GNDA.n2051 1182.8
R62 GNDA.n2037 GNDA.n2036 1182.8
R63 GNDA.n178 GNDA.n177 970.366
R64 GNDA.n1816 GNDA.n506 927.471
R65 GNDA.t366 GNDA.n55 823.313
R66 GNDA.n1819 GNDA.n1818 776.471
R67 GNDA.n1994 GNDA.t379 749.742
R68 GNDA.n1996 GNDA.t458 749.742
R69 GNDA.n2119 GNDA.t425 749.742
R70 GNDA.n2121 GNDA.t439 749.742
R71 GNDA.n504 GNDA.n503 686.79
R72 GNDA.n505 GNDA.n504 686.79
R73 GNDA.n2186 GNDA.n2185 686.717
R74 GNDA.n590 GNDA.n398 686.717
R75 GNDA.n584 GNDA.n577 686.717
R76 GNDA.n2182 GNDA.n392 686.717
R77 GNDA.n503 GNDA.n502 683.336
R78 GNDA.n709 GNDA.n708 669.307
R79 GNDA.n2160 GNDA.n2159 669.307
R80 GNDA.n1910 GNDA.n103 669.307
R81 GNDA.n2084 GNDA.t454 659.367
R82 GNDA.n2059 GNDA.t433 659.367
R83 GNDA.n1813 GNDA.n1812 585.001
R84 GNDA.n1784 GNDA.n1783 585.001
R85 GNDA.n1799 GNDA.n1798 585.001
R86 GNDA.n611 GNDA.n610 585.001
R87 GNDA.n2155 GNDA.n2154 585.001
R88 GNDA.n712 GNDA.n711 585.001
R89 GNDA.n699 GNDA.n698 585.001
R90 GNDA.n2143 GNDA.n2142 585.001
R91 GNDA.n501 GNDA.n500 585
R92 GNDA.n498 GNDA.n497 585
R93 GNDA.n498 GNDA.n487 585
R94 GNDA.n496 GNDA.n488 585
R95 GNDA.n492 GNDA.n488 585
R96 GNDA.n495 GNDA.n494 585
R97 GNDA.n494 GNDA.n493 585
R98 GNDA.n490 GNDA.n489 585
R99 GNDA.n491 GNDA.n490 585
R100 GNDA.n363 GNDA.n362 585
R101 GNDA.n364 GNDA.n363 585
R102 GNDA.n2214 GNDA.n2213 585
R103 GNDA.n2213 GNDA.n2212 585
R104 GNDA.n2215 GNDA.n361 585
R105 GNDA.n361 GNDA.n360 585
R106 GNDA.n2217 GNDA.n2216 585
R107 GNDA.n2218 GNDA.n2217 585
R108 GNDA.n358 GNDA.n357 585
R109 GNDA.n2219 GNDA.n358 585
R110 GNDA.n2222 GNDA.n2221 585
R111 GNDA.n2221 GNDA.n2220 585
R112 GNDA.n2223 GNDA.n356 585
R113 GNDA.n359 GNDA.n356 585
R114 GNDA.n502 GNDA.n486 585
R115 GNDA.n1047 GNDA.n1046 585
R116 GNDA.n1041 GNDA.n987 585
R117 GNDA.n1045 GNDA.n987 585
R118 GNDA.n1043 GNDA.n1042 585
R119 GNDA.n1044 GNDA.n1043 585
R120 GNDA.n1040 GNDA.n989 585
R121 GNDA.n989 GNDA.n988 585
R122 GNDA.n1039 GNDA.n1038 585
R123 GNDA.n1038 GNDA.n1037 585
R124 GNDA.n1036 GNDA.n990 585
R125 GNDA.n1036 GNDA.n61 585
R126 GNDA.n1035 GNDA.n1034 585
R127 GNDA.n1035 GNDA.n60 585
R128 GNDA.n1033 GNDA.n991 585
R129 GNDA.n1029 GNDA.n991 585
R130 GNDA.n1032 GNDA.n1031 585
R131 GNDA.n1031 GNDA.n1030 585
R132 GNDA.n993 GNDA.n992 585
R133 GNDA.n1028 GNDA.n993 585
R134 GNDA.n1026 GNDA.n1025 585
R135 GNDA.n1027 GNDA.n1026 585
R136 GNDA.n1024 GNDA.n995 585
R137 GNDA.n995 GNDA.n994 585
R138 GNDA.n1049 GNDA.n986 585
R139 GNDA.n917 GNDA.n916 585
R140 GNDA.n915 GNDA.n869 585
R141 GNDA.n914 GNDA.n913 585
R142 GNDA.n912 GNDA.n911 585
R143 GNDA.n910 GNDA.n909 585
R144 GNDA.n908 GNDA.n907 585
R145 GNDA.n906 GNDA.n905 585
R146 GNDA.n904 GNDA.n903 585
R147 GNDA.n902 GNDA.n901 585
R148 GNDA.n900 GNDA.n899 585
R149 GNDA.n853 GNDA.n852 585
R150 GNDA.n1776 GNDA.n853 585
R151 GNDA.n1779 GNDA.n1778 585
R152 GNDA.n1779 GNDA.n851 585
R153 GNDA.n1404 GNDA.n1403 585
R154 GNDA.n1402 GNDA.n1401 585
R155 GNDA.n1400 GNDA.n1399 585
R156 GNDA.n1398 GNDA.n1397 585
R157 GNDA.n1396 GNDA.n1395 585
R158 GNDA.n1394 GNDA.n1393 585
R159 GNDA.n1392 GNDA.n1391 585
R160 GNDA.n1390 GNDA.n1389 585
R161 GNDA.n1388 GNDA.n1387 585
R162 GNDA.n1386 GNDA.n1385 585
R163 GNDA.n1384 GNDA.n864 585
R164 GNDA.n1776 GNDA.n864 585
R165 GNDA.n1383 GNDA.n951 585
R166 GNDA.n1383 GNDA.n1382 585
R167 GNDA.n79 GNDA.n77 585
R168 GNDA.n1774 GNDA.n1773 585
R169 GNDA.n1772 GNDA.n920 585
R170 GNDA.n1776 GNDA.n920 585
R171 GNDA.n1771 GNDA.n1770 585
R172 GNDA.n1769 GNDA.n1768 585
R173 GNDA.n1767 GNDA.n1766 585
R174 GNDA.n1765 GNDA.n1764 585
R175 GNDA.n1763 GNDA.n1762 585
R176 GNDA.n1761 GNDA.n1760 585
R177 GNDA.n1759 GNDA.n1758 585
R178 GNDA.n1757 GNDA.n1756 585
R179 GNDA.n1755 GNDA.n1754 585
R180 GNDA.n1754 GNDA.n1753 585
R181 GNDA.n407 GNDA.n406 585
R182 GNDA.n2157 GNDA.n2156 585
R183 GNDA.n2158 GNDA.n2157 585
R184 GNDA.n707 GNDA.n702 585
R185 GNDA.n704 GNDA.n701 585
R186 GNDA.n710 GNDA.n701 585
R187 GNDA.n589 GNDA.n588 585
R188 GNDA.n579 GNDA.n578 585
R189 GNDA.n591 GNDA.n578 585
R190 GNDA.n583 GNDA.n582 585
R191 GNDA.n2175 GNDA.n394 585
R192 GNDA.n2179 GNDA.n393 585
R193 GNDA.n2187 GNDA.n393 585
R194 GNDA.n2178 GNDA.n2177 585
R195 GNDA.n1781 GNDA.n1780 585
R196 GNDA.n1782 GNDA.n1781 585
R197 GNDA.n1787 GNDA.n1786 585
R198 GNDA.n1786 GNDA.n1785 585
R199 GNDA.n1788 GNDA.n539 585
R200 GNDA.n539 GNDA.n538 585
R201 GNDA.n1796 GNDA.n1795 585
R202 GNDA.n1797 GNDA.n1796 585
R203 GNDA.n543 GNDA.n541 585
R204 GNDA.n541 GNDA.n540 585
R205 GNDA.n573 GNDA.n571 585
R206 GNDA.n571 GNDA.n73 585
R207 GNDA.n576 GNDA.n575 585
R208 GNDA.n592 GNDA.n576 585
R209 GNDA.n596 GNDA.n595 585
R210 GNDA.n595 GNDA.n594 585
R211 GNDA.n567 GNDA.n566 585
R212 GNDA.n593 GNDA.n566 585
R213 GNDA.n606 GNDA.n605 585
R214 GNDA.n607 GNDA.n606 585
R215 GNDA.n564 GNDA.n562 585
R216 GNDA.n608 GNDA.n564 585
R217 GNDA.n796 GNDA.n795 585
R218 GNDA.n795 GNDA.n794 585
R219 GNDA.n789 GNDA.n788 585
R220 GNDA.n789 GNDA.n408 585
R221 GNDA.n786 GNDA.n649 585
R222 GNDA.n649 GNDA.n409 585
R223 GNDA.n655 GNDA.n651 585
R224 GNDA.n657 GNDA.n655 585
R225 GNDA.n781 GNDA.n780 585
R226 GNDA.n780 GNDA.n779 585
R227 GNDA.n659 GNDA.n656 585
R228 GNDA.n778 GNDA.n656 585
R229 GNDA.n776 GNDA.n775 585
R230 GNDA.n777 GNDA.n776 585
R231 GNDA.n686 GNDA.n658 585
R232 GNDA.n683 GNDA.n658 585
R233 GNDA.n688 GNDA.n685 585
R234 GNDA.n685 GNDA.n684 585
R235 GNDA.n694 GNDA.n693 585
R236 GNDA.n695 GNDA.n694 585
R237 GNDA.n680 GNDA.n679 585
R238 GNDA.n696 GNDA.n680 585
R239 GNDA.n715 GNDA.n714 585
R240 GNDA.n714 GNDA.n713 585
R241 GNDA.n682 GNDA.n681 585
R242 GNDA.n700 GNDA.n682 585
R243 GNDA.n432 GNDA.n431 585
R244 GNDA.n431 GNDA.n430 585
R245 GNDA.n390 GNDA.n388 585
R246 GNDA.n429 GNDA.n390 585
R247 GNDA.n2202 GNDA.n2201 585
R248 GNDA.n2201 GNDA.n2200 585
R249 GNDA.n2189 GNDA.n391 585
R250 GNDA.n2199 GNDA.n391 585
R251 GNDA.n2197 GNDA.n2196 585
R252 GNDA.n2198 GNDA.n2197 585
R253 GNDA.n2192 GNDA.n365 585
R254 GNDA.n2188 GNDA.n365 585
R255 GNDA.n2210 GNDA.n2209 585
R256 GNDA.n2211 GNDA.n2210 585
R257 GNDA.n367 GNDA.n366 585
R258 GNDA.n418 GNDA.n366 585
R259 GNDA.n424 GNDA.n421 585
R260 GNDA.n421 GNDA.n419 585
R261 GNDA.n2140 GNDA.n2139 585
R262 GNDA.n2141 GNDA.n2140 585
R263 GNDA.n427 GNDA.n422 585
R264 GNDA.n422 GNDA.n420 585
R265 GNDA.n2133 GNDA.n2132 585
R266 GNDA.n2132 GNDA.n2131 585
R267 GNDA.n2225 GNDA.n2224 585
R268 GNDA.n2227 GNDA.n354 585
R269 GNDA.n2229 GNDA.n2228 585
R270 GNDA.n2230 GNDA.n353 585
R271 GNDA.n2232 GNDA.n2231 585
R272 GNDA.n2234 GNDA.n351 585
R273 GNDA.n2236 GNDA.n2235 585
R274 GNDA.n2237 GNDA.n350 585
R275 GNDA.n2239 GNDA.n2238 585
R276 GNDA.n2241 GNDA.n348 585
R277 GNDA.n2243 GNDA.n2242 585
R278 GNDA.n2244 GNDA.n347 585
R279 GNDA.n1381 GNDA.n952 585
R280 GNDA.n1368 GNDA.n953 585
R281 GNDA.n1377 GNDA.n1376 585
R282 GNDA.n1267 GNDA.n1265 585
R283 GNDA.n1293 GNDA.n1292 585
R284 GNDA.n1297 GNDA.n1296 585
R285 GNDA.n1299 GNDA.n1298 585
R286 GNDA.n1306 GNDA.n1305 585
R287 GNDA.n1304 GNDA.n1290 585
R288 GNDA.n1312 GNDA.n1311 585
R289 GNDA.n1314 GNDA.n1313 585
R290 GNDA.n1288 GNDA.n1287 585
R291 GNDA.n1146 GNDA.n311 585
R292 GNDA.n1259 GNDA.n1258 585
R293 GNDA.n1148 GNDA.n1145 585
R294 GNDA.n1253 GNDA.n1252 585
R295 GNDA.n1251 GNDA.n1250 585
R296 GNDA.n1176 GNDA.n1152 585
R297 GNDA.n1178 GNDA.n1177 585
R298 GNDA.n1183 GNDA.n1182 585
R299 GNDA.n1181 GNDA.n1174 585
R300 GNDA.n1189 GNDA.n1188 585
R301 GNDA.n1191 GNDA.n1190 585
R302 GNDA.n1172 GNDA.n1171 585
R303 GNDA.n960 GNDA.n306 585
R304 GNDA.n1138 GNDA.n1137 585
R305 GNDA.n962 GNDA.n959 585
R306 GNDA.n1132 GNDA.n1131 585
R307 GNDA.n1130 GNDA.n1129 585
R308 GNDA.n1055 GNDA.n966 585
R309 GNDA.n1057 GNDA.n1056 585
R310 GNDA.n1062 GNDA.n1061 585
R311 GNDA.n1060 GNDA.n1053 585
R312 GNDA.n1068 GNDA.n1067 585
R313 GNDA.n1070 GNDA.n1069 585
R314 GNDA.n1051 GNDA.n1050 585
R315 GNDA.n1428 GNDA.n945 585
R316 GNDA.n1426 GNDA.n1425 585
R317 GNDA.n1424 GNDA.n946 585
R318 GNDA.n1423 GNDA.n1422 585
R319 GNDA.n1420 GNDA.n947 585
R320 GNDA.n1418 GNDA.n1417 585
R321 GNDA.n1416 GNDA.n948 585
R322 GNDA.n1415 GNDA.n1414 585
R323 GNDA.n1412 GNDA.n949 585
R324 GNDA.n1410 GNDA.n1409 585
R325 GNDA.n1408 GNDA.n950 585
R326 GNDA.n1407 GNDA.n1406 585
R327 GNDA.n1437 GNDA.n278 585
R328 GNDA.n1440 GNDA.n1439 585
R329 GNDA.n1442 GNDA.n1441 585
R330 GNDA.n1444 GNDA.n1435 585
R331 GNDA.n1446 GNDA.n1445 585
R332 GNDA.n1447 GNDA.n1434 585
R333 GNDA.n1449 GNDA.n1448 585
R334 GNDA.n1451 GNDA.n1432 585
R335 GNDA.n1453 GNDA.n1452 585
R336 GNDA.n1454 GNDA.n1431 585
R337 GNDA.n1456 GNDA.n1455 585
R338 GNDA.n1458 GNDA.n944 585
R339 GNDA.n1023 GNDA.n1022 585
R340 GNDA.n1020 GNDA.n996 585
R341 GNDA.n1019 GNDA.n1018 585
R342 GNDA.n1017 GNDA.n1016 585
R343 GNDA.n1015 GNDA.n998 585
R344 GNDA.n1013 GNDA.n1012 585
R345 GNDA.n1011 GNDA.n999 585
R346 GNDA.n1010 GNDA.n1009 585
R347 GNDA.n1007 GNDA.n1000 585
R348 GNDA.n1005 GNDA.n1004 585
R349 GNDA.n1003 GNDA.n1002 585
R350 GNDA.n282 GNDA.n279 585
R351 GNDA.n1752 GNDA.n1751 585
R352 GNDA.n1749 GNDA.n1748 585
R353 GNDA.n1747 GNDA.n1746 585
R354 GNDA.n1663 GNDA.n923 585
R355 GNDA.n1665 GNDA.n1664 585
R356 GNDA.n1669 GNDA.n1668 585
R357 GNDA.n1671 GNDA.n1670 585
R358 GNDA.n1678 GNDA.n1677 585
R359 GNDA.n1676 GNDA.n1661 585
R360 GNDA.n1684 GNDA.n1683 585
R361 GNDA.n1686 GNDA.n1685 585
R362 GNDA.n1659 GNDA.n1658 585
R363 GNDA.n2401 GNDA.n88 585
R364 GNDA.n2401 GNDA.n64 585
R365 GNDA.n2404 GNDA.n2403 585
R366 GNDA.n2403 GNDA.n2402 585
R367 GNDA.n2405 GNDA.n87 585
R368 GNDA.n87 GNDA.n86 585
R369 GNDA.n2407 GNDA.n2406 585
R370 GNDA.n2408 GNDA.n2407 585
R371 GNDA.n85 GNDA.n84 585
R372 GNDA.n2409 GNDA.n85 585
R373 GNDA.n2412 GNDA.n2411 585
R374 GNDA.n2411 GNDA.n2410 585
R375 GNDA.n2413 GNDA.n83 585
R376 GNDA.n83 GNDA.n82 585
R377 GNDA.n2415 GNDA.n2414 585
R378 GNDA.n2416 GNDA.n2415 585
R379 GNDA.n81 GNDA.n80 585
R380 GNDA.n2417 GNDA.n81 585
R381 GNDA.n2420 GNDA.n2419 585
R382 GNDA.n2419 GNDA.n2418 585
R383 GNDA.n2421 GNDA.n78 585
R384 GNDA.n78 GNDA.n76 585
R385 GNDA.n2423 GNDA.n2422 585
R386 GNDA.n2424 GNDA.n2423 585
R387 GNDA.n145 GNDA.n144 585
R388 GNDA.n177 GNDA.n145 585
R389 GNDA.n175 GNDA.n174 585
R390 GNDA.n176 GNDA.n175 585
R391 GNDA.n173 GNDA.n147 585
R392 GNDA.n147 GNDA.n146 585
R393 GNDA.n172 GNDA.n171 585
R394 GNDA.n171 GNDA.n170 585
R395 GNDA.n149 GNDA.n148 585
R396 GNDA.n169 GNDA.n149 585
R397 GNDA.n167 GNDA.n166 585
R398 GNDA.n168 GNDA.n167 585
R399 GNDA.n165 GNDA.n150 585
R400 GNDA.n161 GNDA.n150 585
R401 GNDA.n164 GNDA.n163 585
R402 GNDA.n163 GNDA.n162 585
R403 GNDA.n152 GNDA.n151 585
R404 GNDA.n160 GNDA.n152 585
R405 GNDA.n158 GNDA.n157 585
R406 GNDA.n159 GNDA.n158 585
R407 GNDA.n156 GNDA.n155 585
R408 GNDA.n155 GNDA.n154 585
R409 GNDA.n113 GNDA.n111 585
R410 GNDA.n153 GNDA.n113 585
R411 GNDA.n200 GNDA.n199 585
R412 GNDA.n200 GNDA.n136 585
R413 GNDA.n198 GNDA.n137 585
R414 GNDA.n194 GNDA.n137 585
R415 GNDA.n197 GNDA.n196 585
R416 GNDA.n196 GNDA.n195 585
R417 GNDA.n192 GNDA.n138 585
R418 GNDA.n193 GNDA.n192 585
R419 GNDA.n191 GNDA.n190 585
R420 GNDA.n191 GNDA.n59 585
R421 GNDA.n189 GNDA.n139 585
R422 GNDA.n139 GNDA.n58 585
R423 GNDA.n188 GNDA.n187 585
R424 GNDA.n187 GNDA.n186 585
R425 GNDA.n141 GNDA.n140 585
R426 GNDA.n185 GNDA.n141 585
R427 GNDA.n183 GNDA.n182 585
R428 GNDA.n184 GNDA.n183 585
R429 GNDA.n181 GNDA.n143 585
R430 GNDA.n143 GNDA.n142 585
R431 GNDA.n180 GNDA.n179 585
R432 GNDA.n179 GNDA.n178 585
R433 GNDA.n202 GNDA.n201 585
R434 GNDA.n204 GNDA.n203 585
R435 GNDA.n2340 GNDA.n274 585
R436 GNDA.n24 GNDA.n22 585
R437 GNDA.n2429 GNDA.n2428 585
R438 GNDA.n37 GNDA.n25 585
R439 GNDA.n45 GNDA.n44 585
R440 GNDA.n40 GNDA.n36 585
R441 GNDA.n35 GNDA.n0 585
R442 GNDA.n209 GNDA.n1 585
R443 GNDA.n211 GNDA.n210 585
R444 GNDA.n215 GNDA.n214 585
R445 GNDA.n217 GNDA.n216 585
R446 GNDA.n206 GNDA.n205 585
R447 GNDA.n1654 GNDA.n1653 585
R448 GNDA.n1651 GNDA.n1650 585
R449 GNDA.n1649 GNDA.n1648 585
R450 GNDA.n1565 GNDA.n1543 585
R451 GNDA.n1567 GNDA.n1566 585
R452 GNDA.n1571 GNDA.n1570 585
R453 GNDA.n1573 GNDA.n1572 585
R454 GNDA.n1580 GNDA.n1579 585
R455 GNDA.n1578 GNDA.n1563 585
R456 GNDA.n1586 GNDA.n1585 585
R457 GNDA.n1588 GNDA.n1587 585
R458 GNDA.n276 GNDA.n275 585
R459 GNDA.n2344 GNDA.n133 585
R460 GNDA.n133 GNDA.n57 585
R461 GNDA.n2345 GNDA.n131 585
R462 GNDA.n2347 GNDA.n131 585
R463 GNDA.n130 GNDA.n127 585
R464 GNDA.n2348 GNDA.n130 585
R465 GNDA.n2351 GNDA.n126 585
R466 GNDA.n2349 GNDA.n126 585
R467 GNDA.n2352 GNDA.n125 585
R468 GNDA.n129 GNDA.n125 585
R469 GNDA.n2353 GNDA.n124 585
R470 GNDA.n124 GNDA.n56 585
R471 GNDA.n123 GNDA.n121 585
R472 GNDA.n123 GNDA.n55 585
R473 GNDA.n2358 GNDA.n120 585
R474 GNDA.n2356 GNDA.n120 585
R475 GNDA.n2359 GNDA.n119 585
R476 GNDA.n119 GNDA.n117 585
R477 GNDA.n2360 GNDA.n116 585
R478 GNDA.n2362 GNDA.n116 585
R479 GNDA.n115 GNDA.n112 585
R480 GNDA.n2363 GNDA.n115 585
R481 GNDA.n2366 GNDA.n110 585
R482 GNDA.n2364 GNDA.n110 585
R483 GNDA.n2342 GNDA.n277 585
R484 GNDA.n277 GNDA.n54 585
R485 GNDA.n2366 GNDA.n2365 585
R486 GNDA.n2365 GNDA.n2364 585
R487 GNDA.n114 GNDA.n112 585
R488 GNDA.n2363 GNDA.n114 585
R489 GNDA.n2361 GNDA.n2360 585
R490 GNDA.n2362 GNDA.n2361 585
R491 GNDA.n2359 GNDA.n118 585
R492 GNDA.n118 GNDA.n117 585
R493 GNDA.n2358 GNDA.n2357 585
R494 GNDA.n2357 GNDA.n2356 585
R495 GNDA.n2355 GNDA.n121 585
R496 GNDA.n2355 GNDA.n55 585
R497 GNDA.n2354 GNDA.n2353 585
R498 GNDA.n2354 GNDA.n56 585
R499 GNDA.n2352 GNDA.n122 585
R500 GNDA.n129 GNDA.n122 585
R501 GNDA.n2351 GNDA.n2350 585
R502 GNDA.n2350 GNDA.n2349 585
R503 GNDA.n128 GNDA.n127 585
R504 GNDA.n2348 GNDA.n128 585
R505 GNDA.n2346 GNDA.n2345 585
R506 GNDA.n2347 GNDA.n2346 585
R507 GNDA.n2344 GNDA.n132 585
R508 GNDA.n132 GNDA.n57 585
R509 GNDA.n2342 GNDA.n2341 585
R510 GNDA.n2341 GNDA.n54 585
R511 GNDA.n2317 GNDA.n304 585
R512 GNDA.n2318 GNDA.n302 585
R513 GNDA.n2319 GNDA.n301 585
R514 GNDA.n299 GNDA.n297 585
R515 GNDA.n2325 GNDA.n296 585
R516 GNDA.n2326 GNDA.n294 585
R517 GNDA.n2327 GNDA.n293 585
R518 GNDA.n291 GNDA.n289 585
R519 GNDA.n2332 GNDA.n288 585
R520 GNDA.n2333 GNDA.n286 585
R521 GNDA.n285 GNDA.n281 585
R522 GNDA.n2338 GNDA.n280 585
R523 GNDA.n309 GNDA.n307 585
R524 GNDA.n2313 GNDA.n309 585
R525 GNDA.n2338 GNDA.n2337 585
R526 GNDA.n2335 GNDA.n281 585
R527 GNDA.n2334 GNDA.n2333 585
R528 GNDA.n2332 GNDA.n2331 585
R529 GNDA.n2330 GNDA.n289 585
R530 GNDA.n2328 GNDA.n2327 585
R531 GNDA.n2326 GNDA.n290 585
R532 GNDA.n2325 GNDA.n2324 585
R533 GNDA.n2322 GNDA.n297 585
R534 GNDA.n2320 GNDA.n2319 585
R535 GNDA.n2318 GNDA.n298 585
R536 GNDA.n2317 GNDA.n2316 585
R537 GNDA.n2314 GNDA.n307 585
R538 GNDA.n2314 GNDA.n2313 585
R539 GNDA.n2303 GNDA.n2302 585
R540 GNDA.n332 GNDA.n330 585
R541 GNDA.n338 GNDA.n337 585
R542 GNDA.n2295 GNDA.n2294 585
R543 GNDA.n2293 GNDA.n2292 585
R544 GNDA.n2291 GNDA.n342 585
R545 GNDA.n341 GNDA.n340 585
R546 GNDA.n2285 GNDA.n2284 585
R547 GNDA.n2283 GNDA.n2282 585
R548 GNDA.n2281 GNDA.n346 585
R549 GNDA.n345 GNDA.n344 585
R550 GNDA.n2275 GNDA.n2274 585
R551 GNDA.n334 GNDA.n331 585
R552 GNDA.n697 GNDA.n331 585
R553 GNDA.n2276 GNDA.n2275 585
R554 GNDA.n2278 GNDA.n344 585
R555 GNDA.n2281 GNDA.n2280 585
R556 GNDA.n2282 GNDA.n343 585
R557 GNDA.n2286 GNDA.n2285 585
R558 GNDA.n2288 GNDA.n340 585
R559 GNDA.n2291 GNDA.n2290 585
R560 GNDA.n2292 GNDA.n339 585
R561 GNDA.n2296 GNDA.n2295 585
R562 GNDA.n2298 GNDA.n338 585
R563 GNDA.n2299 GNDA.n332 585
R564 GNDA.n2302 GNDA.n2301 585
R565 GNDA.n335 GNDA.n334 585
R566 GNDA.n428 GNDA.n335 585
R567 GNDA.n2273 GNDA.n2272 585
R568 GNDA.n2271 GNDA.n2270 585
R569 GNDA.n2269 GNDA.n2247 585
R570 GNDA.n2267 GNDA.n2266 585
R571 GNDA.n2265 GNDA.n2248 585
R572 GNDA.n2264 GNDA.n2263 585
R573 GNDA.n2261 GNDA.n2249 585
R574 GNDA.n2259 GNDA.n2258 585
R575 GNDA.n2257 GNDA.n2250 585
R576 GNDA.n2256 GNDA.n2255 585
R577 GNDA.n2253 GNDA.n2251 585
R578 GNDA.n317 GNDA.n313 585
R579 GNDA.n879 GNDA.n314 585
R580 GNDA.n881 GNDA.n877 585
R581 GNDA.n883 GNDA.n882 585
R582 GNDA.n884 GNDA.n876 585
R583 GNDA.n886 GNDA.n885 585
R584 GNDA.n888 GNDA.n874 585
R585 GNDA.n890 GNDA.n889 585
R586 GNDA.n891 GNDA.n873 585
R587 GNDA.n893 GNDA.n892 585
R588 GNDA.n895 GNDA.n871 585
R589 GNDA.n897 GNDA.n896 585
R590 GNDA.n898 GNDA.n870 585
R591 GNDA.n647 GNDA.n646 585
R592 GNDA.n644 GNDA.n612 585
R593 GNDA.n643 GNDA.n642 585
R594 GNDA.n639 GNDA.n636 585
R595 GNDA.n635 GNDA.n614 585
R596 GNDA.n633 GNDA.n632 585
R597 GNDA.n629 GNDA.n615 585
R598 GNDA.n628 GNDA.n625 585
R599 GNDA.n623 GNDA.n616 585
R600 GNDA.n621 GNDA.n620 585
R601 GNDA.n618 GNDA.n316 585
R602 GNDA.n2309 GNDA.n315 585
R603 GNDA.n790 GNDA.n565 585
R604 GNDA.n793 GNDA.n565 585
R605 GNDA.n2309 GNDA.n2308 585
R606 GNDA.n318 GNDA.n316 585
R607 GNDA.n620 GNDA.n619 585
R608 GNDA.n626 GNDA.n616 585
R609 GNDA.n628 GNDA.n627 585
R610 GNDA.n630 GNDA.n629 585
R611 GNDA.n632 GNDA.n631 585
R612 GNDA.n637 GNDA.n614 585
R613 GNDA.n639 GNDA.n638 585
R614 GNDA.n642 GNDA.n641 585
R615 GNDA.n640 GNDA.n612 585
R616 GNDA.n648 GNDA.n647 585
R617 GNDA.n791 GNDA.n790 585
R618 GNDA.n792 GNDA.n791 585
R619 GNDA.n1482 GNDA.n1481 585
R620 GNDA.n1483 GNDA.n1479 585
R621 GNDA.n1484 GNDA.n1478 585
R622 GNDA.n1476 GNDA.n1473 585
R623 GNDA.n1490 GNDA.n1472 585
R624 GNDA.n1491 GNDA.n1470 585
R625 GNDA.n1492 GNDA.n1469 585
R626 GNDA.n1467 GNDA.n1465 585
R627 GNDA.n1497 GNDA.n1464 585
R628 GNDA.n1498 GNDA.n1462 585
R629 GNDA.n1461 GNDA.n1430 585
R630 GNDA.n1503 GNDA.n1429 585
R631 GNDA.n2311 GNDA.n308 585
R632 GNDA.n2313 GNDA.n308 585
R633 GNDA.n1503 GNDA.n1502 585
R634 GNDA.n1500 GNDA.n1430 585
R635 GNDA.n1499 GNDA.n1498 585
R636 GNDA.n1497 GNDA.n1496 585
R637 GNDA.n1495 GNDA.n1465 585
R638 GNDA.n1493 GNDA.n1492 585
R639 GNDA.n1491 GNDA.n1466 585
R640 GNDA.n1490 GNDA.n1489 585
R641 GNDA.n1487 GNDA.n1473 585
R642 GNDA.n1485 GNDA.n1484 585
R643 GNDA.n1483 GNDA.n1475 585
R644 GNDA.n1482 GNDA.n310 585
R645 GNDA.n2312 GNDA.n2311 585
R646 GNDA.n2313 GNDA.n2312 585
R647 GNDA.n1505 GNDA.n943 585
R648 GNDA.n1537 GNDA.n1536 585
R649 GNDA.n1534 GNDA.n1507 585
R650 GNDA.n1532 GNDA.n1531 585
R651 GNDA.n1509 GNDA.n1508 585
R652 GNDA.n1525 GNDA.n1524 585
R653 GNDA.n1522 GNDA.n1511 585
R654 GNDA.n1520 GNDA.n1519 585
R655 GNDA.n1514 GNDA.n1513 585
R656 GNDA.n91 GNDA.n90 585
R657 GNDA.n2398 GNDA.n2397 585
R658 GNDA.n2400 GNDA.n89 585
R659 GNDA.n1657 GNDA.n1656 585
R660 GNDA.n1657 GNDA.n54 585
R661 GNDA.n2394 GNDA.n89 585
R662 GNDA.n2397 GNDA.n2396 585
R663 GNDA.n92 GNDA.n91 585
R664 GNDA.n1516 GNDA.n1514 585
R665 GNDA.n1519 GNDA.n1518 585
R666 GNDA.n1511 GNDA.n1510 585
R667 GNDA.n1526 GNDA.n1525 585
R668 GNDA.n1528 GNDA.n1509 585
R669 GNDA.n1531 GNDA.n1530 585
R670 GNDA.n1507 GNDA.n1506 585
R671 GNDA.n1538 GNDA.n1537 585
R672 GNDA.n1540 GNDA.n1505 585
R673 GNDA.n1656 GNDA.n1655 585
R674 GNDA.n1655 GNDA.n54 585
R675 GNDA.n2369 GNDA.n2368 585
R676 GNDA.n2370 GNDA.n2369 585
R677 GNDA.n107 GNDA.n106 585
R678 GNDA.n2371 GNDA.n107 585
R679 GNDA.n2374 GNDA.n2373 585
R680 GNDA.n2373 GNDA.n2372 585
R681 GNDA.n2375 GNDA.n105 585
R682 GNDA.n108 GNDA.n105 585
R683 GNDA.n2377 GNDA.n2376 585
R684 GNDA.n2377 GNDA.n104 585
R685 GNDA.n2378 GNDA.n100 585
R686 GNDA.n2379 GNDA.n2378 585
R687 GNDA.n2383 GNDA.n99 585
R688 GNDA.n99 GNDA.n98 585
R689 GNDA.n2385 GNDA.n2384 585
R690 GNDA.n2386 GNDA.n2385 585
R691 GNDA.n96 GNDA.n95 585
R692 GNDA.n2387 GNDA.n96 585
R693 GNDA.n2390 GNDA.n2389 585
R694 GNDA.n2389 GNDA.n2388 585
R695 GNDA.n2391 GNDA.n93 585
R696 GNDA.n97 GNDA.n93 585
R697 GNDA.n2393 GNDA.n2392 585
R698 GNDA.n2393 GNDA.n63 585
R699 GNDA.n102 GNDA.n101 585
R700 GNDA.n2381 GNDA.n2380 585
R701 GNDA.n2380 GNDA.t366 585
R702 GNDA.n1990 GNDA.t385 524.808
R703 GNDA.n1983 GNDA.t375 524.808
R704 GNDA.n2114 GNDA.t442 524.808
R705 GNDA.n2107 GNDA.t436 524.808
R706 GNDA.t366 GNDA.n57 512.884
R707 GNDA.n523 GNDA.t445 508.743
R708 GNDA.n2092 GNDA.t388 508.743
R709 GNDA.n2031 GNDA.t393 508.743
R710 GNDA.n2028 GNDA.t401 508.743
R711 GNDA.n2010 GNDA.t415 499.442
R712 GNDA.n2019 GNDA.t423 499.442
R713 GNDA.n2006 GNDA.t407 499.442
R714 GNDA.n522 GNDA.t417 499.442
R715 GNDA.n2008 GNDA.n529 497.837
R716 GNDA.n2117 GNDA.n513 490.517
R717 GNDA.n2015 GNDA.t421 475.976
R718 GNDA.n2015 GNDA.t399 475.976
R719 GNDA.n2021 GNDA.t410 475.976
R720 GNDA.n2021 GNDA.t391 475.976
R721 GNDA.n537 GNDA.t428 425.134
R722 GNDA.n1811 GNDA.t369 409.067
R723 GNDA.n2144 GNDA.t448 409.067
R724 GNDA.n414 GNDA.t404 409.067
R725 GNDA.n413 GNDA.t461 409.067
R726 GNDA.n2153 GNDA.t412 409.067
R727 GNDA.n609 GNDA.t372 409.067
R728 GNDA.n1800 GNDA.t451 409.067
R729 GNDA.t366 GNDA.n56 391.411
R730 GNDA.n504 GNDA.t46 371.606
R731 GNDA.n2050 GNDA.t362 338.034
R732 GNDA.n2038 GNDA.t382 338.034
R733 GNDA.t118 GNDA.t324 333.793
R734 GNDA.t52 GNDA.t118 333.793
R735 GNDA.t26 GNDA.t52 333.793
R736 GNDA.t77 GNDA.t210 333.793
R737 GNDA.t315 GNDA.t77 333.793
R738 GNDA.t551 GNDA.t315 333.793
R739 GNDA.t208 GNDA.t245 333.793
R740 GNDA.t207 GNDA.t245 333.793
R741 GNDA.t366 GNDA.n72 172.876
R742 GNDA.t366 GNDA.n2305 172.876
R743 GNDA.n2306 GNDA.t366 172.615
R744 GNDA.t366 GNDA.n336 172.615
R745 GNDA.n525 GNDA.n524 296.158
R746 GNDA.n2091 GNDA.n2090 296.158
R747 GNDA.n2033 GNDA.n2032 296.158
R748 GNDA.n2027 GNDA.n2026 296.158
R749 GNDA.n2009 GNDA.n2008 292.5
R750 GNDA.n2033 GNDA.n519 292.5
R751 GNDA.n2026 GNDA.n2025 292.5
R752 GNDA.n2018 GNDA.n513 292.5
R753 GNDA.n2008 GNDA.n2007 292.5
R754 GNDA.n521 GNDA.n513 292.5
R755 GNDA.t312 GNDA.t429 273.139
R756 GNDA.n499 GNDA.n485 264.301
R757 GNDA.n1048 GNDA.n985 264.301
R758 GNDA.n1777 GNDA.n1776 264.301
R759 GNDA.n1776 GNDA.n919 264.301
R760 GNDA.n1776 GNDA.n858 264.301
R761 GNDA.n135 GNDA.n134 264.301
R762 GNDA.n2274 GNDA.n2273 259.416
R763 GNDA.n2369 GNDA.n110 259.416
R764 GNDA.n1437 GNDA.n280 259.416
R765 GNDA.n1022 GNDA.n995 259.416
R766 GNDA.n2225 GNDA.n356 259.416
R767 GNDA.n2401 GNDA.n2400 259.416
R768 GNDA.n1429 GNDA.n1428 259.416
R769 GNDA.n879 GNDA.n315 259.416
R770 GNDA.n179 GNDA.n145 259.416
R771 GNDA.n1627 GNDA.n1626 258.334
R772 GNDA.n256 GNDA.n255 258.334
R773 GNDA.n1228 GNDA.n1169 258.334
R774 GNDA.n752 GNDA.n676 258.334
R775 GNDA.n1107 GNDA.n983 258.334
R776 GNDA.n451 GNDA.n450 258.334
R777 GNDA.n1725 GNDA.n1724 258.334
R778 GNDA.n1353 GNDA.n1352 258.334
R779 GNDA.n833 GNDA.n831 258.334
R780 GNDA.n2052 GNDA.t111 257.932
R781 GNDA.n2036 GNDA.t59 257.932
R782 GNDA.n1776 GNDA.n918 254.34
R783 GNDA.n1776 GNDA.n868 254.34
R784 GNDA.n1776 GNDA.n867 254.34
R785 GNDA.n1776 GNDA.n866 254.34
R786 GNDA.n1776 GNDA.n865 254.34
R787 GNDA.n1776 GNDA.n859 254.34
R788 GNDA.n1776 GNDA.n860 254.34
R789 GNDA.n1776 GNDA.n861 254.34
R790 GNDA.n1776 GNDA.n862 254.34
R791 GNDA.n1776 GNDA.n863 254.34
R792 GNDA.n1776 GNDA.n1775 254.34
R793 GNDA.n1776 GNDA.n854 254.34
R794 GNDA.n1776 GNDA.n855 254.34
R795 GNDA.n1776 GNDA.n856 254.34
R796 GNDA.n1776 GNDA.n857 254.34
R797 GNDA.n2226 GNDA.n75 254.34
R798 GNDA.n355 GNDA.n75 254.34
R799 GNDA.n2233 GNDA.n75 254.34
R800 GNDA.n352 GNDA.n75 254.34
R801 GNDA.n2240 GNDA.n75 254.34
R802 GNDA.n349 GNDA.n75 254.34
R803 GNDA.n1380 GNDA.n1379 254.34
R804 GNDA.n1379 GNDA.n1378 254.34
R805 GNDA.n1379 GNDA.n1264 254.34
R806 GNDA.n1379 GNDA.n1263 254.34
R807 GNDA.n1379 GNDA.n1262 254.34
R808 GNDA.n1379 GNDA.n1261 254.34
R809 GNDA.n1379 GNDA.n1260 254.34
R810 GNDA.n1379 GNDA.n1144 254.34
R811 GNDA.n1379 GNDA.n1143 254.34
R812 GNDA.n1379 GNDA.n1142 254.34
R813 GNDA.n1379 GNDA.n1141 254.34
R814 GNDA.n1379 GNDA.n1140 254.34
R815 GNDA.n1379 GNDA.n1139 254.34
R816 GNDA.n1379 GNDA.n958 254.34
R817 GNDA.n1379 GNDA.n957 254.34
R818 GNDA.n1379 GNDA.n956 254.34
R819 GNDA.n1379 GNDA.n955 254.34
R820 GNDA.n1379 GNDA.n954 254.34
R821 GNDA.n1427 GNDA.n67 254.34
R822 GNDA.n1421 GNDA.n67 254.34
R823 GNDA.n1419 GNDA.n67 254.34
R824 GNDA.n1413 GNDA.n67 254.34
R825 GNDA.n1411 GNDA.n67 254.34
R826 GNDA.n1405 GNDA.n67 254.34
R827 GNDA.n1438 GNDA.n67 254.34
R828 GNDA.n1443 GNDA.n67 254.34
R829 GNDA.n1436 GNDA.n67 254.34
R830 GNDA.n1450 GNDA.n67 254.34
R831 GNDA.n1433 GNDA.n67 254.34
R832 GNDA.n1457 GNDA.n67 254.34
R833 GNDA.n1021 GNDA.n67 254.34
R834 GNDA.n997 GNDA.n67 254.34
R835 GNDA.n1014 GNDA.n67 254.34
R836 GNDA.n1008 GNDA.n67 254.34
R837 GNDA.n1006 GNDA.n67 254.34
R838 GNDA.n1001 GNDA.n67 254.34
R839 GNDA.n2426 GNDA.n53 254.34
R840 GNDA.n2426 GNDA.n52 254.34
R841 GNDA.n2426 GNDA.n51 254.34
R842 GNDA.n2426 GNDA.n50 254.34
R843 GNDA.n2426 GNDA.n49 254.34
R844 GNDA.n2426 GNDA.n48 254.34
R845 GNDA.n2426 GNDA.n47 254.34
R846 GNDA.n2427 GNDA.n2426 254.34
R847 GNDA.n2426 GNDA.n46 254.34
R848 GNDA.n2426 GNDA.n34 254.34
R849 GNDA.n2426 GNDA.n33 254.34
R850 GNDA.n2426 GNDA.n32 254.34
R851 GNDA.n2426 GNDA.n31 254.34
R852 GNDA.n2426 GNDA.n30 254.34
R853 GNDA.n2426 GNDA.n29 254.34
R854 GNDA.n2426 GNDA.n28 254.34
R855 GNDA.n2426 GNDA.n27 254.34
R856 GNDA.n2426 GNDA.n26 254.34
R857 GNDA.n303 GNDA.n68 254.34
R858 GNDA.n300 GNDA.n68 254.34
R859 GNDA.n295 GNDA.n68 254.34
R860 GNDA.n292 GNDA.n68 254.34
R861 GNDA.n287 GNDA.n68 254.34
R862 GNDA.n284 GNDA.n68 254.34
R863 GNDA.n2336 GNDA.n70 254.34
R864 GNDA.n283 GNDA.n70 254.34
R865 GNDA.n2329 GNDA.n70 254.34
R866 GNDA.n2323 GNDA.n70 254.34
R867 GNDA.n2321 GNDA.n70 254.34
R868 GNDA.n2315 GNDA.n70 254.34
R869 GNDA.n2305 GNDA.n2304 254.34
R870 GNDA.n2305 GNDA.n329 254.34
R871 GNDA.n2305 GNDA.n328 254.34
R872 GNDA.n2305 GNDA.n327 254.34
R873 GNDA.n2305 GNDA.n326 254.34
R874 GNDA.n2305 GNDA.n325 254.34
R875 GNDA.n2277 GNDA.n336 254.34
R876 GNDA.n2279 GNDA.n336 254.34
R877 GNDA.n2287 GNDA.n336 254.34
R878 GNDA.n2289 GNDA.n336 254.34
R879 GNDA.n2297 GNDA.n336 254.34
R880 GNDA.n2300 GNDA.n336 254.34
R881 GNDA.n2246 GNDA.n75 254.34
R882 GNDA.n2268 GNDA.n75 254.34
R883 GNDA.n2262 GNDA.n75 254.34
R884 GNDA.n2260 GNDA.n75 254.34
R885 GNDA.n2254 GNDA.n75 254.34
R886 GNDA.n2252 GNDA.n75 254.34
R887 GNDA.n880 GNDA.n75 254.34
R888 GNDA.n878 GNDA.n75 254.34
R889 GNDA.n887 GNDA.n75 254.34
R890 GNDA.n875 GNDA.n75 254.34
R891 GNDA.n894 GNDA.n75 254.34
R892 GNDA.n872 GNDA.n75 254.34
R893 GNDA.n645 GNDA.n72 254.34
R894 GNDA.n613 GNDA.n72 254.34
R895 GNDA.n634 GNDA.n72 254.34
R896 GNDA.n624 GNDA.n72 254.34
R897 GNDA.n622 GNDA.n72 254.34
R898 GNDA.n617 GNDA.n72 254.34
R899 GNDA.n2307 GNDA.n2306 254.34
R900 GNDA.n2306 GNDA.n323 254.34
R901 GNDA.n2306 GNDA.n322 254.34
R902 GNDA.n2306 GNDA.n321 254.34
R903 GNDA.n2306 GNDA.n320 254.34
R904 GNDA.n2306 GNDA.n319 254.34
R905 GNDA.n1480 GNDA.n71 254.34
R906 GNDA.n1477 GNDA.n71 254.34
R907 GNDA.n1471 GNDA.n71 254.34
R908 GNDA.n1468 GNDA.n71 254.34
R909 GNDA.n1463 GNDA.n71 254.34
R910 GNDA.n1460 GNDA.n71 254.34
R911 GNDA.n1501 GNDA.n69 254.34
R912 GNDA.n1459 GNDA.n69 254.34
R913 GNDA.n1494 GNDA.n69 254.34
R914 GNDA.n1488 GNDA.n69 254.34
R915 GNDA.n1486 GNDA.n69 254.34
R916 GNDA.n1474 GNDA.n69 254.34
R917 GNDA.n1535 GNDA.n66 254.34
R918 GNDA.n1533 GNDA.n66 254.34
R919 GNDA.n1523 GNDA.n66 254.34
R920 GNDA.n1521 GNDA.n66 254.34
R921 GNDA.n1512 GNDA.n66 254.34
R922 GNDA.n2399 GNDA.n66 254.34
R923 GNDA.n2395 GNDA.n65 254.34
R924 GNDA.n1515 GNDA.n65 254.34
R925 GNDA.n1517 GNDA.n65 254.34
R926 GNDA.n1527 GNDA.n65 254.34
R927 GNDA.n1529 GNDA.n65 254.34
R928 GNDA.n1539 GNDA.n65 254.34
R929 GNDA.n2159 GNDA.n2158 250.349
R930 GNDA.n710 GNDA.n709 250.349
R931 GNDA.t366 GNDA.n103 250.349
R932 GNDA.n2308 GNDA.n317 249.663
R933 GNDA.n2394 GNDA.n2393 249.663
R934 GNDA.n1502 GNDA.n1458 249.663
R935 GNDA.n2337 GNDA.n282 249.663
R936 GNDA.n2276 GNDA.n347 249.663
R937 GNDA.n2423 GNDA.n77 249.663
R938 GNDA.n1406 GNDA.n1404 249.663
R939 GNDA.n917 GNDA.n870 249.663
R940 GNDA.n2365 GNDA.n113 249.663
R941 GNDA.n394 GNDA.n393 246.25
R942 GNDA.n2177 GNDA.n393 246.25
R943 GNDA.n589 GNDA.n578 246.25
R944 GNDA.n582 GNDA.n578 246.25
R945 GNDA.n591 GNDA.n590 241.643
R946 GNDA.n591 GNDA.n577 241.643
R947 GNDA.n2187 GNDA.n2186 241.643
R948 GNDA.n2187 GNDA.n392 241.643
R949 GNDA.n2051 GNDA.t364 233
R950 GNDA.n2037 GNDA.t384 233
R951 GNDA.n2058 GNDA.n2057 199.883
R952 GNDA.n2086 GNDA.n2085 199.883
R953 GNDA.n2048 GNDA.n2047 199.03
R954 GNDA.n2046 GNDA.n2045 199.03
R955 GNDA.n2044 GNDA.n2043 199.03
R956 GNDA.n2042 GNDA.n2041 199.03
R957 GNDA.n2040 GNDA.n2039 199.03
R958 GNDA.n2380 GNDA.n102 197
R959 GNDA.n277 GNDA.n276 197
R960 GNDA.n1171 GNDA.n309 197
R961 GNDA.n682 GNDA.n331 197
R962 GNDA.n702 GNDA.n701 197
R963 GNDA.n2157 GNDA.n407 197
R964 GNDA.n1050 GNDA.n1049 197
R965 GNDA.n2132 GNDA.n486 197
R966 GNDA.n1658 GNDA.n1657 197
R967 GNDA.n1287 GNDA.n308 197
R968 GNDA.n795 GNDA.n565 197
R969 GNDA.n205 GNDA.n204 197
R970 GNDA.n1655 GNDA.n1654 187.249
R971 GNDA.n2312 GNDA.n311 187.249
R972 GNDA.n791 GNDA.n789 187.249
R973 GNDA.n2314 GNDA.n306 187.249
R974 GNDA.n431 GNDA.n335 187.249
R975 GNDA.n1753 GNDA.n1752 187.249
R976 GNDA.n1382 GNDA.n1381 187.249
R977 GNDA.n1781 GNDA.n851 187.249
R978 GNDA.n2341 GNDA.n2340 187.249
R979 GNDA.n1628 GNDA.n1627 185
R980 GNDA.n1630 GNDA.n1629 185
R981 GNDA.n1632 GNDA.n1631 185
R982 GNDA.n1634 GNDA.n1633 185
R983 GNDA.n1636 GNDA.n1635 185
R984 GNDA.n1638 GNDA.n1637 185
R985 GNDA.n1640 GNDA.n1639 185
R986 GNDA.n1642 GNDA.n1641 185
R987 GNDA.n1643 GNDA.n1541 185
R988 GNDA.n1610 GNDA.n1609 185
R989 GNDA.n1612 GNDA.n1611 185
R990 GNDA.n1614 GNDA.n1613 185
R991 GNDA.n1616 GNDA.n1615 185
R992 GNDA.n1618 GNDA.n1617 185
R993 GNDA.n1620 GNDA.n1619 185
R994 GNDA.n1622 GNDA.n1621 185
R995 GNDA.n1624 GNDA.n1623 185
R996 GNDA.n1626 GNDA.n1625 185
R997 GNDA.n1592 GNDA.n1591 185
R998 GNDA.n1594 GNDA.n1593 185
R999 GNDA.n1596 GNDA.n1595 185
R1000 GNDA.n1598 GNDA.n1597 185
R1001 GNDA.n1600 GNDA.n1599 185
R1002 GNDA.n1602 GNDA.n1601 185
R1003 GNDA.n1604 GNDA.n1603 185
R1004 GNDA.n1606 GNDA.n1605 185
R1005 GNDA.n1608 GNDA.n1607 185
R1006 GNDA.n257 GNDA.n256 185
R1007 GNDA.n259 GNDA.n258 185
R1008 GNDA.n261 GNDA.n260 185
R1009 GNDA.n263 GNDA.n262 185
R1010 GNDA.n265 GNDA.n264 185
R1011 GNDA.n267 GNDA.n266 185
R1012 GNDA.n269 GNDA.n268 185
R1013 GNDA.n271 GNDA.n270 185
R1014 GNDA.n272 GNDA.n20 185
R1015 GNDA.n239 GNDA.n238 185
R1016 GNDA.n241 GNDA.n240 185
R1017 GNDA.n243 GNDA.n242 185
R1018 GNDA.n245 GNDA.n244 185
R1019 GNDA.n247 GNDA.n246 185
R1020 GNDA.n249 GNDA.n248 185
R1021 GNDA.n251 GNDA.n250 185
R1022 GNDA.n253 GNDA.n252 185
R1023 GNDA.n255 GNDA.n254 185
R1024 GNDA.n221 GNDA.n220 185
R1025 GNDA.n223 GNDA.n222 185
R1026 GNDA.n225 GNDA.n224 185
R1027 GNDA.n227 GNDA.n226 185
R1028 GNDA.n229 GNDA.n228 185
R1029 GNDA.n231 GNDA.n230 185
R1030 GNDA.n233 GNDA.n232 185
R1031 GNDA.n235 GNDA.n234 185
R1032 GNDA.n237 GNDA.n236 185
R1033 GNDA.n1230 GNDA.n1169 185
R1034 GNDA.n1245 GNDA.n1244 185
R1035 GNDA.n1243 GNDA.n1170 185
R1036 GNDA.n1242 GNDA.n1241 185
R1037 GNDA.n1240 GNDA.n1239 185
R1038 GNDA.n1238 GNDA.n1237 185
R1039 GNDA.n1236 GNDA.n1235 185
R1040 GNDA.n1234 GNDA.n1233 185
R1041 GNDA.n1232 GNDA.n1231 185
R1042 GNDA.n1213 GNDA.n1212 185
R1043 GNDA.n1215 GNDA.n1214 185
R1044 GNDA.n1217 GNDA.n1216 185
R1045 GNDA.n1219 GNDA.n1218 185
R1046 GNDA.n1221 GNDA.n1220 185
R1047 GNDA.n1223 GNDA.n1222 185
R1048 GNDA.n1225 GNDA.n1224 185
R1049 GNDA.n1227 GNDA.n1226 185
R1050 GNDA.n1229 GNDA.n1228 185
R1051 GNDA.n1195 GNDA.n1194 185
R1052 GNDA.n1197 GNDA.n1196 185
R1053 GNDA.n1199 GNDA.n1198 185
R1054 GNDA.n1201 GNDA.n1200 185
R1055 GNDA.n1203 GNDA.n1202 185
R1056 GNDA.n1205 GNDA.n1204 185
R1057 GNDA.n1207 GNDA.n1206 185
R1058 GNDA.n1209 GNDA.n1208 185
R1059 GNDA.n1211 GNDA.n1210 185
R1060 GNDA.n1193 GNDA.n1192 185
R1061 GNDA.n1187 GNDA.n1186 185
R1062 GNDA.n1185 GNDA.n1184 185
R1063 GNDA.n1180 GNDA.n1179 185
R1064 GNDA.n1175 GNDA.n1154 185
R1065 GNDA.n1249 GNDA.n1248 185
R1066 GNDA.n1153 GNDA.n1151 185
R1067 GNDA.n1255 GNDA.n1254 185
R1068 GNDA.n1257 GNDA.n1256 185
R1069 GNDA.n754 GNDA.n676 185
R1070 GNDA.n768 GNDA.n767 185
R1071 GNDA.n766 GNDA.n677 185
R1072 GNDA.n765 GNDA.n764 185
R1073 GNDA.n763 GNDA.n762 185
R1074 GNDA.n761 GNDA.n760 185
R1075 GNDA.n759 GNDA.n758 185
R1076 GNDA.n757 GNDA.n756 185
R1077 GNDA.n755 GNDA.n650 185
R1078 GNDA.n737 GNDA.n736 185
R1079 GNDA.n739 GNDA.n738 185
R1080 GNDA.n741 GNDA.n740 185
R1081 GNDA.n743 GNDA.n742 185
R1082 GNDA.n745 GNDA.n744 185
R1083 GNDA.n747 GNDA.n746 185
R1084 GNDA.n749 GNDA.n748 185
R1085 GNDA.n751 GNDA.n750 185
R1086 GNDA.n753 GNDA.n752 185
R1087 GNDA.n719 GNDA.n718 185
R1088 GNDA.n721 GNDA.n720 185
R1089 GNDA.n723 GNDA.n722 185
R1090 GNDA.n725 GNDA.n724 185
R1091 GNDA.n727 GNDA.n726 185
R1092 GNDA.n729 GNDA.n728 185
R1093 GNDA.n731 GNDA.n730 185
R1094 GNDA.n733 GNDA.n732 185
R1095 GNDA.n735 GNDA.n734 185
R1096 GNDA.n717 GNDA.n716 185
R1097 GNDA.n692 GNDA.n691 185
R1098 GNDA.n690 GNDA.n689 185
R1099 GNDA.n687 GNDA.n661 185
R1100 GNDA.n774 GNDA.n773 185
R1101 GNDA.n771 GNDA.n660 185
R1102 GNDA.n770 GNDA.n654 185
R1103 GNDA.n783 GNDA.n782 185
R1104 GNDA.n785 GNDA.n784 185
R1105 GNDA.n2185 GNDA.n2184 185
R1106 GNDA.n2182 GNDA.n2181 185
R1107 GNDA.n586 GNDA.n398 185
R1108 GNDA.n586 GNDA.n579 185
R1109 GNDA.n580 GNDA.n398 185
R1110 GNDA.n584 GNDA.n580 185
R1111 GNDA.n1109 GNDA.n983 185
R1112 GNDA.n1124 GNDA.n1123 185
R1113 GNDA.n1122 GNDA.n984 185
R1114 GNDA.n1121 GNDA.n1120 185
R1115 GNDA.n1119 GNDA.n1118 185
R1116 GNDA.n1117 GNDA.n1116 185
R1117 GNDA.n1115 GNDA.n1114 185
R1118 GNDA.n1113 GNDA.n1112 185
R1119 GNDA.n1111 GNDA.n1110 185
R1120 GNDA.n1092 GNDA.n1091 185
R1121 GNDA.n1094 GNDA.n1093 185
R1122 GNDA.n1096 GNDA.n1095 185
R1123 GNDA.n1098 GNDA.n1097 185
R1124 GNDA.n1100 GNDA.n1099 185
R1125 GNDA.n1102 GNDA.n1101 185
R1126 GNDA.n1104 GNDA.n1103 185
R1127 GNDA.n1106 GNDA.n1105 185
R1128 GNDA.n1108 GNDA.n1107 185
R1129 GNDA.n1074 GNDA.n1073 185
R1130 GNDA.n1076 GNDA.n1075 185
R1131 GNDA.n1078 GNDA.n1077 185
R1132 GNDA.n1080 GNDA.n1079 185
R1133 GNDA.n1082 GNDA.n1081 185
R1134 GNDA.n1084 GNDA.n1083 185
R1135 GNDA.n1086 GNDA.n1085 185
R1136 GNDA.n1088 GNDA.n1087 185
R1137 GNDA.n1090 GNDA.n1089 185
R1138 GNDA.n1072 GNDA.n1071 185
R1139 GNDA.n1066 GNDA.n1065 185
R1140 GNDA.n1064 GNDA.n1063 185
R1141 GNDA.n1059 GNDA.n1058 185
R1142 GNDA.n1054 GNDA.n968 185
R1143 GNDA.n1128 GNDA.n1127 185
R1144 GNDA.n967 GNDA.n965 185
R1145 GNDA.n1134 GNDA.n1133 185
R1146 GNDA.n1136 GNDA.n1135 185
R1147 GNDA.n450 GNDA.n449 185
R1148 GNDA.n448 GNDA.n447 185
R1149 GNDA.n446 GNDA.n445 185
R1150 GNDA.n444 GNDA.n443 185
R1151 GNDA.n442 GNDA.n441 185
R1152 GNDA.n440 GNDA.n439 185
R1153 GNDA.n438 GNDA.n437 185
R1154 GNDA.n436 GNDA.n435 185
R1155 GNDA.n434 GNDA.n386 185
R1156 GNDA.n468 GNDA.n467 185
R1157 GNDA.n466 GNDA.n465 185
R1158 GNDA.n464 GNDA.n463 185
R1159 GNDA.n462 GNDA.n461 185
R1160 GNDA.n460 GNDA.n459 185
R1161 GNDA.n458 GNDA.n457 185
R1162 GNDA.n456 GNDA.n455 185
R1163 GNDA.n454 GNDA.n453 185
R1164 GNDA.n452 GNDA.n451 185
R1165 GNDA.n2136 GNDA.n2135 185
R1166 GNDA.n484 GNDA.n483 185
R1167 GNDA.n482 GNDA.n481 185
R1168 GNDA.n480 GNDA.n479 185
R1169 GNDA.n478 GNDA.n477 185
R1170 GNDA.n476 GNDA.n475 185
R1171 GNDA.n474 GNDA.n473 185
R1172 GNDA.n472 GNDA.n471 185
R1173 GNDA.n470 GNDA.n469 185
R1174 GNDA.n2138 GNDA.n2137 185
R1175 GNDA.n426 GNDA.n425 185
R1176 GNDA.n423 GNDA.n369 185
R1177 GNDA.n2208 GNDA.n2207 185
R1178 GNDA.n2191 GNDA.n368 185
R1179 GNDA.n2195 GNDA.n2194 185
R1180 GNDA.n2193 GNDA.n2190 185
R1181 GNDA.n389 GNDA.n387 185
R1182 GNDA.n2204 GNDA.n2203 185
R1183 GNDA.n1726 GNDA.n1725 185
R1184 GNDA.n1728 GNDA.n1727 185
R1185 GNDA.n1730 GNDA.n1729 185
R1186 GNDA.n1732 GNDA.n1731 185
R1187 GNDA.n1734 GNDA.n1733 185
R1188 GNDA.n1736 GNDA.n1735 185
R1189 GNDA.n1738 GNDA.n1737 185
R1190 GNDA.n1740 GNDA.n1739 185
R1191 GNDA.n1741 GNDA.n921 185
R1192 GNDA.n1708 GNDA.n1707 185
R1193 GNDA.n1710 GNDA.n1709 185
R1194 GNDA.n1712 GNDA.n1711 185
R1195 GNDA.n1714 GNDA.n1713 185
R1196 GNDA.n1716 GNDA.n1715 185
R1197 GNDA.n1718 GNDA.n1717 185
R1198 GNDA.n1720 GNDA.n1719 185
R1199 GNDA.n1722 GNDA.n1721 185
R1200 GNDA.n1724 GNDA.n1723 185
R1201 GNDA.n1690 GNDA.n1689 185
R1202 GNDA.n1692 GNDA.n1691 185
R1203 GNDA.n1694 GNDA.n1693 185
R1204 GNDA.n1696 GNDA.n1695 185
R1205 GNDA.n1698 GNDA.n1697 185
R1206 GNDA.n1700 GNDA.n1699 185
R1207 GNDA.n1702 GNDA.n1701 185
R1208 GNDA.n1704 GNDA.n1703 185
R1209 GNDA.n1706 GNDA.n1705 185
R1210 GNDA.n1688 GNDA.n1687 185
R1211 GNDA.n1682 GNDA.n1681 185
R1212 GNDA.n1680 GNDA.n1679 185
R1213 GNDA.n1675 GNDA.n1674 185
R1214 GNDA.n1673 GNDA.n1672 185
R1215 GNDA.n1667 GNDA.n1666 185
R1216 GNDA.n1662 GNDA.n925 185
R1217 GNDA.n1745 GNDA.n1744 185
R1218 GNDA.n924 GNDA.n922 185
R1219 GNDA.n1354 GNDA.n1353 185
R1220 GNDA.n1356 GNDA.n1355 185
R1221 GNDA.n1358 GNDA.n1357 185
R1222 GNDA.n1360 GNDA.n1359 185
R1223 GNDA.n1362 GNDA.n1361 185
R1224 GNDA.n1364 GNDA.n1363 185
R1225 GNDA.n1366 GNDA.n1365 185
R1226 GNDA.n1367 GNDA.n1286 185
R1227 GNDA.n1371 GNDA.n1370 185
R1228 GNDA.n1336 GNDA.n1335 185
R1229 GNDA.n1338 GNDA.n1337 185
R1230 GNDA.n1340 GNDA.n1339 185
R1231 GNDA.n1342 GNDA.n1341 185
R1232 GNDA.n1344 GNDA.n1343 185
R1233 GNDA.n1346 GNDA.n1345 185
R1234 GNDA.n1348 GNDA.n1347 185
R1235 GNDA.n1350 GNDA.n1349 185
R1236 GNDA.n1352 GNDA.n1351 185
R1237 GNDA.n1318 GNDA.n1317 185
R1238 GNDA.n1320 GNDA.n1319 185
R1239 GNDA.n1322 GNDA.n1321 185
R1240 GNDA.n1324 GNDA.n1323 185
R1241 GNDA.n1326 GNDA.n1325 185
R1242 GNDA.n1328 GNDA.n1327 185
R1243 GNDA.n1330 GNDA.n1329 185
R1244 GNDA.n1332 GNDA.n1331 185
R1245 GNDA.n1334 GNDA.n1333 185
R1246 GNDA.n1316 GNDA.n1315 185
R1247 GNDA.n1310 GNDA.n1309 185
R1248 GNDA.n1308 GNDA.n1307 185
R1249 GNDA.n1303 GNDA.n1302 185
R1250 GNDA.n1301 GNDA.n1300 185
R1251 GNDA.n1295 GNDA.n1294 185
R1252 GNDA.n1291 GNDA.n1269 185
R1253 GNDA.n1375 GNDA.n1374 185
R1254 GNDA.n1268 GNDA.n1266 185
R1255 GNDA.n834 GNDA.n833 185
R1256 GNDA.n835 GNDA.n549 185
R1257 GNDA.n837 GNDA.n836 185
R1258 GNDA.n839 GNDA.n548 185
R1259 GNDA.n842 GNDA.n841 185
R1260 GNDA.n843 GNDA.n547 185
R1261 GNDA.n845 GNDA.n844 185
R1262 GNDA.n847 GNDA.n546 185
R1263 GNDA.n849 GNDA.n848 185
R1264 GNDA.n815 GNDA.n554 185
R1265 GNDA.n818 GNDA.n817 185
R1266 GNDA.n819 GNDA.n553 185
R1267 GNDA.n821 GNDA.n820 185
R1268 GNDA.n823 GNDA.n552 185
R1269 GNDA.n826 GNDA.n825 185
R1270 GNDA.n827 GNDA.n551 185
R1271 GNDA.n829 GNDA.n828 185
R1272 GNDA.n831 GNDA.n550 185
R1273 GNDA.n799 GNDA.n798 185
R1274 GNDA.n801 GNDA.n559 185
R1275 GNDA.n803 GNDA.n802 185
R1276 GNDA.n804 GNDA.n558 185
R1277 GNDA.n806 GNDA.n805 185
R1278 GNDA.n808 GNDA.n556 185
R1279 GNDA.n810 GNDA.n809 185
R1280 GNDA.n811 GNDA.n555 185
R1281 GNDA.n813 GNDA.n812 185
R1282 GNDA.n604 GNDA.n561 185
R1283 GNDA.n603 GNDA.n602 185
R1284 GNDA.n600 GNDA.n568 185
R1285 GNDA.n598 GNDA.n597 185
R1286 GNDA.n574 GNDA.n570 185
R1287 GNDA.n572 GNDA.n544 185
R1288 GNDA.n1794 GNDA.n1793 185
R1289 GNDA.n1791 GNDA.n542 185
R1290 GNDA.n1790 GNDA.n1789 185
R1291 GNDA.n219 GNDA.n218 185
R1292 GNDA.n213 GNDA.n212 185
R1293 GNDA.n208 GNDA.n3 185
R1294 GNDA.n2435 GNDA.n2434 185
R1295 GNDA.n39 GNDA.n2 185
R1296 GNDA.n43 GNDA.n42 185
R1297 GNDA.n41 GNDA.n38 185
R1298 GNDA.n23 GNDA.n21 185
R1299 GNDA.n2431 GNDA.n2430 185
R1300 GNDA.n1590 GNDA.n1589 185
R1301 GNDA.n1584 GNDA.n1583 185
R1302 GNDA.n1582 GNDA.n1581 185
R1303 GNDA.n1577 GNDA.n1576 185
R1304 GNDA.n1575 GNDA.n1574 185
R1305 GNDA.n1569 GNDA.n1568 185
R1306 GNDA.n1564 GNDA.n1545 185
R1307 GNDA.n1647 GNDA.n1646 185
R1308 GNDA.n1544 GNDA.n1542 185
R1309 GNDA.t130 GNDA.t363 182.07
R1310 GNDA.t394 GNDA.t11 182.07
R1311 GNDA.t30 GNDA.t402 182.07
R1312 GNDA.t383 GNDA.t8 182.07
R1313 GNDA.n619 GNDA.n318 175.546
R1314 GNDA.n627 GNDA.n626 175.546
R1315 GNDA.n631 GNDA.n630 175.546
R1316 GNDA.n638 GNDA.n637 175.546
R1317 GNDA.n641 GNDA.n640 175.546
R1318 GNDA.n2255 GNDA.n2253 175.546
R1319 GNDA.n2259 GNDA.n2250 175.546
R1320 GNDA.n2263 GNDA.n2261 175.546
R1321 GNDA.n2267 GNDA.n2248 175.546
R1322 GNDA.n2270 GNDA.n2269 175.546
R1323 GNDA.n346 GNDA.n345 175.546
R1324 GNDA.n2284 GNDA.n2283 175.546
R1325 GNDA.n342 GNDA.n341 175.546
R1326 GNDA.n2294 GNDA.n2293 175.546
R1327 GNDA.n337 GNDA.n330 175.546
R1328 GNDA.n2396 GNDA.n92 175.546
R1329 GNDA.n1518 GNDA.n1516 175.546
R1330 GNDA.n1526 GNDA.n1510 175.546
R1331 GNDA.n1530 GNDA.n1528 175.546
R1332 GNDA.n1538 GNDA.n1506 175.546
R1333 GNDA.n2393 GNDA.n93 175.546
R1334 GNDA.n2389 GNDA.n93 175.546
R1335 GNDA.n2389 GNDA.n96 175.546
R1336 GNDA.n2385 GNDA.n96 175.546
R1337 GNDA.n2385 GNDA.n99 175.546
R1338 GNDA.n2378 GNDA.n99 175.546
R1339 GNDA.n2378 GNDA.n2377 175.546
R1340 GNDA.n2377 GNDA.n105 175.546
R1341 GNDA.n2373 GNDA.n105 175.546
R1342 GNDA.n2373 GNDA.n107 175.546
R1343 GNDA.n2369 GNDA.n107 175.546
R1344 GNDA.n115 GNDA.n110 175.546
R1345 GNDA.n116 GNDA.n115 175.546
R1346 GNDA.n119 GNDA.n116 175.546
R1347 GNDA.n120 GNDA.n119 175.546
R1348 GNDA.n123 GNDA.n120 175.546
R1349 GNDA.n124 GNDA.n123 175.546
R1350 GNDA.n125 GNDA.n124 175.546
R1351 GNDA.n126 GNDA.n125 175.546
R1352 GNDA.n130 GNDA.n126 175.546
R1353 GNDA.n131 GNDA.n130 175.546
R1354 GNDA.n133 GNDA.n131 175.546
R1355 GNDA.n1650 GNDA.n1649 175.546
R1356 GNDA.n1566 GNDA.n1565 175.546
R1357 GNDA.n1572 GNDA.n1571 175.546
R1358 GNDA.n1579 GNDA.n1578 175.546
R1359 GNDA.n1587 GNDA.n1586 175.546
R1360 GNDA.n286 GNDA.n285 175.546
R1361 GNDA.n291 GNDA.n288 175.546
R1362 GNDA.n294 GNDA.n293 175.546
R1363 GNDA.n299 GNDA.n296 175.546
R1364 GNDA.n302 GNDA.n301 175.546
R1365 GNDA.n1500 GNDA.n1499 175.546
R1366 GNDA.n1496 GNDA.n1495 175.546
R1367 GNDA.n1493 GNDA.n1466 175.546
R1368 GNDA.n1489 GNDA.n1487 175.546
R1369 GNDA.n1485 GNDA.n1475 175.546
R1370 GNDA.n1456 GNDA.n1431 175.546
R1371 GNDA.n1452 GNDA.n1451 175.546
R1372 GNDA.n1449 GNDA.n1434 175.546
R1373 GNDA.n1445 GNDA.n1444 175.546
R1374 GNDA.n1442 GNDA.n1439 175.546
R1375 GNDA.n1259 GNDA.n1145 175.546
R1376 GNDA.n1252 GNDA.n1251 175.546
R1377 GNDA.n1177 GNDA.n1176 175.546
R1378 GNDA.n1182 GNDA.n1181 175.546
R1379 GNDA.n1190 GNDA.n1189 175.546
R1380 GNDA.n789 GNDA.n649 175.546
R1381 GNDA.n655 GNDA.n649 175.546
R1382 GNDA.n780 GNDA.n655 175.546
R1383 GNDA.n780 GNDA.n656 175.546
R1384 GNDA.n776 GNDA.n656 175.546
R1385 GNDA.n776 GNDA.n658 175.546
R1386 GNDA.n685 GNDA.n658 175.546
R1387 GNDA.n694 GNDA.n685 175.546
R1388 GNDA.n694 GNDA.n680 175.546
R1389 GNDA.n714 GNDA.n680 175.546
R1390 GNDA.n714 GNDA.n682 175.546
R1391 GNDA.n2335 GNDA.n2334 175.546
R1392 GNDA.n2331 GNDA.n2330 175.546
R1393 GNDA.n2328 GNDA.n290 175.546
R1394 GNDA.n2324 GNDA.n2322 175.546
R1395 GNDA.n2320 GNDA.n298 175.546
R1396 GNDA.n1005 GNDA.n1002 175.546
R1397 GNDA.n1009 GNDA.n1007 175.546
R1398 GNDA.n1013 GNDA.n999 175.546
R1399 GNDA.n1016 GNDA.n1015 175.546
R1400 GNDA.n1020 GNDA.n1019 175.546
R1401 GNDA.n1138 GNDA.n959 175.546
R1402 GNDA.n1131 GNDA.n1130 175.546
R1403 GNDA.n1056 GNDA.n1055 175.546
R1404 GNDA.n1061 GNDA.n1060 175.546
R1405 GNDA.n1069 GNDA.n1068 175.546
R1406 GNDA.n1026 GNDA.n995 175.546
R1407 GNDA.n1026 GNDA.n993 175.546
R1408 GNDA.n1031 GNDA.n993 175.546
R1409 GNDA.n1031 GNDA.n991 175.546
R1410 GNDA.n1035 GNDA.n991 175.546
R1411 GNDA.n1036 GNDA.n1035 175.546
R1412 GNDA.n1038 GNDA.n1036 175.546
R1413 GNDA.n1038 GNDA.n989 175.546
R1414 GNDA.n1043 GNDA.n989 175.546
R1415 GNDA.n1043 GNDA.n987 175.546
R1416 GNDA.n1047 GNDA.n987 175.546
R1417 GNDA.n2280 GNDA.n2278 175.546
R1418 GNDA.n2286 GNDA.n343 175.546
R1419 GNDA.n2290 GNDA.n2288 175.546
R1420 GNDA.n2296 GNDA.n339 175.546
R1421 GNDA.n2299 GNDA.n2298 175.546
R1422 GNDA.n2242 GNDA.n2241 175.546
R1423 GNDA.n2239 GNDA.n350 175.546
R1424 GNDA.n2235 GNDA.n2234 175.546
R1425 GNDA.n2232 GNDA.n353 175.546
R1426 GNDA.n2228 GNDA.n2227 175.546
R1427 GNDA.n431 GNDA.n390 175.546
R1428 GNDA.n2201 GNDA.n390 175.546
R1429 GNDA.n2201 GNDA.n391 175.546
R1430 GNDA.n2197 GNDA.n391 175.546
R1431 GNDA.n2197 GNDA.n365 175.546
R1432 GNDA.n2210 GNDA.n365 175.546
R1433 GNDA.n2210 GNDA.n366 175.546
R1434 GNDA.n421 GNDA.n366 175.546
R1435 GNDA.n2140 GNDA.n421 175.546
R1436 GNDA.n2140 GNDA.n422 175.546
R1437 GNDA.n2132 GNDA.n422 175.546
R1438 GNDA.n2221 GNDA.n356 175.546
R1439 GNDA.n2221 GNDA.n358 175.546
R1440 GNDA.n2217 GNDA.n358 175.546
R1441 GNDA.n2217 GNDA.n361 175.546
R1442 GNDA.n2213 GNDA.n361 175.546
R1443 GNDA.n2213 GNDA.n363 175.546
R1444 GNDA.n490 GNDA.n363 175.546
R1445 GNDA.n494 GNDA.n490 175.546
R1446 GNDA.n494 GNDA.n488 175.546
R1447 GNDA.n498 GNDA.n488 175.546
R1448 GNDA.n500 GNDA.n498 175.546
R1449 GNDA.n2398 GNDA.n90 175.546
R1450 GNDA.n1520 GNDA.n1513 175.546
R1451 GNDA.n1524 GNDA.n1522 175.546
R1452 GNDA.n1532 GNDA.n1508 175.546
R1453 GNDA.n1536 GNDA.n1534 175.546
R1454 GNDA.n2423 GNDA.n78 175.546
R1455 GNDA.n2419 GNDA.n78 175.546
R1456 GNDA.n2419 GNDA.n81 175.546
R1457 GNDA.n2415 GNDA.n81 175.546
R1458 GNDA.n2415 GNDA.n83 175.546
R1459 GNDA.n2411 GNDA.n83 175.546
R1460 GNDA.n2411 GNDA.n85 175.546
R1461 GNDA.n2407 GNDA.n85 175.546
R1462 GNDA.n2407 GNDA.n87 175.546
R1463 GNDA.n2403 GNDA.n87 175.546
R1464 GNDA.n2403 GNDA.n2401 175.546
R1465 GNDA.n1748 GNDA.n1747 175.546
R1466 GNDA.n1664 GNDA.n1663 175.546
R1467 GNDA.n1670 GNDA.n1669 175.546
R1468 GNDA.n1677 GNDA.n1676 175.546
R1469 GNDA.n1685 GNDA.n1684 175.546
R1470 GNDA.n1774 GNDA.n920 175.546
R1471 GNDA.n1770 GNDA.n920 175.546
R1472 GNDA.n1768 GNDA.n1767 175.546
R1473 GNDA.n1764 GNDA.n1763 175.546
R1474 GNDA.n1760 GNDA.n1759 175.546
R1475 GNDA.n1756 GNDA.n1755 175.546
R1476 GNDA.n1462 GNDA.n1461 175.546
R1477 GNDA.n1467 GNDA.n1464 175.546
R1478 GNDA.n1470 GNDA.n1469 175.546
R1479 GNDA.n1476 GNDA.n1472 175.546
R1480 GNDA.n1479 GNDA.n1478 175.546
R1481 GNDA.n1410 GNDA.n950 175.546
R1482 GNDA.n1414 GNDA.n1412 175.546
R1483 GNDA.n1418 GNDA.n948 175.546
R1484 GNDA.n1422 GNDA.n1420 175.546
R1485 GNDA.n1426 GNDA.n946 175.546
R1486 GNDA.n1377 GNDA.n953 175.546
R1487 GNDA.n1292 GNDA.n1265 175.546
R1488 GNDA.n1298 GNDA.n1297 175.546
R1489 GNDA.n1305 GNDA.n1304 175.546
R1490 GNDA.n1313 GNDA.n1312 175.546
R1491 GNDA.n1401 GNDA.n1400 175.546
R1492 GNDA.n1397 GNDA.n1396 175.546
R1493 GNDA.n1393 GNDA.n1392 175.546
R1494 GNDA.n1389 GNDA.n1388 175.546
R1495 GNDA.n1385 GNDA.n864 175.546
R1496 GNDA.n951 GNDA.n864 175.546
R1497 GNDA.n621 GNDA.n618 175.546
R1498 GNDA.n625 GNDA.n623 175.546
R1499 GNDA.n633 GNDA.n615 175.546
R1500 GNDA.n636 GNDA.n635 175.546
R1501 GNDA.n644 GNDA.n643 175.546
R1502 GNDA.n896 GNDA.n895 175.546
R1503 GNDA.n893 GNDA.n873 175.546
R1504 GNDA.n889 GNDA.n888 175.546
R1505 GNDA.n886 GNDA.n876 175.546
R1506 GNDA.n882 GNDA.n881 175.546
R1507 GNDA.n1786 GNDA.n1781 175.546
R1508 GNDA.n1786 GNDA.n539 175.546
R1509 GNDA.n1796 GNDA.n539 175.546
R1510 GNDA.n1796 GNDA.n541 175.546
R1511 GNDA.n571 GNDA.n541 175.546
R1512 GNDA.n576 GNDA.n571 175.546
R1513 GNDA.n595 GNDA.n576 175.546
R1514 GNDA.n595 GNDA.n566 175.546
R1515 GNDA.n606 GNDA.n566 175.546
R1516 GNDA.n606 GNDA.n564 175.546
R1517 GNDA.n795 GNDA.n564 175.546
R1518 GNDA.n913 GNDA.n869 175.546
R1519 GNDA.n911 GNDA.n910 175.546
R1520 GNDA.n907 GNDA.n906 175.546
R1521 GNDA.n903 GNDA.n902 175.546
R1522 GNDA.n899 GNDA.n853 175.546
R1523 GNDA.n1778 GNDA.n853 175.546
R1524 GNDA.n179 GNDA.n143 175.546
R1525 GNDA.n183 GNDA.n143 175.546
R1526 GNDA.n183 GNDA.n141 175.546
R1527 GNDA.n187 GNDA.n141 175.546
R1528 GNDA.n187 GNDA.n139 175.546
R1529 GNDA.n191 GNDA.n139 175.546
R1530 GNDA.n192 GNDA.n191 175.546
R1531 GNDA.n196 GNDA.n192 175.546
R1532 GNDA.n196 GNDA.n137 175.546
R1533 GNDA.n200 GNDA.n137 175.546
R1534 GNDA.n201 GNDA.n200 175.546
R1535 GNDA.n2428 GNDA.n24 175.546
R1536 GNDA.n45 GNDA.n25 175.546
R1537 GNDA.n36 GNDA.n35 175.546
R1538 GNDA.n210 GNDA.n209 175.546
R1539 GNDA.n216 GNDA.n215 175.546
R1540 GNDA.n2365 GNDA.n114 175.546
R1541 GNDA.n2361 GNDA.n114 175.546
R1542 GNDA.n2361 GNDA.n118 175.546
R1543 GNDA.n2357 GNDA.n118 175.546
R1544 GNDA.n2357 GNDA.n2355 175.546
R1545 GNDA.n2355 GNDA.n2354 175.546
R1546 GNDA.n2354 GNDA.n122 175.546
R1547 GNDA.n2350 GNDA.n122 175.546
R1548 GNDA.n2350 GNDA.n128 175.546
R1549 GNDA.n2346 GNDA.n128 175.546
R1550 GNDA.n2346 GNDA.n132 175.546
R1551 GNDA.n155 GNDA.n113 175.546
R1552 GNDA.n158 GNDA.n155 175.546
R1553 GNDA.n158 GNDA.n152 175.546
R1554 GNDA.n163 GNDA.n152 175.546
R1555 GNDA.n163 GNDA.n150 175.546
R1556 GNDA.n167 GNDA.n150 175.546
R1557 GNDA.n167 GNDA.n149 175.546
R1558 GNDA.n171 GNDA.n149 175.546
R1559 GNDA.n171 GNDA.n147 175.546
R1560 GNDA.n175 GNDA.n147 175.546
R1561 GNDA.n175 GNDA.n145 175.546
R1562 GNDA.t366 GNDA.n71 172.876
R1563 GNDA.t366 GNDA.n68 172.876
R1564 GNDA.t366 GNDA.n66 172.876
R1565 GNDA.t366 GNDA.n69 172.615
R1566 GNDA.t366 GNDA.n70 172.615
R1567 GNDA.t366 GNDA.n65 172.615
R1568 GNDA.t210 GNDA.n2035 166.898
R1569 GNDA.n1591 GNDA.n1590 163.333
R1570 GNDA.n220 GNDA.n219 163.333
R1571 GNDA.n1194 GNDA.n1193 163.333
R1572 GNDA.n718 GNDA.n717 163.333
R1573 GNDA.n1073 GNDA.n1072 163.333
R1574 GNDA.n2137 GNDA.n2136 163.333
R1575 GNDA.n1689 GNDA.n1688 163.333
R1576 GNDA.n1317 GNDA.n1316 163.333
R1577 GNDA.n799 GNDA.n561 163.333
R1578 GNDA.n2016 GNDA.n2015 161.3
R1579 GNDA.n2022 GNDA.n2021 161.3
R1580 GNDA.t366 GNDA.n64 159.365
R1581 GNDA.n2370 GNDA.n109 159.365
R1582 GNDA.t366 GNDA.n63 155.957
R1583 GNDA.n153 GNDA.n109 155.957
R1584 GNDA.t363 GNDA.t111 151.725
R1585 GNDA.t11 GNDA.t130 151.725
R1586 GNDA.t324 GNDA.t394 151.725
R1587 GNDA.n2034 GNDA.t26 151.725
R1588 GNDA.t402 GNDA.t551 151.725
R1589 GNDA.t8 GNDA.t30 151.725
R1590 GNDA.t59 GNDA.t383 151.725
R1591 GNDA.n1623 GNDA.n1622 150
R1592 GNDA.n1619 GNDA.n1618 150
R1593 GNDA.n1615 GNDA.n1614 150
R1594 GNDA.n1611 GNDA.n1610 150
R1595 GNDA.n1607 GNDA.n1606 150
R1596 GNDA.n1603 GNDA.n1602 150
R1597 GNDA.n1599 GNDA.n1598 150
R1598 GNDA.n1595 GNDA.n1594 150
R1599 GNDA.n1646 GNDA.n1544 150
R1600 GNDA.n1568 GNDA.n1545 150
R1601 GNDA.n1576 GNDA.n1575 150
R1602 GNDA.n1583 GNDA.n1582 150
R1603 GNDA.n1631 GNDA.n1630 150
R1604 GNDA.n1635 GNDA.n1634 150
R1605 GNDA.n1639 GNDA.n1638 150
R1606 GNDA.n1643 GNDA.n1642 150
R1607 GNDA.n252 GNDA.n251 150
R1608 GNDA.n248 GNDA.n247 150
R1609 GNDA.n244 GNDA.n243 150
R1610 GNDA.n240 GNDA.n239 150
R1611 GNDA.n236 GNDA.n235 150
R1612 GNDA.n232 GNDA.n231 150
R1613 GNDA.n228 GNDA.n227 150
R1614 GNDA.n224 GNDA.n223 150
R1615 GNDA.n2431 GNDA.n21 150
R1616 GNDA.n42 GNDA.n41 150
R1617 GNDA.n2434 GNDA.n2 150
R1618 GNDA.n212 GNDA.n3 150
R1619 GNDA.n260 GNDA.n259 150
R1620 GNDA.n264 GNDA.n263 150
R1621 GNDA.n268 GNDA.n267 150
R1622 GNDA.n270 GNDA.n20 150
R1623 GNDA.n1226 GNDA.n1225 150
R1624 GNDA.n1222 GNDA.n1221 150
R1625 GNDA.n1218 GNDA.n1217 150
R1626 GNDA.n1214 GNDA.n1213 150
R1627 GNDA.n1210 GNDA.n1209 150
R1628 GNDA.n1206 GNDA.n1205 150
R1629 GNDA.n1202 GNDA.n1201 150
R1630 GNDA.n1198 GNDA.n1197 150
R1631 GNDA.n1256 GNDA.n1255 150
R1632 GNDA.n1248 GNDA.n1153 150
R1633 GNDA.n1179 GNDA.n1154 150
R1634 GNDA.n1186 GNDA.n1185 150
R1635 GNDA.n1245 GNDA.n1170 150
R1636 GNDA.n1241 GNDA.n1240 150
R1637 GNDA.n1237 GNDA.n1236 150
R1638 GNDA.n1233 GNDA.n1232 150
R1639 GNDA.n750 GNDA.n749 150
R1640 GNDA.n746 GNDA.n745 150
R1641 GNDA.n742 GNDA.n741 150
R1642 GNDA.n738 GNDA.n737 150
R1643 GNDA.n734 GNDA.n733 150
R1644 GNDA.n730 GNDA.n729 150
R1645 GNDA.n726 GNDA.n725 150
R1646 GNDA.n722 GNDA.n721 150
R1647 GNDA.n784 GNDA.n783 150
R1648 GNDA.n771 GNDA.n770 150
R1649 GNDA.n773 GNDA.n661 150
R1650 GNDA.n691 GNDA.n690 150
R1651 GNDA.n768 GNDA.n677 150
R1652 GNDA.n764 GNDA.n763 150
R1653 GNDA.n760 GNDA.n759 150
R1654 GNDA.n756 GNDA.n755 150
R1655 GNDA.n1105 GNDA.n1104 150
R1656 GNDA.n1101 GNDA.n1100 150
R1657 GNDA.n1097 GNDA.n1096 150
R1658 GNDA.n1093 GNDA.n1092 150
R1659 GNDA.n1089 GNDA.n1088 150
R1660 GNDA.n1085 GNDA.n1084 150
R1661 GNDA.n1081 GNDA.n1080 150
R1662 GNDA.n1077 GNDA.n1076 150
R1663 GNDA.n1135 GNDA.n1134 150
R1664 GNDA.n1127 GNDA.n967 150
R1665 GNDA.n1058 GNDA.n968 150
R1666 GNDA.n1065 GNDA.n1064 150
R1667 GNDA.n1124 GNDA.n984 150
R1668 GNDA.n1120 GNDA.n1119 150
R1669 GNDA.n1116 GNDA.n1115 150
R1670 GNDA.n1112 GNDA.n1111 150
R1671 GNDA.n455 GNDA.n454 150
R1672 GNDA.n459 GNDA.n458 150
R1673 GNDA.n463 GNDA.n462 150
R1674 GNDA.n467 GNDA.n466 150
R1675 GNDA.n471 GNDA.n470 150
R1676 GNDA.n475 GNDA.n474 150
R1677 GNDA.n479 GNDA.n478 150
R1678 GNDA.n483 GNDA.n482 150
R1679 GNDA.n2204 GNDA.n387 150
R1680 GNDA.n2194 GNDA.n2193 150
R1681 GNDA.n2207 GNDA.n368 150
R1682 GNDA.n425 GNDA.n369 150
R1683 GNDA.n447 GNDA.n446 150
R1684 GNDA.n443 GNDA.n442 150
R1685 GNDA.n439 GNDA.n438 150
R1686 GNDA.n435 GNDA.n386 150
R1687 GNDA.n1721 GNDA.n1720 150
R1688 GNDA.n1717 GNDA.n1716 150
R1689 GNDA.n1713 GNDA.n1712 150
R1690 GNDA.n1709 GNDA.n1708 150
R1691 GNDA.n1705 GNDA.n1704 150
R1692 GNDA.n1701 GNDA.n1700 150
R1693 GNDA.n1697 GNDA.n1696 150
R1694 GNDA.n1693 GNDA.n1692 150
R1695 GNDA.n1744 GNDA.n924 150
R1696 GNDA.n1666 GNDA.n925 150
R1697 GNDA.n1674 GNDA.n1673 150
R1698 GNDA.n1681 GNDA.n1680 150
R1699 GNDA.n1729 GNDA.n1728 150
R1700 GNDA.n1733 GNDA.n1732 150
R1701 GNDA.n1737 GNDA.n1736 150
R1702 GNDA.n1741 GNDA.n1740 150
R1703 GNDA.n1349 GNDA.n1348 150
R1704 GNDA.n1345 GNDA.n1344 150
R1705 GNDA.n1341 GNDA.n1340 150
R1706 GNDA.n1337 GNDA.n1336 150
R1707 GNDA.n1333 GNDA.n1332 150
R1708 GNDA.n1329 GNDA.n1328 150
R1709 GNDA.n1325 GNDA.n1324 150
R1710 GNDA.n1321 GNDA.n1320 150
R1711 GNDA.n1374 GNDA.n1268 150
R1712 GNDA.n1294 GNDA.n1269 150
R1713 GNDA.n1302 GNDA.n1301 150
R1714 GNDA.n1309 GNDA.n1308 150
R1715 GNDA.n1357 GNDA.n1356 150
R1716 GNDA.n1361 GNDA.n1360 150
R1717 GNDA.n1365 GNDA.n1364 150
R1718 GNDA.n1371 GNDA.n1286 150
R1719 GNDA.n829 GNDA.n551 150
R1720 GNDA.n825 GNDA.n823 150
R1721 GNDA.n821 GNDA.n553 150
R1722 GNDA.n817 GNDA.n815 150
R1723 GNDA.n813 GNDA.n555 150
R1724 GNDA.n809 GNDA.n808 150
R1725 GNDA.n806 GNDA.n558 150
R1726 GNDA.n802 GNDA.n801 150
R1727 GNDA.n1791 GNDA.n1790 150
R1728 GNDA.n1793 GNDA.n544 150
R1729 GNDA.n598 GNDA.n570 150
R1730 GNDA.n602 GNDA.n600 150
R1731 GNDA.n837 GNDA.n549 150
R1732 GNDA.n841 GNDA.n839 150
R1733 GNDA.n845 GNDA.n547 150
R1734 GNDA.n848 GNDA.n847 150
R1735 GNDA.n1993 GNDA.n529 148.017
R1736 GNDA.n1998 GNDA.n1997 148.017
R1737 GNDA.n2118 GNDA.n2117 148.017
R1738 GNDA.n2123 GNDA.n2122 148.017
R1739 GNDA.n2145 GNDA.n417 136.145
R1740 GNDA.n2146 GNDA.n416 136.145
R1741 GNDA.n2147 GNDA.n415 136.145
R1742 GNDA.n2150 GNDA.n412 136.145
R1743 GNDA.n2151 GNDA.n411 136.145
R1744 GNDA.n1804 GNDA.n1803 136.145
R1745 GNDA.n1805 GNDA.n1802 136.145
R1746 GNDA.n1806 GNDA.n1801 136.145
R1747 GNDA.n1809 GNDA.n536 136.145
R1748 GNDA.n1810 GNDA.n535 136.145
R1749 GNDA.n587 GNDA.n586 134.268
R1750 GNDA.n587 GNDA.n580 134.268
R1751 GNDA.n2143 GNDA.t450 130.001
R1752 GNDA.n698 GNDA.t406 130.001
R1753 GNDA.n711 GNDA.t463 130.001
R1754 GNDA.n2154 GNDA.t414 130.001
R1755 GNDA.n610 GNDA.t374 130.001
R1756 GNDA.n1799 GNDA.t453 130.001
R1757 GNDA.n1783 GNDA.t431 130.001
R1758 GNDA.n1812 GNDA.t371 130.001
R1759 GNDA.n791 GNDA.n648 124.832
R1760 GNDA.n2303 GNDA.n331 124.832
R1761 GNDA.n1655 GNDA.n1540 124.832
R1762 GNDA.n277 GNDA.n133 124.832
R1763 GNDA.n309 GNDA.n304 124.832
R1764 GNDA.n2312 GNDA.n310 124.832
R1765 GNDA.n2316 GNDA.n2314 124.832
R1766 GNDA.n2301 GNDA.n335 124.832
R1767 GNDA.n1657 GNDA.n943 124.832
R1768 GNDA.n1481 GNDA.n308 124.832
R1769 GNDA.n646 GNDA.n565 124.832
R1770 GNDA.n2341 GNDA.n132 124.832
R1771 GNDA.n2097 GNDA.n2095 124.59
R1772 GNDA.n1823 GNDA.n1821 124.59
R1773 GNDA.n2105 GNDA.n2104 124.028
R1774 GNDA.n2103 GNDA.n2102 124.028
R1775 GNDA.n2101 GNDA.n2100 124.028
R1776 GNDA.n2099 GNDA.n2098 124.028
R1777 GNDA.n2097 GNDA.n2096 124.028
R1778 GNDA.n1831 GNDA.n1830 124.028
R1779 GNDA.n1829 GNDA.n1828 124.028
R1780 GNDA.n1827 GNDA.n1826 124.028
R1781 GNDA.n1825 GNDA.n1824 124.028
R1782 GNDA.n1823 GNDA.n1822 124.028
R1783 GNDA.n1929 GNDA.t282 116.073
R1784 GNDA.n1912 GNDA.t292 115.105
R1785 GNDA.n1911 GNDA.t166 114.635
R1786 GNDA.n1929 GNDA.t256 114.635
R1787 GNDA.n986 GNDA.n359 102.812
R1788 GNDA.n2177 GNDA.n392 101.718
R1789 GNDA.n582 GNDA.n577 101.718
R1790 GNDA.n590 GNDA.n589 101.718
R1791 GNDA.n2186 GNDA.n394 101.718
R1792 GNDA.t366 GNDA.n75 47.6748
R1793 GNDA.n2008 GNDA.t408 98.8358
R1794 GNDA.t418 GNDA.n513 98.8358
R1795 GNDA.t373 GNDA.n792 92.5685
R1796 GNDA.n2184 GNDA.n2176 91.069
R1797 GNDA.n2184 GNDA.n2183 91.069
R1798 GNDA.n2181 GNDA.n2174 91.069
R1799 GNDA.n2181 GNDA.n2180 91.069
R1800 GNDA.n586 GNDA.n585 91.069
R1801 GNDA.n581 GNDA.n580 91.069
R1802 GNDA.n1785 GNDA.n1782 90.5562
R1803 GNDA.n594 GNDA.n593 90.5562
R1804 GNDA.n657 GNDA.n409 90.5562
R1805 GNDA.n713 GNDA.n696 90.5562
R1806 GNDA.n2199 GNDA.n2198 90.5562
R1807 GNDA.n2141 GNDA.n420 90.5562
R1808 GNDA.n2131 GNDA.n420 90.5562
R1809 GNDA.t151 GNDA.t228 89.5224
R1810 GNDA.n1798 GNDA.n538 87.5377
R1811 GNDA.t275 GNDA.n418 87.5377
R1812 GNDA.n697 GNDA.t366 86.5315
R1813 GNDA.n103 GNDA.n102 84.306
R1814 GNDA.n2159 GNDA.n407 84.306
R1815 GNDA.n709 GNDA.n702 84.306
R1816 GNDA.n540 GNDA.t125 83.513
R1817 GNDA.n2142 GNDA.n2141 83.513
R1818 GNDA.t289 GNDA.t229 83.1688
R1819 GNDA.t152 GNDA.n592 82.5068
R1820 GNDA.n778 GNDA.t236 82.5068
R1821 GNDA.n2200 GNDA.t232 82.5068
R1822 GNDA.n2364 GNDA.n109 80.9821
R1823 GNDA.t330 GNDA.t192 80.5329
R1824 GNDA.t302 GNDA.t498 80.5329
R1825 GNDA.t40 GNDA.t493 80.5329
R1826 GNDA.t39 GNDA.t550 80.5329
R1827 GNDA.t193 GNDA.t335 80.5329
R1828 GNDA.t173 GNDA.t171 80.5329
R1829 GNDA.t171 GNDA.t323 80.5329
R1830 GNDA.t590 GNDA.t262 80.5329
R1831 GNDA.t264 GNDA.t17 80.5329
R1832 GNDA.t313 GNDA.t588 80.5329
R1833 GNDA.t326 GNDA.t220 80.5329
R1834 GNDA.t329 GNDA.t199 80.5329
R1835 GNDA.t587 GNDA.t266 80.5329
R1836 GNDA.n607 GNDA.t15 78.4821
R1837 GNDA.n684 GNDA.t13 78.4821
R1838 GNDA.t578 GNDA.n2188 78.4821
R1839 GNDA.t386 GNDA.t459 76.8724
R1840 GNDA.t380 GNDA.t376 76.8724
R1841 GNDA.n525 GNDA.t140 76.8724
R1842 GNDA.t426 GNDA.t443 76.8724
R1843 GNDA.t437 GNDA.t440 76.8724
R1844 GNDA.n2424 GNDA.n76 76.7001
R1845 GNDA.n2418 GNDA.n76 76.7001
R1846 GNDA.n2418 GNDA.n2417 76.7001
R1847 GNDA.n2417 GNDA.n2416 76.7001
R1848 GNDA.n2416 GNDA.n82 76.7001
R1849 GNDA.n2410 GNDA.n2409 76.7001
R1850 GNDA.n2409 GNDA.n2408 76.7001
R1851 GNDA.n2408 GNDA.n86 76.7001
R1852 GNDA.n2402 GNDA.n86 76.7001
R1853 GNDA.n2402 GNDA.n64 76.7001
R1854 GNDA.n97 GNDA.n63 76.7001
R1855 GNDA.n2388 GNDA.n97 76.7001
R1856 GNDA.n2388 GNDA.n2387 76.7001
R1857 GNDA.n2387 GNDA.n2386 76.7001
R1858 GNDA.n2386 GNDA.n98 76.7001
R1859 GNDA.n2379 GNDA.n104 76.7001
R1860 GNDA.n108 GNDA.n104 76.7001
R1861 GNDA.n2372 GNDA.n108 76.7001
R1862 GNDA.n2372 GNDA.n2371 76.7001
R1863 GNDA.n2371 GNDA.n2370 76.7001
R1864 GNDA.n154 GNDA.n153 76.7001
R1865 GNDA.n159 GNDA.n154 76.7001
R1866 GNDA.n160 GNDA.n159 76.7001
R1867 GNDA.n162 GNDA.n160 76.7001
R1868 GNDA.n162 GNDA.n161 76.7001
R1869 GNDA.n169 GNDA.n168 76.7001
R1870 GNDA.n170 GNDA.n169 76.7001
R1871 GNDA.n170 GNDA.n146 76.7001
R1872 GNDA.n176 GNDA.n146 76.7001
R1873 GNDA.n177 GNDA.n176 76.7001
R1874 GNDA.n2308 GNDA.n2307 76.3222
R1875 GNDA.n619 GNDA.n323 76.3222
R1876 GNDA.n627 GNDA.n322 76.3222
R1877 GNDA.n631 GNDA.n321 76.3222
R1878 GNDA.n638 GNDA.n320 76.3222
R1879 GNDA.n640 GNDA.n319 76.3222
R1880 GNDA.n2253 GNDA.n2252 76.3222
R1881 GNDA.n2254 GNDA.n2250 76.3222
R1882 GNDA.n2261 GNDA.n2260 76.3222
R1883 GNDA.n2262 GNDA.n2248 76.3222
R1884 GNDA.n2269 GNDA.n2268 76.3222
R1885 GNDA.n2273 GNDA.n2246 76.3222
R1886 GNDA.n345 GNDA.n325 76.3222
R1887 GNDA.n2283 GNDA.n326 76.3222
R1888 GNDA.n341 GNDA.n327 76.3222
R1889 GNDA.n2293 GNDA.n328 76.3222
R1890 GNDA.n337 GNDA.n329 76.3222
R1891 GNDA.n2304 GNDA.n2303 76.3222
R1892 GNDA.n2395 GNDA.n2394 76.3222
R1893 GNDA.n1515 GNDA.n92 76.3222
R1894 GNDA.n1518 GNDA.n1517 76.3222
R1895 GNDA.n1527 GNDA.n1526 76.3222
R1896 GNDA.n1530 GNDA.n1529 76.3222
R1897 GNDA.n1539 GNDA.n1538 76.3222
R1898 GNDA.n1654 GNDA.n31 76.3222
R1899 GNDA.n1649 GNDA.n30 76.3222
R1900 GNDA.n1566 GNDA.n29 76.3222
R1901 GNDA.n1572 GNDA.n28 76.3222
R1902 GNDA.n1578 GNDA.n27 76.3222
R1903 GNDA.n1587 GNDA.n26 76.3222
R1904 GNDA.n285 GNDA.n284 76.3222
R1905 GNDA.n288 GNDA.n287 76.3222
R1906 GNDA.n293 GNDA.n292 76.3222
R1907 GNDA.n296 GNDA.n295 76.3222
R1908 GNDA.n301 GNDA.n300 76.3222
R1909 GNDA.n304 GNDA.n303 76.3222
R1910 GNDA.n1502 GNDA.n1501 76.3222
R1911 GNDA.n1499 GNDA.n1459 76.3222
R1912 GNDA.n1495 GNDA.n1494 76.3222
R1913 GNDA.n1488 GNDA.n1466 76.3222
R1914 GNDA.n1487 GNDA.n1486 76.3222
R1915 GNDA.n1475 GNDA.n1474 76.3222
R1916 GNDA.n1457 GNDA.n1456 76.3222
R1917 GNDA.n1452 GNDA.n1433 76.3222
R1918 GNDA.n1450 GNDA.n1449 76.3222
R1919 GNDA.n1445 GNDA.n1436 76.3222
R1920 GNDA.n1443 GNDA.n1442 76.3222
R1921 GNDA.n1438 GNDA.n1437 76.3222
R1922 GNDA.n1260 GNDA.n311 76.3222
R1923 GNDA.n1145 GNDA.n1144 76.3222
R1924 GNDA.n1251 GNDA.n1143 76.3222
R1925 GNDA.n1177 GNDA.n1142 76.3222
R1926 GNDA.n1181 GNDA.n1141 76.3222
R1927 GNDA.n1190 GNDA.n1140 76.3222
R1928 GNDA.n2337 GNDA.n2336 76.3222
R1929 GNDA.n2334 GNDA.n283 76.3222
R1930 GNDA.n2330 GNDA.n2329 76.3222
R1931 GNDA.n2323 GNDA.n290 76.3222
R1932 GNDA.n2322 GNDA.n2321 76.3222
R1933 GNDA.n2315 GNDA.n298 76.3222
R1934 GNDA.n1002 GNDA.n1001 76.3222
R1935 GNDA.n1007 GNDA.n1006 76.3222
R1936 GNDA.n1008 GNDA.n999 76.3222
R1937 GNDA.n1015 GNDA.n1014 76.3222
R1938 GNDA.n1019 GNDA.n997 76.3222
R1939 GNDA.n1022 GNDA.n1021 76.3222
R1940 GNDA.n1139 GNDA.n306 76.3222
R1941 GNDA.n959 GNDA.n958 76.3222
R1942 GNDA.n1130 GNDA.n957 76.3222
R1943 GNDA.n1056 GNDA.n956 76.3222
R1944 GNDA.n1060 GNDA.n955 76.3222
R1945 GNDA.n1069 GNDA.n954 76.3222
R1946 GNDA.n2277 GNDA.n2276 76.3222
R1947 GNDA.n2280 GNDA.n2279 76.3222
R1948 GNDA.n2287 GNDA.n2286 76.3222
R1949 GNDA.n2290 GNDA.n2289 76.3222
R1950 GNDA.n2297 GNDA.n2296 76.3222
R1951 GNDA.n2300 GNDA.n2299 76.3222
R1952 GNDA.n2242 GNDA.n349 76.3222
R1953 GNDA.n2240 GNDA.n2239 76.3222
R1954 GNDA.n2235 GNDA.n352 76.3222
R1955 GNDA.n2233 GNDA.n2232 76.3222
R1956 GNDA.n2228 GNDA.n355 76.3222
R1957 GNDA.n2226 GNDA.n2225 76.3222
R1958 GNDA.n2399 GNDA.n2398 76.3222
R1959 GNDA.n1513 GNDA.n1512 76.3222
R1960 GNDA.n1522 GNDA.n1521 76.3222
R1961 GNDA.n1523 GNDA.n1508 76.3222
R1962 GNDA.n1534 GNDA.n1533 76.3222
R1963 GNDA.n1535 GNDA.n943 76.3222
R1964 GNDA.n1752 GNDA.n53 76.3222
R1965 GNDA.n1747 GNDA.n52 76.3222
R1966 GNDA.n1664 GNDA.n51 76.3222
R1967 GNDA.n1670 GNDA.n50 76.3222
R1968 GNDA.n1676 GNDA.n49 76.3222
R1969 GNDA.n1685 GNDA.n48 76.3222
R1970 GNDA.n1775 GNDA.n77 76.3222
R1971 GNDA.n1770 GNDA.n854 76.3222
R1972 GNDA.n1767 GNDA.n855 76.3222
R1973 GNDA.n1763 GNDA.n856 76.3222
R1974 GNDA.n1759 GNDA.n857 76.3222
R1975 GNDA.n1461 GNDA.n1460 76.3222
R1976 GNDA.n1464 GNDA.n1463 76.3222
R1977 GNDA.n1469 GNDA.n1468 76.3222
R1978 GNDA.n1472 GNDA.n1471 76.3222
R1979 GNDA.n1478 GNDA.n1477 76.3222
R1980 GNDA.n1481 GNDA.n1480 76.3222
R1981 GNDA.n1405 GNDA.n950 76.3222
R1982 GNDA.n1412 GNDA.n1411 76.3222
R1983 GNDA.n1413 GNDA.n948 76.3222
R1984 GNDA.n1420 GNDA.n1419 76.3222
R1985 GNDA.n1421 GNDA.n946 76.3222
R1986 GNDA.n1428 GNDA.n1427 76.3222
R1987 GNDA.n1381 GNDA.n1380 76.3222
R1988 GNDA.n1378 GNDA.n1377 76.3222
R1989 GNDA.n1292 GNDA.n1264 76.3222
R1990 GNDA.n1298 GNDA.n1263 76.3222
R1991 GNDA.n1304 GNDA.n1262 76.3222
R1992 GNDA.n1313 GNDA.n1261 76.3222
R1993 GNDA.n1404 GNDA.n859 76.3222
R1994 GNDA.n1400 GNDA.n860 76.3222
R1995 GNDA.n1396 GNDA.n861 76.3222
R1996 GNDA.n1392 GNDA.n862 76.3222
R1997 GNDA.n1388 GNDA.n863 76.3222
R1998 GNDA.n618 GNDA.n617 76.3222
R1999 GNDA.n623 GNDA.n622 76.3222
R2000 GNDA.n624 GNDA.n615 76.3222
R2001 GNDA.n635 GNDA.n634 76.3222
R2002 GNDA.n643 GNDA.n613 76.3222
R2003 GNDA.n646 GNDA.n645 76.3222
R2004 GNDA.n896 GNDA.n872 76.3222
R2005 GNDA.n894 GNDA.n893 76.3222
R2006 GNDA.n889 GNDA.n875 76.3222
R2007 GNDA.n887 GNDA.n886 76.3222
R2008 GNDA.n882 GNDA.n878 76.3222
R2009 GNDA.n880 GNDA.n879 76.3222
R2010 GNDA.n918 GNDA.n917 76.3222
R2011 GNDA.n913 GNDA.n868 76.3222
R2012 GNDA.n910 GNDA.n867 76.3222
R2013 GNDA.n906 GNDA.n866 76.3222
R2014 GNDA.n902 GNDA.n865 76.3222
R2015 GNDA.n918 GNDA.n869 76.3222
R2016 GNDA.n911 GNDA.n868 76.3222
R2017 GNDA.n907 GNDA.n867 76.3222
R2018 GNDA.n903 GNDA.n866 76.3222
R2019 GNDA.n899 GNDA.n865 76.3222
R2020 GNDA.n1401 GNDA.n859 76.3222
R2021 GNDA.n1397 GNDA.n860 76.3222
R2022 GNDA.n1393 GNDA.n861 76.3222
R2023 GNDA.n1389 GNDA.n862 76.3222
R2024 GNDA.n1385 GNDA.n863 76.3222
R2025 GNDA.n1775 GNDA.n1774 76.3222
R2026 GNDA.n1768 GNDA.n854 76.3222
R2027 GNDA.n1764 GNDA.n855 76.3222
R2028 GNDA.n1760 GNDA.n856 76.3222
R2029 GNDA.n1756 GNDA.n857 76.3222
R2030 GNDA.n2227 GNDA.n2226 76.3222
R2031 GNDA.n355 GNDA.n353 76.3222
R2032 GNDA.n2234 GNDA.n2233 76.3222
R2033 GNDA.n352 GNDA.n350 76.3222
R2034 GNDA.n2241 GNDA.n2240 76.3222
R2035 GNDA.n349 GNDA.n347 76.3222
R2036 GNDA.n1380 GNDA.n953 76.3222
R2037 GNDA.n1378 GNDA.n1265 76.3222
R2038 GNDA.n1297 GNDA.n1264 76.3222
R2039 GNDA.n1305 GNDA.n1263 76.3222
R2040 GNDA.n1312 GNDA.n1262 76.3222
R2041 GNDA.n1287 GNDA.n1261 76.3222
R2042 GNDA.n1260 GNDA.n1259 76.3222
R2043 GNDA.n1252 GNDA.n1144 76.3222
R2044 GNDA.n1176 GNDA.n1143 76.3222
R2045 GNDA.n1182 GNDA.n1142 76.3222
R2046 GNDA.n1189 GNDA.n1141 76.3222
R2047 GNDA.n1171 GNDA.n1140 76.3222
R2048 GNDA.n1139 GNDA.n1138 76.3222
R2049 GNDA.n1131 GNDA.n958 76.3222
R2050 GNDA.n1055 GNDA.n957 76.3222
R2051 GNDA.n1061 GNDA.n956 76.3222
R2052 GNDA.n1068 GNDA.n955 76.3222
R2053 GNDA.n1050 GNDA.n954 76.3222
R2054 GNDA.n1427 GNDA.n1426 76.3222
R2055 GNDA.n1422 GNDA.n1421 76.3222
R2056 GNDA.n1419 GNDA.n1418 76.3222
R2057 GNDA.n1414 GNDA.n1413 76.3222
R2058 GNDA.n1411 GNDA.n1410 76.3222
R2059 GNDA.n1406 GNDA.n1405 76.3222
R2060 GNDA.n1439 GNDA.n1438 76.3222
R2061 GNDA.n1444 GNDA.n1443 76.3222
R2062 GNDA.n1436 GNDA.n1434 76.3222
R2063 GNDA.n1451 GNDA.n1450 76.3222
R2064 GNDA.n1433 GNDA.n1431 76.3222
R2065 GNDA.n1458 GNDA.n1457 76.3222
R2066 GNDA.n1021 GNDA.n1020 76.3222
R2067 GNDA.n1016 GNDA.n997 76.3222
R2068 GNDA.n1014 GNDA.n1013 76.3222
R2069 GNDA.n1009 GNDA.n1008 76.3222
R2070 GNDA.n1006 GNDA.n1005 76.3222
R2071 GNDA.n1001 GNDA.n282 76.3222
R2072 GNDA.n1748 GNDA.n53 76.3222
R2073 GNDA.n1663 GNDA.n52 76.3222
R2074 GNDA.n1669 GNDA.n51 76.3222
R2075 GNDA.n1677 GNDA.n50 76.3222
R2076 GNDA.n1684 GNDA.n49 76.3222
R2077 GNDA.n1658 GNDA.n48 76.3222
R2078 GNDA.n2340 GNDA.n47 76.3222
R2079 GNDA.n2428 GNDA.n2427 76.3222
R2080 GNDA.n46 GNDA.n45 76.3222
R2081 GNDA.n35 GNDA.n34 76.3222
R2082 GNDA.n210 GNDA.n33 76.3222
R2083 GNDA.n216 GNDA.n32 76.3222
R2084 GNDA.n47 GNDA.n24 76.3222
R2085 GNDA.n2427 GNDA.n25 76.3222
R2086 GNDA.n46 GNDA.n36 76.3222
R2087 GNDA.n209 GNDA.n34 76.3222
R2088 GNDA.n215 GNDA.n33 76.3222
R2089 GNDA.n205 GNDA.n32 76.3222
R2090 GNDA.n1650 GNDA.n31 76.3222
R2091 GNDA.n1565 GNDA.n30 76.3222
R2092 GNDA.n1571 GNDA.n29 76.3222
R2093 GNDA.n1579 GNDA.n28 76.3222
R2094 GNDA.n1586 GNDA.n27 76.3222
R2095 GNDA.n276 GNDA.n26 76.3222
R2096 GNDA.n303 GNDA.n302 76.3222
R2097 GNDA.n300 GNDA.n299 76.3222
R2098 GNDA.n295 GNDA.n294 76.3222
R2099 GNDA.n292 GNDA.n291 76.3222
R2100 GNDA.n287 GNDA.n286 76.3222
R2101 GNDA.n284 GNDA.n280 76.3222
R2102 GNDA.n2336 GNDA.n2335 76.3222
R2103 GNDA.n2331 GNDA.n283 76.3222
R2104 GNDA.n2329 GNDA.n2328 76.3222
R2105 GNDA.n2324 GNDA.n2323 76.3222
R2106 GNDA.n2321 GNDA.n2320 76.3222
R2107 GNDA.n2316 GNDA.n2315 76.3222
R2108 GNDA.n2304 GNDA.n330 76.3222
R2109 GNDA.n2294 GNDA.n329 76.3222
R2110 GNDA.n342 GNDA.n328 76.3222
R2111 GNDA.n2284 GNDA.n327 76.3222
R2112 GNDA.n346 GNDA.n326 76.3222
R2113 GNDA.n2274 GNDA.n325 76.3222
R2114 GNDA.n2278 GNDA.n2277 76.3222
R2115 GNDA.n2279 GNDA.n343 76.3222
R2116 GNDA.n2288 GNDA.n2287 76.3222
R2117 GNDA.n2289 GNDA.n339 76.3222
R2118 GNDA.n2298 GNDA.n2297 76.3222
R2119 GNDA.n2301 GNDA.n2300 76.3222
R2120 GNDA.n2270 GNDA.n2246 76.3222
R2121 GNDA.n2268 GNDA.n2267 76.3222
R2122 GNDA.n2263 GNDA.n2262 76.3222
R2123 GNDA.n2260 GNDA.n2259 76.3222
R2124 GNDA.n2255 GNDA.n2254 76.3222
R2125 GNDA.n2252 GNDA.n317 76.3222
R2126 GNDA.n881 GNDA.n880 76.3222
R2127 GNDA.n878 GNDA.n876 76.3222
R2128 GNDA.n888 GNDA.n887 76.3222
R2129 GNDA.n875 GNDA.n873 76.3222
R2130 GNDA.n895 GNDA.n894 76.3222
R2131 GNDA.n872 GNDA.n870 76.3222
R2132 GNDA.n645 GNDA.n644 76.3222
R2133 GNDA.n636 GNDA.n613 76.3222
R2134 GNDA.n634 GNDA.n633 76.3222
R2135 GNDA.n625 GNDA.n624 76.3222
R2136 GNDA.n622 GNDA.n621 76.3222
R2137 GNDA.n617 GNDA.n315 76.3222
R2138 GNDA.n2307 GNDA.n318 76.3222
R2139 GNDA.n626 GNDA.n323 76.3222
R2140 GNDA.n630 GNDA.n322 76.3222
R2141 GNDA.n637 GNDA.n321 76.3222
R2142 GNDA.n641 GNDA.n320 76.3222
R2143 GNDA.n648 GNDA.n319 76.3222
R2144 GNDA.n1480 GNDA.n1479 76.3222
R2145 GNDA.n1477 GNDA.n1476 76.3222
R2146 GNDA.n1471 GNDA.n1470 76.3222
R2147 GNDA.n1468 GNDA.n1467 76.3222
R2148 GNDA.n1463 GNDA.n1462 76.3222
R2149 GNDA.n1460 GNDA.n1429 76.3222
R2150 GNDA.n1501 GNDA.n1500 76.3222
R2151 GNDA.n1496 GNDA.n1459 76.3222
R2152 GNDA.n1494 GNDA.n1493 76.3222
R2153 GNDA.n1489 GNDA.n1488 76.3222
R2154 GNDA.n1486 GNDA.n1485 76.3222
R2155 GNDA.n1474 GNDA.n310 76.3222
R2156 GNDA.n1536 GNDA.n1535 76.3222
R2157 GNDA.n1533 GNDA.n1532 76.3222
R2158 GNDA.n1524 GNDA.n1523 76.3222
R2159 GNDA.n1521 GNDA.n1520 76.3222
R2160 GNDA.n1512 GNDA.n90 76.3222
R2161 GNDA.n2400 GNDA.n2399 76.3222
R2162 GNDA.n2396 GNDA.n2395 76.3222
R2163 GNDA.n1516 GNDA.n1515 76.3222
R2164 GNDA.n1517 GNDA.n1510 76.3222
R2165 GNDA.n1528 GNDA.n1527 76.3222
R2166 GNDA.n1529 GNDA.n1506 76.3222
R2167 GNDA.n1540 GNDA.n1539 76.3222
R2168 GNDA.t10 GNDA.n2052 75.8626
R2169 GNDA.n2036 GNDA.t208 75.8626
R2170 GNDA.n1610 GNDA.n1551 74.5978
R2171 GNDA.n1607 GNDA.n1551 74.5978
R2172 GNDA.n239 GNDA.n9 74.5978
R2173 GNDA.n236 GNDA.n9 74.5978
R2174 GNDA.n1213 GNDA.n1159 74.5978
R2175 GNDA.n1210 GNDA.n1159 74.5978
R2176 GNDA.n737 GNDA.n666 74.5978
R2177 GNDA.n734 GNDA.n666 74.5978
R2178 GNDA.n1092 GNDA.n973 74.5978
R2179 GNDA.n1089 GNDA.n973 74.5978
R2180 GNDA.n467 GNDA.n375 74.5978
R2181 GNDA.n470 GNDA.n375 74.5978
R2182 GNDA.n1708 GNDA.n931 74.5978
R2183 GNDA.n1705 GNDA.n931 74.5978
R2184 GNDA.n1336 GNDA.n1275 74.5978
R2185 GNDA.n1333 GNDA.n1275 74.5978
R2186 GNDA.n815 GNDA.n814 74.5978
R2187 GNDA.n814 GNDA.n813 74.5978
R2188 GNDA.n794 GNDA.t64 72.445
R2189 GNDA.t1 GNDA.t589 71.618
R2190 GNDA.n2124 GNDA.t0 69.38
R2191 GNDA.n1644 GNDA.n1544 69.3109
R2192 GNDA.n1644 GNDA.n1643 69.3109
R2193 GNDA.n2432 GNDA.n2431 69.3109
R2194 GNDA.n2432 GNDA.n20 69.3109
R2195 GNDA.n1256 GNDA.n1149 69.3109
R2196 GNDA.n1232 GNDA.n1149 69.3109
R2197 GNDA.n784 GNDA.n652 69.3109
R2198 GNDA.n755 GNDA.n652 69.3109
R2199 GNDA.n1135 GNDA.n963 69.3109
R2200 GNDA.n1111 GNDA.n963 69.3109
R2201 GNDA.n2205 GNDA.n2204 69.3109
R2202 GNDA.n2205 GNDA.n386 69.3109
R2203 GNDA.n1742 GNDA.n924 69.3109
R2204 GNDA.n1742 GNDA.n1741 69.3109
R2205 GNDA.n1372 GNDA.n1268 69.3109
R2206 GNDA.n1372 GNDA.n1371 69.3109
R2207 GNDA.n1790 GNDA.n545 69.3109
R2208 GNDA.n848 GNDA.n545 69.3109
R2209 GNDA.n430 GNDA.t194 68.4204
R2210 GNDA.t368 GNDA.n1561 65.8183
R2211 GNDA.t368 GNDA.n1560 65.8183
R2212 GNDA.t368 GNDA.n1559 65.8183
R2213 GNDA.t368 GNDA.n1558 65.8183
R2214 GNDA.t368 GNDA.n1549 65.8183
R2215 GNDA.t368 GNDA.n1556 65.8183
R2216 GNDA.t368 GNDA.n1546 65.8183
R2217 GNDA.t368 GNDA.n1557 65.8183
R2218 GNDA.t368 GNDA.n1555 65.8183
R2219 GNDA.t368 GNDA.n1554 65.8183
R2220 GNDA.t368 GNDA.n1553 65.8183
R2221 GNDA.t368 GNDA.n1552 65.8183
R2222 GNDA.t398 GNDA.n19 65.8183
R2223 GNDA.t398 GNDA.n18 65.8183
R2224 GNDA.t398 GNDA.n17 65.8183
R2225 GNDA.t398 GNDA.n16 65.8183
R2226 GNDA.t398 GNDA.n7 65.8183
R2227 GNDA.t398 GNDA.n14 65.8183
R2228 GNDA.t398 GNDA.n5 65.8183
R2229 GNDA.t398 GNDA.n15 65.8183
R2230 GNDA.t398 GNDA.n13 65.8183
R2231 GNDA.t398 GNDA.n12 65.8183
R2232 GNDA.t398 GNDA.n11 65.8183
R2233 GNDA.t398 GNDA.n10 65.8183
R2234 GNDA.t378 GNDA.n1246 65.8183
R2235 GNDA.t378 GNDA.n1168 65.8183
R2236 GNDA.t378 GNDA.n1167 65.8183
R2237 GNDA.t378 GNDA.n1166 65.8183
R2238 GNDA.t378 GNDA.n1157 65.8183
R2239 GNDA.t378 GNDA.n1164 65.8183
R2240 GNDA.t378 GNDA.n1155 65.8183
R2241 GNDA.t378 GNDA.n1165 65.8183
R2242 GNDA.t378 GNDA.n1163 65.8183
R2243 GNDA.t378 GNDA.n1162 65.8183
R2244 GNDA.t378 GNDA.n1161 65.8183
R2245 GNDA.t378 GNDA.n1160 65.8183
R2246 GNDA.t378 GNDA.n1158 65.8183
R2247 GNDA.t378 GNDA.n1156 65.8183
R2248 GNDA.n1247 GNDA.t378 65.8183
R2249 GNDA.t378 GNDA.n1150 65.8183
R2250 GNDA.t397 GNDA.n769 65.8183
R2251 GNDA.t397 GNDA.n675 65.8183
R2252 GNDA.t397 GNDA.n674 65.8183
R2253 GNDA.t397 GNDA.n673 65.8183
R2254 GNDA.t397 GNDA.n664 65.8183
R2255 GNDA.t397 GNDA.n671 65.8183
R2256 GNDA.t397 GNDA.n662 65.8183
R2257 GNDA.t397 GNDA.n672 65.8183
R2258 GNDA.t397 GNDA.n670 65.8183
R2259 GNDA.t397 GNDA.n669 65.8183
R2260 GNDA.t397 GNDA.n668 65.8183
R2261 GNDA.t397 GNDA.n667 65.8183
R2262 GNDA.t397 GNDA.n665 65.8183
R2263 GNDA.t397 GNDA.n663 65.8183
R2264 GNDA.n772 GNDA.t397 65.8183
R2265 GNDA.t397 GNDA.n653 65.8183
R2266 GNDA.t396 GNDA.n1125 65.8183
R2267 GNDA.t396 GNDA.n982 65.8183
R2268 GNDA.t396 GNDA.n981 65.8183
R2269 GNDA.t396 GNDA.n980 65.8183
R2270 GNDA.t396 GNDA.n971 65.8183
R2271 GNDA.t396 GNDA.n978 65.8183
R2272 GNDA.t396 GNDA.n969 65.8183
R2273 GNDA.t396 GNDA.n979 65.8183
R2274 GNDA.t396 GNDA.n977 65.8183
R2275 GNDA.t396 GNDA.n976 65.8183
R2276 GNDA.t396 GNDA.n975 65.8183
R2277 GNDA.t396 GNDA.n974 65.8183
R2278 GNDA.t396 GNDA.n972 65.8183
R2279 GNDA.t396 GNDA.n970 65.8183
R2280 GNDA.n1126 GNDA.t396 65.8183
R2281 GNDA.t396 GNDA.n964 65.8183
R2282 GNDA.t432 GNDA.n385 65.8183
R2283 GNDA.t432 GNDA.n384 65.8183
R2284 GNDA.t432 GNDA.n383 65.8183
R2285 GNDA.t432 GNDA.n382 65.8183
R2286 GNDA.t432 GNDA.n373 65.8183
R2287 GNDA.t432 GNDA.n380 65.8183
R2288 GNDA.t432 GNDA.n371 65.8183
R2289 GNDA.t432 GNDA.n381 65.8183
R2290 GNDA.t432 GNDA.n379 65.8183
R2291 GNDA.t432 GNDA.n378 65.8183
R2292 GNDA.t432 GNDA.n377 65.8183
R2293 GNDA.t432 GNDA.n376 65.8183
R2294 GNDA.t432 GNDA.n374 65.8183
R2295 GNDA.n2206 GNDA.t432 65.8183
R2296 GNDA.t432 GNDA.n372 65.8183
R2297 GNDA.t432 GNDA.n370 65.8183
R2298 GNDA.t420 GNDA.n941 65.8183
R2299 GNDA.t420 GNDA.n940 65.8183
R2300 GNDA.t420 GNDA.n939 65.8183
R2301 GNDA.t420 GNDA.n938 65.8183
R2302 GNDA.t420 GNDA.n929 65.8183
R2303 GNDA.t420 GNDA.n936 65.8183
R2304 GNDA.t420 GNDA.n926 65.8183
R2305 GNDA.t420 GNDA.n937 65.8183
R2306 GNDA.t420 GNDA.n935 65.8183
R2307 GNDA.t420 GNDA.n934 65.8183
R2308 GNDA.t420 GNDA.n933 65.8183
R2309 GNDA.t420 GNDA.n932 65.8183
R2310 GNDA.t420 GNDA.n930 65.8183
R2311 GNDA.t420 GNDA.n928 65.8183
R2312 GNDA.t420 GNDA.n927 65.8183
R2313 GNDA.n1743 GNDA.t420 65.8183
R2314 GNDA.t367 GNDA.n1285 65.8183
R2315 GNDA.t367 GNDA.n1284 65.8183
R2316 GNDA.t367 GNDA.n1283 65.8183
R2317 GNDA.t367 GNDA.n1282 65.8183
R2318 GNDA.t367 GNDA.n1273 65.8183
R2319 GNDA.t367 GNDA.n1280 65.8183
R2320 GNDA.t367 GNDA.n1270 65.8183
R2321 GNDA.t367 GNDA.n1281 65.8183
R2322 GNDA.t367 GNDA.n1279 65.8183
R2323 GNDA.t367 GNDA.n1278 65.8183
R2324 GNDA.t367 GNDA.n1277 65.8183
R2325 GNDA.t367 GNDA.n1276 65.8183
R2326 GNDA.t367 GNDA.n1274 65.8183
R2327 GNDA.t367 GNDA.n1272 65.8183
R2328 GNDA.t367 GNDA.n1271 65.8183
R2329 GNDA.n1373 GNDA.t367 65.8183
R2330 GNDA.n832 GNDA.t365 65.8183
R2331 GNDA.n838 GNDA.t365 65.8183
R2332 GNDA.n840 GNDA.t365 65.8183
R2333 GNDA.n846 GNDA.t365 65.8183
R2334 GNDA.n816 GNDA.t365 65.8183
R2335 GNDA.n822 GNDA.t365 65.8183
R2336 GNDA.n824 GNDA.t365 65.8183
R2337 GNDA.n830 GNDA.t365 65.8183
R2338 GNDA.n800 GNDA.t365 65.8183
R2339 GNDA.n560 GNDA.t365 65.8183
R2340 GNDA.n807 GNDA.t365 65.8183
R2341 GNDA.n557 GNDA.t365 65.8183
R2342 GNDA.n601 GNDA.t365 65.8183
R2343 GNDA.n599 GNDA.t365 65.8183
R2344 GNDA.n569 GNDA.t365 65.8183
R2345 GNDA.n1792 GNDA.t365 65.8183
R2346 GNDA.t398 GNDA.n8 65.8183
R2347 GNDA.n2433 GNDA.t398 65.8183
R2348 GNDA.t398 GNDA.n6 65.8183
R2349 GNDA.t398 GNDA.n4 65.8183
R2350 GNDA.t368 GNDA.n1550 65.8183
R2351 GNDA.t368 GNDA.n1548 65.8183
R2352 GNDA.t368 GNDA.n1547 65.8183
R2353 GNDA.n1645 GNDA.t368 65.8183
R2354 GNDA.t408 GNDA.t7 64.8799
R2355 GNDA.t7 GNDA.t222 64.8799
R2356 GNDA.t222 GNDA.t178 64.8799
R2357 GNDA.t9 GNDA.t303 64.8799
R2358 GNDA.t303 GNDA.t418 64.8799
R2359 GNDA.n2130 GNDA.n505 63.891
R2360 GNDA.n779 GNDA.t216 62.3833
R2361 GNDA.n429 GNDA.t154 62.3833
R2362 GNDA.n524 GNDA.t447 62.2505
R2363 GNDA.n2091 GNDA.t390 62.2505
R2364 GNDA.n2009 GNDA.t416 62.2505
R2365 GNDA.n2013 GNDA.t422 62.2505
R2366 GNDA.n2012 GNDA.t400 62.2505
R2367 GNDA.n2024 GNDA.t411 62.2505
R2368 GNDA.n526 GNDA.t392 62.2505
R2369 GNDA.n2018 GNDA.t424 62.2505
R2370 GNDA.n2007 GNDA.t409 62.2505
R2371 GNDA.n2032 GNDA.t395 62.2505
R2372 GNDA.n2027 GNDA.t403 62.2505
R2373 GNDA.n521 GNDA.t419 62.2505
R2374 GNDA.t28 GNDA.t330 62.2301
R2375 GNDA.t335 GNDA.t336 62.2301
R2376 GNDA.n2026 GNDA.t276 62.2301
R2377 GNDA.t17 GNDA.t290 62.2301
R2378 GNDA.t321 GNDA.t587 62.2301
R2379 GNDA.n1982 GNDA.n1981 59.2425
R2380 GNDA.n2116 GNDA.n2115 59.2425
R2381 GNDA.n2106 GNDA.n511 59.2425
R2382 GNDA.n1992 GNDA.n1991 59.2425
R2383 GNDA.n2130 GNDA.t97 58.6335
R2384 GNDA.n608 GNDA.t196 58.3586
R2385 GNDA.n695 GNDA.t585 58.3586
R2386 GNDA.t378 GNDA.n1149 57.8461
R2387 GNDA.t397 GNDA.n652 57.8461
R2388 GNDA.t396 GNDA.n963 57.8461
R2389 GNDA.t432 GNDA.n2205 57.8461
R2390 GNDA.t420 GNDA.n1742 57.8461
R2391 GNDA.t367 GNDA.n1372 57.8461
R2392 GNDA.n545 GNDA.t365 57.8461
R2393 GNDA.t398 GNDA.n2432 57.8461
R2394 GNDA.t368 GNDA.n1644 57.8461
R2395 GNDA.n2158 GNDA.n408 57.3524
R2396 GNDA.n700 GNDA.n699 57.3524
R2397 GNDA.n1048 GNDA.n1047 56.3995
R2398 GNDA.n500 GNDA.n499 56.3995
R2399 GNDA.n499 GNDA.n486 56.3995
R2400 GNDA.n1049 GNDA.n1048 56.3995
R2401 GNDA.n1755 GNDA.n858 56.3995
R2402 GNDA.n951 GNDA.n919 56.3995
R2403 GNDA.n1778 GNDA.n1777 56.3995
R2404 GNDA.n1777 GNDA.n851 56.3995
R2405 GNDA.n1382 GNDA.n919 56.3995
R2406 GNDA.n1753 GNDA.n858 56.3995
R2407 GNDA.n201 GNDA.n135 56.3995
R2408 GNDA.n204 GNDA.n135 56.3995
R2409 GNDA.n994 GNDA.t165 56.1801
R2410 GNDA.t368 GNDA.n1551 55.2026
R2411 GNDA.t398 GNDA.n9 55.2026
R2412 GNDA.t378 GNDA.n1159 55.2026
R2413 GNDA.t397 GNDA.n666 55.2026
R2414 GNDA.t396 GNDA.n973 55.2026
R2415 GNDA.t432 GNDA.n375 55.2026
R2416 GNDA.t420 GNDA.n931 55.2026
R2417 GNDA.t367 GNDA.n1275 55.2026
R2418 GNDA.n814 GNDA.t365 55.2026
R2419 GNDA.n1992 GNDA.t459 54.909
R2420 GNDA.n1981 GNDA.t380 54.909
R2421 GNDA.n2116 GNDA.t426 54.909
R2422 GNDA.t440 GNDA.n511 54.909
R2423 GNDA.t0 GNDA.t1 53.7136
R2424 GNDA.t42 GNDA.t44 53.7136
R2425 GNDA.t44 GNDA.t288 53.7136
R2426 GNDA.t47 GNDA.t200 53.7136
R2427 GNDA.t200 GNDA.t230 53.7136
R2428 GNDA.t228 GNDA.t274 53.7136
R2429 GNDA.n1626 GNDA.n1557 53.3664
R2430 GNDA.n1622 GNDA.n1546 53.3664
R2431 GNDA.n1618 GNDA.n1556 53.3664
R2432 GNDA.n1614 GNDA.n1549 53.3664
R2433 GNDA.n1603 GNDA.n1552 53.3664
R2434 GNDA.n1599 GNDA.n1553 53.3664
R2435 GNDA.n1595 GNDA.n1554 53.3664
R2436 GNDA.n1591 GNDA.n1555 53.3664
R2437 GNDA.n1646 GNDA.n1645 53.3664
R2438 GNDA.n1568 GNDA.n1547 53.3664
R2439 GNDA.n1576 GNDA.n1548 53.3664
R2440 GNDA.n1583 GNDA.n1550 53.3664
R2441 GNDA.n1630 GNDA.n1561 53.3664
R2442 GNDA.n1631 GNDA.n1560 53.3664
R2443 GNDA.n1635 GNDA.n1559 53.3664
R2444 GNDA.n1639 GNDA.n1558 53.3664
R2445 GNDA.n1627 GNDA.n1561 53.3664
R2446 GNDA.n1634 GNDA.n1560 53.3664
R2447 GNDA.n1638 GNDA.n1559 53.3664
R2448 GNDA.n1642 GNDA.n1558 53.3664
R2449 GNDA.n1611 GNDA.n1549 53.3664
R2450 GNDA.n1615 GNDA.n1556 53.3664
R2451 GNDA.n1619 GNDA.n1546 53.3664
R2452 GNDA.n1623 GNDA.n1557 53.3664
R2453 GNDA.n1594 GNDA.n1555 53.3664
R2454 GNDA.n1598 GNDA.n1554 53.3664
R2455 GNDA.n1602 GNDA.n1553 53.3664
R2456 GNDA.n1606 GNDA.n1552 53.3664
R2457 GNDA.n255 GNDA.n15 53.3664
R2458 GNDA.n251 GNDA.n5 53.3664
R2459 GNDA.n247 GNDA.n14 53.3664
R2460 GNDA.n243 GNDA.n7 53.3664
R2461 GNDA.n232 GNDA.n10 53.3664
R2462 GNDA.n228 GNDA.n11 53.3664
R2463 GNDA.n224 GNDA.n12 53.3664
R2464 GNDA.n220 GNDA.n13 53.3664
R2465 GNDA.n21 GNDA.n4 53.3664
R2466 GNDA.n42 GNDA.n6 53.3664
R2467 GNDA.n2434 GNDA.n2433 53.3664
R2468 GNDA.n212 GNDA.n8 53.3664
R2469 GNDA.n259 GNDA.n19 53.3664
R2470 GNDA.n260 GNDA.n18 53.3664
R2471 GNDA.n264 GNDA.n17 53.3664
R2472 GNDA.n268 GNDA.n16 53.3664
R2473 GNDA.n256 GNDA.n19 53.3664
R2474 GNDA.n263 GNDA.n18 53.3664
R2475 GNDA.n267 GNDA.n17 53.3664
R2476 GNDA.n270 GNDA.n16 53.3664
R2477 GNDA.n240 GNDA.n7 53.3664
R2478 GNDA.n244 GNDA.n14 53.3664
R2479 GNDA.n248 GNDA.n5 53.3664
R2480 GNDA.n252 GNDA.n15 53.3664
R2481 GNDA.n223 GNDA.n13 53.3664
R2482 GNDA.n227 GNDA.n12 53.3664
R2483 GNDA.n231 GNDA.n11 53.3664
R2484 GNDA.n235 GNDA.n10 53.3664
R2485 GNDA.n1228 GNDA.n1165 53.3664
R2486 GNDA.n1225 GNDA.n1155 53.3664
R2487 GNDA.n1221 GNDA.n1164 53.3664
R2488 GNDA.n1217 GNDA.n1157 53.3664
R2489 GNDA.n1206 GNDA.n1160 53.3664
R2490 GNDA.n1202 GNDA.n1161 53.3664
R2491 GNDA.n1198 GNDA.n1162 53.3664
R2492 GNDA.n1194 GNDA.n1163 53.3664
R2493 GNDA.n1255 GNDA.n1150 53.3664
R2494 GNDA.n1248 GNDA.n1247 53.3664
R2495 GNDA.n1179 GNDA.n1156 53.3664
R2496 GNDA.n1186 GNDA.n1158 53.3664
R2497 GNDA.n1246 GNDA.n1245 53.3664
R2498 GNDA.n1170 GNDA.n1168 53.3664
R2499 GNDA.n1240 GNDA.n1167 53.3664
R2500 GNDA.n1236 GNDA.n1166 53.3664
R2501 GNDA.n1246 GNDA.n1169 53.3664
R2502 GNDA.n1241 GNDA.n1168 53.3664
R2503 GNDA.n1237 GNDA.n1167 53.3664
R2504 GNDA.n1233 GNDA.n1166 53.3664
R2505 GNDA.n1214 GNDA.n1157 53.3664
R2506 GNDA.n1218 GNDA.n1164 53.3664
R2507 GNDA.n1222 GNDA.n1155 53.3664
R2508 GNDA.n1226 GNDA.n1165 53.3664
R2509 GNDA.n1197 GNDA.n1163 53.3664
R2510 GNDA.n1201 GNDA.n1162 53.3664
R2511 GNDA.n1205 GNDA.n1161 53.3664
R2512 GNDA.n1209 GNDA.n1160 53.3664
R2513 GNDA.n1193 GNDA.n1158 53.3664
R2514 GNDA.n1185 GNDA.n1156 53.3664
R2515 GNDA.n1247 GNDA.n1154 53.3664
R2516 GNDA.n1153 GNDA.n1150 53.3664
R2517 GNDA.n752 GNDA.n672 53.3664
R2518 GNDA.n749 GNDA.n662 53.3664
R2519 GNDA.n745 GNDA.n671 53.3664
R2520 GNDA.n741 GNDA.n664 53.3664
R2521 GNDA.n730 GNDA.n667 53.3664
R2522 GNDA.n726 GNDA.n668 53.3664
R2523 GNDA.n722 GNDA.n669 53.3664
R2524 GNDA.n718 GNDA.n670 53.3664
R2525 GNDA.n783 GNDA.n653 53.3664
R2526 GNDA.n772 GNDA.n771 53.3664
R2527 GNDA.n663 GNDA.n661 53.3664
R2528 GNDA.n691 GNDA.n665 53.3664
R2529 GNDA.n769 GNDA.n768 53.3664
R2530 GNDA.n677 GNDA.n675 53.3664
R2531 GNDA.n763 GNDA.n674 53.3664
R2532 GNDA.n759 GNDA.n673 53.3664
R2533 GNDA.n769 GNDA.n676 53.3664
R2534 GNDA.n764 GNDA.n675 53.3664
R2535 GNDA.n760 GNDA.n674 53.3664
R2536 GNDA.n756 GNDA.n673 53.3664
R2537 GNDA.n738 GNDA.n664 53.3664
R2538 GNDA.n742 GNDA.n671 53.3664
R2539 GNDA.n746 GNDA.n662 53.3664
R2540 GNDA.n750 GNDA.n672 53.3664
R2541 GNDA.n721 GNDA.n670 53.3664
R2542 GNDA.n725 GNDA.n669 53.3664
R2543 GNDA.n729 GNDA.n668 53.3664
R2544 GNDA.n733 GNDA.n667 53.3664
R2545 GNDA.n717 GNDA.n665 53.3664
R2546 GNDA.n690 GNDA.n663 53.3664
R2547 GNDA.n773 GNDA.n772 53.3664
R2548 GNDA.n770 GNDA.n653 53.3664
R2549 GNDA.n1107 GNDA.n979 53.3664
R2550 GNDA.n1104 GNDA.n969 53.3664
R2551 GNDA.n1100 GNDA.n978 53.3664
R2552 GNDA.n1096 GNDA.n971 53.3664
R2553 GNDA.n1085 GNDA.n974 53.3664
R2554 GNDA.n1081 GNDA.n975 53.3664
R2555 GNDA.n1077 GNDA.n976 53.3664
R2556 GNDA.n1073 GNDA.n977 53.3664
R2557 GNDA.n1134 GNDA.n964 53.3664
R2558 GNDA.n1127 GNDA.n1126 53.3664
R2559 GNDA.n1058 GNDA.n970 53.3664
R2560 GNDA.n1065 GNDA.n972 53.3664
R2561 GNDA.n1125 GNDA.n1124 53.3664
R2562 GNDA.n984 GNDA.n982 53.3664
R2563 GNDA.n1119 GNDA.n981 53.3664
R2564 GNDA.n1115 GNDA.n980 53.3664
R2565 GNDA.n1125 GNDA.n983 53.3664
R2566 GNDA.n1120 GNDA.n982 53.3664
R2567 GNDA.n1116 GNDA.n981 53.3664
R2568 GNDA.n1112 GNDA.n980 53.3664
R2569 GNDA.n1093 GNDA.n971 53.3664
R2570 GNDA.n1097 GNDA.n978 53.3664
R2571 GNDA.n1101 GNDA.n969 53.3664
R2572 GNDA.n1105 GNDA.n979 53.3664
R2573 GNDA.n1076 GNDA.n977 53.3664
R2574 GNDA.n1080 GNDA.n976 53.3664
R2575 GNDA.n1084 GNDA.n975 53.3664
R2576 GNDA.n1088 GNDA.n974 53.3664
R2577 GNDA.n1072 GNDA.n972 53.3664
R2578 GNDA.n1064 GNDA.n970 53.3664
R2579 GNDA.n1126 GNDA.n968 53.3664
R2580 GNDA.n967 GNDA.n964 53.3664
R2581 GNDA.n451 GNDA.n381 53.3664
R2582 GNDA.n455 GNDA.n371 53.3664
R2583 GNDA.n459 GNDA.n380 53.3664
R2584 GNDA.n463 GNDA.n373 53.3664
R2585 GNDA.n474 GNDA.n376 53.3664
R2586 GNDA.n478 GNDA.n377 53.3664
R2587 GNDA.n482 GNDA.n378 53.3664
R2588 GNDA.n2136 GNDA.n379 53.3664
R2589 GNDA.n387 GNDA.n370 53.3664
R2590 GNDA.n2194 GNDA.n372 53.3664
R2591 GNDA.n2207 GNDA.n2206 53.3664
R2592 GNDA.n425 GNDA.n374 53.3664
R2593 GNDA.n447 GNDA.n385 53.3664
R2594 GNDA.n446 GNDA.n384 53.3664
R2595 GNDA.n442 GNDA.n383 53.3664
R2596 GNDA.n438 GNDA.n382 53.3664
R2597 GNDA.n450 GNDA.n385 53.3664
R2598 GNDA.n443 GNDA.n384 53.3664
R2599 GNDA.n439 GNDA.n383 53.3664
R2600 GNDA.n435 GNDA.n382 53.3664
R2601 GNDA.n466 GNDA.n373 53.3664
R2602 GNDA.n462 GNDA.n380 53.3664
R2603 GNDA.n458 GNDA.n371 53.3664
R2604 GNDA.n454 GNDA.n381 53.3664
R2605 GNDA.n483 GNDA.n379 53.3664
R2606 GNDA.n479 GNDA.n378 53.3664
R2607 GNDA.n475 GNDA.n377 53.3664
R2608 GNDA.n471 GNDA.n376 53.3664
R2609 GNDA.n2137 GNDA.n374 53.3664
R2610 GNDA.n2206 GNDA.n369 53.3664
R2611 GNDA.n372 GNDA.n368 53.3664
R2612 GNDA.n2193 GNDA.n370 53.3664
R2613 GNDA.n1724 GNDA.n937 53.3664
R2614 GNDA.n1720 GNDA.n926 53.3664
R2615 GNDA.n1716 GNDA.n936 53.3664
R2616 GNDA.n1712 GNDA.n929 53.3664
R2617 GNDA.n1701 GNDA.n932 53.3664
R2618 GNDA.n1697 GNDA.n933 53.3664
R2619 GNDA.n1693 GNDA.n934 53.3664
R2620 GNDA.n1689 GNDA.n935 53.3664
R2621 GNDA.n1744 GNDA.n1743 53.3664
R2622 GNDA.n1666 GNDA.n927 53.3664
R2623 GNDA.n1674 GNDA.n928 53.3664
R2624 GNDA.n1681 GNDA.n930 53.3664
R2625 GNDA.n1728 GNDA.n941 53.3664
R2626 GNDA.n1729 GNDA.n940 53.3664
R2627 GNDA.n1733 GNDA.n939 53.3664
R2628 GNDA.n1737 GNDA.n938 53.3664
R2629 GNDA.n1725 GNDA.n941 53.3664
R2630 GNDA.n1732 GNDA.n940 53.3664
R2631 GNDA.n1736 GNDA.n939 53.3664
R2632 GNDA.n1740 GNDA.n938 53.3664
R2633 GNDA.n1709 GNDA.n929 53.3664
R2634 GNDA.n1713 GNDA.n936 53.3664
R2635 GNDA.n1717 GNDA.n926 53.3664
R2636 GNDA.n1721 GNDA.n937 53.3664
R2637 GNDA.n1692 GNDA.n935 53.3664
R2638 GNDA.n1696 GNDA.n934 53.3664
R2639 GNDA.n1700 GNDA.n933 53.3664
R2640 GNDA.n1704 GNDA.n932 53.3664
R2641 GNDA.n1688 GNDA.n930 53.3664
R2642 GNDA.n1680 GNDA.n928 53.3664
R2643 GNDA.n1673 GNDA.n927 53.3664
R2644 GNDA.n1743 GNDA.n925 53.3664
R2645 GNDA.n1352 GNDA.n1281 53.3664
R2646 GNDA.n1348 GNDA.n1270 53.3664
R2647 GNDA.n1344 GNDA.n1280 53.3664
R2648 GNDA.n1340 GNDA.n1273 53.3664
R2649 GNDA.n1329 GNDA.n1276 53.3664
R2650 GNDA.n1325 GNDA.n1277 53.3664
R2651 GNDA.n1321 GNDA.n1278 53.3664
R2652 GNDA.n1317 GNDA.n1279 53.3664
R2653 GNDA.n1374 GNDA.n1373 53.3664
R2654 GNDA.n1294 GNDA.n1271 53.3664
R2655 GNDA.n1302 GNDA.n1272 53.3664
R2656 GNDA.n1309 GNDA.n1274 53.3664
R2657 GNDA.n1356 GNDA.n1285 53.3664
R2658 GNDA.n1357 GNDA.n1284 53.3664
R2659 GNDA.n1361 GNDA.n1283 53.3664
R2660 GNDA.n1365 GNDA.n1282 53.3664
R2661 GNDA.n1353 GNDA.n1285 53.3664
R2662 GNDA.n1360 GNDA.n1284 53.3664
R2663 GNDA.n1364 GNDA.n1283 53.3664
R2664 GNDA.n1286 GNDA.n1282 53.3664
R2665 GNDA.n1337 GNDA.n1273 53.3664
R2666 GNDA.n1341 GNDA.n1280 53.3664
R2667 GNDA.n1345 GNDA.n1270 53.3664
R2668 GNDA.n1349 GNDA.n1281 53.3664
R2669 GNDA.n1320 GNDA.n1279 53.3664
R2670 GNDA.n1324 GNDA.n1278 53.3664
R2671 GNDA.n1328 GNDA.n1277 53.3664
R2672 GNDA.n1332 GNDA.n1276 53.3664
R2673 GNDA.n1316 GNDA.n1274 53.3664
R2674 GNDA.n1308 GNDA.n1272 53.3664
R2675 GNDA.n1301 GNDA.n1271 53.3664
R2676 GNDA.n1373 GNDA.n1269 53.3664
R2677 GNDA.n831 GNDA.n830 53.3664
R2678 GNDA.n824 GNDA.n551 53.3664
R2679 GNDA.n823 GNDA.n822 53.3664
R2680 GNDA.n816 GNDA.n553 53.3664
R2681 GNDA.n809 GNDA.n557 53.3664
R2682 GNDA.n807 GNDA.n806 53.3664
R2683 GNDA.n802 GNDA.n560 53.3664
R2684 GNDA.n800 GNDA.n799 53.3664
R2685 GNDA.n1792 GNDA.n1791 53.3664
R2686 GNDA.n569 GNDA.n544 53.3664
R2687 GNDA.n599 GNDA.n598 53.3664
R2688 GNDA.n602 GNDA.n601 53.3664
R2689 GNDA.n832 GNDA.n549 53.3664
R2690 GNDA.n838 GNDA.n837 53.3664
R2691 GNDA.n841 GNDA.n840 53.3664
R2692 GNDA.n846 GNDA.n845 53.3664
R2693 GNDA.n833 GNDA.n832 53.3664
R2694 GNDA.n839 GNDA.n838 53.3664
R2695 GNDA.n840 GNDA.n547 53.3664
R2696 GNDA.n847 GNDA.n846 53.3664
R2697 GNDA.n817 GNDA.n816 53.3664
R2698 GNDA.n822 GNDA.n821 53.3664
R2699 GNDA.n825 GNDA.n824 53.3664
R2700 GNDA.n830 GNDA.n829 53.3664
R2701 GNDA.n801 GNDA.n800 53.3664
R2702 GNDA.n560 GNDA.n558 53.3664
R2703 GNDA.n808 GNDA.n807 53.3664
R2704 GNDA.n557 GNDA.n555 53.3664
R2705 GNDA.n601 GNDA.n561 53.3664
R2706 GNDA.n600 GNDA.n599 53.3664
R2707 GNDA.n570 GNDA.n569 53.3664
R2708 GNDA.n1793 GNDA.n1792 53.3664
R2709 GNDA.n219 GNDA.n8 53.3664
R2710 GNDA.n2433 GNDA.n3 53.3664
R2711 GNDA.n6 GNDA.n2 53.3664
R2712 GNDA.n41 GNDA.n4 53.3664
R2713 GNDA.n1590 GNDA.n1550 53.3664
R2714 GNDA.n1582 GNDA.n1548 53.3664
R2715 GNDA.n1575 GNDA.n1547 53.3664
R2716 GNDA.n1645 GNDA.n1545 53.3664
R2717 GNDA.n1784 GNDA.n538 53.3277
R2718 GNDA.n611 GNDA.n408 53.3277
R2719 GNDA.n710 GNDA.n700 53.3277
R2720 GNDA.t260 GNDA.n608 52.3216
R2721 GNDA.t462 GNDA.n695 52.3216
R2722 GNDA.n2211 GNDA.t449 52.3216
R2723 GNDA.n2057 GNDA.t244 50.135
R2724 GNDA.t162 GNDA.n2086 50.135
R2725 GNDA.t452 GNDA.n73 48.2969
R2726 GNDA.n779 GNDA.t413 48.2969
R2727 GNDA.t258 GNDA.n429 48.2969
R2728 GNDA.n2047 GNDA.t12 48.0005
R2729 GNDA.n2047 GNDA.t325 48.0005
R2730 GNDA.n2045 GNDA.t119 48.0005
R2731 GNDA.n2045 GNDA.t53 48.0005
R2732 GNDA.n2043 GNDA.t27 48.0005
R2733 GNDA.n2043 GNDA.t211 48.0005
R2734 GNDA.n2041 GNDA.t78 48.0005
R2735 GNDA.n2041 GNDA.t316 48.0005
R2736 GNDA.n2039 GNDA.t552 48.0005
R2737 GNDA.n2039 GNDA.t31 48.0005
R2738 GNDA.t366 GNDA.n67 47.6748
R2739 GNDA.t297 GNDA.t302 47.5879
R2740 GNDA.t550 GNDA.t218 47.5879
R2741 GNDA.t583 GNDA.t278 47.5879
R2742 GNDA.t588 GNDA.t223 47.5879
R2743 GNDA.t60 GNDA.t329 47.5879
R2744 GNDA.t366 GNDA.n73 47.2907
R2745 GNDA.n428 GNDA.t91 47.2907
R2746 GNDA.t274 GNDA.n1999 46.9995
R2747 GNDA.n793 GNDA.t95 46.2845
R2748 GNDA.n699 GNDA.n697 44.2722
R2749 GNDA.n2126 GNDA.n509 44.0005
R2750 GNDA.n1998 GNDA.n1992 43.9273
R2751 GNDA.n1981 GNDA.n529 43.9273
R2752 GNDA.t111 GNDA.t271 43.9273
R2753 GNDA.t130 GNDA.t319 43.9273
R2754 GNDA.t394 GNDA.t268 43.9273
R2755 GNDA.n2034 GNDA.t140 43.9273
R2756 GNDA.t402 GNDA.t553 43.9273
R2757 GNDA.t8 GNDA.t163 43.9273
R2758 GNDA.t123 GNDA.t59 43.9273
R2759 GNDA.t208 GNDA.t62 43.9273
R2760 GNDA.t245 GNDA.t592 43.9273
R2761 GNDA.n2117 GNDA.n2116 43.9273
R2762 GNDA.n2123 GNDA.n511 43.9273
R2763 GNDA.n2003 GNDA.n2002 43.5649
R2764 GNDA.n792 GNDA.n611 43.266
R2765 GNDA.t366 GNDA.n2211 43.266
R2766 GNDA.t413 GNDA.n657 42.2598
R2767 GNDA.n430 GNDA.t258 42.2598
R2768 GNDA.n777 GNDA.t257 41.2536
R2769 GNDA.n2085 GNDA.t457 40.4338
R2770 GNDA.n2058 GNDA.t435 40.4338
R2771 GNDA.t366 GNDA.n82 40.0547
R2772 GNDA.t366 GNDA.n98 40.0547
R2773 GNDA.n161 GNDA.t366 40.0547
R2774 GNDA.t249 GNDA.t198 39.7296
R2775 GNDA.n794 GNDA.t260 38.2351
R2776 GNDA.n683 GNDA.n324 38.2351
R2777 GNDA.n696 GNDA.t462 38.2351
R2778 GNDA.n2082 GNDA.n2081 37.5297
R2779 GNDA.n2080 GNDA.n2079 37.5297
R2780 GNDA.n2078 GNDA.n2077 37.5297
R2781 GNDA.n2076 GNDA.n2075 37.5297
R2782 GNDA.n2074 GNDA.n2073 37.5297
R2783 GNDA.n2072 GNDA.n2071 37.5297
R2784 GNDA.n2070 GNDA.n2069 37.5297
R2785 GNDA.n2068 GNDA.n2067 37.5297
R2786 GNDA.n2066 GNDA.n2065 37.5297
R2787 GNDA.n2064 GNDA.n2063 37.5297
R2788 GNDA.n2062 GNDA.n2061 37.5297
R2789 GNDA.n1785 GNDA.n1784 37.229
R2790 GNDA.n540 GNDA.t270 37.229
R2791 GNDA.n2410 GNDA.t366 36.6459
R2792 GNDA.t366 GNDA.n2379 36.6459
R2793 GNDA.n168 GNDA.t366 36.6459
R2794 GNDA.t10 GNDA.t271 36.6062
R2795 GNDA.t319 GNDA.t111 36.6062
R2796 GNDA.t130 GNDA.t268 36.6062
R2797 GNDA.t394 GNDA.t583 36.6062
R2798 GNDA.n2034 GNDA.t323 36.6062
R2799 GNDA.t370 GNDA.t250 36.4189
R2800 GNDA.t250 GNDA.t66 36.4189
R2801 GNDA.t66 GNDA.t234 36.4189
R2802 GNDA.n2056 GNDA.t157 35.3897
R2803 GNDA.t300 GNDA.n2088 35.3897
R2804 GNDA.t273 GNDA.n2087 35.3897
R2805 GNDA.n2055 GNDA.t73 35.3897
R2806 GNDA.n2054 GNDA.t179 35.3897
R2807 GNDA.n2053 GNDA.t10 35.3897
R2808 GNDA.t207 GNDA.n2089 35.3897
R2809 GNDA.t95 GNDA.t373 35.2166
R2810 GNDA.t91 GNDA.t405 35.2166
R2811 GNDA.n418 GNDA.t305 33.2043
R2812 GNDA.t285 GNDA.t42 33.1236
R2813 GNDA.t230 GNDA.t43 33.1236
R2814 GNDA.n2170 GNDA.n398 33.0531
R2815 GNDA.n2185 GNDA.n2173 33.0531
R2816 GNDA.n178 GNDA.n142 33.0473
R2817 GNDA.n184 GNDA.n142 33.0473
R2818 GNDA.n185 GNDA.n184 33.0473
R2819 GNDA.n186 GNDA.n185 33.0473
R2820 GNDA.n186 GNDA.n58 33.0473
R2821 GNDA.n193 GNDA.n59 33.0473
R2822 GNDA.n195 GNDA.n193 33.0473
R2823 GNDA.n195 GNDA.n194 33.0473
R2824 GNDA.n194 GNDA.n136 33.0473
R2825 GNDA.n202 GNDA.n136 33.0473
R2826 GNDA.n203 GNDA.n202 33.0473
R2827 GNDA.n203 GNDA.t594 33.0473
R2828 GNDA.n1027 GNDA.n994 33.0473
R2829 GNDA.n1028 GNDA.n1027 33.0473
R2830 GNDA.n1030 GNDA.n1028 33.0473
R2831 GNDA.n1030 GNDA.n1029 33.0473
R2832 GNDA.n1029 GNDA.n60 33.0473
R2833 GNDA.n1037 GNDA.n61 33.0473
R2834 GNDA.n1037 GNDA.n988 33.0473
R2835 GNDA.n1044 GNDA.n988 33.0473
R2836 GNDA.n1045 GNDA.n1044 33.0473
R2837 GNDA.n1046 GNDA.n1045 33.0473
R2838 GNDA.n1046 GNDA.n986 33.0473
R2839 GNDA.n2220 GNDA.n359 33.0473
R2840 GNDA.n2220 GNDA.n2219 33.0473
R2841 GNDA.n2219 GNDA.n2218 33.0473
R2842 GNDA.n2218 GNDA.n360 33.0473
R2843 GNDA.n2212 GNDA.n360 33.0473
R2844 GNDA.n491 GNDA.n364 33.0473
R2845 GNDA.n493 GNDA.n491 33.0473
R2846 GNDA.n493 GNDA.n492 33.0473
R2847 GNDA.n492 GNDA.n487 33.0473
R2848 GNDA.n501 GNDA.n487 33.0473
R2849 GNDA.n502 GNDA.n501 33.0473
R2850 GNDA.t493 GNDA.t297 32.9456
R2851 GNDA.t218 GNDA.t40 32.9456
R2852 GNDA.n2090 GNDA.t592 32.9456
R2853 GNDA.t223 GNDA.t326 32.9456
R2854 GNDA.t220 GNDA.t60 32.9456
R2855 GNDA.n2425 GNDA.t366 32.9056
R2856 GNDA.t366 GNDA.n74 32.9056
R2857 GNDA.n684 GNDA.t585 32.1981
R2858 GNDA.n2019 GNDA.n2018 31.5738
R2859 GNDA.n1993 GNDA.t381 31.1255
R2860 GNDA.n1997 GNDA.t460 31.1255
R2861 GNDA.n2118 GNDA.t427 31.1255
R2862 GNDA.n2122 GNDA.t441 31.1255
R2863 GNDA.n2108 GNDA.n2105 30.8755
R2864 GNDA.n1989 GNDA.n1831 30.813
R2865 GNDA.n2158 GNDA.n2155 30.1857
R2866 GNDA.n712 GNDA.n710 30.1857
R2867 GNDA.n2010 GNDA.n2009 29.8672
R2868 GNDA.n2007 GNDA.n2006 29.8672
R2869 GNDA.n522 GNDA.n521 29.8672
R2870 GNDA.t157 GNDA.n2055 29.4916
R2871 GNDA.t73 GNDA.n2054 29.4916
R2872 GNDA.t179 GNDA.n2053 29.4916
R2873 GNDA.n2089 GNDA.t300 29.4916
R2874 GNDA.t244 GNDA.n2056 29.4916
R2875 GNDA.n2088 GNDA.t273 29.4916
R2876 GNDA.n2087 GNDA.t162 29.4916
R2877 GNDA.t64 GNDA.n793 29.1796
R2878 GNDA.t216 GNDA.n778 28.1734
R2879 GNDA.t194 GNDA.n428 28.1734
R2880 GNDA.n1813 GNDA.t281 28.142
R2881 GNDA.n1628 GNDA.n1625 27.5561
R2882 GNDA.n257 GNDA.n254 27.5561
R2883 GNDA.n1230 GNDA.n1229 27.5561
R2884 GNDA.n754 GNDA.n753 27.5561
R2885 GNDA.n1109 GNDA.n1108 27.5561
R2886 GNDA.n452 GNDA.n449 27.5561
R2887 GNDA.n1726 GNDA.n1723 27.5561
R2888 GNDA.n1354 GNDA.n1351 27.5561
R2889 GNDA.n834 GNDA.n550 27.5561
R2890 GNDA.n2188 GNDA.n2187 27.1672
R2891 GNDA.n1609 GNDA.n1608 26.6672
R2892 GNDA.n238 GNDA.n237 26.6672
R2893 GNDA.n1212 GNDA.n1211 26.6672
R2894 GNDA.n736 GNDA.n735 26.6672
R2895 GNDA.n1091 GNDA.n1090 26.6672
R2896 GNDA.n469 GNDA.n468 26.6672
R2897 GNDA.n1707 GNDA.n1706 26.6672
R2898 GNDA.n1335 GNDA.n1334 26.6672
R2899 GNDA.n812 GNDA.n554 26.6672
R2900 GNDA.n588 GNDA.n587 25.3679
R2901 GNDA.t196 GNDA.t312 25.1549
R2902 GNDA.t154 GNDA.t45 25.1549
R2903 GNDA.n2131 GNDA.n2130 24.1487
R2904 GNDA.n417 GNDA.t579 24.0005
R2905 GNDA.n417 GNDA.t215 24.0005
R2906 GNDA.n416 GNDA.t155 24.0005
R2907 GNDA.n416 GNDA.t233 24.0005
R2908 GNDA.n415 GNDA.t195 24.0005
R2909 GNDA.n415 GNDA.t259 24.0005
R2910 GNDA.n412 GNDA.t14 24.0005
R2911 GNDA.n412 GNDA.t586 24.0005
R2912 GNDA.n411 GNDA.t217 24.0005
R2913 GNDA.n411 GNDA.t237 24.0005
R2914 GNDA.n1803 GNDA.t261 24.0005
R2915 GNDA.n1803 GNDA.t65 24.0005
R2916 GNDA.n1802 GNDA.t16 24.0005
R2917 GNDA.n1802 GNDA.t197 24.0005
R2918 GNDA.n1801 GNDA.t577 24.0005
R2919 GNDA.n1801 GNDA.t153 24.0005
R2920 GNDA.n536 GNDA.t235 24.0005
R2921 GNDA.n536 GNDA.t430 24.0005
R2922 GNDA.n535 GNDA.t251 24.0005
R2923 GNDA.n535 GNDA.t67 24.0005
R2924 GNDA.t156 GNDA.t289 23.7629
R2925 GNDA.t255 GNDA.t156 23.7629
R2926 GNDA.n592 GNDA.n591 23.1425
R2927 GNDA.t366 GNDA.n58 22.3989
R2928 GNDA.t366 GNDA.n60 22.3989
R2929 GNDA.n2212 GNDA.t366 22.3989
R2930 GNDA.t402 GNDA.t54 21.9639
R2931 GNDA.t8 GNDA.t167 21.9639
R2932 GNDA.t59 GNDA.t246 21.9639
R2933 GNDA.t208 GNDA.t144 21.9639
R2934 GNDA.t389 GNDA.t245 21.9639
R2935 GNDA.n1911 GNDA.n1910 21.0192
R2936 GNDA.n1812 GNDA.n1811 20.8233
R2937 GNDA.n2144 GNDA.n2143 20.8233
R2938 GNDA.n698 GNDA.n414 20.8233
R2939 GNDA.n711 GNDA.n413 20.8233
R2940 GNDA.n2154 GNDA.n2153 20.8233
R2941 GNDA.n610 GNDA.n609 20.8233
R2942 GNDA.n1800 GNDA.n1799 20.8233
R2943 GNDA.n1783 GNDA.n537 20.8233
R2944 GNDA.t589 GNDA.t285 20.5905
R2945 GNDA.t43 GNDA.t151 20.5905
R2946 GNDA.n2104 GNDA.t267 19.7005
R2947 GNDA.n2104 GNDA.t532 19.7005
R2948 GNDA.n2102 GNDA.t238 19.7005
R2949 GNDA.n2102 GNDA.t314 19.7005
R2950 GNDA.n2100 GNDA.t241 19.7005
R2951 GNDA.n2100 GNDA.t265 19.7005
R2952 GNDA.n2098 GNDA.t240 19.7005
R2953 GNDA.n2098 GNDA.t231 19.7005
R2954 GNDA.n2096 GNDA.t221 19.7005
R2955 GNDA.n2096 GNDA.t299 19.7005
R2956 GNDA.n2095 GNDA.t540 19.7005
R2957 GNDA.n2095 GNDA.t327 19.7005
R2958 GNDA.n1830 GNDA.t126 19.7005
R2959 GNDA.n1830 GNDA.t348 19.7005
R2960 GNDA.n1828 GNDA.t486 19.7005
R2961 GNDA.n1828 GNDA.t191 19.7005
R2962 GNDA.n1826 GNDA.t328 19.7005
R2963 GNDA.n1826 GNDA.t497 19.7005
R2964 GNDA.n1824 GNDA.t301 19.7005
R2965 GNDA.n1824 GNDA.t347 19.7005
R2966 GNDA.n1822 GNDA.t331 19.7005
R2967 GNDA.n1822 GNDA.t346 19.7005
R2968 GNDA.n1821 GNDA.t304 19.7005
R2969 GNDA.n1821 GNDA.t239 19.7005
R2970 GNDA.t366 GNDA.n62 18.9332
R2971 GNDA.n2382 GNDA.n2381 18.5605
R2972 GNDA.n2020 GNDA.n2019 18.4151
R2973 GNDA.n503 GNDA.t45 18.3598
R2974 GNDA.n505 GNDA.t45 18.3598
R2975 GNDA.t498 GNDA.t28 18.3033
R2976 GNDA.t336 GNDA.t39 18.3033
R2977 GNDA.n2033 GNDA.t173 18.3033
R2978 GNDA.t290 GNDA.t313 18.3033
R2979 GNDA.t199 GNDA.t321 18.3033
R2980 GNDA.n2029 GNDA.n522 18.0922
R2981 GNDA.n1024 GNDA.n1023 17.5843
R2982 GNDA.n2224 GNDA.n2223 17.5843
R2983 GNDA.n180 GNDA.n144 17.5843
R2984 GNDA.t366 GNDA.n2424 17.0449
R2985 GNDA.n2422 GNDA.n79 16.9379
R2986 GNDA.n1407 GNDA.n1403 16.9379
R2987 GNDA.n916 GNDA.n898 16.9379
R2988 GNDA.n2342 GNDA.n2339 16.7709
R2989 GNDA.n2245 GNDA.n307 16.7709
R2990 GNDA.n2311 GNDA.n2310 16.7709
R2991 GNDA.n1656 GNDA.n1504 16.7709
R2992 GNDA.t281 GNDA.t370 16.5543
R2993 GNDA.n1988 GNDA.n1987 16.2608
R2994 GNDA.n1986 GNDA.n1985 16.2608
R2995 GNDA.n2112 GNDA.n2111 16.2608
R2996 GNDA.n2110 GNDA.n2109 16.2608
R2997 GNDA.n1629 GNDA.n1628 16.0005
R2998 GNDA.n1632 GNDA.n1629 16.0005
R2999 GNDA.n1633 GNDA.n1632 16.0005
R3000 GNDA.n1636 GNDA.n1633 16.0005
R3001 GNDA.n1637 GNDA.n1636 16.0005
R3002 GNDA.n1640 GNDA.n1637 16.0005
R3003 GNDA.n1641 GNDA.n1640 16.0005
R3004 GNDA.n1641 GNDA.n1541 16.0005
R3005 GNDA.n1625 GNDA.n1624 16.0005
R3006 GNDA.n1624 GNDA.n1621 16.0005
R3007 GNDA.n1621 GNDA.n1620 16.0005
R3008 GNDA.n1620 GNDA.n1617 16.0005
R3009 GNDA.n1617 GNDA.n1616 16.0005
R3010 GNDA.n1616 GNDA.n1613 16.0005
R3011 GNDA.n1613 GNDA.n1612 16.0005
R3012 GNDA.n1612 GNDA.n1609 16.0005
R3013 GNDA.n1608 GNDA.n1605 16.0005
R3014 GNDA.n1605 GNDA.n1604 16.0005
R3015 GNDA.n1604 GNDA.n1601 16.0005
R3016 GNDA.n1601 GNDA.n1600 16.0005
R3017 GNDA.n1600 GNDA.n1597 16.0005
R3018 GNDA.n1597 GNDA.n1596 16.0005
R3019 GNDA.n1596 GNDA.n1593 16.0005
R3020 GNDA.n1593 GNDA.n1592 16.0005
R3021 GNDA.n258 GNDA.n257 16.0005
R3022 GNDA.n261 GNDA.n258 16.0005
R3023 GNDA.n262 GNDA.n261 16.0005
R3024 GNDA.n265 GNDA.n262 16.0005
R3025 GNDA.n266 GNDA.n265 16.0005
R3026 GNDA.n269 GNDA.n266 16.0005
R3027 GNDA.n271 GNDA.n269 16.0005
R3028 GNDA.n272 GNDA.n271 16.0005
R3029 GNDA.n254 GNDA.n253 16.0005
R3030 GNDA.n253 GNDA.n250 16.0005
R3031 GNDA.n250 GNDA.n249 16.0005
R3032 GNDA.n249 GNDA.n246 16.0005
R3033 GNDA.n246 GNDA.n245 16.0005
R3034 GNDA.n245 GNDA.n242 16.0005
R3035 GNDA.n242 GNDA.n241 16.0005
R3036 GNDA.n241 GNDA.n238 16.0005
R3037 GNDA.n237 GNDA.n234 16.0005
R3038 GNDA.n234 GNDA.n233 16.0005
R3039 GNDA.n233 GNDA.n230 16.0005
R3040 GNDA.n230 GNDA.n229 16.0005
R3041 GNDA.n229 GNDA.n226 16.0005
R3042 GNDA.n226 GNDA.n225 16.0005
R3043 GNDA.n225 GNDA.n222 16.0005
R3044 GNDA.n222 GNDA.n221 16.0005
R3045 GNDA.n1244 GNDA.n1230 16.0005
R3046 GNDA.n1244 GNDA.n1243 16.0005
R3047 GNDA.n1243 GNDA.n1242 16.0005
R3048 GNDA.n1242 GNDA.n1239 16.0005
R3049 GNDA.n1239 GNDA.n1238 16.0005
R3050 GNDA.n1238 GNDA.n1235 16.0005
R3051 GNDA.n1235 GNDA.n1234 16.0005
R3052 GNDA.n1234 GNDA.n1231 16.0005
R3053 GNDA.n1229 GNDA.n1227 16.0005
R3054 GNDA.n1227 GNDA.n1224 16.0005
R3055 GNDA.n1224 GNDA.n1223 16.0005
R3056 GNDA.n1223 GNDA.n1220 16.0005
R3057 GNDA.n1220 GNDA.n1219 16.0005
R3058 GNDA.n1219 GNDA.n1216 16.0005
R3059 GNDA.n1216 GNDA.n1215 16.0005
R3060 GNDA.n1215 GNDA.n1212 16.0005
R3061 GNDA.n1211 GNDA.n1208 16.0005
R3062 GNDA.n1208 GNDA.n1207 16.0005
R3063 GNDA.n1207 GNDA.n1204 16.0005
R3064 GNDA.n1204 GNDA.n1203 16.0005
R3065 GNDA.n1203 GNDA.n1200 16.0005
R3066 GNDA.n1200 GNDA.n1199 16.0005
R3067 GNDA.n1199 GNDA.n1196 16.0005
R3068 GNDA.n1196 GNDA.n1195 16.0005
R3069 GNDA.n767 GNDA.n754 16.0005
R3070 GNDA.n767 GNDA.n766 16.0005
R3071 GNDA.n766 GNDA.n765 16.0005
R3072 GNDA.n765 GNDA.n762 16.0005
R3073 GNDA.n762 GNDA.n761 16.0005
R3074 GNDA.n761 GNDA.n758 16.0005
R3075 GNDA.n758 GNDA.n757 16.0005
R3076 GNDA.n757 GNDA.n650 16.0005
R3077 GNDA.n753 GNDA.n751 16.0005
R3078 GNDA.n751 GNDA.n748 16.0005
R3079 GNDA.n748 GNDA.n747 16.0005
R3080 GNDA.n747 GNDA.n744 16.0005
R3081 GNDA.n744 GNDA.n743 16.0005
R3082 GNDA.n743 GNDA.n740 16.0005
R3083 GNDA.n740 GNDA.n739 16.0005
R3084 GNDA.n739 GNDA.n736 16.0005
R3085 GNDA.n735 GNDA.n732 16.0005
R3086 GNDA.n732 GNDA.n731 16.0005
R3087 GNDA.n731 GNDA.n728 16.0005
R3088 GNDA.n728 GNDA.n727 16.0005
R3089 GNDA.n727 GNDA.n724 16.0005
R3090 GNDA.n724 GNDA.n723 16.0005
R3091 GNDA.n723 GNDA.n720 16.0005
R3092 GNDA.n720 GNDA.n719 16.0005
R3093 GNDA.n1123 GNDA.n1109 16.0005
R3094 GNDA.n1123 GNDA.n1122 16.0005
R3095 GNDA.n1122 GNDA.n1121 16.0005
R3096 GNDA.n1121 GNDA.n1118 16.0005
R3097 GNDA.n1118 GNDA.n1117 16.0005
R3098 GNDA.n1117 GNDA.n1114 16.0005
R3099 GNDA.n1114 GNDA.n1113 16.0005
R3100 GNDA.n1113 GNDA.n1110 16.0005
R3101 GNDA.n1108 GNDA.n1106 16.0005
R3102 GNDA.n1106 GNDA.n1103 16.0005
R3103 GNDA.n1103 GNDA.n1102 16.0005
R3104 GNDA.n1102 GNDA.n1099 16.0005
R3105 GNDA.n1099 GNDA.n1098 16.0005
R3106 GNDA.n1098 GNDA.n1095 16.0005
R3107 GNDA.n1095 GNDA.n1094 16.0005
R3108 GNDA.n1094 GNDA.n1091 16.0005
R3109 GNDA.n1090 GNDA.n1087 16.0005
R3110 GNDA.n1087 GNDA.n1086 16.0005
R3111 GNDA.n1086 GNDA.n1083 16.0005
R3112 GNDA.n1083 GNDA.n1082 16.0005
R3113 GNDA.n1082 GNDA.n1079 16.0005
R3114 GNDA.n1079 GNDA.n1078 16.0005
R3115 GNDA.n1078 GNDA.n1075 16.0005
R3116 GNDA.n1075 GNDA.n1074 16.0005
R3117 GNDA.n449 GNDA.n448 16.0005
R3118 GNDA.n448 GNDA.n445 16.0005
R3119 GNDA.n445 GNDA.n444 16.0005
R3120 GNDA.n444 GNDA.n441 16.0005
R3121 GNDA.n441 GNDA.n440 16.0005
R3122 GNDA.n440 GNDA.n437 16.0005
R3123 GNDA.n437 GNDA.n436 16.0005
R3124 GNDA.n436 GNDA.n434 16.0005
R3125 GNDA.n453 GNDA.n452 16.0005
R3126 GNDA.n456 GNDA.n453 16.0005
R3127 GNDA.n457 GNDA.n456 16.0005
R3128 GNDA.n460 GNDA.n457 16.0005
R3129 GNDA.n461 GNDA.n460 16.0005
R3130 GNDA.n464 GNDA.n461 16.0005
R3131 GNDA.n465 GNDA.n464 16.0005
R3132 GNDA.n468 GNDA.n465 16.0005
R3133 GNDA.n472 GNDA.n469 16.0005
R3134 GNDA.n473 GNDA.n472 16.0005
R3135 GNDA.n476 GNDA.n473 16.0005
R3136 GNDA.n477 GNDA.n476 16.0005
R3137 GNDA.n480 GNDA.n477 16.0005
R3138 GNDA.n481 GNDA.n480 16.0005
R3139 GNDA.n484 GNDA.n481 16.0005
R3140 GNDA.n2135 GNDA.n484 16.0005
R3141 GNDA.n1727 GNDA.n1726 16.0005
R3142 GNDA.n1730 GNDA.n1727 16.0005
R3143 GNDA.n1731 GNDA.n1730 16.0005
R3144 GNDA.n1734 GNDA.n1731 16.0005
R3145 GNDA.n1735 GNDA.n1734 16.0005
R3146 GNDA.n1738 GNDA.n1735 16.0005
R3147 GNDA.n1739 GNDA.n1738 16.0005
R3148 GNDA.n1739 GNDA.n921 16.0005
R3149 GNDA.n1723 GNDA.n1722 16.0005
R3150 GNDA.n1722 GNDA.n1719 16.0005
R3151 GNDA.n1719 GNDA.n1718 16.0005
R3152 GNDA.n1718 GNDA.n1715 16.0005
R3153 GNDA.n1715 GNDA.n1714 16.0005
R3154 GNDA.n1714 GNDA.n1711 16.0005
R3155 GNDA.n1711 GNDA.n1710 16.0005
R3156 GNDA.n1710 GNDA.n1707 16.0005
R3157 GNDA.n1706 GNDA.n1703 16.0005
R3158 GNDA.n1703 GNDA.n1702 16.0005
R3159 GNDA.n1702 GNDA.n1699 16.0005
R3160 GNDA.n1699 GNDA.n1698 16.0005
R3161 GNDA.n1698 GNDA.n1695 16.0005
R3162 GNDA.n1695 GNDA.n1694 16.0005
R3163 GNDA.n1694 GNDA.n1691 16.0005
R3164 GNDA.n1691 GNDA.n1690 16.0005
R3165 GNDA.n1355 GNDA.n1354 16.0005
R3166 GNDA.n1358 GNDA.n1355 16.0005
R3167 GNDA.n1359 GNDA.n1358 16.0005
R3168 GNDA.n1362 GNDA.n1359 16.0005
R3169 GNDA.n1363 GNDA.n1362 16.0005
R3170 GNDA.n1366 GNDA.n1363 16.0005
R3171 GNDA.n1367 GNDA.n1366 16.0005
R3172 GNDA.n1370 GNDA.n1367 16.0005
R3173 GNDA.n1351 GNDA.n1350 16.0005
R3174 GNDA.n1350 GNDA.n1347 16.0005
R3175 GNDA.n1347 GNDA.n1346 16.0005
R3176 GNDA.n1346 GNDA.n1343 16.0005
R3177 GNDA.n1343 GNDA.n1342 16.0005
R3178 GNDA.n1342 GNDA.n1339 16.0005
R3179 GNDA.n1339 GNDA.n1338 16.0005
R3180 GNDA.n1338 GNDA.n1335 16.0005
R3181 GNDA.n1334 GNDA.n1331 16.0005
R3182 GNDA.n1331 GNDA.n1330 16.0005
R3183 GNDA.n1330 GNDA.n1327 16.0005
R3184 GNDA.n1327 GNDA.n1326 16.0005
R3185 GNDA.n1326 GNDA.n1323 16.0005
R3186 GNDA.n1323 GNDA.n1322 16.0005
R3187 GNDA.n1322 GNDA.n1319 16.0005
R3188 GNDA.n1319 GNDA.n1318 16.0005
R3189 GNDA.n835 GNDA.n834 16.0005
R3190 GNDA.n836 GNDA.n835 16.0005
R3191 GNDA.n836 GNDA.n548 16.0005
R3192 GNDA.n842 GNDA.n548 16.0005
R3193 GNDA.n843 GNDA.n842 16.0005
R3194 GNDA.n844 GNDA.n843 16.0005
R3195 GNDA.n844 GNDA.n546 16.0005
R3196 GNDA.n849 GNDA.n546 16.0005
R3197 GNDA.n828 GNDA.n550 16.0005
R3198 GNDA.n828 GNDA.n827 16.0005
R3199 GNDA.n827 GNDA.n826 16.0005
R3200 GNDA.n826 GNDA.n552 16.0005
R3201 GNDA.n820 GNDA.n552 16.0005
R3202 GNDA.n820 GNDA.n819 16.0005
R3203 GNDA.n819 GNDA.n818 16.0005
R3204 GNDA.n818 GNDA.n554 16.0005
R3205 GNDA.n812 GNDA.n811 16.0005
R3206 GNDA.n811 GNDA.n810 16.0005
R3207 GNDA.n810 GNDA.n556 16.0005
R3208 GNDA.n805 GNDA.n556 16.0005
R3209 GNDA.n805 GNDA.n804 16.0005
R3210 GNDA.n804 GNDA.n803 16.0005
R3211 GNDA.n803 GNDA.n559 16.0005
R3212 GNDA.n798 GNDA.n559 16.0005
R3213 GNDA.n1910 GNDA.n101 16.0005
R3214 GNDA.n2381 GNDA.n101 16.0005
R3215 GNDA.n1930 GNDA.n1929 15.3599
R3216 GNDA.n2035 GNDA.n2034 15.1729
R3217 GNDA.t366 GNDA.t576 15.0931
R3218 GNDA.t366 GNDA.t214 15.0931
R3219 GNDA.n2057 GNDA.t178 14.7463
R3220 GNDA.n2086 GNDA.t9 14.7463
R3221 GNDA.t278 GNDA.n2033 14.6428
R3222 GNDA.t446 GNDA.t590 14.6428
R3223 GNDA.t276 GNDA.t54 14.6428
R3224 GNDA.t553 GNDA.t167 14.6428
R3225 GNDA.t163 GNDA.t246 14.6428
R3226 GNDA.t144 GNDA.t123 14.6428
R3227 GNDA.t62 GNDA.t389 14.6428
R3228 GNDA.n1913 GNDA.n1912 14.563
R3229 GNDA.n2426 GNDA.n2425 14.555
R3230 GNDA.n1379 GNDA.n74 14.555
R3231 GNDA.n2011 GNDA.n2010 14.1651
R3232 GNDA.n2006 GNDA.n520 14.0922
R3233 GNDA.n708 GNDA.n707 12.8005
R3234 GNDA.n707 GNDA.n704 12.8005
R3235 GNDA.n2160 GNDA.n406 12.8005
R3236 GNDA.n2156 GNDA.n406 12.8005
R3237 GNDA.n1991 GNDA.t387 12.6791
R3238 GNDA.n1982 GNDA.t377 12.6791
R3239 GNDA.n2115 GNDA.t444 12.6791
R3240 GNDA.n2106 GNDA.t438 12.6791
R3241 GNDA.n2049 GNDA.n516 12.2505
R3242 GNDA.n593 GNDA.t15 12.0746
R3243 GNDA.t13 GNDA.n683 12.0746
R3244 GNDA.n2198 GNDA.t578 12.0746
R3245 GNDA.n1455 GNDA.n944 11.6369
R3246 GNDA.n1455 GNDA.n1454 11.6369
R3247 GNDA.n1454 GNDA.n1453 11.6369
R3248 GNDA.n1453 GNDA.n1432 11.6369
R3249 GNDA.n1448 GNDA.n1432 11.6369
R3250 GNDA.n1448 GNDA.n1447 11.6369
R3251 GNDA.n1447 GNDA.n1446 11.6369
R3252 GNDA.n1446 GNDA.n1435 11.6369
R3253 GNDA.n1441 GNDA.n1435 11.6369
R3254 GNDA.n1441 GNDA.n1440 11.6369
R3255 GNDA.n1440 GNDA.n278 11.6369
R3256 GNDA.n1003 GNDA.n279 11.6369
R3257 GNDA.n1004 GNDA.n1003 11.6369
R3258 GNDA.n1004 GNDA.n1000 11.6369
R3259 GNDA.n1010 GNDA.n1000 11.6369
R3260 GNDA.n1011 GNDA.n1010 11.6369
R3261 GNDA.n1012 GNDA.n1011 11.6369
R3262 GNDA.n1012 GNDA.n998 11.6369
R3263 GNDA.n1017 GNDA.n998 11.6369
R3264 GNDA.n1018 GNDA.n1017 11.6369
R3265 GNDA.n1018 GNDA.n996 11.6369
R3266 GNDA.n1023 GNDA.n996 11.6369
R3267 GNDA.n1025 GNDA.n1024 11.6369
R3268 GNDA.n1025 GNDA.n992 11.6369
R3269 GNDA.n1032 GNDA.n992 11.6369
R3270 GNDA.n1033 GNDA.n1032 11.6369
R3271 GNDA.n1034 GNDA.n1033 11.6369
R3272 GNDA.n1034 GNDA.n990 11.6369
R3273 GNDA.n1039 GNDA.n990 11.6369
R3274 GNDA.n1040 GNDA.n1039 11.6369
R3275 GNDA.n1042 GNDA.n1040 11.6369
R3276 GNDA.n1042 GNDA.n1041 11.6369
R3277 GNDA.n2244 GNDA.n2243 11.6369
R3278 GNDA.n2243 GNDA.n348 11.6369
R3279 GNDA.n2238 GNDA.n348 11.6369
R3280 GNDA.n2238 GNDA.n2237 11.6369
R3281 GNDA.n2237 GNDA.n2236 11.6369
R3282 GNDA.n2236 GNDA.n351 11.6369
R3283 GNDA.n2231 GNDA.n351 11.6369
R3284 GNDA.n2231 GNDA.n2230 11.6369
R3285 GNDA.n2230 GNDA.n2229 11.6369
R3286 GNDA.n2229 GNDA.n354 11.6369
R3287 GNDA.n2224 GNDA.n354 11.6369
R3288 GNDA.n2223 GNDA.n2222 11.6369
R3289 GNDA.n2222 GNDA.n357 11.6369
R3290 GNDA.n2216 GNDA.n357 11.6369
R3291 GNDA.n2216 GNDA.n2215 11.6369
R3292 GNDA.n2215 GNDA.n2214 11.6369
R3293 GNDA.n2214 GNDA.n362 11.6369
R3294 GNDA.n489 GNDA.n362 11.6369
R3295 GNDA.n495 GNDA.n489 11.6369
R3296 GNDA.n496 GNDA.n495 11.6369
R3297 GNDA.n497 GNDA.n496 11.6369
R3298 GNDA.n2422 GNDA.n2421 11.6369
R3299 GNDA.n2421 GNDA.n2420 11.6369
R3300 GNDA.n2420 GNDA.n80 11.6369
R3301 GNDA.n2414 GNDA.n80 11.6369
R3302 GNDA.n2414 GNDA.n2413 11.6369
R3303 GNDA.n2413 GNDA.n2412 11.6369
R3304 GNDA.n2412 GNDA.n84 11.6369
R3305 GNDA.n2406 GNDA.n84 11.6369
R3306 GNDA.n2406 GNDA.n2405 11.6369
R3307 GNDA.n2405 GNDA.n2404 11.6369
R3308 GNDA.n2404 GNDA.n88 11.6369
R3309 GNDA.n1773 GNDA.n79 11.6369
R3310 GNDA.n1773 GNDA.n1772 11.6369
R3311 GNDA.n1772 GNDA.n1771 11.6369
R3312 GNDA.n1771 GNDA.n1769 11.6369
R3313 GNDA.n1769 GNDA.n1766 11.6369
R3314 GNDA.n1766 GNDA.n1765 11.6369
R3315 GNDA.n1765 GNDA.n1762 11.6369
R3316 GNDA.n1762 GNDA.n1761 11.6369
R3317 GNDA.n1761 GNDA.n1758 11.6369
R3318 GNDA.n1758 GNDA.n1757 11.6369
R3319 GNDA.n1408 GNDA.n1407 11.6369
R3320 GNDA.n1409 GNDA.n1408 11.6369
R3321 GNDA.n1409 GNDA.n949 11.6369
R3322 GNDA.n1415 GNDA.n949 11.6369
R3323 GNDA.n1416 GNDA.n1415 11.6369
R3324 GNDA.n1417 GNDA.n1416 11.6369
R3325 GNDA.n1417 GNDA.n947 11.6369
R3326 GNDA.n1423 GNDA.n947 11.6369
R3327 GNDA.n1424 GNDA.n1423 11.6369
R3328 GNDA.n1425 GNDA.n1424 11.6369
R3329 GNDA.n1425 GNDA.n945 11.6369
R3330 GNDA.n1403 GNDA.n1402 11.6369
R3331 GNDA.n1402 GNDA.n1399 11.6369
R3332 GNDA.n1399 GNDA.n1398 11.6369
R3333 GNDA.n1398 GNDA.n1395 11.6369
R3334 GNDA.n1395 GNDA.n1394 11.6369
R3335 GNDA.n1394 GNDA.n1391 11.6369
R3336 GNDA.n1391 GNDA.n1390 11.6369
R3337 GNDA.n1390 GNDA.n1387 11.6369
R3338 GNDA.n1387 GNDA.n1386 11.6369
R3339 GNDA.n1386 GNDA.n1384 11.6369
R3340 GNDA.n916 GNDA.n915 11.6369
R3341 GNDA.n915 GNDA.n914 11.6369
R3342 GNDA.n914 GNDA.n912 11.6369
R3343 GNDA.n912 GNDA.n909 11.6369
R3344 GNDA.n909 GNDA.n908 11.6369
R3345 GNDA.n908 GNDA.n905 11.6369
R3346 GNDA.n905 GNDA.n904 11.6369
R3347 GNDA.n904 GNDA.n901 11.6369
R3348 GNDA.n901 GNDA.n900 11.6369
R3349 GNDA.n900 GNDA.n852 11.6369
R3350 GNDA.n156 GNDA.n111 11.6369
R3351 GNDA.n157 GNDA.n156 11.6369
R3352 GNDA.n157 GNDA.n151 11.6369
R3353 GNDA.n164 GNDA.n151 11.6369
R3354 GNDA.n165 GNDA.n164 11.6369
R3355 GNDA.n166 GNDA.n165 11.6369
R3356 GNDA.n166 GNDA.n148 11.6369
R3357 GNDA.n172 GNDA.n148 11.6369
R3358 GNDA.n173 GNDA.n172 11.6369
R3359 GNDA.n174 GNDA.n173 11.6369
R3360 GNDA.n174 GNDA.n144 11.6369
R3361 GNDA.n181 GNDA.n180 11.6369
R3362 GNDA.n182 GNDA.n181 11.6369
R3363 GNDA.n182 GNDA.n140 11.6369
R3364 GNDA.n188 GNDA.n140 11.6369
R3365 GNDA.n189 GNDA.n188 11.6369
R3366 GNDA.n190 GNDA.n189 11.6369
R3367 GNDA.n190 GNDA.n138 11.6369
R3368 GNDA.n197 GNDA.n138 11.6369
R3369 GNDA.n198 GNDA.n197 11.6369
R3370 GNDA.n199 GNDA.n198 11.6369
R3371 GNDA.n2251 GNDA.n313 11.6369
R3372 GNDA.n2256 GNDA.n2251 11.6369
R3373 GNDA.n2257 GNDA.n2256 11.6369
R3374 GNDA.n2258 GNDA.n2257 11.6369
R3375 GNDA.n2258 GNDA.n2249 11.6369
R3376 GNDA.n2264 GNDA.n2249 11.6369
R3377 GNDA.n2265 GNDA.n2264 11.6369
R3378 GNDA.n2266 GNDA.n2265 11.6369
R3379 GNDA.n2266 GNDA.n2247 11.6369
R3380 GNDA.n2271 GNDA.n2247 11.6369
R3381 GNDA.n2272 GNDA.n2271 11.6369
R3382 GNDA.n898 GNDA.n897 11.6369
R3383 GNDA.n897 GNDA.n871 11.6369
R3384 GNDA.n892 GNDA.n871 11.6369
R3385 GNDA.n892 GNDA.n891 11.6369
R3386 GNDA.n891 GNDA.n890 11.6369
R3387 GNDA.n890 GNDA.n874 11.6369
R3388 GNDA.n885 GNDA.n874 11.6369
R3389 GNDA.n885 GNDA.n884 11.6369
R3390 GNDA.n884 GNDA.n883 11.6369
R3391 GNDA.n883 GNDA.n877 11.6369
R3392 GNDA.n877 GNDA.n314 11.6369
R3393 GNDA.n2392 GNDA.n2391 11.6369
R3394 GNDA.n2391 GNDA.n2390 11.6369
R3395 GNDA.n2390 GNDA.n95 11.6369
R3396 GNDA.n2384 GNDA.n95 11.6369
R3397 GNDA.n2384 GNDA.n2383 11.6369
R3398 GNDA.n2376 GNDA.n100 11.6369
R3399 GNDA.n2376 GNDA.n2375 11.6369
R3400 GNDA.n2375 GNDA.n2374 11.6369
R3401 GNDA.n2374 GNDA.n106 11.6369
R3402 GNDA.n2368 GNDA.n106 11.6369
R3403 GNDA.t198 GNDA.n1813 11.5882
R3404 GNDA.n2145 GNDA.n2144 10.9846
R3405 GNDA.n1811 GNDA.n1810 10.9836
R3406 GNDA.n2148 GNDA.n414 10.87
R3407 GNDA.n2149 GNDA.n413 10.87
R3408 GNDA.n2153 GNDA.n2152 10.87
R3409 GNDA.n609 GNDA.n410 10.87
R3410 GNDA.n1807 GNDA.n1800 10.87
R3411 GNDA.n1808 GNDA.n537 10.87
R3412 GNDA.t366 GNDA.n59 10.6489
R3413 GNDA.t366 GNDA.n61 10.6489
R3414 GNDA.t366 GNDA.n364 10.6489
R3415 GNDA.n1979 GNDA.n1978 9.71925
R3416 GNDA.n2181 GNDA.t98 9.6005
R3417 GNDA.n2184 GNDA.t92 9.6005
R3418 GNDA.n580 GNDA.t94 9.6005
R3419 GNDA.n586 GNDA.t96 9.6005
R3420 GNDA.n2081 GNDA.t213 9.6005
R3421 GNDA.n2081 GNDA.t456 9.6005
R3422 GNDA.n2079 GNDA.t593 9.6005
R3423 GNDA.n2079 GNDA.t309 9.6005
R3424 GNDA.n2077 GNDA.t124 9.6005
R3425 GNDA.n2077 GNDA.t63 9.6005
R3426 GNDA.n2075 GNDA.t554 9.6005
R3427 GNDA.n2075 GNDA.t164 9.6005
R3428 GNDA.n2073 GNDA.t591 9.6005
R3429 GNDA.n2073 GNDA.t277 9.6005
R3430 GNDA.n2071 GNDA.t555 9.6005
R3431 GNDA.n2071 GNDA.t263 9.6005
R3432 GNDA.n2069 GNDA.t172 9.6005
R3433 GNDA.n2069 GNDA.t338 9.6005
R3434 GNDA.n2067 GNDA.t584 9.6005
R3435 GNDA.n2067 GNDA.t174 9.6005
R3436 GNDA.n2065 GNDA.t320 9.6005
R3437 GNDA.n2065 GNDA.t269 9.6005
R3438 GNDA.n2063 GNDA.t311 9.6005
R3439 GNDA.n2063 GNDA.t272 9.6005
R3440 GNDA.n2061 GNDA.t284 9.6005
R3441 GNDA.n2061 GNDA.t318 9.6005
R3442 GNDA.n2051 GNDA.n2050 9.52967
R3443 GNDA.n2038 GNDA.n2037 9.52967
R3444 GNDA.n708 GNDA.n703 9.36264
R3445 GNDA.n2156 GNDA.n404 9.36264
R3446 GNDA.n707 GNDA.n706 9.3005
R3447 GNDA.n705 GNDA.n704 9.3005
R3448 GNDA.n406 GNDA.n405 9.3005
R3449 GNDA.n2161 GNDA.n2160 9.3005
R3450 GNDA.n1996 GNDA.n1995 9.0005
R3451 GNDA.n2121 GNDA.n2120 9.0005
R3452 GNDA.n2120 GNDA.n512 8.90675
R3453 GNDA.n2425 GNDA.n54 8.60107
R3454 GNDA.n2313 GNDA.n74 8.60107
R3455 GNDA.n1782 GNDA.t429 8.04989
R3456 GNDA.n594 GNDA.t152 8.04989
R3457 GNDA.t236 GNDA.n777 8.04989
R3458 GNDA.t232 GNDA.n2199 8.04989
R3459 GNDA.n2094 GNDA.n512 7.46925
R3460 GNDA.n1980 GNDA.n515 7.40675
R3461 GNDA.n2083 GNDA.n512 7.09425
R3462 GNDA.n1797 GNDA.t125 7.04372
R3463 GNDA.t312 GNDA.n607 7.04372
R3464 GNDA.n713 GNDA.n712 7.04372
R3465 GNDA.n2142 GNDA.n419 7.04372
R3466 GNDA.n2060 GNDA.n515 7.03175
R3467 GNDA.n2000 GNDA.t255 6.93119
R3468 GNDA.n2339 GNDA.n278 6.72373
R3469 GNDA.n94 GNDA.n88 6.72373
R3470 GNDA.n1504 GNDA.n945 6.72373
R3471 GNDA.n2272 GNDA.n2245 6.72373
R3472 GNDA.n2310 GNDA.n314 6.72373
R3473 GNDA.n2368 GNDA.n2367 6.72373
R3474 GNDA.n1980 GNDA.n1979 6.313
R3475 GNDA.n1504 GNDA.n944 6.20656
R3476 GNDA.n2339 GNDA.n279 6.20656
R3477 GNDA.n2245 GNDA.n2244 6.20656
R3478 GNDA.n2367 GNDA.n111 6.20656
R3479 GNDA.n2310 GNDA.n313 6.20656
R3480 GNDA.n2392 GNDA.n94 6.20656
R3481 GNDA.n2383 GNDA.n2382 6.07727
R3482 GNDA.t366 GNDA.t257 6.03755
R3483 GNDA.t366 GNDA.t165 5.87549
R3484 GNDA.n588 GNDA.n398 5.81868
R3485 GNDA.n588 GNDA.n579 5.81868
R3486 GNDA.n2382 GNDA.n100 5.5601
R3487 GNDA.n1592 GNDA.n1562 5.51161
R3488 GNDA.n221 GNDA.n207 5.51161
R3489 GNDA.n1195 GNDA.n1173 5.51161
R3490 GNDA.n719 GNDA.n678 5.51161
R3491 GNDA.n1074 GNDA.n1052 5.51161
R3492 GNDA.n2135 GNDA.n2134 5.51161
R3493 GNDA.n1690 GNDA.n1660 5.51161
R3494 GNDA.n1318 GNDA.n1289 5.51161
R3495 GNDA.n798 GNDA.n797 5.51161
R3496 GNDA.t594 GNDA.t41 5.5083
R3497 GNDA.n520 GNDA.n516 5.5005
R3498 GNDA.n1051 GNDA.n985 5.1717
R3499 GNDA.n2133 GNDA.n485 5.1717
R3500 GNDA.n206 GNDA.n134 5.1717
R3501 GNDA.n2040 GNDA.n2038 5.063
R3502 GNDA.t270 GNDA.t452 5.03137
R3503 GNDA.n591 GNDA.t576 5.03137
R3504 GNDA.t366 GNDA.n324 5.03137
R3505 GNDA.t405 GNDA.t366 5.03137
R3506 GNDA.n2187 GNDA.t214 5.03137
R3507 GNDA.t305 GNDA.t449 5.03137
R3508 GNDA.n523 GNDA.n514 5.02133
R3509 GNDA.n2093 GNDA.n2092 5.02133
R3510 GNDA.n1995 GNDA.n1994 5.0005
R3511 GNDA.n2120 GNDA.n2119 5.0005
R3512 GNDA.t234 GNDA.t93 4.96664
R3513 GNDA.n1984 GNDA.n1983 4.91717
R3514 GNDA.n2114 GNDA.n2113 4.91717
R3515 GNDA.n2108 GNDA.n2107 4.91717
R3516 GNDA.n1990 GNDA.n1989 4.91717
R3517 GNDA.n1754 GNDA.n1751 4.9157
R3518 GNDA.n1383 GNDA.n952 4.9157
R3519 GNDA.n1780 GNDA.n1779 4.9157
R3520 GNDA.n2017 GNDA.n2016 4.86508
R3521 GNDA.n2022 GNDA.n2020 4.86508
R3522 GNDA.n2031 GNDA.n2030 4.79217
R3523 GNDA.n2029 GNDA.n2028 4.79217
R3524 GNDA.n397 GNDA.n396 4.5005
R3525 GNDA.n2163 GNDA.n400 4.5005
R3526 GNDA.n2165 GNDA.n2164 4.5005
R3527 GNDA.n2164 GNDA.n2163 4.5005
R3528 GNDA.n705 GNDA.n402 4.5005
R3529 GNDA.n2162 GNDA.n2161 4.5005
R3530 GNDA.n1978 GNDA.n1977 4.5005
R3531 GNDA.n1976 GNDA.n1832 4.5005
R3532 GNDA.n1975 GNDA.n1974 4.5005
R3533 GNDA.n1973 GNDA.n1836 4.5005
R3534 GNDA.n2050 GNDA.n2049 4.5005
R3535 GNDA.n528 GNDA.n527 4.5005
R3536 GNDA.n2060 GNDA.n2059 4.5005
R3537 GNDA.n2084 GNDA.n2083 4.5005
R3538 GNDA.n1904 GNDA.n1900 4.5005
R3539 GNDA.n1908 GNDA.n1907 4.5005
R3540 GNDA.n1909 GNDA.n1899 4.5005
R3541 GNDA.n1914 GNDA.n1913 4.5005
R3542 GNDA.n1923 GNDA.n1919 4.5005
R3543 GNDA.n1927 GNDA.n1926 4.5005
R3544 GNDA.n1928 GNDA.n1918 4.5005
R3545 GNDA.n1931 GNDA.n1930 4.5005
R3546 GNDA.n2366 GNDA.n112 4.26717
R3547 GNDA.n2360 GNDA.n112 4.26717
R3548 GNDA.n2360 GNDA.n2359 4.26717
R3549 GNDA.n2359 GNDA.n2358 4.26717
R3550 GNDA.n2358 GNDA.n121 4.26717
R3551 GNDA.n2353 GNDA.n121 4.26717
R3552 GNDA.n2353 GNDA.n2352 4.26717
R3553 GNDA.n2352 GNDA.n2351 4.26717
R3554 GNDA.n2351 GNDA.n127 4.26717
R3555 GNDA.n2345 GNDA.n127 4.26717
R3556 GNDA.n2345 GNDA.n2344 4.26717
R3557 GNDA.n2338 GNDA.n281 4.26717
R3558 GNDA.n2333 GNDA.n281 4.26717
R3559 GNDA.n2333 GNDA.n2332 4.26717
R3560 GNDA.n2332 GNDA.n289 4.26717
R3561 GNDA.n2327 GNDA.n289 4.26717
R3562 GNDA.n2327 GNDA.n2326 4.26717
R3563 GNDA.n2326 GNDA.n2325 4.26717
R3564 GNDA.n2325 GNDA.n297 4.26717
R3565 GNDA.n2319 GNDA.n297 4.26717
R3566 GNDA.n2319 GNDA.n2318 4.26717
R3567 GNDA.n2318 GNDA.n2317 4.26717
R3568 GNDA.n2275 GNDA.n344 4.26717
R3569 GNDA.n2281 GNDA.n344 4.26717
R3570 GNDA.n2282 GNDA.n2281 4.26717
R3571 GNDA.n2285 GNDA.n2282 4.26717
R3572 GNDA.n2285 GNDA.n340 4.26717
R3573 GNDA.n2291 GNDA.n340 4.26717
R3574 GNDA.n2292 GNDA.n2291 4.26717
R3575 GNDA.n2295 GNDA.n2292 4.26717
R3576 GNDA.n2295 GNDA.n338 4.26717
R3577 GNDA.n338 GNDA.n332 4.26717
R3578 GNDA.n2302 GNDA.n332 4.26717
R3579 GNDA.n2309 GNDA.n316 4.26717
R3580 GNDA.n620 GNDA.n316 4.26717
R3581 GNDA.n620 GNDA.n616 4.26717
R3582 GNDA.n628 GNDA.n616 4.26717
R3583 GNDA.n629 GNDA.n628 4.26717
R3584 GNDA.n632 GNDA.n629 4.26717
R3585 GNDA.n632 GNDA.n614 4.26717
R3586 GNDA.n639 GNDA.n614 4.26717
R3587 GNDA.n642 GNDA.n639 4.26717
R3588 GNDA.n642 GNDA.n612 4.26717
R3589 GNDA.n647 GNDA.n612 4.26717
R3590 GNDA.n1503 GNDA.n1430 4.26717
R3591 GNDA.n1498 GNDA.n1430 4.26717
R3592 GNDA.n1498 GNDA.n1497 4.26717
R3593 GNDA.n1497 GNDA.n1465 4.26717
R3594 GNDA.n1492 GNDA.n1465 4.26717
R3595 GNDA.n1492 GNDA.n1491 4.26717
R3596 GNDA.n1491 GNDA.n1490 4.26717
R3597 GNDA.n1490 GNDA.n1473 4.26717
R3598 GNDA.n1484 GNDA.n1473 4.26717
R3599 GNDA.n1484 GNDA.n1483 4.26717
R3600 GNDA.n1483 GNDA.n1482 4.26717
R3601 GNDA.n2397 GNDA.n89 4.26717
R3602 GNDA.n2397 GNDA.n91 4.26717
R3603 GNDA.n1514 GNDA.n91 4.26717
R3604 GNDA.n1519 GNDA.n1514 4.26717
R3605 GNDA.n1519 GNDA.n1511 4.26717
R3606 GNDA.n1525 GNDA.n1511 4.26717
R3607 GNDA.n1525 GNDA.n1509 4.26717
R3608 GNDA.n1531 GNDA.n1509 4.26717
R3609 GNDA.n1531 GNDA.n1507 4.26717
R3610 GNDA.n1537 GNDA.n1507 4.26717
R3611 GNDA.n1537 GNDA.n1505 4.26717
R3612 GNDA.n2017 GNDA.n2011 4.2505
R3613 GNDA.n2030 GNDA.n520 4.0005
R3614 GNDA.n2367 GNDA.n2366 3.93531
R3615 GNDA.n2339 GNDA.n2338 3.93531
R3616 GNDA.n2275 GNDA.n2245 3.93531
R3617 GNDA.n2310 GNDA.n2309 3.93531
R3618 GNDA.n1504 GNDA.n1503 3.93531
R3619 GNDA.n94 GNDA.n89 3.93531
R3620 GNDA.n2094 GNDA.n2093 3.90675
R3621 GNDA.n2056 GNDA.t434 3.88193
R3622 GNDA.n2055 GNDA.t283 3.88193
R3623 GNDA.n2054 GNDA.t317 3.88193
R3624 GNDA.n2053 GNDA.t310 3.88193
R3625 GNDA.n2089 GNDA.t308 3.88193
R3626 GNDA.n2088 GNDA.t212 3.88193
R3627 GNDA.n2087 GNDA.t455 3.88193
R3628 GNDA.n1258 GNDA.n1257 3.7893
R3629 GNDA.n1254 GNDA.n1148 3.7893
R3630 GNDA.n1253 GNDA.n1151 3.7893
R3631 GNDA.n1250 GNDA.n1249 3.7893
R3632 GNDA.n1175 GNDA.n1152 3.7893
R3633 GNDA.n1184 GNDA.n1183 3.7893
R3634 GNDA.n1187 GNDA.n1174 3.7893
R3635 GNDA.n1192 GNDA.n1188 3.7893
R3636 GNDA.n786 GNDA.n785 3.7893
R3637 GNDA.n782 GNDA.n651 3.7893
R3638 GNDA.n781 GNDA.n654 3.7893
R3639 GNDA.n660 GNDA.n659 3.7893
R3640 GNDA.n775 GNDA.n774 3.7893
R3641 GNDA.n689 GNDA.n688 3.7893
R3642 GNDA.n693 GNDA.n692 3.7893
R3643 GNDA.n716 GNDA.n679 3.7893
R3644 GNDA.n1137 GNDA.n1136 3.7893
R3645 GNDA.n1133 GNDA.n962 3.7893
R3646 GNDA.n1132 GNDA.n965 3.7893
R3647 GNDA.n1129 GNDA.n1128 3.7893
R3648 GNDA.n1054 GNDA.n966 3.7893
R3649 GNDA.n1063 GNDA.n1062 3.7893
R3650 GNDA.n1066 GNDA.n1053 3.7893
R3651 GNDA.n1071 GNDA.n1067 3.7893
R3652 GNDA.n2203 GNDA.n388 3.7893
R3653 GNDA.n2202 GNDA.n389 3.7893
R3654 GNDA.n2190 GNDA.n2189 3.7893
R3655 GNDA.n2196 GNDA.n2195 3.7893
R3656 GNDA.n2192 GNDA.n2191 3.7893
R3657 GNDA.n423 GNDA.n367 3.7893
R3658 GNDA.n426 GNDA.n424 3.7893
R3659 GNDA.n2139 GNDA.n2138 3.7893
R3660 GNDA.n1749 GNDA.n922 3.7893
R3661 GNDA.n1746 GNDA.n1745 3.7893
R3662 GNDA.n1662 GNDA.n923 3.7893
R3663 GNDA.n1667 GNDA.n1665 3.7893
R3664 GNDA.n1672 GNDA.n1668 3.7893
R3665 GNDA.n1679 GNDA.n1678 3.7893
R3666 GNDA.n1682 GNDA.n1661 3.7893
R3667 GNDA.n1687 GNDA.n1683 3.7893
R3668 GNDA.n1368 GNDA.n1266 3.7893
R3669 GNDA.n1376 GNDA.n1375 3.7893
R3670 GNDA.n1291 GNDA.n1267 3.7893
R3671 GNDA.n1295 GNDA.n1293 3.7893
R3672 GNDA.n1300 GNDA.n1296 3.7893
R3673 GNDA.n1307 GNDA.n1306 3.7893
R3674 GNDA.n1310 GNDA.n1290 3.7893
R3675 GNDA.n1315 GNDA.n1311 3.7893
R3676 GNDA.n1789 GNDA.n1787 3.7893
R3677 GNDA.n1788 GNDA.n542 3.7893
R3678 GNDA.n1795 GNDA.n1794 3.7893
R3679 GNDA.n572 GNDA.n543 3.7893
R3680 GNDA.n574 GNDA.n573 3.7893
R3681 GNDA.n596 GNDA.n568 3.7893
R3682 GNDA.n603 GNDA.n567 3.7893
R3683 GNDA.n605 GNDA.n604 3.7893
R3684 GNDA.n2430 GNDA.n22 3.7893
R3685 GNDA.n2429 GNDA.n23 3.7893
R3686 GNDA.n38 GNDA.n37 3.7893
R3687 GNDA.n44 GNDA.n43 3.7893
R3688 GNDA.n40 GNDA.n39 3.7893
R3689 GNDA.n208 GNDA.n1 3.7893
R3690 GNDA.n213 GNDA.n211 3.7893
R3691 GNDA.n218 GNDA.n214 3.7893
R3692 GNDA.n1651 GNDA.n1542 3.7893
R3693 GNDA.n1648 GNDA.n1647 3.7893
R3694 GNDA.n1564 GNDA.n1543 3.7893
R3695 GNDA.n1569 GNDA.n1567 3.7893
R3696 GNDA.n1574 GNDA.n1570 3.7893
R3697 GNDA.n1581 GNDA.n1580 3.7893
R3698 GNDA.n1584 GNDA.n1563 3.7893
R3699 GNDA.n1589 GNDA.n1585 3.7893
R3700 GNDA.n1180 GNDA 3.7381
R3701 GNDA.n687 GNDA 3.7381
R3702 GNDA.n1059 GNDA 3.7381
R3703 GNDA GNDA.n2208 3.7381
R3704 GNDA.n1675 GNDA 3.7381
R3705 GNDA.n1303 GNDA 3.7381
R3706 GNDA.n597 GNDA 3.7381
R3707 GNDA GNDA.n2435 3.7381
R3708 GNDA.n1577 GNDA 3.7381
R3709 GNDA.t192 GNDA.t386 3.66107
R3710 GNDA.t376 GNDA.t193 3.66107
R3711 GNDA.t262 GNDA.n525 3.66107
R3712 GNDA.n2026 GNDA.t446 3.66107
R3713 GNDA.n2090 GNDA.t207 3.66107
R3714 GNDA.t443 GNDA.t264 3.66107
R3715 GNDA.t266 GNDA.t437 3.66107
R3716 GNDA.n2012 GNDA.n519 3.65764
R3717 GNDA.n2013 GNDA.n519 3.65764
R3718 GNDA.n2025 GNDA.n526 3.65764
R3719 GNDA.n2025 GNDA.n2024 3.65764
R3720 GNDA.n527 GNDA.n515 3.53175
R3721 GNDA.n1972 GNDA.n1837 3.50448
R3722 GNDA.n1901 GNDA.n1895 3.47871
R3723 GNDA.n1920 GNDA.n1892 3.47871
R3724 GNDA.n1977 GNDA.n1833 3.43627
R3725 GNDA.n1987 GNDA.t29 3.42907
R3726 GNDA.n1987 GNDA.t298 3.42907
R3727 GNDA.n1985 GNDA.t219 3.42907
R3728 GNDA.n1985 GNDA.t337 3.42907
R3729 GNDA.n2111 GNDA.t291 3.42907
R3730 GNDA.n2111 GNDA.t224 3.42907
R3731 GNDA.n2109 GNDA.t61 3.42907
R3732 GNDA.n2109 GNDA.t322 3.42907
R3733 GNDA.n1971 GNDA.n1970 3.4105
R3734 GNDA.n1969 GNDA.n1836 3.4105
R3735 GNDA.n1975 GNDA.n1835 3.4105
R3736 GNDA.n1976 GNDA.n1834 3.4105
R3737 GNDA.n1899 GNDA.n1898 3.4105
R3738 GNDA.n1907 GNDA.n1906 3.4105
R3739 GNDA.n1905 GNDA.n1904 3.4105
R3740 GNDA.n1903 GNDA.n1902 3.4105
R3741 GNDA.n1915 GNDA.n1914 3.4105
R3742 GNDA.n1918 GNDA.n1917 3.4105
R3743 GNDA.n1926 GNDA.n1925 3.4105
R3744 GNDA.n1924 GNDA.n1923 3.4105
R3745 GNDA.n1922 GNDA.n1921 3.4105
R3746 GNDA.n1932 GNDA.n1931 3.4105
R3747 GNDA.n1933 GNDA.n1892 3.4105
R3748 GNDA.n1933 GNDA.n1932 3.4105
R3749 GNDA.n1916 GNDA.n1895 3.4105
R3750 GNDA.n1916 GNDA.n1915 3.4105
R3751 GNDA.n1934 GNDA.n1887 3.4105
R3752 GNDA.n1887 GNDA.n1884 3.4105
R3753 GNDA.n1939 GNDA.n1887 3.4105
R3754 GNDA.n1938 GNDA.n1937 3.4105
R3755 GNDA.n1939 GNDA.n1938 3.4105
R3756 GNDA.n1937 GNDA.n1885 3.4105
R3757 GNDA.n1885 GNDA.n1881 3.4105
R3758 GNDA.n1885 GNDA.n1883 3.4105
R3759 GNDA.n1885 GNDA.n1880 3.4105
R3760 GNDA.n1885 GNDA.n1884 3.4105
R3761 GNDA.n1939 GNDA.n1885 3.4105
R3762 GNDA.n1940 GNDA.n1881 3.4105
R3763 GNDA.n1940 GNDA.n1883 3.4105
R3764 GNDA.n1940 GNDA.n1880 3.4105
R3765 GNDA.n1940 GNDA.n1884 3.4105
R3766 GNDA.n1940 GNDA.n1939 3.4105
R3767 GNDA.n1966 GNDA.n1949 3.4105
R3768 GNDA.n1962 GNDA.n1949 3.4105
R3769 GNDA.n1964 GNDA.n1949 3.4105
R3770 GNDA.n1963 GNDA.n1962 3.4105
R3771 GNDA.n1964 GNDA.n1963 3.4105
R3772 GNDA.n1966 GNDA.n1839 3.4105
R3773 GNDA.n1954 GNDA.n1839 3.4105
R3774 GNDA.n1952 GNDA.n1839 3.4105
R3775 GNDA.n1955 GNDA.n1839 3.4105
R3776 GNDA.n1962 GNDA.n1839 3.4105
R3777 GNDA.n1964 GNDA.n1839 3.4105
R3778 GNDA.n1966 GNDA.n1965 3.4105
R3779 GNDA.n1965 GNDA.n1954 3.4105
R3780 GNDA.n1965 GNDA.n1952 3.4105
R3781 GNDA.n1965 GNDA.n1955 3.4105
R3782 GNDA.n1965 GNDA.n1964 3.4105
R3783 GNDA.n1943 GNDA.n1853 3.4105
R3784 GNDA.n1946 GNDA.n1853 3.4105
R3785 GNDA.n1946 GNDA.n1841 3.4105
R3786 GNDA.n1946 GNDA.n1945 3.4105
R3787 GNDA.n1947 GNDA.n1946 3.4105
R3788 GNDA.n1853 GNDA.n1845 3.4105
R3789 GNDA.n1845 GNDA.n1843 3.4105
R3790 GNDA.n1945 GNDA.n1845 3.4105
R3791 GNDA.n1947 GNDA.n1845 3.4105
R3792 GNDA.n1948 GNDA.n1841 3.4105
R3793 GNDA.n1948 GNDA.n1843 3.4105
R3794 GNDA.n1948 GNDA.n1947 3.4105
R3795 GNDA.n524 GNDA.n523 3.39217
R3796 GNDA.n2092 GNDA.n2091 3.39217
R3797 GNDA.n2032 GNDA.n2031 3.39217
R3798 GNDA.n2028 GNDA.n2027 3.39217
R3799 GNDA.n2014 GNDA.n2012 3.13621
R3800 GNDA.n2014 GNDA.n2013 3.13621
R3801 GNDA.n2023 GNDA.n526 3.13621
R3802 GNDA.n2024 GNDA.n2023 3.13621
R3803 GNDA.n1798 GNDA.n1797 3.01902
R3804 GNDA.n2155 GNDA.n409 3.01902
R3805 GNDA.n2200 GNDA.t45 3.01902
R3806 GNDA.n419 GNDA.t275 3.01902
R3807 GNDA.t366 GNDA.t429 2.9898
R3808 GNDA.n2175 GNDA.n2174 2.86505
R3809 GNDA.n2176 GNDA.n2175 2.86505
R3810 GNDA.n2180 GNDA.n2178 2.86505
R3811 GNDA.n2183 GNDA.n2178 2.86505
R3812 GNDA.n2179 GNDA.n2176 2.86505
R3813 GNDA.n2183 GNDA.n2182 2.86505
R3814 GNDA.n2185 GNDA.n2174 2.86505
R3815 GNDA.n2180 GNDA.n2179 2.86505
R3816 GNDA.n583 GNDA.n581 2.86505
R3817 GNDA.n585 GNDA.n583 2.86505
R3818 GNDA.n585 GNDA.n584 2.86505
R3819 GNDA.n581 GNDA.n579 2.86505
R3820 GNDA.n527 GNDA.n516 2.813
R3821 GNDA.n1147 GNDA.n1146 2.6629
R3822 GNDA.n1172 GNDA.n305 2.6629
R3823 GNDA.n788 GNDA.n787 2.6629
R3824 GNDA.n681 GNDA.n333 2.6629
R3825 GNDA.n961 GNDA.n960 2.6629
R3826 GNDA.n433 GNDA.n432 2.6629
R3827 GNDA.n1751 GNDA.n1750 2.6629
R3828 GNDA.n1659 GNDA.n942 2.6629
R3829 GNDA.n1369 GNDA.n952 2.6629
R3830 GNDA.n1288 GNDA.n312 2.6629
R3831 GNDA.n1780 GNDA.n850 2.6629
R3832 GNDA.n796 GNDA.n563 2.6629
R3833 GNDA.n274 GNDA.n273 2.6629
R3834 GNDA.n1653 GNDA.n1652 2.6629
R3835 GNDA.n2343 GNDA.n275 2.6629
R3836 GNDA.n1146 GNDA.n312 2.4581
R3837 GNDA.n1173 GNDA.n1172 2.4581
R3838 GNDA.n788 GNDA.n563 2.4581
R3839 GNDA.n681 GNDA.n678 2.4581
R3840 GNDA.n960 GNDA.n305 2.4581
R3841 GNDA.n1052 GNDA.n1051 2.4581
R3842 GNDA.n432 GNDA.n333 2.4581
R3843 GNDA.n2134 GNDA.n2133 2.4581
R3844 GNDA.n1660 GNDA.n1659 2.4581
R3845 GNDA.n1289 GNDA.n1288 2.4581
R3846 GNDA.n797 GNDA.n796 2.4581
R3847 GNDA.n2343 GNDA.n274 2.4581
R3848 GNDA.n207 GNDA.n206 2.4581
R3849 GNDA.n1653 GNDA.n942 2.4581
R3850 GNDA.n1562 GNDA.n275 2.4581
R3851 GNDA.n1973 GNDA.n1972 2.39683
R3852 GNDA.n1901 GNDA.n1900 2.39683
R3853 GNDA.n1920 GNDA.n1919 2.39683
R3854 GNDA.n2172 GNDA.n2171 2.26187
R3855 GNDA.n2030 GNDA.n2029 2.2505
R3856 GNDA.n2170 GNDA.n2169 2.24063
R3857 GNDA.n2168 GNDA.n395 2.24063
R3858 GNDA.n2166 GNDA.n2165 2.24063
R3859 GNDA.n403 GNDA.n401 2.24063
R3860 GNDA.n2173 GNDA.n2172 2.24063
R3861 GNDA.n2167 GNDA.n399 2.24063
R3862 GNDA.n703 GNDA.n402 2.22018
R3863 GNDA.n2162 GNDA.n404 2.22018
R3864 GNDA.t366 GNDA.t41 2.20362
R3865 GNDA.n2059 GNDA.n2058 2.19633
R3866 GNDA.n2344 GNDA.n2343 2.18124
R3867 GNDA.n2317 GNDA.n305 2.18124
R3868 GNDA.n2302 GNDA.n333 2.18124
R3869 GNDA.n647 GNDA.n563 2.18124
R3870 GNDA.n1482 GNDA.n312 2.18124
R3871 GNDA.n1505 GNDA.n942 2.18124
R3872 GNDA.n1191 GNDA.n1173 2.1509
R3873 GNDA.n715 GNDA.n678 2.1509
R3874 GNDA.n1070 GNDA.n1052 2.1509
R3875 GNDA.n2134 GNDA.n427 2.1509
R3876 GNDA.n1686 GNDA.n1660 2.1509
R3877 GNDA.n1314 GNDA.n1289 2.1509
R3878 GNDA.n797 GNDA.n562 2.1509
R3879 GNDA.n217 GNDA.n207 2.1509
R3880 GNDA.n1588 GNDA.n1562 2.1509
R3881 GNDA.n1652 GNDA.n1541 2.13383
R3882 GNDA.n273 GNDA.n272 2.13383
R3883 GNDA.n1231 GNDA.n1147 2.13383
R3884 GNDA.n787 GNDA.n650 2.13383
R3885 GNDA.n1110 GNDA.n961 2.13383
R3886 GNDA.n434 GNDA.n433 2.13383
R3887 GNDA.n1750 GNDA.n921 2.13383
R3888 GNDA.n1370 GNDA.n1369 2.13383
R3889 GNDA.n850 GNDA.n849 2.13383
R3890 GNDA.n1983 GNDA.n1982 2.09414
R3891 GNDA.n2115 GNDA.n2114 2.09414
R3892 GNDA.n2107 GNDA.n2106 2.09414
R3893 GNDA.n1991 GNDA.n1990 2.09414
R3894 GNDA.n2343 GNDA.n2342 2.08643
R3895 GNDA.n307 GNDA.n305 2.08643
R3896 GNDA.n334 GNDA.n333 2.08643
R3897 GNDA.n790 GNDA.n563 2.08643
R3898 GNDA.n2311 GNDA.n312 2.08643
R3899 GNDA.n1656 GNDA.n942 2.08643
R3900 GNDA.n1258 GNDA.n1147 1.9461
R3901 GNDA.n787 GNDA.n786 1.9461
R3902 GNDA.n1137 GNDA.n961 1.9461
R3903 GNDA.n433 GNDA.n388 1.9461
R3904 GNDA.n1750 GNDA.n1749 1.9461
R3905 GNDA.n1369 GNDA.n1368 1.9461
R3906 GNDA.n1787 GNDA.n850 1.9461
R3907 GNDA.n273 GNDA.n22 1.9461
R3908 GNDA.n1652 GNDA.n1651 1.9461
R3909 GNDA.n2093 GNDA.n514 1.938
R3910 GNDA.n1994 GNDA.n1993 1.93383
R3911 GNDA.n1997 GNDA.n1996 1.93383
R3912 GNDA.n2119 GNDA.n2118 1.93383
R3913 GNDA.n2122 GNDA.n2121 1.93383
R3914 GNDA.n2085 GNDA.n2084 1.91062
R3915 GNDA.n1912 GNDA.n1911 1.90675
R3916 GNDA.n2020 GNDA.n2017 1.7505
R3917 GNDA.t93 GNDA.n62 1.74476
R3918 GNDA.n1889 GNDA.n1888 1.70468
R3919 GNDA.n1888 GNDA.n1879 1.70468
R3920 GNDA.n1957 GNDA.n1956 1.70468
R3921 GNDA.n1956 GNDA.n1950 1.70468
R3922 GNDA.n1849 GNDA.n1848 1.70468
R3923 GNDA.n1854 GNDA.n1840 1.70468
R3924 GNDA.n1935 GNDA.n1934 1.70453
R3925 GNDA.n1960 GNDA.n1959 1.70453
R3926 GNDA.n1851 GNDA.n1850 1.70453
R3927 GNDA.n1936 GNDA.n1887 1.70321
R3928 GNDA.n1940 GNDA.n1882 1.70321
R3929 GNDA.n1953 GNDA.n1949 1.70321
R3930 GNDA.n1963 GNDA.n1838 1.70321
R3931 GNDA.n1943 GNDA.n1846 1.70321
R3932 GNDA.n1847 GNDA.n1845 1.70321
R3933 GNDA.n1948 GNDA.n1842 1.70321
R3934 GNDA.n1948 GNDA.n1844 1.70321
R3935 GNDA.n1887 GNDA.n1886 1.70307
R3936 GNDA.n1938 GNDA.n1891 1.70307
R3937 GNDA.n1938 GNDA.n1890 1.70307
R3938 GNDA.n1958 GNDA.n1949 1.70307
R3939 GNDA.n1963 GNDA.n1961 1.70307
R3940 GNDA.n1965 GNDA.n1951 1.70307
R3941 GNDA.n1943 GNDA.n1942 1.70307
R3942 GNDA.n1944 GNDA.n1943 1.70307
R3943 GNDA.n1946 GNDA.n1852 1.70307
R3944 GNDA.n1967 GNDA.n1833 1.69337
R3945 GNDA.n1967 GNDA.n1837 1.69337
R3946 GNDA.n1933 GNDA.n1894 1.6924
R3947 GNDA.n1933 GNDA.n1893 1.6924
R3948 GNDA.n1916 GNDA.n1897 1.6924
R3949 GNDA.n1916 GNDA.n1896 1.6924
R3950 GNDA.n1968 GNDA.n1967 1.6924
R3951 GNDA.n1984 GNDA.n1980 1.563
R3952 GNDA.n1041 GNDA.n985 1.47392
R3953 GNDA.n497 GNDA.n485 1.47392
R3954 GNDA.n1757 GNDA.n1754 1.47392
R3955 GNDA.n1384 GNDA.n1383 1.47392
R3956 GNDA.n1779 GNDA.n852 1.47392
R3957 GNDA.n199 GNDA.n134 1.47392
R3958 GNDA.n1995 GNDA.n528 1.3755
R3959 GNDA.n2110 GNDA.n2108 1.1255
R3960 GNDA.n2112 GNDA.n2110 1.1255
R3961 GNDA.n2113 GNDA.n2112 1.1255
R3962 GNDA.n2113 GNDA.n2094 1.1255
R3963 GNDA.n1986 GNDA.n1984 1.1255
R3964 GNDA.n1988 GNDA.n1986 1.1255
R3965 GNDA.n1989 GNDA.n1988 1.1255
R3966 GNDA.n2011 GNDA.n528 1.0005
R3967 GNDA.n1257 GNDA.n1148 0.8197
R3968 GNDA.n1254 GNDA.n1253 0.8197
R3969 GNDA.n1250 GNDA.n1151 0.8197
R3970 GNDA.n1249 GNDA.n1152 0.8197
R3971 GNDA.n1183 GNDA.n1180 0.8197
R3972 GNDA.n1184 GNDA.n1174 0.8197
R3973 GNDA.n1188 GNDA.n1187 0.8197
R3974 GNDA.n1192 GNDA.n1191 0.8197
R3975 GNDA.n785 GNDA.n651 0.8197
R3976 GNDA.n782 GNDA.n781 0.8197
R3977 GNDA.n659 GNDA.n654 0.8197
R3978 GNDA.n775 GNDA.n660 0.8197
R3979 GNDA.n688 GNDA.n687 0.8197
R3980 GNDA.n693 GNDA.n689 0.8197
R3981 GNDA.n692 GNDA.n679 0.8197
R3982 GNDA.n716 GNDA.n715 0.8197
R3983 GNDA.n1136 GNDA.n962 0.8197
R3984 GNDA.n1133 GNDA.n1132 0.8197
R3985 GNDA.n1129 GNDA.n965 0.8197
R3986 GNDA.n1128 GNDA.n966 0.8197
R3987 GNDA.n1062 GNDA.n1059 0.8197
R3988 GNDA.n1063 GNDA.n1053 0.8197
R3989 GNDA.n1067 GNDA.n1066 0.8197
R3990 GNDA.n1071 GNDA.n1070 0.8197
R3991 GNDA.n2203 GNDA.n2202 0.8197
R3992 GNDA.n2189 GNDA.n389 0.8197
R3993 GNDA.n2196 GNDA.n2190 0.8197
R3994 GNDA.n2195 GNDA.n2192 0.8197
R3995 GNDA.n2208 GNDA.n367 0.8197
R3996 GNDA.n424 GNDA.n423 0.8197
R3997 GNDA.n2139 GNDA.n426 0.8197
R3998 GNDA.n2138 GNDA.n427 0.8197
R3999 GNDA.n1746 GNDA.n922 0.8197
R4000 GNDA.n1745 GNDA.n923 0.8197
R4001 GNDA.n1665 GNDA.n1662 0.8197
R4002 GNDA.n1668 GNDA.n1667 0.8197
R4003 GNDA.n1678 GNDA.n1675 0.8197
R4004 GNDA.n1679 GNDA.n1661 0.8197
R4005 GNDA.n1683 GNDA.n1682 0.8197
R4006 GNDA.n1687 GNDA.n1686 0.8197
R4007 GNDA.n1376 GNDA.n1266 0.8197
R4008 GNDA.n1375 GNDA.n1267 0.8197
R4009 GNDA.n1293 GNDA.n1291 0.8197
R4010 GNDA.n1296 GNDA.n1295 0.8197
R4011 GNDA.n1306 GNDA.n1303 0.8197
R4012 GNDA.n1307 GNDA.n1290 0.8197
R4013 GNDA.n1311 GNDA.n1310 0.8197
R4014 GNDA.n1315 GNDA.n1314 0.8197
R4015 GNDA.n1789 GNDA.n1788 0.8197
R4016 GNDA.n1795 GNDA.n542 0.8197
R4017 GNDA.n1794 GNDA.n543 0.8197
R4018 GNDA.n573 GNDA.n572 0.8197
R4019 GNDA.n597 GNDA.n596 0.8197
R4020 GNDA.n568 GNDA.n567 0.8197
R4021 GNDA.n605 GNDA.n603 0.8197
R4022 GNDA.n604 GNDA.n562 0.8197
R4023 GNDA.n2430 GNDA.n2429 0.8197
R4024 GNDA.n37 GNDA.n23 0.8197
R4025 GNDA.n44 GNDA.n38 0.8197
R4026 GNDA.n43 GNDA.n40 0.8197
R4027 GNDA.n2435 GNDA.n1 0.8197
R4028 GNDA.n211 GNDA.n208 0.8197
R4029 GNDA.n214 GNDA.n213 0.8197
R4030 GNDA.n218 GNDA.n217 0.8197
R4031 GNDA.n1648 GNDA.n1542 0.8197
R4032 GNDA.n1647 GNDA.n1543 0.8197
R4033 GNDA.n1567 GNDA.n1564 0.8197
R4034 GNDA.n1570 GNDA.n1569 0.8197
R4035 GNDA.n1580 GNDA.n1577 0.8197
R4036 GNDA.n1581 GNDA.n1563 0.8197
R4037 GNDA.n1585 GNDA.n1584 0.8197
R4038 GNDA.n1589 GNDA.n1588 0.8197
R4039 GNDA.n2168 GNDA.n2167 0.745292
R4040 GNDA.n1967 GNDA.n1966 0.7384
R4041 GNDA.n1979 GNDA.n514 0.6255
R4042 GNDA GNDA.n1175 0.5637
R4043 GNDA.n774 GNDA 0.5637
R4044 GNDA GNDA.n1054 0.5637
R4045 GNDA.n2191 GNDA 0.5637
R4046 GNDA.n1672 GNDA 0.5637
R4047 GNDA.n1300 GNDA 0.5637
R4048 GNDA GNDA.n574 0.5637
R4049 GNDA.n39 GNDA 0.5637
R4050 GNDA.n1574 GNDA 0.5637
R4051 GNDA.n2042 GNDA.n2040 0.563
R4052 GNDA.n2044 GNDA.n2042 0.563
R4053 GNDA.n2046 GNDA.n2044 0.563
R4054 GNDA.n2048 GNDA.n2046 0.563
R4055 GNDA.n2049 GNDA.n2048 0.563
R4056 GNDA.n2062 GNDA.n2060 0.563
R4057 GNDA.n2064 GNDA.n2062 0.563
R4058 GNDA.n2066 GNDA.n2064 0.563
R4059 GNDA.n2068 GNDA.n2066 0.563
R4060 GNDA.n2070 GNDA.n2068 0.563
R4061 GNDA.n2072 GNDA.n2070 0.563
R4062 GNDA.n2074 GNDA.n2072 0.563
R4063 GNDA.n2076 GNDA.n2074 0.563
R4064 GNDA.n2078 GNDA.n2076 0.563
R4065 GNDA.n2080 GNDA.n2078 0.563
R4066 GNDA.n2082 GNDA.n2080 0.563
R4067 GNDA.n2099 GNDA.n2097 0.563
R4068 GNDA.n2101 GNDA.n2099 0.563
R4069 GNDA.n2103 GNDA.n2101 0.563
R4070 GNDA.n2105 GNDA.n2103 0.563
R4071 GNDA.n1825 GNDA.n1823 0.563
R4072 GNDA.n1827 GNDA.n1825 0.563
R4073 GNDA.n1829 GNDA.n1827 0.563
R4074 GNDA.n1831 GNDA.n1829 0.563
R4075 GNDA.n1776 GNDA.n62 0.526383
R4076 GNDA.n1933 GNDA.n1916 0.513975
R4077 GNDA.n1934 GNDA.n1933 0.476375
R4078 GNDA.n1943 GNDA.n1941 0.466681
R4079 GNDA.n1947 GNDA 0.422325
R4080 GNDA.n1949 GNDA.n1948 0.404112
R4081 GNDA.n1178 GNDA 0.2565
R4082 GNDA.n686 GNDA 0.2565
R4083 GNDA.n1057 GNDA 0.2565
R4084 GNDA.n2209 GNDA 0.2565
R4085 GNDA GNDA.n1671 0.2565
R4086 GNDA GNDA.n1299 0.2565
R4087 GNDA.n575 GNDA 0.2565
R4088 GNDA GNDA.n0 0.2565
R4089 GNDA GNDA.n1573 0.2565
R4090 GNDA.n2083 GNDA.n2082 0.21925
R4091 GNDA.n2016 GNDA.n2014 0.208833
R4092 GNDA.n2023 GNDA.n2022 0.208833
R4093 GNDA.n2163 GNDA.n2162 0.188
R4094 GNDA.n2165 GNDA.n402 0.188
R4095 GNDA.t137 GNDA.t545 0.1603
R4096 GNDA.t109 GNDA.t137 0.1603
R4097 GNDA.t473 GNDA.t109 0.1603
R4098 GNDA.t355 GNDA.t473 0.1603
R4099 GNDA.t508 GNDA.t464 0.1603
R4100 GNDA.t55 GNDA.t508 0.1603
R4101 GNDA.t535 GNDA.t55 0.1603
R4102 GNDA.t474 GNDA.t535 0.1603
R4103 GNDA.t253 GNDA.t561 0.1603
R4104 GNDA.t469 GNDA.t253 0.1603
R4105 GNDA.t71 GNDA.t469 0.1603
R4106 GNDA.t512 GNDA.t71 0.1603
R4107 GNDA.t116 GNDA.t332 0.1603
R4108 GNDA.t499 GNDA.t116 0.1603
R4109 GNDA.t481 GNDA.t499 0.1603
R4110 GNDA.t205 GNDA.t481 0.1603
R4111 GNDA.t307 GNDA.t507 0.1603
R4112 GNDA.t138 GNDA.t307 0.1603
R4113 GNDA.t88 GNDA.t138 0.1603
R4114 GNDA.t101 GNDA.t88 0.1603
R4115 GNDA.t18 GNDA.t353 0.1603
R4116 GNDA.t34 GNDA.t18 0.1603
R4117 GNDA.t541 GNDA.t34 0.1603
R4118 GNDA.t483 GNDA.t541 0.1603
R4119 GNDA.t20 GNDA.t287 0.1603
R4120 GNDA.t503 GNDA.t20 0.1603
R4121 GNDA.t293 GNDA.t503 0.1603
R4122 GNDA.t180 GNDA.t293 0.1603
R4123 GNDA.t295 GNDA.t279 0.1603
R4124 GNDA.t68 GNDA.t295 0.1603
R4125 GNDA.t345 GNDA.t68 0.1603
R4126 GNDA.t83 GNDA.t345 0.1603
R4127 GNDA.t107 GNDA.t158 0.1603
R4128 GNDA.t350 GNDA.t107 0.1603
R4129 GNDA.t519 GNDA.t350 0.1603
R4130 GNDA.t36 GNDA.t519 0.1603
R4131 GNDA.t472 GNDA.t534 0.1603
R4132 GNDA.t354 GNDA.t472 0.1603
R4133 GNDA.t505 GNDA.t354 0.1603
R4134 GNDA.t24 GNDA.t505 0.1603
R4135 GNDA.t548 GNDA.t524 0.1603
R4136 GNDA.t159 GNDA.t548 0.1603
R4137 GNDA.t120 GNDA.t159 0.1603
R4138 GNDA.t202 GNDA.t120 0.1603
R4139 GNDA.t131 GNDA.t482 0.1603
R4140 GNDA.t564 GNDA.t131 0.1603
R4141 GNDA.t573 GNDA.t564 0.1603
R4142 GNDA.t359 GNDA.t573 0.1603
R4143 GNDA.t108 GNDA.t476 0.1603
R4144 GNDA.t296 GNDA.t108 0.1603
R4145 GNDA.t280 GNDA.t296 0.1603
R4146 GNDA.t528 GNDA.t280 0.1603
R4147 GNDA.t484 GNDA.t542 0.1603
R4148 GNDA.t204 GNDA.t484 0.1603
R4149 GNDA.t516 GNDA.t204 0.1603
R4150 GNDA.t100 GNDA.t516 0.1603
R4151 GNDA.t496 GNDA.t539 0.1603
R4152 GNDA.t160 GNDA.t496 0.1603
R4153 GNDA.t530 GNDA.t160 0.1603
R4154 GNDA.t556 GNDA.t530 0.1603
R4155 GNDA.t80 GNDA.t148 0.1603
R4156 GNDA.t489 GNDA.t80 0.1603
R4157 GNDA.t38 GNDA.t489 0.1603
R4158 GNDA.t143 GNDA.t38 0.1603
R4159 GNDA.t333 GNDA.t558 0.1603
R4160 GNDA.t536 GNDA.t333 0.1603
R4161 GNDA.t572 GNDA.t536 0.1603
R4162 GNDA.t177 GNDA.t572 0.1603
R4163 GNDA.t490 GNDA.t86 0.1603
R4164 GNDA.t135 GNDA.t490 0.1603
R4165 GNDA.t522 GNDA.t135 0.1603
R4166 GNDA.t286 GNDA.t522 0.1603
R4167 GNDA.t33 GNDA.t79 0.1603
R4168 GNDA.t485 GNDA.t33 0.1603
R4169 GNDA.t543 GNDA.t485 0.1603
R4170 GNDA.t190 GNDA.t543 0.1603
R4171 GNDA.t361 GNDA.t575 0.1603
R4172 GNDA.t183 GNDA.t361 0.1603
R4173 GNDA.t526 GNDA.t183 0.1603
R4174 GNDA.t114 GNDA.t526 0.1603
R4175 GNDA.t129 GNDA.t51 0.1603
R4176 GNDA.t81 GNDA.t129 0.1603
R4177 GNDA.t149 GNDA.t81 0.1603
R4178 GNDA.t227 GNDA.t149 0.1603
R4179 GNDA.t563 GNDA.t514 0.1603
R4180 GNDA.t90 GNDA.t563 0.1603
R4181 GNDA.t568 GNDA.t90 0.1603
R4182 GNDA.t527 GNDA.t568 0.1603
R4183 GNDA.t358 GNDA.t510 0.1603
R4184 GNDA.t343 GNDA.t358 0.1603
R4185 GNDA.t500 GNDA.t343 0.1603
R4186 GNDA.t117 GNDA.t500 0.1603
R4187 GNDA.t502 GNDA.t466 0.1603
R4188 GNDA.t56 GNDA.t502 0.1603
R4189 GNDA.t537 GNDA.t56 0.1603
R4190 GNDA.t475 GNDA.t537 0.1603
R4191 GNDA.t254 GNDA.t562 0.1603
R4192 GNDA.t470 GNDA.t254 0.1603
R4193 GNDA.t72 GNDA.t470 0.1603
R4194 GNDA.t513 GNDA.t72 0.1603
R4195 GNDA.t349 GNDA.t523 0.1603
R4196 GNDA.t334 GNDA.t349 0.1603
R4197 GNDA.t559 GNDA.t334 0.1603
R4198 GNDA.t538 GNDA.t559 0.1603
R4199 GNDA.t4 GNDA.t181 0.1603
R4200 GNDA.t574 GNDA.t4 0.1603
R4201 GNDA.t511 GNDA.t574 0.1603
R4202 GNDA.t247 GNDA.t511 0.1603
R4203 GNDA.t517 GNDA.t186 0.1603
R4204 GNDA.t99 GNDA.t517 0.1603
R4205 GNDA.t134 GNDA.t99 0.1603
R4206 GNDA.t342 GNDA.t134 0.1603
R4207 GNDA.t478 GNDA.t168 0.1603
R4208 GNDA.t506 GNDA.t478 0.1603
R4209 GNDA.t209 GNDA.t506 0.1603
R4210 GNDA.t19 GNDA.t209 0.1603
R4211 GNDA.t145 GNDA.t565 0.1603
R4212 GNDA.t142 GNDA.t145 0.1603
R4213 GNDA.t182 GNDA.t142 0.1603
R4214 GNDA.t176 GNDA.t182 0.1603
R4215 GNDA.t75 GNDA.t582 0.1603
R4216 GNDA.t169 GNDA.t75 0.1603
R4217 GNDA.t69 GNDA.t169 0.1603
R4218 GNDA.t351 GNDA.t69 0.1603
R4219 GNDA.t521 GNDA.t122 0.1603
R4220 GNDA.t468 GNDA.t521 0.1603
R4221 GNDA.t243 GNDA.t468 0.1603
R4222 GNDA.t189 GNDA.t243 0.1603
R4223 GNDA.t488 GNDA.t37 0.1603
R4224 GNDA.t518 GNDA.t488 0.1603
R4225 GNDA.t187 GNDA.t518 0.1603
R4226 GNDA.t581 GNDA.t187 0.1603
R4227 GNDA.t525 GNDA.t21 0.1603
R4228 GNDA.t113 GNDA.t525 0.1603
R4229 GNDA.t495 GNDA.t113 0.1603
R4230 GNDA.t226 GNDA.t495 0.1603
R4231 GNDA.t82 GNDA.t203 0.1603
R4232 GNDA.t146 GNDA.t82 0.1603
R4233 GNDA.t566 GNDA.t146 0.1603
R4234 GNDA.t132 GNDA.t566 0.1603
R4235 GNDA.t567 GNDA.t136 0.1603
R4236 GNDA.t531 GNDA.t567 0.1603
R4237 GNDA.t49 GNDA.t531 0.1603
R4238 GNDA.t115 GNDA.t49 0.1603
R4239 GNDA.t23 GNDA.t104 0.1603
R4240 GNDA.t252 GNDA.t23 0.1603
R4241 GNDA.t206 GNDA.t252 0.1603
R4242 GNDA.t480 GNDA.t206 0.1603
R4243 GNDA.t533 GNDA.t341 0.1603
R4244 GNDA.t479 GNDA.t533 0.1603
R4245 GNDA.t170 GNDA.t479 0.1603
R4246 GNDA.t509 GNDA.t170 0.1603
R4247 GNDA.t89 GNDA.t557 0.1603
R4248 GNDA.t306 GNDA.t89 0.1603
R4249 GNDA.t22 GNDA.t306 0.1603
R4250 GNDA.t103 GNDA.t22 0.1603
R4251 GNDA.t560 GNDA.t110 0.1603
R4252 GNDA.t76 GNDA.t560 0.1603
R4253 GNDA.t128 GNDA.t76 0.1603
R4254 GNDA.t248 GNDA.t128 0.1603
R4255 GNDA.t294 GNDA.t105 0.1603
R4256 GNDA.t569 GNDA.t294 0.1603
R4257 GNDA.t102 GNDA.t569 0.1603
R4258 GNDA.t492 GNDA.t102 0.1603
R4259 GNDA.t6 GNDA.t57 0.1603
R4260 GNDA.t188 GNDA.t6 0.1603
R4261 GNDA.t357 GNDA.t188 0.1603
R4262 GNDA.t580 GNDA.t357 0.1603
R4263 GNDA.t141 GNDA.t547 0.1603
R4264 GNDA.t106 GNDA.t141 0.1603
R4265 GNDA.t184 GNDA.t106 0.1603
R4266 GNDA.t471 GNDA.t184 0.1603
R4267 GNDA.t344 GNDA.t225 0.1603
R4268 GNDA.t84 GNDA.t344 0.1603
R4269 GNDA.t340 GNDA.t84 0.1603
R4270 GNDA.t58 GNDA.t340 0.1603
R4271 GNDA.t467 GNDA.t5 0.1603
R4272 GNDA.t570 GNDA.t467 0.1603
R4273 GNDA.t175 GNDA.t570 0.1603
R4274 GNDA.t139 GNDA.t175 0.1603
R4275 GNDA.t504 GNDA.t35 0.1603
R4276 GNDA.t25 GNDA.t504 0.1603
R4277 GNDA.t3 GNDA.t25 0.1603
R4278 GNDA.t201 GNDA.t3 0.1603
R4279 GNDA.t112 GNDA.t494 0.1603
R4280 GNDA.t242 GNDA.t112 0.1603
R4281 GNDA.t32 GNDA.t242 0.1603
R4282 GNDA.t544 GNDA.t32 0.1603
R4283 GNDA.t87 GNDA.t50 0.1603
R4284 GNDA.t491 GNDA.t87 0.1603
R4285 GNDA.t147 GNDA.t491 0.1603
R4286 GNDA.t360 GNDA.t147 0.1603
R4287 GNDA.t520 GNDA.n1855 0.159278
R4288 GNDA.t185 GNDA.n1856 0.159278
R4289 GNDA.t515 GNDA.n1857 0.159278
R4290 GNDA.t70 GNDA.n1858 0.159278
R4291 GNDA.t501 GNDA.n1859 0.159278
R4292 GNDA.t150 GNDA.n1860 0.159278
R4293 GNDA.t74 GNDA.n1861 0.159278
R4294 GNDA.t571 GNDA.n1862 0.159278
R4295 GNDA.t529 GNDA.n1863 0.159278
R4296 GNDA.t477 GNDA.n1864 0.159278
R4297 GNDA.t356 GNDA.n1865 0.159278
R4298 GNDA.t161 GNDA.n1866 0.159278
R4299 GNDA.t352 GNDA.n1867 0.159278
R4300 GNDA.t48 GNDA.n1868 0.159278
R4301 GNDA.t465 GNDA.n1869 0.159278
R4302 GNDA.t546 GNDA.n1870 0.159278
R4303 GNDA.t549 GNDA.n1871 0.159278
R4304 GNDA.t85 GNDA.n1872 0.159278
R4305 GNDA.t487 GNDA.n1873 0.159278
R4306 GNDA.t2 GNDA.n1874 0.159278
R4307 GNDA.t339 GNDA.n1875 0.159278
R4308 GNDA.t133 GNDA.n1876 0.159278
R4309 GNDA.t127 GNDA.n1877 0.159278
R4310 GNDA.n2152 GNDA.n410 0.15675
R4311 GNDA.n2149 GNDA.n2148 0.15675
R4312 GNDA.n1808 GNDA.n1807 0.151542
R4313 GNDA.n1976 GNDA.n1975 0.146333
R4314 GNDA.n1975 GNDA.n1836 0.146333
R4315 GNDA.n1971 GNDA.n1836 0.146333
R4316 GNDA.n1974 GNDA.n1832 0.146333
R4317 GNDA.n1974 GNDA.n1973 0.146333
R4318 GNDA.n1908 GNDA.n1900 0.146333
R4319 GNDA.n1909 GNDA.n1908 0.146333
R4320 GNDA.n1904 GNDA.n1903 0.146333
R4321 GNDA.n1907 GNDA.n1904 0.146333
R4322 GNDA.n1907 GNDA.n1899 0.146333
R4323 GNDA.n1927 GNDA.n1919 0.146333
R4324 GNDA.n1928 GNDA.n1927 0.146333
R4325 GNDA.n1923 GNDA.n1922 0.146333
R4326 GNDA.n1926 GNDA.n1923 0.146333
R4327 GNDA.n1926 GNDA.n1918 0.146333
R4328 GNDA.n1878 GNDA.t355 0.1368
R4329 GNDA.n1877 GNDA.t474 0.1368
R4330 GNDA.n1877 GNDA.t512 0.1368
R4331 GNDA.n1876 GNDA.t205 0.1368
R4332 GNDA.n1876 GNDA.t101 0.1368
R4333 GNDA.n1875 GNDA.t483 0.1368
R4334 GNDA.n1875 GNDA.t180 0.1368
R4335 GNDA.n1874 GNDA.t83 0.1368
R4336 GNDA.n1874 GNDA.t36 0.1368
R4337 GNDA.n1873 GNDA.t24 0.1368
R4338 GNDA.n1873 GNDA.t202 0.1368
R4339 GNDA.n1872 GNDA.t359 0.1368
R4340 GNDA.n1872 GNDA.t528 0.1368
R4341 GNDA.n1871 GNDA.t100 0.1368
R4342 GNDA.n1871 GNDA.t556 0.1368
R4343 GNDA.n1870 GNDA.t143 0.1368
R4344 GNDA.n1870 GNDA.t177 0.1368
R4345 GNDA.n1869 GNDA.t286 0.1368
R4346 GNDA.n1869 GNDA.t190 0.1368
R4347 GNDA.n1868 GNDA.t114 0.1368
R4348 GNDA.n1868 GNDA.t227 0.1368
R4349 GNDA.n1867 GNDA.t527 0.1368
R4350 GNDA.n1867 GNDA.t117 0.1368
R4351 GNDA.n1866 GNDA.t475 0.1368
R4352 GNDA.n1866 GNDA.t513 0.1368
R4353 GNDA.n1865 GNDA.t538 0.1368
R4354 GNDA.n1865 GNDA.t247 0.1368
R4355 GNDA.n1864 GNDA.t342 0.1368
R4356 GNDA.n1864 GNDA.t19 0.1368
R4357 GNDA.n1863 GNDA.t176 0.1368
R4358 GNDA.n1863 GNDA.t351 0.1368
R4359 GNDA.n1862 GNDA.t189 0.1368
R4360 GNDA.n1862 GNDA.t581 0.1368
R4361 GNDA.n1861 GNDA.t226 0.1368
R4362 GNDA.n1861 GNDA.t132 0.1368
R4363 GNDA.n1860 GNDA.t115 0.1368
R4364 GNDA.n1860 GNDA.t480 0.1368
R4365 GNDA.n1859 GNDA.t509 0.1368
R4366 GNDA.n1859 GNDA.t103 0.1368
R4367 GNDA.n1858 GNDA.t248 0.1368
R4368 GNDA.n1858 GNDA.t492 0.1368
R4369 GNDA.n1857 GNDA.t580 0.1368
R4370 GNDA.n1857 GNDA.t471 0.1368
R4371 GNDA.n1856 GNDA.t58 0.1368
R4372 GNDA.n1856 GNDA.t139 0.1368
R4373 GNDA.n1855 GNDA.t201 0.1368
R4374 GNDA.n1855 GNDA.t544 0.1368
R4375 GNDA.t50 GNDA.n1878 0.1368
R4376 GNDA.n1941 GNDA.t360 0.1368
R4377 GNDA.n1977 GNDA.n1976 0.135917
R4378 GNDA.n1978 GNDA.n1832 0.135917
R4379 GNDA.n1913 GNDA.n1909 0.135917
R4380 GNDA.n1914 GNDA.n1899 0.135917
R4381 GNDA.n1930 GNDA.n1928 0.135917
R4382 GNDA.n1931 GNDA.n1918 0.135917
R4383 GNDA.n706 GNDA.n705 0.1255
R4384 GNDA.n2161 GNDA.n405 0.1255
R4385 GNDA.n1810 GNDA.n1809 0.115083
R4386 GNDA.n1807 GNDA.n1806 0.115083
R4387 GNDA.n1806 GNDA.n1805 0.115083
R4388 GNDA.n1805 GNDA.n1804 0.115083
R4389 GNDA.n1804 GNDA.n410 0.115083
R4390 GNDA.n2152 GNDA.n2151 0.115083
R4391 GNDA.n2151 GNDA.n2150 0.115083
R4392 GNDA.n2150 GNDA.n2149 0.115083
R4393 GNDA.n2148 GNDA.n2147 0.115083
R4394 GNDA.n2147 GNDA.n2146 0.115083
R4395 GNDA.n2146 GNDA.n2145 0.115083
R4396 GNDA.n1972 GNDA.n1971 0.0667303
R4397 GNDA.n1903 GNDA.n1901 0.0667303
R4398 GNDA.n1922 GNDA.n1920 0.0667303
R4399 GNDA.n1809 GNDA.n1808 0.063
R4400 GNDA.n706 GNDA.n703 0.0626438
R4401 GNDA.n405 GNDA.n404 0.0626438
R4402 GNDA.n1835 GNDA.n1834 0.0553333
R4403 GNDA.n1970 GNDA.n1969 0.0553333
R4404 GNDA.n1906 GNDA.n1905 0.0553333
R4405 GNDA.n1925 GNDA.n1924 0.0553333
R4406 GNDA GNDA.n1178 0.0517
R4407 GNDA GNDA.n686 0.0517
R4408 GNDA GNDA.n1057 0.0517
R4409 GNDA.n2209 GNDA 0.0517
R4410 GNDA.n1671 GNDA 0.0517
R4411 GNDA.n1299 GNDA 0.0517
R4412 GNDA.n575 GNDA 0.0517
R4413 GNDA GNDA.n0 0.0517
R4414 GNDA.n1573 GNDA 0.0517
R4415 GNDA.n1902 GNDA.n1895 0.0514167
R4416 GNDA.n1915 GNDA.n1898 0.0514167
R4417 GNDA.n1921 GNDA.n1892 0.0514167
R4418 GNDA.n1932 GNDA.n1917 0.0514167
R4419 GNDA.n2165 GNDA.n401 0.0421667
R4420 GNDA.n1905 GNDA.n1896 0.028198
R4421 GNDA.n1898 GNDA.n1897 0.028198
R4422 GNDA.n1924 GNDA.n1893 0.028198
R4423 GNDA.n1917 GNDA.n1894 0.028198
R4424 GNDA.n1925 GNDA.n1894 0.028198
R4425 GNDA.n1921 GNDA.n1893 0.028198
R4426 GNDA.n1906 GNDA.n1897 0.028198
R4427 GNDA.n1902 GNDA.n1896 0.028198
R4428 GNDA.n1968 GNDA.n1835 0.028198
R4429 GNDA.n1969 GNDA.n1968 0.028198
R4430 GNDA.n1970 GNDA.n1837 0.0262697
R4431 GNDA.n1834 GNDA.n1833 0.0262697
R4432 GNDA.n2173 GNDA.n395 0.0217373
R4433 GNDA.n2169 GNDA.n396 0.0217373
R4434 GNDA.n2167 GNDA.n2166 0.0217373
R4435 GNDA.n2164 GNDA.n403 0.0217373
R4436 GNDA.n397 GNDA.n395 0.0217373
R4437 GNDA.n2169 GNDA.n2168 0.0217373
R4438 GNDA.n2166 GNDA.n400 0.0217373
R4439 GNDA.n403 GNDA.n400 0.0217373
R4440 GNDA.n2171 GNDA.n397 0.0217373
R4441 GNDA.n2172 GNDA.n396 0.0217373
R4442 GNDA.n2171 GNDA.n2170 0.0217373
R4443 GNDA.n2163 GNDA.n399 0.0217373
R4444 GNDA.n401 GNDA.n399 0.0217373
R4445 GNDA.n1941 GNDA.n1940 0.015775
R4446 GNDA.n1964 GNDA.n1956 0.0116625
R4447 GNDA.n1962 GNDA.n1956 0.0116625
R4448 GNDA.n1939 GNDA.n1888 0.0116625
R4449 GNDA.n1888 GNDA.n1884 0.0116625
R4450 GNDA.n1959 GNDA.n1951 0.0068649
R4451 GNDA.n1959 GNDA.n1958 0.0068649
R4452 GNDA.n1961 GNDA.n1952 0.0068649
R4453 GNDA.n1890 GNDA.n1880 0.0068649
R4454 GNDA.n1886 GNDA.n1880 0.0068649
R4455 GNDA.n1891 GNDA.n1881 0.0068649
R4456 GNDA.n1886 GNDA.n1883 0.0068649
R4457 GNDA.n1891 GNDA.n1883 0.0068649
R4458 GNDA.n1890 GNDA.n1884 0.0068649
R4459 GNDA.n1958 GNDA.n1955 0.0068649
R4460 GNDA.n1961 GNDA.n1955 0.0068649
R4461 GNDA.n1962 GNDA.n1951 0.0068649
R4462 GNDA.n1945 GNDA.n1944 0.0068649
R4463 GNDA.n1854 GNDA.n1852 0.0068649
R4464 GNDA.n1942 GNDA.n1843 0.0068649
R4465 GNDA.n1942 GNDA.n1841 0.0068649
R4466 GNDA.n1944 GNDA.n1854 0.0068649
R4467 GNDA.n1852 GNDA.n1843 0.0068649
R4468 GNDA.n1953 GNDA.n1952 0.00657213
R4469 GNDA.n1966 GNDA.n1838 0.00657213
R4470 GNDA.n1936 GNDA.n1881 0.00657213
R4471 GNDA.n1934 GNDA.n1882 0.00657213
R4472 GNDA.n1937 GNDA.n1936 0.00657213
R4473 GNDA.n1937 GNDA.n1882 0.00657213
R4474 GNDA.n1954 GNDA.n1953 0.00657213
R4475 GNDA.n1954 GNDA.n1838 0.00657213
R4476 GNDA.n1947 GNDA.n1846 0.00657213
R4477 GNDA.n1945 GNDA.n1844 0.00657213
R4478 GNDA.n1847 GNDA.n1841 0.00657213
R4479 GNDA.n1853 GNDA.n1842 0.00657213
R4480 GNDA.n1850 GNDA.n1846 0.00657213
R4481 GNDA.n1848 GNDA.n1847 0.00657213
R4482 GNDA.n1848 GNDA.n1842 0.00657213
R4483 GNDA.n1850 GNDA.n1844 0.00657213
R4484 GNDA.n1935 GNDA.n1885 0.00393497
R4485 GNDA.n1851 GNDA.n1845 0.00393497
R4486 GNDA.n1960 GNDA.n1839 0.00393497
R4487 GNDA.n1938 GNDA.n1935 0.00393497
R4488 GNDA.n1963 GNDA.n1960 0.00393497
R4489 GNDA.n1946 GNDA.n1851 0.00393497
R4490 GNDA.n1938 GNDA.n1889 0.0036417
R4491 GNDA.n1940 GNDA.n1879 0.0036417
R4492 GNDA.n1946 GNDA.n1849 0.0036417
R4493 GNDA.n1948 GNDA.n1840 0.0036417
R4494 GNDA.n1963 GNDA.n1957 0.0036417
R4495 GNDA.n1965 GNDA.n1950 0.0036417
R4496 GNDA.n1889 GNDA.n1887 0.0036417
R4497 GNDA.n1885 GNDA.n1879 0.0036417
R4498 GNDA.n1957 GNDA.n1949 0.0036417
R4499 GNDA.n1950 GNDA.n1839 0.0036417
R4500 GNDA.n1943 GNDA.n1849 0.0036417
R4501 GNDA.n1845 GNDA.n1840 0.0036417
R4502 GNDA.n1855 GNDA.t121 0.00152174
R4503 GNDA.n1856 GNDA.t520 0.00152174
R4504 GNDA.n1857 GNDA.t185 0.00152174
R4505 GNDA.n1858 GNDA.t515 0.00152174
R4506 GNDA.n1859 GNDA.t70 0.00152174
R4507 GNDA.n1860 GNDA.t501 0.00152174
R4508 GNDA.n1861 GNDA.t150 0.00152174
R4509 GNDA.n1862 GNDA.t74 0.00152174
R4510 GNDA.n1863 GNDA.t571 0.00152174
R4511 GNDA.n1864 GNDA.t529 0.00152174
R4512 GNDA.n1865 GNDA.t477 0.00152174
R4513 GNDA.n1866 GNDA.t356 0.00152174
R4514 GNDA.n1867 GNDA.t161 0.00152174
R4515 GNDA.n1868 GNDA.t352 0.00152174
R4516 GNDA.n1869 GNDA.t48 0.00152174
R4517 GNDA.n1870 GNDA.t465 0.00152174
R4518 GNDA.n1871 GNDA.t546 0.00152174
R4519 GNDA.n1872 GNDA.t549 0.00152174
R4520 GNDA.n1873 GNDA.t85 0.00152174
R4521 GNDA.n1874 GNDA.t487 0.00152174
R4522 GNDA.n1875 GNDA.t2 0.00152174
R4523 GNDA.n1876 GNDA.t339 0.00152174
R4524 GNDA.n1877 GNDA.t133 0.00152174
R4525 GNDA.n1878 GNDA.t127 0.00152174
R4526 two_stage_opamp_dummy_magic_23_0.Vb3.n25 two_stage_opamp_dummy_magic_23_0.Vb3.t20 768.551
R4527 two_stage_opamp_dummy_magic_23_0.Vb3.n19 two_stage_opamp_dummy_magic_23_0.Vb3.t8 611.739
R4528 two_stage_opamp_dummy_magic_23_0.Vb3.n15 two_stage_opamp_dummy_magic_23_0.Vb3.t25 611.739
R4529 two_stage_opamp_dummy_magic_23_0.Vb3.n10 two_stage_opamp_dummy_magic_23_0.Vb3.t22 611.739
R4530 two_stage_opamp_dummy_magic_23_0.Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb3.t16 611.739
R4531 two_stage_opamp_dummy_magic_23_0.Vb3.n24 two_stage_opamp_dummy_magic_23_0.Vb3.n23 428.976
R4532 two_stage_opamp_dummy_magic_23_0.Vb3.n24 two_stage_opamp_dummy_magic_23_0.Vb3.n14 428.445
R4533 two_stage_opamp_dummy_magic_23_0.Vb3.n19 two_stage_opamp_dummy_magic_23_0.Vb3.t11 421.75
R4534 two_stage_opamp_dummy_magic_23_0.Vb3.n20 two_stage_opamp_dummy_magic_23_0.Vb3.t28 421.75
R4535 two_stage_opamp_dummy_magic_23_0.Vb3.n21 two_stage_opamp_dummy_magic_23_0.Vb3.t18 421.75
R4536 two_stage_opamp_dummy_magic_23_0.Vb3.n22 two_stage_opamp_dummy_magic_23_0.Vb3.t15 421.75
R4537 two_stage_opamp_dummy_magic_23_0.Vb3.n15 two_stage_opamp_dummy_magic_23_0.Vb3.t27 421.75
R4538 two_stage_opamp_dummy_magic_23_0.Vb3.n16 two_stage_opamp_dummy_magic_23_0.Vb3.t10 421.75
R4539 two_stage_opamp_dummy_magic_23_0.Vb3.n17 two_stage_opamp_dummy_magic_23_0.Vb3.t14 421.75
R4540 two_stage_opamp_dummy_magic_23_0.Vb3.n18 two_stage_opamp_dummy_magic_23_0.Vb3.t12 421.75
R4541 two_stage_opamp_dummy_magic_23_0.Vb3.n10 two_stage_opamp_dummy_magic_23_0.Vb3.t24 421.75
R4542 two_stage_opamp_dummy_magic_23_0.Vb3.n11 two_stage_opamp_dummy_magic_23_0.Vb3.t21 421.75
R4543 two_stage_opamp_dummy_magic_23_0.Vb3.n12 two_stage_opamp_dummy_magic_23_0.Vb3.t17 421.75
R4544 two_stage_opamp_dummy_magic_23_0.Vb3.n13 two_stage_opamp_dummy_magic_23_0.Vb3.t13 421.75
R4545 two_stage_opamp_dummy_magic_23_0.Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb3.t19 421.75
R4546 two_stage_opamp_dummy_magic_23_0.Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb3.t23 421.75
R4547 two_stage_opamp_dummy_magic_23_0.Vb3.n8 two_stage_opamp_dummy_magic_23_0.Vb3.t26 421.75
R4548 two_stage_opamp_dummy_magic_23_0.Vb3.n9 two_stage_opamp_dummy_magic_23_0.Vb3.t9 421.75
R4549 two_stage_opamp_dummy_magic_23_0.Vb3.n20 two_stage_opamp_dummy_magic_23_0.Vb3.n19 167.094
R4550 two_stage_opamp_dummy_magic_23_0.Vb3.n21 two_stage_opamp_dummy_magic_23_0.Vb3.n20 167.094
R4551 two_stage_opamp_dummy_magic_23_0.Vb3.n22 two_stage_opamp_dummy_magic_23_0.Vb3.n21 167.094
R4552 two_stage_opamp_dummy_magic_23_0.Vb3.n16 two_stage_opamp_dummy_magic_23_0.Vb3.n15 167.094
R4553 two_stage_opamp_dummy_magic_23_0.Vb3.n17 two_stage_opamp_dummy_magic_23_0.Vb3.n16 167.094
R4554 two_stage_opamp_dummy_magic_23_0.Vb3.n18 two_stage_opamp_dummy_magic_23_0.Vb3.n17 167.094
R4555 two_stage_opamp_dummy_magic_23_0.Vb3.n11 two_stage_opamp_dummy_magic_23_0.Vb3.n10 167.094
R4556 two_stage_opamp_dummy_magic_23_0.Vb3.n12 two_stage_opamp_dummy_magic_23_0.Vb3.n11 167.094
R4557 two_stage_opamp_dummy_magic_23_0.Vb3.n13 two_stage_opamp_dummy_magic_23_0.Vb3.n12 167.094
R4558 two_stage_opamp_dummy_magic_23_0.Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb3.n6 167.094
R4559 two_stage_opamp_dummy_magic_23_0.Vb3.n8 two_stage_opamp_dummy_magic_23_0.Vb3.n7 167.094
R4560 two_stage_opamp_dummy_magic_23_0.Vb3.n9 two_stage_opamp_dummy_magic_23_0.Vb3.n8 167.094
R4561 two_stage_opamp_dummy_magic_23_0.Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb3.n0 139.639
R4562 two_stage_opamp_dummy_magic_23_0.Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb3.n1 139.638
R4563 two_stage_opamp_dummy_magic_23_0.Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb3.n3 134.577
R4564 two_stage_opamp_dummy_magic_23_0.Vb3.n26 two_stage_opamp_dummy_magic_23_0.Vb3.n5 73.3151
R4565 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb3.n26 51.4318
R4566 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb3.n4 44.313
R4567 two_stage_opamp_dummy_magic_23_0.Vb3.n23 two_stage_opamp_dummy_magic_23_0.Vb3.n22 35.3472
R4568 two_stage_opamp_dummy_magic_23_0.Vb3.n23 two_stage_opamp_dummy_magic_23_0.Vb3.n18 35.3472
R4569 two_stage_opamp_dummy_magic_23_0.Vb3.n14 two_stage_opamp_dummy_magic_23_0.Vb3.n13 35.3472
R4570 two_stage_opamp_dummy_magic_23_0.Vb3.n14 two_stage_opamp_dummy_magic_23_0.Vb3.n9 35.3472
R4571 two_stage_opamp_dummy_magic_23_0.Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb3.t3 24.0005
R4572 two_stage_opamp_dummy_magic_23_0.Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb3.t0 24.0005
R4573 two_stage_opamp_dummy_magic_23_0.Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb3.t7 24.0005
R4574 two_stage_opamp_dummy_magic_23_0.Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb3.t6 24.0005
R4575 two_stage_opamp_dummy_magic_23_0.Vb3.n0 two_stage_opamp_dummy_magic_23_0.Vb3.t5 24.0005
R4576 two_stage_opamp_dummy_magic_23_0.Vb3.n0 two_stage_opamp_dummy_magic_23_0.Vb3.t2 24.0005
R4577 two_stage_opamp_dummy_magic_23_0.Vb3.n25 two_stage_opamp_dummy_magic_23_0.Vb3.n24 14.3443
R4578 two_stage_opamp_dummy_magic_23_0.Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb3.t4 11.2576
R4579 two_stage_opamp_dummy_magic_23_0.Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb3.t1 11.2576
R4580 two_stage_opamp_dummy_magic_23_0.Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb3.n2 4.5005
R4581 two_stage_opamp_dummy_magic_23_0.Vb3.n26 two_stage_opamp_dummy_magic_23_0.Vb3.n25 1.21925
R4582 two_stage_opamp_dummy_magic_23_0.Y.n65 two_stage_opamp_dummy_magic_23_0.Y.t28 1172.87
R4583 two_stage_opamp_dummy_magic_23_0.Y.n63 two_stage_opamp_dummy_magic_23_0.Y.t50 1172.87
R4584 two_stage_opamp_dummy_magic_23_0.Y.n65 two_stage_opamp_dummy_magic_23_0.Y.t44 996.134
R4585 two_stage_opamp_dummy_magic_23_0.Y.n66 two_stage_opamp_dummy_magic_23_0.Y.t30 996.134
R4586 two_stage_opamp_dummy_magic_23_0.Y.n67 two_stage_opamp_dummy_magic_23_0.Y.t38 996.134
R4587 two_stage_opamp_dummy_magic_23_0.Y.n68 two_stage_opamp_dummy_magic_23_0.Y.t53 996.134
R4588 two_stage_opamp_dummy_magic_23_0.Y.n69 two_stage_opamp_dummy_magic_23_0.Y.t40 996.134
R4589 two_stage_opamp_dummy_magic_23_0.Y.n70 two_stage_opamp_dummy_magic_23_0.Y.t25 996.134
R4590 two_stage_opamp_dummy_magic_23_0.Y.n64 two_stage_opamp_dummy_magic_23_0.Y.t42 996.134
R4591 two_stage_opamp_dummy_magic_23_0.Y.n63 two_stage_opamp_dummy_magic_23_0.Y.t35 996.134
R4592 two_stage_opamp_dummy_magic_23_0.Y.n58 two_stage_opamp_dummy_magic_23_0.Y.t54 690.867
R4593 two_stage_opamp_dummy_magic_23_0.Y.n51 two_stage_opamp_dummy_magic_23_0.Y.t47 690.867
R4594 two_stage_opamp_dummy_magic_23_0.Y.n49 two_stage_opamp_dummy_magic_23_0.Y.t49 530.201
R4595 two_stage_opamp_dummy_magic_23_0.Y.n42 two_stage_opamp_dummy_magic_23_0.Y.t43 530.201
R4596 two_stage_opamp_dummy_magic_23_0.Y.n58 two_stage_opamp_dummy_magic_23_0.Y.t41 514.134
R4597 two_stage_opamp_dummy_magic_23_0.Y.n51 two_stage_opamp_dummy_magic_23_0.Y.t32 514.134
R4598 two_stage_opamp_dummy_magic_23_0.Y.n52 two_stage_opamp_dummy_magic_23_0.Y.t39 514.134
R4599 two_stage_opamp_dummy_magic_23_0.Y.n53 two_stage_opamp_dummy_magic_23_0.Y.t51 514.134
R4600 two_stage_opamp_dummy_magic_23_0.Y.n54 two_stage_opamp_dummy_magic_23_0.Y.t36 514.134
R4601 two_stage_opamp_dummy_magic_23_0.Y.n55 two_stage_opamp_dummy_magic_23_0.Y.t48 514.134
R4602 two_stage_opamp_dummy_magic_23_0.Y.n56 two_stage_opamp_dummy_magic_23_0.Y.t33 514.134
R4603 two_stage_opamp_dummy_magic_23_0.Y.n57 two_stage_opamp_dummy_magic_23_0.Y.t26 514.134
R4604 two_stage_opamp_dummy_magic_23_0.Y.n49 two_stage_opamp_dummy_magic_23_0.Y.t37 353.467
R4605 two_stage_opamp_dummy_magic_23_0.Y.n48 two_stage_opamp_dummy_magic_23_0.Y.t52 353.467
R4606 two_stage_opamp_dummy_magic_23_0.Y.n47 two_stage_opamp_dummy_magic_23_0.Y.t29 353.467
R4607 two_stage_opamp_dummy_magic_23_0.Y.n46 two_stage_opamp_dummy_magic_23_0.Y.t45 353.467
R4608 two_stage_opamp_dummy_magic_23_0.Y.n45 two_stage_opamp_dummy_magic_23_0.Y.t31 353.467
R4609 two_stage_opamp_dummy_magic_23_0.Y.n44 two_stage_opamp_dummy_magic_23_0.Y.t46 353.467
R4610 two_stage_opamp_dummy_magic_23_0.Y.n43 two_stage_opamp_dummy_magic_23_0.Y.t34 353.467
R4611 two_stage_opamp_dummy_magic_23_0.Y.n42 two_stage_opamp_dummy_magic_23_0.Y.t27 353.467
R4612 two_stage_opamp_dummy_magic_23_0.Y.n72 two_stage_opamp_dummy_magic_23_0.Y.n71 304.375
R4613 two_stage_opamp_dummy_magic_23_0.Y.n60 two_stage_opamp_dummy_magic_23_0.Y.n50 216.9
R4614 two_stage_opamp_dummy_magic_23_0.Y.n60 two_stage_opamp_dummy_magic_23_0.Y.n59 216.9
R4615 two_stage_opamp_dummy_magic_23_0.Y.n64 two_stage_opamp_dummy_magic_23_0.Y.n63 176.733
R4616 two_stage_opamp_dummy_magic_23_0.Y.n66 two_stage_opamp_dummy_magic_23_0.Y.n65 176.733
R4617 two_stage_opamp_dummy_magic_23_0.Y.n67 two_stage_opamp_dummy_magic_23_0.Y.n66 176.733
R4618 two_stage_opamp_dummy_magic_23_0.Y.n68 two_stage_opamp_dummy_magic_23_0.Y.n67 176.733
R4619 two_stage_opamp_dummy_magic_23_0.Y.n69 two_stage_opamp_dummy_magic_23_0.Y.n68 176.733
R4620 two_stage_opamp_dummy_magic_23_0.Y.n70 two_stage_opamp_dummy_magic_23_0.Y.n69 176.733
R4621 two_stage_opamp_dummy_magic_23_0.Y.n48 two_stage_opamp_dummy_magic_23_0.Y.n47 176.733
R4622 two_stage_opamp_dummy_magic_23_0.Y.n47 two_stage_opamp_dummy_magic_23_0.Y.n46 176.733
R4623 two_stage_opamp_dummy_magic_23_0.Y.n46 two_stage_opamp_dummy_magic_23_0.Y.n45 176.733
R4624 two_stage_opamp_dummy_magic_23_0.Y.n45 two_stage_opamp_dummy_magic_23_0.Y.n44 176.733
R4625 two_stage_opamp_dummy_magic_23_0.Y.n44 two_stage_opamp_dummy_magic_23_0.Y.n43 176.733
R4626 two_stage_opamp_dummy_magic_23_0.Y.n43 two_stage_opamp_dummy_magic_23_0.Y.n42 176.733
R4627 two_stage_opamp_dummy_magic_23_0.Y.n57 two_stage_opamp_dummy_magic_23_0.Y.n56 176.733
R4628 two_stage_opamp_dummy_magic_23_0.Y.n56 two_stage_opamp_dummy_magic_23_0.Y.n55 176.733
R4629 two_stage_opamp_dummy_magic_23_0.Y.n55 two_stage_opamp_dummy_magic_23_0.Y.n54 176.733
R4630 two_stage_opamp_dummy_magic_23_0.Y.n54 two_stage_opamp_dummy_magic_23_0.Y.n53 176.733
R4631 two_stage_opamp_dummy_magic_23_0.Y.n53 two_stage_opamp_dummy_magic_23_0.Y.n52 176.733
R4632 two_stage_opamp_dummy_magic_23_0.Y.n52 two_stage_opamp_dummy_magic_23_0.Y.n51 176.733
R4633 two_stage_opamp_dummy_magic_23_0.Y.n61 two_stage_opamp_dummy_magic_23_0.Y.n60 175.05
R4634 two_stage_opamp_dummy_magic_23_0.Y.n22 two_stage_opamp_dummy_magic_23_0.Y.n21 66.0338
R4635 two_stage_opamp_dummy_magic_23_0.Y.n26 two_stage_opamp_dummy_magic_23_0.Y.n25 66.0338
R4636 two_stage_opamp_dummy_magic_23_0.Y.n28 two_stage_opamp_dummy_magic_23_0.Y.n27 66.0338
R4637 two_stage_opamp_dummy_magic_23_0.Y.n32 two_stage_opamp_dummy_magic_23_0.Y.n31 66.0338
R4638 two_stage_opamp_dummy_magic_23_0.Y.n35 two_stage_opamp_dummy_magic_23_0.Y.n34 66.0338
R4639 two_stage_opamp_dummy_magic_23_0.Y.n39 two_stage_opamp_dummy_magic_23_0.Y.n38 66.0338
R4640 two_stage_opamp_dummy_magic_23_0.Y.t16 two_stage_opamp_dummy_magic_23_0.Y.n72 49.4802
R4641 two_stage_opamp_dummy_magic_23_0.Y.n1 two_stage_opamp_dummy_magic_23_0.Y.n0 49.3505
R4642 two_stage_opamp_dummy_magic_23_0.Y.n6 two_stage_opamp_dummy_magic_23_0.Y.n5 49.3505
R4643 two_stage_opamp_dummy_magic_23_0.Y.n9 two_stage_opamp_dummy_magic_23_0.Y.n8 49.3505
R4644 two_stage_opamp_dummy_magic_23_0.Y.n12 two_stage_opamp_dummy_magic_23_0.Y.n11 49.3505
R4645 two_stage_opamp_dummy_magic_23_0.Y.n4 two_stage_opamp_dummy_magic_23_0.Y.n3 49.3505
R4646 two_stage_opamp_dummy_magic_23_0.Y.n17 two_stage_opamp_dummy_magic_23_0.Y.n16 49.3505
R4647 two_stage_opamp_dummy_magic_23_0.Y.n71 two_stage_opamp_dummy_magic_23_0.Y.n64 40.1672
R4648 two_stage_opamp_dummy_magic_23_0.Y.n71 two_stage_opamp_dummy_magic_23_0.Y.n70 40.1672
R4649 two_stage_opamp_dummy_magic_23_0.Y.n50 two_stage_opamp_dummy_magic_23_0.Y.n48 40.1672
R4650 two_stage_opamp_dummy_magic_23_0.Y.n50 two_stage_opamp_dummy_magic_23_0.Y.n49 40.1672
R4651 two_stage_opamp_dummy_magic_23_0.Y.n59 two_stage_opamp_dummy_magic_23_0.Y.n57 40.1672
R4652 two_stage_opamp_dummy_magic_23_0.Y.n59 two_stage_opamp_dummy_magic_23_0.Y.n58 40.1672
R4653 two_stage_opamp_dummy_magic_23_0.Y.n61 two_stage_opamp_dummy_magic_23_0.Y.n41 17.6567
R4654 two_stage_opamp_dummy_magic_23_0.Y.n0 two_stage_opamp_dummy_magic_23_0.Y.t17 16.0005
R4655 two_stage_opamp_dummy_magic_23_0.Y.n0 two_stage_opamp_dummy_magic_23_0.Y.t12 16.0005
R4656 two_stage_opamp_dummy_magic_23_0.Y.n5 two_stage_opamp_dummy_magic_23_0.Y.t23 16.0005
R4657 two_stage_opamp_dummy_magic_23_0.Y.n5 two_stage_opamp_dummy_magic_23_0.Y.t0 16.0005
R4658 two_stage_opamp_dummy_magic_23_0.Y.n8 two_stage_opamp_dummy_magic_23_0.Y.t11 16.0005
R4659 two_stage_opamp_dummy_magic_23_0.Y.n8 two_stage_opamp_dummy_magic_23_0.Y.t8 16.0005
R4660 two_stage_opamp_dummy_magic_23_0.Y.n11 two_stage_opamp_dummy_magic_23_0.Y.t9 16.0005
R4661 two_stage_opamp_dummy_magic_23_0.Y.n11 two_stage_opamp_dummy_magic_23_0.Y.t7 16.0005
R4662 two_stage_opamp_dummy_magic_23_0.Y.n3 two_stage_opamp_dummy_magic_23_0.Y.t19 16.0005
R4663 two_stage_opamp_dummy_magic_23_0.Y.n3 two_stage_opamp_dummy_magic_23_0.Y.t24 16.0005
R4664 two_stage_opamp_dummy_magic_23_0.Y.n16 two_stage_opamp_dummy_magic_23_0.Y.t18 16.0005
R4665 two_stage_opamp_dummy_magic_23_0.Y.n16 two_stage_opamp_dummy_magic_23_0.Y.t13 16.0005
R4666 two_stage_opamp_dummy_magic_23_0.Y.n21 two_stage_opamp_dummy_magic_23_0.Y.t5 11.2576
R4667 two_stage_opamp_dummy_magic_23_0.Y.n21 two_stage_opamp_dummy_magic_23_0.Y.t10 11.2576
R4668 two_stage_opamp_dummy_magic_23_0.Y.n25 two_stage_opamp_dummy_magic_23_0.Y.t20 11.2576
R4669 two_stage_opamp_dummy_magic_23_0.Y.n25 two_stage_opamp_dummy_magic_23_0.Y.t4 11.2576
R4670 two_stage_opamp_dummy_magic_23_0.Y.n27 two_stage_opamp_dummy_magic_23_0.Y.t2 11.2576
R4671 two_stage_opamp_dummy_magic_23_0.Y.n27 two_stage_opamp_dummy_magic_23_0.Y.t22 11.2576
R4672 two_stage_opamp_dummy_magic_23_0.Y.n31 two_stage_opamp_dummy_magic_23_0.Y.t15 11.2576
R4673 two_stage_opamp_dummy_magic_23_0.Y.n31 two_stage_opamp_dummy_magic_23_0.Y.t3 11.2576
R4674 two_stage_opamp_dummy_magic_23_0.Y.n34 two_stage_opamp_dummy_magic_23_0.Y.t1 11.2576
R4675 two_stage_opamp_dummy_magic_23_0.Y.n34 two_stage_opamp_dummy_magic_23_0.Y.t14 11.2576
R4676 two_stage_opamp_dummy_magic_23_0.Y.n38 two_stage_opamp_dummy_magic_23_0.Y.t6 11.2576
R4677 two_stage_opamp_dummy_magic_23_0.Y.n38 two_stage_opamp_dummy_magic_23_0.Y.t21 11.2576
R4678 two_stage_opamp_dummy_magic_23_0.Y.n62 two_stage_opamp_dummy_magic_23_0.Y.n20 10.2817
R4679 two_stage_opamp_dummy_magic_23_0.Y.n29 two_stage_opamp_dummy_magic_23_0.Y.n26 5.91717
R4680 two_stage_opamp_dummy_magic_23_0.Y.n26 two_stage_opamp_dummy_magic_23_0.Y.n24 5.91717
R4681 two_stage_opamp_dummy_magic_23_0.Y.n37 two_stage_opamp_dummy_magic_23_0.Y.n22 5.91717
R4682 two_stage_opamp_dummy_magic_23_0.Y.n15 two_stage_opamp_dummy_magic_23_0.Y.n4 5.6255
R4683 two_stage_opamp_dummy_magic_23_0.Y.n10 two_stage_opamp_dummy_magic_23_0.Y.n6 5.6255
R4684 two_stage_opamp_dummy_magic_23_0.Y.n18 two_stage_opamp_dummy_magic_23_0.Y.n4 5.438
R4685 two_stage_opamp_dummy_magic_23_0.Y.n7 two_stage_opamp_dummy_magic_23_0.Y.n6 5.438
R4686 two_stage_opamp_dummy_magic_23_0.Y.n28 two_stage_opamp_dummy_magic_23_0.Y.n24 5.29217
R4687 two_stage_opamp_dummy_magic_23_0.Y.n29 two_stage_opamp_dummy_magic_23_0.Y.n28 5.29217
R4688 two_stage_opamp_dummy_magic_23_0.Y.n33 two_stage_opamp_dummy_magic_23_0.Y.n32 5.29217
R4689 two_stage_opamp_dummy_magic_23_0.Y.n32 two_stage_opamp_dummy_magic_23_0.Y.n30 5.29217
R4690 two_stage_opamp_dummy_magic_23_0.Y.n36 two_stage_opamp_dummy_magic_23_0.Y.n35 5.29217
R4691 two_stage_opamp_dummy_magic_23_0.Y.n35 two_stage_opamp_dummy_magic_23_0.Y.n23 5.29217
R4692 two_stage_opamp_dummy_magic_23_0.Y.n39 two_stage_opamp_dummy_magic_23_0.Y.n37 5.29217
R4693 two_stage_opamp_dummy_magic_23_0.Y.n40 two_stage_opamp_dummy_magic_23_0.Y.n39 5.29217
R4694 two_stage_opamp_dummy_magic_23_0.Y.n41 two_stage_opamp_dummy_magic_23_0.Y.n40 5.1255
R4695 two_stage_opamp_dummy_magic_23_0.Y.n10 two_stage_opamp_dummy_magic_23_0.Y.n9 5.063
R4696 two_stage_opamp_dummy_magic_23_0.Y.n13 two_stage_opamp_dummy_magic_23_0.Y.n12 5.063
R4697 two_stage_opamp_dummy_magic_23_0.Y.n17 two_stage_opamp_dummy_magic_23_0.Y.n15 5.063
R4698 two_stage_opamp_dummy_magic_23_0.Y.n14 two_stage_opamp_dummy_magic_23_0.Y.n1 5.063
R4699 two_stage_opamp_dummy_magic_23_0.Y.n9 two_stage_opamp_dummy_magic_23_0.Y.n7 4.8755
R4700 two_stage_opamp_dummy_magic_23_0.Y.n12 two_stage_opamp_dummy_magic_23_0.Y.n2 4.8755
R4701 two_stage_opamp_dummy_magic_23_0.Y.n18 two_stage_opamp_dummy_magic_23_0.Y.n17 4.8755
R4702 two_stage_opamp_dummy_magic_23_0.Y.n20 two_stage_opamp_dummy_magic_23_0.Y.n19 4.5005
R4703 two_stage_opamp_dummy_magic_23_0.Y.n62 two_stage_opamp_dummy_magic_23_0.Y.n61 4.5005
R4704 two_stage_opamp_dummy_magic_23_0.Y.n72 two_stage_opamp_dummy_magic_23_0.Y.n62 3.27133
R4705 two_stage_opamp_dummy_magic_23_0.Y.n41 two_stage_opamp_dummy_magic_23_0.Y.n22 0.792167
R4706 two_stage_opamp_dummy_magic_23_0.Y.n40 two_stage_opamp_dummy_magic_23_0.Y.n23 0.6255
R4707 two_stage_opamp_dummy_magic_23_0.Y.n30 two_stage_opamp_dummy_magic_23_0.Y.n23 0.6255
R4708 two_stage_opamp_dummy_magic_23_0.Y.n30 two_stage_opamp_dummy_magic_23_0.Y.n29 0.6255
R4709 two_stage_opamp_dummy_magic_23_0.Y.n33 two_stage_opamp_dummy_magic_23_0.Y.n24 0.6255
R4710 two_stage_opamp_dummy_magic_23_0.Y.n36 two_stage_opamp_dummy_magic_23_0.Y.n33 0.6255
R4711 two_stage_opamp_dummy_magic_23_0.Y.n37 two_stage_opamp_dummy_magic_23_0.Y.n36 0.6255
R4712 two_stage_opamp_dummy_magic_23_0.Y.n15 two_stage_opamp_dummy_magic_23_0.Y.n14 0.563
R4713 two_stage_opamp_dummy_magic_23_0.Y.n19 two_stage_opamp_dummy_magic_23_0.Y.n18 0.563
R4714 two_stage_opamp_dummy_magic_23_0.Y.n19 two_stage_opamp_dummy_magic_23_0.Y.n2 0.563
R4715 two_stage_opamp_dummy_magic_23_0.Y.n7 two_stage_opamp_dummy_magic_23_0.Y.n2 0.563
R4716 two_stage_opamp_dummy_magic_23_0.Y.n13 two_stage_opamp_dummy_magic_23_0.Y.n10 0.563
R4717 two_stage_opamp_dummy_magic_23_0.Y.n14 two_stage_opamp_dummy_magic_23_0.Y.n13 0.563
R4718 two_stage_opamp_dummy_magic_23_0.Y.n20 two_stage_opamp_dummy_magic_23_0.Y.n1 0.3755
R4719 VDDA.n579 VDDA.t305 1231.74
R4720 VDDA.n582 VDDA.t277 1231.74
R4721 VDDA.n498 VDDA.t366 1231.74
R4722 VDDA.n501 VDDA.t390 1231.74
R4723 VDDA.t372 VDDA.n564 1095.3
R4724 VDDA.n565 VDDA.t186 1095.3
R4725 VDDA.n525 VDDA.t287 1095.3
R4726 VDDA.t269 VDDA.n524 1095.3
R4727 VDDA.n484 VDDA.t381 1095.3
R4728 VDDA.t354 VDDA.n483 1095.3
R4729 VDDA.n427 VDDA.t210 758.64
R4730 VDDA.n536 VDDA.t350 672.293
R4731 VDDA.n539 VDDA.t265 672.293
R4732 VDDA.n455 VDDA.t227 672.293
R4733 VDDA.n458 VDDA.t339 672.293
R4734 VDDA.n564 VDDA.t373 663.801
R4735 VDDA.n565 VDDA.t187 663.801
R4736 VDDA.n525 VDDA.t288 663.801
R4737 VDDA.n524 VDDA.t270 663.801
R4738 VDDA.n484 VDDA.t382 663.801
R4739 VDDA.n483 VDDA.t355 663.801
R4740 VDDA.n597 VDDA.t241 661.375
R4741 VDDA.n600 VDDA.t314 661.375
R4742 VDDA.t275 VDDA.n402 643.037
R4743 VDDA.n403 VDDA.t334 643.037
R4744 VDDA.t249 VDDA.n388 643.037
R4745 VDDA.n389 VDDA.t193 643.037
R4746 VDDA.n397 VDDA.t387 642.992
R4747 VDDA.t328 VDDA.n396 642.992
R4748 VDDA.n381 VDDA.t225 642.992
R4749 VDDA.t362 VDDA.n380 642.992
R4750 VDDA.n504 VDDA.n503 599.342
R4751 VDDA.n506 VDDA.n505 599.342
R4752 VDDA.n508 VDDA.n507 599.342
R4753 VDDA.n510 VDDA.n509 599.342
R4754 VDDA.n512 VDDA.n511 599.342
R4755 VDDA.n514 VDDA.n513 599.342
R4756 VDDA.n516 VDDA.n515 599.342
R4757 VDDA.n518 VDDA.n517 599.342
R4758 VDDA.n520 VDDA.n519 599.342
R4759 VDDA.n522 VDDA.n521 599.342
R4760 VDDA.n351 VDDA.t344 595.842
R4761 VDDA.n557 VDDA.t356 589.076
R4762 VDDA.n560 VDDA.t330 589.076
R4763 VDDA.n476 VDDA.t207 589.076
R4764 VDDA.n479 VDDA.t233 589.076
R4765 VDDA.t396 VDDA.t372 580.557
R4766 VDDA.t421 VDDA.t396 580.557
R4767 VDDA.t12 VDDA.t421 580.557
R4768 VDDA.t34 VDDA.t12 580.557
R4769 VDDA.t10 VDDA.t34 580.557
R4770 VDDA.t414 VDDA.t10 580.557
R4771 VDDA.t65 VDDA.t414 580.557
R4772 VDDA.t92 VDDA.t65 580.557
R4773 VDDA.t33 VDDA.t92 580.557
R4774 VDDA.t420 VDDA.t33 580.557
R4775 VDDA.t186 VDDA.t420 580.557
R4776 VDDA.t287 VDDA.t49 580.557
R4777 VDDA.t49 VDDA.t6 580.557
R4778 VDDA.t6 VDDA.t81 580.557
R4779 VDDA.t81 VDDA.t17 580.557
R4780 VDDA.t17 VDDA.t4 580.557
R4781 VDDA.t4 VDDA.t62 580.557
R4782 VDDA.t62 VDDA.t1 580.557
R4783 VDDA.t1 VDDA.t21 580.557
R4784 VDDA.t21 VDDA.t59 580.557
R4785 VDDA.t59 VDDA.t83 580.557
R4786 VDDA.t83 VDDA.t47 580.557
R4787 VDDA.t47 VDDA.t19 580.557
R4788 VDDA.t19 VDDA.t55 580.557
R4789 VDDA.t55 VDDA.t74 580.557
R4790 VDDA.t74 VDDA.t67 580.557
R4791 VDDA.t67 VDDA.t417 580.557
R4792 VDDA.t417 VDDA.t45 580.557
R4793 VDDA.t45 VDDA.t69 580.557
R4794 VDDA.t69 VDDA.t23 580.557
R4795 VDDA.t23 VDDA.t30 580.557
R4796 VDDA.t30 VDDA.t269 580.557
R4797 VDDA.t381 VDDA.t413 580.557
R4798 VDDA.t413 VDDA.t64 580.557
R4799 VDDA.t64 VDDA.t11 580.557
R4800 VDDA.t11 VDDA.t66 580.557
R4801 VDDA.t66 VDDA.t14 580.557
R4802 VDDA.t14 VDDA.t85 580.557
R4803 VDDA.t85 VDDA.t394 580.557
R4804 VDDA.t394 VDDA.t58 580.557
R4805 VDDA.t58 VDDA.t415 580.557
R4806 VDDA.t415 VDDA.t13 580.557
R4807 VDDA.t13 VDDA.t354 580.557
R4808 VDDA.n329 VDDA.t289 579.775
R4809 VDDA.n417 VDDA.n413 510.991
R4810 VDDA.n439 VDDA.n438 504.726
R4811 VDDA.n340 VDDA.t291 464.281
R4812 VDDA.n337 VDDA.t291 464.281
R4813 VDDA.n346 VDDA.t347 464.281
R4814 VDDA.t347 VDDA.n330 464.281
R4815 VDDA.n589 VDDA.t244 456.526
R4816 VDDA.n592 VDDA.t230 456.526
R4817 VDDA.n395 VDDA.t327 441.2
R4818 VDDA.n398 VDDA.t386 441.2
R4819 VDDA.n379 VDDA.t361 441.2
R4820 VDDA.n382 VDDA.t224 441.2
R4821 VDDA.n399 VDDA.t274 409.067
R4822 VDDA.n404 VDDA.t333 409.067
R4823 VDDA.n591 VDDA.t231 397.784
R4824 VDDA.t245 VDDA.n590 397.784
R4825 VDDA.n387 VDDA.t248 390.322
R4826 VDDA.n390 VDDA.t192 390.322
R4827 VDDA.t205 VDDA.t275 373.214
R4828 VDDA.t337 VDDA.t205 373.214
R4829 VDDA.t272 VDDA.t337 373.214
R4830 VDDA.t202 VDDA.t272 373.214
R4831 VDDA.t334 VDDA.t202 373.214
R4832 VDDA.t263 VDDA.t328 373.214
R4833 VDDA.t199 VDDA.t263 373.214
R4834 VDDA.t325 VDDA.t199 373.214
R4835 VDDA.t260 VDDA.t325 373.214
R4836 VDDA.t384 VDDA.t260 373.214
R4837 VDDA.t309 VDDA.t384 373.214
R4838 VDDA.t312 VDDA.t309 373.214
R4839 VDDA.t237 VDDA.t312 373.214
R4840 VDDA.t387 VDDA.t237 373.214
R4841 VDDA.t255 VDDA.t249 373.214
R4842 VDDA.t196 VDDA.t255 373.214
R4843 VDDA.t322 VDDA.t196 373.214
R4844 VDDA.t252 VDDA.t322 373.214
R4845 VDDA.t193 VDDA.t252 373.214
R4846 VDDA.t293 VDDA.t362 373.214
R4847 VDDA.t220 VDDA.t293 373.214
R4848 VDDA.t225 VDDA.t220 373.214
R4849 VDDA.n0 VDDA.t581 369.534
R4850 VDDA.n435 VDDA.t262 369.534
R4851 VDDA.n432 VDDA.t236 369.534
R4852 VDDA.n415 VDDA.t251 369.534
R4853 VDDA.n414 VDDA.t254 369.534
R4854 VDDA.n429 VDDA.t201 369.534
R4855 VDDA.n428 VDDA.t204 369.534
R4856 VDDA.n300 VDDA.t369 355.293
R4857 VDDA.n397 VDDA.t389 354.154
R4858 VDDA.n396 VDDA.t329 354.154
R4859 VDDA.n381 VDDA.t226 354.154
R4860 VDDA.n380 VDDA.t363 354.154
R4861 VDDA.n523 VDDA.t268 348.325
R4862 VDDA.n526 VDDA.t286 348.325
R4863 VDDA.n563 VDDA.t371 348.075
R4864 VDDA.n566 VDDA.t185 348.075
R4865 VDDA.n482 VDDA.t353 348.075
R4866 VDDA.n485 VDDA.t380 348.075
R4867 VDDA.n310 VDDA.t359 346.8
R4868 VDDA.n559 VDDA.t331 343.882
R4869 VDDA.t357 VDDA.n558 343.882
R4870 VDDA.t208 VDDA.n477 343.882
R4871 VDDA.n478 VDDA.t234 343.882
R4872 VDDA.n376 VDDA.n375 342.197
R4873 VDDA.n385 VDDA.n384 342.197
R4874 VDDA.n405 VDDA.n401 341.769
R4875 VDDA.n406 VDDA.n400 341.769
R4876 VDDA.n639 VDDA.n637 339.961
R4877 VDDA.n309 VDDA.n308 339.522
R4878 VDDA.n300 VDDA.n299 339.522
R4879 VDDA.n639 VDDA.n638 339.272
R4880 VDDA.n425 VDDA.n424 339.272
R4881 VDDA.n423 VDDA.n422 339.272
R4882 VDDA.n421 VDDA.n420 339.272
R4883 VDDA.n419 VDDA.n418 339.272
R4884 VDDA.n635 VDDA.n634 339.272
R4885 VDDA.n643 VDDA.n642 339.272
R4886 VDDA.n645 VDDA.n644 339.272
R4887 VDDA.n409 VDDA.n374 336.341
R4888 VDDA.n410 VDDA.n373 336.341
R4889 VDDA.n372 VDDA.n371 336.341
R4890 VDDA.n393 VDDA.n392 336.341
R4891 VDDA.n378 VDDA.n377 336.341
R4892 VDDA.n304 VDDA.n303 335.022
R4893 VDDA.n412 VDDA.n370 334.894
R4894 VDDA.n640 VDDA.n636 334.772
R4895 VDDA.n388 VDDA.t250 332.267
R4896 VDDA.n389 VDDA.t194 332.267
R4897 VDDA.n402 VDDA.t276 332.084
R4898 VDDA.n403 VDDA.t335 332.084
R4899 VDDA.t290 VDDA.n342 267.188
R4900 VDDA.n348 VDDA.t345 267.188
R4901 VDDA.t231 VDDA.t15 259.091
R4902 VDDA.t15 VDDA.t245 259.091
R4903 VDDA.n413 VDDA.t292 249.034
R4904 VDDA.n413 VDDA.t219 249.034
R4905 VDDA.n347 VDDA.n346 243.698
R4906 VDDA.n350 VDDA.n349 238.367
R4907 VDDA.n655 VDDA.n654 224.934
R4908 VDDA.n654 VDDA.n653 224.934
R4909 VDDA.n653 VDDA.n652 224.934
R4910 VDDA.n652 VDDA.n651 224.934
R4911 VDDA.n651 VDDA.n650 224.934
R4912 VDDA.n650 VDDA.n649 224.934
R4913 VDDA.n649 VDDA.n648 224.934
R4914 VDDA.n1 VDDA.n0 224.934
R4915 VDDA.n2 VDDA.n1 224.934
R4916 VDDA.n3 VDDA.n2 224.934
R4917 VDDA.n4 VDDA.n3 224.934
R4918 VDDA.n5 VDDA.n4 224.934
R4919 VDDA.t331 VDDA.t152 217.708
R4920 VDDA.t152 VDDA.t168 217.708
R4921 VDDA.t168 VDDA.t148 217.708
R4922 VDDA.t148 VDDA.t178 217.708
R4923 VDDA.t178 VDDA.t156 217.708
R4924 VDDA.t156 VDDA.t175 217.708
R4925 VDDA.t175 VDDA.t155 217.708
R4926 VDDA.t155 VDDA.t173 217.708
R4927 VDDA.t173 VDDA.t181 217.708
R4928 VDDA.t181 VDDA.t159 217.708
R4929 VDDA.t159 VDDA.t357 217.708
R4930 VDDA.t96 VDDA.t208 217.708
R4931 VDDA.t398 VDDA.t96 217.708
R4932 VDDA.t36 VDDA.t398 217.708
R4933 VDDA.t86 VDDA.t36 217.708
R4934 VDDA.t406 VDDA.t86 217.708
R4935 VDDA.t72 VDDA.t406 217.708
R4936 VDDA.t95 VDDA.t72 217.708
R4937 VDDA.t88 VDDA.t95 217.708
R4938 VDDA.t94 VDDA.t88 217.708
R4939 VDDA.t76 VDDA.t94 217.708
R4940 VDDA.t234 VDDA.t76 217.708
R4941 VDDA.t211 VDDA.t290 217.708
R4942 VDDA.t345 VDDA.t211 217.708
R4943 VDDA VDDA.t457 214.222
R4944 VDDA.t242 VDDA.n598 213.131
R4945 VDDA.n599 VDDA.t315 213.131
R4946 VDDA.t351 VDDA.n537 213.131
R4947 VDDA.n538 VDDA.t266 213.131
R4948 VDDA.t228 VDDA.n456 213.131
R4949 VDDA.n457 VDDA.t340 213.131
R4950 VDDA.n353 VDDA.n328 201.099
R4951 VDDA.n435 VDDA.t198 192.8
R4952 VDDA.n436 VDDA.t324 192.8
R4953 VDDA.n437 VDDA.t259 192.8
R4954 VDDA.n434 VDDA.t383 192.8
R4955 VDDA.n433 VDDA.t308 192.8
R4956 VDDA.n432 VDDA.t311 192.8
R4957 VDDA.n415 VDDA.t321 192.8
R4958 VDDA.n414 VDDA.t195 192.8
R4959 VDDA.n429 VDDA.t271 192.8
R4960 VDDA.n428 VDDA.t336 192.8
R4961 VDDA.n341 VDDA.n340 190.333
R4962 VDDA.n345 VDDA.n343 185
R4963 VDDA.n344 VDDA.n331 185
R4964 VDDA.n342 VDDA.n341 185
R4965 VDDA.n339 VDDA.n334 185
R4966 VDDA.n338 VDDA.n335 185
R4967 VDDA.n336 VDDA.n333 185
R4968 VDDA.n342 VDDA.n333 185
R4969 VDDA.n306 VDDA.t284 184.097
R4970 VDDA.n306 VDDA.t190 184.097
R4971 VDDA.n301 VDDA.t319 184.097
R4972 VDDA.n301 VDDA.t222 184.097
R4973 VDDA.n434 VDDA.n433 176.733
R4974 VDDA.n433 VDDA.n432 176.733
R4975 VDDA.n436 VDDA.n435 176.733
R4976 VDDA.n437 VDDA.n436 176.733
R4977 VDDA.n591 VDDA.t232 168.139
R4978 VDDA.n590 VDDA.t247 168.139
R4979 VDDA.n431 VDDA.n430 166.541
R4980 VDDA.n417 VDDA.n416 166.343
R4981 VDDA.n307 VDDA.n306 166.05
R4982 VDDA.n302 VDDA.n301 166.05
R4983 VDDA.n647 VDDA.n646 164.113
R4984 VDDA.n588 VDDA.n587 153.576
R4985 VDDA.n343 VDDA.n331 150
R4986 VDDA.n341 VDDA.n334 150
R4987 VDDA.n335 VDDA.n333 150
R4988 VDDA.t119 VDDA.t242 146.155
R4989 VDDA.t315 VDDA.t119 146.155
R4990 VDDA.t143 VDDA.t351 146.155
R4991 VDDA.t137 VDDA.t143 146.155
R4992 VDDA.t103 VDDA.t137 146.155
R4993 VDDA.t123 VDDA.t103 146.155
R4994 VDDA.t129 VDDA.t123 146.155
R4995 VDDA.t135 VDDA.t129 146.155
R4996 VDDA.t131 VDDA.t135 146.155
R4997 VDDA.t139 VDDA.t131 146.155
R4998 VDDA.t105 VDDA.t139 146.155
R4999 VDDA.t109 VDDA.t105 146.155
R5000 VDDA.t266 VDDA.t109 146.155
R5001 VDDA.t115 VDDA.t228 146.155
R5002 VDDA.t111 VDDA.t115 146.155
R5003 VDDA.t117 VDDA.t111 146.155
R5004 VDDA.t125 VDDA.t117 146.155
R5005 VDDA.t133 VDDA.t125 146.155
R5006 VDDA.t141 VDDA.t133 146.155
R5007 VDDA.t107 VDDA.t141 146.155
R5008 VDDA.t113 VDDA.t107 146.155
R5009 VDDA.t121 VDDA.t113 146.155
R5010 VDDA.t127 VDDA.t121 146.155
R5011 VDDA.t340 VDDA.t127 146.155
R5012 VDDA.n655 VDDA.t548 144.601
R5013 VDDA.n654 VDDA.t637 144.601
R5014 VDDA.n653 VDDA.t696 144.601
R5015 VDDA.n652 VDDA.t492 144.601
R5016 VDDA.n651 VDDA.t480 144.601
R5017 VDDA.n650 VDDA.t573 144.601
R5018 VDDA.n649 VDDA.t663 144.601
R5019 VDDA.n648 VDDA.t717 144.601
R5020 VDDA.n0 VDDA.t591 144.601
R5021 VDDA.n1 VDDA.t475 144.601
R5022 VDDA.n2 VDDA.t682 144.601
R5023 VDDA.n3 VDDA.t594 144.601
R5024 VDDA.n4 VDDA.t503 144.601
R5025 VDDA.n5 VDDA.t515 144.601
R5026 VDDA.n559 VDDA.t332 136.701
R5027 VDDA.n558 VDDA.t358 136.701
R5028 VDDA.n477 VDDA.t209 136.701
R5029 VDDA.n478 VDDA.t235 136.701
R5030 VDDA.n581 VDDA.t278 122.829
R5031 VDDA.t306 VDDA.n580 122.829
R5032 VDDA.t367 VDDA.n499 122.829
R5033 VDDA.n500 VDDA.t391 122.829
R5034 VDDA.n426 VDDA.t423 119.087
R5035 VDDA.n632 VDDA.t52 108.424
R5036 VDDA.n304 VDDA.t79 106.558
R5037 VDDA.n419 VDDA.t25 105.671
R5038 VDDA.n646 VDDA.t27 100.766
R5039 VDDA.t278 VDDA.t179 81.6411
R5040 VDDA.t179 VDDA.t157 81.6411
R5041 VDDA.t157 VDDA.t176 81.6411
R5042 VDDA.t176 VDDA.t166 81.6411
R5043 VDDA.t166 VDDA.t146 81.6411
R5044 VDDA.t146 VDDA.t163 81.6411
R5045 VDDA.t163 VDDA.t183 81.6411
R5046 VDDA.t183 VDDA.t160 81.6411
R5047 VDDA.t160 VDDA.t171 81.6411
R5048 VDDA.t171 VDDA.t150 81.6411
R5049 VDDA.t150 VDDA.t306 81.6411
R5050 VDDA.t403 VDDA.t367 81.6411
R5051 VDDA.t77 VDDA.t403 81.6411
R5052 VDDA.t89 VDDA.t77 81.6411
R5053 VDDA.t38 VDDA.t89 81.6411
R5054 VDDA.t409 VDDA.t38 81.6411
R5055 VDDA.t43 VDDA.t409 81.6411
R5056 VDDA.t401 VDDA.t43 81.6411
R5057 VDDA.t41 VDDA.t401 81.6411
R5058 VDDA.t399 VDDA.t41 81.6411
R5059 VDDA.t97 VDDA.t399 81.6411
R5060 VDDA.t391 VDDA.t97 81.6411
R5061 VDDA.n503 VDDA.t50 78.8005
R5062 VDDA.n503 VDDA.t7 78.8005
R5063 VDDA.n505 VDDA.t82 78.8005
R5064 VDDA.n505 VDDA.t18 78.8005
R5065 VDDA.n507 VDDA.t5 78.8005
R5066 VDDA.n507 VDDA.t63 78.8005
R5067 VDDA.n509 VDDA.t2 78.8005
R5068 VDDA.n509 VDDA.t22 78.8005
R5069 VDDA.n511 VDDA.t60 78.8005
R5070 VDDA.n511 VDDA.t84 78.8005
R5071 VDDA.n513 VDDA.t48 78.8005
R5072 VDDA.n513 VDDA.t20 78.8005
R5073 VDDA.n515 VDDA.t56 78.8005
R5074 VDDA.n515 VDDA.t75 78.8005
R5075 VDDA.n517 VDDA.t68 78.8005
R5076 VDDA.n517 VDDA.t418 78.8005
R5077 VDDA.n519 VDDA.t46 78.8005
R5078 VDDA.n519 VDDA.t70 78.8005
R5079 VDDA.n521 VDDA.t24 78.8005
R5080 VDDA.n521 VDDA.t31 78.8005
R5081 VDDA.n598 VDDA.t243 76.2576
R5082 VDDA.n599 VDDA.t316 76.2576
R5083 VDDA.n537 VDDA.t352 76.2576
R5084 VDDA.n538 VDDA.t267 76.2576
R5085 VDDA.n456 VDDA.t229 76.2576
R5086 VDDA.n457 VDDA.t341 76.2576
R5087 VDDA.n533 VDDA.n532 71.513
R5088 VDDA.n535 VDDA.n534 71.513
R5089 VDDA.n541 VDDA.n540 71.513
R5090 VDDA.n543 VDDA.n542 71.513
R5091 VDDA.n452 VDDA.n451 71.513
R5092 VDDA.n454 VDDA.n453 71.513
R5093 VDDA.n460 VDDA.n459 71.513
R5094 VDDA.n462 VDDA.n461 71.513
R5095 VDDA.n596 VDDA.n595 71.388
R5096 VDDA VDDA.n655 69.6227
R5097 VDDA.n648 VDDA.n647 69.6227
R5098 VDDA.n647 VDDA.n5 69.6227
R5099 VDDA.n545 VDDA.n531 67.013
R5100 VDDA.n464 VDDA.n450 67.013
R5101 VDDA.n348 VDDA.n347 65.8183
R5102 VDDA.n349 VDDA.n348 65.8183
R5103 VDDA.n342 VDDA.n332 65.8183
R5104 VDDA.n416 VDDA.n415 56.2338
R5105 VDDA.n416 VDDA.n414 56.2338
R5106 VDDA.n430 VDDA.n429 56.2338
R5107 VDDA.n430 VDDA.n428 56.2338
R5108 VDDA.n438 VDDA.n434 56.2338
R5109 VDDA.n438 VDDA.n437 56.2338
R5110 VDDA.n234 VDDA.t26 54.0032
R5111 VDDA.n347 VDDA.n343 53.3664
R5112 VDDA.n349 VDDA.n331 53.3664
R5113 VDDA.n334 VDDA.n332 53.3664
R5114 VDDA.n335 VDDA.n332 53.3664
R5115 VDDA.n234 VDDA.n233 45.6618
R5116 VDDA.n570 VDDA.n569 41.1393
R5117 VDDA.n572 VDDA.n571 41.1393
R5118 VDDA.n574 VDDA.n573 41.1393
R5119 VDDA.n576 VDDA.n575 41.1393
R5120 VDDA.n578 VDDA.n577 41.1393
R5121 VDDA.n489 VDDA.n488 41.1393
R5122 VDDA.n491 VDDA.n490 41.1393
R5123 VDDA.n493 VDDA.n492 41.1393
R5124 VDDA.n495 VDDA.n494 41.1393
R5125 VDDA.n497 VDDA.n496 41.1393
R5126 VDDA.n581 VDDA.t279 40.9789
R5127 VDDA.n580 VDDA.t307 40.9789
R5128 VDDA.n499 VDDA.t368 40.9789
R5129 VDDA.n500 VDDA.t392 40.9789
R5130 VDDA.n424 VDDA.t360 39.4005
R5131 VDDA.n424 VDDA.t71 39.4005
R5132 VDDA.n422 VDDA.t191 39.4005
R5133 VDDA.n422 VDDA.t285 39.4005
R5134 VDDA.n420 VDDA.t223 39.4005
R5135 VDDA.n420 VDDA.t320 39.4005
R5136 VDDA.n418 VDDA.t412 39.4005
R5137 VDDA.n418 VDDA.t370 39.4005
R5138 VDDA.n401 VDDA.t273 39.4005
R5139 VDDA.n401 VDDA.t203 39.4005
R5140 VDDA.n400 VDDA.t206 39.4005
R5141 VDDA.n400 VDDA.t338 39.4005
R5142 VDDA.n374 VDDA.t238 39.4005
R5143 VDDA.n374 VDDA.t388 39.4005
R5144 VDDA.n373 VDDA.t310 39.4005
R5145 VDDA.n373 VDDA.t313 39.4005
R5146 VDDA.n371 VDDA.t200 39.4005
R5147 VDDA.n371 VDDA.t326 39.4005
R5148 VDDA.n392 VDDA.t329 39.4005
R5149 VDDA.n392 VDDA.t264 39.4005
R5150 VDDA.n375 VDDA.t323 39.4005
R5151 VDDA.n375 VDDA.t253 39.4005
R5152 VDDA.n384 VDDA.t256 39.4005
R5153 VDDA.n384 VDDA.t197 39.4005
R5154 VDDA.n377 VDDA.t294 39.4005
R5155 VDDA.n377 VDDA.t221 39.4005
R5156 VDDA.n370 VDDA.t261 39.4005
R5157 VDDA.n370 VDDA.t385 39.4005
R5158 VDDA.n634 VDDA.t53 39.4005
R5159 VDDA.n634 VDDA.t29 39.4005
R5160 VDDA.n636 VDDA.t51 39.4005
R5161 VDDA.n636 VDDA.t3 39.4005
R5162 VDDA.n638 VDDA.t395 39.4005
R5163 VDDA.n638 VDDA.t397 39.4005
R5164 VDDA.n637 VDDA.t35 39.4005
R5165 VDDA.n637 VDDA.t393 39.4005
R5166 VDDA.n642 VDDA.t80 39.4005
R5167 VDDA.n642 VDDA.t411 39.4005
R5168 VDDA.n644 VDDA.t54 39.4005
R5169 VDDA.n644 VDDA.t416 39.4005
R5170 VDDA.n308 VDDA.t57 39.4005
R5171 VDDA.n308 VDDA.t419 39.4005
R5172 VDDA.n303 VDDA.t422 39.4005
R5173 VDDA.n303 VDDA.t93 39.4005
R5174 VDDA.n299 VDDA.t0 39.4005
R5175 VDDA.n299 VDDA.t32 39.4005
R5176 VDDA.n632 VDDA.n631 37.183
R5177 VDDA.n548 VDDA.n546 30.2255
R5178 VDDA.n467 VDDA.n465 30.2255
R5179 VDDA.n556 VDDA.n555 29.663
R5180 VDDA.n554 VDDA.n553 29.663
R5181 VDDA.n552 VDDA.n551 29.663
R5182 VDDA.n550 VDDA.n549 29.663
R5183 VDDA.n548 VDDA.n547 29.663
R5184 VDDA.n475 VDDA.n474 29.663
R5185 VDDA.n473 VDDA.n472 29.663
R5186 VDDA.n471 VDDA.n470 29.663
R5187 VDDA.n469 VDDA.n468 29.663
R5188 VDDA.n467 VDDA.n466 29.663
R5189 VDDA.n404 VDDA.n403 27.2462
R5190 VDDA.n402 VDDA.n399 27.2462
R5191 VDDA.n390 VDDA.n389 27.2462
R5192 VDDA.n388 VDDA.n387 27.2462
R5193 VDDA.n398 VDDA.n397 24.9931
R5194 VDDA.n396 VDDA.n395 24.9931
R5195 VDDA.n382 VDDA.n381 24.9931
R5196 VDDA.n380 VDDA.n379 24.9931
R5197 VDDA.n351 VDDA.n350 22.8576
R5198 VDDA.n336 VDDA.n329 22.8576
R5199 VDDA.n587 VDDA.t16 21.8894
R5200 VDDA.n587 VDDA.t246 21.8894
R5201 VDDA.n633 VDDA.n632 20.4706
R5202 VDDA.n298 VDDA.t218 20.1258
R5203 VDDA.n328 VDDA.t212 19.7005
R5204 VDDA.n328 VDDA.t346 19.7005
R5205 VDDA.n298 VDDA.n297 18.7759
R5206 VDDA.n235 VDDA.n234 17.3005
R5207 VDDA.n562 VDDA.n556 11.3443
R5208 VDDA.n481 VDDA.n475 11.3443
R5209 VDDA.t243 VDDA.n596 11.2576
R5210 VDDA.n596 VDDA.t120 11.2576
R5211 VDDA.n532 VDDA.t104 11.2576
R5212 VDDA.n532 VDDA.t124 11.2576
R5213 VDDA.n534 VDDA.t144 11.2576
R5214 VDDA.n534 VDDA.t138 11.2576
R5215 VDDA.n540 VDDA.t106 11.2576
R5216 VDDA.n540 VDDA.t110 11.2576
R5217 VDDA.n542 VDDA.t132 11.2576
R5218 VDDA.n542 VDDA.t140 11.2576
R5219 VDDA.n531 VDDA.t130 11.2576
R5220 VDDA.n531 VDDA.t136 11.2576
R5221 VDDA.n451 VDDA.t118 11.2576
R5222 VDDA.n451 VDDA.t126 11.2576
R5223 VDDA.n453 VDDA.t116 11.2576
R5224 VDDA.n453 VDDA.t112 11.2576
R5225 VDDA.n459 VDDA.t122 11.2576
R5226 VDDA.n459 VDDA.t128 11.2576
R5227 VDDA.n461 VDDA.t108 11.2576
R5228 VDDA.n461 VDDA.t114 11.2576
R5229 VDDA.n450 VDDA.t134 11.2576
R5230 VDDA.n450 VDDA.t142 11.2576
R5231 VDDA.n379 VDDA.n378 10.995
R5232 VDDA.n405 VDDA.n404 10.9846
R5233 VDDA.n352 VDDA.n329 10.9846
R5234 VDDA.n352 VDDA.n351 10.9325
R5235 VDDA.n431 VDDA.n427 10.871
R5236 VDDA.n407 VDDA.n399 10.87
R5237 VDDA.n395 VDDA.n394 10.87
R5238 VDDA.n387 VDDA.n386 10.87
R5239 VDDA.n383 VDDA.n382 10.87
R5240 VDDA.n391 VDDA.n390 10.87
R5241 VDDA.n408 VDDA.n398 10.87
R5242 VDDA.n603 VDDA.n602 9.7005
R5243 VDDA.n233 VDDA.t28 9.6005
R5244 VDDA.n233 VDDA.t61 9.6005
R5245 VDDA.n566 VDDA.n565 9.5505
R5246 VDDA.n564 VDDA.n563 9.5505
R5247 VDDA.n485 VDDA.n484 9.5505
R5248 VDDA.n483 VDDA.n482 9.5505
R5249 VDDA.n585 VDDA.n584 9.5005
R5250 VDDA.n530 VDDA.n529 9.5005
R5251 VDDA.n526 VDDA.n525 9.3005
R5252 VDDA.n524 VDDA.n523 9.3005
R5253 VDDA.n640 VDDA.n639 9.2505
R5254 VDDA.n311 VDDA.n310 9.2505
R5255 VDDA.n345 VDDA.n344 9.14336
R5256 VDDA.n339 VDDA.n338 9.14336
R5257 VDDA.n567 VDDA.n563 9.02133
R5258 VDDA.n486 VDDA.n482 9.02133
R5259 VDDA.n311 VDDA.n298 8.85883
R5260 VDDA.n561 VDDA.n557 8.79217
R5261 VDDA.n480 VDDA.n476 8.79217
R5262 VDDA.n555 VDDA.t100 8.0005
R5263 VDDA.n555 VDDA.t145 8.0005
R5264 VDDA.n553 VDDA.t162 8.0005
R5265 VDDA.n553 VDDA.t182 8.0005
R5266 VDDA.n551 VDDA.t174 8.0005
R5267 VDDA.n551 VDDA.t154 8.0005
R5268 VDDA.n549 VDDA.t170 8.0005
R5269 VDDA.n549 VDDA.t149 8.0005
R5270 VDDA.n547 VDDA.t165 8.0005
R5271 VDDA.n547 VDDA.t169 8.0005
R5272 VDDA.n546 VDDA.t153 8.0005
R5273 VDDA.n546 VDDA.t101 8.0005
R5274 VDDA.n474 VDDA.t40 8.0005
R5275 VDDA.n474 VDDA.t99 8.0005
R5276 VDDA.n472 VDDA.t8 8.0005
R5277 VDDA.n472 VDDA.t91 8.0005
R5278 VDDA.n470 VDDA.t9 8.0005
R5279 VDDA.n470 VDDA.t408 8.0005
R5280 VDDA.n468 VDDA.t73 8.0005
R5281 VDDA.n468 VDDA.t405 8.0005
R5282 VDDA.n466 VDDA.t87 8.0005
R5283 VDDA.n466 VDDA.t407 8.0005
R5284 VDDA.n465 VDDA.t102 8.0005
R5285 VDDA.n465 VDDA.t37 8.0005
R5286 VDDA.n585 VDDA.n545 7.71925
R5287 VDDA.n530 VDDA.n464 7.71925
R5288 VDDA.n586 VDDA.n530 6.90675
R5289 VDDA.n586 VDDA.n585 6.8755
R5290 VDDA.n594 VDDA.n586 6.813
R5291 VDDA.n569 VDDA.t180 6.56717
R5292 VDDA.n569 VDDA.t158 6.56717
R5293 VDDA.n571 VDDA.t177 6.56717
R5294 VDDA.n571 VDDA.t167 6.56717
R5295 VDDA.n573 VDDA.t147 6.56717
R5296 VDDA.n573 VDDA.t164 6.56717
R5297 VDDA.n575 VDDA.t184 6.56717
R5298 VDDA.n575 VDDA.t161 6.56717
R5299 VDDA.n577 VDDA.t172 6.56717
R5300 VDDA.n577 VDDA.t151 6.56717
R5301 VDDA.n488 VDDA.t400 6.56717
R5302 VDDA.n488 VDDA.t98 6.56717
R5303 VDDA.n490 VDDA.t402 6.56717
R5304 VDDA.n490 VDDA.t42 6.56717
R5305 VDDA.n492 VDDA.t410 6.56717
R5306 VDDA.n492 VDDA.t44 6.56717
R5307 VDDA.n494 VDDA.t90 6.56717
R5308 VDDA.n494 VDDA.t39 6.56717
R5309 VDDA.n496 VDDA.t404 6.56717
R5310 VDDA.n496 VDDA.t78 6.56717
R5311 VDDA.n426 VDDA.n425 6.15675
R5312 VDDA.n541 VDDA.n539 6.10467
R5313 VDDA.n536 VDDA.n535 6.10467
R5314 VDDA.n460 VDDA.n458 6.10467
R5315 VDDA.n455 VDDA.n454 6.10467
R5316 VDDA.n487 VDDA.n486 6.09425
R5317 VDDA.n568 VDDA.n567 6.063
R5318 VDDA.n312 VDDA.n311 5.98696
R5319 VDDA.n523 VDDA.n522 5.60467
R5320 VDDA.n350 VDDA.n330 5.33286
R5321 VDDA.n337 VDDA.n336 5.33286
R5322 VDDA.n579 VDDA.n578 5.313
R5323 VDDA.n498 VDDA.n497 5.313
R5324 VDDA.n602 VDDA.n601 5.28175
R5325 VDDA.n594 VDDA.n593 5.28175
R5326 VDDA.n584 VDDA.n583 5.28175
R5327 VDDA.n562 VDDA.n561 5.28175
R5328 VDDA.n481 VDDA.n480 5.28175
R5329 VDDA.n633 VDDA.n620 5.27699
R5330 VDDA.n646 VDDA.n645 5.188
R5331 VDDA.n527 VDDA.n526 5.04217
R5332 VDDA.n567 VDDA.n566 5.02133
R5333 VDDA.n486 VDDA.n485 5.02133
R5334 VDDA.n621 VDDA.t282 4.8295
R5335 VDDA.n622 VDDA.t364 4.8295
R5336 VDDA.n623 VDDA.t303 4.8295
R5337 VDDA.n624 VDDA.t213 4.8295
R5338 VDDA.n625 VDDA.t295 4.8295
R5339 VDDA.n626 VDDA.t374 4.8295
R5340 VDDA.n627 VDDA.t348 4.8295
R5341 VDDA.n628 VDDA.t215 4.8295
R5342 VDDA.n629 VDDA.t280 4.8295
R5343 VDDA.n287 VDDA.t513 4.8295
R5344 VDDA.n288 VDDA.t567 4.8295
R5345 VDDA.n289 VDDA.t723 4.8295
R5346 VDDA.n290 VDDA.t481 4.8295
R5347 VDDA.n291 VDDA.t501 4.8295
R5348 VDDA.n292 VDDA.t555 4.8295
R5349 VDDA.n293 VDDA.t712 4.8295
R5350 VDDA.n294 VDDA.t469 4.8295
R5351 VDDA.n295 VDDA.t684 4.8295
R5352 VDDA.n9 VDDA.t436 4.8295
R5353 VDDA.n13 VDDA.t430 4.8295
R5354 VDDA.n18 VDDA.t651 4.8295
R5355 VDDA.n22 VDDA.t642 4.8295
R5356 VDDA.n27 VDDA.t424 4.8295
R5357 VDDA.n31 VDDA.t720 4.8295
R5358 VDDA.n36 VDDA.t638 4.8295
R5359 VDDA.n40 VDDA.t632 4.8295
R5360 VDDA.n45 VDDA.t556 4.8295
R5361 VDDA.n49 VDDA.t549 4.8295
R5362 VDDA.n54 VDDA.t471 4.8295
R5363 VDDA.n58 VDDA.t463 4.8295
R5364 VDDA.n63 VDDA.t542 4.8295
R5365 VDDA.n67 VDDA.t536 4.8295
R5366 VDDA.n72 VDDA.t458 4.8295
R5367 VDDA.n76 VDDA.t451 4.8295
R5368 VDDA.n81 VDDA.t675 4.8295
R5369 VDDA.n85 VDDA.t669 4.8295
R5370 VDDA.n90 VDDA.t447 4.8295
R5371 VDDA.n94 VDDA.t442 4.8295
R5372 VDDA.n99 VDDA.t665 4.8295
R5373 VDDA.n103 VDDA.t656 4.8295
R5374 VDDA.n108 VDDA.t580 4.8295
R5375 VDDA.n112 VDDA.t574 4.8295
R5376 VDDA.n117 VDDA.t652 4.8295
R5377 VDDA.n121 VDDA.t644 4.8295
R5378 VDDA.n126 VDDA.t569 4.8295
R5379 VDDA.n130 VDDA.t560 4.8295
R5380 VDDA.n135 VDDA.t495 4.8295
R5381 VDDA.n139 VDDA.t490 4.8295
R5382 VDDA.n144 VDDA.t707 4.8295
R5383 VDDA.n148 VDDA.t703 4.8295
R5384 VDDA.n153 VDDA.t484 4.8295
R5385 VDDA.n157 VDDA.t479 4.8295
R5386 VDDA.n162 VDDA.t695 4.8295
R5387 VDDA.n166 VDDA.t691 4.8295
R5388 VDDA.n171 VDDA.t611 4.8295
R5389 VDDA.n175 VDDA.t608 4.8295
R5390 VDDA.n180 VDDA.t686 4.8295
R5391 VDDA.n184 VDDA.t681 4.8295
R5392 VDDA.n189 VDDA.t603 4.8295
R5393 VDDA.n193 VDDA.t599 4.8295
R5394 VDDA.n198 VDDA.t519 4.8295
R5395 VDDA.n202 VDDA.t512 4.8295
R5396 VDDA.n207 VDDA.t592 4.8295
R5397 VDDA.n211 VDDA.t588 4.8295
R5398 VDDA.n216 VDDA.t507 4.8295
R5399 VDDA.n561 VDDA.n560 4.79217
R5400 VDDA.n480 VDDA.n479 4.79217
R5401 VDDA.n597 VDDA.n595 4.7505
R5402 VDDA.n589 VDDA.n588 4.7505
R5403 VDDA.n583 VDDA.n582 4.7505
R5404 VDDA.n502 VDDA.n501 4.7505
R5405 VDDA.n439 VDDA 4.5005
R5406 VDDA.n601 VDDA.n600 4.5005
R5407 VDDA.n593 VDDA.n592 4.5005
R5408 VDDA.n545 VDDA.n544 4.5005
R5409 VDDA.n529 VDDA.n528 4.5005
R5410 VDDA.n464 VDDA.n463 4.5005
R5411 VDDA.n440 VDDA.n369 4.5005
R5412 VDDA.n443 VDDA.n441 4.5005
R5413 VDDA.n444 VDDA.n368 4.5005
R5414 VDDA.n448 VDDA.n447 4.5005
R5415 VDDA.n449 VDDA.n367 4.5005
R5416 VDDA.n604 VDDA.n603 4.5005
R5417 VDDA.n641 VDDA.n640 4.5005
R5418 VDDA.n621 VDDA.t239 4.5005
R5419 VDDA.n622 VDDA.t297 4.5005
R5420 VDDA.n623 VDDA.t317 4.5005
R5421 VDDA.n624 VDDA.t342 4.5005
R5422 VDDA.n625 VDDA.t257 4.5005
R5423 VDDA.n626 VDDA.t299 4.5005
R5424 VDDA.n627 VDDA.t301 4.5005
R5425 VDDA.n628 VDDA.t376 4.5005
R5426 VDDA.n631 VDDA.t188 4.5005
R5427 VDDA.n630 VDDA.t378 4.5005
R5428 VDDA.n629 VDDA.t217 4.5005
R5429 VDDA.n620 VDDA.n619 4.5005
R5430 VDDA.n7 VDDA.n6 4.5005
R5431 VDDA.n610 VDDA.n609 4.5005
R5432 VDDA.n614 VDDA.n613 4.5005
R5433 VDDA.n354 VDDA.n327 4.5005
R5434 VDDA.n357 VDDA.n355 4.5005
R5435 VDDA.n358 VDDA.n326 4.5005
R5436 VDDA.n362 VDDA.n361 4.5005
R5437 VDDA.n305 VDDA.n304 4.5005
R5438 VDDA.n287 VDDA.t427 4.5005
R5439 VDDA.n288 VDDA.t645 4.5005
R5440 VDDA.n289 VDDA.t640 4.5005
R5441 VDDA.n290 VDDA.t561 4.5005
R5442 VDDA.n291 VDDA.t715 4.5005
R5443 VDDA.n292 VDDA.t633 4.5005
R5444 VDDA.n293 VDDA.t628 4.5005
R5445 VDDA.n294 VDDA.t550 4.5005
R5446 VDDA.n297 VDDA.t625 4.5005
R5447 VDDA.n296 VDDA.t544 4.5005
R5448 VDDA.n295 VDDA.t464 4.5005
R5449 VDDA.n312 VDDA.n281 4.5005
R5450 VDDA.n315 VDDA.n313 4.5005
R5451 VDDA.n316 VDDA.n280 4.5005
R5452 VDDA.n320 VDDA.n319 4.5005
R5453 VDDA.n235 VDDA.n232 4.5005
R5454 VDDA.n238 VDDA.n236 4.5005
R5455 VDDA.n239 VDDA.n231 4.5005
R5456 VDDA.n243 VDDA.n242 4.5005
R5457 VDDA.n9 VDDA.t488 4.5005
R5458 VDDA.n10 VDDA.t526 4.5005
R5459 VDDA.n11 VDDA.t443 4.5005
R5460 VDDA.n12 VDDA.t664 4.5005
R5461 VDDA.n17 VDDA.t708 4.5005
R5462 VDDA.n16 VDDA.t626 4.5005
R5463 VDDA.n15 VDDA.t545 4.5005
R5464 VDDA.n14 VDDA.t598 4.5005
R5465 VDDA.n13 VDDA.t516 4.5005
R5466 VDDA.n18 VDDA.t700 4.5005
R5467 VDDA.n19 VDDA.t438 4.5005
R5468 VDDA.n20 VDDA.t658 4.5005
R5469 VDDA.n21 VDDA.t577 4.5005
R5470 VDDA.n26 VDDA.t620 4.5005
R5471 VDDA.n25 VDDA.t540 4.5005
R5472 VDDA.n24 VDDA.t459 4.5005
R5473 VDDA.n23 VDDA.t510 4.5005
R5474 VDDA.n22 VDDA.t425 4.5005
R5475 VDDA.n27 VDDA.t476 4.5005
R5476 VDDA.n28 VDDA.t517 4.5005
R5477 VDDA.n29 VDDA.t432 4.5005
R5478 VDDA.n30 VDDA.t650 4.5005
R5479 VDDA.n35 VDDA.t697 4.5005
R5480 VDDA.n34 VDDA.t616 4.5005
R5481 VDDA.n33 VDDA.t535 4.5005
R5482 VDDA.n32 VDDA.t585 4.5005
R5483 VDDA.n31 VDDA.t505 4.5005
R5484 VDDA.n36 VDDA.t690 4.5005
R5485 VDDA.n37 VDDA.t428 4.5005
R5486 VDDA.n38 VDDA.t646 4.5005
R5487 VDDA.n39 VDDA.t568 4.5005
R5488 VDDA.n44 VDDA.t612 4.5005
R5489 VDDA.n43 VDDA.t531 4.5005
R5490 VDDA.n42 VDDA.t450 4.5005
R5491 VDDA.n41 VDDA.t499 4.5005
R5492 VDDA.n40 VDDA.t714 4.5005
R5493 VDDA.n45 VDDA.t605 4.5005
R5494 VDDA.n46 VDDA.t641 4.5005
R5495 VDDA.n47 VDDA.t562 4.5005
R5496 VDDA.n48 VDDA.t483 4.5005
R5497 VDDA.n53 VDDA.t528 4.5005
R5498 VDDA.n52 VDDA.t445 4.5005
R5499 VDDA.n51 VDDA.t668 4.5005
R5500 VDDA.n50 VDDA.t711 4.5005
R5501 VDDA.n49 VDDA.t627 4.5005
R5502 VDDA.n54 VDDA.t520 4.5005
R5503 VDDA.n55 VDDA.t557 4.5005
R5504 VDDA.n56 VDDA.t477 4.5005
R5505 VDDA.n57 VDDA.t694 4.5005
R5506 VDDA.n62 VDDA.t441 4.5005
R5507 VDDA.n61 VDDA.t661 4.5005
R5508 VDDA.n60 VDDA.t583 4.5005
R5509 VDDA.n59 VDDA.t624 4.5005
R5510 VDDA.n58 VDDA.t543 4.5005
R5511 VDDA.n63 VDDA.t597 4.5005
R5512 VDDA.n64 VDDA.t629 4.5005
R5513 VDDA.n65 VDDA.t551 4.5005
R5514 VDDA.n66 VDDA.t470 4.5005
R5515 VDDA.n71 VDDA.t521 4.5005
R5516 VDDA.n70 VDDA.t435 4.5005
R5517 VDDA.n69 VDDA.t654 4.5005
R5518 VDDA.n68 VDDA.t702 4.5005
R5519 VDDA.n67 VDDA.t618 4.5005
R5520 VDDA.n72 VDDA.t509 4.5005
R5521 VDDA.n73 VDDA.t546 4.5005
R5522 VDDA.n74 VDDA.t466 4.5005
R5523 VDDA.n75 VDDA.t685 4.5005
R5524 VDDA.n80 VDDA.t431 4.5005
R5525 VDDA.n79 VDDA.t649 4.5005
R5526 VDDA.n78 VDDA.t570 4.5005
R5527 VDDA.n77 VDDA.t615 4.5005
R5528 VDDA.n76 VDDA.t532 4.5005
R5529 VDDA.n81 VDDA.t721 4.5005
R5530 VDDA.n82 VDDA.t460 4.5005
R5531 VDDA.n83 VDDA.t680 4.5005
R5532 VDDA.n84 VDDA.t602 4.5005
R5533 VDDA.n89 VDDA.t643 4.5005
R5534 VDDA.n88 VDDA.t566 4.5005
R5535 VDDA.n87 VDDA.t485 4.5005
R5536 VDDA.n86 VDDA.t530 4.5005
R5537 VDDA.n85 VDDA.t448 4.5005
R5538 VDDA.n90 VDDA.t498 4.5005
R5539 VDDA.n91 VDDA.t533 4.5005
R5540 VDDA.n92 VDDA.t452 4.5005
R5541 VDDA.n93 VDDA.t674 4.5005
R5542 VDDA.n98 VDDA.t718 4.5005
R5543 VDDA.n97 VDDA.t636 4.5005
R5544 VDDA.n96 VDDA.t559 4.5005
R5545 VDDA.n95 VDDA.t607 4.5005
R5546 VDDA.n94 VDDA.t525 4.5005
R5547 VDDA.n99 VDDA.t710 4.5005
R5548 VDDA.n100 VDDA.t449 4.5005
R5549 VDDA.n101 VDDA.t670 4.5005
R5550 VDDA.n102 VDDA.t590 4.5005
R5551 VDDA.n107 VDDA.t631 4.5005
R5552 VDDA.n106 VDDA.t554 4.5005
R5553 VDDA.n105 VDDA.t473 4.5005
R5554 VDDA.n104 VDDA.t523 4.5005
R5555 VDDA.n103 VDDA.t437 4.5005
R5556 VDDA.n108 VDDA.t623 4.5005
R5557 VDDA.n109 VDDA.t666 4.5005
R5558 VDDA.n110 VDDA.t586 4.5005
R5559 VDDA.n111 VDDA.t506 4.5005
R5560 VDDA.n116 VDDA.t547 4.5005
R5561 VDDA.n115 VDDA.t468 4.5005
R5562 VDDA.n114 VDDA.t688 4.5005
R5563 VDDA.n113 VDDA.t434 4.5005
R5564 VDDA.n112 VDDA.t653 4.5005
R5565 VDDA.n117 VDDA.t701 4.5005
R5566 VDDA.n118 VDDA.t439 4.5005
R5567 VDDA.n119 VDDA.t659 4.5005
R5568 VDDA.n120 VDDA.t578 4.5005
R5569 VDDA.n125 VDDA.t621 4.5005
R5570 VDDA.n124 VDDA.t541 4.5005
R5571 VDDA.n123 VDDA.t461 4.5005
R5572 VDDA.n122 VDDA.t511 4.5005
R5573 VDDA.n121 VDDA.t426 4.5005
R5574 VDDA.n126 VDDA.t614 4.5005
R5575 VDDA.n127 VDDA.t655 4.5005
R5576 VDDA.n128 VDDA.t576 4.5005
R5577 VDDA.n129 VDDA.t493 4.5005
R5578 VDDA.n134 VDDA.t537 4.5005
R5579 VDDA.n133 VDDA.t456 4.5005
R5580 VDDA.n132 VDDA.t676 4.5005
R5581 VDDA.n131 VDDA.t722 4.5005
R5582 VDDA.n130 VDDA.t639 4.5005
R5583 VDDA.n135 VDDA.t538 4.5005
R5584 VDDA.n136 VDDA.t584 4.5005
R5585 VDDA.n137 VDDA.t502 4.5005
R5586 VDDA.n138 VDDA.t716 4.5005
R5587 VDDA.n143 VDDA.t465 4.5005
R5588 VDDA.n142 VDDA.t683 4.5005
R5589 VDDA.n141 VDDA.t606 4.5005
R5590 VDDA.n140 VDDA.t648 4.5005
R5591 VDDA.n139 VDDA.t571 4.5005
R5592 VDDA.n144 VDDA.t454 4.5005
R5593 VDDA.n145 VDDA.t496 4.5005
R5594 VDDA.n146 VDDA.t713 4.5005
R5595 VDDA.n147 VDDA.t630 4.5005
R5596 VDDA.n152 VDDA.t679 4.5005
R5597 VDDA.n151 VDDA.t601 4.5005
R5598 VDDA.n150 VDDA.t522 4.5005
R5599 VDDA.n149 VDDA.t565 4.5005
R5600 VDDA.n148 VDDA.t486 4.5005
R5601 VDDA.n153 VDDA.t529 4.5005
R5602 VDDA.n154 VDDA.t572 4.5005
R5603 VDDA.n155 VDDA.t491 4.5005
R5604 VDDA.n156 VDDA.t706 4.5005
R5605 VDDA.n161 VDDA.t453 4.5005
R5606 VDDA.n160 VDDA.t673 4.5005
R5607 VDDA.n159 VDDA.t596 4.5005
R5608 VDDA.n158 VDDA.t635 4.5005
R5609 VDDA.n157 VDDA.t558 4.5005
R5610 VDDA.n162 VDDA.t444 4.5005
R5611 VDDA.n163 VDDA.t487 4.5005
R5612 VDDA.n164 VDDA.t704 4.5005
R5613 VDDA.n165 VDDA.t619 4.5005
R5614 VDDA.n170 VDDA.t671 4.5005
R5615 VDDA.n169 VDDA.t589 4.5005
R5616 VDDA.n168 VDDA.t508 4.5005
R5617 VDDA.n167 VDDA.t553 4.5005
R5618 VDDA.n166 VDDA.t472 4.5005
R5619 VDDA.n171 VDDA.t660 4.5005
R5620 VDDA.n172 VDDA.t699 4.5005
R5621 VDDA.n173 VDDA.t617 4.5005
R5622 VDDA.n174 VDDA.t534 4.5005
R5623 VDDA.n179 VDDA.t587 4.5005
R5624 VDDA.n178 VDDA.t504 4.5005
R5625 VDDA.n177 VDDA.t719 4.5005
R5626 VDDA.n176 VDDA.t467 4.5005
R5627 VDDA.n175 VDDA.t687 4.5005
R5628 VDDA.n180 VDDA.t433 4.5005
R5629 VDDA.n181 VDDA.t474 4.5005
R5630 VDDA.n182 VDDA.t692 4.5005
R5631 VDDA.n183 VDDA.t610 4.5005
R5632 VDDA.n188 VDDA.t657 4.5005
R5633 VDDA.n187 VDDA.t579 4.5005
R5634 VDDA.n186 VDDA.t497 4.5005
R5635 VDDA.n185 VDDA.t539 4.5005
R5636 VDDA.n184 VDDA.t462 4.5005
R5637 VDDA.n189 VDDA.t647 4.5005
R5638 VDDA.n190 VDDA.t689 4.5005
R5639 VDDA.n191 VDDA.t609 4.5005
R5640 VDDA.n192 VDDA.t527 4.5005
R5641 VDDA.n197 VDDA.t575 4.5005
R5642 VDDA.n196 VDDA.t494 4.5005
R5643 VDDA.n195 VDDA.t709 4.5005
R5644 VDDA.n194 VDDA.t455 4.5005
R5645 VDDA.n193 VDDA.t677 4.5005
R5646 VDDA.n198 VDDA.t564 4.5005
R5647 VDDA.n199 VDDA.t604 4.5005
R5648 VDDA.n200 VDDA.t524 4.5005
R5649 VDDA.n201 VDDA.t440 4.5005
R5650 VDDA.n206 VDDA.t489 4.5005
R5651 VDDA.n205 VDDA.t705 4.5005
R5652 VDDA.n204 VDDA.t622 4.5005
R5653 VDDA.n203 VDDA.t672 4.5005
R5654 VDDA.n202 VDDA.t593 4.5005
R5655 VDDA.n207 VDDA.t634 4.5005
R5656 VDDA.n208 VDDA.t678 4.5005
R5657 VDDA.n209 VDDA.t600 4.5005
R5658 VDDA.n210 VDDA.t518 4.5005
R5659 VDDA.n215 VDDA.t563 4.5005
R5660 VDDA.n214 VDDA.t482 4.5005
R5661 VDDA.n213 VDDA.t698 4.5005
R5662 VDDA.n212 VDDA.t446 4.5005
R5663 VDDA.n211 VDDA.t667 4.5005
R5664 VDDA.n216 VDDA.t552 4.5005
R5665 VDDA.n217 VDDA.t595 4.5005
R5666 VDDA.n218 VDDA.t514 4.5005
R5667 VDDA.n219 VDDA.t429 4.5005
R5668 VDDA.n220 VDDA.t478 4.5005
R5669 VDDA.n221 VDDA.t693 4.5005
R5670 VDDA.n222 VDDA.t613 4.5005
R5671 VDDA.n223 VDDA.t662 4.5005
R5672 VDDA.n224 VDDA.t582 4.5005
R5673 VDDA.n225 VDDA.t500 4.5005
R5674 VDDA.n584 VDDA.n568 3.84425
R5675 VDDA.n529 VDDA.n487 3.84425
R5676 VDDA.n346 VDDA.n345 3.75335
R5677 VDDA.n344 VDDA.n330 3.75335
R5678 VDDA.n340 VDDA.n339 3.75335
R5679 VDDA.n338 VDDA.n337 3.75335
R5680 VDDA.n635 VDDA.n633 3.7212
R5681 VDDA.n616 VDDA.n615 3.47871
R5682 VDDA.n364 VDDA.n363 3.47871
R5683 VDDA.n322 VDDA.n321 3.47871
R5684 VDDA.n245 VDDA.n244 3.47871
R5685 VDDA.n367 VDDA.n366 3.4105
R5686 VDDA.n447 VDDA.n446 3.4105
R5687 VDDA.n445 VDDA.n444 3.4105
R5688 VDDA.n443 VDDA.n442 3.4105
R5689 VDDA.n369 VDDA.n249 3.4105
R5690 VDDA.n605 VDDA.n604 3.4105
R5691 VDDA.n608 VDDA.n607 3.4105
R5692 VDDA.n613 VDDA.n612 3.4105
R5693 VDDA.n611 VDDA.n610 3.4105
R5694 VDDA.n8 VDDA.n7 3.4105
R5695 VDDA.n619 VDDA.n618 3.4105
R5696 VDDA.n325 VDDA.n324 3.4105
R5697 VDDA.n361 VDDA.n360 3.4105
R5698 VDDA.n359 VDDA.n358 3.4105
R5699 VDDA.n357 VDDA.n356 3.4105
R5700 VDDA.n327 VDDA.n252 3.4105
R5701 VDDA.n279 VDDA.n278 3.4105
R5702 VDDA.n319 VDDA.n318 3.4105
R5703 VDDA.n317 VDDA.n316 3.4105
R5704 VDDA.n315 VDDA.n314 3.4105
R5705 VDDA.n281 VDDA.n255 3.4105
R5706 VDDA.n230 VDDA.n229 3.4105
R5707 VDDA.n242 VDDA.n241 3.4105
R5708 VDDA.n240 VDDA.n239 3.4105
R5709 VDDA.n238 VDDA.n237 3.4105
R5710 VDDA.n232 VDDA.n226 3.4105
R5711 VDDA.n246 VDDA.n226 3.4105
R5712 VDDA.n246 VDDA.n245 3.4105
R5713 VDDA.n323 VDDA.n255 3.4105
R5714 VDDA.n323 VDDA.n322 3.4105
R5715 VDDA.n365 VDDA.n252 3.4105
R5716 VDDA.n365 VDDA.n364 3.4105
R5717 VDDA.n618 VDDA.n617 3.4105
R5718 VDDA.n617 VDDA.n616 3.4105
R5719 VDDA.n606 VDDA.n249 3.4105
R5720 VDDA.n606 VDDA.n605 3.4105
R5721 VDDA.n269 VDDA.n259 3.4105
R5722 VDDA.n275 VDDA.n259 3.4105
R5723 VDDA.n277 VDDA.n259 3.4105
R5724 VDDA.n267 VDDA.n262 3.4105
R5725 VDDA.n277 VDDA.n262 3.4105
R5726 VDDA.n267 VDDA.n258 3.4105
R5727 VDDA.n265 VDDA.n258 3.4105
R5728 VDDA.n273 VDDA.n258 3.4105
R5729 VDDA.n264 VDDA.n258 3.4105
R5730 VDDA.n275 VDDA.n258 3.4105
R5731 VDDA.n277 VDDA.n258 3.4105
R5732 VDDA.n276 VDDA.n265 3.4105
R5733 VDDA.n276 VDDA.n273 3.4105
R5734 VDDA.n276 VDDA.n264 3.4105
R5735 VDDA.n276 VDDA.n275 3.4105
R5736 VDDA.n277 VDDA.n276 3.4105
R5737 VDDA.n528 VDDA.n527 3.1255
R5738 VDDA.n592 VDDA.n591 2.8255
R5739 VDDA.n590 VDDA.n589 2.8255
R5740 VDDA.n354 VDDA.n353 2.52468
R5741 VDDA.n560 VDDA.n559 2.423
R5742 VDDA.n558 VDDA.n557 2.423
R5743 VDDA.n479 VDDA.n478 2.423
R5744 VDDA.n477 VDDA.n476 2.423
R5745 VDDA.n615 VDDA.n614 2.39683
R5746 VDDA.n363 VDDA.n362 2.39683
R5747 VDDA.n321 VDDA.n320 2.39683
R5748 VDDA.n244 VDDA.n243 2.39683
R5749 VDDA VDDA.n431 2.29514
R5750 VDDA VDDA.n417 2.28175
R5751 VDDA.n645 VDDA.n643 2.1255
R5752 VDDA.n643 VDDA.n641 2.1255
R5753 VDDA.n641 VDDA.n635 2.1255
R5754 VDDA.n582 VDDA.n581 1.97758
R5755 VDDA.n580 VDDA.n579 1.97758
R5756 VDDA.n501 VDDA.n500 1.97758
R5757 VDDA.n499 VDDA.n498 1.97758
R5758 VDDA.n600 VDDA.n599 1.888
R5759 VDDA.n598 VDDA.n597 1.888
R5760 VDDA.n261 VDDA.n260 1.70468
R5761 VDDA.n263 VDDA.n260 1.70468
R5762 VDDA.n269 VDDA.n268 1.70453
R5763 VDDA.n266 VDDA.n259 1.70321
R5764 VDDA.n276 VDDA.n270 1.70321
R5765 VDDA.n271 VDDA.n259 1.70307
R5766 VDDA.n272 VDDA.n262 1.70307
R5767 VDDA.n274 VDDA.n262 1.70307
R5768 VDDA.n246 VDDA.n228 1.6924
R5769 VDDA.n246 VDDA.n227 1.6924
R5770 VDDA.n323 VDDA.n257 1.6924
R5771 VDDA.n323 VDDA.n256 1.6924
R5772 VDDA.n365 VDDA.n254 1.6924
R5773 VDDA.n365 VDDA.n253 1.6924
R5774 VDDA.n617 VDDA.n248 1.6924
R5775 VDDA.n617 VDDA.n247 1.6924
R5776 VDDA.n606 VDDA.n251 1.68971
R5777 VDDA.n606 VDDA.n250 1.68971
R5778 VDDA.n427 VDDA.n426 1.59425
R5779 VDDA.n353 VDDA.n352 1.45302
R5780 VDDA.n412 VDDA.n411 1.44719
R5781 VDDA.n568 VDDA.n562 1.438
R5782 VDDA.n487 VDDA.n481 1.438
R5783 VDDA.n302 VDDA.n300 1.3755
R5784 VDDA.n307 VDDA.n305 1.3755
R5785 VDDA.n310 VDDA.n309 1.188
R5786 VDDA.n421 VDDA.n419 1.1255
R5787 VDDA.n423 VDDA.n421 1.1255
R5788 VDDA.n425 VDDA.n423 1.1255
R5789 VDDA.n539 VDDA.n538 1.03383
R5790 VDDA.n537 VDDA.n536 1.03383
R5791 VDDA.n458 VDDA.n457 1.03383
R5792 VDDA.n456 VDDA.n455 1.03383
R5793 VDDA.n602 VDDA.n594 0.938
R5794 VDDA.n440 VDDA.n439 0.809875
R5795 VDDA.n528 VDDA.n502 0.78175
R5796 VDDA.n601 VDDA.n595 0.6255
R5797 VDDA.n593 VDDA.n588 0.6255
R5798 VDDA.n544 VDDA.n543 0.6255
R5799 VDDA.n543 VDDA.n541 0.6255
R5800 VDDA.n535 VDDA.n533 0.6255
R5801 VDDA.n544 VDDA.n533 0.6255
R5802 VDDA.n463 VDDA.n462 0.6255
R5803 VDDA.n462 VDDA.n460 0.6255
R5804 VDDA.n454 VDDA.n452 0.6255
R5805 VDDA.n463 VDDA.n452 0.6255
R5806 VDDA.n305 VDDA.n302 0.6255
R5807 VDDA.n309 VDDA.n307 0.6255
R5808 VDDA.n578 VDDA.n576 0.563
R5809 VDDA.n576 VDDA.n574 0.563
R5810 VDDA.n574 VDDA.n572 0.563
R5811 VDDA.n572 VDDA.n570 0.563
R5812 VDDA.n583 VDDA.n570 0.563
R5813 VDDA.n550 VDDA.n548 0.563
R5814 VDDA.n552 VDDA.n550 0.563
R5815 VDDA.n554 VDDA.n552 0.563
R5816 VDDA.n556 VDDA.n554 0.563
R5817 VDDA.n522 VDDA.n520 0.563
R5818 VDDA.n520 VDDA.n518 0.563
R5819 VDDA.n518 VDDA.n516 0.563
R5820 VDDA.n516 VDDA.n514 0.563
R5821 VDDA.n514 VDDA.n512 0.563
R5822 VDDA.n512 VDDA.n510 0.563
R5823 VDDA.n510 VDDA.n508 0.563
R5824 VDDA.n508 VDDA.n506 0.563
R5825 VDDA.n506 VDDA.n504 0.563
R5826 VDDA.n527 VDDA.n504 0.563
R5827 VDDA.n497 VDDA.n495 0.563
R5828 VDDA.n495 VDDA.n493 0.563
R5829 VDDA.n493 VDDA.n491 0.563
R5830 VDDA.n491 VDDA.n489 0.563
R5831 VDDA.n502 VDDA.n489 0.563
R5832 VDDA.n469 VDDA.n467 0.563
R5833 VDDA.n471 VDDA.n469 0.563
R5834 VDDA.n473 VDDA.n471 0.563
R5835 VDDA.n475 VDDA.n473 0.563
R5836 VDDA.n323 VDDA.n277 0.482838
R5837 VDDA.n622 VDDA.n621 0.3295
R5838 VDDA.n624 VDDA.n623 0.3295
R5839 VDDA.n626 VDDA.n625 0.3295
R5840 VDDA.n628 VDDA.n627 0.3295
R5841 VDDA.n631 VDDA.n630 0.3295
R5842 VDDA.n630 VDDA.n629 0.3295
R5843 VDDA.n288 VDDA.n287 0.3295
R5844 VDDA.n290 VDDA.n289 0.3295
R5845 VDDA.n292 VDDA.n291 0.3295
R5846 VDDA.n294 VDDA.n293 0.3295
R5847 VDDA.n297 VDDA.n296 0.3295
R5848 VDDA.n296 VDDA.n295 0.3295
R5849 VDDA.n10 VDDA.n9 0.3295
R5850 VDDA.n11 VDDA.n10 0.3295
R5851 VDDA.n12 VDDA.n11 0.3295
R5852 VDDA.n17 VDDA.n12 0.3295
R5853 VDDA.n17 VDDA.n16 0.3295
R5854 VDDA.n16 VDDA.n15 0.3295
R5855 VDDA.n15 VDDA.n14 0.3295
R5856 VDDA.n14 VDDA.n13 0.3295
R5857 VDDA.n19 VDDA.n18 0.3295
R5858 VDDA.n20 VDDA.n19 0.3295
R5859 VDDA.n21 VDDA.n20 0.3295
R5860 VDDA.n26 VDDA.n21 0.3295
R5861 VDDA.n26 VDDA.n25 0.3295
R5862 VDDA.n25 VDDA.n24 0.3295
R5863 VDDA.n24 VDDA.n23 0.3295
R5864 VDDA.n23 VDDA.n22 0.3295
R5865 VDDA.n28 VDDA.n27 0.3295
R5866 VDDA.n29 VDDA.n28 0.3295
R5867 VDDA.n30 VDDA.n29 0.3295
R5868 VDDA.n35 VDDA.n30 0.3295
R5869 VDDA.n35 VDDA.n34 0.3295
R5870 VDDA.n34 VDDA.n33 0.3295
R5871 VDDA.n33 VDDA.n32 0.3295
R5872 VDDA.n32 VDDA.n31 0.3295
R5873 VDDA.n37 VDDA.n36 0.3295
R5874 VDDA.n38 VDDA.n37 0.3295
R5875 VDDA.n39 VDDA.n38 0.3295
R5876 VDDA.n44 VDDA.n39 0.3295
R5877 VDDA.n44 VDDA.n43 0.3295
R5878 VDDA.n43 VDDA.n42 0.3295
R5879 VDDA.n42 VDDA.n41 0.3295
R5880 VDDA.n41 VDDA.n40 0.3295
R5881 VDDA.n46 VDDA.n45 0.3295
R5882 VDDA.n47 VDDA.n46 0.3295
R5883 VDDA.n48 VDDA.n47 0.3295
R5884 VDDA.n53 VDDA.n48 0.3295
R5885 VDDA.n53 VDDA.n52 0.3295
R5886 VDDA.n52 VDDA.n51 0.3295
R5887 VDDA.n51 VDDA.n50 0.3295
R5888 VDDA.n50 VDDA.n49 0.3295
R5889 VDDA.n55 VDDA.n54 0.3295
R5890 VDDA.n56 VDDA.n55 0.3295
R5891 VDDA.n57 VDDA.n56 0.3295
R5892 VDDA.n62 VDDA.n57 0.3295
R5893 VDDA.n62 VDDA.n61 0.3295
R5894 VDDA.n61 VDDA.n60 0.3295
R5895 VDDA.n60 VDDA.n59 0.3295
R5896 VDDA.n59 VDDA.n58 0.3295
R5897 VDDA.n64 VDDA.n63 0.3295
R5898 VDDA.n65 VDDA.n64 0.3295
R5899 VDDA.n66 VDDA.n65 0.3295
R5900 VDDA.n71 VDDA.n66 0.3295
R5901 VDDA.n71 VDDA.n70 0.3295
R5902 VDDA.n70 VDDA.n69 0.3295
R5903 VDDA.n69 VDDA.n68 0.3295
R5904 VDDA.n68 VDDA.n67 0.3295
R5905 VDDA.n73 VDDA.n72 0.3295
R5906 VDDA.n74 VDDA.n73 0.3295
R5907 VDDA.n75 VDDA.n74 0.3295
R5908 VDDA.n80 VDDA.n75 0.3295
R5909 VDDA.n80 VDDA.n79 0.3295
R5910 VDDA.n79 VDDA.n78 0.3295
R5911 VDDA.n78 VDDA.n77 0.3295
R5912 VDDA.n77 VDDA.n76 0.3295
R5913 VDDA.n82 VDDA.n81 0.3295
R5914 VDDA.n83 VDDA.n82 0.3295
R5915 VDDA.n84 VDDA.n83 0.3295
R5916 VDDA.n89 VDDA.n84 0.3295
R5917 VDDA.n89 VDDA.n88 0.3295
R5918 VDDA.n88 VDDA.n87 0.3295
R5919 VDDA.n87 VDDA.n86 0.3295
R5920 VDDA.n86 VDDA.n85 0.3295
R5921 VDDA.n91 VDDA.n90 0.3295
R5922 VDDA.n92 VDDA.n91 0.3295
R5923 VDDA.n93 VDDA.n92 0.3295
R5924 VDDA.n98 VDDA.n93 0.3295
R5925 VDDA.n98 VDDA.n97 0.3295
R5926 VDDA.n97 VDDA.n96 0.3295
R5927 VDDA.n96 VDDA.n95 0.3295
R5928 VDDA.n95 VDDA.n94 0.3295
R5929 VDDA.n100 VDDA.n99 0.3295
R5930 VDDA.n101 VDDA.n100 0.3295
R5931 VDDA.n102 VDDA.n101 0.3295
R5932 VDDA.n107 VDDA.n102 0.3295
R5933 VDDA.n107 VDDA.n106 0.3295
R5934 VDDA.n106 VDDA.n105 0.3295
R5935 VDDA.n105 VDDA.n104 0.3295
R5936 VDDA.n104 VDDA.n103 0.3295
R5937 VDDA.n109 VDDA.n108 0.3295
R5938 VDDA.n110 VDDA.n109 0.3295
R5939 VDDA.n111 VDDA.n110 0.3295
R5940 VDDA.n116 VDDA.n111 0.3295
R5941 VDDA.n116 VDDA.n115 0.3295
R5942 VDDA.n115 VDDA.n114 0.3295
R5943 VDDA.n114 VDDA.n113 0.3295
R5944 VDDA.n113 VDDA.n112 0.3295
R5945 VDDA.n118 VDDA.n117 0.3295
R5946 VDDA.n119 VDDA.n118 0.3295
R5947 VDDA.n120 VDDA.n119 0.3295
R5948 VDDA.n125 VDDA.n120 0.3295
R5949 VDDA.n125 VDDA.n124 0.3295
R5950 VDDA.n124 VDDA.n123 0.3295
R5951 VDDA.n123 VDDA.n122 0.3295
R5952 VDDA.n122 VDDA.n121 0.3295
R5953 VDDA.n127 VDDA.n126 0.3295
R5954 VDDA.n128 VDDA.n127 0.3295
R5955 VDDA.n129 VDDA.n128 0.3295
R5956 VDDA.n134 VDDA.n129 0.3295
R5957 VDDA.n134 VDDA.n133 0.3295
R5958 VDDA.n133 VDDA.n132 0.3295
R5959 VDDA.n132 VDDA.n131 0.3295
R5960 VDDA.n131 VDDA.n130 0.3295
R5961 VDDA.n136 VDDA.n135 0.3295
R5962 VDDA.n137 VDDA.n136 0.3295
R5963 VDDA.n138 VDDA.n137 0.3295
R5964 VDDA.n143 VDDA.n138 0.3295
R5965 VDDA.n143 VDDA.n142 0.3295
R5966 VDDA.n142 VDDA.n141 0.3295
R5967 VDDA.n141 VDDA.n140 0.3295
R5968 VDDA.n140 VDDA.n139 0.3295
R5969 VDDA.n145 VDDA.n144 0.3295
R5970 VDDA.n146 VDDA.n145 0.3295
R5971 VDDA.n147 VDDA.n146 0.3295
R5972 VDDA.n152 VDDA.n147 0.3295
R5973 VDDA.n152 VDDA.n151 0.3295
R5974 VDDA.n151 VDDA.n150 0.3295
R5975 VDDA.n150 VDDA.n149 0.3295
R5976 VDDA.n149 VDDA.n148 0.3295
R5977 VDDA.n154 VDDA.n153 0.3295
R5978 VDDA.n155 VDDA.n154 0.3295
R5979 VDDA.n156 VDDA.n155 0.3295
R5980 VDDA.n161 VDDA.n156 0.3295
R5981 VDDA.n161 VDDA.n160 0.3295
R5982 VDDA.n160 VDDA.n159 0.3295
R5983 VDDA.n159 VDDA.n158 0.3295
R5984 VDDA.n158 VDDA.n157 0.3295
R5985 VDDA.n163 VDDA.n162 0.3295
R5986 VDDA.n164 VDDA.n163 0.3295
R5987 VDDA.n165 VDDA.n164 0.3295
R5988 VDDA.n170 VDDA.n165 0.3295
R5989 VDDA.n170 VDDA.n169 0.3295
R5990 VDDA.n169 VDDA.n168 0.3295
R5991 VDDA.n168 VDDA.n167 0.3295
R5992 VDDA.n167 VDDA.n166 0.3295
R5993 VDDA.n172 VDDA.n171 0.3295
R5994 VDDA.n173 VDDA.n172 0.3295
R5995 VDDA.n174 VDDA.n173 0.3295
R5996 VDDA.n179 VDDA.n174 0.3295
R5997 VDDA.n179 VDDA.n178 0.3295
R5998 VDDA.n178 VDDA.n177 0.3295
R5999 VDDA.n177 VDDA.n176 0.3295
R6000 VDDA.n176 VDDA.n175 0.3295
R6001 VDDA.n181 VDDA.n180 0.3295
R6002 VDDA.n182 VDDA.n181 0.3295
R6003 VDDA.n183 VDDA.n182 0.3295
R6004 VDDA.n188 VDDA.n183 0.3295
R6005 VDDA.n188 VDDA.n187 0.3295
R6006 VDDA.n187 VDDA.n186 0.3295
R6007 VDDA.n186 VDDA.n185 0.3295
R6008 VDDA.n185 VDDA.n184 0.3295
R6009 VDDA.n190 VDDA.n189 0.3295
R6010 VDDA.n191 VDDA.n190 0.3295
R6011 VDDA.n192 VDDA.n191 0.3295
R6012 VDDA.n197 VDDA.n192 0.3295
R6013 VDDA.n197 VDDA.n196 0.3295
R6014 VDDA.n196 VDDA.n195 0.3295
R6015 VDDA.n195 VDDA.n194 0.3295
R6016 VDDA.n194 VDDA.n193 0.3295
R6017 VDDA.n199 VDDA.n198 0.3295
R6018 VDDA.n200 VDDA.n199 0.3295
R6019 VDDA.n201 VDDA.n200 0.3295
R6020 VDDA.n206 VDDA.n201 0.3295
R6021 VDDA.n206 VDDA.n205 0.3295
R6022 VDDA.n205 VDDA.n204 0.3295
R6023 VDDA.n204 VDDA.n203 0.3295
R6024 VDDA.n203 VDDA.n202 0.3295
R6025 VDDA.n208 VDDA.n207 0.3295
R6026 VDDA.n209 VDDA.n208 0.3295
R6027 VDDA.n210 VDDA.n209 0.3295
R6028 VDDA.n215 VDDA.n210 0.3295
R6029 VDDA.n215 VDDA.n214 0.3295
R6030 VDDA.n214 VDDA.n213 0.3295
R6031 VDDA.n213 VDDA.n212 0.3295
R6032 VDDA.n212 VDDA.n211 0.3295
R6033 VDDA.n217 VDDA.n216 0.3295
R6034 VDDA.n218 VDDA.n217 0.3295
R6035 VDDA.n219 VDDA.n218 0.3295
R6036 VDDA.n220 VDDA.n219 0.3295
R6037 VDDA.n221 VDDA.n220 0.3295
R6038 VDDA.n222 VDDA.n221 0.3295
R6039 VDDA.n223 VDDA.n222 0.3295
R6040 VDDA.n224 VDDA.n223 0.3295
R6041 VDDA.n225 VDDA.n224 0.3295
R6042 VDDA.n246 VDDA.n225 0.318925
R6043 VDDA.n439 VDDA.n412 0.294805
R6044 VDDA.n386 VDDA.n383 0.292167
R6045 VDDA.n394 VDDA.n391 0.292167
R6046 VDDA.n408 VDDA.n407 0.292167
R6047 VDDA.n624 VDDA.n622 0.2825
R6048 VDDA.n626 VDDA.n624 0.2825
R6049 VDDA.n628 VDDA.n626 0.2825
R6050 VDDA.n629 VDDA.n628 0.2825
R6051 VDDA.n290 VDDA.n288 0.2825
R6052 VDDA.n292 VDDA.n290 0.2825
R6053 VDDA.n294 VDDA.n292 0.2825
R6054 VDDA.n295 VDDA.n294 0.2825
R6055 VDDA.n26 VDDA.n17 0.2825
R6056 VDDA.n35 VDDA.n26 0.2825
R6057 VDDA.n44 VDDA.n35 0.2825
R6058 VDDA.n53 VDDA.n44 0.2825
R6059 VDDA.n62 VDDA.n53 0.2825
R6060 VDDA.n71 VDDA.n62 0.2825
R6061 VDDA.n80 VDDA.n71 0.2825
R6062 VDDA.n89 VDDA.n80 0.2825
R6063 VDDA.n98 VDDA.n89 0.2825
R6064 VDDA.n107 VDDA.n98 0.2825
R6065 VDDA.n116 VDDA.n107 0.2825
R6066 VDDA.n125 VDDA.n116 0.2825
R6067 VDDA.n134 VDDA.n125 0.2825
R6068 VDDA.n143 VDDA.n134 0.2825
R6069 VDDA.n152 VDDA.n143 0.2825
R6070 VDDA.n161 VDDA.n152 0.2825
R6071 VDDA.n170 VDDA.n161 0.2825
R6072 VDDA.n179 VDDA.n170 0.2825
R6073 VDDA.n188 VDDA.n179 0.2825
R6074 VDDA.n197 VDDA.n188 0.2825
R6075 VDDA.n206 VDDA.n197 0.2825
R6076 VDDA.n215 VDDA.n206 0.2825
R6077 VDDA.n220 VDDA.n215 0.2825
R6078 VDDA.n617 VDDA.n606 0.215525
R6079 VDDA.n441 VDDA.n368 0.1755
R6080 VDDA.n448 VDDA.n368 0.1755
R6081 VDDA.n449 VDDA.n448 0.1755
R6082 VDDA.n444 VDDA.n443 0.1755
R6083 VDDA.n447 VDDA.n444 0.1755
R6084 VDDA.n447 VDDA.n367 0.1755
R6085 VDDA.n441 VDDA.n440 0.163
R6086 VDDA.n603 VDDA.n449 0.163
R6087 VDDA.n443 VDDA.n369 0.163
R6088 VDDA.n604 VDDA.n367 0.163
R6089 VDDA.t379 VDDA.t189 0.1603
R6090 VDDA.t302 VDDA.t349 0.1603
R6091 VDDA.t258 VDDA.t296 0.1603
R6092 VDDA.t318 VDDA.t304 0.1603
R6093 VDDA.t240 VDDA.t283 0.1603
R6094 VDDA.n283 VDDA.t298 0.159278
R6095 VDDA.n284 VDDA.t343 0.159278
R6096 VDDA.n285 VDDA.t300 0.159278
R6097 VDDA.n286 VDDA.t377 0.159278
R6098 VDDA.n609 VDDA.n6 0.146333
R6099 VDDA.n614 VDDA.n609 0.146333
R6100 VDDA.n610 VDDA.n7 0.146333
R6101 VDDA.n613 VDDA.n610 0.146333
R6102 VDDA.n613 VDDA.n608 0.146333
R6103 VDDA.n355 VDDA.n326 0.146333
R6104 VDDA.n362 VDDA.n326 0.146333
R6105 VDDA.n358 VDDA.n357 0.146333
R6106 VDDA.n361 VDDA.n358 0.146333
R6107 VDDA.n361 VDDA.n325 0.146333
R6108 VDDA.n313 VDDA.n280 0.146333
R6109 VDDA.n320 VDDA.n280 0.146333
R6110 VDDA.n316 VDDA.n315 0.146333
R6111 VDDA.n319 VDDA.n316 0.146333
R6112 VDDA.n319 VDDA.n279 0.146333
R6113 VDDA.n236 VDDA.n231 0.146333
R6114 VDDA.n243 VDDA.n231 0.146333
R6115 VDDA.n239 VDDA.n238 0.146333
R6116 VDDA.n242 VDDA.n239 0.146333
R6117 VDDA.n242 VDDA.n230 0.146333
R6118 VDDA.n606 VDDA.n365 0.145025
R6119 VDDA.n286 VDDA.t281 0.1368
R6120 VDDA.n286 VDDA.t379 0.1368
R6121 VDDA.n285 VDDA.t216 0.1368
R6122 VDDA.n285 VDDA.t302 0.1368
R6123 VDDA.n284 VDDA.t375 0.1368
R6124 VDDA.n284 VDDA.t258 0.1368
R6125 VDDA.n283 VDDA.t214 0.1368
R6126 VDDA.n283 VDDA.t318 0.1368
R6127 VDDA.n282 VDDA.t365 0.1368
R6128 VDDA.n282 VDDA.t240 0.1368
R6129 VDDA.n620 VDDA.n6 0.135917
R6130 VDDA.n619 VDDA.n7 0.135917
R6131 VDDA.n355 VDDA.n354 0.135917
R6132 VDDA.n357 VDDA.n327 0.135917
R6133 VDDA.n313 VDDA.n312 0.135917
R6134 VDDA.n315 VDDA.n281 0.135917
R6135 VDDA.n236 VDDA.n235 0.135917
R6136 VDDA.n238 VDDA.n232 0.135917
R6137 VDDA.n383 VDDA.n378 0.1255
R6138 VDDA.n386 VDDA.n385 0.115083
R6139 VDDA.n385 VDDA.n376 0.115083
R6140 VDDA.n391 VDDA.n376 0.115083
R6141 VDDA.n393 VDDA.n372 0.115083
R6142 VDDA.n411 VDDA.n372 0.115083
R6143 VDDA.n411 VDDA.n410 0.115083
R6144 VDDA.n410 VDDA.n409 0.115083
R6145 VDDA.n407 VDDA.n406 0.115083
R6146 VDDA.n406 VDDA.n405 0.115083
R6147 VDDA.n365 VDDA.n323 0.100963
R6148 VDDA.n259 VDDA 0.0806938
R6149 VDDA.n394 VDDA.n393 0.0682083
R6150 VDDA.n409 VDDA.n408 0.0682083
R6151 VDDA.n615 VDDA.n608 0.0667303
R6152 VDDA.n363 VDDA.n325 0.0667303
R6153 VDDA.n321 VDDA.n279 0.0667303
R6154 VDDA.n244 VDDA.n230 0.0667303
R6155 VDDA.n446 VDDA.n445 0.0663
R6156 VDDA.n442 VDDA.n249 0.0616
R6157 VDDA.n605 VDDA.n366 0.0616
R6158 VDDA.n612 VDDA.n611 0.0553333
R6159 VDDA.n360 VDDA.n359 0.0553333
R6160 VDDA.n318 VDDA.n317 0.0553333
R6161 VDDA.n241 VDDA.n240 0.0553333
R6162 VDDA.n618 VDDA.n8 0.0514167
R6163 VDDA.n616 VDDA.n607 0.0514167
R6164 VDDA.n356 VDDA.n252 0.0514167
R6165 VDDA.n364 VDDA.n324 0.0514167
R6166 VDDA.n314 VDDA.n255 0.0514167
R6167 VDDA.n322 VDDA.n278 0.0514167
R6168 VDDA.n237 VDDA.n226 0.0514167
R6169 VDDA.n245 VDDA.n229 0.0514167
R6170 VDDA.n617 VDDA.n246 0.034575
R6171 VDDA.n445 VDDA.n250 0.0335856
R6172 VDDA.n366 VDDA.n251 0.0335856
R6173 VDDA.n446 VDDA.n251 0.0335856
R6174 VDDA.n442 VDDA.n250 0.0335856
R6175 VDDA.n611 VDDA.n247 0.028198
R6176 VDDA.n607 VDDA.n248 0.028198
R6177 VDDA.n359 VDDA.n253 0.028198
R6178 VDDA.n324 VDDA.n254 0.028198
R6179 VDDA.n317 VDDA.n256 0.028198
R6180 VDDA.n278 VDDA.n257 0.028198
R6181 VDDA.n240 VDDA.n227 0.028198
R6182 VDDA.n229 VDDA.n228 0.028198
R6183 VDDA.n241 VDDA.n228 0.028198
R6184 VDDA.n237 VDDA.n227 0.028198
R6185 VDDA.n318 VDDA.n257 0.028198
R6186 VDDA.n314 VDDA.n256 0.028198
R6187 VDDA.n360 VDDA.n254 0.028198
R6188 VDDA.n356 VDDA.n253 0.028198
R6189 VDDA.n612 VDDA.n248 0.028198
R6190 VDDA.n247 VDDA.n8 0.028198
R6191 VDDA.n277 VDDA.n260 0.0116625
R6192 VDDA.n275 VDDA.n260 0.0116625
R6193 VDDA.n274 VDDA.n264 0.0068649
R6194 VDDA.n271 VDDA.n264 0.0068649
R6195 VDDA.n272 VDDA.n265 0.0068649
R6196 VDDA.n273 VDDA.n271 0.0068649
R6197 VDDA.n273 VDDA.n272 0.0068649
R6198 VDDA.n275 VDDA.n274 0.0068649
R6199 VDDA.n266 VDDA.n265 0.00657213
R6200 VDDA.n270 VDDA.n269 0.00657213
R6201 VDDA.n267 VDDA.n266 0.00657213
R6202 VDDA.n270 VDDA.n267 0.00657213
R6203 VDDA.n268 VDDA.n258 0.00393497
R6204 VDDA.n268 VDDA.n262 0.00393497
R6205 VDDA.n262 VDDA.n261 0.0036417
R6206 VDDA.n276 VDDA.n263 0.0036417
R6207 VDDA.n261 VDDA.n259 0.0036417
R6208 VDDA.n263 VDDA.n258 0.0036417
R6209 VDDA.t298 VDDA.n282 0.00152174
R6210 VDDA.t343 VDDA.n283 0.00152174
R6211 VDDA.t300 VDDA.n284 0.00152174
R6212 VDDA.t377 VDDA.n285 0.00152174
R6213 VDDA.t218 VDDA.n286 0.00152174
R6214 VOUT+.n9 VOUT+.t0 113.192
R6215 VOUT+.n11 VOUT+.n10 34.9935
R6216 VOUT+.n13 VOUT+.n12 34.9935
R6217 VOUT+.n17 VOUT+.n16 34.9935
R6218 VOUT+.n20 VOUT+.n19 34.9935
R6219 VOUT+.n23 VOUT+.n22 34.9935
R6220 VOUT+.n27 VOUT+.n26 34.9935
R6221 VOUT+.n110 VOUT+.n30 20.5005
R6222 VOUT+.n110 VOUT+.n109 11.6871
R6223 VOUT+.n2 VOUT+.n1 9.73997
R6224 VOUT+.n4 VOUT+.n3 9.73997
R6225 VOUT+.n7 VOUT+.n6 9.73997
R6226 VOUT+ VOUT+.n110 9.34425
R6227 VOUT+.n7 VOUT+.n5 7.14633
R6228 VOUT+.n5 VOUT+.n2 7.14633
R6229 VOUT+.n2 VOUT+.n0 7.14633
R6230 VOUT+.n10 VOUT+.t9 6.56717
R6231 VOUT+.n10 VOUT+.t14 6.56717
R6232 VOUT+.n12 VOUT+.t17 6.56717
R6233 VOUT+.n12 VOUT+.t15 6.56717
R6234 VOUT+.n16 VOUT+.t8 6.56717
R6235 VOUT+.n16 VOUT+.t18 6.56717
R6236 VOUT+.n19 VOUT+.t10 6.56717
R6237 VOUT+.n19 VOUT+.t13 6.56717
R6238 VOUT+.n22 VOUT+.t11 6.56717
R6239 VOUT+.n22 VOUT+.t16 6.56717
R6240 VOUT+.n26 VOUT+.t12 6.56717
R6241 VOUT+.n26 VOUT+.t7 6.56717
R6242 VOUT+.n21 VOUT+.n17 6.3755
R6243 VOUT+.n18 VOUT+.n17 6.3755
R6244 VOUT+.n29 VOUT+.n13 6.3755
R6245 VOUT+.n15 VOUT+.n13 6.3755
R6246 VOUT+.n4 VOUT+.n0 6.02133
R6247 VOUT+.n5 VOUT+.n4 6.02133
R6248 VOUT+.n8 VOUT+.n7 6.02133
R6249 VOUT+.n20 VOUT+.n18 5.813
R6250 VOUT+.n21 VOUT+.n20 5.813
R6251 VOUT+.n23 VOUT+.n14 5.813
R6252 VOUT+.n24 VOUT+.n23 5.813
R6253 VOUT+.n28 VOUT+.n27 5.813
R6254 VOUT+.n27 VOUT+.n25 5.813
R6255 VOUT+.n15 VOUT+.n11 5.813
R6256 VOUT+.n57 VOUT+.t66 4.8295
R6257 VOUT+.n59 VOUT+.t137 4.8295
R6258 VOUT+.n61 VOUT+.t27 4.8295
R6259 VOUT+.n63 VOUT+.t81 4.8295
R6260 VOUT+.n65 VOUT+.t114 4.8295
R6261 VOUT+.n77 VOUT+.t105 4.8295
R6262 VOUT+.n79 VOUT+.t48 4.8295
R6263 VOUT+.n80 VOUT+.t62 4.8295
R6264 VOUT+.n82 VOUT+.t139 4.8295
R6265 VOUT+.n83 VOUT+.t26 4.8295
R6266 VOUT+.n85 VOUT+.t104 4.8295
R6267 VOUT+.n86 VOUT+.t129 4.8295
R6268 VOUT+.n88 VOUT+.t135 4.8295
R6269 VOUT+.n89 VOUT+.t23 4.8295
R6270 VOUT+.n91 VOUT+.t97 4.8295
R6271 VOUT+.n92 VOUT+.t123 4.8295
R6272 VOUT+.n94 VOUT+.t57 4.8295
R6273 VOUT+.n95 VOUT+.t85 4.8295
R6274 VOUT+.n97 VOUT+.t89 4.8295
R6275 VOUT+.n98 VOUT+.t118 4.8295
R6276 VOUT+.n100 VOUT+.t52 4.8295
R6277 VOUT+.n101 VOUT+.t80 4.8295
R6278 VOUT+.n103 VOUT+.t151 4.8295
R6279 VOUT+.n104 VOUT+.t41 4.8295
R6280 VOUT+.n31 VOUT+.t35 4.8295
R6281 VOUT+.n43 VOUT+.t58 4.8295
R6282 VOUT+.n45 VOUT+.t103 4.8295
R6283 VOUT+.n46 VOUT+.t130 4.8295
R6284 VOUT+.n48 VOUT+.t67 4.8295
R6285 VOUT+.n49 VOUT+.t98 4.8295
R6286 VOUT+.n51 VOUT+.t109 4.8295
R6287 VOUT+.n52 VOUT+.t136 4.8295
R6288 VOUT+.n54 VOUT+.t145 4.8295
R6289 VOUT+.n55 VOUT+.t32 4.8295
R6290 VOUT+.n106 VOUT+.t74 4.8295
R6291 VOUT+.n70 VOUT+.t37 4.8154
R6292 VOUT+.n69 VOUT+.t76 4.8154
R6293 VOUT+.n68 VOUT+.t56 4.8154
R6294 VOUT+.n67 VOUT+.t91 4.8154
R6295 VOUT+.n76 VOUT+.t75 4.806
R6296 VOUT+.n75 VOUT+.t53 4.806
R6297 VOUT+.n74 VOUT+.t90 4.806
R6298 VOUT+.n73 VOUT+.t126 4.806
R6299 VOUT+.n72 VOUT+.t110 4.806
R6300 VOUT+.n71 VOUT+.t148 4.806
R6301 VOUT+.n70 VOUT+.t44 4.806
R6302 VOUT+.n69 VOUT+.t82 4.806
R6303 VOUT+.n68 VOUT+.t61 4.806
R6304 VOUT+.n67 VOUT+.t100 4.806
R6305 VOUT+.n42 VOUT+.t99 4.806
R6306 VOUT+.n41 VOUT+.t149 4.806
R6307 VOUT+.n40 VOUT+.t43 4.806
R6308 VOUT+.n39 VOUT+.t77 4.806
R6309 VOUT+.n38 VOUT+.t125 4.806
R6310 VOUT+.n37 VOUT+.t20 4.806
R6311 VOUT+.n36 VOUT+.t59 4.806
R6312 VOUT+.n35 VOUT+.t92 4.806
R6313 VOUT+.n34 VOUT+.t143 4.806
R6314 VOUT+.n33 VOUT+.t39 4.806
R6315 VOUT+.n58 VOUT+.t36 4.5005
R6316 VOUT+.n57 VOUT+.t28 4.5005
R6317 VOUT+.n59 VOUT+.t33 4.5005
R6318 VOUT+.n60 VOUT+.t86 4.5005
R6319 VOUT+.n61 VOUT+.t69 4.5005
R6320 VOUT+.n62 VOUT+.t122 4.5005
R6321 VOUT+.n63 VOUT+.t119 4.5005
R6322 VOUT+.n64 VOUT+.t106 4.5005
R6323 VOUT+.n65 VOUT+.t156 4.5005
R6324 VOUT+.n66 VOUT+.t140 4.5005
R6325 VOUT+.n67 VOUT+.t131 4.5005
R6326 VOUT+.n68 VOUT+.t94 4.5005
R6327 VOUT+.n69 VOUT+.t115 4.5005
R6328 VOUT+.n70 VOUT+.t78 4.5005
R6329 VOUT+.n71 VOUT+.t42 4.5005
R6330 VOUT+.n72 VOUT+.t141 4.5005
R6331 VOUT+.n73 VOUT+.t22 4.5005
R6332 VOUT+.n74 VOUT+.t124 4.5005
R6333 VOUT+.n75 VOUT+.t87 4.5005
R6334 VOUT+.n76 VOUT+.t112 4.5005
R6335 VOUT+.n78 VOUT+.t71 4.5005
R6336 VOUT+.n77 VOUT+.t68 4.5005
R6337 VOUT+.n79 VOUT+.t70 4.5005
R6338 VOUT+.n81 VOUT+.t29 4.5005
R6339 VOUT+.n80 VOUT+.t24 4.5005
R6340 VOUT+.n82 VOUT+.t88 4.5005
R6341 VOUT+.n84 VOUT+.t54 4.5005
R6342 VOUT+.n83 VOUT+.t25 4.5005
R6343 VOUT+.n85 VOUT+.t51 4.5005
R6344 VOUT+.n87 VOUT+.t154 4.5005
R6345 VOUT+.n86 VOUT+.t128 4.5005
R6346 VOUT+.n88 VOUT+.t83 4.5005
R6347 VOUT+.n90 VOUT+.t50 4.5005
R6348 VOUT+.n89 VOUT+.t21 4.5005
R6349 VOUT+.n91 VOUT+.t46 4.5005
R6350 VOUT+.n93 VOUT+.t150 4.5005
R6351 VOUT+.n92 VOUT+.t121 4.5005
R6352 VOUT+.n94 VOUT+.t144 4.5005
R6353 VOUT+.n96 VOUT+.t111 4.5005
R6354 VOUT+.n95 VOUT+.t84 4.5005
R6355 VOUT+.n97 VOUT+.t38 4.5005
R6356 VOUT+.n99 VOUT+.t142 4.5005
R6357 VOUT+.n98 VOUT+.t117 4.5005
R6358 VOUT+.n100 VOUT+.t138 4.5005
R6359 VOUT+.n102 VOUT+.t108 4.5005
R6360 VOUT+.n101 VOUT+.t79 4.5005
R6361 VOUT+.n103 VOUT+.t102 4.5005
R6362 VOUT+.n105 VOUT+.t64 4.5005
R6363 VOUT+.n104 VOUT+.t40 4.5005
R6364 VOUT+.n32 VOUT+.t63 4.5005
R6365 VOUT+.n31 VOUT+.t34 4.5005
R6366 VOUT+.n33 VOUT+.t95 4.5005
R6367 VOUT+.n34 VOUT+.t146 4.5005
R6368 VOUT+.n35 VOUT+.t107 4.5005
R6369 VOUT+.n36 VOUT+.t153 4.5005
R6370 VOUT+.n37 VOUT+.t65 4.5005
R6371 VOUT+.n38 VOUT+.t113 4.5005
R6372 VOUT+.n39 VOUT+.t72 4.5005
R6373 VOUT+.n40 VOUT+.t120 4.5005
R6374 VOUT+.n41 VOUT+.t31 4.5005
R6375 VOUT+.n42 VOUT+.t132 4.5005
R6376 VOUT+.n44 VOUT+.t45 4.5005
R6377 VOUT+.n43 VOUT+.t147 4.5005
R6378 VOUT+.n45 VOUT+.t49 4.5005
R6379 VOUT+.n47 VOUT+.t152 4.5005
R6380 VOUT+.n46 VOUT+.t127 4.5005
R6381 VOUT+.n48 VOUT+.t155 4.5005
R6382 VOUT+.n50 VOUT+.t116 4.5005
R6383 VOUT+.n49 VOUT+.t96 4.5005
R6384 VOUT+.n51 VOUT+.t55 4.5005
R6385 VOUT+.n53 VOUT+.t19 4.5005
R6386 VOUT+.n52 VOUT+.t134 4.5005
R6387 VOUT+.n54 VOUT+.t93 4.5005
R6388 VOUT+.n56 VOUT+.t60 4.5005
R6389 VOUT+.n55 VOUT+.t30 4.5005
R6390 VOUT+.n109 VOUT+.t47 4.5005
R6391 VOUT+.n108 VOUT+.t133 4.5005
R6392 VOUT+.n107 VOUT+.t101 4.5005
R6393 VOUT+.n106 VOUT+.t73 4.5005
R6394 VOUT+.n30 VOUT+.n29 4.5005
R6395 VOUT+.n1 VOUT+.t6 3.42907
R6396 VOUT+.n1 VOUT+.t3 3.42907
R6397 VOUT+.n3 VOUT+.t2 3.42907
R6398 VOUT+.n3 VOUT+.t1 3.42907
R6399 VOUT+.n6 VOUT+.t4 3.42907
R6400 VOUT+.n6 VOUT+.t5 3.42907
R6401 VOUT+ VOUT+.n9 1.938
R6402 VOUT+.n9 VOUT+.n8 1.84425
R6403 VOUT+.n30 VOUT+.n11 1.313
R6404 VOUT+.n8 VOUT+.n0 1.1255
R6405 VOUT+.n25 VOUT+.n15 0.563
R6406 VOUT+.n25 VOUT+.n24 0.563
R6407 VOUT+.n24 VOUT+.n21 0.563
R6408 VOUT+.n18 VOUT+.n14 0.563
R6409 VOUT+.n28 VOUT+.n14 0.563
R6410 VOUT+.n29 VOUT+.n28 0.563
R6411 VOUT+.n58 VOUT+.n57 0.3295
R6412 VOUT+.n60 VOUT+.n59 0.3295
R6413 VOUT+.n62 VOUT+.n61 0.3295
R6414 VOUT+.n64 VOUT+.n63 0.3295
R6415 VOUT+.n66 VOUT+.n65 0.3295
R6416 VOUT+.n68 VOUT+.n67 0.3295
R6417 VOUT+.n69 VOUT+.n68 0.3295
R6418 VOUT+.n70 VOUT+.n69 0.3295
R6419 VOUT+.n71 VOUT+.n70 0.3295
R6420 VOUT+.n72 VOUT+.n71 0.3295
R6421 VOUT+.n73 VOUT+.n72 0.3295
R6422 VOUT+.n74 VOUT+.n73 0.3295
R6423 VOUT+.n75 VOUT+.n74 0.3295
R6424 VOUT+.n76 VOUT+.n75 0.3295
R6425 VOUT+.n78 VOUT+.n76 0.3295
R6426 VOUT+.n78 VOUT+.n77 0.3295
R6427 VOUT+.n81 VOUT+.n79 0.3295
R6428 VOUT+.n81 VOUT+.n80 0.3295
R6429 VOUT+.n84 VOUT+.n82 0.3295
R6430 VOUT+.n84 VOUT+.n83 0.3295
R6431 VOUT+.n87 VOUT+.n85 0.3295
R6432 VOUT+.n87 VOUT+.n86 0.3295
R6433 VOUT+.n90 VOUT+.n88 0.3295
R6434 VOUT+.n90 VOUT+.n89 0.3295
R6435 VOUT+.n93 VOUT+.n91 0.3295
R6436 VOUT+.n93 VOUT+.n92 0.3295
R6437 VOUT+.n96 VOUT+.n94 0.3295
R6438 VOUT+.n96 VOUT+.n95 0.3295
R6439 VOUT+.n99 VOUT+.n97 0.3295
R6440 VOUT+.n99 VOUT+.n98 0.3295
R6441 VOUT+.n102 VOUT+.n100 0.3295
R6442 VOUT+.n102 VOUT+.n101 0.3295
R6443 VOUT+.n105 VOUT+.n103 0.3295
R6444 VOUT+.n105 VOUT+.n104 0.3295
R6445 VOUT+.n32 VOUT+.n31 0.3295
R6446 VOUT+.n34 VOUT+.n33 0.3295
R6447 VOUT+.n35 VOUT+.n34 0.3295
R6448 VOUT+.n36 VOUT+.n35 0.3295
R6449 VOUT+.n37 VOUT+.n36 0.3295
R6450 VOUT+.n38 VOUT+.n37 0.3295
R6451 VOUT+.n39 VOUT+.n38 0.3295
R6452 VOUT+.n40 VOUT+.n39 0.3295
R6453 VOUT+.n41 VOUT+.n40 0.3295
R6454 VOUT+.n42 VOUT+.n41 0.3295
R6455 VOUT+.n44 VOUT+.n42 0.3295
R6456 VOUT+.n44 VOUT+.n43 0.3295
R6457 VOUT+.n47 VOUT+.n45 0.3295
R6458 VOUT+.n47 VOUT+.n46 0.3295
R6459 VOUT+.n50 VOUT+.n48 0.3295
R6460 VOUT+.n50 VOUT+.n49 0.3295
R6461 VOUT+.n53 VOUT+.n51 0.3295
R6462 VOUT+.n53 VOUT+.n52 0.3295
R6463 VOUT+.n56 VOUT+.n54 0.3295
R6464 VOUT+.n56 VOUT+.n55 0.3295
R6465 VOUT+.n109 VOUT+.n108 0.3295
R6466 VOUT+.n108 VOUT+.n107 0.3295
R6467 VOUT+.n107 VOUT+.n106 0.3295
R6468 VOUT+.n74 VOUT+.n60 0.306
R6469 VOUT+.n73 VOUT+.n62 0.306
R6470 VOUT+.n72 VOUT+.n64 0.306
R6471 VOUT+.n71 VOUT+.n66 0.306
R6472 VOUT+.n78 VOUT+.n58 0.2825
R6473 VOUT+.n81 VOUT+.n78 0.2825
R6474 VOUT+.n84 VOUT+.n81 0.2825
R6475 VOUT+.n87 VOUT+.n84 0.2825
R6476 VOUT+.n90 VOUT+.n87 0.2825
R6477 VOUT+.n93 VOUT+.n90 0.2825
R6478 VOUT+.n96 VOUT+.n93 0.2825
R6479 VOUT+.n99 VOUT+.n96 0.2825
R6480 VOUT+.n102 VOUT+.n99 0.2825
R6481 VOUT+.n105 VOUT+.n102 0.2825
R6482 VOUT+.n44 VOUT+.n32 0.2825
R6483 VOUT+.n47 VOUT+.n44 0.2825
R6484 VOUT+.n50 VOUT+.n47 0.2825
R6485 VOUT+.n53 VOUT+.n50 0.2825
R6486 VOUT+.n56 VOUT+.n53 0.2825
R6487 VOUT+.n107 VOUT+.n56 0.2825
R6488 VOUT+.n107 VOUT+.n105 0.2825
R6489 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t19 369.534
R6490 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t21 369.534
R6491 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t5 369.534
R6492 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.t20 369.534
R6493 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t13 369.534
R6494 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.t11 369.534
R6495 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.t0 369.534
R6496 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n0 360.678
R6497 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t7 249.034
R6498 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t18 192.8
R6499 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t6 192.8
R6500 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t12 192.8
R6501 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t9 192.8
R6502 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t15 192.8
R6503 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.t8 192.8
R6504 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t10 192.8
R6505 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.t17 192.8
R6506 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t16 192.8
R6507 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t22 192.8
R6508 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.t14 192.8
R6509 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R6510 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.n2 176.733
R6511 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n10 176.733
R6512 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.n11 176.733
R6513 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n5 167.843
R6514 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 166.343
R6515 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n14 166.343
R6516 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n17 166.343
R6517 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n18 141.752
R6518 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 56.2338
R6519 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n1 56.2338
R6520 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R6521 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.n6 56.2338
R6522 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n13 56.2338
R6523 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n12 56.2338
R6524 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n16 56.2338
R6525 bgr_11_0.NFET_GATE_10uA.t4 bgr_11_0.NFET_GATE_10uA.n19 39.4005
R6526 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t3 39.4005
R6527 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t2 24.0005
R6528 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t1 24.0005
R6529 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n15 2.01612
R6530 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n9 1.5005
R6531 bgr_11_0.cap_res2.t20 bgr_11_0.cap_res2.t18 121.245
R6532 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.t8 0.1603
R6533 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.t2 0.1603
R6534 bgr_11_0.cap_res2.t1 bgr_11_0.cap_res2.t15 0.1603
R6535 bgr_11_0.cap_res2.t5 bgr_11_0.cap_res2.t0 0.1603
R6536 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.t14 0.1603
R6537 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t4 0.159278
R6538 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t10 0.159278
R6539 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t6 0.159278
R6540 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t12 0.159278
R6541 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t3 0.1368
R6542 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t13 0.1368
R6543 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t17 0.1368
R6544 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t7 0.1368
R6545 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t11 0.1368
R6546 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t1 0.1368
R6547 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t16 0.1368
R6548 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t5 0.1368
R6549 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t9 0.1368
R6550 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t19 0.1368
R6551 bgr_11_0.cap_res2.t4 bgr_11_0.cap_res2.n0 0.00152174
R6552 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.n1 0.00152174
R6553 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.n2 0.00152174
R6554 bgr_11_0.cap_res2.t12 bgr_11_0.cap_res2.n3 0.00152174
R6555 bgr_11_0.cap_res2.t18 bgr_11_0.cap_res2.n4 0.00152174
R6556 VOUT-.n110 VOUT-.t5 113.16
R6557 VOUT-.n1 VOUT-.n0 34.9935
R6558 VOUT-.n5 VOUT-.n4 34.9935
R6559 VOUT-.n7 VOUT-.n6 34.9935
R6560 VOUT-.n11 VOUT-.n10 34.9935
R6561 VOUT-.n14 VOUT-.n13 34.9935
R6562 VOUT-.n18 VOUT-.n17 34.9935
R6563 VOUT-.n100 VOUT-.n20 20.4693
R6564 VOUT-.n100 VOUT-.n99 11.6871
R6565 VOUT-.n103 VOUT-.n102 9.73997
R6566 VOUT-.n105 VOUT-.n104 9.73997
R6567 VOUT-.n108 VOUT-.n107 9.73997
R6568 VOUT- VOUT-.n100 9.6255
R6569 VOUT-.n108 VOUT-.n106 7.14633
R6570 VOUT-.n106 VOUT-.n103 7.14633
R6571 VOUT-.n103 VOUT-.n101 7.14633
R6572 VOUT-.n0 VOUT-.t2 6.56717
R6573 VOUT-.n0 VOUT-.t15 6.56717
R6574 VOUT-.n4 VOUT-.t13 6.56717
R6575 VOUT-.n4 VOUT-.t17 6.56717
R6576 VOUT-.n6 VOUT-.t7 6.56717
R6577 VOUT-.n6 VOUT-.t8 6.56717
R6578 VOUT-.n10 VOUT-.t1 6.56717
R6579 VOUT-.n10 VOUT-.t18 6.56717
R6580 VOUT-.n13 VOUT-.t3 6.56717
R6581 VOUT-.n13 VOUT-.t16 6.56717
R6582 VOUT-.n17 VOUT-.t10 6.56717
R6583 VOUT-.n17 VOUT-.t14 6.56717
R6584 VOUT-.n18 VOUT-.n16 6.3755
R6585 VOUT-.n19 VOUT-.n18 6.3755
R6586 VOUT-.n8 VOUT-.n5 6.3755
R6587 VOUT-.n5 VOUT-.n3 6.3755
R6588 VOUT-.n105 VOUT-.n101 6.02133
R6589 VOUT-.n106 VOUT-.n105 6.02133
R6590 VOUT-.n109 VOUT-.n108 6.02133
R6591 VOUT-.n7 VOUT-.n3 5.813
R6592 VOUT-.n8 VOUT-.n7 5.813
R6593 VOUT-.n12 VOUT-.n11 5.813
R6594 VOUT-.n11 VOUT-.n9 5.813
R6595 VOUT-.n15 VOUT-.n14 5.813
R6596 VOUT-.n14 VOUT-.n2 5.813
R6597 VOUT-.n16 VOUT-.n1 5.813
R6598 VOUT-.n47 VOUT-.t56 4.8295
R6599 VOUT-.n56 VOUT-.t88 4.8295
R6600 VOUT-.n54 VOUT-.t117 4.8295
R6601 VOUT-.n52 VOUT-.t156 4.8295
R6602 VOUT-.n50 VOUT-.t57 4.8295
R6603 VOUT-.n49 VOUT-.t87 4.8295
R6604 VOUT-.n69 VOUT-.t50 4.8295
R6605 VOUT-.n70 VOUT-.t95 4.8295
R6606 VOUT-.n72 VOUT-.t19 4.8295
R6607 VOUT-.n73 VOUT-.t144 4.8295
R6608 VOUT-.n75 VOUT-.t114 4.8295
R6609 VOUT-.n76 VOUT-.t100 4.8295
R6610 VOUT-.n78 VOUT-.t154 4.8295
R6611 VOUT-.n79 VOUT-.t138 4.8295
R6612 VOUT-.n81 VOUT-.t108 4.8295
R6613 VOUT-.n82 VOUT-.t96 4.8295
R6614 VOUT-.n84 VOUT-.t72 4.8295
R6615 VOUT-.n85 VOUT-.t60 4.8295
R6616 VOUT-.n87 VOUT-.t105 4.8295
R6617 VOUT-.n88 VOUT-.t93 4.8295
R6618 VOUT-.n90 VOUT-.t68 4.8295
R6619 VOUT-.n91 VOUT-.t58 4.8295
R6620 VOUT-.n93 VOUT-.t28 4.8295
R6621 VOUT-.n94 VOUT-.t152 4.8295
R6622 VOUT-.n21 VOUT-.t24 4.8295
R6623 VOUT-.n23 VOUT-.t61 4.8295
R6624 VOUT-.n35 VOUT-.t113 4.8295
R6625 VOUT-.n36 VOUT-.t102 4.8295
R6626 VOUT-.n38 VOUT-.t85 4.8295
R6627 VOUT-.n39 VOUT-.t66 4.8295
R6628 VOUT-.n41 VOUT-.t120 4.8295
R6629 VOUT-.n42 VOUT-.t103 4.8295
R6630 VOUT-.n44 VOUT-.t22 4.8295
R6631 VOUT-.n45 VOUT-.t147 4.8295
R6632 VOUT-.n96 VOUT-.t62 4.8295
R6633 VOUT-.n58 VOUT-.t128 4.8154
R6634 VOUT-.n59 VOUT-.t104 4.8154
R6635 VOUT-.n60 VOUT-.t122 4.8154
R6636 VOUT-.n61 VOUT-.t23 4.8154
R6637 VOUT-.n58 VOUT-.t136 4.806
R6638 VOUT-.n59 VOUT-.t107 4.806
R6639 VOUT-.n60 VOUT-.t130 4.806
R6640 VOUT-.n61 VOUT-.t30 4.806
R6641 VOUT-.n62 VOUT-.t146 4.806
R6642 VOUT-.n63 VOUT-.t49 4.806
R6643 VOUT-.n64 VOUT-.t82 4.806
R6644 VOUT-.n65 VOUT-.t116 4.806
R6645 VOUT-.n66 VOUT-.t99 4.806
R6646 VOUT-.n67 VOUT-.t137 4.806
R6647 VOUT-.n24 VOUT-.t73 4.806
R6648 VOUT-.n25 VOUT-.t121 4.806
R6649 VOUT-.n26 VOUT-.t52 4.806
R6650 VOUT-.n27 VOUT-.t81 4.806
R6651 VOUT-.n28 VOUT-.t134 4.806
R6652 VOUT-.n29 VOUT-.t29 4.806
R6653 VOUT-.n30 VOUT-.t63 4.806
R6654 VOUT-.n31 VOUT-.t98 4.806
R6655 VOUT-.n32 VOUT-.t151 4.806
R6656 VOUT-.n33 VOUT-.t48 4.806
R6657 VOUT-.n47 VOUT-.t153 4.5005
R6658 VOUT-.n48 VOUT-.t39 4.5005
R6659 VOUT-.n56 VOUT-.t123 4.5005
R6660 VOUT-.n57 VOUT-.t143 4.5005
R6661 VOUT-.n54 VOUT-.t20 4.5005
R6662 VOUT-.n55 VOUT-.t44 4.5005
R6663 VOUT-.n52 VOUT-.t59 4.5005
R6664 VOUT-.n53 VOUT-.t75 4.5005
R6665 VOUT-.n50 VOUT-.t92 4.5005
R6666 VOUT-.n51 VOUT-.t109 4.5005
R6667 VOUT-.n49 VOUT-.t54 4.5005
R6668 VOUT-.n68 VOUT-.t69 4.5005
R6669 VOUT-.n67 VOUT-.t34 4.5005
R6670 VOUT-.n66 VOUT-.t135 4.5005
R6671 VOUT-.n65 VOUT-.t155 4.5005
R6672 VOUT-.n64 VOUT-.t111 4.5005
R6673 VOUT-.n63 VOUT-.t78 4.5005
R6674 VOUT-.n62 VOUT-.t45 4.5005
R6675 VOUT-.n61 VOUT-.t64 4.5005
R6676 VOUT-.n60 VOUT-.t25 4.5005
R6677 VOUT-.n59 VOUT-.t149 4.5005
R6678 VOUT-.n58 VOUT-.t33 4.5005
R6679 VOUT-.n69 VOUT-.t148 4.5005
R6680 VOUT-.n71 VOUT-.t32 4.5005
R6681 VOUT-.n70 VOUT-.t131 4.5005
R6682 VOUT-.n72 VOUT-.t119 4.5005
R6683 VOUT-.n74 VOUT-.t70 4.5005
R6684 VOUT-.n73 VOUT-.t40 4.5005
R6685 VOUT-.n75 VOUT-.t84 4.5005
R6686 VOUT-.n77 VOUT-.t37 4.5005
R6687 VOUT-.n76 VOUT-.t140 4.5005
R6688 VOUT-.n78 VOUT-.t112 4.5005
R6689 VOUT-.n80 VOUT-.t65 4.5005
R6690 VOUT-.n79 VOUT-.t35 4.5005
R6691 VOUT-.n81 VOUT-.t76 4.5005
R6692 VOUT-.n83 VOUT-.t26 4.5005
R6693 VOUT-.n82 VOUT-.t132 4.5005
R6694 VOUT-.n84 VOUT-.t43 4.5005
R6695 VOUT-.n86 VOUT-.t125 4.5005
R6696 VOUT-.n85 VOUT-.t94 4.5005
R6697 VOUT-.n87 VOUT-.t71 4.5005
R6698 VOUT-.n89 VOUT-.t21 4.5005
R6699 VOUT-.n88 VOUT-.t124 4.5005
R6700 VOUT-.n90 VOUT-.t38 4.5005
R6701 VOUT-.n92 VOUT-.t118 4.5005
R6702 VOUT-.n91 VOUT-.t89 4.5005
R6703 VOUT-.n93 VOUT-.t133 4.5005
R6704 VOUT-.n95 VOUT-.t80 4.5005
R6705 VOUT-.n94 VOUT-.t53 4.5005
R6706 VOUT-.n21 VOUT-.t129 4.5005
R6707 VOUT-.n22 VOUT-.t77 4.5005
R6708 VOUT-.n23 VOUT-.t106 4.5005
R6709 VOUT-.n34 VOUT-.t67 4.5005
R6710 VOUT-.n33 VOUT-.t115 4.5005
R6711 VOUT-.n32 VOUT-.t31 4.5005
R6712 VOUT-.n31 VOUT-.t126 4.5005
R6713 VOUT-.n30 VOUT-.t42 4.5005
R6714 VOUT-.n29 VOUT-.t91 4.5005
R6715 VOUT-.n28 VOUT-.t142 4.5005
R6716 VOUT-.n27 VOUT-.t97 4.5005
R6717 VOUT-.n26 VOUT-.t150 4.5005
R6718 VOUT-.n25 VOUT-.t86 4.5005
R6719 VOUT-.n24 VOUT-.t47 4.5005
R6720 VOUT-.n35 VOUT-.t83 4.5005
R6721 VOUT-.n37 VOUT-.t36 4.5005
R6722 VOUT-.n36 VOUT-.t139 4.5005
R6723 VOUT-.n38 VOUT-.t55 4.5005
R6724 VOUT-.n40 VOUT-.t141 4.5005
R6725 VOUT-.n39 VOUT-.t101 4.5005
R6726 VOUT-.n41 VOUT-.t90 4.5005
R6727 VOUT-.n43 VOUT-.t41 4.5005
R6728 VOUT-.n42 VOUT-.t145 4.5005
R6729 VOUT-.n44 VOUT-.t127 4.5005
R6730 VOUT-.n46 VOUT-.t74 4.5005
R6731 VOUT-.n45 VOUT-.t46 4.5005
R6732 VOUT-.n96 VOUT-.t27 4.5005
R6733 VOUT-.n97 VOUT-.t110 4.5005
R6734 VOUT-.n98 VOUT-.t79 4.5005
R6735 VOUT-.n99 VOUT-.t51 4.5005
R6736 VOUT-.n20 VOUT-.n19 4.5005
R6737 VOUT-.n102 VOUT-.t9 3.42907
R6738 VOUT-.n102 VOUT-.t11 3.42907
R6739 VOUT-.n104 VOUT-.t6 3.42907
R6740 VOUT-.n104 VOUT-.t4 3.42907
R6741 VOUT-.n107 VOUT-.t12 3.42907
R6742 VOUT-.n107 VOUT-.t0 3.42907
R6743 VOUT- VOUT-.n110 1.78175
R6744 VOUT-.n110 VOUT-.n109 1.69693
R6745 VOUT-.n20 VOUT-.n1 1.313
R6746 VOUT-.n109 VOUT-.n101 1.13443
R6747 VOUT-.n19 VOUT-.n2 0.563
R6748 VOUT-.n9 VOUT-.n2 0.563
R6749 VOUT-.n9 VOUT-.n8 0.563
R6750 VOUT-.n12 VOUT-.n3 0.563
R6751 VOUT-.n15 VOUT-.n12 0.563
R6752 VOUT-.n16 VOUT-.n15 0.563
R6753 VOUT-.n48 VOUT-.n47 0.3295
R6754 VOUT-.n57 VOUT-.n56 0.3295
R6755 VOUT-.n55 VOUT-.n54 0.3295
R6756 VOUT-.n53 VOUT-.n52 0.3295
R6757 VOUT-.n51 VOUT-.n50 0.3295
R6758 VOUT-.n68 VOUT-.n49 0.3295
R6759 VOUT-.n68 VOUT-.n67 0.3295
R6760 VOUT-.n67 VOUT-.n66 0.3295
R6761 VOUT-.n66 VOUT-.n65 0.3295
R6762 VOUT-.n65 VOUT-.n64 0.3295
R6763 VOUT-.n64 VOUT-.n63 0.3295
R6764 VOUT-.n63 VOUT-.n62 0.3295
R6765 VOUT-.n62 VOUT-.n61 0.3295
R6766 VOUT-.n61 VOUT-.n60 0.3295
R6767 VOUT-.n60 VOUT-.n59 0.3295
R6768 VOUT-.n59 VOUT-.n58 0.3295
R6769 VOUT-.n71 VOUT-.n69 0.3295
R6770 VOUT-.n71 VOUT-.n70 0.3295
R6771 VOUT-.n74 VOUT-.n72 0.3295
R6772 VOUT-.n74 VOUT-.n73 0.3295
R6773 VOUT-.n77 VOUT-.n75 0.3295
R6774 VOUT-.n77 VOUT-.n76 0.3295
R6775 VOUT-.n80 VOUT-.n78 0.3295
R6776 VOUT-.n80 VOUT-.n79 0.3295
R6777 VOUT-.n83 VOUT-.n81 0.3295
R6778 VOUT-.n83 VOUT-.n82 0.3295
R6779 VOUT-.n86 VOUT-.n84 0.3295
R6780 VOUT-.n86 VOUT-.n85 0.3295
R6781 VOUT-.n89 VOUT-.n87 0.3295
R6782 VOUT-.n89 VOUT-.n88 0.3295
R6783 VOUT-.n92 VOUT-.n90 0.3295
R6784 VOUT-.n92 VOUT-.n91 0.3295
R6785 VOUT-.n95 VOUT-.n93 0.3295
R6786 VOUT-.n95 VOUT-.n94 0.3295
R6787 VOUT-.n22 VOUT-.n21 0.3295
R6788 VOUT-.n34 VOUT-.n23 0.3295
R6789 VOUT-.n34 VOUT-.n33 0.3295
R6790 VOUT-.n33 VOUT-.n32 0.3295
R6791 VOUT-.n32 VOUT-.n31 0.3295
R6792 VOUT-.n31 VOUT-.n30 0.3295
R6793 VOUT-.n30 VOUT-.n29 0.3295
R6794 VOUT-.n29 VOUT-.n28 0.3295
R6795 VOUT-.n28 VOUT-.n27 0.3295
R6796 VOUT-.n27 VOUT-.n26 0.3295
R6797 VOUT-.n26 VOUT-.n25 0.3295
R6798 VOUT-.n25 VOUT-.n24 0.3295
R6799 VOUT-.n37 VOUT-.n35 0.3295
R6800 VOUT-.n37 VOUT-.n36 0.3295
R6801 VOUT-.n40 VOUT-.n38 0.3295
R6802 VOUT-.n40 VOUT-.n39 0.3295
R6803 VOUT-.n43 VOUT-.n41 0.3295
R6804 VOUT-.n43 VOUT-.n42 0.3295
R6805 VOUT-.n46 VOUT-.n44 0.3295
R6806 VOUT-.n46 VOUT-.n45 0.3295
R6807 VOUT-.n97 VOUT-.n96 0.3295
R6808 VOUT-.n98 VOUT-.n97 0.3295
R6809 VOUT-.n99 VOUT-.n98 0.3295
R6810 VOUT-.n62 VOUT-.n57 0.306
R6811 VOUT-.n63 VOUT-.n55 0.306
R6812 VOUT-.n64 VOUT-.n53 0.306
R6813 VOUT-.n65 VOUT-.n51 0.306
R6814 VOUT-.n68 VOUT-.n48 0.2825
R6815 VOUT-.n71 VOUT-.n68 0.2825
R6816 VOUT-.n74 VOUT-.n71 0.2825
R6817 VOUT-.n77 VOUT-.n74 0.2825
R6818 VOUT-.n80 VOUT-.n77 0.2825
R6819 VOUT-.n83 VOUT-.n80 0.2825
R6820 VOUT-.n86 VOUT-.n83 0.2825
R6821 VOUT-.n89 VOUT-.n86 0.2825
R6822 VOUT-.n92 VOUT-.n89 0.2825
R6823 VOUT-.n95 VOUT-.n92 0.2825
R6824 VOUT-.n34 VOUT-.n22 0.2825
R6825 VOUT-.n37 VOUT-.n34 0.2825
R6826 VOUT-.n40 VOUT-.n37 0.2825
R6827 VOUT-.n43 VOUT-.n40 0.2825
R6828 VOUT-.n46 VOUT-.n43 0.2825
R6829 VOUT-.n97 VOUT-.n46 0.2825
R6830 VOUT-.n97 VOUT-.n95 0.2825
R6831 two_stage_opamp_dummy_magic_23_0.cap_res_X.t0 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 50.1603
R6832 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 two_stage_opamp_dummy_magic_23_0.cap_res_X.t29 0.1603
R6833 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 two_stage_opamp_dummy_magic_23_0.cap_res_X.t53 0.1603
R6834 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 two_stage_opamp_dummy_magic_23_0.cap_res_X.t35 0.1603
R6835 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 two_stage_opamp_dummy_magic_23_0.cap_res_X.t134 0.1603
R6836 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t69 0.1603
R6837 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 0.1603
R6838 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 0.1603
R6839 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 two_stage_opamp_dummy_magic_23_0.cap_res_X.t40 0.1603
R6840 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 0.1603
R6841 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 0.1603
R6842 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 two_stage_opamp_dummy_magic_23_0.cap_res_X.t70 0.1603
R6843 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 two_stage_opamp_dummy_magic_23_0.cap_res_X.t101 0.1603
R6844 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t62 0.1603
R6845 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 two_stage_opamp_dummy_magic_23_0.cap_res_X.t107 0.1603
R6846 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 two_stage_opamp_dummy_magic_23_0.cap_res_X.t13 0.1603
R6847 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 two_stage_opamp_dummy_magic_23_0.cap_res_X.t138 0.1603
R6848 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t57 0.1603
R6849 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 two_stage_opamp_dummy_magic_23_0.cap_res_X.t43 0.1603
R6850 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 two_stage_opamp_dummy_magic_23_0.cap_res_X.t19 0.1603
R6851 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 two_stage_opamp_dummy_magic_23_0.cap_res_X.t3 0.1603
R6852 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t61 0.1603
R6853 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 two_stage_opamp_dummy_magic_23_0.cap_res_X.t49 0.1603
R6854 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 two_stage_opamp_dummy_magic_23_0.cap_res_X.t97 0.1603
R6855 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 two_stage_opamp_dummy_magic_23_0.cap_res_X.t85 0.1603
R6856 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t64 0.1603
R6857 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 two_stage_opamp_dummy_magic_23_0.cap_res_X.t52 0.1603
R6858 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 two_stage_opamp_dummy_magic_23_0.cap_res_X.t99 0.1603
R6859 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 two_stage_opamp_dummy_magic_23_0.cap_res_X.t89 0.1603
R6860 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 two_stage_opamp_dummy_magic_23_0.cap_res_X.t5 0.1603
R6861 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t129 0.1603
R6862 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 two_stage_opamp_dummy_magic_23_0.cap_res_X.t106 0.1603
R6863 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 two_stage_opamp_dummy_magic_23_0.cap_res_X.t95 0.1603
R6864 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 two_stage_opamp_dummy_magic_23_0.cap_res_X.t10 0.1603
R6865 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t135 0.1603
R6866 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t54 0.1603
R6867 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 two_stage_opamp_dummy_magic_23_0.cap_res_X.t37 0.1603
R6868 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 two_stage_opamp_dummy_magic_23_0.cap_res_X.t91 0.1603
R6869 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 two_stage_opamp_dummy_magic_23_0.cap_res_X.t72 0.1603
R6870 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t55 0.1603
R6871 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 two_stage_opamp_dummy_magic_23_0.cap_res_X.t44 0.1603
R6872 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 two_stage_opamp_dummy_magic_23_0.cap_res_X.t84 0.1603
R6873 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 two_stage_opamp_dummy_magic_23_0.cap_res_X.t36 0.1603
R6874 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 two_stage_opamp_dummy_magic_23_0.cap_res_X.t105 0.1603
R6875 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 two_stage_opamp_dummy_magic_23_0.cap_res_X.t76 0.1603
R6876 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t23 0.1603
R6877 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 two_stage_opamp_dummy_magic_23_0.cap_res_X.t128 0.1603
R6878 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 two_stage_opamp_dummy_magic_23_0.cap_res_X.t94 0.1603
R6879 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t59 0.1603
R6880 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 two_stage_opamp_dummy_magic_23_0.cap_res_X.t6 0.1603
R6881 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 two_stage_opamp_dummy_magic_23_0.cap_res_X.t109 0.1603
R6882 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 two_stage_opamp_dummy_magic_23_0.cap_res_X.t96 0.1603
R6883 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t133 0.1603
R6884 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 two_stage_opamp_dummy_magic_23_0.cap_res_X.t100 0.1603
R6885 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 0.1603
R6886 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 0.1603
R6887 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 0.1603
R6888 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 0.1603
R6889 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 0.1603
R6890 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 two_stage_opamp_dummy_magic_23_0.cap_res_X.t21 0.159278
R6891 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t50 0.159278
R6892 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t27 0.159278
R6893 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 two_stage_opamp_dummy_magic_23_0.cap_res_X.t127 0.159278
R6894 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t11 0.159278
R6895 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t108 0.159278
R6896 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 0.159278
R6897 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 0.159278
R6898 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 0.159278
R6899 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 0.159278
R6900 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 0.159278
R6901 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 0.159278
R6902 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 0.159278
R6903 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 0.159278
R6904 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 0.159278
R6905 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 0.159278
R6906 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 0.159278
R6907 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 0.159278
R6908 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 0.159278
R6909 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 0.159278
R6910 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 0.159278
R6911 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 0.159278
R6912 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 0.159278
R6913 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t20 0.159278
R6914 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 two_stage_opamp_dummy_magic_23_0.cap_res_X.t58 0.159278
R6915 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t41 0.159278
R6916 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 two_stage_opamp_dummy_magic_23_0.cap_res_X.t75 0.159278
R6917 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 0.137822
R6918 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 0.1368
R6919 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 0.1368
R6920 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 0.1368
R6921 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 0.1368
R6922 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 0.1368
R6923 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 0.1368
R6924 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 0.1368
R6925 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 0.1368
R6926 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 0.1368
R6927 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 0.1368
R6928 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 0.1368
R6929 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 0.1368
R6930 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 0.1368
R6931 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 0.1368
R6932 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 0.1368
R6933 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 0.1368
R6934 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 0.1368
R6935 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 0.1368
R6936 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 0.1368
R6937 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 0.1368
R6938 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 0.1368
R6939 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 0.1368
R6940 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 0.1368
R6941 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 0.1368
R6942 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 0.1368
R6943 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 0.1368
R6944 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 0.1368
R6945 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 0.1368
R6946 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 0.1368
R6947 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 0.1368
R6948 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 0.1368
R6949 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 0.114322
R6950 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 0.1133
R6951 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 0.1133
R6952 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 0.1133
R6953 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 0.1133
R6954 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 0.1133
R6955 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 0.1133
R6956 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 0.1133
R6957 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 0.1133
R6958 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 0.1133
R6959 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 0.1133
R6960 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 0.1133
R6961 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 0.1133
R6962 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 0.1133
R6963 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 0.1133
R6964 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 0.1133
R6965 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 0.1133
R6966 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 0.1133
R6967 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 0.1133
R6968 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 0.1133
R6969 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 0.00152174
R6970 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 0.00152174
R6971 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 0.00152174
R6972 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 0.00152174
R6973 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 0.00152174
R6974 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 0.00152174
R6975 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 0.00152174
R6976 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 0.00152174
R6977 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 0.00152174
R6978 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 0.00152174
R6979 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 0.00152174
R6980 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 0.00152174
R6981 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 0.00152174
R6982 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 0.00152174
R6983 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 0.00152174
R6984 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 two_stage_opamp_dummy_magic_23_0.cap_res_X.t80 0.00152174
R6985 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 0.00152174
R6986 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 0.00152174
R6987 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 0.00152174
R6988 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 0.00152174
R6989 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 0.00152174
R6990 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 0.00152174
R6991 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 0.00152174
R6992 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 0.00152174
R6993 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 0.00152174
R6994 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 0.00152174
R6995 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 0.00152174
R6996 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 0.00152174
R6997 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 0.00152174
R6998 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 0.00152174
R6999 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 0.00152174
R7000 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 0.00152174
R7001 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t123 0.00152174
R7002 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 two_stage_opamp_dummy_magic_23_0.cap_res_X.t22 0.00152174
R7003 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 0.00152174
R7004 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 0.00152174
R7005 two_stage_opamp_dummy_magic_23_0.Vb1.n24 two_stage_opamp_dummy_magic_23_0.Vb1.n23 611.782
R7006 two_stage_opamp_dummy_magic_23_0.Vb1.n15 two_stage_opamp_dummy_magic_23_0.Vb1.t16 449.868
R7007 two_stage_opamp_dummy_magic_23_0.Vb1.n6 two_stage_opamp_dummy_magic_23_0.Vb1.t6 449.868
R7008 two_stage_opamp_dummy_magic_23_0.Vb1.n5 two_stage_opamp_dummy_magic_23_0.Vb1.t0 449.868
R7009 two_stage_opamp_dummy_magic_23_0.Vb1.n34 two_stage_opamp_dummy_magic_23_0.Vb1.n33 310.392
R7010 two_stage_opamp_dummy_magic_23_0.Vb1.n33 two_stage_opamp_dummy_magic_23_0.Vb1.t31 273.134
R7011 two_stage_opamp_dummy_magic_23_0.Vb1.n24 two_stage_opamp_dummy_magic_23_0.Vb1.t17 273.134
R7012 two_stage_opamp_dummy_magic_23_0.Vb1.n23 two_stage_opamp_dummy_magic_23_0.Vb1.t15 273.134
R7013 two_stage_opamp_dummy_magic_23_0.Vb1.n22 two_stage_opamp_dummy_magic_23_0.Vb1.t25 273.134
R7014 two_stage_opamp_dummy_magic_23_0.Vb1.n21 two_stage_opamp_dummy_magic_23_0.Vb1.t14 273.134
R7015 two_stage_opamp_dummy_magic_23_0.Vb1.n20 two_stage_opamp_dummy_magic_23_0.Vb1.t23 273.134
R7016 two_stage_opamp_dummy_magic_23_0.Vb1.n19 two_stage_opamp_dummy_magic_23_0.Vb1.t32 273.134
R7017 two_stage_opamp_dummy_magic_23_0.Vb1.n18 two_stage_opamp_dummy_magic_23_0.Vb1.t24 273.134
R7018 two_stage_opamp_dummy_magic_23_0.Vb1.n17 two_stage_opamp_dummy_magic_23_0.Vb1.t12 273.134
R7019 two_stage_opamp_dummy_magic_23_0.Vb1.n16 two_stage_opamp_dummy_magic_23_0.Vb1.t22 273.134
R7020 two_stage_opamp_dummy_magic_23_0.Vb1.n15 two_stage_opamp_dummy_magic_23_0.Vb1.t30 273.134
R7021 two_stage_opamp_dummy_magic_23_0.Vb1.n32 two_stage_opamp_dummy_magic_23_0.Vb1.t21 273.134
R7022 two_stage_opamp_dummy_magic_23_0.Vb1.n31 two_stage_opamp_dummy_magic_23_0.Vb1.t29 273.134
R7023 two_stage_opamp_dummy_magic_23_0.Vb1.n30 two_stage_opamp_dummy_magic_23_0.Vb1.t20 273.134
R7024 two_stage_opamp_dummy_magic_23_0.Vb1.n29 two_stage_opamp_dummy_magic_23_0.Vb1.t28 273.134
R7025 two_stage_opamp_dummy_magic_23_0.Vb1.n28 two_stage_opamp_dummy_magic_23_0.Vb1.t18 273.134
R7026 two_stage_opamp_dummy_magic_23_0.Vb1.n27 two_stage_opamp_dummy_magic_23_0.Vb1.t13 273.134
R7027 two_stage_opamp_dummy_magic_23_0.Vb1.n26 two_stage_opamp_dummy_magic_23_0.Vb1.t19 273.134
R7028 two_stage_opamp_dummy_magic_23_0.Vb1.n25 two_stage_opamp_dummy_magic_23_0.Vb1.t27 273.134
R7029 two_stage_opamp_dummy_magic_23_0.Vb1.n6 two_stage_opamp_dummy_magic_23_0.Vb1.t2 273.134
R7030 two_stage_opamp_dummy_magic_23_0.Vb1.n5 two_stage_opamp_dummy_magic_23_0.Vb1.t4 273.134
R7031 bgr_11_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb1.n0 218.364
R7032 two_stage_opamp_dummy_magic_23_0.Vb1.n16 two_stage_opamp_dummy_magic_23_0.Vb1.n15 176.733
R7033 two_stage_opamp_dummy_magic_23_0.Vb1.n17 two_stage_opamp_dummy_magic_23_0.Vb1.n16 176.733
R7034 two_stage_opamp_dummy_magic_23_0.Vb1.n18 two_stage_opamp_dummy_magic_23_0.Vb1.n17 176.733
R7035 two_stage_opamp_dummy_magic_23_0.Vb1.n19 two_stage_opamp_dummy_magic_23_0.Vb1.n18 176.733
R7036 two_stage_opamp_dummy_magic_23_0.Vb1.n20 two_stage_opamp_dummy_magic_23_0.Vb1.n19 176.733
R7037 two_stage_opamp_dummy_magic_23_0.Vb1.n21 two_stage_opamp_dummy_magic_23_0.Vb1.n20 176.733
R7038 two_stage_opamp_dummy_magic_23_0.Vb1.n22 two_stage_opamp_dummy_magic_23_0.Vb1.n21 176.733
R7039 two_stage_opamp_dummy_magic_23_0.Vb1.n23 two_stage_opamp_dummy_magic_23_0.Vb1.n22 176.733
R7040 two_stage_opamp_dummy_magic_23_0.Vb1.n25 two_stage_opamp_dummy_magic_23_0.Vb1.n24 176.733
R7041 two_stage_opamp_dummy_magic_23_0.Vb1.n26 two_stage_opamp_dummy_magic_23_0.Vb1.n25 176.733
R7042 two_stage_opamp_dummy_magic_23_0.Vb1.n27 two_stage_opamp_dummy_magic_23_0.Vb1.n26 176.733
R7043 two_stage_opamp_dummy_magic_23_0.Vb1.n28 two_stage_opamp_dummy_magic_23_0.Vb1.n27 176.733
R7044 two_stage_opamp_dummy_magic_23_0.Vb1.n29 two_stage_opamp_dummy_magic_23_0.Vb1.n28 176.733
R7045 two_stage_opamp_dummy_magic_23_0.Vb1.n30 two_stage_opamp_dummy_magic_23_0.Vb1.n29 176.733
R7046 two_stage_opamp_dummy_magic_23_0.Vb1.n31 two_stage_opamp_dummy_magic_23_0.Vb1.n30 176.733
R7047 two_stage_opamp_dummy_magic_23_0.Vb1.n32 two_stage_opamp_dummy_magic_23_0.Vb1.n31 176.733
R7048 two_stage_opamp_dummy_magic_23_0.Vb1.n33 two_stage_opamp_dummy_magic_23_0.Vb1.n32 176.733
R7049 two_stage_opamp_dummy_magic_23_0.Vb1.n2 two_stage_opamp_dummy_magic_23_0.Vb1.t26 167.769
R7050 two_stage_opamp_dummy_magic_23_0.Vb1.n8 two_stage_opamp_dummy_magic_23_0.Vb1.n7 161.3
R7051 two_stage_opamp_dummy_magic_23_0.Vb1.n4 two_stage_opamp_dummy_magic_23_0.Vb1.n3 49.3505
R7052 two_stage_opamp_dummy_magic_23_0.Vb1.n10 two_stage_opamp_dummy_magic_23_0.Vb1.n9 49.3505
R7053 two_stage_opamp_dummy_magic_23_0.Vb1.n13 two_stage_opamp_dummy_magic_23_0.Vb1.n12 49.3505
R7054 two_stage_opamp_dummy_magic_23_0.Vb1.n7 two_stage_opamp_dummy_magic_23_0.Vb1.n6 45.5227
R7055 two_stage_opamp_dummy_magic_23_0.Vb1.n7 two_stage_opamp_dummy_magic_23_0.Vb1.n5 45.5227
R7056 bgr_11_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb1.n34 39.5734
R7057 two_stage_opamp_dummy_magic_23_0.Vb1.n0 two_stage_opamp_dummy_magic_23_0.Vb1.t11 19.7005
R7058 two_stage_opamp_dummy_magic_23_0.Vb1.n0 two_stage_opamp_dummy_magic_23_0.Vb1.t10 19.7005
R7059 two_stage_opamp_dummy_magic_23_0.Vb1.n34 two_stage_opamp_dummy_magic_23_0.Vb1.n14 17.8547
R7060 two_stage_opamp_dummy_magic_23_0.Vb1.n3 two_stage_opamp_dummy_magic_23_0.Vb1.t9 16.0005
R7061 two_stage_opamp_dummy_magic_23_0.Vb1.n3 two_stage_opamp_dummy_magic_23_0.Vb1.t1 16.0005
R7062 two_stage_opamp_dummy_magic_23_0.Vb1.n9 two_stage_opamp_dummy_magic_23_0.Vb1.t5 16.0005
R7063 two_stage_opamp_dummy_magic_23_0.Vb1.n9 two_stage_opamp_dummy_magic_23_0.Vb1.t3 16.0005
R7064 two_stage_opamp_dummy_magic_23_0.Vb1.n12 two_stage_opamp_dummy_magic_23_0.Vb1.t7 16.0005
R7065 two_stage_opamp_dummy_magic_23_0.Vb1.n12 two_stage_opamp_dummy_magic_23_0.Vb1.t8 16.0005
R7066 two_stage_opamp_dummy_magic_23_0.Vb1.n13 two_stage_opamp_dummy_magic_23_0.Vb1.n11 5.6255
R7067 two_stage_opamp_dummy_magic_23_0.Vb1.n11 two_stage_opamp_dummy_magic_23_0.Vb1.n4 5.6255
R7068 two_stage_opamp_dummy_magic_23_0.Vb1.n11 two_stage_opamp_dummy_magic_23_0.Vb1.n10 5.063
R7069 two_stage_opamp_dummy_magic_23_0.Vb1.n14 two_stage_opamp_dummy_magic_23_0.Vb1.n13 4.938
R7070 two_stage_opamp_dummy_magic_23_0.Vb1.n4 two_stage_opamp_dummy_magic_23_0.Vb1.n2 4.938
R7071 two_stage_opamp_dummy_magic_23_0.Vb1.n8 two_stage_opamp_dummy_magic_23_0.Vb1.n1 4.5005
R7072 two_stage_opamp_dummy_magic_23_0.Vb1.n2 two_stage_opamp_dummy_magic_23_0.Vb1.n1 0.563
R7073 two_stage_opamp_dummy_magic_23_0.Vb1.n14 two_stage_opamp_dummy_magic_23_0.Vb1.n1 0.563
R7074 two_stage_opamp_dummy_magic_23_0.Vb1.n10 two_stage_opamp_dummy_magic_23_0.Vb1.n8 0.438
R7075 two_stage_opamp_dummy_magic_23_0.X.n27 two_stage_opamp_dummy_magic_23_0.X.t46 1172.87
R7076 two_stage_opamp_dummy_magic_23_0.X.n21 two_stage_opamp_dummy_magic_23_0.X.t39 1172.87
R7077 two_stage_opamp_dummy_magic_23_0.X.n27 two_stage_opamp_dummy_magic_23_0.X.t31 996.134
R7078 two_stage_opamp_dummy_magic_23_0.X.n28 two_stage_opamp_dummy_magic_23_0.X.t48 996.134
R7079 two_stage_opamp_dummy_magic_23_0.X.n26 two_stage_opamp_dummy_magic_23_0.X.t34 996.134
R7080 two_stage_opamp_dummy_magic_23_0.X.n25 two_stage_opamp_dummy_magic_23_0.X.t51 996.134
R7081 two_stage_opamp_dummy_magic_23_0.X.n24 two_stage_opamp_dummy_magic_23_0.X.t37 996.134
R7082 two_stage_opamp_dummy_magic_23_0.X.n23 two_stage_opamp_dummy_magic_23_0.X.t53 996.134
R7083 two_stage_opamp_dummy_magic_23_0.X.n22 two_stage_opamp_dummy_magic_23_0.X.t36 996.134
R7084 two_stage_opamp_dummy_magic_23_0.X.n21 two_stage_opamp_dummy_magic_23_0.X.t52 996.134
R7085 two_stage_opamp_dummy_magic_23_0.X.n62 two_stage_opamp_dummy_magic_23_0.X.t41 690.867
R7086 two_stage_opamp_dummy_magic_23_0.X.n61 two_stage_opamp_dummy_magic_23_0.X.t35 690.867
R7087 two_stage_opamp_dummy_magic_23_0.X.n53 two_stage_opamp_dummy_magic_23_0.X.t38 530.201
R7088 two_stage_opamp_dummy_magic_23_0.X.n52 two_stage_opamp_dummy_magic_23_0.X.t30 530.201
R7089 two_stage_opamp_dummy_magic_23_0.X.n68 two_stage_opamp_dummy_magic_23_0.X.t32 514.134
R7090 two_stage_opamp_dummy_magic_23_0.X.n67 two_stage_opamp_dummy_magic_23_0.X.t50 514.134
R7091 two_stage_opamp_dummy_magic_23_0.X.n66 two_stage_opamp_dummy_magic_23_0.X.t33 514.134
R7092 two_stage_opamp_dummy_magic_23_0.X.n65 two_stage_opamp_dummy_magic_23_0.X.t47 514.134
R7093 two_stage_opamp_dummy_magic_23_0.X.n64 two_stage_opamp_dummy_magic_23_0.X.t29 514.134
R7094 two_stage_opamp_dummy_magic_23_0.X.n63 two_stage_opamp_dummy_magic_23_0.X.t43 514.134
R7095 two_stage_opamp_dummy_magic_23_0.X.n62 two_stage_opamp_dummy_magic_23_0.X.t26 514.134
R7096 two_stage_opamp_dummy_magic_23_0.X.n61 two_stage_opamp_dummy_magic_23_0.X.t49 514.134
R7097 two_stage_opamp_dummy_magic_23_0.X.n53 two_stage_opamp_dummy_magic_23_0.X.t54 353.467
R7098 two_stage_opamp_dummy_magic_23_0.X.n54 two_stage_opamp_dummy_magic_23_0.X.t40 353.467
R7099 two_stage_opamp_dummy_magic_23_0.X.n55 two_stage_opamp_dummy_magic_23_0.X.t25 353.467
R7100 two_stage_opamp_dummy_magic_23_0.X.n56 two_stage_opamp_dummy_magic_23_0.X.t42 353.467
R7101 two_stage_opamp_dummy_magic_23_0.X.n57 two_stage_opamp_dummy_magic_23_0.X.t28 353.467
R7102 two_stage_opamp_dummy_magic_23_0.X.n58 two_stage_opamp_dummy_magic_23_0.X.t45 353.467
R7103 two_stage_opamp_dummy_magic_23_0.X.n59 two_stage_opamp_dummy_magic_23_0.X.t27 353.467
R7104 two_stage_opamp_dummy_magic_23_0.X.n52 two_stage_opamp_dummy_magic_23_0.X.t44 353.467
R7105 two_stage_opamp_dummy_magic_23_0.X.n30 two_stage_opamp_dummy_magic_23_0.X.n29 304.375
R7106 two_stage_opamp_dummy_magic_23_0.X.n70 two_stage_opamp_dummy_magic_23_0.X.n60 216.9
R7107 two_stage_opamp_dummy_magic_23_0.X.n70 two_stage_opamp_dummy_magic_23_0.X.n69 216.9
R7108 two_stage_opamp_dummy_magic_23_0.X.n26 two_stage_opamp_dummy_magic_23_0.X.n25 176.733
R7109 two_stage_opamp_dummy_magic_23_0.X.n25 two_stage_opamp_dummy_magic_23_0.X.n24 176.733
R7110 two_stage_opamp_dummy_magic_23_0.X.n24 two_stage_opamp_dummy_magic_23_0.X.n23 176.733
R7111 two_stage_opamp_dummy_magic_23_0.X.n23 two_stage_opamp_dummy_magic_23_0.X.n22 176.733
R7112 two_stage_opamp_dummy_magic_23_0.X.n22 two_stage_opamp_dummy_magic_23_0.X.n21 176.733
R7113 two_stage_opamp_dummy_magic_23_0.X.n28 two_stage_opamp_dummy_magic_23_0.X.n27 176.733
R7114 two_stage_opamp_dummy_magic_23_0.X.n54 two_stage_opamp_dummy_magic_23_0.X.n53 176.733
R7115 two_stage_opamp_dummy_magic_23_0.X.n55 two_stage_opamp_dummy_magic_23_0.X.n54 176.733
R7116 two_stage_opamp_dummy_magic_23_0.X.n56 two_stage_opamp_dummy_magic_23_0.X.n55 176.733
R7117 two_stage_opamp_dummy_magic_23_0.X.n57 two_stage_opamp_dummy_magic_23_0.X.n56 176.733
R7118 two_stage_opamp_dummy_magic_23_0.X.n58 two_stage_opamp_dummy_magic_23_0.X.n57 176.733
R7119 two_stage_opamp_dummy_magic_23_0.X.n59 two_stage_opamp_dummy_magic_23_0.X.n58 176.733
R7120 two_stage_opamp_dummy_magic_23_0.X.n63 two_stage_opamp_dummy_magic_23_0.X.n62 176.733
R7121 two_stage_opamp_dummy_magic_23_0.X.n64 two_stage_opamp_dummy_magic_23_0.X.n63 176.733
R7122 two_stage_opamp_dummy_magic_23_0.X.n65 two_stage_opamp_dummy_magic_23_0.X.n64 176.733
R7123 two_stage_opamp_dummy_magic_23_0.X.n66 two_stage_opamp_dummy_magic_23_0.X.n65 176.733
R7124 two_stage_opamp_dummy_magic_23_0.X.n67 two_stage_opamp_dummy_magic_23_0.X.n66 176.733
R7125 two_stage_opamp_dummy_magic_23_0.X.n68 two_stage_opamp_dummy_magic_23_0.X.n67 176.733
R7126 two_stage_opamp_dummy_magic_23_0.X.n71 two_stage_opamp_dummy_magic_23_0.X.n70 175.05
R7127 two_stage_opamp_dummy_magic_23_0.X.n32 two_stage_opamp_dummy_magic_23_0.X.n31 66.0338
R7128 two_stage_opamp_dummy_magic_23_0.X.n36 two_stage_opamp_dummy_magic_23_0.X.n35 66.0338
R7129 two_stage_opamp_dummy_magic_23_0.X.n38 two_stage_opamp_dummy_magic_23_0.X.n37 66.0338
R7130 two_stage_opamp_dummy_magic_23_0.X.n42 two_stage_opamp_dummy_magic_23_0.X.n41 66.0338
R7131 two_stage_opamp_dummy_magic_23_0.X.n45 two_stage_opamp_dummy_magic_23_0.X.n44 66.0338
R7132 two_stage_opamp_dummy_magic_23_0.X.n49 two_stage_opamp_dummy_magic_23_0.X.n48 66.0338
R7133 two_stage_opamp_dummy_magic_23_0.X.n30 two_stage_opamp_dummy_magic_23_0.X.t3 49.4481
R7134 two_stage_opamp_dummy_magic_23_0.X.n1 two_stage_opamp_dummy_magic_23_0.X.n0 49.3505
R7135 two_stage_opamp_dummy_magic_23_0.X.n5 two_stage_opamp_dummy_magic_23_0.X.n4 49.3505
R7136 two_stage_opamp_dummy_magic_23_0.X.n7 two_stage_opamp_dummy_magic_23_0.X.n6 49.3505
R7137 two_stage_opamp_dummy_magic_23_0.X.n11 two_stage_opamp_dummy_magic_23_0.X.n10 49.3505
R7138 two_stage_opamp_dummy_magic_23_0.X.n13 two_stage_opamp_dummy_magic_23_0.X.n12 49.3505
R7139 two_stage_opamp_dummy_magic_23_0.X.n17 two_stage_opamp_dummy_magic_23_0.X.n16 49.3505
R7140 two_stage_opamp_dummy_magic_23_0.X.n29 two_stage_opamp_dummy_magic_23_0.X.n26 40.1672
R7141 two_stage_opamp_dummy_magic_23_0.X.n29 two_stage_opamp_dummy_magic_23_0.X.n28 40.1672
R7142 two_stage_opamp_dummy_magic_23_0.X.n60 two_stage_opamp_dummy_magic_23_0.X.n52 40.1672
R7143 two_stage_opamp_dummy_magic_23_0.X.n60 two_stage_opamp_dummy_magic_23_0.X.n59 40.1672
R7144 two_stage_opamp_dummy_magic_23_0.X.n69 two_stage_opamp_dummy_magic_23_0.X.n61 40.1672
R7145 two_stage_opamp_dummy_magic_23_0.X.n69 two_stage_opamp_dummy_magic_23_0.X.n68 40.1672
R7146 two_stage_opamp_dummy_magic_23_0.X.n71 two_stage_opamp_dummy_magic_23_0.X.n51 17.688
R7147 two_stage_opamp_dummy_magic_23_0.X.n0 two_stage_opamp_dummy_magic_23_0.X.t4 16.0005
R7148 two_stage_opamp_dummy_magic_23_0.X.n0 two_stage_opamp_dummy_magic_23_0.X.t10 16.0005
R7149 two_stage_opamp_dummy_magic_23_0.X.n4 two_stage_opamp_dummy_magic_23_0.X.t24 16.0005
R7150 two_stage_opamp_dummy_magic_23_0.X.n4 two_stage_opamp_dummy_magic_23_0.X.t13 16.0005
R7151 two_stage_opamp_dummy_magic_23_0.X.n6 two_stage_opamp_dummy_magic_23_0.X.t8 16.0005
R7152 two_stage_opamp_dummy_magic_23_0.X.n6 two_stage_opamp_dummy_magic_23_0.X.t12 16.0005
R7153 two_stage_opamp_dummy_magic_23_0.X.n10 two_stage_opamp_dummy_magic_23_0.X.t5 16.0005
R7154 two_stage_opamp_dummy_magic_23_0.X.n10 two_stage_opamp_dummy_magic_23_0.X.t23 16.0005
R7155 two_stage_opamp_dummy_magic_23_0.X.n12 two_stage_opamp_dummy_magic_23_0.X.t6 16.0005
R7156 two_stage_opamp_dummy_magic_23_0.X.n12 two_stage_opamp_dummy_magic_23_0.X.t9 16.0005
R7157 two_stage_opamp_dummy_magic_23_0.X.n16 two_stage_opamp_dummy_magic_23_0.X.t7 16.0005
R7158 two_stage_opamp_dummy_magic_23_0.X.n16 two_stage_opamp_dummy_magic_23_0.X.t11 16.0005
R7159 two_stage_opamp_dummy_magic_23_0.X.n31 two_stage_opamp_dummy_magic_23_0.X.t15 11.2576
R7160 two_stage_opamp_dummy_magic_23_0.X.n31 two_stage_opamp_dummy_magic_23_0.X.t17 11.2576
R7161 two_stage_opamp_dummy_magic_23_0.X.n35 two_stage_opamp_dummy_magic_23_0.X.t18 11.2576
R7162 two_stage_opamp_dummy_magic_23_0.X.n35 two_stage_opamp_dummy_magic_23_0.X.t20 11.2576
R7163 two_stage_opamp_dummy_magic_23_0.X.n37 two_stage_opamp_dummy_magic_23_0.X.t0 11.2576
R7164 two_stage_opamp_dummy_magic_23_0.X.n37 two_stage_opamp_dummy_magic_23_0.X.t21 11.2576
R7165 two_stage_opamp_dummy_magic_23_0.X.n41 two_stage_opamp_dummy_magic_23_0.X.t16 11.2576
R7166 two_stage_opamp_dummy_magic_23_0.X.n41 two_stage_opamp_dummy_magic_23_0.X.t22 11.2576
R7167 two_stage_opamp_dummy_magic_23_0.X.n44 two_stage_opamp_dummy_magic_23_0.X.t1 11.2576
R7168 two_stage_opamp_dummy_magic_23_0.X.n44 two_stage_opamp_dummy_magic_23_0.X.t14 11.2576
R7169 two_stage_opamp_dummy_magic_23_0.X.n48 two_stage_opamp_dummy_magic_23_0.X.t2 11.2576
R7170 two_stage_opamp_dummy_magic_23_0.X.n48 two_stage_opamp_dummy_magic_23_0.X.t19 11.2576
R7171 two_stage_opamp_dummy_magic_23_0.X.n73 two_stage_opamp_dummy_magic_23_0.X.n72 8.09425
R7172 two_stage_opamp_dummy_magic_23_0.X.n39 two_stage_opamp_dummy_magic_23_0.X.n36 5.91717
R7173 two_stage_opamp_dummy_magic_23_0.X.n36 two_stage_opamp_dummy_magic_23_0.X.n34 5.91717
R7174 two_stage_opamp_dummy_magic_23_0.X.n47 two_stage_opamp_dummy_magic_23_0.X.n32 5.91717
R7175 two_stage_opamp_dummy_magic_23_0.X.n14 two_stage_opamp_dummy_magic_23_0.X.n11 5.6255
R7176 two_stage_opamp_dummy_magic_23_0.X.n8 two_stage_opamp_dummy_magic_23_0.X.n5 5.6255
R7177 two_stage_opamp_dummy_magic_23_0.X.n11 two_stage_opamp_dummy_magic_23_0.X.n3 5.438
R7178 two_stage_opamp_dummy_magic_23_0.X.n5 two_stage_opamp_dummy_magic_23_0.X.n2 5.438
R7179 two_stage_opamp_dummy_magic_23_0.X.n38 two_stage_opamp_dummy_magic_23_0.X.n34 5.29217
R7180 two_stage_opamp_dummy_magic_23_0.X.n39 two_stage_opamp_dummy_magic_23_0.X.n38 5.29217
R7181 two_stage_opamp_dummy_magic_23_0.X.n43 two_stage_opamp_dummy_magic_23_0.X.n42 5.29217
R7182 two_stage_opamp_dummy_magic_23_0.X.n42 two_stage_opamp_dummy_magic_23_0.X.n40 5.29217
R7183 two_stage_opamp_dummy_magic_23_0.X.n46 two_stage_opamp_dummy_magic_23_0.X.n45 5.29217
R7184 two_stage_opamp_dummy_magic_23_0.X.n45 two_stage_opamp_dummy_magic_23_0.X.n33 5.29217
R7185 two_stage_opamp_dummy_magic_23_0.X.n49 two_stage_opamp_dummy_magic_23_0.X.n47 5.29217
R7186 two_stage_opamp_dummy_magic_23_0.X.n50 two_stage_opamp_dummy_magic_23_0.X.n49 5.29217
R7187 two_stage_opamp_dummy_magic_23_0.X.n51 two_stage_opamp_dummy_magic_23_0.X.n50 5.1255
R7188 two_stage_opamp_dummy_magic_23_0.X.n8 two_stage_opamp_dummy_magic_23_0.X.n7 5.063
R7189 two_stage_opamp_dummy_magic_23_0.X.n14 two_stage_opamp_dummy_magic_23_0.X.n13 5.063
R7190 two_stage_opamp_dummy_magic_23_0.X.n17 two_stage_opamp_dummy_magic_23_0.X.n15 5.063
R7191 two_stage_opamp_dummy_magic_23_0.X.n9 two_stage_opamp_dummy_magic_23_0.X.n1 5.063
R7192 two_stage_opamp_dummy_magic_23_0.X.n7 two_stage_opamp_dummy_magic_23_0.X.n2 4.8755
R7193 two_stage_opamp_dummy_magic_23_0.X.n13 two_stage_opamp_dummy_magic_23_0.X.n3 4.8755
R7194 two_stage_opamp_dummy_magic_23_0.X.n18 two_stage_opamp_dummy_magic_23_0.X.n17 4.8755
R7195 two_stage_opamp_dummy_magic_23_0.X.n20 two_stage_opamp_dummy_magic_23_0.X.n19 4.5005
R7196 two_stage_opamp_dummy_magic_23_0.X.n72 two_stage_opamp_dummy_magic_23_0.X.n71 4.5005
R7197 two_stage_opamp_dummy_magic_23_0.X.n72 two_stage_opamp_dummy_magic_23_0.X.n30 3.27133
R7198 two_stage_opamp_dummy_magic_23_0.X.n73 two_stage_opamp_dummy_magic_23_0.X.n20 2.15675
R7199 two_stage_opamp_dummy_magic_23_0.X.n51 two_stage_opamp_dummy_magic_23_0.X.n32 0.792167
R7200 two_stage_opamp_dummy_magic_23_0.X.n50 two_stage_opamp_dummy_magic_23_0.X.n33 0.6255
R7201 two_stage_opamp_dummy_magic_23_0.X.n40 two_stage_opamp_dummy_magic_23_0.X.n33 0.6255
R7202 two_stage_opamp_dummy_magic_23_0.X.n40 two_stage_opamp_dummy_magic_23_0.X.n39 0.6255
R7203 two_stage_opamp_dummy_magic_23_0.X.n43 two_stage_opamp_dummy_magic_23_0.X.n34 0.6255
R7204 two_stage_opamp_dummy_magic_23_0.X.n46 two_stage_opamp_dummy_magic_23_0.X.n43 0.6255
R7205 two_stage_opamp_dummy_magic_23_0.X.n47 two_stage_opamp_dummy_magic_23_0.X.n46 0.6255
R7206 two_stage_opamp_dummy_magic_23_0.X.n15 two_stage_opamp_dummy_magic_23_0.X.n9 0.563
R7207 two_stage_opamp_dummy_magic_23_0.X.n15 two_stage_opamp_dummy_magic_23_0.X.n14 0.563
R7208 two_stage_opamp_dummy_magic_23_0.X.n18 two_stage_opamp_dummy_magic_23_0.X.n3 0.563
R7209 two_stage_opamp_dummy_magic_23_0.X.n19 two_stage_opamp_dummy_magic_23_0.X.n18 0.563
R7210 two_stage_opamp_dummy_magic_23_0.X.n19 two_stage_opamp_dummy_magic_23_0.X.n2 0.563
R7211 two_stage_opamp_dummy_magic_23_0.X.n9 two_stage_opamp_dummy_magic_23_0.X.n8 0.563
R7212 two_stage_opamp_dummy_magic_23_0.X.n20 two_stage_opamp_dummy_magic_23_0.X.n1 0.3755
R7213 two_stage_opamp_dummy_magic_23_0.X two_stage_opamp_dummy_magic_23_0.X.n73 0.063
R7214 two_stage_opamp_dummy_magic_23_0.VD1.n2 two_stage_opamp_dummy_magic_23_0.VD1.n1 49.3505
R7215 two_stage_opamp_dummy_magic_23_0.VD1.n5 two_stage_opamp_dummy_magic_23_0.VD1.n4 49.3505
R7216 two_stage_opamp_dummy_magic_23_0.VD1.n7 two_stage_opamp_dummy_magic_23_0.VD1.n6 49.3505
R7217 two_stage_opamp_dummy_magic_23_0.VD1.n11 two_stage_opamp_dummy_magic_23_0.VD1.n10 49.3505
R7218 two_stage_opamp_dummy_magic_23_0.VD1.n15 two_stage_opamp_dummy_magic_23_0.VD1.n14 49.3505
R7219 two_stage_opamp_dummy_magic_23_0.VD1.n18 two_stage_opamp_dummy_magic_23_0.VD1.n17 49.3505
R7220 two_stage_opamp_dummy_magic_23_0.VD1.n21 two_stage_opamp_dummy_magic_23_0.VD1.n20 49.3505
R7221 two_stage_opamp_dummy_magic_23_0.VD1.n24 two_stage_opamp_dummy_magic_23_0.VD1.n23 49.3505
R7222 two_stage_opamp_dummy_magic_23_0.VD1.n26 two_stage_opamp_dummy_magic_23_0.VD1.n25 49.3505
R7223 two_stage_opamp_dummy_magic_23_0.VD1.n30 two_stage_opamp_dummy_magic_23_0.VD1.n29 49.3505
R7224 two_stage_opamp_dummy_magic_23_0.VD1.n37 two_stage_opamp_dummy_magic_23_0.VD1.n36 49.3505
R7225 two_stage_opamp_dummy_magic_23_0.VD1.n1 two_stage_opamp_dummy_magic_23_0.VD1.t7 16.0005
R7226 two_stage_opamp_dummy_magic_23_0.VD1.n1 two_stage_opamp_dummy_magic_23_0.VD1.t2 16.0005
R7227 two_stage_opamp_dummy_magic_23_0.VD1.n4 two_stage_opamp_dummy_magic_23_0.VD1.t3 16.0005
R7228 two_stage_opamp_dummy_magic_23_0.VD1.n4 two_stage_opamp_dummy_magic_23_0.VD1.t8 16.0005
R7229 two_stage_opamp_dummy_magic_23_0.VD1.n6 two_stage_opamp_dummy_magic_23_0.VD1.t5 16.0005
R7230 two_stage_opamp_dummy_magic_23_0.VD1.n6 two_stage_opamp_dummy_magic_23_0.VD1.t9 16.0005
R7231 two_stage_opamp_dummy_magic_23_0.VD1.n10 two_stage_opamp_dummy_magic_23_0.VD1.t4 16.0005
R7232 two_stage_opamp_dummy_magic_23_0.VD1.n10 two_stage_opamp_dummy_magic_23_0.VD1.t1 16.0005
R7233 two_stage_opamp_dummy_magic_23_0.VD1.n14 two_stage_opamp_dummy_magic_23_0.VD1.t20 16.0005
R7234 two_stage_opamp_dummy_magic_23_0.VD1.n14 two_stage_opamp_dummy_magic_23_0.VD1.t15 16.0005
R7235 two_stage_opamp_dummy_magic_23_0.VD1.n17 two_stage_opamp_dummy_magic_23_0.VD1.t14 16.0005
R7236 two_stage_opamp_dummy_magic_23_0.VD1.n17 two_stage_opamp_dummy_magic_23_0.VD1.t16 16.0005
R7237 two_stage_opamp_dummy_magic_23_0.VD1.n20 two_stage_opamp_dummy_magic_23_0.VD1.t21 16.0005
R7238 two_stage_opamp_dummy_magic_23_0.VD1.n20 two_stage_opamp_dummy_magic_23_0.VD1.t18 16.0005
R7239 two_stage_opamp_dummy_magic_23_0.VD1.n23 two_stage_opamp_dummy_magic_23_0.VD1.t13 16.0005
R7240 two_stage_opamp_dummy_magic_23_0.VD1.n23 two_stage_opamp_dummy_magic_23_0.VD1.t19 16.0005
R7241 two_stage_opamp_dummy_magic_23_0.VD1.n25 two_stage_opamp_dummy_magic_23_0.VD1.t0 16.0005
R7242 two_stage_opamp_dummy_magic_23_0.VD1.n25 two_stage_opamp_dummy_magic_23_0.VD1.t12 16.0005
R7243 two_stage_opamp_dummy_magic_23_0.VD1.n29 two_stage_opamp_dummy_magic_23_0.VD1.t11 16.0005
R7244 two_stage_opamp_dummy_magic_23_0.VD1.n29 two_stage_opamp_dummy_magic_23_0.VD1.t17 16.0005
R7245 two_stage_opamp_dummy_magic_23_0.VD1.n37 two_stage_opamp_dummy_magic_23_0.VD1.t6 16.0005
R7246 two_stage_opamp_dummy_magic_23_0.VD1.t10 two_stage_opamp_dummy_magic_23_0.VD1.n37 16.0005
R7247 two_stage_opamp_dummy_magic_23_0.VD1.n33 two_stage_opamp_dummy_magic_23_0.VD1.n32 5.77133
R7248 two_stage_opamp_dummy_magic_23_0.VD1.n24 two_stage_opamp_dummy_magic_23_0.VD1.n13 5.64633
R7249 two_stage_opamp_dummy_magic_23_0.VD1.n16 two_stage_opamp_dummy_magic_23_0.VD1.n15 5.64633
R7250 two_stage_opamp_dummy_magic_23_0.VD1.n8 two_stage_opamp_dummy_magic_23_0.VD1.n5 5.6255
R7251 two_stage_opamp_dummy_magic_23_0.VD1.n2 two_stage_opamp_dummy_magic_23_0.VD1.n0 5.6255
R7252 two_stage_opamp_dummy_magic_23_0.VD1.n27 two_stage_opamp_dummy_magic_23_0.VD1.n24 5.438
R7253 two_stage_opamp_dummy_magic_23_0.VD1.n19 two_stage_opamp_dummy_magic_23_0.VD1.n15 5.438
R7254 two_stage_opamp_dummy_magic_23_0.VD1.n5 two_stage_opamp_dummy_magic_23_0.VD1.n3 5.438
R7255 two_stage_opamp_dummy_magic_23_0.VD1.n35 two_stage_opamp_dummy_magic_23_0.VD1.n2 5.438
R7256 two_stage_opamp_dummy_magic_23_0.VD1.n18 two_stage_opamp_dummy_magic_23_0.VD1.n16 5.08383
R7257 two_stage_opamp_dummy_magic_23_0.VD1.n21 two_stage_opamp_dummy_magic_23_0.VD1.n12 5.08383
R7258 two_stage_opamp_dummy_magic_23_0.VD1.n26 two_stage_opamp_dummy_magic_23_0.VD1.n13 5.08383
R7259 two_stage_opamp_dummy_magic_23_0.VD1.n31 two_stage_opamp_dummy_magic_23_0.VD1.n30 5.08383
R7260 two_stage_opamp_dummy_magic_23_0.VD1.n36 two_stage_opamp_dummy_magic_23_0.VD1.n0 5.063
R7261 two_stage_opamp_dummy_magic_23_0.VD1.n8 two_stage_opamp_dummy_magic_23_0.VD1.n7 5.063
R7262 two_stage_opamp_dummy_magic_23_0.VD1.n11 two_stage_opamp_dummy_magic_23_0.VD1.n9 5.063
R7263 two_stage_opamp_dummy_magic_23_0.VD1.n7 two_stage_opamp_dummy_magic_23_0.VD1.n3 4.8755
R7264 two_stage_opamp_dummy_magic_23_0.VD1.n19 two_stage_opamp_dummy_magic_23_0.VD1.n18 4.8755
R7265 two_stage_opamp_dummy_magic_23_0.VD1.n22 two_stage_opamp_dummy_magic_23_0.VD1.n21 4.8755
R7266 two_stage_opamp_dummy_magic_23_0.VD1.n27 two_stage_opamp_dummy_magic_23_0.VD1.n26 4.8755
R7267 two_stage_opamp_dummy_magic_23_0.VD1.n30 two_stage_opamp_dummy_magic_23_0.VD1.n28 4.8755
R7268 two_stage_opamp_dummy_magic_23_0.VD1.n36 two_stage_opamp_dummy_magic_23_0.VD1.n35 4.8755
R7269 two_stage_opamp_dummy_magic_23_0.VD1.n34 two_stage_opamp_dummy_magic_23_0.VD1.n33 4.5005
R7270 two_stage_opamp_dummy_magic_23_0.VD1.n31 two_stage_opamp_dummy_magic_23_0.VD1.n13 0.563
R7271 two_stage_opamp_dummy_magic_23_0.VD1.n28 two_stage_opamp_dummy_magic_23_0.VD1.n27 0.563
R7272 two_stage_opamp_dummy_magic_23_0.VD1.n28 two_stage_opamp_dummy_magic_23_0.VD1.n22 0.563
R7273 two_stage_opamp_dummy_magic_23_0.VD1.n22 two_stage_opamp_dummy_magic_23_0.VD1.n19 0.563
R7274 two_stage_opamp_dummy_magic_23_0.VD1.n16 two_stage_opamp_dummy_magic_23_0.VD1.n12 0.563
R7275 two_stage_opamp_dummy_magic_23_0.VD1.n35 two_stage_opamp_dummy_magic_23_0.VD1.n34 0.563
R7276 two_stage_opamp_dummy_magic_23_0.VD1.n34 two_stage_opamp_dummy_magic_23_0.VD1.n3 0.563
R7277 two_stage_opamp_dummy_magic_23_0.VD1.n9 two_stage_opamp_dummy_magic_23_0.VD1.n8 0.563
R7278 two_stage_opamp_dummy_magic_23_0.VD1.n9 two_stage_opamp_dummy_magic_23_0.VD1.n0 0.563
R7279 two_stage_opamp_dummy_magic_23_0.VD1.n33 two_stage_opamp_dummy_magic_23_0.VD1.n11 0.3755
R7280 two_stage_opamp_dummy_magic_23_0.VD1.n32 two_stage_opamp_dummy_magic_23_0.VD1.n31 0.234875
R7281 two_stage_opamp_dummy_magic_23_0.VD1.n32 two_stage_opamp_dummy_magic_23_0.VD1.n12 0.234875
R7282 two_stage_opamp_dummy_magic_23_0.Vb2.n23 two_stage_opamp_dummy_magic_23_0.Vb2.t15 746.673
R7283 two_stage_opamp_dummy_magic_23_0.Vb2.n1 two_stage_opamp_dummy_magic_23_0.Vb2.t9 721.625
R7284 two_stage_opamp_dummy_magic_23_0.Vb2.n16 two_stage_opamp_dummy_magic_23_0.Vb2.t30 611.739
R7285 two_stage_opamp_dummy_magic_23_0.Vb2.n12 two_stage_opamp_dummy_magic_23_0.Vb2.t24 611.739
R7286 two_stage_opamp_dummy_magic_23_0.Vb2.n7 two_stage_opamp_dummy_magic_23_0.Vb2.t19 611.739
R7287 two_stage_opamp_dummy_magic_23_0.Vb2.n3 two_stage_opamp_dummy_magic_23_0.Vb2.t16 611.739
R7288 two_stage_opamp_dummy_magic_23_0.Vb2.n2 two_stage_opamp_dummy_magic_23_0.Vb2.t31 563.451
R7289 two_stage_opamp_dummy_magic_23_0.Vb2.n16 two_stage_opamp_dummy_magic_23_0.Vb2.t27 421.75
R7290 two_stage_opamp_dummy_magic_23_0.Vb2.n17 two_stage_opamp_dummy_magic_23_0.Vb2.t22 421.75
R7291 two_stage_opamp_dummy_magic_23_0.Vb2.n18 two_stage_opamp_dummy_magic_23_0.Vb2.t18 421.75
R7292 two_stage_opamp_dummy_magic_23_0.Vb2.n19 two_stage_opamp_dummy_magic_23_0.Vb2.t12 421.75
R7293 two_stage_opamp_dummy_magic_23_0.Vb2.n12 two_stage_opamp_dummy_magic_23_0.Vb2.t20 421.75
R7294 two_stage_opamp_dummy_magic_23_0.Vb2.n13 two_stage_opamp_dummy_magic_23_0.Vb2.t25 421.75
R7295 two_stage_opamp_dummy_magic_23_0.Vb2.n14 two_stage_opamp_dummy_magic_23_0.Vb2.t29 421.75
R7296 two_stage_opamp_dummy_magic_23_0.Vb2.n15 two_stage_opamp_dummy_magic_23_0.Vb2.t32 421.75
R7297 two_stage_opamp_dummy_magic_23_0.Vb2.n7 two_stage_opamp_dummy_magic_23_0.Vb2.t14 421.75
R7298 two_stage_opamp_dummy_magic_23_0.Vb2.n8 two_stage_opamp_dummy_magic_23_0.Vb2.t17 421.75
R7299 two_stage_opamp_dummy_magic_23_0.Vb2.n9 two_stage_opamp_dummy_magic_23_0.Vb2.t13 421.75
R7300 two_stage_opamp_dummy_magic_23_0.Vb2.n10 two_stage_opamp_dummy_magic_23_0.Vb2.t11 421.75
R7301 two_stage_opamp_dummy_magic_23_0.Vb2.n3 two_stage_opamp_dummy_magic_23_0.Vb2.t21 421.75
R7302 two_stage_opamp_dummy_magic_23_0.Vb2.n4 two_stage_opamp_dummy_magic_23_0.Vb2.t26 421.75
R7303 two_stage_opamp_dummy_magic_23_0.Vb2.n5 two_stage_opamp_dummy_magic_23_0.Vb2.t23 421.75
R7304 two_stage_opamp_dummy_magic_23_0.Vb2.n6 two_stage_opamp_dummy_magic_23_0.Vb2.t28 421.75
R7305 two_stage_opamp_dummy_magic_23_0.Vb2.n21 two_stage_opamp_dummy_magic_23_0.Vb2.n11 313.776
R7306 two_stage_opamp_dummy_magic_23_0.Vb2.n21 two_stage_opamp_dummy_magic_23_0.Vb2.n20 313.212
R7307 two_stage_opamp_dummy_magic_23_0.Vb2.n17 two_stage_opamp_dummy_magic_23_0.Vb2.n16 167.094
R7308 two_stage_opamp_dummy_magic_23_0.Vb2.n18 two_stage_opamp_dummy_magic_23_0.Vb2.n17 167.094
R7309 two_stage_opamp_dummy_magic_23_0.Vb2.n19 two_stage_opamp_dummy_magic_23_0.Vb2.n18 167.094
R7310 two_stage_opamp_dummy_magic_23_0.Vb2.n13 two_stage_opamp_dummy_magic_23_0.Vb2.n12 167.094
R7311 two_stage_opamp_dummy_magic_23_0.Vb2.n14 two_stage_opamp_dummy_magic_23_0.Vb2.n13 167.094
R7312 two_stage_opamp_dummy_magic_23_0.Vb2.n15 two_stage_opamp_dummy_magic_23_0.Vb2.n14 167.094
R7313 two_stage_opamp_dummy_magic_23_0.Vb2.n8 two_stage_opamp_dummy_magic_23_0.Vb2.n7 167.094
R7314 two_stage_opamp_dummy_magic_23_0.Vb2.n9 two_stage_opamp_dummy_magic_23_0.Vb2.n8 167.094
R7315 two_stage_opamp_dummy_magic_23_0.Vb2.n10 two_stage_opamp_dummy_magic_23_0.Vb2.n9 167.094
R7316 two_stage_opamp_dummy_magic_23_0.Vb2.n4 two_stage_opamp_dummy_magic_23_0.Vb2.n3 167.094
R7317 two_stage_opamp_dummy_magic_23_0.Vb2.n5 two_stage_opamp_dummy_magic_23_0.Vb2.n4 167.094
R7318 two_stage_opamp_dummy_magic_23_0.Vb2.n6 two_stage_opamp_dummy_magic_23_0.Vb2.n5 167.094
R7319 two_stage_opamp_dummy_magic_23_0.Vb2.n29 two_stage_opamp_dummy_magic_23_0.Vb2.n28 140.546
R7320 two_stage_opamp_dummy_magic_23_0.Vb2.n27 two_stage_opamp_dummy_magic_23_0.Vb2.n26 139.297
R7321 two_stage_opamp_dummy_magic_23_0.Vb2.n25 two_stage_opamp_dummy_magic_23_0.Vb2.n24 139.297
R7322 two_stage_opamp_dummy_magic_23_0.Vb2.n30 two_stage_opamp_dummy_magic_23_0.Vb2.n29 139.297
R7323 two_stage_opamp_dummy_magic_23_0.Vb2.n25 two_stage_opamp_dummy_magic_23_0.Vb2.n23 67.8536
R7324 two_stage_opamp_dummy_magic_23_0.Vb2.n1 two_stage_opamp_dummy_magic_23_0.Vb2.n0 67.013
R7325 two_stage_opamp_dummy_magic_23_0.Vb2.n20 two_stage_opamp_dummy_magic_23_0.Vb2.n19 35.3472
R7326 two_stage_opamp_dummy_magic_23_0.Vb2.n20 two_stage_opamp_dummy_magic_23_0.Vb2.n15 35.3472
R7327 two_stage_opamp_dummy_magic_23_0.Vb2.n11 two_stage_opamp_dummy_magic_23_0.Vb2.n10 35.3472
R7328 two_stage_opamp_dummy_magic_23_0.Vb2.n11 two_stage_opamp_dummy_magic_23_0.Vb2.n6 35.3472
R7329 two_stage_opamp_dummy_magic_23_0.Vb2.n28 two_stage_opamp_dummy_magic_23_0.Vb2.t2 24.0005
R7330 two_stage_opamp_dummy_magic_23_0.Vb2.n28 two_stage_opamp_dummy_magic_23_0.Vb2.t7 24.0005
R7331 two_stage_opamp_dummy_magic_23_0.Vb2.n26 two_stage_opamp_dummy_magic_23_0.Vb2.t1 24.0005
R7332 two_stage_opamp_dummy_magic_23_0.Vb2.n26 two_stage_opamp_dummy_magic_23_0.Vb2.t5 24.0005
R7333 two_stage_opamp_dummy_magic_23_0.Vb2.n24 two_stage_opamp_dummy_magic_23_0.Vb2.t8 24.0005
R7334 two_stage_opamp_dummy_magic_23_0.Vb2.n24 two_stage_opamp_dummy_magic_23_0.Vb2.t4 24.0005
R7335 two_stage_opamp_dummy_magic_23_0.Vb2.t6 two_stage_opamp_dummy_magic_23_0.Vb2.n30 24.0005
R7336 two_stage_opamp_dummy_magic_23_0.Vb2.n30 two_stage_opamp_dummy_magic_23_0.Vb2.t3 24.0005
R7337 two_stage_opamp_dummy_magic_23_0.Vb2.n22 two_stage_opamp_dummy_magic_23_0.Vb2.n21 13.2817
R7338 two_stage_opamp_dummy_magic_23_0.Vb2.n0 two_stage_opamp_dummy_magic_23_0.Vb2.t10 11.2576
R7339 two_stage_opamp_dummy_magic_23_0.Vb2.n0 two_stage_opamp_dummy_magic_23_0.Vb2.t0 11.2576
R7340 two_stage_opamp_dummy_magic_23_0.Vb2.n2 two_stage_opamp_dummy_magic_23_0.Vb2.n1 7.35988
R7341 two_stage_opamp_dummy_magic_23_0.Vb2.n29 two_stage_opamp_dummy_magic_23_0.Vb2.n27 5.8755
R7342 two_stage_opamp_dummy_magic_23_0.Vb2.n23 two_stage_opamp_dummy_magic_23_0.Vb2.n22 4.55362
R7343 two_stage_opamp_dummy_magic_23_0.Vb2.n27 two_stage_opamp_dummy_magic_23_0.Vb2.n25 1.2505
R7344 two_stage_opamp_dummy_magic_23_0.Vb2.n22 two_stage_opamp_dummy_magic_23_0.Vb2.n2 1.14112
R7345 two_stage_opamp_dummy_magic_23_0.VD3.n26 two_stage_opamp_dummy_magic_23_0.VD3.t32 672.293
R7346 two_stage_opamp_dummy_magic_23_0.VD3.n29 two_stage_opamp_dummy_magic_23_0.VD3.t35 672.293
R7347 two_stage_opamp_dummy_magic_23_0.VD3.t33 two_stage_opamp_dummy_magic_23_0.VD3.n27 213.131
R7348 two_stage_opamp_dummy_magic_23_0.VD3.n28 two_stage_opamp_dummy_magic_23_0.VD3.t36 213.131
R7349 two_stage_opamp_dummy_magic_23_0.VD3.t20 two_stage_opamp_dummy_magic_23_0.VD3.t33 146.155
R7350 two_stage_opamp_dummy_magic_23_0.VD3.t26 two_stage_opamp_dummy_magic_23_0.VD3.t20 146.155
R7351 two_stage_opamp_dummy_magic_23_0.VD3.t22 two_stage_opamp_dummy_magic_23_0.VD3.t26 146.155
R7352 two_stage_opamp_dummy_magic_23_0.VD3.t28 two_stage_opamp_dummy_magic_23_0.VD3.t22 146.155
R7353 two_stage_opamp_dummy_magic_23_0.VD3.t30 two_stage_opamp_dummy_magic_23_0.VD3.t28 146.155
R7354 two_stage_opamp_dummy_magic_23_0.VD3.t12 two_stage_opamp_dummy_magic_23_0.VD3.t30 146.155
R7355 two_stage_opamp_dummy_magic_23_0.VD3.t16 two_stage_opamp_dummy_magic_23_0.VD3.t12 146.155
R7356 two_stage_opamp_dummy_magic_23_0.VD3.t14 two_stage_opamp_dummy_magic_23_0.VD3.t16 146.155
R7357 two_stage_opamp_dummy_magic_23_0.VD3.t18 two_stage_opamp_dummy_magic_23_0.VD3.t14 146.155
R7358 two_stage_opamp_dummy_magic_23_0.VD3.t24 two_stage_opamp_dummy_magic_23_0.VD3.t18 146.155
R7359 two_stage_opamp_dummy_magic_23_0.VD3.t36 two_stage_opamp_dummy_magic_23_0.VD3.t24 146.155
R7360 two_stage_opamp_dummy_magic_23_0.VD3.n27 two_stage_opamp_dummy_magic_23_0.VD3.t34 76.2576
R7361 two_stage_opamp_dummy_magic_23_0.VD3.n28 two_stage_opamp_dummy_magic_23_0.VD3.t37 76.2576
R7362 two_stage_opamp_dummy_magic_23_0.VD3.n1 two_stage_opamp_dummy_magic_23_0.VD3.n0 71.513
R7363 two_stage_opamp_dummy_magic_23_0.VD3.n24 two_stage_opamp_dummy_magic_23_0.VD3.n23 71.513
R7364 two_stage_opamp_dummy_magic_23_0.VD3.n31 two_stage_opamp_dummy_magic_23_0.VD3.n30 71.513
R7365 two_stage_opamp_dummy_magic_23_0.VD3.n33 two_stage_opamp_dummy_magic_23_0.VD3.n32 71.513
R7366 two_stage_opamp_dummy_magic_23_0.VD3.n35 two_stage_opamp_dummy_magic_23_0.VD3.n34 71.513
R7367 two_stage_opamp_dummy_magic_23_0.VD3.n5 two_stage_opamp_dummy_magic_23_0.VD3.n4 66.0338
R7368 two_stage_opamp_dummy_magic_23_0.VD3.n8 two_stage_opamp_dummy_magic_23_0.VD3.n7 66.0338
R7369 two_stage_opamp_dummy_magic_23_0.VD3.n11 two_stage_opamp_dummy_magic_23_0.VD3.n10 66.0338
R7370 two_stage_opamp_dummy_magic_23_0.VD3.n15 two_stage_opamp_dummy_magic_23_0.VD3.n14 66.0338
R7371 two_stage_opamp_dummy_magic_23_0.VD3.n18 two_stage_opamp_dummy_magic_23_0.VD3.n17 66.0338
R7372 two_stage_opamp_dummy_magic_23_0.VD3.n21 two_stage_opamp_dummy_magic_23_0.VD3.n20 66.0338
R7373 two_stage_opamp_dummy_magic_23_0.VD3.n25 two_stage_opamp_dummy_magic_23_0.VD3.n22 14.0005
R7374 two_stage_opamp_dummy_magic_23_0.VD3.n0 two_stage_opamp_dummy_magic_23_0.VD3.t23 11.2576
R7375 two_stage_opamp_dummy_magic_23_0.VD3.n0 two_stage_opamp_dummy_magic_23_0.VD3.t29 11.2576
R7376 two_stage_opamp_dummy_magic_23_0.VD3.n23 two_stage_opamp_dummy_magic_23_0.VD3.t21 11.2576
R7377 two_stage_opamp_dummy_magic_23_0.VD3.n23 two_stage_opamp_dummy_magic_23_0.VD3.t27 11.2576
R7378 two_stage_opamp_dummy_magic_23_0.VD3.n30 two_stage_opamp_dummy_magic_23_0.VD3.t19 11.2576
R7379 two_stage_opamp_dummy_magic_23_0.VD3.n30 two_stage_opamp_dummy_magic_23_0.VD3.t25 11.2576
R7380 two_stage_opamp_dummy_magic_23_0.VD3.n32 two_stage_opamp_dummy_magic_23_0.VD3.t17 11.2576
R7381 two_stage_opamp_dummy_magic_23_0.VD3.n32 two_stage_opamp_dummy_magic_23_0.VD3.t15 11.2576
R7382 two_stage_opamp_dummy_magic_23_0.VD3.n4 two_stage_opamp_dummy_magic_23_0.VD3.t10 11.2576
R7383 two_stage_opamp_dummy_magic_23_0.VD3.n4 two_stage_opamp_dummy_magic_23_0.VD3.t3 11.2576
R7384 two_stage_opamp_dummy_magic_23_0.VD3.n7 two_stage_opamp_dummy_magic_23_0.VD3.t1 11.2576
R7385 two_stage_opamp_dummy_magic_23_0.VD3.n7 two_stage_opamp_dummy_magic_23_0.VD3.t4 11.2576
R7386 two_stage_opamp_dummy_magic_23_0.VD3.n10 two_stage_opamp_dummy_magic_23_0.VD3.t6 11.2576
R7387 two_stage_opamp_dummy_magic_23_0.VD3.n10 two_stage_opamp_dummy_magic_23_0.VD3.t8 11.2576
R7388 two_stage_opamp_dummy_magic_23_0.VD3.n14 two_stage_opamp_dummy_magic_23_0.VD3.t9 11.2576
R7389 two_stage_opamp_dummy_magic_23_0.VD3.n14 two_stage_opamp_dummy_magic_23_0.VD3.t0 11.2576
R7390 two_stage_opamp_dummy_magic_23_0.VD3.n17 two_stage_opamp_dummy_magic_23_0.VD3.t2 11.2576
R7391 two_stage_opamp_dummy_magic_23_0.VD3.n17 two_stage_opamp_dummy_magic_23_0.VD3.t5 11.2576
R7392 two_stage_opamp_dummy_magic_23_0.VD3.n20 two_stage_opamp_dummy_magic_23_0.VD3.t7 11.2576
R7393 two_stage_opamp_dummy_magic_23_0.VD3.n20 two_stage_opamp_dummy_magic_23_0.VD3.t11 11.2576
R7394 two_stage_opamp_dummy_magic_23_0.VD3.t31 two_stage_opamp_dummy_magic_23_0.VD3.n35 11.2576
R7395 two_stage_opamp_dummy_magic_23_0.VD3.n35 two_stage_opamp_dummy_magic_23_0.VD3.t13 11.2576
R7396 two_stage_opamp_dummy_magic_23_0.VD3.n31 two_stage_opamp_dummy_magic_23_0.VD3.n29 6.10467
R7397 two_stage_opamp_dummy_magic_23_0.VD3.n21 two_stage_opamp_dummy_magic_23_0.VD3.n19 5.91717
R7398 two_stage_opamp_dummy_magic_23_0.VD3.n6 two_stage_opamp_dummy_magic_23_0.VD3.n5 5.91717
R7399 two_stage_opamp_dummy_magic_23_0.VD3.n9 two_stage_opamp_dummy_magic_23_0.VD3.n5 5.91717
R7400 two_stage_opamp_dummy_magic_23_0.VD3.n26 two_stage_opamp_dummy_magic_23_0.VD3.n25 5.47967
R7401 two_stage_opamp_dummy_magic_23_0.VD3.n9 two_stage_opamp_dummy_magic_23_0.VD3.n8 5.29217
R7402 two_stage_opamp_dummy_magic_23_0.VD3.n8 two_stage_opamp_dummy_magic_23_0.VD3.n6 5.29217
R7403 two_stage_opamp_dummy_magic_23_0.VD3.n12 two_stage_opamp_dummy_magic_23_0.VD3.n11 5.29217
R7404 two_stage_opamp_dummy_magic_23_0.VD3.n11 two_stage_opamp_dummy_magic_23_0.VD3.n3 5.29217
R7405 two_stage_opamp_dummy_magic_23_0.VD3.n15 two_stage_opamp_dummy_magic_23_0.VD3.n13 5.29217
R7406 two_stage_opamp_dummy_magic_23_0.VD3.n16 two_stage_opamp_dummy_magic_23_0.VD3.n15 5.29217
R7407 two_stage_opamp_dummy_magic_23_0.VD3.n18 two_stage_opamp_dummy_magic_23_0.VD3.n2 5.29217
R7408 two_stage_opamp_dummy_magic_23_0.VD3.n19 two_stage_opamp_dummy_magic_23_0.VD3.n18 5.29217
R7409 two_stage_opamp_dummy_magic_23_0.VD3.n22 two_stage_opamp_dummy_magic_23_0.VD3.n21 5.29217
R7410 two_stage_opamp_dummy_magic_23_0.VD3.n29 two_stage_opamp_dummy_magic_23_0.VD3.n28 1.03383
R7411 two_stage_opamp_dummy_magic_23_0.VD3.n27 two_stage_opamp_dummy_magic_23_0.VD3.n26 1.03383
R7412 two_stage_opamp_dummy_magic_23_0.VD3.n34 two_stage_opamp_dummy_magic_23_0.VD3.n33 0.6255
R7413 two_stage_opamp_dummy_magic_23_0.VD3.n33 two_stage_opamp_dummy_magic_23_0.VD3.n31 0.6255
R7414 two_stage_opamp_dummy_magic_23_0.VD3.n19 two_stage_opamp_dummy_magic_23_0.VD3.n16 0.6255
R7415 two_stage_opamp_dummy_magic_23_0.VD3.n16 two_stage_opamp_dummy_magic_23_0.VD3.n3 0.6255
R7416 two_stage_opamp_dummy_magic_23_0.VD3.n6 two_stage_opamp_dummy_magic_23_0.VD3.n3 0.6255
R7417 two_stage_opamp_dummy_magic_23_0.VD3.n12 two_stage_opamp_dummy_magic_23_0.VD3.n9 0.6255
R7418 two_stage_opamp_dummy_magic_23_0.VD3.n13 two_stage_opamp_dummy_magic_23_0.VD3.n12 0.6255
R7419 two_stage_opamp_dummy_magic_23_0.VD3.n13 two_stage_opamp_dummy_magic_23_0.VD3.n2 0.6255
R7420 two_stage_opamp_dummy_magic_23_0.VD3.n22 two_stage_opamp_dummy_magic_23_0.VD3.n2 0.6255
R7421 two_stage_opamp_dummy_magic_23_0.VD3.n25 two_stage_opamp_dummy_magic_23_0.VD3.n24 0.6255
R7422 two_stage_opamp_dummy_magic_23_0.VD3.n24 two_stage_opamp_dummy_magic_23_0.VD3.n1 0.6255
R7423 two_stage_opamp_dummy_magic_23_0.VD3.n34 two_stage_opamp_dummy_magic_23_0.VD3.n1 0.6255
R7424 a_5820_23644.t0 a_5820_23644.t1 178.133
R7425 two_stage_opamp_dummy_magic_23_0.cap_res_Y two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 49.2388
R7426 two_stage_opamp_dummy_magic_23_0.cap_res_Y two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 0.922875
R7427 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 0.1603
R7428 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t90 0.1603
R7429 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t94 0.1603
R7430 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 0.1603
R7431 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 0.1603
R7432 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 0.1603
R7433 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t27 0.1603
R7434 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t52 0.1603
R7435 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 0.1603
R7436 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t21 0.1603
R7437 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 0.1603
R7438 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t59 0.1603
R7439 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 0.1603
R7440 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t99 0.1603
R7441 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 0.1603
R7442 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t67 0.1603
R7443 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t76 0.1603
R7444 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t104 0.1603
R7445 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 0.1603
R7446 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 0.1603
R7447 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t82 0.1603
R7448 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t109 0.1603
R7449 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 0.1603
R7450 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 0.1603
R7451 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t20 0.1603
R7452 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t47 0.1603
R7453 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t58 0.1603
R7454 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 0.1603
R7455 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 0.1603
R7456 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t53 0.1603
R7457 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t98 0.1603
R7458 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 0.1603
R7459 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 0.1603
R7460 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 0.1603
R7461 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 0.1603
R7462 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 0.1603
R7463 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t31 0.1603
R7464 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 0.1603
R7465 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t113 0.1603
R7466 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 0.1603
R7467 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t57 0.1603
R7468 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 0.1603
R7469 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 0.1603
R7470 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 0.1603
R7471 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 0.1603
R7472 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t65 0.1603
R7473 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t100 0.1603
R7474 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t80 0.1603
R7475 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 0.1603
R7476 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 0.1603
R7477 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 0.1603
R7478 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 0.1603
R7479 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t75 0.1603
R7480 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 0.1603
R7481 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 0.1603
R7482 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 0.1603
R7483 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 0.1603
R7484 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 0.1603
R7485 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 0.159278
R7486 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 0.159278
R7487 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 0.159278
R7488 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 0.159278
R7489 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 0.159278
R7490 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 0.159278
R7491 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 0.159278
R7492 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 0.159278
R7493 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 0.159278
R7494 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 0.159278
R7495 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 0.159278
R7496 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 0.159278
R7497 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 0.159278
R7498 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 0.159278
R7499 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 0.159278
R7500 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 0.159278
R7501 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 0.159278
R7502 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t81 0.159278
R7503 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 0.159278
R7504 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t66 0.159278
R7505 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 0.159278
R7506 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t95 0.159278
R7507 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 0.159278
R7508 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 0.159278
R7509 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t8 0.159278
R7510 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 0.159278
R7511 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 0.159278
R7512 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 0.137822
R7513 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 0.1368
R7514 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 0.1368
R7515 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 0.1368
R7516 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 0.1368
R7517 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 0.1368
R7518 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 0.1368
R7519 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 0.1368
R7520 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 0.1368
R7521 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 0.1368
R7522 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 0.1368
R7523 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 0.1368
R7524 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 0.1368
R7525 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 0.1368
R7526 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 0.1368
R7527 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 0.1368
R7528 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 0.1368
R7529 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 0.1368
R7530 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 0.1368
R7531 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 0.1368
R7532 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 0.1368
R7533 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 0.1368
R7534 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 0.1368
R7535 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 0.1368
R7536 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 0.1368
R7537 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 0.1368
R7538 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 0.1368
R7539 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 0.1368
R7540 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 0.1368
R7541 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 0.1368
R7542 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 0.1368
R7543 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 0.1368
R7544 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 0.114322
R7545 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 0.1133
R7546 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 0.1133
R7547 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 0.1133
R7548 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 0.1133
R7549 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 0.1133
R7550 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 0.1133
R7551 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 0.1133
R7552 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 0.1133
R7553 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 0.1133
R7554 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 0.1133
R7555 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 0.1133
R7556 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 0.1133
R7557 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 0.1133
R7558 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 0.1133
R7559 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 0.1133
R7560 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 0.1133
R7561 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 0.1133
R7562 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 0.1133
R7563 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 0.1133
R7564 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 0.00152174
R7565 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 0.00152174
R7566 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 0.00152174
R7567 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 0.00152174
R7568 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 0.00152174
R7569 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 0.00152174
R7570 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 0.00152174
R7571 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 0.00152174
R7572 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 0.00152174
R7573 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 0.00152174
R7574 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 0.00152174
R7575 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 0.00152174
R7576 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 0.00152174
R7577 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 0.00152174
R7578 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 0.00152174
R7579 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 0.00152174
R7580 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 0.00152174
R7581 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 0.00152174
R7582 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 0.00152174
R7583 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 0.00152174
R7584 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 0.00152174
R7585 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 0.00152174
R7586 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 0.00152174
R7587 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 0.00152174
R7588 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 0.00152174
R7589 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 0.00152174
R7590 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 0.00152174
R7591 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 0.00152174
R7592 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 0.00152174
R7593 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 0.00152174
R7594 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 0.00152174
R7595 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 0.00152174
R7596 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 0.00152174
R7597 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 0.00152174
R7598 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 0.00152174
R7599 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 0.00152174
R7600 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 325.473
R7601 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 325.473
R7602 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 325.473
R7603 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t18 310.488
R7604 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t16 310.488
R7605 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t17 310.488
R7606 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t8 184.097
R7607 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t10 184.097
R7608 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t2 184.097
R7609 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.n11 167.094
R7610 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R7611 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R7612 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n13 152
R7613 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 152
R7614 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 152
R7615 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t14 120.501
R7616 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t6 120.501
R7617 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t15 120.501
R7618 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t4 120.501
R7619 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t13 120.501
R7620 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t0 120.501
R7621 bgr_11_0.V_mir1.t12 bgr_11_0.V_mir1.n16 106.931
R7622 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 40.7027
R7623 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R7624 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R7625 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.t9 39.4005
R7626 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.t7 39.4005
R7627 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t11 39.4005
R7628 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t5 39.4005
R7629 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t3 39.4005
R7630 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t1 39.4005
R7631 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 15.9255
R7632 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n4 15.9255
R7633 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.n15 9.3005
R7634 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.n10 4.5005
R7635 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t10 354.854
R7636 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t23 346.8
R7637 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n11 339.522
R7638 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n6 339.522
R7639 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 335.022
R7640 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t25 184.097
R7641 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t9 184.097
R7642 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t19 184.097
R7643 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t12 184.097
R7644 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n10 166.05
R7645 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n7 166.05
R7646 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t6 106.556
R7647 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.n0 54.5884
R7648 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t2 39.4005
R7649 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t1 39.4005
R7650 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t4 39.4005
R7651 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t0 39.4005
R7652 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t5 39.4005
R7653 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t3 39.4005
R7654 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t7 4.8295
R7655 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t24 4.8295
R7656 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t28 4.8295
R7657 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t15 4.8295
R7658 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t32 4.8295
R7659 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t21 4.8295
R7660 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t26 4.8295
R7661 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t14 4.8295
R7662 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t16 4.8295
R7663 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t29 4.5005
R7664 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t31 4.5005
R7665 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R7666 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t22 4.5005
R7667 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t27 4.5005
R7668 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t30 4.5005
R7669 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t17 4.5005
R7670 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t20 4.5005
R7671 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t11 4.5005
R7672 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t13 4.5005
R7673 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t8 4.5005
R7674 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n9 4.5005
R7675 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n2 2.2095
R7676 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n4 2.0005
R7677 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n3 1.813
R7678 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n5 1.813
R7679 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.8935
R7680 w_6100_17280.n27 w_6100_17280.t44 708.125
R7681 w_6100_17280.t44 w_6100_17280.n12 708.125
R7682 w_6100_17280.n35 w_6100_17280.t47 708.125
R7683 w_6100_17280.t47 w_6100_17280.n29 708.125
R7684 w_6100_17280.n37 w_6100_17280.t40 660.001
R7685 w_6100_17280.n26 w_6100_17280.t43 657.76
R7686 w_6100_17280.t46 w_6100_17280.n36 657.76
R7687 w_6100_17280.t37 w_6100_17280.n25 540.818
R7688 w_6100_17280.t43 w_6100_17280.t76 407.144
R7689 w_6100_17280.t76 w_6100_17280.t0 407.144
R7690 w_6100_17280.t0 w_6100_17280.t32 407.144
R7691 w_6100_17280.t32 w_6100_17280.t78 407.144
R7692 w_6100_17280.t78 w_6100_17280.t30 407.144
R7693 w_6100_17280.t30 w_6100_17280.t68 407.144
R7694 w_6100_17280.t68 w_6100_17280.t72 407.144
R7695 w_6100_17280.t72 w_6100_17280.t82 407.144
R7696 w_6100_17280.t82 w_6100_17280.t64 407.144
R7697 w_6100_17280.t64 w_6100_17280.t2 407.144
R7698 w_6100_17280.t2 w_6100_17280.t28 407.144
R7699 w_6100_17280.t28 w_6100_17280.t66 407.144
R7700 w_6100_17280.t66 w_6100_17280.t70 407.144
R7701 w_6100_17280.t70 w_6100_17280.t48 407.144
R7702 w_6100_17280.t48 w_6100_17280.t80 407.144
R7703 w_6100_17280.t80 w_6100_17280.t34 407.144
R7704 w_6100_17280.t34 w_6100_17280.t62 407.144
R7705 w_6100_17280.t62 w_6100_17280.t74 407.144
R7706 w_6100_17280.t74 w_6100_17280.t37 407.144
R7707 w_6100_17280.t52 w_6100_17280.t46 407.144
R7708 w_6100_17280.t4 w_6100_17280.t52 407.144
R7709 w_6100_17280.t16 w_6100_17280.t4 407.144
R7710 w_6100_17280.t26 w_6100_17280.t16 407.144
R7711 w_6100_17280.t12 w_6100_17280.t26 407.144
R7712 w_6100_17280.t56 w_6100_17280.t12 407.144
R7713 w_6100_17280.t54 w_6100_17280.t56 407.144
R7714 w_6100_17280.t24 w_6100_17280.t54 407.144
R7715 w_6100_17280.t10 w_6100_17280.t24 407.144
R7716 w_6100_17280.t20 w_6100_17280.t10 407.144
R7717 w_6100_17280.t6 w_6100_17280.t20 407.144
R7718 w_6100_17280.t60 w_6100_17280.t6 407.144
R7719 w_6100_17280.t50 w_6100_17280.t60 407.144
R7720 w_6100_17280.t22 w_6100_17280.t50 407.144
R7721 w_6100_17280.t8 w_6100_17280.t22 407.144
R7722 w_6100_17280.t18 w_6100_17280.t8 407.144
R7723 w_6100_17280.t14 w_6100_17280.t18 407.144
R7724 w_6100_17280.t58 w_6100_17280.t14 407.144
R7725 w_6100_17280.t40 w_6100_17280.t58 407.144
R7726 w_6100_17280.t42 w_6100_17280.n27 379.582
R7727 w_6100_17280.n35 w_6100_17280.t45 379.582
R7728 w_6100_17280.n24 w_6100_17280.t36 379.277
R7729 w_6100_17280.t36 w_6100_17280.n22 358.858
R7730 w_6100_17280.n28 w_6100_17280.t42 358.858
R7731 w_6100_17280.n38 w_6100_17280.t39 358.858
R7732 w_6100_17280.t45 w_6100_17280.n34 358.858
R7733 w_6100_17280.n37 w_6100_17280.t41 354.065
R7734 w_6100_17280.n23 w_6100_17280.t38 351.793
R7735 w_6100_17280.n9 w_6100_17280.n21 339.214
R7736 w_6100_17280.n9 w_6100_17280.n20 339.214
R7737 w_6100_17280.n8 w_6100_17280.n19 339.214
R7738 w_6100_17280.n8 w_6100_17280.n18 339.214
R7739 w_6100_17280.n7 w_6100_17280.n17 339.214
R7740 w_6100_17280.n7 w_6100_17280.n16 339.214
R7741 w_6100_17280.n6 w_6100_17280.n15 339.214
R7742 w_6100_17280.n6 w_6100_17280.n14 339.214
R7743 w_6100_17280.n5 w_6100_17280.n11 339.214
R7744 w_6100_17280.n4 w_6100_17280.n39 339.214
R7745 w_6100_17280.n3 w_6100_17280.n40 339.214
R7746 w_6100_17280.n3 w_6100_17280.n41 339.214
R7747 w_6100_17280.n2 w_6100_17280.n10 339.214
R7748 w_6100_17280.n0 w_6100_17280.n30 339.214
R7749 w_6100_17280.n0 w_6100_17280.n31 339.214
R7750 w_6100_17280.n1 w_6100_17280.n32 339.214
R7751 w_6100_17280.n1 w_6100_17280.n33 339.214
R7752 w_6100_17280.n42 w_6100_17280.n2 339.214
R7753 w_6100_17280.n25 w_6100_17280.n24 238.367
R7754 w_6100_17280.n25 w_6100_17280.n13 238.367
R7755 w_6100_17280.n21 w_6100_17280.t63 39.4005
R7756 w_6100_17280.n21 w_6100_17280.t75 39.4005
R7757 w_6100_17280.n20 w_6100_17280.t81 39.4005
R7758 w_6100_17280.n20 w_6100_17280.t35 39.4005
R7759 w_6100_17280.n19 w_6100_17280.t71 39.4005
R7760 w_6100_17280.n19 w_6100_17280.t49 39.4005
R7761 w_6100_17280.n18 w_6100_17280.t29 39.4005
R7762 w_6100_17280.n18 w_6100_17280.t67 39.4005
R7763 w_6100_17280.n17 w_6100_17280.t65 39.4005
R7764 w_6100_17280.n17 w_6100_17280.t3 39.4005
R7765 w_6100_17280.n16 w_6100_17280.t73 39.4005
R7766 w_6100_17280.n16 w_6100_17280.t83 39.4005
R7767 w_6100_17280.n15 w_6100_17280.t31 39.4005
R7768 w_6100_17280.n15 w_6100_17280.t69 39.4005
R7769 w_6100_17280.n14 w_6100_17280.t33 39.4005
R7770 w_6100_17280.n14 w_6100_17280.t79 39.4005
R7771 w_6100_17280.n11 w_6100_17280.t77 39.4005
R7772 w_6100_17280.n11 w_6100_17280.t1 39.4005
R7773 w_6100_17280.n39 w_6100_17280.t15 39.4005
R7774 w_6100_17280.n39 w_6100_17280.t59 39.4005
R7775 w_6100_17280.n40 w_6100_17280.t9 39.4005
R7776 w_6100_17280.n40 w_6100_17280.t19 39.4005
R7777 w_6100_17280.n41 w_6100_17280.t51 39.4005
R7778 w_6100_17280.n41 w_6100_17280.t23 39.4005
R7779 w_6100_17280.n10 w_6100_17280.t11 39.4005
R7780 w_6100_17280.n10 w_6100_17280.t21 39.4005
R7781 w_6100_17280.n30 w_6100_17280.t55 39.4005
R7782 w_6100_17280.n30 w_6100_17280.t25 39.4005
R7783 w_6100_17280.n31 w_6100_17280.t13 39.4005
R7784 w_6100_17280.n31 w_6100_17280.t57 39.4005
R7785 w_6100_17280.n32 w_6100_17280.t17 39.4005
R7786 w_6100_17280.n32 w_6100_17280.t27 39.4005
R7787 w_6100_17280.n33 w_6100_17280.t53 39.4005
R7788 w_6100_17280.n33 w_6100_17280.t5 39.4005
R7789 w_6100_17280.n42 w_6100_17280.t7 39.4005
R7790 w_6100_17280.t61 w_6100_17280.n42 39.4005
R7791 w_6100_17280.n38 w_6100_17280.n37 22.9536
R7792 w_6100_17280.n22 w_6100_17280.n13 20.7243
R7793 w_6100_17280.n28 w_6100_17280.n12 20.7243
R7794 w_6100_17280.n34 w_6100_17280.n29 20.7243
R7795 w_6100_17280.n34 w_6100_17280.n1 11.7346
R7796 w_6100_17280.n22 w_6100_17280.n9 11.7346
R7797 w_6100_17280.n5 w_6100_17280.n28 11.6096
R7798 w_6100_17280.n4 w_6100_17280.n38 11.6096
R7799 w_6100_17280.n23 w_6100_17280.n13 4.54311
R7800 w_6100_17280.n24 w_6100_17280.n23 4.54311
R7801 w_6100_17280.n26 w_6100_17280.n12 4.48641
R7802 w_6100_17280.n27 w_6100_17280.n26 4.48641
R7803 w_6100_17280.n36 w_6100_17280.n29 4.48641
R7804 w_6100_17280.n36 w_6100_17280.n35 4.48641
R7805 w_6100_17280.n6 w_6100_17280.n5 0.3755
R7806 w_6100_17280.n1 w_6100_17280.n0 0.3755
R7807 w_6100_17280.n4 w_6100_17280.n5 0.333833
R7808 w_6100_17280.n9 w_6100_17280.n8 0.2505
R7809 w_6100_17280.n8 w_6100_17280.n7 0.2505
R7810 w_6100_17280.n7 w_6100_17280.n6 0.2505
R7811 w_6100_17280.n3 w_6100_17280.n4 0.2505
R7812 w_6100_17280.n2 w_6100_17280.n3 0.2505
R7813 w_6100_17280.n0 w_6100_17280.n2 0.2505
R7814 bgr_11_0.cap_res1.t0 bgr_11_0.cap_res1.t18 121.245
R7815 bgr_11_0.cap_res1.t17 bgr_11_0.cap_res1.t19 0.1603
R7816 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.t16 0.1603
R7817 bgr_11_0.cap_res1.t3 bgr_11_0.cap_res1.t10 0.1603
R7818 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t15 0.1603
R7819 bgr_11_0.cap_res1.t2 bgr_11_0.cap_res1.t8 0.1603
R7820 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t4 0.159278
R7821 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t12 0.159278
R7822 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t6 0.159278
R7823 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t13 0.159278
R7824 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t17 0.1368
R7825 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t14 0.1368
R7826 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t11 0.1368
R7827 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t7 0.1368
R7828 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t3 0.1368
R7829 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t1 0.1368
R7830 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t9 0.1368
R7831 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t5 0.1368
R7832 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t2 0.1368
R7833 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t20 0.1368
R7834 bgr_11_0.cap_res1.t4 bgr_11_0.cap_res1.n0 0.00152174
R7835 bgr_11_0.cap_res1.t12 bgr_11_0.cap_res1.n1 0.00152174
R7836 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.n2 0.00152174
R7837 bgr_11_0.cap_res1.t13 bgr_11_0.cap_res1.n3 0.00152174
R7838 bgr_11_0.cap_res1.t18 bgr_11_0.cap_res1.n4 0.00152174
R7839 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t3 536.909
R7840 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 371.678
R7841 bgr_11_0.V_CUR_REF_REG.t0 bgr_11_0.V_CUR_REF_REG.n1 153.099
R7842 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t1 39.4005
R7843 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R7844 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t0 201.28
R7845 bgr_11_0.V_p_2.t1 bgr_11_0.V_p_2.n0 9.6005
R7846 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 9.6005
R7847 two_stage_opamp_dummy_magic_23_0.VD2.n6 two_stage_opamp_dummy_magic_23_0.VD2.n5 49.3505
R7848 two_stage_opamp_dummy_magic_23_0.VD2.n4 two_stage_opamp_dummy_magic_23_0.VD2.n3 49.3505
R7849 two_stage_opamp_dummy_magic_23_0.VD2.n13 two_stage_opamp_dummy_magic_23_0.VD2.n12 49.3505
R7850 two_stage_opamp_dummy_magic_23_0.VD2.n1 two_stage_opamp_dummy_magic_23_0.VD2.n0 49.3505
R7851 two_stage_opamp_dummy_magic_23_0.VD2.n20 two_stage_opamp_dummy_magic_23_0.VD2.n19 49.3505
R7852 two_stage_opamp_dummy_magic_23_0.VD2.n23 two_stage_opamp_dummy_magic_23_0.VD2.n22 49.3505
R7853 two_stage_opamp_dummy_magic_23_0.VD2.n26 two_stage_opamp_dummy_magic_23_0.VD2.n25 49.3505
R7854 two_stage_opamp_dummy_magic_23_0.VD2.n29 two_stage_opamp_dummy_magic_23_0.VD2.n28 49.3505
R7855 two_stage_opamp_dummy_magic_23_0.VD2.n31 two_stage_opamp_dummy_magic_23_0.VD2.n30 49.3505
R7856 two_stage_opamp_dummy_magic_23_0.VD2.n35 two_stage_opamp_dummy_magic_23_0.VD2.n34 49.3505
R7857 two_stage_opamp_dummy_magic_23_0.VD2.n8 two_stage_opamp_dummy_magic_23_0.VD2.n7 49.3505
R7858 two_stage_opamp_dummy_magic_23_0.VD2.n5 two_stage_opamp_dummy_magic_23_0.VD2.t9 16.0005
R7859 two_stage_opamp_dummy_magic_23_0.VD2.n5 two_stage_opamp_dummy_magic_23_0.VD2.t4 16.0005
R7860 two_stage_opamp_dummy_magic_23_0.VD2.n3 two_stage_opamp_dummy_magic_23_0.VD2.t5 16.0005
R7861 two_stage_opamp_dummy_magic_23_0.VD2.n3 two_stage_opamp_dummy_magic_23_0.VD2.t1 16.0005
R7862 two_stage_opamp_dummy_magic_23_0.VD2.n12 two_stage_opamp_dummy_magic_23_0.VD2.t6 16.0005
R7863 two_stage_opamp_dummy_magic_23_0.VD2.n12 two_stage_opamp_dummy_magic_23_0.VD2.t2 16.0005
R7864 two_stage_opamp_dummy_magic_23_0.VD2.n0 two_stage_opamp_dummy_magic_23_0.VD2.t8 16.0005
R7865 two_stage_opamp_dummy_magic_23_0.VD2.n0 two_stage_opamp_dummy_magic_23_0.VD2.t3 16.0005
R7866 two_stage_opamp_dummy_magic_23_0.VD2.n19 two_stage_opamp_dummy_magic_23_0.VD2.t19 16.0005
R7867 two_stage_opamp_dummy_magic_23_0.VD2.n19 two_stage_opamp_dummy_magic_23_0.VD2.t21 16.0005
R7868 two_stage_opamp_dummy_magic_23_0.VD2.n22 two_stage_opamp_dummy_magic_23_0.VD2.t11 16.0005
R7869 two_stage_opamp_dummy_magic_23_0.VD2.n22 two_stage_opamp_dummy_magic_23_0.VD2.t18 16.0005
R7870 two_stage_opamp_dummy_magic_23_0.VD2.n25 two_stage_opamp_dummy_magic_23_0.VD2.t15 16.0005
R7871 two_stage_opamp_dummy_magic_23_0.VD2.n25 two_stage_opamp_dummy_magic_23_0.VD2.t14 16.0005
R7872 two_stage_opamp_dummy_magic_23_0.VD2.n28 two_stage_opamp_dummy_magic_23_0.VD2.t16 16.0005
R7873 two_stage_opamp_dummy_magic_23_0.VD2.n28 two_stage_opamp_dummy_magic_23_0.VD2.t20 16.0005
R7874 two_stage_opamp_dummy_magic_23_0.VD2.n30 two_stage_opamp_dummy_magic_23_0.VD2.t12 16.0005
R7875 two_stage_opamp_dummy_magic_23_0.VD2.n30 two_stage_opamp_dummy_magic_23_0.VD2.t0 16.0005
R7876 two_stage_opamp_dummy_magic_23_0.VD2.n34 two_stage_opamp_dummy_magic_23_0.VD2.t17 16.0005
R7877 two_stage_opamp_dummy_magic_23_0.VD2.n34 two_stage_opamp_dummy_magic_23_0.VD2.t13 16.0005
R7878 two_stage_opamp_dummy_magic_23_0.VD2.n7 two_stage_opamp_dummy_magic_23_0.VD2.t7 16.0005
R7879 two_stage_opamp_dummy_magic_23_0.VD2.n7 two_stage_opamp_dummy_magic_23_0.VD2.t10 16.0005
R7880 two_stage_opamp_dummy_magic_23_0.VD2.n29 two_stage_opamp_dummy_magic_23_0.VD2.n18 5.64633
R7881 two_stage_opamp_dummy_magic_23_0.VD2.n21 two_stage_opamp_dummy_magic_23_0.VD2.n20 5.64633
R7882 two_stage_opamp_dummy_magic_23_0.VD2.n11 two_stage_opamp_dummy_magic_23_0.VD2.n4 5.6255
R7883 two_stage_opamp_dummy_magic_23_0.VD2.n9 two_stage_opamp_dummy_magic_23_0.VD2.n6 5.6255
R7884 two_stage_opamp_dummy_magic_23_0.VD2.n32 two_stage_opamp_dummy_magic_23_0.VD2.n29 5.438
R7885 two_stage_opamp_dummy_magic_23_0.VD2.n24 two_stage_opamp_dummy_magic_23_0.VD2.n20 5.438
R7886 two_stage_opamp_dummy_magic_23_0.VD2.n14 two_stage_opamp_dummy_magic_23_0.VD2.n4 5.438
R7887 two_stage_opamp_dummy_magic_23_0.VD2.n6 two_stage_opamp_dummy_magic_23_0.VD2.n2 5.438
R7888 two_stage_opamp_dummy_magic_23_0.VD2.n23 two_stage_opamp_dummy_magic_23_0.VD2.n21 5.08383
R7889 two_stage_opamp_dummy_magic_23_0.VD2.n26 two_stage_opamp_dummy_magic_23_0.VD2.n17 5.08383
R7890 two_stage_opamp_dummy_magic_23_0.VD2.n31 two_stage_opamp_dummy_magic_23_0.VD2.n18 5.08383
R7891 two_stage_opamp_dummy_magic_23_0.VD2.n36 two_stage_opamp_dummy_magic_23_0.VD2.n35 5.08383
R7892 two_stage_opamp_dummy_magic_23_0.VD2.n9 two_stage_opamp_dummy_magic_23_0.VD2.n8 5.063
R7893 two_stage_opamp_dummy_magic_23_0.VD2.n13 two_stage_opamp_dummy_magic_23_0.VD2.n11 5.063
R7894 two_stage_opamp_dummy_magic_23_0.VD2.n10 two_stage_opamp_dummy_magic_23_0.VD2.n1 5.063
R7895 two_stage_opamp_dummy_magic_23_0.VD2 two_stage_opamp_dummy_magic_23_0.VD2.n37 5.02133
R7896 two_stage_opamp_dummy_magic_23_0.VD2.n14 two_stage_opamp_dummy_magic_23_0.VD2.n13 4.8755
R7897 two_stage_opamp_dummy_magic_23_0.VD2.n24 two_stage_opamp_dummy_magic_23_0.VD2.n23 4.8755
R7898 two_stage_opamp_dummy_magic_23_0.VD2.n27 two_stage_opamp_dummy_magic_23_0.VD2.n26 4.8755
R7899 two_stage_opamp_dummy_magic_23_0.VD2.n32 two_stage_opamp_dummy_magic_23_0.VD2.n31 4.8755
R7900 two_stage_opamp_dummy_magic_23_0.VD2.n35 two_stage_opamp_dummy_magic_23_0.VD2.n33 4.8755
R7901 two_stage_opamp_dummy_magic_23_0.VD2.n8 two_stage_opamp_dummy_magic_23_0.VD2.n2 4.8755
R7902 two_stage_opamp_dummy_magic_23_0.VD2.n16 two_stage_opamp_dummy_magic_23_0.VD2.n15 4.5005
R7903 two_stage_opamp_dummy_magic_23_0.VD2 two_stage_opamp_dummy_magic_23_0.VD2.n16 0.7505
R7904 two_stage_opamp_dummy_magic_23_0.VD2.n36 two_stage_opamp_dummy_magic_23_0.VD2.n18 0.563
R7905 two_stage_opamp_dummy_magic_23_0.VD2.n33 two_stage_opamp_dummy_magic_23_0.VD2.n32 0.563
R7906 two_stage_opamp_dummy_magic_23_0.VD2.n33 two_stage_opamp_dummy_magic_23_0.VD2.n27 0.563
R7907 two_stage_opamp_dummy_magic_23_0.VD2.n27 two_stage_opamp_dummy_magic_23_0.VD2.n24 0.563
R7908 two_stage_opamp_dummy_magic_23_0.VD2.n21 two_stage_opamp_dummy_magic_23_0.VD2.n17 0.563
R7909 two_stage_opamp_dummy_magic_23_0.VD2.n15 two_stage_opamp_dummy_magic_23_0.VD2.n2 0.563
R7910 two_stage_opamp_dummy_magic_23_0.VD2.n15 two_stage_opamp_dummy_magic_23_0.VD2.n14 0.563
R7911 two_stage_opamp_dummy_magic_23_0.VD2.n11 two_stage_opamp_dummy_magic_23_0.VD2.n10 0.563
R7912 two_stage_opamp_dummy_magic_23_0.VD2.n10 two_stage_opamp_dummy_magic_23_0.VD2.n9 0.563
R7913 two_stage_opamp_dummy_magic_23_0.VD2.n16 two_stage_opamp_dummy_magic_23_0.VD2.n1 0.3755
R7914 two_stage_opamp_dummy_magic_23_0.VD2.n37 two_stage_opamp_dummy_magic_23_0.VD2.n36 0.234875
R7915 two_stage_opamp_dummy_magic_23_0.VD2.n37 two_stage_opamp_dummy_magic_23_0.VD2.n17 0.234875
R7916 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t21 610.534
R7917 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t19 610.534
R7918 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t30 433.8
R7919 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t27 433.8
R7920 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t16 433.8
R7921 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t24 433.8
R7922 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t13 433.8
R7923 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t23 433.8
R7924 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t12 433.8
R7925 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t22 433.8
R7926 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t25 433.8
R7927 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t14 433.8
R7928 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t31 433.8
R7929 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t20 433.8
R7930 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t29 433.8
R7931 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t18 433.8
R7932 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t28 433.8
R7933 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t17 433.8
R7934 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t26 433.8
R7935 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t15 433.8
R7936 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 339.836
R7937 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 339.834
R7938 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 339.272
R7939 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 287.264
R7940 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 176.733
R7941 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 176.733
R7942 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 176.733
R7943 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 176.733
R7944 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 176.733
R7945 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 176.733
R7946 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 176.733
R7947 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 176.733
R7948 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 176.733
R7949 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 176.733
R7950 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 176.733
R7951 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 176.733
R7952 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 176.733
R7953 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 176.733
R7954 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 176.733
R7955 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 176.733
R7956 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 162.508
R7957 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 107.689
R7958 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 56.2338
R7959 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 56.2338
R7960 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 52.01
R7961 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 50.5797
R7962 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 49.3505
R7963 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t9 39.4005
R7964 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t5 39.4005
R7965 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t10 39.4005
R7966 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t6 39.4005
R7967 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t7 39.4005
R7968 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t4 39.4005
R7969 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t11 39.4005
R7970 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t8 39.4005
R7971 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t3 16.0005
R7972 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t1 16.0005
R7973 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t0 16.0005
R7974 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t2 16.0005
R7975 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 10.7922
R7976 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 1.04217
R7977 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 0.563
R7978 two_stage_opamp_dummy_magic_23_0.V_source.n48 two_stage_opamp_dummy_magic_23_0.V_source.t2 66.2047
R7979 two_stage_opamp_dummy_magic_23_0.V_source.n5 two_stage_opamp_dummy_magic_23_0.V_source.n4 49.3505
R7980 two_stage_opamp_dummy_magic_23_0.V_source.n8 two_stage_opamp_dummy_magic_23_0.V_source.n7 49.3505
R7981 two_stage_opamp_dummy_magic_23_0.V_source.n11 two_stage_opamp_dummy_magic_23_0.V_source.n10 49.3505
R7982 two_stage_opamp_dummy_magic_23_0.V_source.n14 two_stage_opamp_dummy_magic_23_0.V_source.n13 49.3505
R7983 two_stage_opamp_dummy_magic_23_0.V_source.n18 two_stage_opamp_dummy_magic_23_0.V_source.n17 49.3505
R7984 two_stage_opamp_dummy_magic_23_0.V_source.n23 two_stage_opamp_dummy_magic_23_0.V_source.n22 49.3505
R7985 two_stage_opamp_dummy_magic_23_0.V_source.n25 two_stage_opamp_dummy_magic_23_0.V_source.n24 49.3505
R7986 two_stage_opamp_dummy_magic_23_0.V_source.n29 two_stage_opamp_dummy_magic_23_0.V_source.n28 49.3505
R7987 two_stage_opamp_dummy_magic_23_0.V_source.n32 two_stage_opamp_dummy_magic_23_0.V_source.n31 49.3505
R7988 two_stage_opamp_dummy_magic_23_0.V_source.n35 two_stage_opamp_dummy_magic_23_0.V_source.n34 49.3505
R7989 two_stage_opamp_dummy_magic_23_0.V_source.n40 two_stage_opamp_dummy_magic_23_0.V_source.n39 32.3838
R7990 two_stage_opamp_dummy_magic_23_0.V_source.n42 two_stage_opamp_dummy_magic_23_0.V_source.n41 32.3838
R7991 two_stage_opamp_dummy_magic_23_0.V_source.n47 two_stage_opamp_dummy_magic_23_0.V_source.n46 32.3838
R7992 two_stage_opamp_dummy_magic_23_0.V_source.n51 two_stage_opamp_dummy_magic_23_0.V_source.n50 32.3838
R7993 two_stage_opamp_dummy_magic_23_0.V_source.n55 two_stage_opamp_dummy_magic_23_0.V_source.n54 32.3838
R7994 two_stage_opamp_dummy_magic_23_0.V_source.n58 two_stage_opamp_dummy_magic_23_0.V_source.n57 32.3838
R7995 two_stage_opamp_dummy_magic_23_0.V_source.n62 two_stage_opamp_dummy_magic_23_0.V_source.n61 32.3838
R7996 two_stage_opamp_dummy_magic_23_0.V_source.n65 two_stage_opamp_dummy_magic_23_0.V_source.n64 32.3838
R7997 two_stage_opamp_dummy_magic_23_0.V_source.n68 two_stage_opamp_dummy_magic_23_0.V_source.n67 32.3838
R7998 two_stage_opamp_dummy_magic_23_0.V_source.n72 two_stage_opamp_dummy_magic_23_0.V_source.n71 32.3838
R7999 two_stage_opamp_dummy_magic_23_0.V_source.n4 two_stage_opamp_dummy_magic_23_0.V_source.t5 16.0005
R8000 two_stage_opamp_dummy_magic_23_0.V_source.n4 two_stage_opamp_dummy_magic_23_0.V_source.t6 16.0005
R8001 two_stage_opamp_dummy_magic_23_0.V_source.n7 two_stage_opamp_dummy_magic_23_0.V_source.t9 16.0005
R8002 two_stage_opamp_dummy_magic_23_0.V_source.n7 two_stage_opamp_dummy_magic_23_0.V_source.t8 16.0005
R8003 two_stage_opamp_dummy_magic_23_0.V_source.n10 two_stage_opamp_dummy_magic_23_0.V_source.t13 16.0005
R8004 two_stage_opamp_dummy_magic_23_0.V_source.n10 two_stage_opamp_dummy_magic_23_0.V_source.t40 16.0005
R8005 two_stage_opamp_dummy_magic_23_0.V_source.n13 two_stage_opamp_dummy_magic_23_0.V_source.t17 16.0005
R8006 two_stage_opamp_dummy_magic_23_0.V_source.n13 two_stage_opamp_dummy_magic_23_0.V_source.t4 16.0005
R8007 two_stage_opamp_dummy_magic_23_0.V_source.n17 two_stage_opamp_dummy_magic_23_0.V_source.t16 16.0005
R8008 two_stage_opamp_dummy_magic_23_0.V_source.n17 two_stage_opamp_dummy_magic_23_0.V_source.t1 16.0005
R8009 two_stage_opamp_dummy_magic_23_0.V_source.n22 two_stage_opamp_dummy_magic_23_0.V_source.t0 16.0005
R8010 two_stage_opamp_dummy_magic_23_0.V_source.n22 two_stage_opamp_dummy_magic_23_0.V_source.t15 16.0005
R8011 two_stage_opamp_dummy_magic_23_0.V_source.n24 two_stage_opamp_dummy_magic_23_0.V_source.t10 16.0005
R8012 two_stage_opamp_dummy_magic_23_0.V_source.n24 two_stage_opamp_dummy_magic_23_0.V_source.t7 16.0005
R8013 two_stage_opamp_dummy_magic_23_0.V_source.n28 two_stage_opamp_dummy_magic_23_0.V_source.t11 16.0005
R8014 two_stage_opamp_dummy_magic_23_0.V_source.n28 two_stage_opamp_dummy_magic_23_0.V_source.t18 16.0005
R8015 two_stage_opamp_dummy_magic_23_0.V_source.n31 two_stage_opamp_dummy_magic_23_0.V_source.t19 16.0005
R8016 two_stage_opamp_dummy_magic_23_0.V_source.n31 two_stage_opamp_dummy_magic_23_0.V_source.t12 16.0005
R8017 two_stage_opamp_dummy_magic_23_0.V_source.n34 two_stage_opamp_dummy_magic_23_0.V_source.t21 16.0005
R8018 two_stage_opamp_dummy_magic_23_0.V_source.n34 two_stage_opamp_dummy_magic_23_0.V_source.t3 16.0005
R8019 two_stage_opamp_dummy_magic_23_0.V_source.n39 two_stage_opamp_dummy_magic_23_0.V_source.t20 9.6005
R8020 two_stage_opamp_dummy_magic_23_0.V_source.n39 two_stage_opamp_dummy_magic_23_0.V_source.t14 9.6005
R8021 two_stage_opamp_dummy_magic_23_0.V_source.n41 two_stage_opamp_dummy_magic_23_0.V_source.t32 9.6005
R8022 two_stage_opamp_dummy_magic_23_0.V_source.n41 two_stage_opamp_dummy_magic_23_0.V_source.t36 9.6005
R8023 two_stage_opamp_dummy_magic_23_0.V_source.n46 two_stage_opamp_dummy_magic_23_0.V_source.t26 9.6005
R8024 two_stage_opamp_dummy_magic_23_0.V_source.n46 two_stage_opamp_dummy_magic_23_0.V_source.t34 9.6005
R8025 two_stage_opamp_dummy_magic_23_0.V_source.n50 two_stage_opamp_dummy_magic_23_0.V_source.t24 9.6005
R8026 two_stage_opamp_dummy_magic_23_0.V_source.n50 two_stage_opamp_dummy_magic_23_0.V_source.t33 9.6005
R8027 two_stage_opamp_dummy_magic_23_0.V_source.n54 two_stage_opamp_dummy_magic_23_0.V_source.t23 9.6005
R8028 two_stage_opamp_dummy_magic_23_0.V_source.n54 two_stage_opamp_dummy_magic_23_0.V_source.t31 9.6005
R8029 two_stage_opamp_dummy_magic_23_0.V_source.n57 two_stage_opamp_dummy_magic_23_0.V_source.t22 9.6005
R8030 two_stage_opamp_dummy_magic_23_0.V_source.n57 two_stage_opamp_dummy_magic_23_0.V_source.t37 9.6005
R8031 two_stage_opamp_dummy_magic_23_0.V_source.n61 two_stage_opamp_dummy_magic_23_0.V_source.t27 9.6005
R8032 two_stage_opamp_dummy_magic_23_0.V_source.n61 two_stage_opamp_dummy_magic_23_0.V_source.t30 9.6005
R8033 two_stage_opamp_dummy_magic_23_0.V_source.n64 two_stage_opamp_dummy_magic_23_0.V_source.t35 9.6005
R8034 two_stage_opamp_dummy_magic_23_0.V_source.n64 two_stage_opamp_dummy_magic_23_0.V_source.t25 9.6005
R8035 two_stage_opamp_dummy_magic_23_0.V_source.n67 two_stage_opamp_dummy_magic_23_0.V_source.t38 9.6005
R8036 two_stage_opamp_dummy_magic_23_0.V_source.n67 two_stage_opamp_dummy_magic_23_0.V_source.t28 9.6005
R8037 two_stage_opamp_dummy_magic_23_0.V_source.t39 two_stage_opamp_dummy_magic_23_0.V_source.n72 9.6005
R8038 two_stage_opamp_dummy_magic_23_0.V_source.n72 two_stage_opamp_dummy_magic_23_0.V_source.t29 9.6005
R8039 two_stage_opamp_dummy_magic_23_0.V_source.n69 two_stage_opamp_dummy_magic_23_0.V_source.n65 5.89633
R8040 two_stage_opamp_dummy_magic_23_0.V_source.n40 two_stage_opamp_dummy_magic_23_0.V_source.n3 5.89633
R8041 two_stage_opamp_dummy_magic_23_0.V_source.n66 two_stage_opamp_dummy_magic_23_0.V_source.n65 5.70883
R8042 two_stage_opamp_dummy_magic_23_0.V_source.n43 two_stage_opamp_dummy_magic_23_0.V_source.n40 5.70883
R8043 two_stage_opamp_dummy_magic_23_0.V_source.n26 two_stage_opamp_dummy_magic_23_0.V_source.n23 5.6255
R8044 two_stage_opamp_dummy_magic_23_0.V_source.n9 two_stage_opamp_dummy_magic_23_0.V_source.n8 5.6255
R8045 two_stage_opamp_dummy_magic_23_0.V_source.n35 two_stage_opamp_dummy_magic_23_0.V_source.n33 5.45883
R8046 two_stage_opamp_dummy_magic_23_0.V_source.n23 two_stage_opamp_dummy_magic_23_0.V_source.n21 5.45883
R8047 two_stage_opamp_dummy_magic_23_0.V_source.n12 two_stage_opamp_dummy_magic_23_0.V_source.n8 5.45883
R8048 two_stage_opamp_dummy_magic_23_0.V_source.n16 two_stage_opamp_dummy_magic_23_0.V_source.n5 5.45883
R8049 two_stage_opamp_dummy_magic_23_0.V_source.n42 two_stage_opamp_dummy_magic_23_0.V_source.n3 5.33383
R8050 two_stage_opamp_dummy_magic_23_0.V_source.n52 two_stage_opamp_dummy_magic_23_0.V_source.n51 5.33383
R8051 two_stage_opamp_dummy_magic_23_0.V_source.n55 two_stage_opamp_dummy_magic_23_0.V_source.n53 5.33383
R8052 two_stage_opamp_dummy_magic_23_0.V_source.n58 two_stage_opamp_dummy_magic_23_0.V_source.n1 5.33383
R8053 two_stage_opamp_dummy_magic_23_0.V_source.n63 two_stage_opamp_dummy_magic_23_0.V_source.n62 5.33383
R8054 two_stage_opamp_dummy_magic_23_0.V_source.n69 two_stage_opamp_dummy_magic_23_0.V_source.n68 5.33383
R8055 two_stage_opamp_dummy_magic_23_0.V_source.n71 two_stage_opamp_dummy_magic_23_0.V_source.n70 5.33383
R8056 two_stage_opamp_dummy_magic_23_0.V_source.n43 two_stage_opamp_dummy_magic_23_0.V_source.n42 5.14633
R8057 two_stage_opamp_dummy_magic_23_0.V_source.n51 two_stage_opamp_dummy_magic_23_0.V_source.n2 5.14633
R8058 two_stage_opamp_dummy_magic_23_0.V_source.n56 two_stage_opamp_dummy_magic_23_0.V_source.n55 5.14633
R8059 two_stage_opamp_dummy_magic_23_0.V_source.n59 two_stage_opamp_dummy_magic_23_0.V_source.n58 5.14633
R8060 two_stage_opamp_dummy_magic_23_0.V_source.n62 two_stage_opamp_dummy_magic_23_0.V_source.n60 5.14633
R8061 two_stage_opamp_dummy_magic_23_0.V_source.n71 two_stage_opamp_dummy_magic_23_0.V_source.n0 5.14633
R8062 two_stage_opamp_dummy_magic_23_0.V_source.n68 two_stage_opamp_dummy_magic_23_0.V_source.n66 5.14633
R8063 two_stage_opamp_dummy_magic_23_0.V_source.n11 two_stage_opamp_dummy_magic_23_0.V_source.n9 5.063
R8064 two_stage_opamp_dummy_magic_23_0.V_source.n14 two_stage_opamp_dummy_magic_23_0.V_source.n6 5.063
R8065 two_stage_opamp_dummy_magic_23_0.V_source.n19 two_stage_opamp_dummy_magic_23_0.V_source.n18 5.063
R8066 two_stage_opamp_dummy_magic_23_0.V_source.n26 two_stage_opamp_dummy_magic_23_0.V_source.n25 5.063
R8067 two_stage_opamp_dummy_magic_23_0.V_source.n29 two_stage_opamp_dummy_magic_23_0.V_source.n27 5.063
R8068 two_stage_opamp_dummy_magic_23_0.V_source.n32 two_stage_opamp_dummy_magic_23_0.V_source.n20 5.063
R8069 two_stage_opamp_dummy_magic_23_0.V_source.n36 two_stage_opamp_dummy_magic_23_0.V_source.n35 5.063
R8070 two_stage_opamp_dummy_magic_23_0.V_source.n12 two_stage_opamp_dummy_magic_23_0.V_source.n11 4.89633
R8071 two_stage_opamp_dummy_magic_23_0.V_source.n15 two_stage_opamp_dummy_magic_23_0.V_source.n14 4.89633
R8072 two_stage_opamp_dummy_magic_23_0.V_source.n18 two_stage_opamp_dummy_magic_23_0.V_source.n16 4.89633
R8073 two_stage_opamp_dummy_magic_23_0.V_source.n25 two_stage_opamp_dummy_magic_23_0.V_source.n21 4.89633
R8074 two_stage_opamp_dummy_magic_23_0.V_source.n30 two_stage_opamp_dummy_magic_23_0.V_source.n29 4.89633
R8075 two_stage_opamp_dummy_magic_23_0.V_source.n33 two_stage_opamp_dummy_magic_23_0.V_source.n32 4.89633
R8076 two_stage_opamp_dummy_magic_23_0.V_source.n38 two_stage_opamp_dummy_magic_23_0.V_source.n37 4.5005
R8077 two_stage_opamp_dummy_magic_23_0.V_source.n45 two_stage_opamp_dummy_magic_23_0.V_source.n44 4.5005
R8078 two_stage_opamp_dummy_magic_23_0.V_source.n49 two_stage_opamp_dummy_magic_23_0.V_source.n48 4.5005
R8079 two_stage_opamp_dummy_magic_23_0.V_source.n37 two_stage_opamp_dummy_magic_23_0.V_source.n36 3.6255
R8080 two_stage_opamp_dummy_magic_23_0.V_source.n45 two_stage_opamp_dummy_magic_23_0.V_source.n38 1.738
R8081 two_stage_opamp_dummy_magic_23_0.V_source.n48 two_stage_opamp_dummy_magic_23_0.V_source.n47 0.833833
R8082 two_stage_opamp_dummy_magic_23_0.V_source.n47 two_stage_opamp_dummy_magic_23_0.V_source.n45 0.633833
R8083 two_stage_opamp_dummy_magic_23_0.V_source.n33 two_stage_opamp_dummy_magic_23_0.V_source.n30 0.563
R8084 two_stage_opamp_dummy_magic_23_0.V_source.n30 two_stage_opamp_dummy_magic_23_0.V_source.n21 0.563
R8085 two_stage_opamp_dummy_magic_23_0.V_source.n27 two_stage_opamp_dummy_magic_23_0.V_source.n26 0.563
R8086 two_stage_opamp_dummy_magic_23_0.V_source.n27 two_stage_opamp_dummy_magic_23_0.V_source.n20 0.563
R8087 two_stage_opamp_dummy_magic_23_0.V_source.n36 two_stage_opamp_dummy_magic_23_0.V_source.n20 0.563
R8088 two_stage_opamp_dummy_magic_23_0.V_source.n37 two_stage_opamp_dummy_magic_23_0.V_source.n19 0.563
R8089 two_stage_opamp_dummy_magic_23_0.V_source.n19 two_stage_opamp_dummy_magic_23_0.V_source.n6 0.563
R8090 two_stage_opamp_dummy_magic_23_0.V_source.n9 two_stage_opamp_dummy_magic_23_0.V_source.n6 0.563
R8091 two_stage_opamp_dummy_magic_23_0.V_source.n15 two_stage_opamp_dummy_magic_23_0.V_source.n12 0.563
R8092 two_stage_opamp_dummy_magic_23_0.V_source.n16 two_stage_opamp_dummy_magic_23_0.V_source.n15 0.563
R8093 two_stage_opamp_dummy_magic_23_0.V_source.n38 two_stage_opamp_dummy_magic_23_0.V_source.n5 0.563
R8094 two_stage_opamp_dummy_magic_23_0.V_source.n70 two_stage_opamp_dummy_magic_23_0.V_source.n69 0.563
R8095 two_stage_opamp_dummy_magic_23_0.V_source.n66 two_stage_opamp_dummy_magic_23_0.V_source.n0 0.563
R8096 two_stage_opamp_dummy_magic_23_0.V_source.n60 two_stage_opamp_dummy_magic_23_0.V_source.n0 0.563
R8097 two_stage_opamp_dummy_magic_23_0.V_source.n60 two_stage_opamp_dummy_magic_23_0.V_source.n59 0.563
R8098 two_stage_opamp_dummy_magic_23_0.V_source.n59 two_stage_opamp_dummy_magic_23_0.V_source.n56 0.563
R8099 two_stage_opamp_dummy_magic_23_0.V_source.n56 two_stage_opamp_dummy_magic_23_0.V_source.n2 0.563
R8100 two_stage_opamp_dummy_magic_23_0.V_source.n44 two_stage_opamp_dummy_magic_23_0.V_source.n2 0.563
R8101 two_stage_opamp_dummy_magic_23_0.V_source.n44 two_stage_opamp_dummy_magic_23_0.V_source.n43 0.563
R8102 two_stage_opamp_dummy_magic_23_0.V_source.n49 two_stage_opamp_dummy_magic_23_0.V_source.n3 0.563
R8103 two_stage_opamp_dummy_magic_23_0.V_source.n52 two_stage_opamp_dummy_magic_23_0.V_source.n49 0.563
R8104 two_stage_opamp_dummy_magic_23_0.V_source.n53 two_stage_opamp_dummy_magic_23_0.V_source.n52 0.563
R8105 two_stage_opamp_dummy_magic_23_0.V_source.n53 two_stage_opamp_dummy_magic_23_0.V_source.n1 0.563
R8106 two_stage_opamp_dummy_magic_23_0.V_source.n63 two_stage_opamp_dummy_magic_23_0.V_source.n1 0.563
R8107 two_stage_opamp_dummy_magic_23_0.V_source.n70 two_stage_opamp_dummy_magic_23_0.V_source.n63 0.563
R8108 two_stage_opamp_dummy_magic_23_0.VD4.n10 two_stage_opamp_dummy_magic_23_0.VD4.t0 672.293
R8109 two_stage_opamp_dummy_magic_23_0.VD4.n13 two_stage_opamp_dummy_magic_23_0.VD4.t3 672.293
R8110 two_stage_opamp_dummy_magic_23_0.VD4.t1 two_stage_opamp_dummy_magic_23_0.VD4.n11 213.131
R8111 two_stage_opamp_dummy_magic_23_0.VD4.n12 two_stage_opamp_dummy_magic_23_0.VD4.t4 213.131
R8112 two_stage_opamp_dummy_magic_23_0.VD4.t20 two_stage_opamp_dummy_magic_23_0.VD4.t1 146.155
R8113 two_stage_opamp_dummy_magic_23_0.VD4.t24 two_stage_opamp_dummy_magic_23_0.VD4.t20 146.155
R8114 two_stage_opamp_dummy_magic_23_0.VD4.t30 two_stage_opamp_dummy_magic_23_0.VD4.t24 146.155
R8115 two_stage_opamp_dummy_magic_23_0.VD4.t34 two_stage_opamp_dummy_magic_23_0.VD4.t30 146.155
R8116 two_stage_opamp_dummy_magic_23_0.VD4.t36 two_stage_opamp_dummy_magic_23_0.VD4.t34 146.155
R8117 two_stage_opamp_dummy_magic_23_0.VD4.t18 two_stage_opamp_dummy_magic_23_0.VD4.t36 146.155
R8118 two_stage_opamp_dummy_magic_23_0.VD4.t22 two_stage_opamp_dummy_magic_23_0.VD4.t18 146.155
R8119 two_stage_opamp_dummy_magic_23_0.VD4.t26 two_stage_opamp_dummy_magic_23_0.VD4.t22 146.155
R8120 two_stage_opamp_dummy_magic_23_0.VD4.t32 two_stage_opamp_dummy_magic_23_0.VD4.t26 146.155
R8121 two_stage_opamp_dummy_magic_23_0.VD4.t28 two_stage_opamp_dummy_magic_23_0.VD4.t32 146.155
R8122 two_stage_opamp_dummy_magic_23_0.VD4.t4 two_stage_opamp_dummy_magic_23_0.VD4.t28 146.155
R8123 two_stage_opamp_dummy_magic_23_0.VD4.n11 two_stage_opamp_dummy_magic_23_0.VD4.t2 76.2576
R8124 two_stage_opamp_dummy_magic_23_0.VD4.n12 two_stage_opamp_dummy_magic_23_0.VD4.t5 76.2576
R8125 two_stage_opamp_dummy_magic_23_0.VD4.n7 two_stage_opamp_dummy_magic_23_0.VD4.n6 71.513
R8126 two_stage_opamp_dummy_magic_23_0.VD4.n9 two_stage_opamp_dummy_magic_23_0.VD4.n8 71.513
R8127 two_stage_opamp_dummy_magic_23_0.VD4.n1 two_stage_opamp_dummy_magic_23_0.VD4.n0 71.513
R8128 two_stage_opamp_dummy_magic_23_0.VD4.n3 two_stage_opamp_dummy_magic_23_0.VD4.n2 71.513
R8129 two_stage_opamp_dummy_magic_23_0.VD4.n5 two_stage_opamp_dummy_magic_23_0.VD4.n4 71.513
R8130 two_stage_opamp_dummy_magic_23_0.VD4.n18 two_stage_opamp_dummy_magic_23_0.VD4.n17 66.0338
R8131 two_stage_opamp_dummy_magic_23_0.VD4.n21 two_stage_opamp_dummy_magic_23_0.VD4.n20 66.0338
R8132 two_stage_opamp_dummy_magic_23_0.VD4.n24 two_stage_opamp_dummy_magic_23_0.VD4.n23 66.0338
R8133 two_stage_opamp_dummy_magic_23_0.VD4.n28 two_stage_opamp_dummy_magic_23_0.VD4.n27 66.0338
R8134 two_stage_opamp_dummy_magic_23_0.VD4.n31 two_stage_opamp_dummy_magic_23_0.VD4.n30 66.0338
R8135 two_stage_opamp_dummy_magic_23_0.VD4.n34 two_stage_opamp_dummy_magic_23_0.VD4.n33 66.0338
R8136 two_stage_opamp_dummy_magic_23_0.VD4.n6 two_stage_opamp_dummy_magic_23_0.VD4.t31 11.2576
R8137 two_stage_opamp_dummy_magic_23_0.VD4.n6 two_stage_opamp_dummy_magic_23_0.VD4.t35 11.2576
R8138 two_stage_opamp_dummy_magic_23_0.VD4.n8 two_stage_opamp_dummy_magic_23_0.VD4.t21 11.2576
R8139 two_stage_opamp_dummy_magic_23_0.VD4.n8 two_stage_opamp_dummy_magic_23_0.VD4.t25 11.2576
R8140 two_stage_opamp_dummy_magic_23_0.VD4.n17 two_stage_opamp_dummy_magic_23_0.VD4.t8 11.2576
R8141 two_stage_opamp_dummy_magic_23_0.VD4.n17 two_stage_opamp_dummy_magic_23_0.VD4.t16 11.2576
R8142 two_stage_opamp_dummy_magic_23_0.VD4.n20 two_stage_opamp_dummy_magic_23_0.VD4.t14 11.2576
R8143 two_stage_opamp_dummy_magic_23_0.VD4.n20 two_stage_opamp_dummy_magic_23_0.VD4.t7 11.2576
R8144 two_stage_opamp_dummy_magic_23_0.VD4.n23 two_stage_opamp_dummy_magic_23_0.VD4.t12 11.2576
R8145 two_stage_opamp_dummy_magic_23_0.VD4.n23 two_stage_opamp_dummy_magic_23_0.VD4.t11 11.2576
R8146 two_stage_opamp_dummy_magic_23_0.VD4.n27 two_stage_opamp_dummy_magic_23_0.VD4.t9 11.2576
R8147 two_stage_opamp_dummy_magic_23_0.VD4.n27 two_stage_opamp_dummy_magic_23_0.VD4.t10 11.2576
R8148 two_stage_opamp_dummy_magic_23_0.VD4.n30 two_stage_opamp_dummy_magic_23_0.VD4.t13 11.2576
R8149 two_stage_opamp_dummy_magic_23_0.VD4.n30 two_stage_opamp_dummy_magic_23_0.VD4.t6 11.2576
R8150 two_stage_opamp_dummy_magic_23_0.VD4.n33 two_stage_opamp_dummy_magic_23_0.VD4.t17 11.2576
R8151 two_stage_opamp_dummy_magic_23_0.VD4.n33 two_stage_opamp_dummy_magic_23_0.VD4.t15 11.2576
R8152 two_stage_opamp_dummy_magic_23_0.VD4.n0 two_stage_opamp_dummy_magic_23_0.VD4.t33 11.2576
R8153 two_stage_opamp_dummy_magic_23_0.VD4.n0 two_stage_opamp_dummy_magic_23_0.VD4.t29 11.2576
R8154 two_stage_opamp_dummy_magic_23_0.VD4.n2 two_stage_opamp_dummy_magic_23_0.VD4.t23 11.2576
R8155 two_stage_opamp_dummy_magic_23_0.VD4.n2 two_stage_opamp_dummy_magic_23_0.VD4.t27 11.2576
R8156 two_stage_opamp_dummy_magic_23_0.VD4.n4 two_stage_opamp_dummy_magic_23_0.VD4.t37 11.2576
R8157 two_stage_opamp_dummy_magic_23_0.VD4.n4 two_stage_opamp_dummy_magic_23_0.VD4.t19 11.2576
R8158 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.VD4.n35 8.59425
R8159 two_stage_opamp_dummy_magic_23_0.VD4.n10 two_stage_opamp_dummy_magic_23_0.VD4.n9 6.10467
R8160 two_stage_opamp_dummy_magic_23_0.VD4.n34 two_stage_opamp_dummy_magic_23_0.VD4.n32 5.91717
R8161 two_stage_opamp_dummy_magic_23_0.VD4.n19 two_stage_opamp_dummy_magic_23_0.VD4.n18 5.91717
R8162 two_stage_opamp_dummy_magic_23_0.VD4.n22 two_stage_opamp_dummy_magic_23_0.VD4.n18 5.91717
R8163 two_stage_opamp_dummy_magic_23_0.VD4.n14 two_stage_opamp_dummy_magic_23_0.VD4.n13 5.47967
R8164 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.VD4.n14 5.3755
R8165 two_stage_opamp_dummy_magic_23_0.VD4.n22 two_stage_opamp_dummy_magic_23_0.VD4.n21 5.29217
R8166 two_stage_opamp_dummy_magic_23_0.VD4.n21 two_stage_opamp_dummy_magic_23_0.VD4.n19 5.29217
R8167 two_stage_opamp_dummy_magic_23_0.VD4.n25 two_stage_opamp_dummy_magic_23_0.VD4.n24 5.29217
R8168 two_stage_opamp_dummy_magic_23_0.VD4.n24 two_stage_opamp_dummy_magic_23_0.VD4.n16 5.29217
R8169 two_stage_opamp_dummy_magic_23_0.VD4.n28 two_stage_opamp_dummy_magic_23_0.VD4.n26 5.29217
R8170 two_stage_opamp_dummy_magic_23_0.VD4.n29 two_stage_opamp_dummy_magic_23_0.VD4.n28 5.29217
R8171 two_stage_opamp_dummy_magic_23_0.VD4.n31 two_stage_opamp_dummy_magic_23_0.VD4.n15 5.29217
R8172 two_stage_opamp_dummy_magic_23_0.VD4.n32 two_stage_opamp_dummy_magic_23_0.VD4.n31 5.29217
R8173 two_stage_opamp_dummy_magic_23_0.VD4.n35 two_stage_opamp_dummy_magic_23_0.VD4.n34 5.29217
R8174 two_stage_opamp_dummy_magic_23_0.VD4.n13 two_stage_opamp_dummy_magic_23_0.VD4.n12 1.03383
R8175 two_stage_opamp_dummy_magic_23_0.VD4.n11 two_stage_opamp_dummy_magic_23_0.VD4.n10 1.03383
R8176 two_stage_opamp_dummy_magic_23_0.VD4.n32 two_stage_opamp_dummy_magic_23_0.VD4.n29 0.6255
R8177 two_stage_opamp_dummy_magic_23_0.VD4.n29 two_stage_opamp_dummy_magic_23_0.VD4.n16 0.6255
R8178 two_stage_opamp_dummy_magic_23_0.VD4.n19 two_stage_opamp_dummy_magic_23_0.VD4.n16 0.6255
R8179 two_stage_opamp_dummy_magic_23_0.VD4.n25 two_stage_opamp_dummy_magic_23_0.VD4.n22 0.6255
R8180 two_stage_opamp_dummy_magic_23_0.VD4.n26 two_stage_opamp_dummy_magic_23_0.VD4.n25 0.6255
R8181 two_stage_opamp_dummy_magic_23_0.VD4.n26 two_stage_opamp_dummy_magic_23_0.VD4.n15 0.6255
R8182 two_stage_opamp_dummy_magic_23_0.VD4.n35 two_stage_opamp_dummy_magic_23_0.VD4.n15 0.6255
R8183 two_stage_opamp_dummy_magic_23_0.VD4.n5 two_stage_opamp_dummy_magic_23_0.VD4.n3 0.6255
R8184 two_stage_opamp_dummy_magic_23_0.VD4.n3 two_stage_opamp_dummy_magic_23_0.VD4.n1 0.6255
R8185 two_stage_opamp_dummy_magic_23_0.VD4.n14 two_stage_opamp_dummy_magic_23_0.VD4.n1 0.6255
R8186 two_stage_opamp_dummy_magic_23_0.VD4.n9 two_stage_opamp_dummy_magic_23_0.VD4.n7 0.6255
R8187 two_stage_opamp_dummy_magic_23_0.VD4.n7 two_stage_opamp_dummy_magic_23_0.VD4.n5 0.6255
R8188 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 129.005
R8189 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 118.861
R8190 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 118.861
R8191 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 118.861
R8192 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 118.861
R8193 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 118.861
R8194 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t3 19.7005
R8195 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t7 19.7005
R8196 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t2 19.7005
R8197 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t9 19.7005
R8198 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t4 19.7005
R8199 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t8 19.7005
R8200 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t5 19.7005
R8201 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t10 19.7005
R8202 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t6 19.7005
R8203 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t1 19.7005
R8204 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 5.60467
R8205 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 5.54217
R8206 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 5.54217
R8207 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 5.04217
R8208 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 5.04217
R8209 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 5.04217
R8210 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 5.04217
R8211 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 4.97967
R8212 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 4.97967
R8213 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 4.97967
R8214 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 0.563
R8215 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 0.563
R8216 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 0.563
R8217 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 0.563
R8218 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 0.563
R8219 two_stage_opamp_dummy_magic_23_0.Vb2_2.n2 two_stage_opamp_dummy_magic_23_0.Vb2_2.t3 661.375
R8220 two_stage_opamp_dummy_magic_23_0.Vb2_2.n4 two_stage_opamp_dummy_magic_23_0.Vb2_2.t0 661.375
R8221 two_stage_opamp_dummy_magic_23_0.Vb2_2.t4 two_stage_opamp_dummy_magic_23_0.Vb2_2.n0 213.131
R8222 two_stage_opamp_dummy_magic_23_0.Vb2_2.n3 two_stage_opamp_dummy_magic_23_0.Vb2_2.t1 213.131
R8223 two_stage_opamp_dummy_magic_23_0.Vb2_2.n6 two_stage_opamp_dummy_magic_23_0.Vb2_2.n1 154.983
R8224 two_stage_opamp_dummy_magic_23_0.Vb2_2.t7 two_stage_opamp_dummy_magic_23_0.Vb2_2.t4 146.155
R8225 two_stage_opamp_dummy_magic_23_0.Vb2_2.t1 two_stage_opamp_dummy_magic_23_0.Vb2_2.t7 146.155
R8226 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n0 76.2576
R8227 two_stage_opamp_dummy_magic_23_0.Vb2_2.n3 two_stage_opamp_dummy_magic_23_0.Vb2_2.t2 76.2576
R8228 two_stage_opamp_dummy_magic_23_0.Vb2_2.n7 two_stage_opamp_dummy_magic_23_0.Vb2_2.n6 66.4421
R8229 two_stage_opamp_dummy_magic_23_0.Vb2_2.n1 two_stage_opamp_dummy_magic_23_0.Vb2_2.t6 21.8894
R8230 two_stage_opamp_dummy_magic_23_0.Vb2_2.n1 two_stage_opamp_dummy_magic_23_0.Vb2_2.t9 21.8894
R8231 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n7 11.2576
R8232 two_stage_opamp_dummy_magic_23_0.Vb2_2.n7 two_stage_opamp_dummy_magic_23_0.Vb2_2.t8 11.2576
R8233 two_stage_opamp_dummy_magic_23_0.Vb2_2.n5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n4 5.1255
R8234 two_stage_opamp_dummy_magic_23_0.Vb2_2.n6 two_stage_opamp_dummy_magic_23_0.Vb2_2.n5 4.92067
R8235 two_stage_opamp_dummy_magic_23_0.Vb2_2.n5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n2 4.7505
R8236 two_stage_opamp_dummy_magic_23_0.Vb2_2.n4 two_stage_opamp_dummy_magic_23_0.Vb2_2.n3 1.888
R8237 two_stage_opamp_dummy_magic_23_0.Vb2_2.n2 two_stage_opamp_dummy_magic_23_0.Vb2_2.n0 1.888
R8238 a_6470_23450.t0 a_6470_23450.t1 178.133
R8239 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t14 120.504
R8240 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 107.121
R8241 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 97.4332
R8242 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 40.5317
R8243 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 39.2193
R8244 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 24.288
R8245 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 24.288
R8246 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 24.288
R8247 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 24.288
R8248 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 24.288
R8249 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t3 24.0005
R8250 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t0 24.0005
R8251 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t2 24.0005
R8252 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t1 24.0005
R8253 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t4 8.0005
R8254 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t8 8.0005
R8255 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t13 8.0005
R8256 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t11 8.0005
R8257 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t6 8.0005
R8258 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t10 8.0005
R8259 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t5 8.0005
R8260 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t9 8.0005
R8261 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t12 8.0005
R8262 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t7 8.0005
R8263 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 6.0005
R8264 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 5.7505
R8265 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 5.7505
R8266 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 5.7505
R8267 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 5.188
R8268 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 5.188
R8269 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 5.188
R8270 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 5.188
R8271 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 5.188
R8272 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 5.188
R8273 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 5.188
R8274 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 0.563
R8275 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 0.563
R8276 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 0.563
R8277 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 0.563
R8278 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 0.563
R8279 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t15 739.067
R8280 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 724.936
R8281 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t10 540.458
R8282 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 530.201
R8283 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 530.201
R8284 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 530.201
R8285 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 361.5
R8286 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t12 208.868
R8287 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t8 208.868
R8288 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t13 208.868
R8289 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t7 208.868
R8290 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t14 208.868
R8291 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t9 208.868
R8292 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t16 208.868
R8293 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t11 208.868
R8294 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t17 208.868
R8295 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 176.733
R8296 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 176.733
R8297 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 176.733
R8298 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 176.733
R8299 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 173.654
R8300 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 169.279
R8301 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 169.279
R8302 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t6 126.361
R8303 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 50.2817
R8304 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t3 13.1338
R8305 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t1 13.1338
R8306 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t2 13.1338
R8307 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t5 13.1338
R8308 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t0 13.1338
R8309 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t4 13.1338
R8310 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 10.0317
R8311 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 4.3755
R8312 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 3.6255
R8313 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 594.301
R8314 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 594.301
R8315 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 594.301
R8316 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 594.301
R8317 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 594.301
R8318 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 594.301
R8319 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 594.301
R8320 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 594.301
R8321 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 594.301
R8322 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 594.301
R8323 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 594.301
R8324 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 two_stage_opamp_dummy_magic_23_0.V_err_p.t6 78.8005
R8325 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 two_stage_opamp_dummy_magic_23_0.V_err_p.t18 78.8005
R8326 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 two_stage_opamp_dummy_magic_23_0.V_err_p.t21 78.8005
R8327 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 two_stage_opamp_dummy_magic_23_0.V_err_p.t7 78.8005
R8328 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 two_stage_opamp_dummy_magic_23_0.V_err_p.t4 78.8005
R8329 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 two_stage_opamp_dummy_magic_23_0.V_err_p.t9 78.8005
R8330 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 two_stage_opamp_dummy_magic_23_0.V_err_p.t5 78.8005
R8331 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 two_stage_opamp_dummy_magic_23_0.V_err_p.t10 78.8005
R8332 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 two_stage_opamp_dummy_magic_23_0.V_err_p.t3 78.8005
R8333 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 two_stage_opamp_dummy_magic_23_0.V_err_p.t0 78.8005
R8334 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 two_stage_opamp_dummy_magic_23_0.V_err_p.t13 78.8005
R8335 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 two_stage_opamp_dummy_magic_23_0.V_err_p.t2 78.8005
R8336 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 two_stage_opamp_dummy_magic_23_0.V_err_p.t15 78.8005
R8337 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 two_stage_opamp_dummy_magic_23_0.V_err_p.t11 78.8005
R8338 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 two_stage_opamp_dummy_magic_23_0.V_err_p.t1 78.8005
R8339 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 two_stage_opamp_dummy_magic_23_0.V_err_p.t16 78.8005
R8340 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 two_stage_opamp_dummy_magic_23_0.V_err_p.t12 78.8005
R8341 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 two_stage_opamp_dummy_magic_23_0.V_err_p.t17 78.8005
R8342 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 two_stage_opamp_dummy_magic_23_0.V_err_p.t20 78.8005
R8343 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 two_stage_opamp_dummy_magic_23_0.V_err_p.t14 78.8005
R8344 two_stage_opamp_dummy_magic_23_0.V_err_p.t19 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 78.8005
R8345 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 two_stage_opamp_dummy_magic_23_0.V_err_p.t8 78.8005
R8346 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 6.10467
R8347 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 6.10467
R8348 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 5.97967
R8349 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 5.94842
R8350 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 5.91717
R8351 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 5.91717
R8352 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 5.79217
R8353 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 5.41717
R8354 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 5.22967
R8355 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 5.22967
R8356 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 5.063
R8357 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 4.85467
R8358 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 4.85467
R8359 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 4.85467
R8360 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 4.85467
R8361 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 4.85467
R8362 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 4.85467
R8363 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 4.66717
R8364 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 4.66717
R8365 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 4.66717
R8366 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 4.66717
R8367 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 4.66717
R8368 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 3.7505
R8369 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 3.7505
R8370 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 two_stage_opamp_dummy_magic_23_0.err_amp_out.t12 840.595
R8371 two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 601.051
R8372 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 599.801
R8373 two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 599.801
R8374 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 194.3
R8375 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 194.3
R8376 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 194.3
R8377 two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 two_stage_opamp_dummy_magic_23_0.err_amp_out.t5 78.8005
R8378 two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 two_stage_opamp_dummy_magic_23_0.err_amp_out.t7 78.8005
R8379 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 two_stage_opamp_dummy_magic_23_0.err_amp_out.t11 78.8005
R8380 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 two_stage_opamp_dummy_magic_23_0.err_amp_out.t4 78.8005
R8381 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 two_stage_opamp_dummy_magic_23_0.err_amp_out.t6 78.8005
R8382 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 two_stage_opamp_dummy_magic_23_0.err_amp_out.t8 78.8005
R8383 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 two_stage_opamp_dummy_magic_23_0.err_amp_out.t0 48.0005
R8384 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 two_stage_opamp_dummy_magic_23_0.err_amp_out.t10 48.0005
R8385 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 two_stage_opamp_dummy_magic_23_0.err_amp_out.t3 48.0005
R8386 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 two_stage_opamp_dummy_magic_23_0.err_amp_out.t1 48.0005
R8387 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 two_stage_opamp_dummy_magic_23_0.err_amp_out.t9 48.0005
R8388 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 two_stage_opamp_dummy_magic_23_0.err_amp_out.t2 48.0005
R8389 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 6.20883
R8390 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 6.20883
R8391 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 4.95883
R8392 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 4.95883
R8393 two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 4.95883
R8394 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 4.95883
R8395 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 1.2505
R8396 two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 1.2505
R8397 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 1.2505
R8398 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 1.063
R8399 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 594.301
R8400 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 594.301
R8401 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 594.301
R8402 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 594.301
R8403 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 594.301
R8404 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 594.301
R8405 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t16 289.2
R8406 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 two_stage_opamp_dummy_magic_23_0.V_err_gate.t14 224.934
R8407 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 176.733
R8408 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 176.733
R8409 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 176.733
R8410 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 176.733
R8411 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 176.733
R8412 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 176.733
R8413 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 176.733
R8414 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 176.733
R8415 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 176.733
R8416 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 176.733
R8417 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 176.733
R8418 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 176.733
R8419 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 176.733
R8420 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 176.733
R8421 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 176.733
R8422 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 176.733
R8423 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 171.638
R8424 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 161.869
R8425 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 two_stage_opamp_dummy_magic_23_0.V_err_gate.t29 112.468
R8426 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 two_stage_opamp_dummy_magic_23_0.V_err_gate.t26 112.468
R8427 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 two_stage_opamp_dummy_magic_23_0.V_err_gate.t17 112.468
R8428 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 two_stage_opamp_dummy_magic_23_0.V_err_gate.t27 112.468
R8429 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 two_stage_opamp_dummy_magic_23_0.V_err_gate.t18 112.468
R8430 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 two_stage_opamp_dummy_magic_23_0.V_err_gate.t28 112.468
R8431 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 two_stage_opamp_dummy_magic_23_0.V_err_gate.t21 112.468
R8432 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 two_stage_opamp_dummy_magic_23_0.V_err_gate.t31 112.468
R8433 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t24 112.468
R8434 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 two_stage_opamp_dummy_magic_23_0.V_err_gate.t20 112.468
R8435 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 two_stage_opamp_dummy_magic_23_0.V_err_gate.t30 112.468
R8436 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 two_stage_opamp_dummy_magic_23_0.V_err_gate.t22 112.468
R8437 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 two_stage_opamp_dummy_magic_23_0.V_err_gate.t32 112.468
R8438 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 two_stage_opamp_dummy_magic_23_0.V_err_gate.t23 112.468
R8439 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 two_stage_opamp_dummy_magic_23_0.V_err_gate.t33 112.468
R8440 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 two_stage_opamp_dummy_magic_23_0.V_err_gate.t25 112.468
R8441 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 two_stage_opamp_dummy_magic_23_0.V_err_gate.t15 112.468
R8442 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 two_stage_opamp_dummy_magic_23_0.V_err_gate.t19 112.468
R8443 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 two_stage_opamp_dummy_magic_23_0.V_err_gate.t6 78.8005
R8444 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 two_stage_opamp_dummy_magic_23_0.V_err_gate.t11 78.8005
R8445 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 two_stage_opamp_dummy_magic_23_0.V_err_gate.t10 78.8005
R8446 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 two_stage_opamp_dummy_magic_23_0.V_err_gate.t1 78.8005
R8447 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 two_stage_opamp_dummy_magic_23_0.V_err_gate.t9 78.8005
R8448 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 two_stage_opamp_dummy_magic_23_0.V_err_gate.t8 78.8005
R8449 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 two_stage_opamp_dummy_magic_23_0.V_err_gate.t2 78.8005
R8450 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 two_stage_opamp_dummy_magic_23_0.V_err_gate.t0 78.8005
R8451 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 two_stage_opamp_dummy_magic_23_0.V_err_gate.t5 78.8005
R8452 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 two_stage_opamp_dummy_magic_23_0.V_err_gate.t7 78.8005
R8453 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 two_stage_opamp_dummy_magic_23_0.V_err_gate.t12 78.8005
R8454 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 two_stage_opamp_dummy_magic_23_0.V_err_gate.t13 78.8005
R8455 two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 56.2338
R8456 two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 56.2338
R8457 two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 two_stage_opamp_dummy_magic_23_0.V_err_gate.t3 24.0005
R8458 two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 two_stage_opamp_dummy_magic_23_0.V_err_gate.t4 24.0005
R8459 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 6.89112
R8460 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 5.41717
R8461 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 5.22967
R8462 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 5.22967
R8463 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 4.85467
R8464 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 4.85467
R8465 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 4.85467
R8466 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 4.85467
R8467 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 4.85467
R8468 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 4.66717
R8469 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 4.66717
R8470 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 4.66717
R8471 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 4.66717
R8472 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 1.688
R8473 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 1.1255
R8474 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 1.1255
R8475 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 594.301
R8476 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 594.301
R8477 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 594.301
R8478 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t18 289.2
R8479 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t11 289.2
R8480 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 194.3
R8481 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 194.3
R8482 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 194.3
R8483 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 176.733
R8484 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 176.733
R8485 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 176.733
R8486 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 176.733
R8487 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 176.733
R8488 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 161.3
R8489 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 161.3
R8490 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t7 112.468
R8491 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t15 112.468
R8492 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t20 112.468
R8493 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t17 112.468
R8494 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t13 112.468
R8495 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t19 112.468
R8496 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t21 112.468
R8497 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t9 112.468
R8498 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t3 78.8005
R8499 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t6 78.8005
R8500 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t2 78.8005
R8501 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t0 78.8005
R8502 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t1 78.8005
R8503 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t5 78.8005
R8504 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t4 48.0005
R8505 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t12 48.0005
R8506 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t14 48.0005
R8507 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t8 48.0005
R8508 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t16 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 48.0005
R8509 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t10 48.0005
R8510 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 45.5227
R8511 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 45.5227
R8512 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 45.5227
R8513 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 45.5227
R8514 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 6.39633
R8515 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 6.39633
R8516 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 6.39633
R8517 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 6.10467
R8518 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 6.10467
R8519 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 5.97967
R8520 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 5.91717
R8521 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 5.91717
R8522 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 5.14633
R8523 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 4.85467
R8524 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 4.72967
R8525 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 4.72967
R8526 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 4.66717
R8527 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 1.2505
R8528 a_7460_6300.n2 a_7460_6300.n1 594.301
R8529 a_7460_6300.n5 a_7460_6300.n4 594.301
R8530 a_7460_6300.n26 a_7460_6300.n25 594.301
R8531 a_7460_6300.n29 a_7460_6300.n28 594.301
R8532 a_7460_6300.n8 a_7460_6300.n7 594.301
R8533 a_7460_6300.n10 a_7460_6300.n9 594.301
R8534 a_7460_6300.n14 a_7460_6300.n13 594.301
R8535 a_7460_6300.n16 a_7460_6300.n15 594.301
R8536 a_7460_6300.n20 a_7460_6300.n19 594.301
R8537 a_7460_6300.n33 a_7460_6300.n32 594.301
R8538 a_7460_6300.n1 a_7460_6300.t4 78.8005
R8539 a_7460_6300.n1 a_7460_6300.t7 78.8005
R8540 a_7460_6300.n4 a_7460_6300.t1 78.8005
R8541 a_7460_6300.n4 a_7460_6300.t5 78.8005
R8542 a_7460_6300.n25 a_7460_6300.t6 78.8005
R8543 a_7460_6300.n25 a_7460_6300.t2 78.8005
R8544 a_7460_6300.n28 a_7460_6300.t9 78.8005
R8545 a_7460_6300.n28 a_7460_6300.t3 78.8005
R8546 a_7460_6300.n7 a_7460_6300.t14 78.8005
R8547 a_7460_6300.n7 a_7460_6300.t12 78.8005
R8548 a_7460_6300.n9 a_7460_6300.t19 78.8005
R8549 a_7460_6300.n9 a_7460_6300.t17 78.8005
R8550 a_7460_6300.n13 a_7460_6300.t11 78.8005
R8551 a_7460_6300.n13 a_7460_6300.t15 78.8005
R8552 a_7460_6300.n15 a_7460_6300.t13 78.8005
R8553 a_7460_6300.n15 a_7460_6300.t18 78.8005
R8554 a_7460_6300.n19 a_7460_6300.t0 78.8005
R8555 a_7460_6300.n19 a_7460_6300.t16 78.8005
R8556 a_7460_6300.t10 a_7460_6300.n33 78.8005
R8557 a_7460_6300.n33 a_7460_6300.t8 78.8005
R8558 a_7460_6300.n6 a_7460_6300.n2 6.20883
R8559 a_7460_6300.n27 a_7460_6300.n26 5.91717
R8560 a_7460_6300.n3 a_7460_6300.n2 5.91717
R8561 a_7460_6300.n30 a_7460_6300.n24 5.7505
R8562 a_7460_6300.n14 a_7460_6300.n11 5.41717
R8563 a_7460_6300.n22 a_7460_6300.n10 5.41717
R8564 a_7460_6300.n17 a_7460_6300.n14 5.22967
R8565 a_7460_6300.n12 a_7460_6300.n10 5.22967
R8566 a_7460_6300.n6 a_7460_6300.n5 4.95883
R8567 a_7460_6300.n30 a_7460_6300.n29 4.95883
R8568 a_7460_6300.n32 a_7460_6300.n31 4.95883
R8569 a_7460_6300.n16 a_7460_6300.n11 4.85467
R8570 a_7460_6300.n21 a_7460_6300.n20 4.85467
R8571 a_7460_6300.n5 a_7460_6300.n3 4.66717
R8572 a_7460_6300.n32 a_7460_6300.n0 4.66717
R8573 a_7460_6300.n29 a_7460_6300.n27 4.66717
R8574 a_7460_6300.n17 a_7460_6300.n16 4.66717
R8575 a_7460_6300.n20 a_7460_6300.n18 4.66717
R8576 a_7460_6300.n12 a_7460_6300.n8 4.66717
R8577 a_7460_6300.n23 a_7460_6300.n22 4.5005
R8578 a_7460_6300.n31 a_7460_6300.n30 1.2505
R8579 a_7460_6300.n27 a_7460_6300.n0 1.2505
R8580 a_7460_6300.n3 a_7460_6300.n0 1.2505
R8581 a_7460_6300.n31 a_7460_6300.n6 1.2505
R8582 a_7460_6300.n18 a_7460_6300.n12 0.563
R8583 a_7460_6300.n18 a_7460_6300.n17 0.563
R8584 a_7460_6300.n21 a_7460_6300.n11 0.563
R8585 a_7460_6300.n22 a_7460_6300.n21 0.563
R8586 a_7460_6300.n24 a_7460_6300.n23 0.51925
R8587 a_7460_6300.n26 a_7460_6300.n24 0.446333
R8588 a_7460_6300.n23 a_7460_6300.n8 0.354667
R8589 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 128.724
R8590 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 118.861
R8591 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 118.861
R8592 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 118.861
R8593 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 118.861
R8594 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 118.861
R8595 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t2 19.7005
R8596 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t6 19.7005
R8597 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t1 19.7005
R8598 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t9 19.7005
R8599 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t4 19.7005
R8600 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t8 19.7005
R8601 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t3 19.7005
R8602 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t7 19.7005
R8603 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t10 19.7005
R8604 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t5 19.7005
R8605 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 5.60467
R8606 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 5.54217
R8607 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 5.54217
R8608 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 5.04217
R8609 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 5.04217
R8610 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 5.04217
R8611 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 5.04217
R8612 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 4.97967
R8613 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 4.97967
R8614 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 4.97967
R8615 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 0.563
R8616 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 0.563
R8617 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 0.563
R8618 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 0.563
R8619 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 0.563
R8620 VIN-.n0 VIN-.t9 1000.38
R8621 VIN- VIN-.n9 433.019
R8622 VIN-.n9 VIN-.t1 273.134
R8623 VIN-.n0 VIN-.t0 273.134
R8624 VIN-.n1 VIN-.t5 273.134
R8625 VIN-.n2 VIN-.t10 273.134
R8626 VIN-.n3 VIN-.t3 273.134
R8627 VIN-.n4 VIN-.t7 273.134
R8628 VIN-.n5 VIN-.t4 273.134
R8629 VIN-.n6 VIN-.t8 273.134
R8630 VIN-.n7 VIN-.t2 273.134
R8631 VIN-.n8 VIN-.t6 273.134
R8632 VIN-.n9 VIN-.n8 176.733
R8633 VIN-.n8 VIN-.n7 176.733
R8634 VIN-.n7 VIN-.n6 176.733
R8635 VIN-.n6 VIN-.n5 176.733
R8636 VIN-.n5 VIN-.n4 176.733
R8637 VIN-.n4 VIN-.n3 176.733
R8638 VIN-.n3 VIN-.n2 176.733
R8639 VIN-.n2 VIN-.n1 176.733
R8640 VIN-.n1 VIN-.n0 176.733
R8641 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 120.817
R8642 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 107.121
R8643 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 97.4332
R8644 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 70.8161
R8645 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 24.288
R8646 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 24.288
R8647 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 24.288
R8648 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 24.288
R8649 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 24.288
R8650 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t3 24.0005
R8651 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t14 24.0005
R8652 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t1 24.0005
R8653 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t2 24.0005
R8654 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t5 8.0005
R8655 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t9 8.0005
R8656 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t4 8.0005
R8657 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t11 8.0005
R8658 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t6 8.0005
R8659 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t10 8.0005
R8660 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t7 8.0005
R8661 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t12 8.0005
R8662 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t8 8.0005
R8663 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t13 8.0005
R8664 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 5.96925
R8665 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 5.7505
R8666 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 5.7505
R8667 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 5.7505
R8668 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 5.188
R8669 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 5.188
R8670 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 5.188
R8671 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 5.188
R8672 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 5.188
R8673 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 5.188
R8674 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 5.188
R8675 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 0.563
R8676 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 0.563
R8677 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 0.563
R8678 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 0.563
R8679 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 0.563
R8680 VIN+.n0 VIN+.t3 1001.28
R8681 VIN+ VIN+.n9 433.019
R8682 VIN+.n9 VIN+.t9 273.134
R8683 VIN+.n0 VIN+.t0 273.134
R8684 VIN+.n8 VIN+.t5 273.134
R8685 VIN+.n7 VIN+.t8 273.134
R8686 VIN+.n6 VIN+.t4 273.134
R8687 VIN+.n5 VIN+.t7 273.134
R8688 VIN+.n4 VIN+.t1 273.134
R8689 VIN+.n3 VIN+.t10 273.134
R8690 VIN+.n2 VIN+.t2 273.134
R8691 VIN+.n1 VIN+.t6 273.134
R8692 VIN+.n1 VIN+.n0 176.733
R8693 VIN+.n2 VIN+.n1 176.733
R8694 VIN+.n3 VIN+.n2 176.733
R8695 VIN+.n4 VIN+.n3 176.733
R8696 VIN+.n5 VIN+.n4 176.733
R8697 VIN+.n6 VIN+.n5 176.733
R8698 VIN+.n7 VIN+.n6 176.733
R8699 VIN+.n8 VIN+.n7 176.733
R8700 VIN+.n9 VIN+.n8 176.733
R8701 w_7200_15600.t45 w_7200_15600.n3 698.638
R8702 w_7200_15600.t45 w_7200_15600.n52 694.444
R8703 w_7200_15600.t44 w_7200_15600.n3 674.87
R8704 w_7200_15600.n4 w_7200_15600.t38 643.038
R8705 w_7200_15600.n31 w_7200_15600.n20 587.407
R8706 w_7200_15600.n27 w_7200_15600.n26 587.407
R8707 w_7200_15600.n43 w_7200_15600.n42 587.407
R8708 w_7200_15600.n44 w_7200_15600.n15 587.407
R8709 w_7200_15600.n43 w_7200_15600.n36 585
R8710 w_7200_15600.n45 w_7200_15600.n44 585
R8711 w_7200_15600.n29 w_7200_15600.n20 585
R8712 w_7200_15600.n28 w_7200_15600.n27 585
R8713 w_7200_15600.n51 w_7200_15600.t43 413.084
R8714 w_7200_15600.n5 w_7200_15600.t37 413.084
R8715 w_7200_15600.t38 w_7200_15600.t32 373.214
R8716 w_7200_15600.t32 w_7200_15600.t33 373.214
R8717 w_7200_15600.t33 w_7200_15600.t44 373.214
R8718 w_7200_15600.n6 w_7200_15600.t34 360.868
R8719 w_7200_15600.n50 w_7200_15600.t40 360.868
R8720 w_7200_15600.n4 w_7200_15600.t39 354.063
R8721 w_7200_15600.t14 w_7200_15600.t35 251.471
R8722 w_7200_15600.t10 w_7200_15600.t14 251.471
R8723 w_7200_15600.t28 w_7200_15600.t10 251.471
R8724 w_7200_15600.t2 w_7200_15600.t28 251.471
R8725 w_7200_15600.t12 w_7200_15600.t2 251.471
R8726 w_7200_15600.t22 w_7200_15600.t12 251.471
R8727 w_7200_15600.t20 w_7200_15600.t22 251.471
R8728 w_7200_15600.t0 w_7200_15600.t20 251.471
R8729 w_7200_15600.t6 w_7200_15600.t0 251.471
R8730 w_7200_15600.t16 w_7200_15600.t6 251.471
R8731 w_7200_15600.t26 w_7200_15600.t16 251.471
R8732 w_7200_15600.t24 w_7200_15600.t26 251.471
R8733 w_7200_15600.t4 w_7200_15600.t24 251.471
R8734 w_7200_15600.t8 w_7200_15600.t4 251.471
R8735 w_7200_15600.t18 w_7200_15600.t8 251.471
R8736 w_7200_15600.t30 w_7200_15600.t18 251.471
R8737 w_7200_15600.t41 w_7200_15600.t30 251.471
R8738 w_7200_15600.n42 w_7200_15600.n37 243.698
R8739 w_7200_15600.n49 w_7200_15600.n48 238.367
R8740 w_7200_15600.t35 w_7200_15600.n33 237.5
R8741 w_7200_15600.n34 w_7200_15600.t41 237.5
R8742 w_7200_15600.n32 w_7200_15600.n31 190.333
R8743 w_7200_15600.n41 w_7200_15600.n40 185
R8744 w_7200_15600.n39 w_7200_15600.n36 185
R8745 w_7200_15600.n45 w_7200_15600.n35 185
R8746 w_7200_15600.n47 w_7200_15600.n46 185
R8747 w_7200_15600.n33 w_7200_15600.n32 185
R8748 w_7200_15600.n30 w_7200_15600.n19 185
R8749 w_7200_15600.n29 w_7200_15600.n21 185
R8750 w_7200_15600.n28 w_7200_15600.n22 185
R8751 w_7200_15600.n24 w_7200_15600.n23 185
R8752 w_7200_15600.n25 w_7200_15600.n18 185
R8753 w_7200_15600.n33 w_7200_15600.n18 185
R8754 w_7200_15600.n0 w_7200_15600.n14 165.505
R8755 w_7200_15600.n0 w_7200_15600.n13 165.505
R8756 w_7200_15600.n0 w_7200_15600.n12 165.505
R8757 w_7200_15600.n0 w_7200_15600.n11 165.505
R8758 w_7200_15600.n1 w_7200_15600.n10 165.505
R8759 w_7200_15600.n1 w_7200_15600.n9 165.505
R8760 w_7200_15600.n1 w_7200_15600.n8 165.505
R8761 w_7200_15600.n1 w_7200_15600.n7 165.505
R8762 w_7200_15600.n40 w_7200_15600.n39 150
R8763 w_7200_15600.n47 w_7200_15600.n35 150
R8764 w_7200_15600.n32 w_7200_15600.n19 150
R8765 w_7200_15600.n22 w_7200_15600.n21 150
R8766 w_7200_15600.n23 w_7200_15600.n18 150
R8767 w_7200_15600.t36 w_7200_15600.n20 123.126
R8768 w_7200_15600.n27 w_7200_15600.t36 123.126
R8769 w_7200_15600.t42 w_7200_15600.n43 123.126
R8770 w_7200_15600.n44 w_7200_15600.t42 123.126
R8771 w_7200_15600.n37 w_7200_15600.n34 65.8183
R8772 w_7200_15600.n38 w_7200_15600.n34 65.8183
R8773 w_7200_15600.n48 w_7200_15600.n34 65.8183
R8774 w_7200_15600.n33 w_7200_15600.n16 65.8183
R8775 w_7200_15600.n33 w_7200_15600.n17 65.8183
R8776 w_7200_15600.n40 w_7200_15600.n37 53.3664
R8777 w_7200_15600.n39 w_7200_15600.n38 53.3664
R8778 w_7200_15600.n48 w_7200_15600.n47 53.3664
R8779 w_7200_15600.n38 w_7200_15600.n35 53.3664
R8780 w_7200_15600.n19 w_7200_15600.n16 53.3664
R8781 w_7200_15600.n22 w_7200_15600.n17 53.3664
R8782 w_7200_15600.n21 w_7200_15600.n16 53.3664
R8783 w_7200_15600.n23 w_7200_15600.n17 53.3664
R8784 w_7200_15600.n5 w_7200_15600.n4 22.9536
R8785 w_7200_15600.n50 w_7200_15600.n49 22.8576
R8786 w_7200_15600.n25 w_7200_15600.n6 22.8576
R8787 w_7200_15600.n52 w_7200_15600.n51 18.3472
R8788 w_7200_15600.n14 w_7200_15600.t19 13.1338
R8789 w_7200_15600.n14 w_7200_15600.t31 13.1338
R8790 w_7200_15600.n13 w_7200_15600.t5 13.1338
R8791 w_7200_15600.n13 w_7200_15600.t9 13.1338
R8792 w_7200_15600.n12 w_7200_15600.t27 13.1338
R8793 w_7200_15600.n12 w_7200_15600.t25 13.1338
R8794 w_7200_15600.n11 w_7200_15600.t7 13.1338
R8795 w_7200_15600.n11 w_7200_15600.t17 13.1338
R8796 w_7200_15600.n10 w_7200_15600.t21 13.1338
R8797 w_7200_15600.n10 w_7200_15600.t1 13.1338
R8798 w_7200_15600.n9 w_7200_15600.t13 13.1338
R8799 w_7200_15600.n9 w_7200_15600.t23 13.1338
R8800 w_7200_15600.n8 w_7200_15600.t29 13.1338
R8801 w_7200_15600.n8 w_7200_15600.t3 13.1338
R8802 w_7200_15600.n7 w_7200_15600.t15 13.1338
R8803 w_7200_15600.n7 w_7200_15600.t11 13.1338
R8804 w_7200_15600.n2 w_7200_15600.n5 11.5991
R8805 w_7200_15600.n51 w_7200_15600.n2 11.3696
R8806 w_7200_15600.n0 w_7200_15600.n50 11.0575
R8807 w_7200_15600.n2 w_7200_15600.n6 10.87
R8808 w_7200_15600.n41 w_7200_15600.n36 9.14336
R8809 w_7200_15600.n45 w_7200_15600.n36 9.14336
R8810 w_7200_15600.n46 w_7200_15600.n45 9.14336
R8811 w_7200_15600.n30 w_7200_15600.n29 9.14336
R8812 w_7200_15600.n29 w_7200_15600.n28 9.14336
R8813 w_7200_15600.n28 w_7200_15600.n24 9.14336
R8814 w_7200_15600.n49 w_7200_15600.n15 5.33286
R8815 w_7200_15600.n26 w_7200_15600.n25 5.33286
R8816 w_7200_15600.n52 w_7200_15600.n3 4.19264
R8817 w_7200_15600.n42 w_7200_15600.n41 3.75335
R8818 w_7200_15600.n46 w_7200_15600.n15 3.75335
R8819 w_7200_15600.n31 w_7200_15600.n30 3.75335
R8820 w_7200_15600.n26 w_7200_15600.n24 3.75335
R8821 w_7200_15600.n1 w_7200_15600.n0 1.1255
R8822 w_7200_15600.n2 w_7200_15600.n1 0.703625
R8823 a_12070_24908.t0 a_12070_24908.t1 178.133
R8824 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t3 661.375
R8825 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t0 661.375
R8826 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n6 213.131
R8827 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t4 213.131
R8828 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t1 146.155
R8829 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t9 146.155
R8830 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t2 76.2576
R8831 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n7 76.2576
R8832 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n1 72.4424
R8833 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n2 66.4532
R8834 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t10 11.2576
R8835 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t5 11.2576
R8836 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t7 11.2576
R8837 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t8 11.2576
R8838 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n4 5.1255
R8839 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n3 4.9096
R8840 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n0 4.7505
R8841 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n5 1.888
R8842 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n0 1.888
R8843 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R8844 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R8845 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 175.623
R8846 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 169
R8847 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 166.988
R8848 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t1 130.001
R8849 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t0 81.7074
R8850 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.8552
R8851 bgr_11_0.START_UP bgr_11_0.START_UP.n5 15.4067
R8852 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t2 13.1338
R8853 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t4 13.1338
R8854 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t3 13.1338
R8855 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t5 13.1338
R8856 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R8857 a_5700_24908.t0 a_5700_24908.t1 178.133
R8858 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 528.612
R8859 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n1 169.56
R8860 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 168.435
R8861 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t0 148.653
R8862 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t1 125.418
R8863 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n0 17.871
R8864 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t2 13.1338
R8865 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t5 13.1338
R8866 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t4 13.1338
R8867 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t3 13.1338
R8868 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 11.8755
R8869 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 5.54738
R8870 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.n15 325.473
R8871 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.n8 325.473
R8872 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.n3 325.473
R8873 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t17 310.488
R8874 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t18 310.488
R8875 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t13 310.488
R8876 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.t10 184.097
R8877 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.t8 184.097
R8878 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.t6 184.097
R8879 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.n12 167.094
R8880 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.n5 167.094
R8881 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.n0 167.094
R8882 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.n7 152
R8883 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.n2 152
R8884 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n14 152
R8885 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t14 120.501
R8886 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.t2 120.501
R8887 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t16 120.501
R8888 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.t4 120.501
R8889 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t15 120.501
R8890 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.t0 120.501
R8891 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.t12 106.933
R8892 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.n13 40.7027
R8893 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.n6 40.7027
R8894 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.n1 40.7027
R8895 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.t5 39.4005
R8896 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.t9 39.4005
R8897 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.t1 39.4005
R8898 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.t7 39.4005
R8899 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.t3 39.4005
R8900 bgr_11_0.V_mir2.t11 bgr_11_0.V_mir2.n16 39.4005
R8901 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n4 15.9255
R8902 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n11 15.9255
R8903 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.n9 9.3005
R8904 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n10 4.5005
R8905 bgr_11_0.Vin- bgr_11_0.Vin-.t8 531.89
R8906 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 351.522
R8907 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n10 170.904
R8908 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n11 168.654
R8909 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.t2 115.442
R8910 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.n2 83.5719
R8911 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n4 83.5719
R8912 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n1 73.8495
R8913 bgr_11_0.Vin-.t3 bgr_11_0.Vin-.n0 65.0341
R8914 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.t1 39.4005
R8915 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.t0 39.4005
R8916 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n3 26.074
R8917 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 20.7036
R8918 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.t7 13.1338
R8919 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.t4 13.1338
R8920 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t5 13.1338
R8921 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t6 13.1338
R8922 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n9 11.4067
R8923 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 8.313
R8924 bgr_11_0.Vin- bgr_11_0.Vin-.n15 5.70362
R8925 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n12 2.0005
R8926 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.n0 1.56483
R8927 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 1.5505
R8928 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n5 0.885803
R8929 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n2 0.77514
R8930 bgr_11_0.Vin-.n5 bgr_11_0.Vin- 0.756696
R8931 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n1 0.711459
R8932 bgr_11_0.Vin- bgr_11_0.Vin-.n1 0.576566
R8933 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n0 0.531499
R8934 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t3 0.290206
R8935 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 0.00817857
R8936 two_stage_opamp_dummy_magic_23_0.V_p_mir.n1 two_stage_opamp_dummy_magic_23_0.V_p_mir.n0 97.1193
R8937 two_stage_opamp_dummy_magic_23_0.V_p_mir.n0 two_stage_opamp_dummy_magic_23_0.V_p_mir.t1 16.0005
R8938 two_stage_opamp_dummy_magic_23_0.V_p_mir.n0 two_stage_opamp_dummy_magic_23_0.V_p_mir.t0 16.0005
R8939 two_stage_opamp_dummy_magic_23_0.V_p_mir.t2 two_stage_opamp_dummy_magic_23_0.V_p_mir.n1 9.6005
R8940 two_stage_opamp_dummy_magic_23_0.V_p_mir.n1 two_stage_opamp_dummy_magic_23_0.V_p_mir.t3 9.6005
R8941 a_6350_25058.t0 a_6350_25058.t1 178.133
R8942 a_8260_1600.n1 a_8260_1600.t4 65.3505
R8943 a_8260_1600.n3 a_8260_1600.n2 49.3505
R8944 a_8260_1600.n6 a_8260_1600.n5 49.3505
R8945 a_8260_1600.n2 a_8260_1600.t0 16.0005
R8946 a_8260_1600.n2 a_8260_1600.t2 16.0005
R8947 a_8260_1600.n6 a_8260_1600.t1 16.0005
R8948 a_8260_1600.t3 a_8260_1600.n6 16.0005
R8949 a_8260_1600.n1 a_8260_1600.n0 6.3755
R8950 a_8260_1600.n4 a_8260_1600.n1 6.1255
R8951 a_8260_1600.n3 a_8260_1600.n0 5.688
R8952 a_8260_1600.n4 a_8260_1600.n3 5.438
R8953 a_8260_1600.n5 a_8260_1600.n0 5.1255
R8954 a_8260_1600.n5 a_8260_1600.n4 4.8755
R8955 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 172.969
R8956 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R8957 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R8958 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R8959 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R8960 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R8961 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R8962 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R8963 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R8964 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R8965 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R8966 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R8967 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R8968 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R8969 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R8970 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R8971 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R8972 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R8973 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R8974 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R8975 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R8976 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R8977 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R8978 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R8979 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R8980 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R8981 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R8982 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R8983 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R8984 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R8985 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R8986 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R8987 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R8988 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R8989 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R8990 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R8991 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R8992 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 65.0299
R8993 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R8994 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R8995 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R8996 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R8997 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R8998 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R8999 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R9000 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R9001 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R9002 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R9003 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R9004 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R9005 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R9006 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R9007 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R9008 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R9009 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9010 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9011 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R9012 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9013 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9014 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9015 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R9016 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9017 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9018 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9019 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9020 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R9021 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R9022 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9023 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9024 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9025 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R9026 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9027 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9028 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9029 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R9030 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9031 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9032 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9033 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R9034 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R9035 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R9036 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9037 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9038 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9039 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R9040 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9041 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9042 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9043 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R9044 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9045 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9046 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9047 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9048 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9049 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9050 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9051 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9052 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9053 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9054 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9055 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9056 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R9057 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R9058 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9059 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9060 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9061 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9062 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R9063 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R9064 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R9065 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R9066 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R9067 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R9068 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R9069 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R9070 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R9071 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R9072 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R9073 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R9074 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R9075 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R9076 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R9077 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R9078 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R9079 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R9080 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R9081 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R9082 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R9083 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R9084 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R9085 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R9086 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R9087 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R9088 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R9089 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R9090 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R9091 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R9092 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R9093 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R9094 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R9095 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R9096 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R9097 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R9098 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R9099 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R9100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R9101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R9102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R9103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R9104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R9105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R9106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R9107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R9108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R9109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R9110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R9111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R9112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R9113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R9114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R9115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R9116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R9117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R9118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R9119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R9120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R9121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R9122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R9123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R9124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R9125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R9126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R9127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R9128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R9129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R9130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R9131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R9132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R9133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R9134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R9135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R9136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R9137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R9138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R9139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R9140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R9141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R9142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R9143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R9144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R9145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R9146 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R9147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R9148 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R9149 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R9150 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R9151 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R9152 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R9153 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R9154 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R9155 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R9156 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R9157 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R9158 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R9159 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R9160 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R9161 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R9162 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R9163 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R9164 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R9165 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R9166 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R9167 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R9168 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R9169 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R9170 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R9171 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9172 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9173 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9174 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R9175 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9176 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R9177 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R9178 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R9179 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R9180 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R9181 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R9182 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R9183 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R9184 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R9185 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R9186 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R9187 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R9188 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R9189 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R9190 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R9191 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R9192 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R9193 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R9194 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R9195 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R9196 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R9197 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R9198 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R9199 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R9200 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R9201 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R9202 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R9203 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R9204 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R9205 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R9206 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R9207 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R9208 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R9209 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R9210 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R9211 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R9212 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R9213 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R9214 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R9215 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R9216 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R9217 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R9218 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R9219 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R9220 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R9221 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R9222 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R9223 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R9224 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R9225 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R9226 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R9227 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R9228 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R9229 bgr_11_0.V_CMFB_S3.n2 bgr_11_0.V_CMFB_S3.n0 345.264
R9230 bgr_11_0.V_CMFB_S3.n3 bgr_11_0.V_CMFB_S3.n2 345.264
R9231 bgr_11_0.V_CMFB_S3.n2 bgr_11_0.V_CMFB_S3.n1 344.7
R9232 bgr_11_0.V_CMFB_S3.n1 bgr_11_0.V_CMFB_S3.t5 39.4005
R9233 bgr_11_0.V_CMFB_S3.n1 bgr_11_0.V_CMFB_S3.t2 39.4005
R9234 bgr_11_0.V_CMFB_S3.n0 bgr_11_0.V_CMFB_S3.t3 39.4005
R9235 bgr_11_0.V_CMFB_S3.n0 bgr_11_0.V_CMFB_S3.t1 39.4005
R9236 bgr_11_0.V_CMFB_S3.n3 bgr_11_0.V_CMFB_S3.t0 39.4005
R9237 bgr_11_0.V_CMFB_S3.t4 bgr_11_0.V_CMFB_S3.n3 39.4005
R9238 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R9239 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t8 525.38
R9240 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t3 525.38
R9241 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t5 483.608
R9242 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t6 360.43
R9243 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t2 291.209
R9244 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t4 281.168
R9245 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t9 281.168
R9246 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t7 281.168
R9247 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 244.214
R9248 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 202.44
R9249 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 202.159
R9250 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 165.972
R9251 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 117.754
R9252 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t1 117.254
R9253 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 79.2627
R9254 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 18.9067
R9255 a_4200_4468.t0 a_4200_4468.t1 169.905
R9256 two_stage_opamp_dummy_magic_23_0.V_tot.n6 two_stage_opamp_dummy_magic_23_0.V_tot.n5 771.76
R9257 two_stage_opamp_dummy_magic_23_0.V_tot.n11 two_stage_opamp_dummy_magic_23_0.V_tot.n10 595.444
R9258 two_stage_opamp_dummy_magic_23_0.V_tot.n1 two_stage_opamp_dummy_magic_23_0.V_tot.n0 595.131
R9259 two_stage_opamp_dummy_magic_23_0.V_tot.n3 two_stage_opamp_dummy_magic_23_0.V_tot.n2 530.201
R9260 two_stage_opamp_dummy_magic_23_0.V_tot.n5 two_stage_opamp_dummy_magic_23_0.V_tot.n4 530.201
R9261 two_stage_opamp_dummy_magic_23_0.V_tot.n7 two_stage_opamp_dummy_magic_23_0.V_tot.n6 530.201
R9262 two_stage_opamp_dummy_magic_23_0.V_tot.n9 two_stage_opamp_dummy_magic_23_0.V_tot.n8 530.201
R9263 two_stage_opamp_dummy_magic_23_0.V_tot.n5 two_stage_opamp_dummy_magic_23_0.V_tot.t8 208.868
R9264 two_stage_opamp_dummy_magic_23_0.V_tot.n4 two_stage_opamp_dummy_magic_23_0.V_tot.t13 208.868
R9265 two_stage_opamp_dummy_magic_23_0.V_tot.n3 two_stage_opamp_dummy_magic_23_0.V_tot.t6 208.868
R9266 two_stage_opamp_dummy_magic_23_0.V_tot.n2 two_stage_opamp_dummy_magic_23_0.V_tot.t12 208.868
R9267 two_stage_opamp_dummy_magic_23_0.V_tot.n1 two_stage_opamp_dummy_magic_23_0.V_tot.t5 208.868
R9268 two_stage_opamp_dummy_magic_23_0.V_tot.n10 two_stage_opamp_dummy_magic_23_0.V_tot.t11 208.868
R9269 two_stage_opamp_dummy_magic_23_0.V_tot.n9 two_stage_opamp_dummy_magic_23_0.V_tot.t4 208.868
R9270 two_stage_opamp_dummy_magic_23_0.V_tot.n8 two_stage_opamp_dummy_magic_23_0.V_tot.t10 208.868
R9271 two_stage_opamp_dummy_magic_23_0.V_tot.n7 two_stage_opamp_dummy_magic_23_0.V_tot.t7 208.868
R9272 two_stage_opamp_dummy_magic_23_0.V_tot.n6 two_stage_opamp_dummy_magic_23_0.V_tot.t9 208.868
R9273 two_stage_opamp_dummy_magic_23_0.V_tot.n2 two_stage_opamp_dummy_magic_23_0.V_tot.n1 176.733
R9274 two_stage_opamp_dummy_magic_23_0.V_tot.n4 two_stage_opamp_dummy_magic_23_0.V_tot.n3 176.733
R9275 two_stage_opamp_dummy_magic_23_0.V_tot.n8 two_stage_opamp_dummy_magic_23_0.V_tot.n7 176.733
R9276 two_stage_opamp_dummy_magic_23_0.V_tot.n10 two_stage_opamp_dummy_magic_23_0.V_tot.n9 176.733
R9277 two_stage_opamp_dummy_magic_23_0.V_tot.n0 two_stage_opamp_dummy_magic_23_0.V_tot.t2 117.591
R9278 two_stage_opamp_dummy_magic_23_0.V_tot.t0 two_stage_opamp_dummy_magic_23_0.V_tot.n11 117.591
R9279 two_stage_opamp_dummy_magic_23_0.V_tot.n11 two_stage_opamp_dummy_magic_23_0.V_tot.t3 108.424
R9280 two_stage_opamp_dummy_magic_23_0.V_tot.n0 two_stage_opamp_dummy_magic_23_0.V_tot.t1 108.424
R9281 bgr_11_0.V_CMFB_S1.n2 bgr_11_0.V_CMFB_S1.n0 344.837
R9282 bgr_11_0.V_CMFB_S1.n3 bgr_11_0.V_CMFB_S1.n2 344.837
R9283 bgr_11_0.V_CMFB_S1.n2 bgr_11_0.V_CMFB_S1.n1 344.274
R9284 bgr_11_0.V_CMFB_S1.n1 bgr_11_0.V_CMFB_S1.t1 39.4005
R9285 bgr_11_0.V_CMFB_S1.n1 bgr_11_0.V_CMFB_S1.t5 39.4005
R9286 bgr_11_0.V_CMFB_S1.n0 bgr_11_0.V_CMFB_S1.t3 39.4005
R9287 bgr_11_0.V_CMFB_S1.n0 bgr_11_0.V_CMFB_S1.t0 39.4005
R9288 bgr_11_0.V_CMFB_S1.n3 bgr_11_0.V_CMFB_S1.t2 39.4005
R9289 bgr_11_0.V_CMFB_S1.t4 bgr_11_0.V_CMFB_S1.n3 39.4005
R9290 a_11420_25058.t0 a_11420_25058.t1 178.133
R9291 a_11950_23700.t0 a_11950_23700.t1 178.133
R9292 a_4600_1446.t0 a_4600_1446.t1 169.905
R9293 a_4080_4468.t0 a_4080_4468.t1 294.339
R9294 a_13130_1456.t0 a_13130_1456.t1 169.905
R9295 a_11300_23450.t0 a_11300_23450.t1 178.133
R9296 a_13450_4368.t0 a_13450_4368.t1 294.339
R9297 a_13570_4368.t0 a_13570_4368.t1 169.905
C0 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.Vin- 1.06389f
C1 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_tail_gate 1.43091f
C2 a_6520_18930# bgr_11_0.1st_Vout_1 0.067812f
C3 two_stage_opamp_dummy_magic_23_0.V_err_gate VDDA 2.4373f
C4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref bgr_11_0.Vin+ 0.303835f
C5 VIN+ VIN- 0.151796f
C6 bgr_11_0.START_UP VDDA 0.893209f
C7 VIN+ two_stage_opamp_dummy_magic_23_0.VD2 0.510937f
C8 VDDA bgr_11_0.Vin- 1.17623f
C9 two_stage_opamp_dummy_magic_23_0.X two_stage_opamp_dummy_magic_23_0.err_amp_out 0.20522f
C10 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.01235f
C11 two_stage_opamp_dummy_magic_23_0.V_tail_gate VOUT+ 0.010408f
C12 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.289292f
C13 bgr_11_0.1st_Vout_1 VDDA 3.19163f
C14 VDDA VOUT+ 13.4377f
C15 VDDA two_stage_opamp_dummy_magic_23_0.VD4 8.479321f
C16 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.cap_res_Y 0.03128f
C17 two_stage_opamp_dummy_magic_23_0.cap_res_Y VDDA 0.533063f
C18 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.X 0.18001f
C19 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.START_UP 0.751706f
C20 two_stage_opamp_dummy_magic_23_0.V_tail_gate VOUT- 0.02527f
C21 two_stage_opamp_dummy_magic_23_0.X VDDA 5.01789f
C22 a_6520_18930# bgr_11_0.Vin+ 0.037147f
C23 VDDA VOUT- 13.403299f
C24 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.Vin- 0.285566f
C25 VDDA two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 4.79436f
C26 bgr_11_0.START_UP_NFET1 a_6520_18930# 0.203967f
C27 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.24593f
C28 two_stage_opamp_dummy_magic_23_0.V_tail_gate VIN+ 0.056847f
C29 bgr_11_0.START_UP bgr_11_0.Vin- 3.75854f
C30 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.1st_Vout_1 0.043095f
C31 two_stage_opamp_dummy_magic_23_0.V_tail_gate VIN- 0.135101f
C32 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.042777f
C33 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.X 0.161254f
C34 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.VD2 0.02379f
C35 two_stage_opamp_dummy_magic_23_0.V_err_gate VOUT- 0.038404f
C36 VDDA bgr_11_0.Vin+ 1.80899f
C37 VDDA two_stage_opamp_dummy_magic_23_0.VD2 0.027746f
C38 bgr_11_0.1st_Vout_1 bgr_11_0.Vin- 0.85607f
C39 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.492517f
C40 bgr_11_0.START_UP_NFET1 VDDA 0.010695f
C41 bgr_11_0.START_UP two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 1.37084f
C42 a_6520_18930# VDDA 1.51775f
C43 VOUT+ two_stage_opamp_dummy_magic_23_0.VD4 0.028865f
C44 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref bgr_11_0.Vin- 0.126816f
C45 VDDA bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.112096f
C46 two_stage_opamp_dummy_magic_23_0.cap_res_Y VOUT+ 50.8462f
C47 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.err_amp_out 0.343731f
C48 two_stage_opamp_dummy_magic_23_0.cap_res_Y two_stage_opamp_dummy_magic_23_0.VD4 0.054393f
C49 two_stage_opamp_dummy_magic_23_0.err_amp_out VDDA 1.0994f
C50 VOUT+ VOUT- 0.305434f
C51 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.Vin+ 0.097188f
C52 VOUT+ two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.039549f
C53 two_stage_opamp_dummy_magic_23_0.cap_res_Y VOUT- 0.028842f
C54 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.04352f
C55 bgr_11_0.START_UP bgr_11_0.Vin+ 0.315805f
C56 two_stage_opamp_dummy_magic_23_0.X VOUT- 2.33193f
C57 two_stage_opamp_dummy_magic_23_0.cap_res_Y two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.243261f
C58 two_stage_opamp_dummy_magic_23_0.V_tail_gate VDDA 7.06141f
C59 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C60 bgr_11_0.Vin+ bgr_11_0.Vin- 5.51003f
C61 bgr_11_0.START_UP a_6520_18930# 0.322861f
C62 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.err_amp_out 0.026461f
C63 bgr_11_0.1st_Vout_1 bgr_11_0.Vin+ 0.168603f
C64 a_6520_18930# bgr_11_0.Vin- 0.010578f
C65 VIN- GNDA 1.92317f
C66 VIN+ GNDA 1.90963f
C67 VOUT- GNDA 20.532288f
C68 VOUT+ GNDA 20.582405f
C69 VDDA GNDA 0.230761p
C70 two_stage_opamp_dummy_magic_23_0.VD2 GNDA 2.003606f
C71 two_stage_opamp_dummy_magic_23_0.err_amp_out GNDA 5.194764f
C72 two_stage_opamp_dummy_magic_23_0.cap_res_Y GNDA 33.372776f
C73 two_stage_opamp_dummy_magic_23_0.X GNDA 7.15177f
C74 two_stage_opamp_dummy_magic_23_0.V_tail_gate GNDA 10.119929f
C75 bgr_11_0.1st_Vout_1 GNDA 7.227168f
C76 a_6520_18930# GNDA 9.62462f
C77 bgr_11_0.START_UP GNDA 6.80373f
C78 bgr_11_0.START_UP_NFET1 GNDA 4.94893f
C79 two_stage_opamp_dummy_magic_23_0.V_err_gate GNDA 11.45712f
C80 bgr_11_0.Vin- GNDA 5.178825f
C81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.1884f
C82 bgr_11_0.Vin+ GNDA 4.851241f
C83 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref GNDA 8.26348f
C84 two_stage_opamp_dummy_magic_23_0.VD4 GNDA 5.12103f
C85 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t1 GNDA 0.124526f
C86 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t5 GNDA 0.365905f
C87 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t7 GNDA 0.313782f
C88 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t3 GNDA 0.37241f
C89 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 GNDA 0.195093f
C90 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t2 GNDA 0.317627f
C91 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 GNDA 0.210094f
C92 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 GNDA 0.585951f
C93 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t6 GNDA 0.340499f
C94 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t9 GNDA 0.313782f
C95 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t4 GNDA 0.313782f
C96 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t8 GNDA 0.37241f
C97 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 GNDA 0.196704f
C98 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 GNDA 0.124569f
C99 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 GNDA 0.118809f
C100 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 GNDA 0.608541f
C101 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t0 GNDA 0.125517f
C102 a_8260_1600.t1 GNDA 0.047649f
C103 a_8260_1600.n0 GNDA 0.318351f
C104 a_8260_1600.t4 GNDA 0.161927f
C105 a_8260_1600.n1 GNDA 0.491746f
C106 a_8260_1600.t0 GNDA 0.047649f
C107 a_8260_1600.t2 GNDA 0.047649f
C108 a_8260_1600.n2 GNDA 0.103679f
C109 a_8260_1600.n3 GNDA 0.42438f
C110 a_8260_1600.n4 GNDA 0.297965f
C111 a_8260_1600.n5 GNDA 0.407675f
C112 a_8260_1600.n6 GNDA 0.103679f
C113 a_8260_1600.t3 GNDA 0.047649f
C114 bgr_11_0.Vin-.n0 GNDA 0.593347f
C115 bgr_11_0.Vin-.n1 GNDA 0.450957f
C116 bgr_11_0.Vin-.n2 GNDA 0.150555f
C117 bgr_11_0.Vin-.t3 GNDA 0.329365f
C118 bgr_11_0.Vin-.n3 GNDA 0.087966f
C119 bgr_11_0.Vin-.n4 GNDA 0.397997f
C120 bgr_11_0.Vin-.n5 GNDA 0.087803f
C121 bgr_11_0.Vin-.n6 GNDA 0.08879f
C122 bgr_11_0.Vin-.n7 GNDA 0.728936f
C123 bgr_11_0.Vin-.n8 GNDA 1.56103f
C124 bgr_11_0.Vin-.t2 GNDA 0.149853f
C125 bgr_11_0.Vin-.n9 GNDA 1.3499f
C126 bgr_11_0.Vin-.t7 GNDA 0.034117f
C127 bgr_11_0.Vin-.t4 GNDA 0.034117f
C128 bgr_11_0.Vin-.n10 GNDA 0.117222f
C129 bgr_11_0.Vin-.t5 GNDA 0.034117f
C130 bgr_11_0.Vin-.t6 GNDA 0.034117f
C131 bgr_11_0.Vin-.n11 GNDA 0.113415f
C132 bgr_11_0.Vin-.n12 GNDA 0.710998f
C133 bgr_11_0.Vin-.t1 GNDA 0.011372f
C134 bgr_11_0.Vin-.t0 GNDA 0.011372f
C135 bgr_11_0.Vin-.n13 GNDA 0.034848f
C136 bgr_11_0.Vin-.n14 GNDA 0.652105f
C137 bgr_11_0.Vin-.n15 GNDA 0.994698f
C138 bgr_11_0.Vin-.t8 GNDA 0.052355f
C139 bgr_11_0.Vin+.t1 GNDA 0.249571f
C140 bgr_11_0.Vin+.t0 GNDA 0.108169f
C141 bgr_11_0.Vin+.n0 GNDA 1.7947f
C142 bgr_11_0.Vin+.t2 GNDA 0.037179f
C143 bgr_11_0.Vin+.t5 GNDA 0.037179f
C144 bgr_11_0.Vin+.n1 GNDA 0.124175f
C145 bgr_11_0.Vin+.t4 GNDA 0.037179f
C146 bgr_11_0.Vin+.t3 GNDA 0.037179f
C147 bgr_11_0.Vin+.n2 GNDA 0.122828f
C148 bgr_11_0.Vin+.n3 GNDA 1.00899f
C149 bgr_11_0.Vin+.n4 GNDA 1.45475f
C150 bgr_11_0.Vin+.t6 GNDA 0.05926f
C151 bgr_11_0.START_UP.t0 GNDA 1.24502f
C152 bgr_11_0.START_UP.t1 GNDA 0.032728f
C153 bgr_11_0.START_UP.n0 GNDA 0.833376f
C154 bgr_11_0.START_UP.t2 GNDA 0.031233f
C155 bgr_11_0.START_UP.t4 GNDA 0.031233f
C156 bgr_11_0.START_UP.n1 GNDA 0.113473f
C157 bgr_11_0.START_UP.t3 GNDA 0.031233f
C158 bgr_11_0.START_UP.t5 GNDA 0.031233f
C159 bgr_11_0.START_UP.n2 GNDA 0.10433f
C160 bgr_11_0.START_UP.n3 GNDA 0.543759f
C161 bgr_11_0.START_UP.t6 GNDA 0.011737f
C162 bgr_11_0.START_UP.t7 GNDA 0.011737f
C163 bgr_11_0.START_UP.n4 GNDA 0.033214f
C164 bgr_11_0.START_UP.n5 GNDA 0.333711f
C165 w_7200_15600.n0 GNDA 0.337884f
C166 w_7200_15600.n1 GNDA 0.299565f
C167 w_7200_15600.n2 GNDA 0.211497f
C168 w_7200_15600.n3 GNDA 0.032403f
C169 w_7200_15600.t44 GNDA 0.027783f
C170 w_7200_15600.t33 GNDA 0.017313f
C171 w_7200_15600.t32 GNDA 0.017313f
C172 w_7200_15600.t38 GNDA 0.027282f
C173 w_7200_15600.n4 GNDA 0.039398f
C174 w_7200_15600.n5 GNDA 0.010281f
C175 w_7200_15600.t34 GNDA 0.032163f
C176 w_7200_15600.n6 GNDA 0.012329f
C177 w_7200_15600.n7 GNDA 0.022014f
C178 w_7200_15600.n8 GNDA 0.022014f
C179 w_7200_15600.n9 GNDA 0.022014f
C180 w_7200_15600.n10 GNDA 0.022014f
C181 w_7200_15600.n11 GNDA 0.022014f
C182 w_7200_15600.n12 GNDA 0.022014f
C183 w_7200_15600.n13 GNDA 0.022014f
C184 w_7200_15600.n14 GNDA 0.022014f
C185 w_7200_15600.n31 GNDA 0.011391f
C186 w_7200_15600.n33 GNDA 0.063067f
C187 w_7200_15600.t35 GNDA 0.066889f
C188 w_7200_15600.t14 GNDA 0.0688f
C189 w_7200_15600.t10 GNDA 0.0688f
C190 w_7200_15600.t28 GNDA 0.0688f
C191 w_7200_15600.t2 GNDA 0.0688f
C192 w_7200_15600.t12 GNDA 0.0688f
C193 w_7200_15600.t22 GNDA 0.0688f
C194 w_7200_15600.t20 GNDA 0.0688f
C195 w_7200_15600.t0 GNDA 0.0688f
C196 w_7200_15600.t6 GNDA 0.0688f
C197 w_7200_15600.t16 GNDA 0.0688f
C198 w_7200_15600.t26 GNDA 0.0688f
C199 w_7200_15600.t24 GNDA 0.0688f
C200 w_7200_15600.t4 GNDA 0.0688f
C201 w_7200_15600.t8 GNDA 0.0688f
C202 w_7200_15600.t18 GNDA 0.0688f
C203 w_7200_15600.t30 GNDA 0.0688f
C204 w_7200_15600.t41 GNDA 0.066889f
C205 w_7200_15600.n34 GNDA 0.063067f
C206 w_7200_15600.n42 GNDA 0.012427f
C207 w_7200_15600.t40 GNDA 0.032163f
C208 w_7200_15600.n50 GNDA 0.01299f
C209 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t3 GNDA 0.025303f
C210 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t14 GNDA 0.025303f
C211 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 GNDA 0.079574f
C212 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t1 GNDA 0.025303f
C213 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t2 GNDA 0.025303f
C214 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 GNDA 0.054277f
C215 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 GNDA 4.14756f
C216 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 GNDA 0.088012f
C217 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 GNDA 0.151434f
C218 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t5 GNDA 0.075909f
C219 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t9 GNDA 0.075909f
C220 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 GNDA 0.162355f
C221 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 GNDA 0.507845f
C222 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t4 GNDA 0.075909f
C223 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t11 GNDA 0.075909f
C224 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 GNDA 0.162355f
C225 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 GNDA 0.494091f
C226 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 GNDA 0.151434f
C227 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 GNDA 0.088012f
C228 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t6 GNDA 0.075909f
C229 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t10 GNDA 0.075909f
C230 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 GNDA 0.162355f
C231 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 GNDA 0.494091f
C232 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 GNDA 0.088012f
C233 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t7 GNDA 0.075909f
C234 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t12 GNDA 0.075909f
C235 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 GNDA 0.162355f
C236 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 GNDA 0.494091f
C237 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 GNDA 0.151434f
C238 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t8 GNDA 0.075909f
C239 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t13 GNDA 0.075909f
C240 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 GNDA 0.162355f
C241 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 GNDA 0.500968f
C242 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 GNDA 0.196238f
C243 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 GNDA 3.42529f
C244 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t0 GNDA 0.31557f
C245 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 GNDA 0.057368f
C246 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 GNDA 0.101473f
C247 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t2 GNDA 0.036321f
C248 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t6 GNDA 0.036321f
C249 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 GNDA 0.074261f
C250 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 GNDA 0.249441f
C251 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t1 GNDA 0.036321f
C252 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t9 GNDA 0.036321f
C253 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 GNDA 0.074261f
C254 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 GNDA 0.240213f
C255 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 GNDA 0.097542f
C256 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 GNDA 0.057368f
C257 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t4 GNDA 0.036321f
C258 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t8 GNDA 0.036321f
C259 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 GNDA 0.074261f
C260 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 GNDA 0.240213f
C261 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 GNDA 0.059466f
C262 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t3 GNDA 0.036321f
C263 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t7 GNDA 0.036321f
C264 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 GNDA 0.074261f
C265 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 GNDA 0.240213f
C266 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 GNDA 0.101473f
C267 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t10 GNDA 0.036321f
C268 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t5 GNDA 0.036321f
C269 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 GNDA 0.074261f
C270 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 GNDA 0.244959f
C271 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 GNDA 2.23639f
C272 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t0 GNDA 0.339365f
C273 a_7460_6300.t8 GNDA 0.020006f
C274 a_7460_6300.n0 GNDA 0.210468f
C275 a_7460_6300.t4 GNDA 0.020006f
C276 a_7460_6300.t7 GNDA 0.020006f
C277 a_7460_6300.n1 GNDA 0.040763f
C278 a_7460_6300.n2 GNDA 0.365375f
C279 a_7460_6300.n3 GNDA 0.319666f
C280 a_7460_6300.t1 GNDA 0.020006f
C281 a_7460_6300.t5 GNDA 0.020006f
C282 a_7460_6300.n4 GNDA 0.040763f
C283 a_7460_6300.n5 GNDA 0.306668f
C284 a_7460_6300.n6 GNDA 0.335179f
C285 a_7460_6300.t14 GNDA 0.020006f
C286 a_7460_6300.t12 GNDA 0.020006f
C287 a_7460_6300.n7 GNDA 0.040763f
C288 a_7460_6300.n8 GNDA 0.191134f
C289 a_7460_6300.t19 GNDA 0.020006f
C290 a_7460_6300.t17 GNDA 0.020006f
C291 a_7460_6300.n9 GNDA 0.040763f
C292 a_7460_6300.n10 GNDA 0.300378f
C293 a_7460_6300.n11 GNDA 0.215758f
C294 a_7460_6300.n12 GNDA 0.206718f
C295 a_7460_6300.t11 GNDA 0.020006f
C296 a_7460_6300.t15 GNDA 0.020006f
C297 a_7460_6300.n13 GNDA 0.040763f
C298 a_7460_6300.n14 GNDA 0.300378f
C299 a_7460_6300.t13 GNDA 0.020006f
C300 a_7460_6300.t18 GNDA 0.020006f
C301 a_7460_6300.n15 GNDA 0.040763f
C302 a_7460_6300.n16 GNDA 0.279938f
C303 a_7460_6300.n17 GNDA 0.206718f
C304 a_7460_6300.n18 GNDA 0.122442f
C305 a_7460_6300.t0 GNDA 0.020006f
C306 a_7460_6300.t16 GNDA 0.020006f
C307 a_7460_6300.n19 GNDA 0.040763f
C308 a_7460_6300.n20 GNDA 0.279938f
C309 a_7460_6300.n21 GNDA 0.127024f
C310 a_7460_6300.n22 GNDA 0.208769f
C311 a_7460_6300.n23 GNDA 0.121174f
C312 a_7460_6300.n24 GNDA 0.18461f
C313 a_7460_6300.t6 GNDA 0.020006f
C314 a_7460_6300.t2 GNDA 0.020006f
C315 a_7460_6300.n25 GNDA 0.040763f
C316 a_7460_6300.n26 GNDA 0.233788f
C317 a_7460_6300.n27 GNDA 0.319666f
C318 a_7460_6300.t9 GNDA 0.020006f
C319 a_7460_6300.t3 GNDA 0.020006f
C320 a_7460_6300.n28 GNDA 0.040763f
C321 a_7460_6300.n29 GNDA 0.306668f
C322 a_7460_6300.n30 GNDA 0.324795f
C323 a_7460_6300.n31 GNDA 0.218329f
C324 a_7460_6300.n32 GNDA 0.306668f
C325 a_7460_6300.n33 GNDA 0.040763f
C326 a_7460_6300.t10 GNDA 0.020006f
C327 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 GNDA 0.408216f
C328 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 GNDA 0.318908f
C329 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 GNDA 0.362794f
C330 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t10 GNDA 0.014742f
C331 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t4 GNDA 0.014742f
C332 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t12 GNDA 0.014742f
C333 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 GNDA 0.031178f
C334 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 GNDA 0.293793f
C335 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t13 GNDA 0.012162f
C336 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t19 GNDA 0.012162f
C337 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t21 GNDA 0.012162f
C338 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t9 GNDA 0.012162f
C339 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t15 GNDA 0.012162f
C340 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t20 GNDA 0.012162f
C341 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t17 GNDA 0.012162f
C342 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t11 GNDA 0.026351f
C343 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 GNDA 0.041093f
C344 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 GNDA 0.032064f
C345 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 GNDA 0.028584f
C346 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 GNDA 0.04506f
C347 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 GNDA 0.028584f
C348 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 GNDA 0.032064f
C349 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 GNDA 0.032064f
C350 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 GNDA 0.028584f
C351 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t7 GNDA 0.012162f
C352 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t18 GNDA 0.026351f
C353 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 GNDA 0.037614f
C354 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 GNDA 0.04506f
C355 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t3 GNDA 0.014742f
C356 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t6 GNDA 0.014742f
C357 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 GNDA 0.030038f
C358 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t2 GNDA 0.014742f
C359 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t0 GNDA 0.014742f
C360 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 GNDA 0.030038f
C361 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 GNDA 0.249418f
C362 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 GNDA 0.316023f
C363 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t1 GNDA 0.014742f
C364 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t5 GNDA 0.014742f
C365 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 GNDA 0.030038f
C366 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 GNDA 0.249418f
C367 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 GNDA 0.320943f
C368 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 GNDA 0.239385f
C369 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 GNDA 0.23177f
C370 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t14 GNDA 0.014742f
C371 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t8 GNDA 0.014742f
C372 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 GNDA 0.031178f
C373 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 GNDA 0.348011f
C374 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 GNDA 0.031178f
C375 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t16 GNDA 0.014742f
C376 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 GNDA 0.20958f
C377 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 GNDA 0.20958f
C378 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 GNDA 0.191254f
C379 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 GNDA 0.265929f
C380 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 GNDA 0.137376f
C381 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 GNDA 0.161756f
C382 two_stage_opamp_dummy_magic_23_0.V_err_gate.t3 GNDA 0.025476f
C383 two_stage_opamp_dummy_magic_23_0.V_err_gate.t4 GNDA 0.025476f
C384 two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 GNDA 0.329843f
C385 two_stage_opamp_dummy_magic_23_0.V_err_gate.t19 GNDA 0.010509f
C386 two_stage_opamp_dummy_magic_23_0.V_err_gate.t15 GNDA 0.010509f
C387 two_stage_opamp_dummy_magic_23_0.V_err_gate.t25 GNDA 0.010509f
C388 two_stage_opamp_dummy_magic_23_0.V_err_gate.t33 GNDA 0.010509f
C389 two_stage_opamp_dummy_magic_23_0.V_err_gate.t23 GNDA 0.010509f
C390 two_stage_opamp_dummy_magic_23_0.V_err_gate.t32 GNDA 0.010509f
C391 two_stage_opamp_dummy_magic_23_0.V_err_gate.t22 GNDA 0.010509f
C392 two_stage_opamp_dummy_magic_23_0.V_err_gate.t30 GNDA 0.010509f
C393 two_stage_opamp_dummy_magic_23_0.V_err_gate.t20 GNDA 0.010509f
C394 two_stage_opamp_dummy_magic_23_0.V_err_gate.t24 GNDA 0.010509f
C395 two_stage_opamp_dummy_magic_23_0.V_err_gate.t16 GNDA 0.022769f
C396 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 GNDA 0.035507f
C397 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 GNDA 0.027705f
C398 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 GNDA 0.027705f
C399 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 GNDA 0.027705f
C400 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 GNDA 0.027705f
C401 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 GNDA 0.027705f
C402 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 GNDA 0.027705f
C403 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 GNDA 0.027705f
C404 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 GNDA 0.027705f
C405 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 GNDA 0.022724f
C406 two_stage_opamp_dummy_magic_23_0.V_err_gate.t29 GNDA 0.010509f
C407 two_stage_opamp_dummy_magic_23_0.V_err_gate.t26 GNDA 0.010509f
C408 two_stage_opamp_dummy_magic_23_0.V_err_gate.t17 GNDA 0.010509f
C409 two_stage_opamp_dummy_magic_23_0.V_err_gate.t27 GNDA 0.010509f
C410 two_stage_opamp_dummy_magic_23_0.V_err_gate.t18 GNDA 0.010509f
C411 two_stage_opamp_dummy_magic_23_0.V_err_gate.t28 GNDA 0.010509f
C412 two_stage_opamp_dummy_magic_23_0.V_err_gate.t21 GNDA 0.010509f
C413 two_stage_opamp_dummy_magic_23_0.V_err_gate.t31 GNDA 0.010509f
C414 two_stage_opamp_dummy_magic_23_0.V_err_gate.t14 GNDA 0.026272f
C415 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 GNDA 0.054932f
C416 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 GNDA 0.027705f
C417 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 GNDA 0.027705f
C418 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 GNDA 0.027705f
C419 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 GNDA 0.027705f
C420 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 GNDA 0.027705f
C421 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 GNDA 0.027705f
C422 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 GNDA 0.022724f
C423 two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 GNDA 0.034919f
C424 two_stage_opamp_dummy_magic_23_0.V_err_gate.t6 GNDA 0.012738f
C425 two_stage_opamp_dummy_magic_23_0.V_err_gate.t11 GNDA 0.012738f
C426 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 GNDA 0.025954f
C427 two_stage_opamp_dummy_magic_23_0.V_err_gate.t10 GNDA 0.012738f
C428 two_stage_opamp_dummy_magic_23_0.V_err_gate.t1 GNDA 0.012738f
C429 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 GNDA 0.025954f
C430 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 GNDA 0.178239f
C431 two_stage_opamp_dummy_magic_23_0.V_err_gate.t9 GNDA 0.012738f
C432 two_stage_opamp_dummy_magic_23_0.V_err_gate.t8 GNDA 0.012738f
C433 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 GNDA 0.025954f
C434 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 GNDA 0.178239f
C435 two_stage_opamp_dummy_magic_23_0.V_err_gate.t2 GNDA 0.012738f
C436 two_stage_opamp_dummy_magic_23_0.V_err_gate.t0 GNDA 0.012738f
C437 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 GNDA 0.025954f
C438 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 GNDA 0.178239f
C439 two_stage_opamp_dummy_magic_23_0.V_err_gate.t5 GNDA 0.012738f
C440 two_stage_opamp_dummy_magic_23_0.V_err_gate.t7 GNDA 0.012738f
C441 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 GNDA 0.025954f
C442 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 GNDA 0.178239f
C443 two_stage_opamp_dummy_magic_23_0.V_err_gate.t12 GNDA 0.012738f
C444 two_stage_opamp_dummy_magic_23_0.V_err_gate.t13 GNDA 0.012738f
C445 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 GNDA 0.025954f
C446 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 GNDA 0.184707f
C447 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 GNDA 0.095072f
C448 two_stage_opamp_dummy_magic_23_0.err_amp_out.t12 GNDA 0.054088f
C449 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 GNDA 0.012001f
C450 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 GNDA 0.124861f
C451 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 GNDA 0.012001f
C452 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 GNDA 0.10815f
C453 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 GNDA 0.095072f
C454 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 GNDA 0.719147f
C455 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 GNDA 0.012001f
C456 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 GNDA 0.10815f
C457 two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 GNDA 0.057175f
C458 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 GNDA 0.012844f
C459 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 GNDA 0.012527f
C460 two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 GNDA 0.325317f
C461 two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 GNDA 0.012527f
C462 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 GNDA 0.845522f
C463 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 GNDA 0.630165f
C464 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 GNDA 0.630165f
C465 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 GNDA 0.392203f
C466 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 GNDA 0.614283f
C467 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 GNDA 0.611494f
C468 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 GNDA 0.620939f
C469 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 GNDA 0.639167f
C470 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 GNDA 0.348058f
C471 two_stage_opamp_dummy_magic_23_0.V_err_p.t8 GNDA 0.023181f
C472 two_stage_opamp_dummy_magic_23_0.V_err_p.t6 GNDA 0.023181f
C473 two_stage_opamp_dummy_magic_23_0.V_err_p.t18 GNDA 0.023181f
C474 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 GNDA 0.047234f
C475 two_stage_opamp_dummy_magic_23_0.V_err_p.t21 GNDA 0.023181f
C476 two_stage_opamp_dummy_magic_23_0.V_err_p.t7 GNDA 0.023181f
C477 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 GNDA 0.047234f
C478 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 GNDA 0.324373f
C479 two_stage_opamp_dummy_magic_23_0.V_err_p.t4 GNDA 0.023181f
C480 two_stage_opamp_dummy_magic_23_0.V_err_p.t9 GNDA 0.023181f
C481 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 GNDA 0.047234f
C482 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 GNDA 0.324373f
C483 two_stage_opamp_dummy_magic_23_0.V_err_p.t5 GNDA 0.023181f
C484 two_stage_opamp_dummy_magic_23_0.V_err_p.t10 GNDA 0.023181f
C485 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 GNDA 0.047234f
C486 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 GNDA 0.324373f
C487 two_stage_opamp_dummy_magic_23_0.V_err_p.t3 GNDA 0.023181f
C488 two_stage_opamp_dummy_magic_23_0.V_err_p.t0 GNDA 0.023181f
C489 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 GNDA 0.047234f
C490 two_stage_opamp_dummy_magic_23_0.V_err_p.t13 GNDA 0.023181f
C491 two_stage_opamp_dummy_magic_23_0.V_err_p.t2 GNDA 0.023181f
C492 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 GNDA 0.047234f
C493 two_stage_opamp_dummy_magic_23_0.V_err_p.t15 GNDA 0.023181f
C494 two_stage_opamp_dummy_magic_23_0.V_err_p.t11 GNDA 0.023181f
C495 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 GNDA 0.047234f
C496 two_stage_opamp_dummy_magic_23_0.V_err_p.t1 GNDA 0.023181f
C497 two_stage_opamp_dummy_magic_23_0.V_err_p.t16 GNDA 0.023181f
C498 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 GNDA 0.047234f
C499 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 GNDA 0.324373f
C500 two_stage_opamp_dummy_magic_23_0.V_err_p.t12 GNDA 0.023181f
C501 two_stage_opamp_dummy_magic_23_0.V_err_p.t17 GNDA 0.023181f
C502 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 GNDA 0.047234f
C503 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 GNDA 0.324373f
C504 two_stage_opamp_dummy_magic_23_0.V_err_p.t20 GNDA 0.023181f
C505 two_stage_opamp_dummy_magic_23_0.V_err_p.t14 GNDA 0.023181f
C506 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 GNDA 0.047234f
C507 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 GNDA 0.324373f
C508 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 GNDA 0.392203f
C509 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 GNDA 0.047234f
C510 two_stage_opamp_dummy_magic_23_0.V_err_p.t19 GNDA 0.023181f
C511 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t12 GNDA 0.011605f
C512 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t17 GNDA 0.011605f
C513 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t11 GNDA 0.011605f
C514 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t16 GNDA 0.011605f
C515 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t9 GNDA 0.011605f
C516 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t8 GNDA 0.011605f
C517 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t14 GNDA 0.011605f
C518 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t7 GNDA 0.011605f
C519 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t13 GNDA 0.011605f
C520 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t15 GNDA 0.035602f
C521 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 GNDA 0.048365f
C522 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 GNDA 0.038911f
C523 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 GNDA 0.038911f
C524 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 GNDA 0.229146f
C525 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 GNDA 0.229146f
C526 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 GNDA 0.038911f
C527 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 GNDA 0.038911f
C528 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 GNDA 0.038911f
C529 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 GNDA 0.057863f
C530 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t6 GNDA 0.293124f
C531 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t10 GNDA 0.089212f
C532 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 GNDA 1.59901f
C533 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t0 GNDA 0.054613f
C534 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t4 GNDA 0.054613f
C535 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 GNDA 0.192596f
C536 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t2 GNDA 0.054613f
C537 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t5 GNDA 0.054613f
C538 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 GNDA 0.183176f
C539 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 GNDA 0.862116f
C540 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t3 GNDA 0.054613f
C541 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t1 GNDA 0.054613f
C542 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 GNDA 0.183176f
C543 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 GNDA 0.615045f
C544 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 GNDA 1.41464f
C545 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t3 GNDA 0.032304f
C546 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t0 GNDA 0.032304f
C547 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 GNDA 0.101592f
C548 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t2 GNDA 0.032304f
C549 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t1 GNDA 0.032304f
C550 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 GNDA 0.069296f
C551 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 GNDA 2.19459f
C552 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t14 GNDA 0.401158f
C553 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 GNDA 0.112365f
C554 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 GNDA 0.193336f
C555 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t4 GNDA 0.096913f
C556 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t8 GNDA 0.096913f
C557 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 GNDA 0.207278f
C558 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 GNDA 0.648366f
C559 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t13 GNDA 0.096913f
C560 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t11 GNDA 0.096913f
C561 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 GNDA 0.207278f
C562 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 GNDA 0.630805f
C563 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 GNDA 0.193336f
C564 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 GNDA 0.112365f
C565 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t6 GNDA 0.096913f
C566 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t10 GNDA 0.096913f
C567 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 GNDA 0.207278f
C568 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 GNDA 0.630805f
C569 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 GNDA 0.112365f
C570 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t5 GNDA 0.096913f
C571 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t9 GNDA 0.096913f
C572 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 GNDA 0.207278f
C573 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 GNDA 0.630805f
C574 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 GNDA 0.193336f
C575 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t12 GNDA 0.096913f
C576 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t7 GNDA 0.096913f
C577 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 GNDA 0.207278f
C578 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 GNDA 0.639586f
C579 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 GNDA 0.252889f
C580 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 GNDA 2.58687f
C581 bgr_11_0.V_CMFB_S4 GNDA 3.3614f
C582 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 GNDA 0.057181f
C583 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 GNDA 0.101143f
C584 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t3 GNDA 0.036202f
C585 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t7 GNDA 0.036202f
C586 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 GNDA 0.074019f
C587 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 GNDA 0.248628f
C588 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t2 GNDA 0.036202f
C589 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t9 GNDA 0.036202f
C590 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 GNDA 0.074019f
C591 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 GNDA 0.23943f
C592 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 GNDA 0.097224f
C593 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 GNDA 0.057181f
C594 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t4 GNDA 0.036202f
C595 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t8 GNDA 0.036202f
C596 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 GNDA 0.074019f
C597 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 GNDA 0.23943f
C598 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 GNDA 0.059272f
C599 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t5 GNDA 0.036202f
C600 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t10 GNDA 0.036202f
C601 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 GNDA 0.074019f
C602 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 GNDA 0.23943f
C603 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 GNDA 0.101143f
C604 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t6 GNDA 0.036202f
C605 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t1 GNDA 0.036202f
C606 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 GNDA 0.074019f
C607 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 GNDA 0.244161f
C608 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 GNDA 2.24416f
C609 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t0 GNDA 0.339492f
C610 two_stage_opamp_dummy_magic_23_0.VD4.t33 GNDA 0.060801f
C611 two_stage_opamp_dummy_magic_23_0.VD4.t29 GNDA 0.060801f
C612 two_stage_opamp_dummy_magic_23_0.VD4.n0 GNDA 0.154331f
C613 two_stage_opamp_dummy_magic_23_0.VD4.n1 GNDA 0.431096f
C614 two_stage_opamp_dummy_magic_23_0.VD4.t3 GNDA 0.106612f
C615 two_stage_opamp_dummy_magic_23_0.VD4.t2 GNDA 0.216278f
C616 two_stage_opamp_dummy_magic_23_0.VD4.t23 GNDA 0.060801f
C617 two_stage_opamp_dummy_magic_23_0.VD4.t27 GNDA 0.060801f
C618 two_stage_opamp_dummy_magic_23_0.VD4.n2 GNDA 0.154331f
C619 two_stage_opamp_dummy_magic_23_0.VD4.n3 GNDA 0.431096f
C620 two_stage_opamp_dummy_magic_23_0.VD4.t37 GNDA 0.060801f
C621 two_stage_opamp_dummy_magic_23_0.VD4.t19 GNDA 0.060801f
C622 two_stage_opamp_dummy_magic_23_0.VD4.n4 GNDA 0.154331f
C623 two_stage_opamp_dummy_magic_23_0.VD4.n5 GNDA 0.431096f
C624 two_stage_opamp_dummy_magic_23_0.VD4.t31 GNDA 0.060801f
C625 two_stage_opamp_dummy_magic_23_0.VD4.t35 GNDA 0.060801f
C626 two_stage_opamp_dummy_magic_23_0.VD4.n6 GNDA 0.154331f
C627 two_stage_opamp_dummy_magic_23_0.VD4.n7 GNDA 0.431096f
C628 two_stage_opamp_dummy_magic_23_0.VD4.t21 GNDA 0.060801f
C629 two_stage_opamp_dummy_magic_23_0.VD4.t25 GNDA 0.060801f
C630 two_stage_opamp_dummy_magic_23_0.VD4.n8 GNDA 0.154331f
C631 two_stage_opamp_dummy_magic_23_0.VD4.n9 GNDA 0.481515f
C632 two_stage_opamp_dummy_magic_23_0.VD4.t0 GNDA 0.106612f
C633 two_stage_opamp_dummy_magic_23_0.VD4.n10 GNDA 0.316782f
C634 two_stage_opamp_dummy_magic_23_0.VD4.n11 GNDA 0.627403f
C635 two_stage_opamp_dummy_magic_23_0.VD4.t1 GNDA 0.518263f
C636 two_stage_opamp_dummy_magic_23_0.VD4.t20 GNDA 0.406498f
C637 two_stage_opamp_dummy_magic_23_0.VD4.t24 GNDA 0.406498f
C638 two_stage_opamp_dummy_magic_23_0.VD4.t30 GNDA 0.406498f
C639 two_stage_opamp_dummy_magic_23_0.VD4.t34 GNDA 0.406498f
C640 two_stage_opamp_dummy_magic_23_0.VD4.t36 GNDA 0.406498f
C641 two_stage_opamp_dummy_magic_23_0.VD4.t18 GNDA 0.406498f
C642 two_stage_opamp_dummy_magic_23_0.VD4.t22 GNDA 0.406498f
C643 two_stage_opamp_dummy_magic_23_0.VD4.t26 GNDA 0.406498f
C644 two_stage_opamp_dummy_magic_23_0.VD4.t32 GNDA 0.406498f
C645 two_stage_opamp_dummy_magic_23_0.VD4.t28 GNDA 0.406498f
C646 two_stage_opamp_dummy_magic_23_0.VD4.t4 GNDA 0.518263f
C647 two_stage_opamp_dummy_magic_23_0.VD4.t5 GNDA 0.216278f
C648 two_stage_opamp_dummy_magic_23_0.VD4.n12 GNDA 0.627403f
C649 two_stage_opamp_dummy_magic_23_0.VD4.n13 GNDA 0.311031f
C650 two_stage_opamp_dummy_magic_23_0.VD4.n14 GNDA 0.102448f
C651 two_stage_opamp_dummy_magic_23_0.VD4.n15 GNDA 0.065949f
C652 two_stage_opamp_dummy_magic_23_0.VD4.n16 GNDA 0.065949f
C653 two_stage_opamp_dummy_magic_23_0.VD4.t8 GNDA 0.060801f
C654 two_stage_opamp_dummy_magic_23_0.VD4.t16 GNDA 0.060801f
C655 two_stage_opamp_dummy_magic_23_0.VD4.n17 GNDA 0.124375f
C656 two_stage_opamp_dummy_magic_23_0.VD4.n18 GNDA 0.402689f
C657 two_stage_opamp_dummy_magic_23_0.VD4.n19 GNDA 0.112503f
C658 two_stage_opamp_dummy_magic_23_0.VD4.t14 GNDA 0.060801f
C659 two_stage_opamp_dummy_magic_23_0.VD4.t7 GNDA 0.060801f
C660 two_stage_opamp_dummy_magic_23_0.VD4.n20 GNDA 0.124375f
C661 two_stage_opamp_dummy_magic_23_0.VD4.n21 GNDA 0.391692f
C662 two_stage_opamp_dummy_magic_23_0.VD4.n22 GNDA 0.112503f
C663 two_stage_opamp_dummy_magic_23_0.VD4.t12 GNDA 0.060801f
C664 two_stage_opamp_dummy_magic_23_0.VD4.t11 GNDA 0.060801f
C665 two_stage_opamp_dummy_magic_23_0.VD4.n23 GNDA 0.124375f
C666 two_stage_opamp_dummy_magic_23_0.VD4.n24 GNDA 0.391692f
C667 two_stage_opamp_dummy_magic_23_0.VD4.n25 GNDA 0.065949f
C668 two_stage_opamp_dummy_magic_23_0.VD4.n26 GNDA 0.065949f
C669 two_stage_opamp_dummy_magic_23_0.VD4.t9 GNDA 0.060801f
C670 two_stage_opamp_dummy_magic_23_0.VD4.t10 GNDA 0.060801f
C671 two_stage_opamp_dummy_magic_23_0.VD4.n27 GNDA 0.124375f
C672 two_stage_opamp_dummy_magic_23_0.VD4.n28 GNDA 0.391692f
C673 two_stage_opamp_dummy_magic_23_0.VD4.n29 GNDA 0.065949f
C674 two_stage_opamp_dummy_magic_23_0.VD4.t13 GNDA 0.060801f
C675 two_stage_opamp_dummy_magic_23_0.VD4.t6 GNDA 0.060801f
C676 two_stage_opamp_dummy_magic_23_0.VD4.n30 GNDA 0.124375f
C677 two_stage_opamp_dummy_magic_23_0.VD4.n31 GNDA 0.391692f
C678 two_stage_opamp_dummy_magic_23_0.VD4.n32 GNDA 0.112503f
C679 two_stage_opamp_dummy_magic_23_0.VD4.t17 GNDA 0.060801f
C680 two_stage_opamp_dummy_magic_23_0.VD4.t15 GNDA 0.060801f
C681 two_stage_opamp_dummy_magic_23_0.VD4.n33 GNDA 0.124375f
C682 two_stage_opamp_dummy_magic_23_0.VD4.n34 GNDA 0.39719f
C683 two_stage_opamp_dummy_magic_23_0.VD4.n35 GNDA 0.183347f
C684 two_stage_opamp_dummy_magic_23_0.V_source.t29 GNDA 0.038168f
C685 two_stage_opamp_dummy_magic_23_0.V_source.n0 GNDA 0.052428f
C686 two_stage_opamp_dummy_magic_23_0.V_source.n1 GNDA 0.05567f
C687 two_stage_opamp_dummy_magic_23_0.V_source.n2 GNDA 0.052428f
C688 two_stage_opamp_dummy_magic_23_0.V_source.n3 GNDA 0.096361f
C689 two_stage_opamp_dummy_magic_23_0.V_source.t5 GNDA 0.022901f
C690 two_stage_opamp_dummy_magic_23_0.V_source.t6 GNDA 0.022901f
C691 two_stage_opamp_dummy_magic_23_0.V_source.n4 GNDA 0.049829f
C692 two_stage_opamp_dummy_magic_23_0.V_source.n5 GNDA 0.153174f
C693 two_stage_opamp_dummy_magic_23_0.V_source.n6 GNDA 0.051154f
C694 two_stage_opamp_dummy_magic_23_0.V_source.t9 GNDA 0.022901f
C695 two_stage_opamp_dummy_magic_23_0.V_source.t8 GNDA 0.022901f
C696 two_stage_opamp_dummy_magic_23_0.V_source.n7 GNDA 0.049829f
C697 two_stage_opamp_dummy_magic_23_0.V_source.n8 GNDA 0.200044f
C698 two_stage_opamp_dummy_magic_23_0.V_source.n9 GNDA 0.087575f
C699 two_stage_opamp_dummy_magic_23_0.V_source.t13 GNDA 0.022901f
C700 two_stage_opamp_dummy_magic_23_0.V_source.t40 GNDA 0.022901f
C701 two_stage_opamp_dummy_magic_23_0.V_source.n10 GNDA 0.049829f
C702 two_stage_opamp_dummy_magic_23_0.V_source.n11 GNDA 0.192055f
C703 two_stage_opamp_dummy_magic_23_0.V_source.n12 GNDA 0.083262f
C704 two_stage_opamp_dummy_magic_23_0.V_source.t17 GNDA 0.022901f
C705 two_stage_opamp_dummy_magic_23_0.V_source.t4 GNDA 0.022901f
C706 two_stage_opamp_dummy_magic_23_0.V_source.n13 GNDA 0.049829f
C707 two_stage_opamp_dummy_magic_23_0.V_source.n14 GNDA 0.192055f
C708 two_stage_opamp_dummy_magic_23_0.V_source.n15 GNDA 0.048946f
C709 two_stage_opamp_dummy_magic_23_0.V_source.n16 GNDA 0.083262f
C710 two_stage_opamp_dummy_magic_23_0.V_source.t16 GNDA 0.022901f
C711 two_stage_opamp_dummy_magic_23_0.V_source.t1 GNDA 0.022901f
C712 two_stage_opamp_dummy_magic_23_0.V_source.n17 GNDA 0.049829f
C713 two_stage_opamp_dummy_magic_23_0.V_source.n18 GNDA 0.192055f
C714 two_stage_opamp_dummy_magic_23_0.V_source.n19 GNDA 0.051154f
C715 two_stage_opamp_dummy_magic_23_0.V_source.n20 GNDA 0.051154f
C716 two_stage_opamp_dummy_magic_23_0.V_source.n21 GNDA 0.083262f
C717 two_stage_opamp_dummy_magic_23_0.V_source.t0 GNDA 0.022901f
C718 two_stage_opamp_dummy_magic_23_0.V_source.t15 GNDA 0.022901f
C719 two_stage_opamp_dummy_magic_23_0.V_source.n22 GNDA 0.049829f
C720 two_stage_opamp_dummy_magic_23_0.V_source.n23 GNDA 0.200044f
C721 two_stage_opamp_dummy_magic_23_0.V_source.t10 GNDA 0.022901f
C722 two_stage_opamp_dummy_magic_23_0.V_source.t7 GNDA 0.022901f
C723 two_stage_opamp_dummy_magic_23_0.V_source.n24 GNDA 0.049829f
C724 two_stage_opamp_dummy_magic_23_0.V_source.n25 GNDA 0.192055f
C725 two_stage_opamp_dummy_magic_23_0.V_source.n26 GNDA 0.087575f
C726 two_stage_opamp_dummy_magic_23_0.V_source.n27 GNDA 0.051154f
C727 two_stage_opamp_dummy_magic_23_0.V_source.t11 GNDA 0.022901f
C728 two_stage_opamp_dummy_magic_23_0.V_source.t18 GNDA 0.022901f
C729 two_stage_opamp_dummy_magic_23_0.V_source.n28 GNDA 0.049829f
C730 two_stage_opamp_dummy_magic_23_0.V_source.n29 GNDA 0.192055f
C731 two_stage_opamp_dummy_magic_23_0.V_source.n30 GNDA 0.048946f
C732 two_stage_opamp_dummy_magic_23_0.V_source.t19 GNDA 0.022901f
C733 two_stage_opamp_dummy_magic_23_0.V_source.t12 GNDA 0.022901f
C734 two_stage_opamp_dummy_magic_23_0.V_source.n31 GNDA 0.049829f
C735 two_stage_opamp_dummy_magic_23_0.V_source.n32 GNDA 0.192055f
C736 two_stage_opamp_dummy_magic_23_0.V_source.n33 GNDA 0.083262f
C737 two_stage_opamp_dummy_magic_23_0.V_source.t21 GNDA 0.022901f
C738 two_stage_opamp_dummy_magic_23_0.V_source.t3 GNDA 0.022901f
C739 two_stage_opamp_dummy_magic_23_0.V_source.n34 GNDA 0.049829f
C740 two_stage_opamp_dummy_magic_23_0.V_source.n35 GNDA 0.195998f
C741 two_stage_opamp_dummy_magic_23_0.V_source.n36 GNDA 0.125964f
C742 two_stage_opamp_dummy_magic_23_0.V_source.n37 GNDA 0.120611f
C743 two_stage_opamp_dummy_magic_23_0.V_source.n38 GNDA 0.087586f
C744 two_stage_opamp_dummy_magic_23_0.V_source.t20 GNDA 0.038168f
C745 two_stage_opamp_dummy_magic_23_0.V_source.t14 GNDA 0.038168f
C746 two_stage_opamp_dummy_magic_23_0.V_source.n39 GNDA 0.081597f
C747 two_stage_opamp_dummy_magic_23_0.V_source.n40 GNDA 0.294282f
C748 two_stage_opamp_dummy_magic_23_0.V_source.t32 GNDA 0.038168f
C749 two_stage_opamp_dummy_magic_23_0.V_source.t36 GNDA 0.038168f
C750 two_stage_opamp_dummy_magic_23_0.V_source.n41 GNDA 0.081597f
C751 two_stage_opamp_dummy_magic_23_0.V_source.n42 GNDA 0.285878f
C752 two_stage_opamp_dummy_magic_23_0.V_source.n43 GNDA 0.090055f
C753 two_stage_opamp_dummy_magic_23_0.V_source.n44 GNDA 0.045802f
C754 two_stage_opamp_dummy_magic_23_0.V_source.n45 GNDA 0.099442f
C755 two_stage_opamp_dummy_magic_23_0.V_source.t26 GNDA 0.038168f
C756 two_stage_opamp_dummy_magic_23_0.V_source.t34 GNDA 0.038168f
C757 two_stage_opamp_dummy_magic_23_0.V_source.n46 GNDA 0.081597f
C758 two_stage_opamp_dummy_magic_23_0.V_source.n47 GNDA 0.185859f
C759 two_stage_opamp_dummy_magic_23_0.V_source.t2 GNDA 0.079851f
C760 two_stage_opamp_dummy_magic_23_0.V_source.n48 GNDA 0.258116f
C761 two_stage_opamp_dummy_magic_23_0.V_source.n49 GNDA 0.045802f
C762 two_stage_opamp_dummy_magic_23_0.V_source.t24 GNDA 0.038168f
C763 two_stage_opamp_dummy_magic_23_0.V_source.t33 GNDA 0.038168f
C764 two_stage_opamp_dummy_magic_23_0.V_source.n50 GNDA 0.081597f
C765 two_stage_opamp_dummy_magic_23_0.V_source.n51 GNDA 0.285878f
C766 two_stage_opamp_dummy_magic_23_0.V_source.n52 GNDA 0.05567f
C767 two_stage_opamp_dummy_magic_23_0.V_source.n53 GNDA 0.05567f
C768 two_stage_opamp_dummy_magic_23_0.V_source.t23 GNDA 0.038168f
C769 two_stage_opamp_dummy_magic_23_0.V_source.t31 GNDA 0.038168f
C770 two_stage_opamp_dummy_magic_23_0.V_source.n54 GNDA 0.081597f
C771 two_stage_opamp_dummy_magic_23_0.V_source.n55 GNDA 0.285878f
C772 two_stage_opamp_dummy_magic_23_0.V_source.n56 GNDA 0.052428f
C773 two_stage_opamp_dummy_magic_23_0.V_source.t22 GNDA 0.038168f
C774 two_stage_opamp_dummy_magic_23_0.V_source.t37 GNDA 0.038168f
C775 two_stage_opamp_dummy_magic_23_0.V_source.n57 GNDA 0.081597f
C776 two_stage_opamp_dummy_magic_23_0.V_source.n58 GNDA 0.285878f
C777 two_stage_opamp_dummy_magic_23_0.V_source.n59 GNDA 0.052428f
C778 two_stage_opamp_dummy_magic_23_0.V_source.n60 GNDA 0.052428f
C779 two_stage_opamp_dummy_magic_23_0.V_source.t27 GNDA 0.038168f
C780 two_stage_opamp_dummy_magic_23_0.V_source.t30 GNDA 0.038168f
C781 two_stage_opamp_dummy_magic_23_0.V_source.n61 GNDA 0.081597f
C782 two_stage_opamp_dummy_magic_23_0.V_source.n62 GNDA 0.285878f
C783 two_stage_opamp_dummy_magic_23_0.V_source.n63 GNDA 0.05567f
C784 two_stage_opamp_dummy_magic_23_0.V_source.t35 GNDA 0.038168f
C785 two_stage_opamp_dummy_magic_23_0.V_source.t25 GNDA 0.038168f
C786 two_stage_opamp_dummy_magic_23_0.V_source.n64 GNDA 0.081597f
C787 two_stage_opamp_dummy_magic_23_0.V_source.n65 GNDA 0.294282f
C788 two_stage_opamp_dummy_magic_23_0.V_source.n66 GNDA 0.090055f
C789 two_stage_opamp_dummy_magic_23_0.V_source.t38 GNDA 0.038168f
C790 two_stage_opamp_dummy_magic_23_0.V_source.t28 GNDA 0.038168f
C791 two_stage_opamp_dummy_magic_23_0.V_source.n67 GNDA 0.081597f
C792 two_stage_opamp_dummy_magic_23_0.V_source.n68 GNDA 0.285878f
C793 two_stage_opamp_dummy_magic_23_0.V_source.n69 GNDA 0.096361f
C794 two_stage_opamp_dummy_magic_23_0.V_source.n70 GNDA 0.05567f
C795 two_stage_opamp_dummy_magic_23_0.V_source.n71 GNDA 0.285878f
C796 two_stage_opamp_dummy_magic_23_0.V_source.n72 GNDA 0.081597f
C797 two_stage_opamp_dummy_magic_23_0.V_source.t39 GNDA 0.038168f
C798 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t7 GNDA 0.021693f
C799 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t4 GNDA 0.021693f
C800 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 GNDA 0.025108f
C801 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t9 GNDA 0.021693f
C802 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t5 GNDA 0.021693f
C803 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 GNDA 0.025108f
C804 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t11 GNDA 0.021693f
C805 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t8 GNDA 0.021693f
C806 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 GNDA 0.025081f
C807 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 GNDA 0.047428f
C808 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 GNDA 0.148528f
C809 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t10 GNDA 0.021693f
C810 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t6 GNDA 0.021693f
C811 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 GNDA 0.043385f
C812 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 GNDA 1.17574f
C813 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t0 GNDA 0.032539f
C814 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t2 GNDA 0.032539f
C815 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 GNDA 0.07557f
C816 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t14 GNDA 0.057757f
C817 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t31 GNDA 0.057757f
C818 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t20 GNDA 0.057757f
C819 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t29 GNDA 0.057757f
C820 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t18 GNDA 0.057757f
C821 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t28 GNDA 0.057757f
C822 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t17 GNDA 0.057757f
C823 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t26 GNDA 0.057757f
C824 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t15 GNDA 0.057757f
C825 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t19 GNDA 0.067411f
C826 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 GNDA 0.063558f
C827 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 GNDA 0.03986f
C828 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 GNDA 0.03986f
C829 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 GNDA 0.03986f
C830 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 GNDA 0.03986f
C831 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 GNDA 0.03986f
C832 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 GNDA 0.03986f
C833 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 GNDA 0.03986f
C834 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 GNDA 0.035618f
C835 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t25 GNDA 0.057757f
C836 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t22 GNDA 0.057757f
C837 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t12 GNDA 0.057757f
C838 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t23 GNDA 0.057757f
C839 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t13 GNDA 0.057757f
C840 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t24 GNDA 0.057757f
C841 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t16 GNDA 0.057757f
C842 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t27 GNDA 0.057757f
C843 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t30 GNDA 0.057757f
C844 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t21 GNDA 0.067411f
C845 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 GNDA 0.063558f
C846 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 GNDA 0.03986f
C847 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 GNDA 0.03986f
C848 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 GNDA 0.03986f
C849 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 GNDA 0.03986f
C850 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 GNDA 0.03986f
C851 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 GNDA 0.03986f
C852 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 GNDA 0.03986f
C853 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 GNDA 0.035618f
C854 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 GNDA 0.030153f
C855 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 GNDA 0.455043f
C856 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t3 GNDA 0.032539f
C857 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t1 GNDA 0.032539f
C858 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 GNDA 0.070801f
C859 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 GNDA 0.319895f
C860 two_stage_opamp_dummy_magic_23_0.VD2.t8 GNDA 0.053331f
C861 two_stage_opamp_dummy_magic_23_0.VD2.t3 GNDA 0.053331f
C862 two_stage_opamp_dummy_magic_23_0.VD2.n0 GNDA 0.116042f
C863 two_stage_opamp_dummy_magic_23_0.VD2.n1 GNDA 0.361396f
C864 two_stage_opamp_dummy_magic_23_0.VD2.n2 GNDA 0.192793f
C865 two_stage_opamp_dummy_magic_23_0.VD2.t5 GNDA 0.053331f
C866 two_stage_opamp_dummy_magic_23_0.VD2.t1 GNDA 0.053331f
C867 two_stage_opamp_dummy_magic_23_0.VD2.n3 GNDA 0.116042f
C868 two_stage_opamp_dummy_magic_23_0.VD2.n4 GNDA 0.461069f
C869 two_stage_opamp_dummy_magic_23_0.VD2.t9 GNDA 0.053331f
C870 two_stage_opamp_dummy_magic_23_0.VD2.t4 GNDA 0.053331f
C871 two_stage_opamp_dummy_magic_23_0.VD2.n5 GNDA 0.116042f
C872 two_stage_opamp_dummy_magic_23_0.VD2.n6 GNDA 0.461069f
C873 two_stage_opamp_dummy_magic_23_0.VD2.t7 GNDA 0.053331f
C874 two_stage_opamp_dummy_magic_23_0.VD2.t10 GNDA 0.053331f
C875 two_stage_opamp_dummy_magic_23_0.VD2.n7 GNDA 0.116042f
C876 two_stage_opamp_dummy_magic_23_0.VD2.n8 GNDA 0.442486f
C877 two_stage_opamp_dummy_magic_23_0.VD2.n9 GNDA 0.203944f
C878 two_stage_opamp_dummy_magic_23_0.VD2.n10 GNDA 0.119128f
C879 two_stage_opamp_dummy_magic_23_0.VD2.n11 GNDA 0.203944f
C880 two_stage_opamp_dummy_magic_23_0.VD2.t6 GNDA 0.053331f
C881 two_stage_opamp_dummy_magic_23_0.VD2.t2 GNDA 0.053331f
C882 two_stage_opamp_dummy_magic_23_0.VD2.n12 GNDA 0.116042f
C883 two_stage_opamp_dummy_magic_23_0.VD2.n13 GNDA 0.442486f
C884 two_stage_opamp_dummy_magic_23_0.VD2.n14 GNDA 0.192793f
C885 two_stage_opamp_dummy_magic_23_0.VD2.n15 GNDA 0.106662f
C886 two_stage_opamp_dummy_magic_23_0.VD2.n16 GNDA 0.122513f
C887 two_stage_opamp_dummy_magic_23_0.VD2.n17 GNDA 0.099935f
C888 two_stage_opamp_dummy_magic_23_0.VD2.n18 GNDA 0.205342f
C889 two_stage_opamp_dummy_magic_23_0.VD2.t19 GNDA 0.053331f
C890 two_stage_opamp_dummy_magic_23_0.VD2.t21 GNDA 0.053331f
C891 two_stage_opamp_dummy_magic_23_0.VD2.n19 GNDA 0.116042f
C892 two_stage_opamp_dummy_magic_23_0.VD2.n20 GNDA 0.465721f
C893 two_stage_opamp_dummy_magic_23_0.VD2.n21 GNDA 0.205342f
C894 two_stage_opamp_dummy_magic_23_0.VD2.t11 GNDA 0.053331f
C895 two_stage_opamp_dummy_magic_23_0.VD2.t18 GNDA 0.053331f
C896 two_stage_opamp_dummy_magic_23_0.VD2.n22 GNDA 0.116042f
C897 two_stage_opamp_dummy_magic_23_0.VD2.n23 GNDA 0.447102f
C898 two_stage_opamp_dummy_magic_23_0.VD2.n24 GNDA 0.192793f
C899 two_stage_opamp_dummy_magic_23_0.VD2.t15 GNDA 0.053331f
C900 two_stage_opamp_dummy_magic_23_0.VD2.t14 GNDA 0.053331f
C901 two_stage_opamp_dummy_magic_23_0.VD2.n25 GNDA 0.116042f
C902 two_stage_opamp_dummy_magic_23_0.VD2.n26 GNDA 0.447102f
C903 two_stage_opamp_dummy_magic_23_0.VD2.n27 GNDA 0.113419f
C904 two_stage_opamp_dummy_magic_23_0.VD2.t16 GNDA 0.053331f
C905 two_stage_opamp_dummy_magic_23_0.VD2.t20 GNDA 0.053331f
C906 two_stage_opamp_dummy_magic_23_0.VD2.n28 GNDA 0.116042f
C907 two_stage_opamp_dummy_magic_23_0.VD2.n29 GNDA 0.465721f
C908 two_stage_opamp_dummy_magic_23_0.VD2.t12 GNDA 0.053331f
C909 two_stage_opamp_dummy_magic_23_0.VD2.t0 GNDA 0.053331f
C910 two_stage_opamp_dummy_magic_23_0.VD2.n30 GNDA 0.116042f
C911 two_stage_opamp_dummy_magic_23_0.VD2.n31 GNDA 0.447102f
C912 two_stage_opamp_dummy_magic_23_0.VD2.n32 GNDA 0.192793f
C913 two_stage_opamp_dummy_magic_23_0.VD2.n33 GNDA 0.113419f
C914 two_stage_opamp_dummy_magic_23_0.VD2.t17 GNDA 0.053331f
C915 two_stage_opamp_dummy_magic_23_0.VD2.t13 GNDA 0.053331f
C916 two_stage_opamp_dummy_magic_23_0.VD2.n34 GNDA 0.116042f
C917 two_stage_opamp_dummy_magic_23_0.VD2.n35 GNDA 0.447102f
C918 two_stage_opamp_dummy_magic_23_0.VD2.n36 GNDA 0.099935f
C919 two_stage_opamp_dummy_magic_23_0.VD2.n37 GNDA 0.06757f
C920 bgr_11_0.cap_res1.t14 GNDA 0.331712f
C921 bgr_11_0.cap_res1.t19 GNDA 0.349187f
C922 bgr_11_0.cap_res1.t17 GNDA 0.350452f
C923 bgr_11_0.cap_res1.t7 GNDA 0.331712f
C924 bgr_11_0.cap_res1.t16 GNDA 0.349187f
C925 bgr_11_0.cap_res1.t11 GNDA 0.350452f
C926 bgr_11_0.cap_res1.t1 GNDA 0.331712f
C927 bgr_11_0.cap_res1.t10 GNDA 0.349187f
C928 bgr_11_0.cap_res1.t3 GNDA 0.350452f
C929 bgr_11_0.cap_res1.t5 GNDA 0.331712f
C930 bgr_11_0.cap_res1.t15 GNDA 0.349187f
C931 bgr_11_0.cap_res1.t9 GNDA 0.350452f
C932 bgr_11_0.cap_res1.t20 GNDA 0.331712f
C933 bgr_11_0.cap_res1.t8 GNDA 0.349187f
C934 bgr_11_0.cap_res1.t2 GNDA 0.350452f
C935 bgr_11_0.cap_res1.n0 GNDA 0.23406f
C936 bgr_11_0.cap_res1.t4 GNDA 0.186395f
C937 bgr_11_0.cap_res1.n1 GNDA 0.253961f
C938 bgr_11_0.cap_res1.t12 GNDA 0.186395f
C939 bgr_11_0.cap_res1.n2 GNDA 0.253961f
C940 bgr_11_0.cap_res1.t6 GNDA 0.186395f
C941 bgr_11_0.cap_res1.n3 GNDA 0.253961f
C942 bgr_11_0.cap_res1.t13 GNDA 0.186395f
C943 bgr_11_0.cap_res1.n4 GNDA 0.253961f
C944 bgr_11_0.cap_res1.t18 GNDA 0.363549f
C945 bgr_11_0.cap_res1.t0 GNDA 0.08421f
C946 w_6100_17280.n0 GNDA 0.296479f
C947 w_6100_17280.n1 GNDA 0.388831f
C948 w_6100_17280.n2 GNDA 0.296479f
C949 w_6100_17280.n3 GNDA 0.296479f
C950 w_6100_17280.n4 GNDA 0.336948f
C951 w_6100_17280.n5 GNDA 0.336948f
C952 w_6100_17280.n6 GNDA 0.296479f
C953 w_6100_17280.n7 GNDA 0.296479f
C954 w_6100_17280.n8 GNDA 0.296479f
C955 w_6100_17280.n9 GNDA 0.388831f
C956 w_6100_17280.n10 GNDA 0.014102f
C957 w_6100_17280.n11 GNDA 0.014102f
C958 w_6100_17280.n12 GNDA 0.024006f
C959 w_6100_17280.n13 GNDA 0.024006f
C960 w_6100_17280.n14 GNDA 0.014102f
C961 w_6100_17280.n15 GNDA 0.014102f
C962 w_6100_17280.n16 GNDA 0.014102f
C963 w_6100_17280.n17 GNDA 0.014102f
C964 w_6100_17280.n18 GNDA 0.014102f
C965 w_6100_17280.n19 GNDA 0.014102f
C966 w_6100_17280.n20 GNDA 0.014102f
C967 w_6100_17280.n21 GNDA 0.014102f
C968 w_6100_17280.n22 GNDA 0.022473f
C969 w_6100_17280.t36 GNDA 0.020943f
C970 w_6100_17280.t38 GNDA 0.019744f
C971 w_6100_17280.n24 GNDA 0.037999f
C972 w_6100_17280.n25 GNDA 0.069969f
C973 w_6100_17280.t37 GNDA 0.058908f
C974 w_6100_17280.t74 GNDA 0.047681f
C975 w_6100_17280.t62 GNDA 0.047681f
C976 w_6100_17280.t34 GNDA 0.047681f
C977 w_6100_17280.t80 GNDA 0.047681f
C978 w_6100_17280.t48 GNDA 0.047681f
C979 w_6100_17280.t70 GNDA 0.047681f
C980 w_6100_17280.t66 GNDA 0.047681f
C981 w_6100_17280.t28 GNDA 0.047681f
C982 w_6100_17280.t2 GNDA 0.047681f
C983 w_6100_17280.t64 GNDA 0.047681f
C984 w_6100_17280.t82 GNDA 0.047681f
C985 w_6100_17280.t72 GNDA 0.047681f
C986 w_6100_17280.t68 GNDA 0.047681f
C987 w_6100_17280.t30 GNDA 0.047681f
C988 w_6100_17280.t78 GNDA 0.047681f
C989 w_6100_17280.t32 GNDA 0.047681f
C990 w_6100_17280.t0 GNDA 0.047681f
C991 w_6100_17280.t76 GNDA 0.047681f
C992 w_6100_17280.t43 GNDA 0.071347f
C993 w_6100_17280.n26 GNDA 0.05753f
C994 w_6100_17280.t44 GNDA 0.019744f
C995 w_6100_17280.n27 GNDA 0.037846f
C996 w_6100_17280.t42 GNDA 0.020954f
C997 w_6100_17280.n28 GNDA 0.021479f
C998 w_6100_17280.t41 GNDA 0.019882f
C999 w_6100_17280.n29 GNDA 0.024006f
C1000 w_6100_17280.n30 GNDA 0.014102f
C1001 w_6100_17280.n31 GNDA 0.014102f
C1002 w_6100_17280.n32 GNDA 0.014102f
C1003 w_6100_17280.n33 GNDA 0.014102f
C1004 w_6100_17280.n34 GNDA 0.022473f
C1005 w_6100_17280.t45 GNDA 0.020954f
C1006 w_6100_17280.t47 GNDA 0.019744f
C1007 w_6100_17280.n35 GNDA 0.037846f
C1008 w_6100_17280.n36 GNDA 0.05753f
C1009 w_6100_17280.t46 GNDA 0.071347f
C1010 w_6100_17280.t52 GNDA 0.047681f
C1011 w_6100_17280.t4 GNDA 0.047681f
C1012 w_6100_17280.t16 GNDA 0.047681f
C1013 w_6100_17280.t26 GNDA 0.047681f
C1014 w_6100_17280.t12 GNDA 0.047681f
C1015 w_6100_17280.t56 GNDA 0.047681f
C1016 w_6100_17280.t54 GNDA 0.047681f
C1017 w_6100_17280.t24 GNDA 0.047681f
C1018 w_6100_17280.t10 GNDA 0.047681f
C1019 w_6100_17280.t20 GNDA 0.047681f
C1020 w_6100_17280.t6 GNDA 0.047681f
C1021 w_6100_17280.t60 GNDA 0.047681f
C1022 w_6100_17280.t50 GNDA 0.047681f
C1023 w_6100_17280.t22 GNDA 0.047681f
C1024 w_6100_17280.t8 GNDA 0.047681f
C1025 w_6100_17280.t18 GNDA 0.047681f
C1026 w_6100_17280.t14 GNDA 0.047681f
C1027 w_6100_17280.t58 GNDA 0.047681f
C1028 w_6100_17280.t40 GNDA 0.07273f
C1029 w_6100_17280.n37 GNDA 0.103559f
C1030 w_6100_17280.t39 GNDA 0.014051f
C1031 w_6100_17280.n38 GNDA 0.02381f
C1032 w_6100_17280.n39 GNDA 0.014102f
C1033 w_6100_17280.n40 GNDA 0.014102f
C1034 w_6100_17280.n41 GNDA 0.014102f
C1035 w_6100_17280.n42 GNDA 0.014102f
C1036 bgr_11_0.1st_Vout_1.n0 GNDA 1.57339f
C1037 bgr_11_0.1st_Vout_1.n1 GNDA 0.470087f
C1038 bgr_11_0.1st_Vout_1.n2 GNDA 1.05551f
C1039 bgr_11_0.1st_Vout_1.n3 GNDA 0.105834f
C1040 bgr_11_0.1st_Vout_1.n4 GNDA 0.163342f
C1041 bgr_11_0.1st_Vout_1.t7 GNDA 0.312799f
C1042 bgr_11_0.1st_Vout_1.t29 GNDA 0.307561f
C1043 bgr_11_0.1st_Vout_1.t24 GNDA 0.312799f
C1044 bgr_11_0.1st_Vout_1.t31 GNDA 0.307561f
C1045 bgr_11_0.1st_Vout_1.t28 GNDA 0.312799f
C1046 bgr_11_0.1st_Vout_1.t18 GNDA 0.307561f
C1047 bgr_11_0.1st_Vout_1.t15 GNDA 0.312799f
C1048 bgr_11_0.1st_Vout_1.t22 GNDA 0.307561f
C1049 bgr_11_0.1st_Vout_1.t32 GNDA 0.312799f
C1050 bgr_11_0.1st_Vout_1.t27 GNDA 0.307561f
C1051 bgr_11_0.1st_Vout_1.t21 GNDA 0.312799f
C1052 bgr_11_0.1st_Vout_1.t30 GNDA 0.307561f
C1053 bgr_11_0.1st_Vout_1.t26 GNDA 0.312799f
C1054 bgr_11_0.1st_Vout_1.t17 GNDA 0.307561f
C1055 bgr_11_0.1st_Vout_1.t14 GNDA 0.312799f
C1056 bgr_11_0.1st_Vout_1.t20 GNDA 0.307561f
C1057 bgr_11_0.1st_Vout_1.t16 GNDA 0.312799f
C1058 bgr_11_0.1st_Vout_1.t11 GNDA 0.307561f
C1059 bgr_11_0.1st_Vout_1.t13 GNDA 0.307561f
C1060 bgr_11_0.1st_Vout_1.t8 GNDA 0.307561f
C1061 bgr_11_0.1st_Vout_1.t23 GNDA 0.020092f
C1062 bgr_11_0.1st_Vout_1.n5 GNDA 0.628306f
C1063 bgr_11_0.1st_Vout_1.n6 GNDA 0.019383f
C1064 bgr_11_0.1st_Vout_1.t12 GNDA 0.011713f
C1065 bgr_11_0.1st_Vout_1.t19 GNDA 0.011713f
C1066 bgr_11_0.1st_Vout_1.n7 GNDA 0.026058f
C1067 bgr_11_0.1st_Vout_1.t6 GNDA 0.104485f
C1068 bgr_11_0.1st_Vout_1.n8 GNDA 0.018579f
C1069 bgr_11_0.1st_Vout_1.n9 GNDA 0.11222f
C1070 bgr_11_0.1st_Vout_1.t9 GNDA 0.011713f
C1071 bgr_11_0.1st_Vout_1.t25 GNDA 0.011713f
C1072 bgr_11_0.1st_Vout_1.n10 GNDA 0.026058f
C1073 bgr_11_0.1st_Vout_1.n11 GNDA 0.019383f
C1074 bgr_11_0.1st_Vout_1.t10 GNDA 0.018385f
C1075 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 GNDA 0.343734f
C1076 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t65 GNDA 0.344881f
C1077 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 GNDA 0.185242f
C1078 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 GNDA 0.197802f
C1079 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t95 GNDA 0.343734f
C1080 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t100 GNDA 0.344881f
C1081 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 GNDA 0.185242f
C1082 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 GNDA 0.216311f
C1083 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 GNDA 0.343734f
C1084 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t80 GNDA 0.344881f
C1085 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 GNDA 0.185242f
C1086 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 GNDA 0.216311f
C1087 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 GNDA 0.343734f
C1088 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 GNDA 0.344881f
C1089 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 GNDA 0.185242f
C1090 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 GNDA 0.216311f
C1091 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t8 GNDA 0.343734f
C1092 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 GNDA 0.344881f
C1093 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 GNDA 0.36339f
C1094 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 GNDA 0.36339f
C1095 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 GNDA 0.185242f
C1096 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 GNDA 0.216311f
C1097 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 GNDA 0.343734f
C1098 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t75 GNDA 0.344881f
C1099 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 GNDA 0.36339f
C1100 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 GNDA 0.36339f
C1101 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 GNDA 0.185242f
C1102 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 GNDA 0.216311f
C1103 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 GNDA 0.344881f
C1104 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 GNDA 0.346131f
C1105 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t90 GNDA 0.344881f
C1106 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 GNDA 0.347585f
C1107 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 GNDA 0.378048f
C1108 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 GNDA 0.344881f
C1109 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 GNDA 0.346131f
C1110 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t94 GNDA 0.344881f
C1111 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 GNDA 0.346131f
C1112 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 GNDA 0.344881f
C1113 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 GNDA 0.346131f
C1114 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 GNDA 0.344881f
C1115 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 GNDA 0.346131f
C1116 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t52 GNDA 0.344881f
C1117 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 GNDA 0.346131f
C1118 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t27 GNDA 0.344881f
C1119 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 GNDA 0.346131f
C1120 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t21 GNDA 0.344881f
C1121 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 GNDA 0.346131f
C1122 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 GNDA 0.344881f
C1123 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 GNDA 0.346131f
C1124 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t59 GNDA 0.344881f
C1125 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 GNDA 0.346131f
C1126 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 GNDA 0.344881f
C1127 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 GNDA 0.346131f
C1128 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t99 GNDA 0.344881f
C1129 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 GNDA 0.346131f
C1130 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 GNDA 0.344881f
C1131 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 GNDA 0.346131f
C1132 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t67 GNDA 0.344881f
C1133 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 GNDA 0.346131f
C1134 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 GNDA 0.344881f
C1135 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 GNDA 0.346131f
C1136 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t104 GNDA 0.344881f
C1137 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 GNDA 0.346131f
C1138 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t76 GNDA 0.344881f
C1139 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 GNDA 0.346131f
C1140 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 GNDA 0.344881f
C1141 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 GNDA 0.346131f
C1142 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 GNDA 0.344881f
C1143 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 GNDA 0.346131f
C1144 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t109 GNDA 0.344881f
C1145 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 GNDA 0.346131f
C1146 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t82 GNDA 0.344881f
C1147 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 GNDA 0.346131f
C1148 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 GNDA 0.344881f
C1149 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 GNDA 0.346131f
C1150 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 GNDA 0.344881f
C1151 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 GNDA 0.346131f
C1152 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t47 GNDA 0.344881f
C1153 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 GNDA 0.346131f
C1154 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t20 GNDA 0.344881f
C1155 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 GNDA 0.346131f
C1156 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 GNDA 0.344881f
C1157 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 GNDA 0.346131f
C1158 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t58 GNDA 0.344881f
C1159 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 GNDA 0.346131f
C1160 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t53 GNDA 0.344881f
C1161 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 GNDA 0.346131f
C1162 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 GNDA 0.344881f
C1163 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 GNDA 0.346131f
C1164 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 GNDA 0.344881f
C1165 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 GNDA 0.36179f
C1166 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 GNDA 0.344881f
C1167 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 GNDA 0.185242f
C1168 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 GNDA 0.198255f
C1169 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 GNDA 0.344881f
C1170 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 GNDA 0.185242f
C1171 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 GNDA 0.196656f
C1172 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 GNDA 0.344881f
C1173 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 GNDA 0.185242f
C1174 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 GNDA 0.196656f
C1175 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 GNDA 0.344881f
C1176 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 GNDA 0.185242f
C1177 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 GNDA 0.196656f
C1178 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t31 GNDA 0.344881f
C1179 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 GNDA 0.185242f
C1180 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 GNDA 0.196656f
C1181 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 GNDA 0.344881f
C1182 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 GNDA 0.185242f
C1183 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 GNDA 0.196656f
C1184 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t113 GNDA 0.344881f
C1185 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 GNDA 0.185242f
C1186 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 GNDA 0.196656f
C1187 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 GNDA 0.344881f
C1188 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 GNDA 0.185242f
C1189 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 GNDA 0.196656f
C1190 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t57 GNDA 0.344881f
C1191 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 GNDA 0.185242f
C1192 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 GNDA 0.196656f
C1193 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t98 GNDA 0.344881f
C1194 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 GNDA 0.346131f
C1195 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 GNDA 0.344881f
C1196 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 GNDA 0.346131f
C1197 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 GNDA 0.166734f
C1198 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 GNDA 0.215061f
C1199 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 GNDA 0.184096f
C1200 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 GNDA 0.23357f
C1201 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 GNDA 0.184096f
C1202 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 GNDA 0.250829f
C1203 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 GNDA 0.184096f
C1204 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 GNDA 0.250829f
C1205 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 GNDA 0.184096f
C1206 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 GNDA 0.250829f
C1207 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 GNDA 0.184096f
C1208 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 GNDA 0.250829f
C1209 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 GNDA 0.184096f
C1210 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 GNDA 0.250829f
C1211 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 GNDA 0.184096f
C1212 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 GNDA 0.250829f
C1213 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 GNDA 0.184096f
C1214 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 GNDA 0.250829f
C1215 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 GNDA 0.184096f
C1216 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 GNDA 0.250829f
C1217 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 GNDA 0.184096f
C1218 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 GNDA 0.250829f
C1219 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 GNDA 0.184096f
C1220 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 GNDA 0.250829f
C1221 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 GNDA 0.184096f
C1222 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 GNDA 0.250829f
C1223 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 GNDA 0.184096f
C1224 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 GNDA 0.250829f
C1225 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 GNDA 0.184096f
C1226 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 GNDA 0.250829f
C1227 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 GNDA 0.184096f
C1228 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 GNDA 0.250829f
C1229 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 GNDA 0.184096f
C1230 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 GNDA 0.23357f
C1231 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t81 GNDA 0.343734f
C1232 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 GNDA 0.166734f
C1233 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 GNDA 0.216311f
C1234 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 GNDA 0.343734f
C1235 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 GNDA 0.166734f
C1236 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 GNDA 0.216311f
C1237 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t66 GNDA 0.343734f
C1238 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 GNDA 0.344881f
C1239 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 GNDA 0.36339f
C1240 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 GNDA 0.36339f
C1241 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 GNDA 0.185242f
C1242 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 GNDA 0.216311f
C1243 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 GNDA 0.343734f
C1244 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 GNDA 0.216311f
C1245 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 GNDA 0.185242f
C1246 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 GNDA 0.36339f
C1247 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 GNDA 0.36339f
C1248 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 GNDA 0.434792f
C1249 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 GNDA 0.291879f
C1250 two_stage_opamp_dummy_magic_23_0.VD3.t13 GNDA 0.060837f
C1251 two_stage_opamp_dummy_magic_23_0.VD3.t23 GNDA 0.060837f
C1252 two_stage_opamp_dummy_magic_23_0.VD3.t29 GNDA 0.060837f
C1253 two_stage_opamp_dummy_magic_23_0.VD3.n0 GNDA 0.154422f
C1254 two_stage_opamp_dummy_magic_23_0.VD3.n1 GNDA 0.43135f
C1255 two_stage_opamp_dummy_magic_23_0.VD3.t35 GNDA 0.106675f
C1256 two_stage_opamp_dummy_magic_23_0.VD3.t34 GNDA 0.216405f
C1257 two_stage_opamp_dummy_magic_23_0.VD3.n2 GNDA 0.065988f
C1258 two_stage_opamp_dummy_magic_23_0.VD3.n3 GNDA 0.065988f
C1259 two_stage_opamp_dummy_magic_23_0.VD3.t10 GNDA 0.060837f
C1260 two_stage_opamp_dummy_magic_23_0.VD3.t3 GNDA 0.060837f
C1261 two_stage_opamp_dummy_magic_23_0.VD3.n4 GNDA 0.124448f
C1262 two_stage_opamp_dummy_magic_23_0.VD3.n5 GNDA 0.402926f
C1263 two_stage_opamp_dummy_magic_23_0.VD3.n6 GNDA 0.112569f
C1264 two_stage_opamp_dummy_magic_23_0.VD3.t1 GNDA 0.060837f
C1265 two_stage_opamp_dummy_magic_23_0.VD3.t4 GNDA 0.060837f
C1266 two_stage_opamp_dummy_magic_23_0.VD3.n7 GNDA 0.124448f
C1267 two_stage_opamp_dummy_magic_23_0.VD3.n8 GNDA 0.391923f
C1268 two_stage_opamp_dummy_magic_23_0.VD3.n9 GNDA 0.112569f
C1269 two_stage_opamp_dummy_magic_23_0.VD3.t6 GNDA 0.060837f
C1270 two_stage_opamp_dummy_magic_23_0.VD3.t8 GNDA 0.060837f
C1271 two_stage_opamp_dummy_magic_23_0.VD3.n10 GNDA 0.124448f
C1272 two_stage_opamp_dummy_magic_23_0.VD3.n11 GNDA 0.391923f
C1273 two_stage_opamp_dummy_magic_23_0.VD3.n12 GNDA 0.065988f
C1274 two_stage_opamp_dummy_magic_23_0.VD3.n13 GNDA 0.065988f
C1275 two_stage_opamp_dummy_magic_23_0.VD3.t9 GNDA 0.060837f
C1276 two_stage_opamp_dummy_magic_23_0.VD3.t0 GNDA 0.060837f
C1277 two_stage_opamp_dummy_magic_23_0.VD3.n14 GNDA 0.124448f
C1278 two_stage_opamp_dummy_magic_23_0.VD3.n15 GNDA 0.391923f
C1279 two_stage_opamp_dummy_magic_23_0.VD3.n16 GNDA 0.065988f
C1280 two_stage_opamp_dummy_magic_23_0.VD3.t2 GNDA 0.060837f
C1281 two_stage_opamp_dummy_magic_23_0.VD3.t5 GNDA 0.060837f
C1282 two_stage_opamp_dummy_magic_23_0.VD3.n17 GNDA 0.124448f
C1283 two_stage_opamp_dummy_magic_23_0.VD3.n18 GNDA 0.391923f
C1284 two_stage_opamp_dummy_magic_23_0.VD3.n19 GNDA 0.112569f
C1285 two_stage_opamp_dummy_magic_23_0.VD3.t7 GNDA 0.060837f
C1286 two_stage_opamp_dummy_magic_23_0.VD3.t11 GNDA 0.060837f
C1287 two_stage_opamp_dummy_magic_23_0.VD3.n20 GNDA 0.124448f
C1288 two_stage_opamp_dummy_magic_23_0.VD3.n21 GNDA 0.397425f
C1289 two_stage_opamp_dummy_magic_23_0.VD3.n22 GNDA 0.257485f
C1290 two_stage_opamp_dummy_magic_23_0.VD3.t21 GNDA 0.060837f
C1291 two_stage_opamp_dummy_magic_23_0.VD3.t27 GNDA 0.060837f
C1292 two_stage_opamp_dummy_magic_23_0.VD3.n23 GNDA 0.154422f
C1293 two_stage_opamp_dummy_magic_23_0.VD3.n24 GNDA 0.43135f
C1294 two_stage_opamp_dummy_magic_23_0.VD3.n25 GNDA 0.2193f
C1295 two_stage_opamp_dummy_magic_23_0.VD3.t32 GNDA 0.106675f
C1296 two_stage_opamp_dummy_magic_23_0.VD3.n26 GNDA 0.311214f
C1297 two_stage_opamp_dummy_magic_23_0.VD3.n27 GNDA 0.627773f
C1298 two_stage_opamp_dummy_magic_23_0.VD3.t33 GNDA 0.518568f
C1299 two_stage_opamp_dummy_magic_23_0.VD3.t20 GNDA 0.406738f
C1300 two_stage_opamp_dummy_magic_23_0.VD3.t26 GNDA 0.406738f
C1301 two_stage_opamp_dummy_magic_23_0.VD3.t22 GNDA 0.406738f
C1302 two_stage_opamp_dummy_magic_23_0.VD3.t28 GNDA 0.402972f
C1303 two_stage_opamp_dummy_magic_23_0.VD3.t30 GNDA 0.399206f
C1304 two_stage_opamp_dummy_magic_23_0.VD3.t12 GNDA 0.406738f
C1305 two_stage_opamp_dummy_magic_23_0.VD3.t16 GNDA 0.406738f
C1306 two_stage_opamp_dummy_magic_23_0.VD3.t14 GNDA 0.406738f
C1307 two_stage_opamp_dummy_magic_23_0.VD3.t18 GNDA 0.406738f
C1308 two_stage_opamp_dummy_magic_23_0.VD3.t24 GNDA 0.406738f
C1309 two_stage_opamp_dummy_magic_23_0.VD3.t36 GNDA 0.518568f
C1310 two_stage_opamp_dummy_magic_23_0.VD3.t37 GNDA 0.216405f
C1311 two_stage_opamp_dummy_magic_23_0.VD3.n28 GNDA 0.627773f
C1312 two_stage_opamp_dummy_magic_23_0.VD3.n29 GNDA 0.316969f
C1313 two_stage_opamp_dummy_magic_23_0.VD3.t19 GNDA 0.060837f
C1314 two_stage_opamp_dummy_magic_23_0.VD3.t25 GNDA 0.060837f
C1315 two_stage_opamp_dummy_magic_23_0.VD3.n30 GNDA 0.154422f
C1316 two_stage_opamp_dummy_magic_23_0.VD3.n31 GNDA 0.481799f
C1317 two_stage_opamp_dummy_magic_23_0.VD3.t17 GNDA 0.060837f
C1318 two_stage_opamp_dummy_magic_23_0.VD3.t15 GNDA 0.060837f
C1319 two_stage_opamp_dummy_magic_23_0.VD3.n32 GNDA 0.154422f
C1320 two_stage_opamp_dummy_magic_23_0.VD3.n33 GNDA 0.43135f
C1321 two_stage_opamp_dummy_magic_23_0.VD3.n34 GNDA 0.43135f
C1322 two_stage_opamp_dummy_magic_23_0.VD3.n35 GNDA 0.154422f
C1323 two_stage_opamp_dummy_magic_23_0.VD3.t31 GNDA 0.060837f
C1324 two_stage_opamp_dummy_magic_23_0.Vb2.t10 GNDA 0.05533f
C1325 two_stage_opamp_dummy_magic_23_0.Vb2.t0 GNDA 0.05533f
C1326 two_stage_opamp_dummy_magic_23_0.Vb2.n0 GNDA 0.117497f
C1327 two_stage_opamp_dummy_magic_23_0.Vb2.t9 GNDA 0.103286f
C1328 two_stage_opamp_dummy_magic_23_0.Vb2.n1 GNDA 0.478278f
C1329 two_stage_opamp_dummy_magic_23_0.Vb2.t31 GNDA 0.062028f
C1330 two_stage_opamp_dummy_magic_23_0.Vb2.n2 GNDA 0.238127f
C1331 two_stage_opamp_dummy_magic_23_0.Vb2.t28 GNDA 0.078252f
C1332 two_stage_opamp_dummy_magic_23_0.Vb2.t23 GNDA 0.078252f
C1333 two_stage_opamp_dummy_magic_23_0.Vb2.t26 GNDA 0.078252f
C1334 two_stage_opamp_dummy_magic_23_0.Vb2.t21 GNDA 0.078252f
C1335 two_stage_opamp_dummy_magic_23_0.Vb2.t16 GNDA 0.090303f
C1336 two_stage_opamp_dummy_magic_23_0.Vb2.n3 GNDA 0.073316f
C1337 two_stage_opamp_dummy_magic_23_0.Vb2.n4 GNDA 0.045054f
C1338 two_stage_opamp_dummy_magic_23_0.Vb2.n5 GNDA 0.045054f
C1339 two_stage_opamp_dummy_magic_23_0.Vb2.n6 GNDA 0.039504f
C1340 two_stage_opamp_dummy_magic_23_0.Vb2.t11 GNDA 0.078252f
C1341 two_stage_opamp_dummy_magic_23_0.Vb2.t13 GNDA 0.078252f
C1342 two_stage_opamp_dummy_magic_23_0.Vb2.t17 GNDA 0.078252f
C1343 two_stage_opamp_dummy_magic_23_0.Vb2.t14 GNDA 0.078252f
C1344 two_stage_opamp_dummy_magic_23_0.Vb2.t19 GNDA 0.090303f
C1345 two_stage_opamp_dummy_magic_23_0.Vb2.n7 GNDA 0.073316f
C1346 two_stage_opamp_dummy_magic_23_0.Vb2.n8 GNDA 0.045054f
C1347 two_stage_opamp_dummy_magic_23_0.Vb2.n9 GNDA 0.045054f
C1348 two_stage_opamp_dummy_magic_23_0.Vb2.n10 GNDA 0.039504f
C1349 two_stage_opamp_dummy_magic_23_0.Vb2.n11 GNDA 0.029278f
C1350 two_stage_opamp_dummy_magic_23_0.Vb2.t32 GNDA 0.078252f
C1351 two_stage_opamp_dummy_magic_23_0.Vb2.t29 GNDA 0.078252f
C1352 two_stage_opamp_dummy_magic_23_0.Vb2.t25 GNDA 0.078252f
C1353 two_stage_opamp_dummy_magic_23_0.Vb2.t20 GNDA 0.078252f
C1354 two_stage_opamp_dummy_magic_23_0.Vb2.t24 GNDA 0.090303f
C1355 two_stage_opamp_dummy_magic_23_0.Vb2.n12 GNDA 0.073316f
C1356 two_stage_opamp_dummy_magic_23_0.Vb2.n13 GNDA 0.045054f
C1357 two_stage_opamp_dummy_magic_23_0.Vb2.n14 GNDA 0.045054f
C1358 two_stage_opamp_dummy_magic_23_0.Vb2.n15 GNDA 0.039504f
C1359 two_stage_opamp_dummy_magic_23_0.Vb2.t12 GNDA 0.078252f
C1360 two_stage_opamp_dummy_magic_23_0.Vb2.t18 GNDA 0.078252f
C1361 two_stage_opamp_dummy_magic_23_0.Vb2.t22 GNDA 0.078252f
C1362 two_stage_opamp_dummy_magic_23_0.Vb2.t27 GNDA 0.078252f
C1363 two_stage_opamp_dummy_magic_23_0.Vb2.t30 GNDA 0.090303f
C1364 two_stage_opamp_dummy_magic_23_0.Vb2.n16 GNDA 0.073316f
C1365 two_stage_opamp_dummy_magic_23_0.Vb2.n17 GNDA 0.045054f
C1366 two_stage_opamp_dummy_magic_23_0.Vb2.n18 GNDA 0.045054f
C1367 two_stage_opamp_dummy_magic_23_0.Vb2.n19 GNDA 0.039504f
C1368 two_stage_opamp_dummy_magic_23_0.Vb2.n20 GNDA 0.028848f
C1369 two_stage_opamp_dummy_magic_23_0.Vb2.n21 GNDA 0.628828f
C1370 two_stage_opamp_dummy_magic_23_0.Vb2.n22 GNDA 0.293265f
C1371 two_stage_opamp_dummy_magic_23_0.Vb2.t15 GNDA 0.101693f
C1372 two_stage_opamp_dummy_magic_23_0.Vb2.n23 GNDA 1.46665f
C1373 two_stage_opamp_dummy_magic_23_0.Vb2.t8 GNDA 0.015809f
C1374 two_stage_opamp_dummy_magic_23_0.Vb2.t4 GNDA 0.015809f
C1375 two_stage_opamp_dummy_magic_23_0.Vb2.n24 GNDA 0.05155f
C1376 two_stage_opamp_dummy_magic_23_0.Vb2.n25 GNDA 1.60272f
C1377 two_stage_opamp_dummy_magic_23_0.Vb2.t1 GNDA 0.015809f
C1378 two_stage_opamp_dummy_magic_23_0.Vb2.t5 GNDA 0.015809f
C1379 two_stage_opamp_dummy_magic_23_0.Vb2.n26 GNDA 0.05155f
C1380 two_stage_opamp_dummy_magic_23_0.Vb2.n27 GNDA 0.308885f
C1381 two_stage_opamp_dummy_magic_23_0.Vb2.t2 GNDA 0.015809f
C1382 two_stage_opamp_dummy_magic_23_0.Vb2.t7 GNDA 0.015809f
C1383 two_stage_opamp_dummy_magic_23_0.Vb2.n28 GNDA 0.053004f
C1384 two_stage_opamp_dummy_magic_23_0.Vb2.n29 GNDA 0.470878f
C1385 two_stage_opamp_dummy_magic_23_0.Vb2.t3 GNDA 0.015809f
C1386 two_stage_opamp_dummy_magic_23_0.Vb2.n30 GNDA 0.05155f
C1387 two_stage_opamp_dummy_magic_23_0.Vb2.t6 GNDA 0.015809f
C1388 two_stage_opamp_dummy_magic_23_0.VD1.t6 GNDA 0.053331f
C1389 two_stage_opamp_dummy_magic_23_0.VD1.n0 GNDA 0.203944f
C1390 two_stage_opamp_dummy_magic_23_0.VD1.t7 GNDA 0.053331f
C1391 two_stage_opamp_dummy_magic_23_0.VD1.t2 GNDA 0.053331f
C1392 two_stage_opamp_dummy_magic_23_0.VD1.n1 GNDA 0.116042f
C1393 two_stage_opamp_dummy_magic_23_0.VD1.n2 GNDA 0.461069f
C1394 two_stage_opamp_dummy_magic_23_0.VD1.n3 GNDA 0.192793f
C1395 two_stage_opamp_dummy_magic_23_0.VD1.t3 GNDA 0.053331f
C1396 two_stage_opamp_dummy_magic_23_0.VD1.t8 GNDA 0.053331f
C1397 two_stage_opamp_dummy_magic_23_0.VD1.n4 GNDA 0.116042f
C1398 two_stage_opamp_dummy_magic_23_0.VD1.n5 GNDA 0.461069f
C1399 two_stage_opamp_dummy_magic_23_0.VD1.t5 GNDA 0.053331f
C1400 two_stage_opamp_dummy_magic_23_0.VD1.t9 GNDA 0.053331f
C1401 two_stage_opamp_dummy_magic_23_0.VD1.n6 GNDA 0.116042f
C1402 two_stage_opamp_dummy_magic_23_0.VD1.n7 GNDA 0.442486f
C1403 two_stage_opamp_dummy_magic_23_0.VD1.n8 GNDA 0.203944f
C1404 two_stage_opamp_dummy_magic_23_0.VD1.n9 GNDA 0.119128f
C1405 two_stage_opamp_dummy_magic_23_0.VD1.t4 GNDA 0.053331f
C1406 two_stage_opamp_dummy_magic_23_0.VD1.t1 GNDA 0.053331f
C1407 two_stage_opamp_dummy_magic_23_0.VD1.n10 GNDA 0.116042f
C1408 two_stage_opamp_dummy_magic_23_0.VD1.n11 GNDA 0.361396f
C1409 two_stage_opamp_dummy_magic_23_0.VD1.n12 GNDA 0.099935f
C1410 two_stage_opamp_dummy_magic_23_0.VD1.n13 GNDA 0.205342f
C1411 two_stage_opamp_dummy_magic_23_0.VD1.t20 GNDA 0.053331f
C1412 two_stage_opamp_dummy_magic_23_0.VD1.t15 GNDA 0.053331f
C1413 two_stage_opamp_dummy_magic_23_0.VD1.n14 GNDA 0.116042f
C1414 two_stage_opamp_dummy_magic_23_0.VD1.n15 GNDA 0.465721f
C1415 two_stage_opamp_dummy_magic_23_0.VD1.n16 GNDA 0.205342f
C1416 two_stage_opamp_dummy_magic_23_0.VD1.t14 GNDA 0.053331f
C1417 two_stage_opamp_dummy_magic_23_0.VD1.t16 GNDA 0.053331f
C1418 two_stage_opamp_dummy_magic_23_0.VD1.n17 GNDA 0.116042f
C1419 two_stage_opamp_dummy_magic_23_0.VD1.n18 GNDA 0.447102f
C1420 two_stage_opamp_dummy_magic_23_0.VD1.n19 GNDA 0.192793f
C1421 two_stage_opamp_dummy_magic_23_0.VD1.t21 GNDA 0.053331f
C1422 two_stage_opamp_dummy_magic_23_0.VD1.t18 GNDA 0.053331f
C1423 two_stage_opamp_dummy_magic_23_0.VD1.n20 GNDA 0.116042f
C1424 two_stage_opamp_dummy_magic_23_0.VD1.n21 GNDA 0.447102f
C1425 two_stage_opamp_dummy_magic_23_0.VD1.n22 GNDA 0.113419f
C1426 two_stage_opamp_dummy_magic_23_0.VD1.t13 GNDA 0.053331f
C1427 two_stage_opamp_dummy_magic_23_0.VD1.t19 GNDA 0.053331f
C1428 two_stage_opamp_dummy_magic_23_0.VD1.n23 GNDA 0.116042f
C1429 two_stage_opamp_dummy_magic_23_0.VD1.n24 GNDA 0.465721f
C1430 two_stage_opamp_dummy_magic_23_0.VD1.t0 GNDA 0.053331f
C1431 two_stage_opamp_dummy_magic_23_0.VD1.t12 GNDA 0.053331f
C1432 two_stage_opamp_dummy_magic_23_0.VD1.n25 GNDA 0.116042f
C1433 two_stage_opamp_dummy_magic_23_0.VD1.n26 GNDA 0.447102f
C1434 two_stage_opamp_dummy_magic_23_0.VD1.n27 GNDA 0.192793f
C1435 two_stage_opamp_dummy_magic_23_0.VD1.n28 GNDA 0.113419f
C1436 two_stage_opamp_dummy_magic_23_0.VD1.t11 GNDA 0.053331f
C1437 two_stage_opamp_dummy_magic_23_0.VD1.t17 GNDA 0.053331f
C1438 two_stage_opamp_dummy_magic_23_0.VD1.n29 GNDA 0.116042f
C1439 two_stage_opamp_dummy_magic_23_0.VD1.n30 GNDA 0.447102f
C1440 two_stage_opamp_dummy_magic_23_0.VD1.n31 GNDA 0.099935f
C1441 two_stage_opamp_dummy_magic_23_0.VD1.n32 GNDA 0.08441f
C1442 two_stage_opamp_dummy_magic_23_0.VD1.n33 GNDA 0.235249f
C1443 two_stage_opamp_dummy_magic_23_0.VD1.n34 GNDA 0.106662f
C1444 two_stage_opamp_dummy_magic_23_0.VD1.n35 GNDA 0.192793f
C1445 two_stage_opamp_dummy_magic_23_0.VD1.n36 GNDA 0.442486f
C1446 two_stage_opamp_dummy_magic_23_0.VD1.n37 GNDA 0.116042f
C1447 two_stage_opamp_dummy_magic_23_0.VD1.t10 GNDA 0.053331f
C1448 two_stage_opamp_dummy_magic_23_0.X.t4 GNDA 0.038289f
C1449 two_stage_opamp_dummy_magic_23_0.X.t10 GNDA 0.038289f
C1450 two_stage_opamp_dummy_magic_23_0.X.n0 GNDA 0.083312f
C1451 two_stage_opamp_dummy_magic_23_0.X.n1 GNDA 0.259463f
C1452 two_stage_opamp_dummy_magic_23_0.X.n2 GNDA 0.138415f
C1453 two_stage_opamp_dummy_magic_23_0.X.n3 GNDA 0.138415f
C1454 two_stage_opamp_dummy_magic_23_0.X.t24 GNDA 0.038289f
C1455 two_stage_opamp_dummy_magic_23_0.X.t13 GNDA 0.038289f
C1456 two_stage_opamp_dummy_magic_23_0.X.n4 GNDA 0.083312f
C1457 two_stage_opamp_dummy_magic_23_0.X.n5 GNDA 0.331023f
C1458 two_stage_opamp_dummy_magic_23_0.X.t8 GNDA 0.038289f
C1459 two_stage_opamp_dummy_magic_23_0.X.t12 GNDA 0.038289f
C1460 two_stage_opamp_dummy_magic_23_0.X.n6 GNDA 0.083312f
C1461 two_stage_opamp_dummy_magic_23_0.X.n7 GNDA 0.317681f
C1462 two_stage_opamp_dummy_magic_23_0.X.n8 GNDA 0.146421f
C1463 two_stage_opamp_dummy_magic_23_0.X.n9 GNDA 0.085527f
C1464 two_stage_opamp_dummy_magic_23_0.X.t5 GNDA 0.038289f
C1465 two_stage_opamp_dummy_magic_23_0.X.t23 GNDA 0.038289f
C1466 two_stage_opamp_dummy_magic_23_0.X.n10 GNDA 0.083312f
C1467 two_stage_opamp_dummy_magic_23_0.X.n11 GNDA 0.331023f
C1468 two_stage_opamp_dummy_magic_23_0.X.t6 GNDA 0.038289f
C1469 two_stage_opamp_dummy_magic_23_0.X.t9 GNDA 0.038289f
C1470 two_stage_opamp_dummy_magic_23_0.X.n12 GNDA 0.083312f
C1471 two_stage_opamp_dummy_magic_23_0.X.n13 GNDA 0.317681f
C1472 two_stage_opamp_dummy_magic_23_0.X.n14 GNDA 0.146421f
C1473 two_stage_opamp_dummy_magic_23_0.X.n15 GNDA 0.085527f
C1474 two_stage_opamp_dummy_magic_23_0.X.t7 GNDA 0.038289f
C1475 two_stage_opamp_dummy_magic_23_0.X.t11 GNDA 0.038289f
C1476 two_stage_opamp_dummy_magic_23_0.X.n16 GNDA 0.083312f
C1477 two_stage_opamp_dummy_magic_23_0.X.n17 GNDA 0.317681f
C1478 two_stage_opamp_dummy_magic_23_0.X.n18 GNDA 0.081429f
C1479 two_stage_opamp_dummy_magic_23_0.X.n19 GNDA 0.076577f
C1480 two_stage_opamp_dummy_magic_23_0.X.n20 GNDA 0.145807f
C1481 two_stage_opamp_dummy_magic_23_0.X.t3 GNDA 1.22341f
C1482 two_stage_opamp_dummy_magic_23_0.X.t34 GNDA 0.16847f
C1483 two_stage_opamp_dummy_magic_23_0.X.t51 GNDA 0.16847f
C1484 two_stage_opamp_dummy_magic_23_0.X.t37 GNDA 0.16847f
C1485 two_stage_opamp_dummy_magic_23_0.X.t53 GNDA 0.16847f
C1486 two_stage_opamp_dummy_magic_23_0.X.t36 GNDA 0.16847f
C1487 two_stage_opamp_dummy_magic_23_0.X.t52 GNDA 0.16847f
C1488 two_stage_opamp_dummy_magic_23_0.X.t39 GNDA 0.179433f
C1489 two_stage_opamp_dummy_magic_23_0.X.n21 GNDA 0.142193f
C1490 two_stage_opamp_dummy_magic_23_0.X.n22 GNDA 0.080406f
C1491 two_stage_opamp_dummy_magic_23_0.X.n23 GNDA 0.080406f
C1492 two_stage_opamp_dummy_magic_23_0.X.n24 GNDA 0.080406f
C1493 two_stage_opamp_dummy_magic_23_0.X.n25 GNDA 0.080406f
C1494 two_stage_opamp_dummy_magic_23_0.X.n26 GNDA 0.07227f
C1495 two_stage_opamp_dummy_magic_23_0.X.t48 GNDA 0.16847f
C1496 two_stage_opamp_dummy_magic_23_0.X.t31 GNDA 0.16847f
C1497 two_stage_opamp_dummy_magic_23_0.X.t46 GNDA 0.179433f
C1498 two_stage_opamp_dummy_magic_23_0.X.n27 GNDA 0.142193f
C1499 two_stage_opamp_dummy_magic_23_0.X.n28 GNDA 0.07227f
C1500 two_stage_opamp_dummy_magic_23_0.X.n29 GNDA 0.036557f
C1501 two_stage_opamp_dummy_magic_23_0.X.n30 GNDA 1.2754f
C1502 two_stage_opamp_dummy_magic_23_0.X.t15 GNDA 0.08934f
C1503 two_stage_opamp_dummy_magic_23_0.X.t17 GNDA 0.08934f
C1504 two_stage_opamp_dummy_magic_23_0.X.n31 GNDA 0.182755f
C1505 two_stage_opamp_dummy_magic_23_0.X.n32 GNDA 0.497099f
C1506 two_stage_opamp_dummy_magic_23_0.X.n33 GNDA 0.096905f
C1507 two_stage_opamp_dummy_magic_23_0.X.n34 GNDA 0.16531f
C1508 two_stage_opamp_dummy_magic_23_0.X.t18 GNDA 0.08934f
C1509 two_stage_opamp_dummy_magic_23_0.X.t20 GNDA 0.08934f
C1510 two_stage_opamp_dummy_magic_23_0.X.n35 GNDA 0.182755f
C1511 two_stage_opamp_dummy_magic_23_0.X.n36 GNDA 0.591707f
C1512 two_stage_opamp_dummy_magic_23_0.X.t0 GNDA 0.08934f
C1513 two_stage_opamp_dummy_magic_23_0.X.t21 GNDA 0.08934f
C1514 two_stage_opamp_dummy_magic_23_0.X.n37 GNDA 0.182755f
C1515 two_stage_opamp_dummy_magic_23_0.X.n38 GNDA 0.575548f
C1516 two_stage_opamp_dummy_magic_23_0.X.n39 GNDA 0.16531f
C1517 two_stage_opamp_dummy_magic_23_0.X.n40 GNDA 0.096905f
C1518 two_stage_opamp_dummy_magic_23_0.X.t16 GNDA 0.08934f
C1519 two_stage_opamp_dummy_magic_23_0.X.t22 GNDA 0.08934f
C1520 two_stage_opamp_dummy_magic_23_0.X.n41 GNDA 0.182755f
C1521 two_stage_opamp_dummy_magic_23_0.X.n42 GNDA 0.575548f
C1522 two_stage_opamp_dummy_magic_23_0.X.n43 GNDA 0.096905f
C1523 two_stage_opamp_dummy_magic_23_0.X.t1 GNDA 0.08934f
C1524 two_stage_opamp_dummy_magic_23_0.X.t14 GNDA 0.08934f
C1525 two_stage_opamp_dummy_magic_23_0.X.n44 GNDA 0.182755f
C1526 two_stage_opamp_dummy_magic_23_0.X.n45 GNDA 0.575548f
C1527 two_stage_opamp_dummy_magic_23_0.X.n46 GNDA 0.096905f
C1528 two_stage_opamp_dummy_magic_23_0.X.n47 GNDA 0.16531f
C1529 two_stage_opamp_dummy_magic_23_0.X.t2 GNDA 0.08934f
C1530 two_stage_opamp_dummy_magic_23_0.X.t19 GNDA 0.08934f
C1531 two_stage_opamp_dummy_magic_23_0.X.n48 GNDA 0.182755f
C1532 two_stage_opamp_dummy_magic_23_0.X.n49 GNDA 0.575548f
C1533 two_stage_opamp_dummy_magic_23_0.X.n50 GNDA 0.150696f
C1534 two_stage_opamp_dummy_magic_23_0.X.n51 GNDA 0.491162f
C1535 two_stage_opamp_dummy_magic_23_0.X.t44 GNDA 0.053604f
C1536 two_stage_opamp_dummy_magic_23_0.X.t30 GNDA 0.065091f
C1537 two_stage_opamp_dummy_magic_23_0.X.n52 GNDA 0.056954f
C1538 two_stage_opamp_dummy_magic_23_0.X.t27 GNDA 0.053604f
C1539 two_stage_opamp_dummy_magic_23_0.X.t45 GNDA 0.053604f
C1540 two_stage_opamp_dummy_magic_23_0.X.t28 GNDA 0.053604f
C1541 two_stage_opamp_dummy_magic_23_0.X.t42 GNDA 0.053604f
C1542 two_stage_opamp_dummy_magic_23_0.X.t25 GNDA 0.053604f
C1543 two_stage_opamp_dummy_magic_23_0.X.t40 GNDA 0.053604f
C1544 two_stage_opamp_dummy_magic_23_0.X.t54 GNDA 0.053604f
C1545 two_stage_opamp_dummy_magic_23_0.X.t38 GNDA 0.065091f
C1546 two_stage_opamp_dummy_magic_23_0.X.n53 GNDA 0.065091f
C1547 two_stage_opamp_dummy_magic_23_0.X.n54 GNDA 0.042118f
C1548 two_stage_opamp_dummy_magic_23_0.X.n55 GNDA 0.042118f
C1549 two_stage_opamp_dummy_magic_23_0.X.n56 GNDA 0.042118f
C1550 two_stage_opamp_dummy_magic_23_0.X.n57 GNDA 0.042118f
C1551 two_stage_opamp_dummy_magic_23_0.X.n58 GNDA 0.042118f
C1552 two_stage_opamp_dummy_magic_23_0.X.n59 GNDA 0.033981f
C1553 two_stage_opamp_dummy_magic_23_0.X.n60 GNDA 0.021431f
C1554 two_stage_opamp_dummy_magic_23_0.X.t49 GNDA 0.082321f
C1555 two_stage_opamp_dummy_magic_23_0.X.t35 GNDA 0.093585f
C1556 two_stage_opamp_dummy_magic_23_0.X.n61 GNDA 0.076321f
C1557 two_stage_opamp_dummy_magic_23_0.X.t32 GNDA 0.082321f
C1558 two_stage_opamp_dummy_magic_23_0.X.t50 GNDA 0.082321f
C1559 two_stage_opamp_dummy_magic_23_0.X.t33 GNDA 0.082321f
C1560 two_stage_opamp_dummy_magic_23_0.X.t47 GNDA 0.082321f
C1561 two_stage_opamp_dummy_magic_23_0.X.t29 GNDA 0.082321f
C1562 two_stage_opamp_dummy_magic_23_0.X.t43 GNDA 0.082321f
C1563 two_stage_opamp_dummy_magic_23_0.X.t26 GNDA 0.082321f
C1564 two_stage_opamp_dummy_magic_23_0.X.t41 GNDA 0.093585f
C1565 two_stage_opamp_dummy_magic_23_0.X.n62 GNDA 0.084458f
C1566 two_stage_opamp_dummy_magic_23_0.X.n63 GNDA 0.05169f
C1567 two_stage_opamp_dummy_magic_23_0.X.n64 GNDA 0.05169f
C1568 two_stage_opamp_dummy_magic_23_0.X.n65 GNDA 0.05169f
C1569 two_stage_opamp_dummy_magic_23_0.X.n66 GNDA 0.05169f
C1570 two_stage_opamp_dummy_magic_23_0.X.n67 GNDA 0.05169f
C1571 two_stage_opamp_dummy_magic_23_0.X.n68 GNDA 0.043554f
C1572 two_stage_opamp_dummy_magic_23_0.X.n69 GNDA 0.021431f
C1573 two_stage_opamp_dummy_magic_23_0.X.n70 GNDA 0.092553f
C1574 two_stage_opamp_dummy_magic_23_0.X.n71 GNDA 1.05185f
C1575 two_stage_opamp_dummy_magic_23_0.X.n72 GNDA 0.412424f
C1576 two_stage_opamp_dummy_magic_23_0.X.n73 GNDA 0.199954f
C1577 two_stage_opamp_dummy_magic_23_0.Vb1.t11 GNDA 0.025704f
C1578 two_stage_opamp_dummy_magic_23_0.Vb1.t10 GNDA 0.025704f
C1579 two_stage_opamp_dummy_magic_23_0.Vb1.n0 GNDA 0.091378f
C1580 two_stage_opamp_dummy_magic_23_0.Vb1.n1 GNDA 0.038556f
C1581 two_stage_opamp_dummy_magic_23_0.Vb1.t26 GNDA 0.602322f
C1582 two_stage_opamp_dummy_magic_23_0.Vb1.n2 GNDA 0.166741f
C1583 two_stage_opamp_dummy_magic_23_0.Vb1.t9 GNDA 0.019278f
C1584 two_stage_opamp_dummy_magic_23_0.Vb1.t1 GNDA 0.019278f
C1585 two_stage_opamp_dummy_magic_23_0.Vb1.n3 GNDA 0.041947f
C1586 two_stage_opamp_dummy_magic_23_0.Vb1.n4 GNDA 0.168509f
C1587 two_stage_opamp_dummy_magic_23_0.Vb1.t4 GNDA 0.01976f
C1588 two_stage_opamp_dummy_magic_23_0.Vb1.t0 GNDA 0.02563f
C1589 two_stage_opamp_dummy_magic_23_0.Vb1.n5 GNDA 0.026351f
C1590 two_stage_opamp_dummy_magic_23_0.Vb1.t2 GNDA 0.01976f
C1591 two_stage_opamp_dummy_magic_23_0.Vb1.t6 GNDA 0.02563f
C1592 two_stage_opamp_dummy_magic_23_0.Vb1.n6 GNDA 0.026351f
C1593 two_stage_opamp_dummy_magic_23_0.Vb1.n7 GNDA 0.019642f
C1594 two_stage_opamp_dummy_magic_23_0.Vb1.n8 GNDA 0.054079f
C1595 two_stage_opamp_dummy_magic_23_0.Vb1.t5 GNDA 0.019278f
C1596 two_stage_opamp_dummy_magic_23_0.Vb1.t3 GNDA 0.019278f
C1597 two_stage_opamp_dummy_magic_23_0.Vb1.n9 GNDA 0.041947f
C1598 two_stage_opamp_dummy_magic_23_0.Vb1.n10 GNDA 0.133477f
C1599 two_stage_opamp_dummy_magic_23_0.Vb1.n11 GNDA 0.104382f
C1600 two_stage_opamp_dummy_magic_23_0.Vb1.t7 GNDA 0.019278f
C1601 two_stage_opamp_dummy_magic_23_0.Vb1.t8 GNDA 0.019278f
C1602 two_stage_opamp_dummy_magic_23_0.Vb1.n12 GNDA 0.041947f
C1603 two_stage_opamp_dummy_magic_23_0.Vb1.n13 GNDA 0.168509f
C1604 two_stage_opamp_dummy_magic_23_0.Vb1.n14 GNDA 0.300052f
C1605 two_stage_opamp_dummy_magic_23_0.Vb1.t31 GNDA 0.01976f
C1606 two_stage_opamp_dummy_magic_23_0.Vb1.t21 GNDA 0.01976f
C1607 two_stage_opamp_dummy_magic_23_0.Vb1.t29 GNDA 0.01976f
C1608 two_stage_opamp_dummy_magic_23_0.Vb1.t20 GNDA 0.01976f
C1609 two_stage_opamp_dummy_magic_23_0.Vb1.t28 GNDA 0.01976f
C1610 two_stage_opamp_dummy_magic_23_0.Vb1.t18 GNDA 0.01976f
C1611 two_stage_opamp_dummy_magic_23_0.Vb1.t13 GNDA 0.01976f
C1612 two_stage_opamp_dummy_magic_23_0.Vb1.t19 GNDA 0.01976f
C1613 two_stage_opamp_dummy_magic_23_0.Vb1.t27 GNDA 0.01976f
C1614 two_stage_opamp_dummy_magic_23_0.Vb1.t15 GNDA 0.01976f
C1615 two_stage_opamp_dummy_magic_23_0.Vb1.t25 GNDA 0.01976f
C1616 two_stage_opamp_dummy_magic_23_0.Vb1.t14 GNDA 0.01976f
C1617 two_stage_opamp_dummy_magic_23_0.Vb1.t23 GNDA 0.01976f
C1618 two_stage_opamp_dummy_magic_23_0.Vb1.t32 GNDA 0.01976f
C1619 two_stage_opamp_dummy_magic_23_0.Vb1.t24 GNDA 0.01976f
C1620 two_stage_opamp_dummy_magic_23_0.Vb1.t12 GNDA 0.01976f
C1621 two_stage_opamp_dummy_magic_23_0.Vb1.t22 GNDA 0.01976f
C1622 two_stage_opamp_dummy_magic_23_0.Vb1.t30 GNDA 0.01976f
C1623 two_stage_opamp_dummy_magic_23_0.Vb1.t16 GNDA 0.02563f
C1624 two_stage_opamp_dummy_magic_23_0.Vb1.n15 GNDA 0.027867f
C1625 two_stage_opamp_dummy_magic_23_0.Vb1.n16 GNDA 0.018796f
C1626 two_stage_opamp_dummy_magic_23_0.Vb1.n17 GNDA 0.018796f
C1627 two_stage_opamp_dummy_magic_23_0.Vb1.n18 GNDA 0.018796f
C1628 two_stage_opamp_dummy_magic_23_0.Vb1.n19 GNDA 0.018796f
C1629 two_stage_opamp_dummy_magic_23_0.Vb1.n20 GNDA 0.018796f
C1630 two_stage_opamp_dummy_magic_23_0.Vb1.n21 GNDA 0.018796f
C1631 two_stage_opamp_dummy_magic_23_0.Vb1.n22 GNDA 0.018796f
C1632 two_stage_opamp_dummy_magic_23_0.Vb1.n23 GNDA 0.145711f
C1633 two_stage_opamp_dummy_magic_23_0.Vb1.t17 GNDA 0.01976f
C1634 two_stage_opamp_dummy_magic_23_0.Vb1.n24 GNDA 0.145711f
C1635 two_stage_opamp_dummy_magic_23_0.Vb1.n25 GNDA 0.018796f
C1636 two_stage_opamp_dummy_magic_23_0.Vb1.n26 GNDA 0.018796f
C1637 two_stage_opamp_dummy_magic_23_0.Vb1.n27 GNDA 0.018796f
C1638 two_stage_opamp_dummy_magic_23_0.Vb1.n28 GNDA 0.018796f
C1639 two_stage_opamp_dummy_magic_23_0.Vb1.n29 GNDA 0.018796f
C1640 two_stage_opamp_dummy_magic_23_0.Vb1.n30 GNDA 0.018796f
C1641 two_stage_opamp_dummy_magic_23_0.Vb1.n31 GNDA 0.018796f
C1642 two_stage_opamp_dummy_magic_23_0.Vb1.n32 GNDA 0.018796f
C1643 two_stage_opamp_dummy_magic_23_0.Vb1.n33 GNDA 0.033499f
C1644 two_stage_opamp_dummy_magic_23_0.Vb1.n34 GNDA 1.20347f
C1645 bgr_11_0.VB1_CUR_BIAS GNDA 1.07668f
C1646 two_stage_opamp_dummy_magic_23_0.cap_res_X.t70 GNDA 0.344881f
C1647 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 GNDA 0.346131f
C1648 two_stage_opamp_dummy_magic_23_0.cap_res_X.t101 GNDA 0.344881f
C1649 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 GNDA 0.347585f
C1650 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 GNDA 0.378048f
C1651 two_stage_opamp_dummy_magic_23_0.cap_res_X.t107 GNDA 0.344881f
C1652 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 GNDA 0.346131f
C1653 two_stage_opamp_dummy_magic_23_0.cap_res_X.t62 GNDA 0.344881f
C1654 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 GNDA 0.346131f
C1655 two_stage_opamp_dummy_magic_23_0.cap_res_X.t138 GNDA 0.344881f
C1656 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 GNDA 0.346131f
C1657 two_stage_opamp_dummy_magic_23_0.cap_res_X.t13 GNDA 0.344881f
C1658 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 GNDA 0.346131f
C1659 two_stage_opamp_dummy_magic_23_0.cap_res_X.t43 GNDA 0.344881f
C1660 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 GNDA 0.346131f
C1661 two_stage_opamp_dummy_magic_23_0.cap_res_X.t57 GNDA 0.344881f
C1662 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 GNDA 0.346131f
C1663 two_stage_opamp_dummy_magic_23_0.cap_res_X.t3 GNDA 0.344881f
C1664 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 GNDA 0.346131f
C1665 two_stage_opamp_dummy_magic_23_0.cap_res_X.t19 GNDA 0.344881f
C1666 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 GNDA 0.346131f
C1667 two_stage_opamp_dummy_magic_23_0.cap_res_X.t49 GNDA 0.344881f
C1668 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 GNDA 0.346131f
C1669 two_stage_opamp_dummy_magic_23_0.cap_res_X.t61 GNDA 0.344881f
C1670 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 GNDA 0.346131f
C1671 two_stage_opamp_dummy_magic_23_0.cap_res_X.t85 GNDA 0.344881f
C1672 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 GNDA 0.346131f
C1673 two_stage_opamp_dummy_magic_23_0.cap_res_X.t97 GNDA 0.344881f
C1674 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 GNDA 0.346131f
C1675 two_stage_opamp_dummy_magic_23_0.cap_res_X.t52 GNDA 0.344881f
C1676 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 GNDA 0.346131f
C1677 two_stage_opamp_dummy_magic_23_0.cap_res_X.t64 GNDA 0.344881f
C1678 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 GNDA 0.346131f
C1679 two_stage_opamp_dummy_magic_23_0.cap_res_X.t89 GNDA 0.344881f
C1680 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 GNDA 0.346131f
C1681 two_stage_opamp_dummy_magic_23_0.cap_res_X.t99 GNDA 0.344881f
C1682 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 GNDA 0.346131f
C1683 two_stage_opamp_dummy_magic_23_0.cap_res_X.t129 GNDA 0.344881f
C1684 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 GNDA 0.346131f
C1685 two_stage_opamp_dummy_magic_23_0.cap_res_X.t5 GNDA 0.344881f
C1686 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 GNDA 0.346131f
C1687 two_stage_opamp_dummy_magic_23_0.cap_res_X.t95 GNDA 0.344881f
C1688 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 GNDA 0.346131f
C1689 two_stage_opamp_dummy_magic_23_0.cap_res_X.t106 GNDA 0.344881f
C1690 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 GNDA 0.346131f
C1691 two_stage_opamp_dummy_magic_23_0.cap_res_X.t135 GNDA 0.344881f
C1692 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 GNDA 0.346131f
C1693 two_stage_opamp_dummy_magic_23_0.cap_res_X.t10 GNDA 0.344881f
C1694 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 GNDA 0.346131f
C1695 two_stage_opamp_dummy_magic_23_0.cap_res_X.t37 GNDA 0.344881f
C1696 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 GNDA 0.346131f
C1697 two_stage_opamp_dummy_magic_23_0.cap_res_X.t54 GNDA 0.344881f
C1698 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 GNDA 0.346131f
C1699 two_stage_opamp_dummy_magic_23_0.cap_res_X.t72 GNDA 0.344881f
C1700 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 GNDA 0.346131f
C1701 two_stage_opamp_dummy_magic_23_0.cap_res_X.t91 GNDA 0.344881f
C1702 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 GNDA 0.346131f
C1703 two_stage_opamp_dummy_magic_23_0.cap_res_X.t44 GNDA 0.344881f
C1704 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 GNDA 0.346131f
C1705 two_stage_opamp_dummy_magic_23_0.cap_res_X.t55 GNDA 0.344881f
C1706 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 GNDA 0.346131f
C1707 two_stage_opamp_dummy_magic_23_0.cap_res_X.t96 GNDA 0.344881f
C1708 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 GNDA 0.346131f
C1709 two_stage_opamp_dummy_magic_23_0.cap_res_X.t84 GNDA 0.344881f
C1710 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 GNDA 0.361791f
C1711 two_stage_opamp_dummy_magic_23_0.cap_res_X.t36 GNDA 0.344881f
C1712 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 GNDA 0.185242f
C1713 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 GNDA 0.198255f
C1714 two_stage_opamp_dummy_magic_23_0.cap_res_X.t105 GNDA 0.344881f
C1715 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 GNDA 0.185242f
C1716 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 GNDA 0.196656f
C1717 two_stage_opamp_dummy_magic_23_0.cap_res_X.t76 GNDA 0.344881f
C1718 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 GNDA 0.185242f
C1719 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 GNDA 0.196656f
C1720 two_stage_opamp_dummy_magic_23_0.cap_res_X.t23 GNDA 0.344881f
C1721 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 GNDA 0.185242f
C1722 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 GNDA 0.196656f
C1723 two_stage_opamp_dummy_magic_23_0.cap_res_X.t128 GNDA 0.344881f
C1724 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 GNDA 0.185242f
C1725 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 GNDA 0.196656f
C1726 two_stage_opamp_dummy_magic_23_0.cap_res_X.t94 GNDA 0.344881f
C1727 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 GNDA 0.185242f
C1728 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 GNDA 0.196656f
C1729 two_stage_opamp_dummy_magic_23_0.cap_res_X.t59 GNDA 0.344881f
C1730 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 GNDA 0.185242f
C1731 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 GNDA 0.196656f
C1732 two_stage_opamp_dummy_magic_23_0.cap_res_X.t6 GNDA 0.344881f
C1733 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 GNDA 0.185242f
C1734 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 GNDA 0.196656f
C1735 two_stage_opamp_dummy_magic_23_0.cap_res_X.t109 GNDA 0.344881f
C1736 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 GNDA 0.185242f
C1737 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 GNDA 0.196656f
C1738 two_stage_opamp_dummy_magic_23_0.cap_res_X.t133 GNDA 0.344881f
C1739 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 GNDA 0.346131f
C1740 two_stage_opamp_dummy_magic_23_0.cap_res_X.t80 GNDA 0.166734f
C1741 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 GNDA 0.215061f
C1742 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 GNDA 0.184096f
C1743 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 GNDA 0.23357f
C1744 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 GNDA 0.184096f
C1745 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 GNDA 0.250829f
C1746 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 GNDA 0.184096f
C1747 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 GNDA 0.250829f
C1748 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 GNDA 0.184096f
C1749 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 GNDA 0.250829f
C1750 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 GNDA 0.184096f
C1751 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 GNDA 0.250829f
C1752 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 GNDA 0.184096f
C1753 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 GNDA 0.250829f
C1754 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 GNDA 0.184096f
C1755 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 GNDA 0.250829f
C1756 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 GNDA 0.184096f
C1757 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 GNDA 0.250829f
C1758 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 GNDA 0.184096f
C1759 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 GNDA 0.250829f
C1760 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 GNDA 0.184096f
C1761 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 GNDA 0.250829f
C1762 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 GNDA 0.184096f
C1763 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 GNDA 0.250829f
C1764 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 GNDA 0.184096f
C1765 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 GNDA 0.250829f
C1766 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 GNDA 0.184096f
C1767 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 GNDA 0.250829f
C1768 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 GNDA 0.184096f
C1769 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 GNDA 0.250829f
C1770 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 GNDA 0.184096f
C1771 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 GNDA 0.250829f
C1772 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 GNDA 0.184096f
C1773 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 GNDA 0.23357f
C1774 two_stage_opamp_dummy_magic_23_0.cap_res_X.t20 GNDA 0.343735f
C1775 two_stage_opamp_dummy_magic_23_0.cap_res_X.t123 GNDA 0.166734f
C1776 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 GNDA 0.216311f
C1777 two_stage_opamp_dummy_magic_23_0.cap_res_X.t58 GNDA 0.343735f
C1778 two_stage_opamp_dummy_magic_23_0.cap_res_X.t22 GNDA 0.166734f
C1779 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 GNDA 0.216311f
C1780 two_stage_opamp_dummy_magic_23_0.cap_res_X.t41 GNDA 0.343735f
C1781 two_stage_opamp_dummy_magic_23_0.cap_res_X.t100 GNDA 0.344881f
C1782 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 GNDA 0.36339f
C1783 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 GNDA 0.36339f
C1784 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 GNDA 0.185242f
C1785 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 GNDA 0.216311f
C1786 two_stage_opamp_dummy_magic_23_0.cap_res_X.t21 GNDA 0.343735f
C1787 two_stage_opamp_dummy_magic_23_0.cap_res_X.t29 GNDA 0.344881f
C1788 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 GNDA 0.185242f
C1789 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 GNDA 0.197803f
C1790 two_stage_opamp_dummy_magic_23_0.cap_res_X.t50 GNDA 0.343735f
C1791 two_stage_opamp_dummy_magic_23_0.cap_res_X.t53 GNDA 0.344881f
C1792 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 GNDA 0.185242f
C1793 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 GNDA 0.216311f
C1794 two_stage_opamp_dummy_magic_23_0.cap_res_X.t27 GNDA 0.343735f
C1795 two_stage_opamp_dummy_magic_23_0.cap_res_X.t35 GNDA 0.344881f
C1796 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 GNDA 0.185242f
C1797 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 GNDA 0.216311f
C1798 two_stage_opamp_dummy_magic_23_0.cap_res_X.t127 GNDA 0.343735f
C1799 two_stage_opamp_dummy_magic_23_0.cap_res_X.t134 GNDA 0.344881f
C1800 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 GNDA 0.185242f
C1801 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 GNDA 0.216311f
C1802 two_stage_opamp_dummy_magic_23_0.cap_res_X.t11 GNDA 0.343735f
C1803 two_stage_opamp_dummy_magic_23_0.cap_res_X.t69 GNDA 0.344881f
C1804 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 GNDA 0.36339f
C1805 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 GNDA 0.36339f
C1806 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 GNDA 0.185242f
C1807 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 GNDA 0.216311f
C1808 two_stage_opamp_dummy_magic_23_0.cap_res_X.t108 GNDA 0.343735f
C1809 two_stage_opamp_dummy_magic_23_0.cap_res_X.t40 GNDA 0.344881f
C1810 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 GNDA 0.36339f
C1811 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 GNDA 0.36339f
C1812 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 GNDA 0.185242f
C1813 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 GNDA 0.216311f
C1814 two_stage_opamp_dummy_magic_23_0.cap_res_X.t75 GNDA 0.343735f
C1815 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 GNDA 0.216311f
C1816 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 GNDA 0.185242f
C1817 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 GNDA 0.36339f
C1818 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 GNDA 0.36339f
C1819 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 GNDA 0.736617f
C1820 two_stage_opamp_dummy_magic_23_0.cap_res_X.t0 GNDA 0.297532f
C1821 VOUT-.t2 GNDA 0.047629f
C1822 VOUT-.t15 GNDA 0.047629f
C1823 VOUT-.n0 GNDA 0.097592f
C1824 VOUT-.n1 GNDA 0.249374f
C1825 VOUT-.n2 GNDA 0.03433f
C1826 VOUT-.n3 GNDA 0.060565f
C1827 VOUT-.t13 GNDA 0.047629f
C1828 VOUT-.t17 GNDA 0.047629f
C1829 VOUT-.n4 GNDA 0.097592f
C1830 VOUT-.n5 GNDA 0.290507f
C1831 VOUT-.t7 GNDA 0.047629f
C1832 VOUT-.t8 GNDA 0.047629f
C1833 VOUT-.n6 GNDA 0.097592f
C1834 VOUT-.n7 GNDA 0.285429f
C1835 VOUT-.n8 GNDA 0.060565f
C1836 VOUT-.n9 GNDA 0.03433f
C1837 VOUT-.t1 GNDA 0.047629f
C1838 VOUT-.t18 GNDA 0.047629f
C1839 VOUT-.n10 GNDA 0.097592f
C1840 VOUT-.n11 GNDA 0.285429f
C1841 VOUT-.n12 GNDA 0.03433f
C1842 VOUT-.t3 GNDA 0.047629f
C1843 VOUT-.t16 GNDA 0.047629f
C1844 VOUT-.n13 GNDA 0.097592f
C1845 VOUT-.n14 GNDA 0.285429f
C1846 VOUT-.n15 GNDA 0.03433f
C1847 VOUT-.n16 GNDA 0.060565f
C1848 VOUT-.t10 GNDA 0.047629f
C1849 VOUT-.t14 GNDA 0.047629f
C1850 VOUT-.n17 GNDA 0.097592f
C1851 VOUT-.n18 GNDA 0.290507f
C1852 VOUT-.n19 GNDA 0.050049f
C1853 VOUT-.n20 GNDA 0.198401f
C1854 VOUT-.t24 GNDA 0.322935f
C1855 VOUT-.t129 GNDA 0.317527f
C1856 VOUT-.n21 GNDA 0.212891f
C1857 VOUT-.t77 GNDA 0.317527f
C1858 VOUT-.n22 GNDA 0.138918f
C1859 VOUT-.t61 GNDA 0.322935f
C1860 VOUT-.t106 GNDA 0.317527f
C1861 VOUT-.n23 GNDA 0.212891f
C1862 VOUT-.t67 GNDA 0.317527f
C1863 VOUT-.t48 GNDA 0.322258f
C1864 VOUT-.t151 GNDA 0.322258f
C1865 VOUT-.t98 GNDA 0.322258f
C1866 VOUT-.t63 GNDA 0.322258f
C1867 VOUT-.t29 GNDA 0.322258f
C1868 VOUT-.t134 GNDA 0.322258f
C1869 VOUT-.t81 GNDA 0.322258f
C1870 VOUT-.t52 GNDA 0.322258f
C1871 VOUT-.t121 GNDA 0.322258f
C1872 VOUT-.t73 GNDA 0.322258f
C1873 VOUT-.t47 GNDA 0.317527f
C1874 VOUT-.n24 GNDA 0.213569f
C1875 VOUT-.t86 GNDA 0.317527f
C1876 VOUT-.n25 GNDA 0.273105f
C1877 VOUT-.t150 GNDA 0.317527f
C1878 VOUT-.n26 GNDA 0.273105f
C1879 VOUT-.t97 GNDA 0.317527f
C1880 VOUT-.n27 GNDA 0.273105f
C1881 VOUT-.t142 GNDA 0.317527f
C1882 VOUT-.n28 GNDA 0.273105f
C1883 VOUT-.t91 GNDA 0.317527f
C1884 VOUT-.n29 GNDA 0.273105f
C1885 VOUT-.t42 GNDA 0.317527f
C1886 VOUT-.n30 GNDA 0.273105f
C1887 VOUT-.t126 GNDA 0.317527f
C1888 VOUT-.n31 GNDA 0.273105f
C1889 VOUT-.t31 GNDA 0.317527f
C1890 VOUT-.n32 GNDA 0.273105f
C1891 VOUT-.t115 GNDA 0.317527f
C1892 VOUT-.n33 GNDA 0.273105f
C1893 VOUT-.n34 GNDA 0.257991f
C1894 VOUT-.t113 GNDA 0.322935f
C1895 VOUT-.t83 GNDA 0.317527f
C1896 VOUT-.n35 GNDA 0.212891f
C1897 VOUT-.t36 GNDA 0.317527f
C1898 VOUT-.t102 GNDA 0.322935f
C1899 VOUT-.t139 GNDA 0.317527f
C1900 VOUT-.n36 GNDA 0.212891f
C1901 VOUT-.n37 GNDA 0.257991f
C1902 VOUT-.t85 GNDA 0.322935f
C1903 VOUT-.t55 GNDA 0.317527f
C1904 VOUT-.n38 GNDA 0.212891f
C1905 VOUT-.t141 GNDA 0.317527f
C1906 VOUT-.t66 GNDA 0.322935f
C1907 VOUT-.t101 GNDA 0.317527f
C1908 VOUT-.n39 GNDA 0.212891f
C1909 VOUT-.n40 GNDA 0.257991f
C1910 VOUT-.t120 GNDA 0.322935f
C1911 VOUT-.t90 GNDA 0.317527f
C1912 VOUT-.n41 GNDA 0.212891f
C1913 VOUT-.t41 GNDA 0.317527f
C1914 VOUT-.t103 GNDA 0.322935f
C1915 VOUT-.t145 GNDA 0.317527f
C1916 VOUT-.n42 GNDA 0.212891f
C1917 VOUT-.n43 GNDA 0.257991f
C1918 VOUT-.t22 GNDA 0.322935f
C1919 VOUT-.t127 GNDA 0.317527f
C1920 VOUT-.n44 GNDA 0.212891f
C1921 VOUT-.t74 GNDA 0.317527f
C1922 VOUT-.t147 GNDA 0.322935f
C1923 VOUT-.t46 GNDA 0.317527f
C1924 VOUT-.n45 GNDA 0.212891f
C1925 VOUT-.n46 GNDA 0.257991f
C1926 VOUT-.t56 GNDA 0.322935f
C1927 VOUT-.t153 GNDA 0.317527f
C1928 VOUT-.n47 GNDA 0.212891f
C1929 VOUT-.t39 GNDA 0.317527f
C1930 VOUT-.n48 GNDA 0.138918f
C1931 VOUT-.t87 GNDA 0.322935f
C1932 VOUT-.t54 GNDA 0.317527f
C1933 VOUT-.n49 GNDA 0.212891f
C1934 VOUT-.t69 GNDA 0.317527f
C1935 VOUT-.t137 GNDA 0.322258f
C1936 VOUT-.t99 GNDA 0.322258f
C1937 VOUT-.t57 GNDA 0.322935f
C1938 VOUT-.t92 GNDA 0.317527f
C1939 VOUT-.n50 GNDA 0.212891f
C1940 VOUT-.t109 GNDA 0.317527f
C1941 VOUT-.n51 GNDA 0.133957f
C1942 VOUT-.t116 GNDA 0.322258f
C1943 VOUT-.t156 GNDA 0.322935f
C1944 VOUT-.t59 GNDA 0.317527f
C1945 VOUT-.n52 GNDA 0.212891f
C1946 VOUT-.t75 GNDA 0.317527f
C1947 VOUT-.n53 GNDA 0.133957f
C1948 VOUT-.t82 GNDA 0.322258f
C1949 VOUT-.t117 GNDA 0.322935f
C1950 VOUT-.t20 GNDA 0.317527f
C1951 VOUT-.n54 GNDA 0.212891f
C1952 VOUT-.t44 GNDA 0.317527f
C1953 VOUT-.n55 GNDA 0.133957f
C1954 VOUT-.t49 GNDA 0.322258f
C1955 VOUT-.t88 GNDA 0.322935f
C1956 VOUT-.t123 GNDA 0.317527f
C1957 VOUT-.n56 GNDA 0.212891f
C1958 VOUT-.t143 GNDA 0.317527f
C1959 VOUT-.n57 GNDA 0.133957f
C1960 VOUT-.t146 GNDA 0.322258f
C1961 VOUT-.t23 GNDA 0.322524f
C1962 VOUT-.t30 GNDA 0.322258f
C1963 VOUT-.t122 GNDA 0.322524f
C1964 VOUT-.t130 GNDA 0.322258f
C1965 VOUT-.t104 GNDA 0.322524f
C1966 VOUT-.t107 GNDA 0.322258f
C1967 VOUT-.t128 GNDA 0.322524f
C1968 VOUT-.t136 GNDA 0.322258f
C1969 VOUT-.t33 GNDA 0.317527f
C1970 VOUT-.n58 GNDA 0.351459f
C1971 VOUT-.t149 GNDA 0.317527f
C1972 VOUT-.n59 GNDA 0.410995f
C1973 VOUT-.t25 GNDA 0.317527f
C1974 VOUT-.n60 GNDA 0.410995f
C1975 VOUT-.t64 GNDA 0.317527f
C1976 VOUT-.n61 GNDA 0.410995f
C1977 VOUT-.t45 GNDA 0.317527f
C1978 VOUT-.n62 GNDA 0.337603f
C1979 VOUT-.t78 GNDA 0.317527f
C1980 VOUT-.n63 GNDA 0.337603f
C1981 VOUT-.t111 GNDA 0.317527f
C1982 VOUT-.n64 GNDA 0.337603f
C1983 VOUT-.t155 GNDA 0.317527f
C1984 VOUT-.n65 GNDA 0.337603f
C1985 VOUT-.t135 GNDA 0.317527f
C1986 VOUT-.n66 GNDA 0.273105f
C1987 VOUT-.t34 GNDA 0.317527f
C1988 VOUT-.n67 GNDA 0.273105f
C1989 VOUT-.n68 GNDA 0.257991f
C1990 VOUT-.t50 GNDA 0.322935f
C1991 VOUT-.t148 GNDA 0.317527f
C1992 VOUT-.n69 GNDA 0.212891f
C1993 VOUT-.t32 GNDA 0.317527f
C1994 VOUT-.t95 GNDA 0.322935f
C1995 VOUT-.t131 GNDA 0.317527f
C1996 VOUT-.n70 GNDA 0.212891f
C1997 VOUT-.n71 GNDA 0.257991f
C1998 VOUT-.t19 GNDA 0.322935f
C1999 VOUT-.t119 GNDA 0.317527f
C2000 VOUT-.n72 GNDA 0.212891f
C2001 VOUT-.t70 GNDA 0.317527f
C2002 VOUT-.t144 GNDA 0.322935f
C2003 VOUT-.t40 GNDA 0.317527f
C2004 VOUT-.n73 GNDA 0.212891f
C2005 VOUT-.n74 GNDA 0.257991f
C2006 VOUT-.t114 GNDA 0.322935f
C2007 VOUT-.t84 GNDA 0.317527f
C2008 VOUT-.n75 GNDA 0.212891f
C2009 VOUT-.t37 GNDA 0.317527f
C2010 VOUT-.t100 GNDA 0.322935f
C2011 VOUT-.t140 GNDA 0.317527f
C2012 VOUT-.n76 GNDA 0.212891f
C2013 VOUT-.n77 GNDA 0.257991f
C2014 VOUT-.t154 GNDA 0.322935f
C2015 VOUT-.t112 GNDA 0.317527f
C2016 VOUT-.n78 GNDA 0.212891f
C2017 VOUT-.t65 GNDA 0.317527f
C2018 VOUT-.t138 GNDA 0.322935f
C2019 VOUT-.t35 GNDA 0.317527f
C2020 VOUT-.n79 GNDA 0.212891f
C2021 VOUT-.n80 GNDA 0.257991f
C2022 VOUT-.t108 GNDA 0.322935f
C2023 VOUT-.t76 GNDA 0.317527f
C2024 VOUT-.n81 GNDA 0.212891f
C2025 VOUT-.t26 GNDA 0.317527f
C2026 VOUT-.t96 GNDA 0.322935f
C2027 VOUT-.t132 GNDA 0.317527f
C2028 VOUT-.n82 GNDA 0.212891f
C2029 VOUT-.n83 GNDA 0.257991f
C2030 VOUT-.t72 GNDA 0.322935f
C2031 VOUT-.t43 GNDA 0.317527f
C2032 VOUT-.n84 GNDA 0.212891f
C2033 VOUT-.t125 GNDA 0.317527f
C2034 VOUT-.t60 GNDA 0.322935f
C2035 VOUT-.t94 GNDA 0.317527f
C2036 VOUT-.n85 GNDA 0.212891f
C2037 VOUT-.n86 GNDA 0.257991f
C2038 VOUT-.t105 GNDA 0.322935f
C2039 VOUT-.t71 GNDA 0.317527f
C2040 VOUT-.n87 GNDA 0.212891f
C2041 VOUT-.t21 GNDA 0.317527f
C2042 VOUT-.t93 GNDA 0.322935f
C2043 VOUT-.t124 GNDA 0.317527f
C2044 VOUT-.n88 GNDA 0.212891f
C2045 VOUT-.n89 GNDA 0.257991f
C2046 VOUT-.t68 GNDA 0.322935f
C2047 VOUT-.t38 GNDA 0.317527f
C2048 VOUT-.n90 GNDA 0.212891f
C2049 VOUT-.t118 GNDA 0.317527f
C2050 VOUT-.t58 GNDA 0.322935f
C2051 VOUT-.t89 GNDA 0.317527f
C2052 VOUT-.n91 GNDA 0.212891f
C2053 VOUT-.n92 GNDA 0.257991f
C2054 VOUT-.t28 GNDA 0.322935f
C2055 VOUT-.t133 GNDA 0.317527f
C2056 VOUT-.n93 GNDA 0.212891f
C2057 VOUT-.t80 GNDA 0.317527f
C2058 VOUT-.t152 GNDA 0.322935f
C2059 VOUT-.t53 GNDA 0.317527f
C2060 VOUT-.n94 GNDA 0.212891f
C2061 VOUT-.n95 GNDA 0.257991f
C2062 VOUT-.t62 GNDA 0.322935f
C2063 VOUT-.t27 GNDA 0.317527f
C2064 VOUT-.n96 GNDA 0.212891f
C2065 VOUT-.t110 GNDA 0.317527f
C2066 VOUT-.n97 GNDA 0.257991f
C2067 VOUT-.t79 GNDA 0.317527f
C2068 VOUT-.n98 GNDA 0.138918f
C2069 VOUT-.t51 GNDA 0.317527f
C2070 VOUT-.n99 GNDA 0.252511f
C2071 VOUT-.n100 GNDA 0.309727f
C2072 VOUT-.n101 GNDA 0.084056f
C2073 VOUT-.t9 GNDA 0.055567f
C2074 VOUT-.t11 GNDA 0.055567f
C2075 VOUT-.n102 GNDA 0.119393f
C2076 VOUT-.n103 GNDA 0.333803f
C2077 VOUT-.t6 GNDA 0.055567f
C2078 VOUT-.t4 GNDA 0.055567f
C2079 VOUT-.n104 GNDA 0.119393f
C2080 VOUT-.n105 GNDA 0.321626f
C2081 VOUT-.n106 GNDA 0.11654f
C2082 VOUT-.t12 GNDA 0.055567f
C2083 VOUT-.t0 GNDA 0.055567f
C2084 VOUT-.n107 GNDA 0.119393f
C2085 VOUT-.n108 GNDA 0.326528f
C2086 VOUT-.n109 GNDA 0.056324f
C2087 VOUT-.t5 GNDA 0.091827f
C2088 VOUT-.n110 GNDA 0.111609f
C2089 bgr_11_0.cap_res2.t8 GNDA 0.399727f
C2090 bgr_11_0.cap_res2.t13 GNDA 0.401176f
C2091 bgr_11_0.cap_res2.t3 GNDA 0.379724f
C2092 bgr_11_0.cap_res2.t2 GNDA 0.399727f
C2093 bgr_11_0.cap_res2.t7 GNDA 0.401176f
C2094 bgr_11_0.cap_res2.t17 GNDA 0.379724f
C2095 bgr_11_0.cap_res2.t15 GNDA 0.399727f
C2096 bgr_11_0.cap_res2.t1 GNDA 0.401176f
C2097 bgr_11_0.cap_res2.t11 GNDA 0.379724f
C2098 bgr_11_0.cap_res2.t0 GNDA 0.399727f
C2099 bgr_11_0.cap_res2.t5 GNDA 0.401176f
C2100 bgr_11_0.cap_res2.t16 GNDA 0.379724f
C2101 bgr_11_0.cap_res2.t14 GNDA 0.399727f
C2102 bgr_11_0.cap_res2.t19 GNDA 0.401176f
C2103 bgr_11_0.cap_res2.t9 GNDA 0.379724f
C2104 bgr_11_0.cap_res2.n0 GNDA 0.267938f
C2105 bgr_11_0.cap_res2.t4 GNDA 0.213373f
C2106 bgr_11_0.cap_res2.n1 GNDA 0.290719f
C2107 bgr_11_0.cap_res2.t10 GNDA 0.213373f
C2108 bgr_11_0.cap_res2.n2 GNDA 0.290719f
C2109 bgr_11_0.cap_res2.t6 GNDA 0.213373f
C2110 bgr_11_0.cap_res2.n3 GNDA 0.290719f
C2111 bgr_11_0.cap_res2.t12 GNDA 0.213373f
C2112 bgr_11_0.cap_res2.n4 GNDA 0.290719f
C2113 bgr_11_0.cap_res2.t18 GNDA 0.416168f
C2114 bgr_11_0.cap_res2.t20 GNDA 0.096398f
C2115 bgr_11_0.NFET_GATE_10uA.n0 GNDA 1.79799f
C2116 bgr_11_0.NFET_GATE_10uA.t21 GNDA 0.01337f
C2117 bgr_11_0.NFET_GATE_10uA.n1 GNDA 0.014733f
C2118 bgr_11_0.NFET_GATE_10uA.t19 GNDA 0.01337f
C2119 bgr_11_0.NFET_GATE_10uA.n2 GNDA 0.016546f
C2120 bgr_11_0.NFET_GATE_10uA.n3 GNDA 0.011828f
C2121 bgr_11_0.NFET_GATE_10uA.n4 GNDA 0.010014f
C2122 bgr_11_0.NFET_GATE_10uA.n5 GNDA 0.01584f
C2123 bgr_11_0.NFET_GATE_10uA.t20 GNDA 0.01337f
C2124 bgr_11_0.NFET_GATE_10uA.n6 GNDA 0.014733f
C2125 bgr_11_0.NFET_GATE_10uA.t5 GNDA 0.01337f
C2126 bgr_11_0.NFET_GATE_10uA.n7 GNDA 0.014733f
C2127 bgr_11_0.NFET_GATE_10uA.n8 GNDA 0.014432f
C2128 bgr_11_0.NFET_GATE_10uA.n9 GNDA 0.395351f
C2129 bgr_11_0.NFET_GATE_10uA.t11 GNDA 0.01337f
C2130 bgr_11_0.NFET_GATE_10uA.n10 GNDA 0.016546f
C2131 bgr_11_0.NFET_GATE_10uA.n11 GNDA 0.011828f
C2132 bgr_11_0.NFET_GATE_10uA.n12 GNDA 0.010014f
C2133 bgr_11_0.NFET_GATE_10uA.t13 GNDA 0.01337f
C2134 bgr_11_0.NFET_GATE_10uA.n13 GNDA 0.014733f
C2135 bgr_11_0.NFET_GATE_10uA.n14 GNDA 0.014432f
C2136 bgr_11_0.NFET_GATE_10uA.n15 GNDA 0.2494f
C2137 bgr_11_0.NFET_GATE_10uA.t0 GNDA 0.01337f
C2138 bgr_11_0.NFET_GATE_10uA.n16 GNDA 0.014733f
C2139 bgr_11_0.NFET_GATE_10uA.t7 GNDA 0.010677f
C2140 bgr_11_0.NFET_GATE_10uA.n17 GNDA 0.02003f
C2141 bgr_11_0.NFET_GATE_10uA.n18 GNDA 0.030903f
C2142 bgr_11_0.NFET_GATE_10uA.n19 GNDA 0.070319f
C2143 VOUT+.n0 GNDA 0.08395f
C2144 VOUT+.t6 GNDA 0.055563f
C2145 VOUT+.t3 GNDA 0.055563f
C2146 VOUT+.n1 GNDA 0.119383f
C2147 VOUT+.n2 GNDA 0.333776f
C2148 VOUT+.t2 GNDA 0.055563f
C2149 VOUT+.t1 GNDA 0.055563f
C2150 VOUT+.n3 GNDA 0.119383f
C2151 VOUT+.n4 GNDA 0.321601f
C2152 VOUT+.n5 GNDA 0.116531f
C2153 VOUT+.t4 GNDA 0.055563f
C2154 VOUT+.t5 GNDA 0.055563f
C2155 VOUT+.n6 GNDA 0.119383f
C2156 VOUT+.n7 GNDA 0.327689f
C2157 VOUT+.n8 GNDA 0.060497f
C2158 VOUT+.t0 GNDA 0.091865f
C2159 VOUT+.n9 GNDA 0.11622f
C2160 VOUT+.t9 GNDA 0.047625f
C2161 VOUT+.t14 GNDA 0.047625f
C2162 VOUT+.n10 GNDA 0.097584f
C2163 VOUT+.n11 GNDA 0.249355f
C2164 VOUT+.t17 GNDA 0.047625f
C2165 VOUT+.t15 GNDA 0.047625f
C2166 VOUT+.n12 GNDA 0.097584f
C2167 VOUT+.n13 GNDA 0.290484f
C2168 VOUT+.n14 GNDA 0.034328f
C2169 VOUT+.n15 GNDA 0.06056f
C2170 VOUT+.t8 GNDA 0.047625f
C2171 VOUT+.t18 GNDA 0.047625f
C2172 VOUT+.n16 GNDA 0.097584f
C2173 VOUT+.n17 GNDA 0.290484f
C2174 VOUT+.n18 GNDA 0.06056f
C2175 VOUT+.t10 GNDA 0.047625f
C2176 VOUT+.t13 GNDA 0.047625f
C2177 VOUT+.n19 GNDA 0.097584f
C2178 VOUT+.n20 GNDA 0.285406f
C2179 VOUT+.n21 GNDA 0.06056f
C2180 VOUT+.t11 GNDA 0.047625f
C2181 VOUT+.t16 GNDA 0.047625f
C2182 VOUT+.n22 GNDA 0.097584f
C2183 VOUT+.n23 GNDA 0.285406f
C2184 VOUT+.n24 GNDA 0.034328f
C2185 VOUT+.n25 GNDA 0.034328f
C2186 VOUT+.t12 GNDA 0.047625f
C2187 VOUT+.t7 GNDA 0.047625f
C2188 VOUT+.n26 GNDA 0.097584f
C2189 VOUT+.n27 GNDA 0.285406f
C2190 VOUT+.n28 GNDA 0.034328f
C2191 VOUT+.n29 GNDA 0.050045f
C2192 VOUT+.n30 GNDA 0.198804f
C2193 VOUT+.t63 GNDA 0.317501f
C2194 VOUT+.t35 GNDA 0.322909f
C2195 VOUT+.t34 GNDA 0.317501f
C2196 VOUT+.n31 GNDA 0.212874f
C2197 VOUT+.n32 GNDA 0.138907f
C2198 VOUT+.t99 GNDA 0.322232f
C2199 VOUT+.t149 GNDA 0.322232f
C2200 VOUT+.t43 GNDA 0.322232f
C2201 VOUT+.t77 GNDA 0.322232f
C2202 VOUT+.t125 GNDA 0.322232f
C2203 VOUT+.t20 GNDA 0.322232f
C2204 VOUT+.t59 GNDA 0.322232f
C2205 VOUT+.t92 GNDA 0.322232f
C2206 VOUT+.t143 GNDA 0.322232f
C2207 VOUT+.t39 GNDA 0.322232f
C2208 VOUT+.t95 GNDA 0.317501f
C2209 VOUT+.n33 GNDA 0.213552f
C2210 VOUT+.t146 GNDA 0.317501f
C2211 VOUT+.n34 GNDA 0.273083f
C2212 VOUT+.t107 GNDA 0.317501f
C2213 VOUT+.n35 GNDA 0.273083f
C2214 VOUT+.t153 GNDA 0.317501f
C2215 VOUT+.n36 GNDA 0.273083f
C2216 VOUT+.t65 GNDA 0.317501f
C2217 VOUT+.n37 GNDA 0.273083f
C2218 VOUT+.t113 GNDA 0.317501f
C2219 VOUT+.n38 GNDA 0.273083f
C2220 VOUT+.t72 GNDA 0.317501f
C2221 VOUT+.n39 GNDA 0.273083f
C2222 VOUT+.t120 GNDA 0.317501f
C2223 VOUT+.n40 GNDA 0.273083f
C2224 VOUT+.t31 GNDA 0.317501f
C2225 VOUT+.n41 GNDA 0.273083f
C2226 VOUT+.t132 GNDA 0.317501f
C2227 VOUT+.n42 GNDA 0.273083f
C2228 VOUT+.t45 GNDA 0.317501f
C2229 VOUT+.t58 GNDA 0.322909f
C2230 VOUT+.t147 GNDA 0.317501f
C2231 VOUT+.n43 GNDA 0.212874f
C2232 VOUT+.n44 GNDA 0.25797f
C2233 VOUT+.t103 GNDA 0.322909f
C2234 VOUT+.t49 GNDA 0.317501f
C2235 VOUT+.n45 GNDA 0.212874f
C2236 VOUT+.t152 GNDA 0.317501f
C2237 VOUT+.t130 GNDA 0.322909f
C2238 VOUT+.t127 GNDA 0.317501f
C2239 VOUT+.n46 GNDA 0.212874f
C2240 VOUT+.n47 GNDA 0.25797f
C2241 VOUT+.t67 GNDA 0.322909f
C2242 VOUT+.t155 GNDA 0.317501f
C2243 VOUT+.n48 GNDA 0.212874f
C2244 VOUT+.t116 GNDA 0.317501f
C2245 VOUT+.t98 GNDA 0.322909f
C2246 VOUT+.t96 GNDA 0.317501f
C2247 VOUT+.n49 GNDA 0.212874f
C2248 VOUT+.n50 GNDA 0.25797f
C2249 VOUT+.t109 GNDA 0.322909f
C2250 VOUT+.t55 GNDA 0.317501f
C2251 VOUT+.n51 GNDA 0.212874f
C2252 VOUT+.t19 GNDA 0.317501f
C2253 VOUT+.t136 GNDA 0.322909f
C2254 VOUT+.t134 GNDA 0.317501f
C2255 VOUT+.n52 GNDA 0.212874f
C2256 VOUT+.n53 GNDA 0.25797f
C2257 VOUT+.t145 GNDA 0.322909f
C2258 VOUT+.t93 GNDA 0.317501f
C2259 VOUT+.n54 GNDA 0.212874f
C2260 VOUT+.t60 GNDA 0.317501f
C2261 VOUT+.t32 GNDA 0.322909f
C2262 VOUT+.t30 GNDA 0.317501f
C2263 VOUT+.n55 GNDA 0.212874f
C2264 VOUT+.n56 GNDA 0.25797f
C2265 VOUT+.t36 GNDA 0.317501f
C2266 VOUT+.t66 GNDA 0.322909f
C2267 VOUT+.t28 GNDA 0.317501f
C2268 VOUT+.n57 GNDA 0.212874f
C2269 VOUT+.n58 GNDA 0.138907f
C2270 VOUT+.t75 GNDA 0.322232f
C2271 VOUT+.t53 GNDA 0.322232f
C2272 VOUT+.t137 GNDA 0.322909f
C2273 VOUT+.t33 GNDA 0.317501f
C2274 VOUT+.n59 GNDA 0.212874f
C2275 VOUT+.t86 GNDA 0.317501f
C2276 VOUT+.n60 GNDA 0.133946f
C2277 VOUT+.t90 GNDA 0.322232f
C2278 VOUT+.t27 GNDA 0.322909f
C2279 VOUT+.t69 GNDA 0.317501f
C2280 VOUT+.n61 GNDA 0.212874f
C2281 VOUT+.t122 GNDA 0.317501f
C2282 VOUT+.n62 GNDA 0.133946f
C2283 VOUT+.t126 GNDA 0.322232f
C2284 VOUT+.t81 GNDA 0.322909f
C2285 VOUT+.t119 GNDA 0.317501f
C2286 VOUT+.n63 GNDA 0.212874f
C2287 VOUT+.t106 GNDA 0.317501f
C2288 VOUT+.n64 GNDA 0.133946f
C2289 VOUT+.t110 GNDA 0.322232f
C2290 VOUT+.t114 GNDA 0.322909f
C2291 VOUT+.t156 GNDA 0.317501f
C2292 VOUT+.n65 GNDA 0.212874f
C2293 VOUT+.t140 GNDA 0.317501f
C2294 VOUT+.n66 GNDA 0.133946f
C2295 VOUT+.t148 GNDA 0.322232f
C2296 VOUT+.t37 GNDA 0.322498f
C2297 VOUT+.t44 GNDA 0.322232f
C2298 VOUT+.t76 GNDA 0.322498f
C2299 VOUT+.t82 GNDA 0.322232f
C2300 VOUT+.t56 GNDA 0.322498f
C2301 VOUT+.t61 GNDA 0.322232f
C2302 VOUT+.t91 GNDA 0.322498f
C2303 VOUT+.t100 GNDA 0.322232f
C2304 VOUT+.t131 GNDA 0.317501f
C2305 VOUT+.n67 GNDA 0.351431f
C2306 VOUT+.t94 GNDA 0.317501f
C2307 VOUT+.n68 GNDA 0.410962f
C2308 VOUT+.t115 GNDA 0.317501f
C2309 VOUT+.n69 GNDA 0.410962f
C2310 VOUT+.t78 GNDA 0.317501f
C2311 VOUT+.n70 GNDA 0.410962f
C2312 VOUT+.t42 GNDA 0.317501f
C2313 VOUT+.n71 GNDA 0.337576f
C2314 VOUT+.t141 GNDA 0.317501f
C2315 VOUT+.n72 GNDA 0.337576f
C2316 VOUT+.t22 GNDA 0.317501f
C2317 VOUT+.n73 GNDA 0.337576f
C2318 VOUT+.t124 GNDA 0.317501f
C2319 VOUT+.n74 GNDA 0.337576f
C2320 VOUT+.t87 GNDA 0.317501f
C2321 VOUT+.n75 GNDA 0.273083f
C2322 VOUT+.t112 GNDA 0.317501f
C2323 VOUT+.n76 GNDA 0.273083f
C2324 VOUT+.t71 GNDA 0.317501f
C2325 VOUT+.t105 GNDA 0.322909f
C2326 VOUT+.t68 GNDA 0.317501f
C2327 VOUT+.n77 GNDA 0.212874f
C2328 VOUT+.n78 GNDA 0.25797f
C2329 VOUT+.t48 GNDA 0.322909f
C2330 VOUT+.t70 GNDA 0.317501f
C2331 VOUT+.n79 GNDA 0.212874f
C2332 VOUT+.t29 GNDA 0.317501f
C2333 VOUT+.t62 GNDA 0.322909f
C2334 VOUT+.t24 GNDA 0.317501f
C2335 VOUT+.n80 GNDA 0.212874f
C2336 VOUT+.n81 GNDA 0.25797f
C2337 VOUT+.t139 GNDA 0.322909f
C2338 VOUT+.t88 GNDA 0.317501f
C2339 VOUT+.n82 GNDA 0.212874f
C2340 VOUT+.t54 GNDA 0.317501f
C2341 VOUT+.t26 GNDA 0.322909f
C2342 VOUT+.t25 GNDA 0.317501f
C2343 VOUT+.n83 GNDA 0.212874f
C2344 VOUT+.n84 GNDA 0.25797f
C2345 VOUT+.t104 GNDA 0.322909f
C2346 VOUT+.t51 GNDA 0.317501f
C2347 VOUT+.n85 GNDA 0.212874f
C2348 VOUT+.t154 GNDA 0.317501f
C2349 VOUT+.t129 GNDA 0.322909f
C2350 VOUT+.t128 GNDA 0.317501f
C2351 VOUT+.n86 GNDA 0.212874f
C2352 VOUT+.n87 GNDA 0.25797f
C2353 VOUT+.t135 GNDA 0.322909f
C2354 VOUT+.t83 GNDA 0.317501f
C2355 VOUT+.n88 GNDA 0.212874f
C2356 VOUT+.t50 GNDA 0.317501f
C2357 VOUT+.t23 GNDA 0.322909f
C2358 VOUT+.t21 GNDA 0.317501f
C2359 VOUT+.n89 GNDA 0.212874f
C2360 VOUT+.n90 GNDA 0.25797f
C2361 VOUT+.t97 GNDA 0.322909f
C2362 VOUT+.t46 GNDA 0.317501f
C2363 VOUT+.n91 GNDA 0.212874f
C2364 VOUT+.t150 GNDA 0.317501f
C2365 VOUT+.t123 GNDA 0.322909f
C2366 VOUT+.t121 GNDA 0.317501f
C2367 VOUT+.n92 GNDA 0.212874f
C2368 VOUT+.n93 GNDA 0.25797f
C2369 VOUT+.t57 GNDA 0.322909f
C2370 VOUT+.t144 GNDA 0.317501f
C2371 VOUT+.n94 GNDA 0.212874f
C2372 VOUT+.t111 GNDA 0.317501f
C2373 VOUT+.t85 GNDA 0.322909f
C2374 VOUT+.t84 GNDA 0.317501f
C2375 VOUT+.n95 GNDA 0.212874f
C2376 VOUT+.n96 GNDA 0.25797f
C2377 VOUT+.t89 GNDA 0.322909f
C2378 VOUT+.t38 GNDA 0.317501f
C2379 VOUT+.n97 GNDA 0.212874f
C2380 VOUT+.t142 GNDA 0.317501f
C2381 VOUT+.t118 GNDA 0.322909f
C2382 VOUT+.t117 GNDA 0.317501f
C2383 VOUT+.n98 GNDA 0.212874f
C2384 VOUT+.n99 GNDA 0.25797f
C2385 VOUT+.t52 GNDA 0.322909f
C2386 VOUT+.t138 GNDA 0.317501f
C2387 VOUT+.n100 GNDA 0.212874f
C2388 VOUT+.t108 GNDA 0.317501f
C2389 VOUT+.t80 GNDA 0.322909f
C2390 VOUT+.t79 GNDA 0.317501f
C2391 VOUT+.n101 GNDA 0.212874f
C2392 VOUT+.n102 GNDA 0.25797f
C2393 VOUT+.t151 GNDA 0.322909f
C2394 VOUT+.t102 GNDA 0.317501f
C2395 VOUT+.n103 GNDA 0.212874f
C2396 VOUT+.t64 GNDA 0.317501f
C2397 VOUT+.t41 GNDA 0.322909f
C2398 VOUT+.t40 GNDA 0.317501f
C2399 VOUT+.n104 GNDA 0.212874f
C2400 VOUT+.n105 GNDA 0.25797f
C2401 VOUT+.t74 GNDA 0.322909f
C2402 VOUT+.t73 GNDA 0.317501f
C2403 VOUT+.n106 GNDA 0.212874f
C2404 VOUT+.t101 GNDA 0.317501f
C2405 VOUT+.n107 GNDA 0.25797f
C2406 VOUT+.t133 GNDA 0.317501f
C2407 VOUT+.n108 GNDA 0.138907f
C2408 VOUT+.t47 GNDA 0.317501f
C2409 VOUT+.n109 GNDA 0.252491f
C2410 VOUT+.n110 GNDA 0.308286f
C2411 VDDA.t548 GNDA 0.040257f
C2412 VDDA.t637 GNDA 0.040257f
C2413 VDDA.t696 GNDA 0.040257f
C2414 VDDA.t492 GNDA 0.040257f
C2415 VDDA.t480 GNDA 0.040257f
C2416 VDDA.t573 GNDA 0.040257f
C2417 VDDA.t663 GNDA 0.040257f
C2418 VDDA.t717 GNDA 0.040257f
C2419 VDDA.t515 GNDA 0.040257f
C2420 VDDA.t503 GNDA 0.040257f
C2421 VDDA.t594 GNDA 0.040257f
C2422 VDDA.t682 GNDA 0.040257f
C2423 VDDA.t475 GNDA 0.040257f
C2424 VDDA.t591 GNDA 0.040257f
C2425 VDDA.t581 GNDA 0.052626f
C2426 VDDA.n0 GNDA 0.029422f
C2427 VDDA.n1 GNDA 0.02147f
C2428 VDDA.n2 GNDA 0.02147f
C2429 VDDA.n3 GNDA 0.02147f
C2430 VDDA.n4 GNDA 0.02147f
C2431 VDDA.n5 GNDA 0.020022f
C2432 VDDA.t27 GNDA 0.053053f
C2433 VDDA.n6 GNDA 0.015528f
C2434 VDDA.n7 GNDA 0.015528f
C2435 VDDA.n8 GNDA 0.015528f
C2436 VDDA.t436 GNDA 0.155972f
C2437 VDDA.t488 GNDA 0.15336f
C2438 VDDA.n9 GNDA 0.102823f
C2439 VDDA.t526 GNDA 0.15336f
C2440 VDDA.n10 GNDA 0.067095f
C2441 VDDA.t443 GNDA 0.15336f
C2442 VDDA.n11 GNDA 0.067095f
C2443 VDDA.t664 GNDA 0.15336f
C2444 VDDA.n12 GNDA 0.067095f
C2445 VDDA.t708 GNDA 0.15336f
C2446 VDDA.t430 GNDA 0.155972f
C2447 VDDA.t516 GNDA 0.15336f
C2448 VDDA.n13 GNDA 0.102823f
C2449 VDDA.t598 GNDA 0.15336f
C2450 VDDA.n14 GNDA 0.067095f
C2451 VDDA.t545 GNDA 0.15336f
C2452 VDDA.n15 GNDA 0.067095f
C2453 VDDA.t626 GNDA 0.15336f
C2454 VDDA.n16 GNDA 0.067095f
C2455 VDDA.n17 GNDA 0.09585f
C2456 VDDA.t651 GNDA 0.155972f
C2457 VDDA.t700 GNDA 0.15336f
C2458 VDDA.n18 GNDA 0.102823f
C2459 VDDA.t438 GNDA 0.15336f
C2460 VDDA.n19 GNDA 0.067095f
C2461 VDDA.t658 GNDA 0.15336f
C2462 VDDA.n20 GNDA 0.067095f
C2463 VDDA.t577 GNDA 0.15336f
C2464 VDDA.n21 GNDA 0.067095f
C2465 VDDA.t620 GNDA 0.15336f
C2466 VDDA.t642 GNDA 0.155972f
C2467 VDDA.t425 GNDA 0.15336f
C2468 VDDA.n22 GNDA 0.102823f
C2469 VDDA.t510 GNDA 0.15336f
C2470 VDDA.n23 GNDA 0.067095f
C2471 VDDA.t459 GNDA 0.15336f
C2472 VDDA.n24 GNDA 0.067095f
C2473 VDDA.t540 GNDA 0.15336f
C2474 VDDA.n25 GNDA 0.067095f
C2475 VDDA.n26 GNDA 0.124605f
C2476 VDDA.t424 GNDA 0.155972f
C2477 VDDA.t476 GNDA 0.15336f
C2478 VDDA.n27 GNDA 0.102823f
C2479 VDDA.t517 GNDA 0.15336f
C2480 VDDA.n28 GNDA 0.067095f
C2481 VDDA.t432 GNDA 0.15336f
C2482 VDDA.n29 GNDA 0.067095f
C2483 VDDA.t650 GNDA 0.15336f
C2484 VDDA.n30 GNDA 0.067095f
C2485 VDDA.t697 GNDA 0.15336f
C2486 VDDA.t720 GNDA 0.155972f
C2487 VDDA.t505 GNDA 0.15336f
C2488 VDDA.n31 GNDA 0.102823f
C2489 VDDA.t585 GNDA 0.15336f
C2490 VDDA.n32 GNDA 0.067095f
C2491 VDDA.t535 GNDA 0.15336f
C2492 VDDA.n33 GNDA 0.067095f
C2493 VDDA.t616 GNDA 0.15336f
C2494 VDDA.n34 GNDA 0.067095f
C2495 VDDA.n35 GNDA 0.124605f
C2496 VDDA.t638 GNDA 0.155972f
C2497 VDDA.t690 GNDA 0.15336f
C2498 VDDA.n36 GNDA 0.102823f
C2499 VDDA.t428 GNDA 0.15336f
C2500 VDDA.n37 GNDA 0.067095f
C2501 VDDA.t646 GNDA 0.15336f
C2502 VDDA.n38 GNDA 0.067095f
C2503 VDDA.t568 GNDA 0.15336f
C2504 VDDA.n39 GNDA 0.067095f
C2505 VDDA.t612 GNDA 0.15336f
C2506 VDDA.t632 GNDA 0.155972f
C2507 VDDA.t714 GNDA 0.15336f
C2508 VDDA.n40 GNDA 0.102823f
C2509 VDDA.t499 GNDA 0.15336f
C2510 VDDA.n41 GNDA 0.067095f
C2511 VDDA.t450 GNDA 0.15336f
C2512 VDDA.n42 GNDA 0.067095f
C2513 VDDA.t531 GNDA 0.15336f
C2514 VDDA.n43 GNDA 0.067095f
C2515 VDDA.n44 GNDA 0.124605f
C2516 VDDA.t556 GNDA 0.155972f
C2517 VDDA.t605 GNDA 0.15336f
C2518 VDDA.n45 GNDA 0.102823f
C2519 VDDA.t641 GNDA 0.15336f
C2520 VDDA.n46 GNDA 0.067095f
C2521 VDDA.t562 GNDA 0.15336f
C2522 VDDA.n47 GNDA 0.067095f
C2523 VDDA.t483 GNDA 0.15336f
C2524 VDDA.n48 GNDA 0.067095f
C2525 VDDA.t528 GNDA 0.15336f
C2526 VDDA.t549 GNDA 0.155972f
C2527 VDDA.t627 GNDA 0.15336f
C2528 VDDA.n49 GNDA 0.102823f
C2529 VDDA.t711 GNDA 0.15336f
C2530 VDDA.n50 GNDA 0.067095f
C2531 VDDA.t668 GNDA 0.15336f
C2532 VDDA.n51 GNDA 0.067095f
C2533 VDDA.t445 GNDA 0.15336f
C2534 VDDA.n52 GNDA 0.067095f
C2535 VDDA.n53 GNDA 0.124605f
C2536 VDDA.t471 GNDA 0.155972f
C2537 VDDA.t520 GNDA 0.15336f
C2538 VDDA.n54 GNDA 0.102823f
C2539 VDDA.t557 GNDA 0.15336f
C2540 VDDA.n55 GNDA 0.067095f
C2541 VDDA.t477 GNDA 0.15336f
C2542 VDDA.n56 GNDA 0.067095f
C2543 VDDA.t694 GNDA 0.15336f
C2544 VDDA.n57 GNDA 0.067095f
C2545 VDDA.t441 GNDA 0.15336f
C2546 VDDA.t463 GNDA 0.155972f
C2547 VDDA.t543 GNDA 0.15336f
C2548 VDDA.n58 GNDA 0.102823f
C2549 VDDA.t624 GNDA 0.15336f
C2550 VDDA.n59 GNDA 0.067095f
C2551 VDDA.t583 GNDA 0.15336f
C2552 VDDA.n60 GNDA 0.067095f
C2553 VDDA.t661 GNDA 0.15336f
C2554 VDDA.n61 GNDA 0.067095f
C2555 VDDA.n62 GNDA 0.124605f
C2556 VDDA.t542 GNDA 0.155972f
C2557 VDDA.t597 GNDA 0.15336f
C2558 VDDA.n63 GNDA 0.102823f
C2559 VDDA.t629 GNDA 0.15336f
C2560 VDDA.n64 GNDA 0.067095f
C2561 VDDA.t551 GNDA 0.15336f
C2562 VDDA.n65 GNDA 0.067095f
C2563 VDDA.t470 GNDA 0.15336f
C2564 VDDA.n66 GNDA 0.067095f
C2565 VDDA.t521 GNDA 0.15336f
C2566 VDDA.t536 GNDA 0.155972f
C2567 VDDA.t618 GNDA 0.15336f
C2568 VDDA.n67 GNDA 0.102823f
C2569 VDDA.t702 GNDA 0.15336f
C2570 VDDA.n68 GNDA 0.067095f
C2571 VDDA.t654 GNDA 0.15336f
C2572 VDDA.n69 GNDA 0.067095f
C2573 VDDA.t435 GNDA 0.15336f
C2574 VDDA.n70 GNDA 0.067095f
C2575 VDDA.n71 GNDA 0.124605f
C2576 VDDA.t458 GNDA 0.155972f
C2577 VDDA.t509 GNDA 0.15336f
C2578 VDDA.n72 GNDA 0.102823f
C2579 VDDA.t546 GNDA 0.15336f
C2580 VDDA.n73 GNDA 0.067095f
C2581 VDDA.t466 GNDA 0.15336f
C2582 VDDA.n74 GNDA 0.067095f
C2583 VDDA.t685 GNDA 0.15336f
C2584 VDDA.n75 GNDA 0.067095f
C2585 VDDA.t431 GNDA 0.15336f
C2586 VDDA.t451 GNDA 0.155972f
C2587 VDDA.t532 GNDA 0.15336f
C2588 VDDA.n76 GNDA 0.102823f
C2589 VDDA.t615 GNDA 0.15336f
C2590 VDDA.n77 GNDA 0.067095f
C2591 VDDA.t570 GNDA 0.15336f
C2592 VDDA.n78 GNDA 0.067095f
C2593 VDDA.t649 GNDA 0.15336f
C2594 VDDA.n79 GNDA 0.067095f
C2595 VDDA.n80 GNDA 0.124605f
C2596 VDDA.t675 GNDA 0.155972f
C2597 VDDA.t721 GNDA 0.15336f
C2598 VDDA.n81 GNDA 0.102823f
C2599 VDDA.t460 GNDA 0.15336f
C2600 VDDA.n82 GNDA 0.067095f
C2601 VDDA.t680 GNDA 0.15336f
C2602 VDDA.n83 GNDA 0.067095f
C2603 VDDA.t602 GNDA 0.15336f
C2604 VDDA.n84 GNDA 0.067095f
C2605 VDDA.t643 GNDA 0.15336f
C2606 VDDA.t669 GNDA 0.155972f
C2607 VDDA.t448 GNDA 0.15336f
C2608 VDDA.n85 GNDA 0.102823f
C2609 VDDA.t530 GNDA 0.15336f
C2610 VDDA.n86 GNDA 0.067095f
C2611 VDDA.t485 GNDA 0.15336f
C2612 VDDA.n87 GNDA 0.067095f
C2613 VDDA.t566 GNDA 0.15336f
C2614 VDDA.n88 GNDA 0.067095f
C2615 VDDA.n89 GNDA 0.124605f
C2616 VDDA.t447 GNDA 0.155972f
C2617 VDDA.t498 GNDA 0.15336f
C2618 VDDA.n90 GNDA 0.102823f
C2619 VDDA.t533 GNDA 0.15336f
C2620 VDDA.n91 GNDA 0.067095f
C2621 VDDA.t452 GNDA 0.15336f
C2622 VDDA.n92 GNDA 0.067095f
C2623 VDDA.t674 GNDA 0.15336f
C2624 VDDA.n93 GNDA 0.067095f
C2625 VDDA.t718 GNDA 0.15336f
C2626 VDDA.t442 GNDA 0.155972f
C2627 VDDA.t525 GNDA 0.15336f
C2628 VDDA.n94 GNDA 0.102823f
C2629 VDDA.t607 GNDA 0.15336f
C2630 VDDA.n95 GNDA 0.067095f
C2631 VDDA.t559 GNDA 0.15336f
C2632 VDDA.n96 GNDA 0.067095f
C2633 VDDA.t636 GNDA 0.15336f
C2634 VDDA.n97 GNDA 0.067095f
C2635 VDDA.n98 GNDA 0.124605f
C2636 VDDA.t665 GNDA 0.155972f
C2637 VDDA.t710 GNDA 0.15336f
C2638 VDDA.n99 GNDA 0.102823f
C2639 VDDA.t449 GNDA 0.15336f
C2640 VDDA.n100 GNDA 0.067095f
C2641 VDDA.t670 GNDA 0.15336f
C2642 VDDA.n101 GNDA 0.067095f
C2643 VDDA.t590 GNDA 0.15336f
C2644 VDDA.n102 GNDA 0.067095f
C2645 VDDA.t631 GNDA 0.15336f
C2646 VDDA.t656 GNDA 0.155972f
C2647 VDDA.t437 GNDA 0.15336f
C2648 VDDA.n103 GNDA 0.102823f
C2649 VDDA.t523 GNDA 0.15336f
C2650 VDDA.n104 GNDA 0.067095f
C2651 VDDA.t473 GNDA 0.15336f
C2652 VDDA.n105 GNDA 0.067095f
C2653 VDDA.t554 GNDA 0.15336f
C2654 VDDA.n106 GNDA 0.067095f
C2655 VDDA.n107 GNDA 0.124605f
C2656 VDDA.t580 GNDA 0.155972f
C2657 VDDA.t623 GNDA 0.15336f
C2658 VDDA.n108 GNDA 0.102823f
C2659 VDDA.t666 GNDA 0.15336f
C2660 VDDA.n109 GNDA 0.067095f
C2661 VDDA.t586 GNDA 0.15336f
C2662 VDDA.n110 GNDA 0.067095f
C2663 VDDA.t506 GNDA 0.15336f
C2664 VDDA.n111 GNDA 0.067095f
C2665 VDDA.t547 GNDA 0.15336f
C2666 VDDA.t574 GNDA 0.155972f
C2667 VDDA.t653 GNDA 0.15336f
C2668 VDDA.n112 GNDA 0.102823f
C2669 VDDA.t434 GNDA 0.15336f
C2670 VDDA.n113 GNDA 0.067095f
C2671 VDDA.t688 GNDA 0.15336f
C2672 VDDA.n114 GNDA 0.067095f
C2673 VDDA.t468 GNDA 0.15336f
C2674 VDDA.n115 GNDA 0.067095f
C2675 VDDA.n116 GNDA 0.124605f
C2676 VDDA.t652 GNDA 0.155972f
C2677 VDDA.t701 GNDA 0.15336f
C2678 VDDA.n117 GNDA 0.102823f
C2679 VDDA.t439 GNDA 0.15336f
C2680 VDDA.n118 GNDA 0.067095f
C2681 VDDA.t659 GNDA 0.15336f
C2682 VDDA.n119 GNDA 0.067095f
C2683 VDDA.t578 GNDA 0.15336f
C2684 VDDA.n120 GNDA 0.067095f
C2685 VDDA.t621 GNDA 0.15336f
C2686 VDDA.t644 GNDA 0.155972f
C2687 VDDA.t426 GNDA 0.15336f
C2688 VDDA.n121 GNDA 0.102823f
C2689 VDDA.t511 GNDA 0.15336f
C2690 VDDA.n122 GNDA 0.067095f
C2691 VDDA.t461 GNDA 0.15336f
C2692 VDDA.n123 GNDA 0.067095f
C2693 VDDA.t541 GNDA 0.15336f
C2694 VDDA.n124 GNDA 0.067095f
C2695 VDDA.n125 GNDA 0.124605f
C2696 VDDA.t569 GNDA 0.155972f
C2697 VDDA.t614 GNDA 0.15336f
C2698 VDDA.n126 GNDA 0.102823f
C2699 VDDA.t655 GNDA 0.15336f
C2700 VDDA.n127 GNDA 0.067095f
C2701 VDDA.t576 GNDA 0.15336f
C2702 VDDA.n128 GNDA 0.067095f
C2703 VDDA.t493 GNDA 0.15336f
C2704 VDDA.n129 GNDA 0.067095f
C2705 VDDA.t537 GNDA 0.15336f
C2706 VDDA.t560 GNDA 0.155972f
C2707 VDDA.t639 GNDA 0.15336f
C2708 VDDA.n130 GNDA 0.102823f
C2709 VDDA.t722 GNDA 0.15336f
C2710 VDDA.n131 GNDA 0.067095f
C2711 VDDA.t676 GNDA 0.15336f
C2712 VDDA.n132 GNDA 0.067095f
C2713 VDDA.t456 GNDA 0.15336f
C2714 VDDA.n133 GNDA 0.067095f
C2715 VDDA.n134 GNDA 0.124605f
C2716 VDDA.t495 GNDA 0.155972f
C2717 VDDA.t538 GNDA 0.15336f
C2718 VDDA.n135 GNDA 0.102823f
C2719 VDDA.t584 GNDA 0.15336f
C2720 VDDA.n136 GNDA 0.067095f
C2721 VDDA.t502 GNDA 0.15336f
C2722 VDDA.n137 GNDA 0.067095f
C2723 VDDA.t716 GNDA 0.15336f
C2724 VDDA.n138 GNDA 0.067095f
C2725 VDDA.t465 GNDA 0.15336f
C2726 VDDA.t490 GNDA 0.155972f
C2727 VDDA.t571 GNDA 0.15336f
C2728 VDDA.n139 GNDA 0.102823f
C2729 VDDA.t648 GNDA 0.15336f
C2730 VDDA.n140 GNDA 0.067095f
C2731 VDDA.t606 GNDA 0.15336f
C2732 VDDA.n141 GNDA 0.067095f
C2733 VDDA.t683 GNDA 0.15336f
C2734 VDDA.n142 GNDA 0.067095f
C2735 VDDA.n143 GNDA 0.124605f
C2736 VDDA.t707 GNDA 0.155972f
C2737 VDDA.t454 GNDA 0.15336f
C2738 VDDA.n144 GNDA 0.102823f
C2739 VDDA.t496 GNDA 0.15336f
C2740 VDDA.n145 GNDA 0.067095f
C2741 VDDA.t713 GNDA 0.15336f
C2742 VDDA.n146 GNDA 0.067095f
C2743 VDDA.t630 GNDA 0.15336f
C2744 VDDA.n147 GNDA 0.067095f
C2745 VDDA.t679 GNDA 0.15336f
C2746 VDDA.t703 GNDA 0.155972f
C2747 VDDA.t486 GNDA 0.15336f
C2748 VDDA.n148 GNDA 0.102823f
C2749 VDDA.t565 GNDA 0.15336f
C2750 VDDA.n149 GNDA 0.067095f
C2751 VDDA.t522 GNDA 0.15336f
C2752 VDDA.n150 GNDA 0.067095f
C2753 VDDA.t601 GNDA 0.15336f
C2754 VDDA.n151 GNDA 0.067095f
C2755 VDDA.n152 GNDA 0.124605f
C2756 VDDA.t484 GNDA 0.155972f
C2757 VDDA.t529 GNDA 0.15336f
C2758 VDDA.n153 GNDA 0.102823f
C2759 VDDA.t572 GNDA 0.15336f
C2760 VDDA.n154 GNDA 0.067095f
C2761 VDDA.t491 GNDA 0.15336f
C2762 VDDA.n155 GNDA 0.067095f
C2763 VDDA.t706 GNDA 0.15336f
C2764 VDDA.n156 GNDA 0.067095f
C2765 VDDA.t453 GNDA 0.15336f
C2766 VDDA.t479 GNDA 0.155972f
C2767 VDDA.t558 GNDA 0.15336f
C2768 VDDA.n157 GNDA 0.102823f
C2769 VDDA.t635 GNDA 0.15336f
C2770 VDDA.n158 GNDA 0.067095f
C2771 VDDA.t596 GNDA 0.15336f
C2772 VDDA.n159 GNDA 0.067095f
C2773 VDDA.t673 GNDA 0.15336f
C2774 VDDA.n160 GNDA 0.067095f
C2775 VDDA.n161 GNDA 0.124605f
C2776 VDDA.t695 GNDA 0.155972f
C2777 VDDA.t444 GNDA 0.15336f
C2778 VDDA.n162 GNDA 0.102823f
C2779 VDDA.t487 GNDA 0.15336f
C2780 VDDA.n163 GNDA 0.067095f
C2781 VDDA.t704 GNDA 0.15336f
C2782 VDDA.n164 GNDA 0.067095f
C2783 VDDA.t619 GNDA 0.15336f
C2784 VDDA.n165 GNDA 0.067095f
C2785 VDDA.t671 GNDA 0.15336f
C2786 VDDA.t691 GNDA 0.155972f
C2787 VDDA.t472 GNDA 0.15336f
C2788 VDDA.n166 GNDA 0.102823f
C2789 VDDA.t553 GNDA 0.15336f
C2790 VDDA.n167 GNDA 0.067095f
C2791 VDDA.t508 GNDA 0.15336f
C2792 VDDA.n168 GNDA 0.067095f
C2793 VDDA.t589 GNDA 0.15336f
C2794 VDDA.n169 GNDA 0.067095f
C2795 VDDA.n170 GNDA 0.124605f
C2796 VDDA.t611 GNDA 0.155972f
C2797 VDDA.t660 GNDA 0.15336f
C2798 VDDA.n171 GNDA 0.102823f
C2799 VDDA.t699 GNDA 0.15336f
C2800 VDDA.n172 GNDA 0.067095f
C2801 VDDA.t617 GNDA 0.15336f
C2802 VDDA.n173 GNDA 0.067095f
C2803 VDDA.t534 GNDA 0.15336f
C2804 VDDA.n174 GNDA 0.067095f
C2805 VDDA.t587 GNDA 0.15336f
C2806 VDDA.t608 GNDA 0.155972f
C2807 VDDA.t687 GNDA 0.15336f
C2808 VDDA.n175 GNDA 0.102823f
C2809 VDDA.t467 GNDA 0.15336f
C2810 VDDA.n176 GNDA 0.067095f
C2811 VDDA.t719 GNDA 0.15336f
C2812 VDDA.n177 GNDA 0.067095f
C2813 VDDA.t504 GNDA 0.15336f
C2814 VDDA.n178 GNDA 0.067095f
C2815 VDDA.n179 GNDA 0.124605f
C2816 VDDA.t686 GNDA 0.155972f
C2817 VDDA.t433 GNDA 0.15336f
C2818 VDDA.n180 GNDA 0.102823f
C2819 VDDA.t474 GNDA 0.15336f
C2820 VDDA.n181 GNDA 0.067095f
C2821 VDDA.t692 GNDA 0.15336f
C2822 VDDA.n182 GNDA 0.067095f
C2823 VDDA.t610 GNDA 0.15336f
C2824 VDDA.n183 GNDA 0.067095f
C2825 VDDA.t657 GNDA 0.15336f
C2826 VDDA.t681 GNDA 0.155972f
C2827 VDDA.t462 GNDA 0.15336f
C2828 VDDA.n184 GNDA 0.102823f
C2829 VDDA.t539 GNDA 0.15336f
C2830 VDDA.n185 GNDA 0.067095f
C2831 VDDA.t497 GNDA 0.15336f
C2832 VDDA.n186 GNDA 0.067095f
C2833 VDDA.t579 GNDA 0.15336f
C2834 VDDA.n187 GNDA 0.067095f
C2835 VDDA.n188 GNDA 0.124605f
C2836 VDDA.t603 GNDA 0.155972f
C2837 VDDA.t647 GNDA 0.15336f
C2838 VDDA.n189 GNDA 0.102823f
C2839 VDDA.t689 GNDA 0.15336f
C2840 VDDA.n190 GNDA 0.067095f
C2841 VDDA.t609 GNDA 0.15336f
C2842 VDDA.n191 GNDA 0.067095f
C2843 VDDA.t527 GNDA 0.15336f
C2844 VDDA.n192 GNDA 0.067095f
C2845 VDDA.t575 GNDA 0.15336f
C2846 VDDA.t599 GNDA 0.155972f
C2847 VDDA.t677 GNDA 0.15336f
C2848 VDDA.n193 GNDA 0.102823f
C2849 VDDA.t455 GNDA 0.15336f
C2850 VDDA.n194 GNDA 0.067095f
C2851 VDDA.t709 GNDA 0.15336f
C2852 VDDA.n195 GNDA 0.067095f
C2853 VDDA.t494 GNDA 0.15336f
C2854 VDDA.n196 GNDA 0.067095f
C2855 VDDA.n197 GNDA 0.124605f
C2856 VDDA.t519 GNDA 0.155972f
C2857 VDDA.t564 GNDA 0.15336f
C2858 VDDA.n198 GNDA 0.102823f
C2859 VDDA.t604 GNDA 0.15336f
C2860 VDDA.n199 GNDA 0.067095f
C2861 VDDA.t524 GNDA 0.15336f
C2862 VDDA.n200 GNDA 0.067095f
C2863 VDDA.t440 GNDA 0.15336f
C2864 VDDA.n201 GNDA 0.067095f
C2865 VDDA.t489 GNDA 0.15336f
C2866 VDDA.t512 GNDA 0.155972f
C2867 VDDA.t593 GNDA 0.15336f
C2868 VDDA.n202 GNDA 0.102823f
C2869 VDDA.t672 GNDA 0.15336f
C2870 VDDA.n203 GNDA 0.067095f
C2871 VDDA.t622 GNDA 0.15336f
C2872 VDDA.n204 GNDA 0.067095f
C2873 VDDA.t705 GNDA 0.15336f
C2874 VDDA.n205 GNDA 0.067095f
C2875 VDDA.n206 GNDA 0.124605f
C2876 VDDA.t592 GNDA 0.155972f
C2877 VDDA.t634 GNDA 0.15336f
C2878 VDDA.n207 GNDA 0.102823f
C2879 VDDA.t678 GNDA 0.15336f
C2880 VDDA.n208 GNDA 0.067095f
C2881 VDDA.t600 GNDA 0.15336f
C2882 VDDA.n209 GNDA 0.067095f
C2883 VDDA.t518 GNDA 0.15336f
C2884 VDDA.n210 GNDA 0.067095f
C2885 VDDA.t563 GNDA 0.15336f
C2886 VDDA.t588 GNDA 0.155972f
C2887 VDDA.t667 GNDA 0.15336f
C2888 VDDA.n211 GNDA 0.102823f
C2889 VDDA.t446 GNDA 0.15336f
C2890 VDDA.n212 GNDA 0.067095f
C2891 VDDA.t698 GNDA 0.15336f
C2892 VDDA.n213 GNDA 0.067095f
C2893 VDDA.t482 GNDA 0.15336f
C2894 VDDA.n214 GNDA 0.067095f
C2895 VDDA.n215 GNDA 0.124605f
C2896 VDDA.t507 GNDA 0.155972f
C2897 VDDA.t552 GNDA 0.15336f
C2898 VDDA.n216 GNDA 0.102823f
C2899 VDDA.t595 GNDA 0.15336f
C2900 VDDA.n217 GNDA 0.067095f
C2901 VDDA.t514 GNDA 0.15336f
C2902 VDDA.n218 GNDA 0.067095f
C2903 VDDA.t429 GNDA 0.15336f
C2904 VDDA.n219 GNDA 0.067095f
C2905 VDDA.t478 GNDA 0.15336f
C2906 VDDA.n220 GNDA 0.09585f
C2907 VDDA.t693 GNDA 0.15336f
C2908 VDDA.n221 GNDA 0.067095f
C2909 VDDA.t613 GNDA 0.15336f
C2910 VDDA.n222 GNDA 0.067095f
C2911 VDDA.t662 GNDA 0.15336f
C2912 VDDA.n223 GNDA 0.067095f
C2913 VDDA.t582 GNDA 0.15336f
C2914 VDDA.n224 GNDA 0.067095f
C2915 VDDA.t500 GNDA 0.15336f
C2916 VDDA.n225 GNDA 0.066267f
C2917 VDDA.n226 GNDA 0.014377f
C2918 VDDA.n229 GNDA 0.015528f
C2919 VDDA.n230 GNDA 0.015528f
C2920 VDDA.n231 GNDA 0.016103f
C2921 VDDA.n232 GNDA 0.014377f
C2922 VDDA.n233 GNDA 0.032195f
C2923 VDDA.t26 GNDA 0.041968f
C2924 VDDA.n234 GNDA 0.359389f
C2925 VDDA.n235 GNDA 0.312927f
C2926 VDDA.n236 GNDA 0.015528f
C2927 VDDA.n237 GNDA 0.015528f
C2928 VDDA.n238 GNDA 0.015528f
C2929 VDDA.n239 GNDA 0.016103f
C2930 VDDA.n240 GNDA 0.016103f
C2931 VDDA.n241 GNDA 0.016103f
C2932 VDDA.n242 GNDA 0.016103f
C2933 VDDA.n243 GNDA 0.043793f
C2934 VDDA.n244 GNDA 0.016302f
C2935 VDDA.n245 GNDA 0.014668f
C2936 VDDA.n246 GNDA 0.299879f
C2937 VDDA.n249 GNDA 0.011981f
C2938 VDDA.n252 GNDA 0.014377f
C2939 VDDA.n255 GNDA 0.014377f
C2940 VDDA.n258 GNDA 0.291383f
C2941 VDDA.n259 GNDA 2.23138f
C2942 VDDA.n260 GNDA 0.145692f
C2943 VDDA.n262 GNDA 0.291383f
C2944 VDDA.n264 GNDA 0.15336f
C2945 VDDA.n265 GNDA 0.149526f
C2946 VDDA.n267 GNDA 0.145692f
C2947 VDDA.n269 GNDA 0.164862f
C2948 VDDA.n273 GNDA 0.15336f
C2949 VDDA.n275 GNDA 0.149526f
C2950 VDDA.n276 GNDA 0.322055f
C2951 VDDA.n277 GNDA 3.22055f
C2952 VDDA.n278 GNDA 0.015528f
C2953 VDDA.n279 GNDA 0.015528f
C2954 VDDA.n280 GNDA 0.016103f
C2955 VDDA.n281 GNDA 0.014377f
C2956 VDDA.t189 GNDA 0.21432f
C2957 VDDA.t379 GNDA 0.215097f
C2958 VDDA.t281 GNDA 0.203595f
C2959 VDDA.t349 GNDA 0.21432f
C2960 VDDA.t302 GNDA 0.215097f
C2961 VDDA.t216 GNDA 0.203595f
C2962 VDDA.t296 GNDA 0.21432f
C2963 VDDA.t258 GNDA 0.215097f
C2964 VDDA.t375 GNDA 0.203595f
C2965 VDDA.t304 GNDA 0.21432f
C2966 VDDA.t318 GNDA 0.215097f
C2967 VDDA.t214 GNDA 0.203595f
C2968 VDDA.t283 GNDA 0.21432f
C2969 VDDA.t240 GNDA 0.215097f
C2970 VDDA.t365 GNDA 0.203595f
C2971 VDDA.n282 GNDA 0.143659f
C2972 VDDA.t298 GNDA 0.114403f
C2973 VDDA.n283 GNDA 0.155873f
C2974 VDDA.t343 GNDA 0.114403f
C2975 VDDA.n284 GNDA 0.155873f
C2976 VDDA.t300 GNDA 0.114403f
C2977 VDDA.n285 GNDA 0.155873f
C2978 VDDA.t377 GNDA 0.114403f
C2979 VDDA.n286 GNDA 0.155873f
C2980 VDDA.t218 GNDA 0.198749f
C2981 VDDA.t625 GNDA 0.15336f
C2982 VDDA.t513 GNDA 0.155972f
C2983 VDDA.t427 GNDA 0.15336f
C2984 VDDA.n287 GNDA 0.102823f
C2985 VDDA.t645 GNDA 0.15336f
C2986 VDDA.t567 GNDA 0.155972f
C2987 VDDA.n288 GNDA 0.131578f
C2988 VDDA.t723 GNDA 0.155972f
C2989 VDDA.t640 GNDA 0.15336f
C2990 VDDA.n289 GNDA 0.102823f
C2991 VDDA.t561 GNDA 0.15336f
C2992 VDDA.t481 GNDA 0.155972f
C2993 VDDA.n290 GNDA 0.160333f
C2994 VDDA.t501 GNDA 0.155972f
C2995 VDDA.t715 GNDA 0.15336f
C2996 VDDA.n291 GNDA 0.102823f
C2997 VDDA.t633 GNDA 0.15336f
C2998 VDDA.t555 GNDA 0.155972f
C2999 VDDA.n292 GNDA 0.160333f
C3000 VDDA.t712 GNDA 0.155972f
C3001 VDDA.t628 GNDA 0.15336f
C3002 VDDA.n293 GNDA 0.102823f
C3003 VDDA.t550 GNDA 0.15336f
C3004 VDDA.t469 GNDA 0.155972f
C3005 VDDA.n294 GNDA 0.160333f
C3006 VDDA.t684 GNDA 0.155972f
C3007 VDDA.t464 GNDA 0.15336f
C3008 VDDA.n295 GNDA 0.131578f
C3009 VDDA.t544 GNDA 0.15336f
C3010 VDDA.n296 GNDA 0.067095f
C3011 VDDA.n297 GNDA 0.143836f
C3012 VDDA.n298 GNDA 0.63978f
C3013 VDDA.n300 GNDA 0.073533f
C3014 VDDA.n301 GNDA 0.012993f
C3015 VDDA.n302 GNDA 0.035903f
C3016 VDDA.t79 GNDA 0.0521f
C3017 VDDA.n304 GNDA 0.055956f
C3018 VDDA.n305 GNDA 0.01687f
C3019 VDDA.n306 GNDA 0.012993f
C3020 VDDA.n307 GNDA 0.035903f
C3021 VDDA.n309 GNDA 0.045545f
C3022 VDDA.t359 GNDA 0.010019f
C3023 VDDA.n310 GNDA 0.081531f
C3024 VDDA.n311 GNDA 0.65987f
C3025 VDDA.n312 GNDA 0.158195f
C3026 VDDA.n313 GNDA 0.015528f
C3027 VDDA.n314 GNDA 0.015528f
C3028 VDDA.n315 GNDA 0.015528f
C3029 VDDA.n316 GNDA 0.016103f
C3030 VDDA.n317 GNDA 0.016103f
C3031 VDDA.n318 GNDA 0.016103f
C3032 VDDA.n319 GNDA 0.016103f
C3033 VDDA.n320 GNDA 0.043793f
C3034 VDDA.n321 GNDA 0.016302f
C3035 VDDA.n322 GNDA 0.014668f
C3036 VDDA.n323 GNDA 3.80332f
C3037 VDDA.n324 GNDA 0.015528f
C3038 VDDA.n325 GNDA 0.015528f
C3039 VDDA.n326 GNDA 0.016103f
C3040 VDDA.n327 GNDA 0.014377f
C3041 VDDA.n328 GNDA 0.021759f
C3042 VDDA.t289 GNDA 0.011028f
C3043 VDDA.n329 GNDA 0.016101f
C3044 VDDA.t291 GNDA 0.020216f
C3045 VDDA.n336 GNDA 0.015208f
C3046 VDDA.n338 GNDA 0.013419f
C3047 VDDA.n339 GNDA 0.013419f
C3048 VDDA.n340 GNDA 0.016903f
C3049 VDDA.n342 GNDA 0.067862f
C3050 VDDA.t290 GNDA 0.05636f
C3051 VDDA.t211 GNDA 0.050609f
C3052 VDDA.t345 GNDA 0.05636f
C3053 VDDA.n344 GNDA 0.013419f
C3054 VDDA.n345 GNDA 0.013419f
C3055 VDDA.t347 GNDA 0.020216f
C3056 VDDA.n346 GNDA 0.01867f
C3057 VDDA.n348 GNDA 0.067862f
C3058 VDDA.n350 GNDA 0.016924f
C3059 VDDA.t344 GNDA 0.011158f
C3060 VDDA.n351 GNDA 0.015955f
C3061 VDDA.n352 GNDA 0.127592f
C3062 VDDA.n353 GNDA 0.072223f
C3063 VDDA.n354 GNDA 0.073372f
C3064 VDDA.n355 GNDA 0.015528f
C3065 VDDA.n356 GNDA 0.015528f
C3066 VDDA.n357 GNDA 0.015528f
C3067 VDDA.n358 GNDA 0.016103f
C3068 VDDA.n359 GNDA 0.016103f
C3069 VDDA.n360 GNDA 0.016103f
C3070 VDDA.n361 GNDA 0.016103f
C3071 VDDA.n362 GNDA 0.043793f
C3072 VDDA.n363 GNDA 0.016302f
C3073 VDDA.n364 GNDA 0.014668f
C3074 VDDA.n365 GNDA 1.59877f
C3075 VDDA.n366 GNDA 0.01294f
C3076 VDDA.n367 GNDA 0.01294f
C3077 VDDA.n368 GNDA 0.013419f
C3078 VDDA.n369 GNDA 0.011981f
C3079 VDDA.n372 GNDA 0.085294f
C3080 VDDA.t389 GNDA 0.013435f
C3081 VDDA.t329 GNDA 0.017269f
C3082 VDDA.n376 GNDA 0.08527f
C3083 VDDA.t194 GNDA 0.013985f
C3084 VDDA.t250 GNDA 0.013985f
C3085 VDDA.n378 GNDA 0.141964f
C3086 VDDA.t226 GNDA 0.013435f
C3087 VDDA.t363 GNDA 0.013435f
C3088 VDDA.n379 GNDA 0.016896f
C3089 VDDA.n380 GNDA 0.066813f
C3090 VDDA.t362 GNDA 0.04652f
C3091 VDDA.t293 GNDA 0.029522f
C3092 VDDA.t220 GNDA 0.029522f
C3093 VDDA.t225 GNDA 0.04652f
C3094 VDDA.n381 GNDA 0.066813f
C3095 VDDA.n382 GNDA 0.016297f
C3096 VDDA.n383 GNDA 0.107877f
C3097 VDDA.n385 GNDA 0.08527f
C3098 VDDA.n386 GNDA 0.105577f
C3099 VDDA.n387 GNDA 0.01631f
C3100 VDDA.n388 GNDA 0.039909f
C3101 VDDA.t249 GNDA 0.042059f
C3102 VDDA.t255 GNDA 0.029522f
C3103 VDDA.t196 GNDA 0.029522f
C3104 VDDA.t322 GNDA 0.029522f
C3105 VDDA.t252 GNDA 0.029522f
C3106 VDDA.t193 GNDA 0.042059f
C3107 VDDA.n389 GNDA 0.039909f
C3108 VDDA.n390 GNDA 0.01631f
C3109 VDDA.n391 GNDA 0.105577f
C3110 VDDA.n393 GNDA 0.074942f
C3111 VDDA.n394 GNDA 0.095225f
C3112 VDDA.n395 GNDA 0.016297f
C3113 VDDA.n396 GNDA 0.066813f
C3114 VDDA.t328 GNDA 0.04652f
C3115 VDDA.t263 GNDA 0.029522f
C3116 VDDA.t199 GNDA 0.029522f
C3117 VDDA.t325 GNDA 0.029522f
C3118 VDDA.t260 GNDA 0.029522f
C3119 VDDA.t384 GNDA 0.029522f
C3120 VDDA.t309 GNDA 0.029522f
C3121 VDDA.t312 GNDA 0.029522f
C3122 VDDA.t237 GNDA 0.029522f
C3123 VDDA.t387 GNDA 0.04652f
C3124 VDDA.n397 GNDA 0.066813f
C3125 VDDA.n398 GNDA 0.016297f
C3126 VDDA.n399 GNDA 0.01607f
C3127 VDDA.t335 GNDA 0.013978f
C3128 VDDA.t276 GNDA 0.013978f
C3129 VDDA.n402 GNDA 0.039917f
C3130 VDDA.t275 GNDA 0.042059f
C3131 VDDA.t205 GNDA 0.029522f
C3132 VDDA.t337 GNDA 0.029522f
C3133 VDDA.t272 GNDA 0.029522f
C3134 VDDA.t202 GNDA 0.029522f
C3135 VDDA.t334 GNDA 0.042059f
C3136 VDDA.n403 GNDA 0.039917f
C3137 VDDA.n404 GNDA 0.016595f
C3138 VDDA.n405 GNDA 0.135116f
C3139 VDDA.n406 GNDA 0.085274f
C3140 VDDA.n407 GNDA 0.105577f
C3141 VDDA.n408 GNDA 0.095225f
C3142 VDDA.n409 GNDA 0.074942f
C3143 VDDA.n410 GNDA 0.085294f
C3144 VDDA.n411 GNDA 0.050609f
C3145 VDDA.n412 GNDA 0.057403f
C3146 VDDA.n413 GNDA 0.015192f
C3147 VDDA.n417 GNDA 0.190011f
C3148 VDDA.t423 GNDA 0.066643f
C3149 VDDA.t25 GNDA 0.057271f
C3150 VDDA.n419 GNDA 0.15843f
C3151 VDDA.n421 GNDA 0.077485f
C3152 VDDA.n423 GNDA 0.077485f
C3153 VDDA.n425 GNDA 0.12247f
C3154 VDDA.n426 GNDA 0.551021f
C3155 VDDA.t210 GNDA 0.013632f
C3156 VDDA.n427 GNDA 0.312364f
C3157 VDDA.n431 GNDA 0.238506f
C3158 VDDA.n438 GNDA 0.010674f
C3159 VDDA.n439 GNDA 0.041387f
C3160 VDDA.n440 GNDA 0.028065f
C3161 VDDA.n441 GNDA 0.01294f
C3162 VDDA.n442 GNDA 0.01294f
C3163 VDDA.n443 GNDA 0.01294f
C3164 VDDA.n444 GNDA 0.013419f
C3165 VDDA.n445 GNDA 0.013419f
C3166 VDDA.n446 GNDA 0.013419f
C3167 VDDA.n447 GNDA 0.013419f
C3168 VDDA.n448 GNDA 0.013419f
C3169 VDDA.n449 GNDA 0.01294f
C3170 VDDA.t134 GNDA 0.013419f
C3171 VDDA.t142 GNDA 0.013419f
C3172 VDDA.n450 GNDA 0.028496f
C3173 VDDA.t118 GNDA 0.013419f
C3174 VDDA.t126 GNDA 0.013419f
C3175 VDDA.n451 GNDA 0.034061f
C3176 VDDA.n452 GNDA 0.095144f
C3177 VDDA.t339 GNDA 0.02353f
C3178 VDDA.t229 GNDA 0.047733f
C3179 VDDA.t116 GNDA 0.013419f
C3180 VDDA.t112 GNDA 0.013419f
C3181 VDDA.n453 GNDA 0.034061f
C3182 VDDA.n454 GNDA 0.106272f
C3183 VDDA.t227 GNDA 0.02353f
C3184 VDDA.n455 GNDA 0.069915f
C3185 VDDA.n456 GNDA 0.13847f
C3186 VDDA.t228 GNDA 0.114382f
C3187 VDDA.t115 GNDA 0.089715f
C3188 VDDA.t111 GNDA 0.089715f
C3189 VDDA.t117 GNDA 0.089715f
C3190 VDDA.t125 GNDA 0.089715f
C3191 VDDA.t133 GNDA 0.089715f
C3192 VDDA.t141 GNDA 0.089715f
C3193 VDDA.t107 GNDA 0.089715f
C3194 VDDA.t113 GNDA 0.089715f
C3195 VDDA.t121 GNDA 0.089715f
C3196 VDDA.t127 GNDA 0.089715f
C3197 VDDA.t340 GNDA 0.115877f
C3198 VDDA.t341 GNDA 0.047733f
C3199 VDDA.n457 GNDA 0.144451f
C3200 VDDA.n458 GNDA 0.069915f
C3201 VDDA.t122 GNDA 0.013419f
C3202 VDDA.t128 GNDA 0.013419f
C3203 VDDA.n459 GNDA 0.034061f
C3204 VDDA.n460 GNDA 0.106272f
C3205 VDDA.t108 GNDA 0.013419f
C3206 VDDA.t114 GNDA 0.013419f
C3207 VDDA.n461 GNDA 0.034061f
C3208 VDDA.n462 GNDA 0.095144f
C3209 VDDA.n463 GNDA 0.012269f
C3210 VDDA.n464 GNDA 0.105674f
C3211 VDDA.t102 GNDA 0.011502f
C3212 VDDA.t37 GNDA 0.011502f
C3213 VDDA.n465 GNDA 0.039415f
C3214 VDDA.t87 GNDA 0.011502f
C3215 VDDA.t407 GNDA 0.011502f
C3216 VDDA.n466 GNDA 0.038068f
C3217 VDDA.n467 GNDA 0.146038f
C3218 VDDA.t73 GNDA 0.011502f
C3219 VDDA.t405 GNDA 0.011502f
C3220 VDDA.n468 GNDA 0.038068f
C3221 VDDA.n469 GNDA 0.075034f
C3222 VDDA.t9 GNDA 0.011502f
C3223 VDDA.t408 GNDA 0.011502f
C3224 VDDA.n470 GNDA 0.038068f
C3225 VDDA.n471 GNDA 0.075034f
C3226 VDDA.t8 GNDA 0.011502f
C3227 VDDA.t91 GNDA 0.011502f
C3228 VDDA.n472 GNDA 0.038068f
C3229 VDDA.n473 GNDA 0.075034f
C3230 VDDA.t40 GNDA 0.011502f
C3231 VDDA.t99 GNDA 0.011502f
C3232 VDDA.n474 GNDA 0.038068f
C3233 VDDA.n475 GNDA 0.109928f
C3234 VDDA.t207 GNDA 0.011199f
C3235 VDDA.n476 GNDA 0.058561f
C3236 VDDA.t209 GNDA 0.027357f
C3237 VDDA.n477 GNDA 0.084043f
C3238 VDDA.t208 GNDA 0.068154f
C3239 VDDA.t96 GNDA 0.050609f
C3240 VDDA.t398 GNDA 0.050609f
C3241 VDDA.t36 GNDA 0.050609f
C3242 VDDA.t86 GNDA 0.050609f
C3243 VDDA.t406 GNDA 0.050609f
C3244 VDDA.t72 GNDA 0.050609f
C3245 VDDA.t95 GNDA 0.050609f
C3246 VDDA.t88 GNDA 0.050609f
C3247 VDDA.t94 GNDA 0.050609f
C3248 VDDA.t76 GNDA 0.050609f
C3249 VDDA.t234 GNDA 0.068154f
C3250 VDDA.t235 GNDA 0.027357f
C3251 VDDA.n478 GNDA 0.084043f
C3252 VDDA.t233 GNDA 0.011199f
C3253 VDDA.n479 GNDA 0.044725f
C3254 VDDA.n480 GNDA 0.059667f
C3255 VDDA.n481 GNDA 0.071277f
C3256 VDDA.n482 GNDA 0.048211f
C3257 VDDA.n483 GNDA 0.021777f
C3258 VDDA.t354 GNDA 0.028707f
C3259 VDDA.t13 GNDA 0.018978f
C3260 VDDA.t415 GNDA 0.018978f
C3261 VDDA.t58 GNDA 0.018978f
C3262 VDDA.t394 GNDA 0.018978f
C3263 VDDA.t85 GNDA 0.018978f
C3264 VDDA.t14 GNDA 0.018978f
C3265 VDDA.t66 GNDA 0.018978f
C3266 VDDA.t11 GNDA 0.018978f
C3267 VDDA.t64 GNDA 0.018978f
C3268 VDDA.t413 GNDA 0.018978f
C3269 VDDA.t381 GNDA 0.028707f
C3270 VDDA.n484 GNDA 0.021777f
C3271 VDDA.n485 GNDA 0.034421f
C3272 VDDA.n486 GNDA 0.068603f
C3273 VDDA.n487 GNDA 0.040959f
C3274 VDDA.t400 GNDA 0.023004f
C3275 VDDA.t98 GNDA 0.023004f
C3276 VDDA.n488 GNDA 0.068536f
C3277 VDDA.n489 GNDA 0.140609f
C3278 VDDA.t368 GNDA 0.080957f
C3279 VDDA.t402 GNDA 0.023004f
C3280 VDDA.t42 GNDA 0.023004f
C3281 VDDA.n490 GNDA 0.068536f
C3282 VDDA.n491 GNDA 0.140609f
C3283 VDDA.t410 GNDA 0.023004f
C3284 VDDA.t44 GNDA 0.023004f
C3285 VDDA.n492 GNDA 0.068536f
C3286 VDDA.n493 GNDA 0.140609f
C3287 VDDA.t90 GNDA 0.023004f
C3288 VDDA.t39 GNDA 0.023004f
C3289 VDDA.n494 GNDA 0.068536f
C3290 VDDA.n495 GNDA 0.140609f
C3291 VDDA.t404 GNDA 0.023004f
C3292 VDDA.t78 GNDA 0.023004f
C3293 VDDA.n496 GNDA 0.068536f
C3294 VDDA.n497 GNDA 0.148855f
C3295 VDDA.t366 GNDA 0.02791f
C3296 VDDA.n498 GNDA 0.063735f
C3297 VDDA.n499 GNDA 0.270807f
C3298 VDDA.t367 GNDA 0.175394f
C3299 VDDA.t403 GNDA 0.134957f
C3300 VDDA.t77 GNDA 0.134957f
C3301 VDDA.t89 GNDA 0.134957f
C3302 VDDA.t38 GNDA 0.134957f
C3303 VDDA.t409 GNDA 0.134957f
C3304 VDDA.t43 GNDA 0.134957f
C3305 VDDA.t401 GNDA 0.134957f
C3306 VDDA.t41 GNDA 0.134957f
C3307 VDDA.t399 GNDA 0.134957f
C3308 VDDA.t97 GNDA 0.134957f
C3309 VDDA.t391 GNDA 0.175394f
C3310 VDDA.t392 GNDA 0.080957f
C3311 VDDA.n500 GNDA 0.270807f
C3312 VDDA.t390 GNDA 0.02791f
C3313 VDDA.n501 GNDA 0.062758f
C3314 VDDA.n502 GNDA 0.013249f
C3315 VDDA.n504 GNDA 0.037483f
C3316 VDDA.n506 GNDA 0.037483f
C3317 VDDA.n508 GNDA 0.037483f
C3318 VDDA.n510 GNDA 0.037483f
C3319 VDDA.n512 GNDA 0.037483f
C3320 VDDA.n514 GNDA 0.037483f
C3321 VDDA.n516 GNDA 0.037483f
C3322 VDDA.n518 GNDA 0.037483f
C3323 VDDA.n520 GNDA 0.037483f
C3324 VDDA.n522 GNDA 0.046558f
C3325 VDDA.n523 GNDA 0.036075f
C3326 VDDA.n524 GNDA 0.021626f
C3327 VDDA.t269 GNDA 0.028707f
C3328 VDDA.t30 GNDA 0.018978f
C3329 VDDA.t23 GNDA 0.018978f
C3330 VDDA.t69 GNDA 0.018978f
C3331 VDDA.t45 GNDA 0.018978f
C3332 VDDA.t417 GNDA 0.018978f
C3333 VDDA.t67 GNDA 0.018978f
C3334 VDDA.t74 GNDA 0.018978f
C3335 VDDA.t55 GNDA 0.018978f
C3336 VDDA.t19 GNDA 0.018978f
C3337 VDDA.t47 GNDA 0.018978f
C3338 VDDA.t83 GNDA 0.018978f
C3339 VDDA.t59 GNDA 0.018978f
C3340 VDDA.t21 GNDA 0.018978f
C3341 VDDA.t1 GNDA 0.018978f
C3342 VDDA.t62 GNDA 0.018978f
C3343 VDDA.t4 GNDA 0.018978f
C3344 VDDA.t17 GNDA 0.018978f
C3345 VDDA.t81 GNDA 0.018978f
C3346 VDDA.t6 GNDA 0.018978f
C3347 VDDA.t49 GNDA 0.018978f
C3348 VDDA.t287 GNDA 0.028707f
C3349 VDDA.n525 GNDA 0.021626f
C3350 VDDA.n526 GNDA 0.035063f
C3351 VDDA.n527 GNDA 0.02849f
C3352 VDDA.n528 GNDA 0.028563f
C3353 VDDA.n529 GNDA 0.075923f
C3354 VDDA.n530 GNDA 0.098159f
C3355 VDDA.t130 GNDA 0.013419f
C3356 VDDA.t136 GNDA 0.013419f
C3357 VDDA.n531 GNDA 0.028496f
C3358 VDDA.t104 GNDA 0.013419f
C3359 VDDA.t124 GNDA 0.013419f
C3360 VDDA.n532 GNDA 0.034061f
C3361 VDDA.n533 GNDA 0.095144f
C3362 VDDA.t265 GNDA 0.02353f
C3363 VDDA.t352 GNDA 0.047733f
C3364 VDDA.t144 GNDA 0.013419f
C3365 VDDA.t138 GNDA 0.013419f
C3366 VDDA.n534 GNDA 0.034061f
C3367 VDDA.n535 GNDA 0.106272f
C3368 VDDA.t350 GNDA 0.02353f
C3369 VDDA.n536 GNDA 0.069915f
C3370 VDDA.n537 GNDA 0.13847f
C3371 VDDA.t351 GNDA 0.114382f
C3372 VDDA.t143 GNDA 0.089715f
C3373 VDDA.t137 GNDA 0.089715f
C3374 VDDA.t103 GNDA 0.089715f
C3375 VDDA.t123 GNDA 0.089715f
C3376 VDDA.t129 GNDA 0.089715f
C3377 VDDA.t135 GNDA 0.089715f
C3378 VDDA.t131 GNDA 0.089715f
C3379 VDDA.t139 GNDA 0.089715f
C3380 VDDA.t105 GNDA 0.089715f
C3381 VDDA.t109 GNDA 0.089715f
C3382 VDDA.t266 GNDA 0.114382f
C3383 VDDA.t267 GNDA 0.047733f
C3384 VDDA.n538 GNDA 0.13847f
C3385 VDDA.n539 GNDA 0.069915f
C3386 VDDA.t106 GNDA 0.013419f
C3387 VDDA.t110 GNDA 0.013419f
C3388 VDDA.n540 GNDA 0.034061f
C3389 VDDA.n541 GNDA 0.106272f
C3390 VDDA.t132 GNDA 0.013419f
C3391 VDDA.t140 GNDA 0.013419f
C3392 VDDA.n542 GNDA 0.034061f
C3393 VDDA.n543 GNDA 0.095144f
C3394 VDDA.n544 GNDA 0.012269f
C3395 VDDA.n545 GNDA 0.105674f
C3396 VDDA.t153 GNDA 0.011502f
C3397 VDDA.t101 GNDA 0.011502f
C3398 VDDA.n546 GNDA 0.039415f
C3399 VDDA.t165 GNDA 0.011502f
C3400 VDDA.t169 GNDA 0.011502f
C3401 VDDA.n547 GNDA 0.038068f
C3402 VDDA.n548 GNDA 0.146038f
C3403 VDDA.t170 GNDA 0.011502f
C3404 VDDA.t149 GNDA 0.011502f
C3405 VDDA.n549 GNDA 0.038068f
C3406 VDDA.n550 GNDA 0.075034f
C3407 VDDA.t174 GNDA 0.011502f
C3408 VDDA.t154 GNDA 0.011502f
C3409 VDDA.n551 GNDA 0.038068f
C3410 VDDA.n552 GNDA 0.075034f
C3411 VDDA.t162 GNDA 0.011502f
C3412 VDDA.t182 GNDA 0.011502f
C3413 VDDA.n553 GNDA 0.038068f
C3414 VDDA.n554 GNDA 0.075034f
C3415 VDDA.t100 GNDA 0.011502f
C3416 VDDA.t145 GNDA 0.011502f
C3417 VDDA.n555 GNDA 0.038068f
C3418 VDDA.n556 GNDA 0.109928f
C3419 VDDA.t356 GNDA 0.011199f
C3420 VDDA.n557 GNDA 0.058561f
C3421 VDDA.t358 GNDA 0.027357f
C3422 VDDA.n558 GNDA 0.084043f
C3423 VDDA.t357 GNDA 0.068154f
C3424 VDDA.t159 GNDA 0.050609f
C3425 VDDA.t181 GNDA 0.050609f
C3426 VDDA.t173 GNDA 0.050609f
C3427 VDDA.t155 GNDA 0.050609f
C3428 VDDA.t175 GNDA 0.050609f
C3429 VDDA.t156 GNDA 0.050609f
C3430 VDDA.t178 GNDA 0.050609f
C3431 VDDA.t148 GNDA 0.050609f
C3432 VDDA.t168 GNDA 0.050609f
C3433 VDDA.t152 GNDA 0.050609f
C3434 VDDA.t331 GNDA 0.068154f
C3435 VDDA.t332 GNDA 0.027357f
C3436 VDDA.n559 GNDA 0.084043f
C3437 VDDA.t330 GNDA 0.011199f
C3438 VDDA.n560 GNDA 0.044725f
C3439 VDDA.n561 GNDA 0.059667f
C3440 VDDA.n562 GNDA 0.071277f
C3441 VDDA.n563 GNDA 0.048211f
C3442 VDDA.n564 GNDA 0.021777f
C3443 VDDA.t372 GNDA 0.028707f
C3444 VDDA.t396 GNDA 0.018978f
C3445 VDDA.t421 GNDA 0.018978f
C3446 VDDA.t12 GNDA 0.018978f
C3447 VDDA.t34 GNDA 0.018978f
C3448 VDDA.t10 GNDA 0.018978f
C3449 VDDA.t414 GNDA 0.018978f
C3450 VDDA.t65 GNDA 0.018978f
C3451 VDDA.t92 GNDA 0.018978f
C3452 VDDA.t33 GNDA 0.018978f
C3453 VDDA.t420 GNDA 0.018978f
C3454 VDDA.t186 GNDA 0.028707f
C3455 VDDA.n565 GNDA 0.021777f
C3456 VDDA.n566 GNDA 0.034421f
C3457 VDDA.n567 GNDA 0.068327f
C3458 VDDA.n568 GNDA 0.040852f
C3459 VDDA.t180 GNDA 0.023004f
C3460 VDDA.t158 GNDA 0.023004f
C3461 VDDA.n569 GNDA 0.068536f
C3462 VDDA.n570 GNDA 0.140609f
C3463 VDDA.t307 GNDA 0.080957f
C3464 VDDA.t177 GNDA 0.023004f
C3465 VDDA.t167 GNDA 0.023004f
C3466 VDDA.n571 GNDA 0.068536f
C3467 VDDA.n572 GNDA 0.140609f
C3468 VDDA.t147 GNDA 0.023004f
C3469 VDDA.t164 GNDA 0.023004f
C3470 VDDA.n573 GNDA 0.068536f
C3471 VDDA.n574 GNDA 0.140609f
C3472 VDDA.t184 GNDA 0.023004f
C3473 VDDA.t161 GNDA 0.023004f
C3474 VDDA.n575 GNDA 0.068536f
C3475 VDDA.n576 GNDA 0.140609f
C3476 VDDA.t172 GNDA 0.023004f
C3477 VDDA.t151 GNDA 0.023004f
C3478 VDDA.n577 GNDA 0.068536f
C3479 VDDA.n578 GNDA 0.148855f
C3480 VDDA.t305 GNDA 0.02791f
C3481 VDDA.n579 GNDA 0.063735f
C3482 VDDA.n580 GNDA 0.270807f
C3483 VDDA.t306 GNDA 0.175394f
C3484 VDDA.t150 GNDA 0.134957f
C3485 VDDA.t171 GNDA 0.134957f
C3486 VDDA.t160 GNDA 0.134957f
C3487 VDDA.t183 GNDA 0.134957f
C3488 VDDA.t163 GNDA 0.134957f
C3489 VDDA.t146 GNDA 0.134957f
C3490 VDDA.t166 GNDA 0.134957f
C3491 VDDA.t176 GNDA 0.134957f
C3492 VDDA.t157 GNDA 0.134957f
C3493 VDDA.t179 GNDA 0.134957f
C3494 VDDA.t278 GNDA 0.175394f
C3495 VDDA.t279 GNDA 0.080957f
C3496 VDDA.n581 GNDA 0.270807f
C3497 VDDA.t277 GNDA 0.02791f
C3498 VDDA.n582 GNDA 0.062758f
C3499 VDDA.n583 GNDA 0.021906f
C3500 VDDA.n584 GNDA 0.077426f
C3501 VDDA.n585 GNDA 0.097968f
C3502 VDDA.n586 GNDA 0.095778f
C3503 VDDA.n587 GNDA 0.01561f
C3504 VDDA.n588 GNDA 0.062241f
C3505 VDDA.t230 GNDA 0.014423f
C3506 VDDA.t247 GNDA 0.02491f
C3507 VDDA.t244 GNDA 0.014423f
C3508 VDDA.n589 GNDA 0.038183f
C3509 VDDA.n590 GNDA 0.074999f
C3510 VDDA.t245 GNDA 0.06677f
C3511 VDDA.t15 GNDA 0.050609f
C3512 VDDA.t231 GNDA 0.06677f
C3513 VDDA.t232 GNDA 0.02491f
C3514 VDDA.n591 GNDA 0.074999f
C3515 VDDA.n592 GNDA 0.03782f
C3516 VDDA.n593 GNDA 0.021884f
C3517 VDDA.n594 GNDA 0.038957f
C3518 VDDA.n595 GNDA 0.096283f
C3519 VDDA.t314 GNDA 0.023763f
C3520 VDDA.t120 GNDA 0.013419f
C3521 VDDA.n596 GNDA 0.033709f
C3522 VDDA.t243 GNDA 0.061152f
C3523 VDDA.t241 GNDA 0.023763f
C3524 VDDA.n597 GNDA 0.050193f
C3525 VDDA.n598 GNDA 0.152676f
C3526 VDDA.t242 GNDA 0.114382f
C3527 VDDA.t119 GNDA 0.089715f
C3528 VDDA.t315 GNDA 0.114382f
C3529 VDDA.t316 GNDA 0.047733f
C3530 VDDA.n599 GNDA 0.152676f
C3531 VDDA.n600 GNDA 0.049829f
C3532 VDDA.n601 GNDA 0.021884f
C3533 VDDA.n602 GNDA 0.07137f
C3534 VDDA.n603 GNDA 0.070553f
C3535 VDDA.n604 GNDA 0.011981f
C3536 VDDA.n605 GNDA 0.011981f
C3537 VDDA.n606 GNDA 2.3464f
C3538 VDDA.n607 GNDA 0.015528f
C3539 VDDA.n608 GNDA 0.015528f
C3540 VDDA.n609 GNDA 0.016103f
C3541 VDDA.n610 GNDA 0.016103f
C3542 VDDA.n611 GNDA 0.016103f
C3543 VDDA.n612 GNDA 0.016103f
C3544 VDDA.n613 GNDA 0.016103f
C3545 VDDA.n614 GNDA 0.043793f
C3546 VDDA.n615 GNDA 0.016302f
C3547 VDDA.n616 GNDA 0.014668f
C3548 VDDA.n617 GNDA 1.62561f
C3549 VDDA.n618 GNDA 0.014377f
C3550 VDDA.n619 GNDA 0.014377f
C3551 VDDA.n620 GNDA 0.140769f
C3552 VDDA.t188 GNDA 0.15336f
C3553 VDDA.t282 GNDA 0.155972f
C3554 VDDA.t239 GNDA 0.15336f
C3555 VDDA.n621 GNDA 0.102823f
C3556 VDDA.t297 GNDA 0.15336f
C3557 VDDA.t364 GNDA 0.155972f
C3558 VDDA.n622 GNDA 0.131578f
C3559 VDDA.t303 GNDA 0.155972f
C3560 VDDA.t317 GNDA 0.15336f
C3561 VDDA.n623 GNDA 0.102823f
C3562 VDDA.t342 GNDA 0.15336f
C3563 VDDA.t213 GNDA 0.155972f
C3564 VDDA.n624 GNDA 0.160333f
C3565 VDDA.t295 GNDA 0.155972f
C3566 VDDA.t257 GNDA 0.15336f
C3567 VDDA.n625 GNDA 0.102823f
C3568 VDDA.t299 GNDA 0.15336f
C3569 VDDA.t374 GNDA 0.155972f
C3570 VDDA.n626 GNDA 0.160333f
C3571 VDDA.t348 GNDA 0.155972f
C3572 VDDA.t301 GNDA 0.15336f
C3573 VDDA.n627 GNDA 0.102823f
C3574 VDDA.t376 GNDA 0.15336f
C3575 VDDA.t215 GNDA 0.155972f
C3576 VDDA.n628 GNDA 0.160333f
C3577 VDDA.t280 GNDA 0.155972f
C3578 VDDA.t217 GNDA 0.15336f
C3579 VDDA.n629 GNDA 0.131578f
C3580 VDDA.t378 GNDA 0.15336f
C3581 VDDA.n630 GNDA 0.067095f
C3582 VDDA.n631 GNDA 0.229746f
C3583 VDDA.t52 GNDA 0.043154f
C3584 VDDA.n632 GNDA 0.269283f
C3585 VDDA.n633 GNDA 0.279962f
C3586 VDDA.n635 GNDA 0.078745f
C3587 VDDA.n639 GNDA 0.092288f
C3588 VDDA.n640 GNDA 0.061423f
C3589 VDDA.n641 GNDA 0.030672f
C3590 VDDA.n643 GNDA 0.052948f
C3591 VDDA.n645 GNDA 0.052444f
C3592 VDDA.n646 GNDA 0.135434f
C3593 VDDA.n648 GNDA 0.020022f
C3594 VDDA.n649 GNDA 0.02147f
C3595 VDDA.n650 GNDA 0.02147f
C3596 VDDA.n651 GNDA 0.02147f
C3597 VDDA.n652 GNDA 0.02147f
C3598 VDDA.n653 GNDA 0.02147f
C3599 VDDA.n654 GNDA 0.02147f
C3600 VDDA.n655 GNDA 0.020022f
C3601 VDDA.t457 GNDA 0.04639f
C3602 two_stage_opamp_dummy_magic_23_0.Y.t17 GNDA 0.037911f
C3603 two_stage_opamp_dummy_magic_23_0.Y.t12 GNDA 0.037911f
C3604 two_stage_opamp_dummy_magic_23_0.Y.n0 GNDA 0.082489f
C3605 two_stage_opamp_dummy_magic_23_0.Y.n1 GNDA 0.256901f
C3606 two_stage_opamp_dummy_magic_23_0.Y.n2 GNDA 0.080625f
C3607 two_stage_opamp_dummy_magic_23_0.Y.t19 GNDA 0.037911f
C3608 two_stage_opamp_dummy_magic_23_0.Y.t24 GNDA 0.037911f
C3609 two_stage_opamp_dummy_magic_23_0.Y.n3 GNDA 0.082489f
C3610 two_stage_opamp_dummy_magic_23_0.Y.n4 GNDA 0.327754f
C3611 two_stage_opamp_dummy_magic_23_0.Y.t23 GNDA 0.037911f
C3612 two_stage_opamp_dummy_magic_23_0.Y.t0 GNDA 0.037911f
C3613 two_stage_opamp_dummy_magic_23_0.Y.n5 GNDA 0.082489f
C3614 two_stage_opamp_dummy_magic_23_0.Y.n6 GNDA 0.327754f
C3615 two_stage_opamp_dummy_magic_23_0.Y.n7 GNDA 0.137048f
C3616 two_stage_opamp_dummy_magic_23_0.Y.t11 GNDA 0.037911f
C3617 two_stage_opamp_dummy_magic_23_0.Y.t8 GNDA 0.037911f
C3618 two_stage_opamp_dummy_magic_23_0.Y.n8 GNDA 0.082489f
C3619 two_stage_opamp_dummy_magic_23_0.Y.n9 GNDA 0.314545f
C3620 two_stage_opamp_dummy_magic_23_0.Y.n10 GNDA 0.144975f
C3621 two_stage_opamp_dummy_magic_23_0.Y.t9 GNDA 0.037911f
C3622 two_stage_opamp_dummy_magic_23_0.Y.t7 GNDA 0.037911f
C3623 two_stage_opamp_dummy_magic_23_0.Y.n11 GNDA 0.082489f
C3624 two_stage_opamp_dummy_magic_23_0.Y.n12 GNDA 0.314545f
C3625 two_stage_opamp_dummy_magic_23_0.Y.n13 GNDA 0.084683f
C3626 two_stage_opamp_dummy_magic_23_0.Y.n14 GNDA 0.084683f
C3627 two_stage_opamp_dummy_magic_23_0.Y.n15 GNDA 0.144975f
C3628 two_stage_opamp_dummy_magic_23_0.Y.t18 GNDA 0.037911f
C3629 two_stage_opamp_dummy_magic_23_0.Y.t13 GNDA 0.037911f
C3630 two_stage_opamp_dummy_magic_23_0.Y.n16 GNDA 0.082489f
C3631 two_stage_opamp_dummy_magic_23_0.Y.n17 GNDA 0.314545f
C3632 two_stage_opamp_dummy_magic_23_0.Y.n18 GNDA 0.137048f
C3633 two_stage_opamp_dummy_magic_23_0.Y.n19 GNDA 0.075821f
C3634 two_stage_opamp_dummy_magic_23_0.Y.n20 GNDA 0.3074f
C3635 two_stage_opamp_dummy_magic_23_0.Y.t5 GNDA 0.088458f
C3636 two_stage_opamp_dummy_magic_23_0.Y.t10 GNDA 0.088458f
C3637 two_stage_opamp_dummy_magic_23_0.Y.n21 GNDA 0.180951f
C3638 two_stage_opamp_dummy_magic_23_0.Y.n22 GNDA 0.492191f
C3639 two_stage_opamp_dummy_magic_23_0.Y.n23 GNDA 0.095948f
C3640 two_stage_opamp_dummy_magic_23_0.Y.n24 GNDA 0.163678f
C3641 two_stage_opamp_dummy_magic_23_0.Y.t20 GNDA 0.088458f
C3642 two_stage_opamp_dummy_magic_23_0.Y.t4 GNDA 0.088458f
C3643 two_stage_opamp_dummy_magic_23_0.Y.n25 GNDA 0.180951f
C3644 two_stage_opamp_dummy_magic_23_0.Y.n26 GNDA 0.585864f
C3645 two_stage_opamp_dummy_magic_23_0.Y.t2 GNDA 0.088458f
C3646 two_stage_opamp_dummy_magic_23_0.Y.t22 GNDA 0.088458f
C3647 two_stage_opamp_dummy_magic_23_0.Y.n27 GNDA 0.180951f
C3648 two_stage_opamp_dummy_magic_23_0.Y.n28 GNDA 0.569865f
C3649 two_stage_opamp_dummy_magic_23_0.Y.n29 GNDA 0.163678f
C3650 two_stage_opamp_dummy_magic_23_0.Y.n30 GNDA 0.095948f
C3651 two_stage_opamp_dummy_magic_23_0.Y.t15 GNDA 0.088458f
C3652 two_stage_opamp_dummy_magic_23_0.Y.t3 GNDA 0.088458f
C3653 two_stage_opamp_dummy_magic_23_0.Y.n31 GNDA 0.180951f
C3654 two_stage_opamp_dummy_magic_23_0.Y.n32 GNDA 0.569865f
C3655 two_stage_opamp_dummy_magic_23_0.Y.n33 GNDA 0.095948f
C3656 two_stage_opamp_dummy_magic_23_0.Y.t1 GNDA 0.088458f
C3657 two_stage_opamp_dummy_magic_23_0.Y.t14 GNDA 0.088458f
C3658 two_stage_opamp_dummy_magic_23_0.Y.n34 GNDA 0.180951f
C3659 two_stage_opamp_dummy_magic_23_0.Y.n35 GNDA 0.569865f
C3660 two_stage_opamp_dummy_magic_23_0.Y.n36 GNDA 0.095948f
C3661 two_stage_opamp_dummy_magic_23_0.Y.n37 GNDA 0.163678f
C3662 two_stage_opamp_dummy_magic_23_0.Y.t6 GNDA 0.088458f
C3663 two_stage_opamp_dummy_magic_23_0.Y.t21 GNDA 0.088458f
C3664 two_stage_opamp_dummy_magic_23_0.Y.n38 GNDA 0.180951f
C3665 two_stage_opamp_dummy_magic_23_0.Y.n39 GNDA 0.569865f
C3666 two_stage_opamp_dummy_magic_23_0.Y.n40 GNDA 0.149208f
C3667 two_stage_opamp_dummy_magic_23_0.Y.n41 GNDA 0.48498f
C3668 two_stage_opamp_dummy_magic_23_0.Y.t52 GNDA 0.053075f
C3669 two_stage_opamp_dummy_magic_23_0.Y.t29 GNDA 0.053075f
C3670 two_stage_opamp_dummy_magic_23_0.Y.t45 GNDA 0.053075f
C3671 two_stage_opamp_dummy_magic_23_0.Y.t31 GNDA 0.053075f
C3672 two_stage_opamp_dummy_magic_23_0.Y.t46 GNDA 0.053075f
C3673 two_stage_opamp_dummy_magic_23_0.Y.t34 GNDA 0.053075f
C3674 two_stage_opamp_dummy_magic_23_0.Y.t27 GNDA 0.053075f
C3675 two_stage_opamp_dummy_magic_23_0.Y.t43 GNDA 0.064448f
C3676 two_stage_opamp_dummy_magic_23_0.Y.n42 GNDA 0.064448f
C3677 two_stage_opamp_dummy_magic_23_0.Y.n43 GNDA 0.041702f
C3678 two_stage_opamp_dummy_magic_23_0.Y.n44 GNDA 0.041702f
C3679 two_stage_opamp_dummy_magic_23_0.Y.n45 GNDA 0.041702f
C3680 two_stage_opamp_dummy_magic_23_0.Y.n46 GNDA 0.041702f
C3681 two_stage_opamp_dummy_magic_23_0.Y.n47 GNDA 0.041702f
C3682 two_stage_opamp_dummy_magic_23_0.Y.n48 GNDA 0.033646f
C3683 two_stage_opamp_dummy_magic_23_0.Y.t37 GNDA 0.053075f
C3684 two_stage_opamp_dummy_magic_23_0.Y.t49 GNDA 0.064448f
C3685 two_stage_opamp_dummy_magic_23_0.Y.n49 GNDA 0.056392f
C3686 two_stage_opamp_dummy_magic_23_0.Y.n50 GNDA 0.021219f
C3687 two_stage_opamp_dummy_magic_23_0.Y.t26 GNDA 0.081508f
C3688 two_stage_opamp_dummy_magic_23_0.Y.t33 GNDA 0.081508f
C3689 two_stage_opamp_dummy_magic_23_0.Y.t48 GNDA 0.081508f
C3690 two_stage_opamp_dummy_magic_23_0.Y.t36 GNDA 0.081508f
C3691 two_stage_opamp_dummy_magic_23_0.Y.t51 GNDA 0.081508f
C3692 two_stage_opamp_dummy_magic_23_0.Y.t39 GNDA 0.081508f
C3693 two_stage_opamp_dummy_magic_23_0.Y.t32 GNDA 0.081508f
C3694 two_stage_opamp_dummy_magic_23_0.Y.t47 GNDA 0.092661f
C3695 two_stage_opamp_dummy_magic_23_0.Y.n51 GNDA 0.083624f
C3696 two_stage_opamp_dummy_magic_23_0.Y.n52 GNDA 0.05118f
C3697 two_stage_opamp_dummy_magic_23_0.Y.n53 GNDA 0.05118f
C3698 two_stage_opamp_dummy_magic_23_0.Y.n54 GNDA 0.05118f
C3699 two_stage_opamp_dummy_magic_23_0.Y.n55 GNDA 0.05118f
C3700 two_stage_opamp_dummy_magic_23_0.Y.n56 GNDA 0.05118f
C3701 two_stage_opamp_dummy_magic_23_0.Y.n57 GNDA 0.043123f
C3702 two_stage_opamp_dummy_magic_23_0.Y.t41 GNDA 0.081508f
C3703 two_stage_opamp_dummy_magic_23_0.Y.t54 GNDA 0.092661f
C3704 two_stage_opamp_dummy_magic_23_0.Y.n58 GNDA 0.075568f
C3705 two_stage_opamp_dummy_magic_23_0.Y.n59 GNDA 0.021219f
C3706 two_stage_opamp_dummy_magic_23_0.Y.n60 GNDA 0.091639f
C3707 two_stage_opamp_dummy_magic_23_0.Y.n61 GNDA 1.04027f
C3708 two_stage_opamp_dummy_magic_23_0.Y.n62 GNDA 0.450882f
C3709 two_stage_opamp_dummy_magic_23_0.Y.t42 GNDA 0.166807f
C3710 two_stage_opamp_dummy_magic_23_0.Y.t35 GNDA 0.166807f
C3711 two_stage_opamp_dummy_magic_23_0.Y.t50 GNDA 0.177661f
C3712 two_stage_opamp_dummy_magic_23_0.Y.n63 GNDA 0.140789f
C3713 two_stage_opamp_dummy_magic_23_0.Y.n64 GNDA 0.071557f
C3714 two_stage_opamp_dummy_magic_23_0.Y.t25 GNDA 0.166807f
C3715 two_stage_opamp_dummy_magic_23_0.Y.t40 GNDA 0.166807f
C3716 two_stage_opamp_dummy_magic_23_0.Y.t53 GNDA 0.166807f
C3717 two_stage_opamp_dummy_magic_23_0.Y.t38 GNDA 0.166807f
C3718 two_stage_opamp_dummy_magic_23_0.Y.t30 GNDA 0.166807f
C3719 two_stage_opamp_dummy_magic_23_0.Y.t44 GNDA 0.166807f
C3720 two_stage_opamp_dummy_magic_23_0.Y.t28 GNDA 0.177661f
C3721 two_stage_opamp_dummy_magic_23_0.Y.n65 GNDA 0.140789f
C3722 two_stage_opamp_dummy_magic_23_0.Y.n66 GNDA 0.079613f
C3723 two_stage_opamp_dummy_magic_23_0.Y.n67 GNDA 0.079613f
C3724 two_stage_opamp_dummy_magic_23_0.Y.n68 GNDA 0.079613f
C3725 two_stage_opamp_dummy_magic_23_0.Y.n69 GNDA 0.079613f
C3726 two_stage_opamp_dummy_magic_23_0.Y.n70 GNDA 0.071557f
C3727 two_stage_opamp_dummy_magic_23_0.Y.n71 GNDA 0.036197f
C3728 two_stage_opamp_dummy_magic_23_0.Y.n72 GNDA 1.26467f
C3729 two_stage_opamp_dummy_magic_23_0.Y.t16 GNDA 1.21199f
C3730 two_stage_opamp_dummy_magic_23_0.Vb3.t5 GNDA 0.01662f
C3731 two_stage_opamp_dummy_magic_23_0.Vb3.t2 GNDA 0.01662f
C3732 two_stage_opamp_dummy_magic_23_0.Vb3.n0 GNDA 0.053535f
C3733 two_stage_opamp_dummy_magic_23_0.Vb3.t7 GNDA 0.01662f
C3734 two_stage_opamp_dummy_magic_23_0.Vb3.t6 GNDA 0.01662f
C3735 two_stage_opamp_dummy_magic_23_0.Vb3.n1 GNDA 0.053535f
C3736 two_stage_opamp_dummy_magic_23_0.Vb3.n2 GNDA 0.295139f
C3737 two_stage_opamp_dummy_magic_23_0.Vb3.t3 GNDA 0.01662f
C3738 two_stage_opamp_dummy_magic_23_0.Vb3.t0 GNDA 0.01662f
C3739 two_stage_opamp_dummy_magic_23_0.Vb3.n3 GNDA 0.0502f
C3740 two_stage_opamp_dummy_magic_23_0.Vb3.n4 GNDA 0.975504f
C3741 two_stage_opamp_dummy_magic_23_0.Vb3.t4 GNDA 0.058171f
C3742 two_stage_opamp_dummy_magic_23_0.Vb3.t1 GNDA 0.058171f
C3743 two_stage_opamp_dummy_magic_23_0.Vb3.n5 GNDA 0.160478f
C3744 two_stage_opamp_dummy_magic_23_0.Vb3.t9 GNDA 0.08227f
C3745 two_stage_opamp_dummy_magic_23_0.Vb3.t26 GNDA 0.08227f
C3746 two_stage_opamp_dummy_magic_23_0.Vb3.t23 GNDA 0.08227f
C3747 two_stage_opamp_dummy_magic_23_0.Vb3.t19 GNDA 0.08227f
C3748 two_stage_opamp_dummy_magic_23_0.Vb3.t16 GNDA 0.094939f
C3749 two_stage_opamp_dummy_magic_23_0.Vb3.n6 GNDA 0.07708f
C3750 two_stage_opamp_dummy_magic_23_0.Vb3.n7 GNDA 0.047368f
C3751 two_stage_opamp_dummy_magic_23_0.Vb3.n8 GNDA 0.047368f
C3752 two_stage_opamp_dummy_magic_23_0.Vb3.n9 GNDA 0.041532f
C3753 two_stage_opamp_dummy_magic_23_0.Vb3.t13 GNDA 0.08227f
C3754 two_stage_opamp_dummy_magic_23_0.Vb3.t17 GNDA 0.08227f
C3755 two_stage_opamp_dummy_magic_23_0.Vb3.t21 GNDA 0.08227f
C3756 two_stage_opamp_dummy_magic_23_0.Vb3.t24 GNDA 0.08227f
C3757 two_stage_opamp_dummy_magic_23_0.Vb3.t22 GNDA 0.094939f
C3758 two_stage_opamp_dummy_magic_23_0.Vb3.n10 GNDA 0.07708f
C3759 two_stage_opamp_dummy_magic_23_0.Vb3.n11 GNDA 0.047368f
C3760 two_stage_opamp_dummy_magic_23_0.Vb3.n12 GNDA 0.047368f
C3761 two_stage_opamp_dummy_magic_23_0.Vb3.n13 GNDA 0.041532f
C3762 two_stage_opamp_dummy_magic_23_0.Vb3.n14 GNDA 0.041916f
C3763 two_stage_opamp_dummy_magic_23_0.Vb3.t12 GNDA 0.08227f
C3764 two_stage_opamp_dummy_magic_23_0.Vb3.t14 GNDA 0.08227f
C3765 two_stage_opamp_dummy_magic_23_0.Vb3.t10 GNDA 0.08227f
C3766 two_stage_opamp_dummy_magic_23_0.Vb3.t27 GNDA 0.08227f
C3767 two_stage_opamp_dummy_magic_23_0.Vb3.t25 GNDA 0.094939f
C3768 two_stage_opamp_dummy_magic_23_0.Vb3.n15 GNDA 0.07708f
C3769 two_stage_opamp_dummy_magic_23_0.Vb3.n16 GNDA 0.047368f
C3770 two_stage_opamp_dummy_magic_23_0.Vb3.n17 GNDA 0.047368f
C3771 two_stage_opamp_dummy_magic_23_0.Vb3.n18 GNDA 0.041532f
C3772 two_stage_opamp_dummy_magic_23_0.Vb3.t15 GNDA 0.08227f
C3773 two_stage_opamp_dummy_magic_23_0.Vb3.t18 GNDA 0.08227f
C3774 two_stage_opamp_dummy_magic_23_0.Vb3.t28 GNDA 0.08227f
C3775 two_stage_opamp_dummy_magic_23_0.Vb3.t11 GNDA 0.08227f
C3776 two_stage_opamp_dummy_magic_23_0.Vb3.t8 GNDA 0.094939f
C3777 two_stage_opamp_dummy_magic_23_0.Vb3.n19 GNDA 0.07708f
C3778 two_stage_opamp_dummy_magic_23_0.Vb3.n20 GNDA 0.047368f
C3779 two_stage_opamp_dummy_magic_23_0.Vb3.n21 GNDA 0.047368f
C3780 two_stage_opamp_dummy_magic_23_0.Vb3.n22 GNDA 0.041532f
C3781 two_stage_opamp_dummy_magic_23_0.Vb3.n23 GNDA 0.042678f
C3782 two_stage_opamp_dummy_magic_23_0.Vb3.n24 GNDA 1.40034f
C3783 two_stage_opamp_dummy_magic_23_0.Vb3.t20 GNDA 0.107472f
C3784 two_stage_opamp_dummy_magic_23_0.Vb3.n25 GNDA 0.377587f
C3785 two_stage_opamp_dummy_magic_23_0.Vb3.n26 GNDA 1.2975f
C3786 bgr_11_0.VB3_CUR_BIAS GNDA 2.07858f
.ends

