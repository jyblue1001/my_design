* PEX produced on Sun Feb 23 05:28:58 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from full_pll_magic_2.ext - technology: sky130A

.subckt full_pll_magic V_OSC VDDA GNDA F_REF I_IN
X0 GNDA.t168 a_6200_5250.t4 a_6200_5250.t5 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X1 a_5970_4630.t7 V_CONT.t8 a_6200_5250.t0 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 GNDA.t210 GNDA.t208 GNDA.t210 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X3 a_7630_n1440.t0 VCO_FD_magic_0.div120_2_0.div2.t2 GNDA.t265 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 a_870_1400.t1 pfd_8_0.QA_b.t3 VDDA.t214 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X5 pfd_8_0.DOWN_b.t1 VDDA.t221 pfd_8_0.DOWN_PFD_b.t2 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 GNDA.t241 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t1 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t0 VCO_FD_magic_0.div120_2_0.div24.t3 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 GNDA.t85 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t1 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X9 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t2 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X10 pfd_8_0.UP_input.t3 pfd_8_0.UP_b.t1 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X11 VDDA.t100 VCO_FD_magic_0.vco2_3_0.V1.t3 VCO_FD_magic_0.vco2_3_0.V4.t0 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X12 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t3 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 VDDA.t92 pfd_8_0.opamp_out.t10 opamp_cell_4_0.VIN+.t3 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X14 opamp_cell_4_0.n_right.t2 opamp_cell_4_0.VIN+.t6 a_6320_5840.t3 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X15 opamp_cell_4_0.n_right.t0 opamp_cell_4_0.n_left.t6 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X16 pfd_8_0.opamp_out.t5 opamp_cell_4_0.n_right.t5 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X17 GNDA.t56 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t4 VCO_FD_magic_0.div120_2_0.div8.t0 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 pfd_8_0.opamp_out.t9 a_6490_4630.t5 GNDA.t158 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X19 a_2350_1400.t0 pfd_8_0.before_Reset.t3 GNDA.t239 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X20 VDDA.t152 GNDA.t270 VCO_FD_magic_0.vco2_3_0.V4.t2 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X21 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t3 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X22 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t0 a_7630_n1440.t3 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t0 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X23 VDDA.t141 opamp_cell_4_0.p_bias.t6 opamp_cell_4_0.p_bias.t7 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X24 a_n30_1400.t0 F_REF.t0 VDDA.t132 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X25 GNDA.t136 I_IN.t2 I_IN.t3 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X26 VDDA.t66 VCO_FD_magic_0.div120_2_0.div4.t2 a_6330_n1440.t2 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 GNDA.t246 pfd_8_0.QA.t3 pfd_8_0.QA_b.t2 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 a_6200_5250.t3 a_6200_5250.t2 GNDA.t166 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X29 a_6200_5250.t1 V_CONT.t9 a_5970_4630.t6 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X30 VDDA.t139 opamp_cell_4_0.p_bias.t9 a_5970_4630.t5 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X31 VDDA.t191 VDDA.t188 VDDA.t190 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X32 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t3 a_8930_n1440.t3 GNDA.t248 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X33 VDDA.t187 VDDA.t185 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X34 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t4 I_IN.t5 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X35 VDDA.t195 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t0 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X36 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t0 VCO_FD_magic_0.div120_2_0.div8.t2 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X37 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t4 GNDA.t212 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X38 a_1910_2020.t1 pfd_8_0.QB.t3 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X39 VDDA.t204 pfd_8_0.UP_input.t4 V_CONT.t7 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X40 a_6220_5810.t7 a_6220_5810.t6 GNDA.t251 GNDA.t250 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X41 GNDA.t20 a_7630_n1440.t4 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t2 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X42 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t2 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X43 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t2 VCO_FD_magic_0.div120_2_0.div8.t3 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X44 GNDA.t223 F_VCO.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t1 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X45 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t2 VCO_FD_magic_0.div120_2_0.div24.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 a_8930_n1440.t0 V_OSC.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 VDDA.t82 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t2 F_VCO.t1 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X48 a_8930_n1440.t2 V_OSC.t3 GNDA.t140 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X49 GNDA.t74 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t1 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X50 a_6320_5840.t9 a_6220_5810.t9 GNDA.t89 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X51 pfd_8_0.QA.t2 pfd_8_0.QA_b.t4 GNDA.t235 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X52 pfd_8_0.UP_input.t1 pfd_8_0.UP.t2 pfd_8_0.opamp_out.t4 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X53 VDDA.t117 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t2 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X54 a_5970_4630.t3 opamp_cell_4_0.p_bias.t10 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X55 a_1390_1400.t1 pfd_8_0.E.t3 pfd_8_0.E_b.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X56 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN.t3 I_IN.t4 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X57 a_870_640.t1 pfd_8_0.QB_b.t3 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X58 I_IN.t1 I_IN.t0 GNDA.t126 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X59 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t1 F_VCO.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t0 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X60 VDDA.t184 VDDA.t181 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X61 VDDA.t84 a_2530_190.t2 a_2200_190.t1 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X62 V_CONT.t1 loop_filter_2_0.R1_C1.t0 GNDA.t67 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X63 pfd_8_0.opamp_out.t11 a_9360_3514.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X64 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t4 VDDA.t202 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X65 GNDA.t207 GNDA.t205 GNDA.t207 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X66 GNDA.t204 GNDA.t201 GNDA.t203 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X67 opamp_cell_4_0.p_bias.t5 opamp_cell_4_0.p_bias.t4 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X68 VCO_FD_magic_0.vco2_3_0.V1.t2 V_CONT.t10 GNDA.t6 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X69 VCO_FD_magic_0.vco2_3_0.V8.t1 VCO_FD_magic_0.vco2_3_0.V9.t2 VCO_FD_magic_0.vco2_3_0.V4.t1 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X70 V_CONT.t2 pfd_8_0.UP_input.t5 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X71 VDDA.t180 VDDA.t178 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X72 V_OSC.t0 VCO_FD_magic_0.vco2_3_0.V8.t2 VCO_FD_magic_0.vco2_3_0.V3.t0 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X73 GNDA.t200 GNDA.t197 GNDA.t199 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X74 pfd_8_0.F.t1 pfd_8_0.QB_b.t4 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X75 GNDA.t82 a_2530_190.t3 a_2200_190.t0 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X76 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN_b.t5 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X77 GNDA.t144 VCO_FD_magic_0.div120_2_0.div24.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t2 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X78 GNDA.t50 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t4 VCO_FD_magic_0.div120_2_0.div4.t1 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X79 GNDA.t196 GNDA.t193 GNDA.t195 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X80 VDDA.t211 a_8930_n1440.t4 VCO_FD_magic_0.div120_2_0.div2.t1 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X81 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t0 a_8930_n1440.t5 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t0 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X82 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t2 GNDA.t138 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X83 GNDA.t225 pfd_8_0.E_b.t3 pfd_8_0.E.t2 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X84 pfd_8_0.UP_b.t0 pfd_8_0.UP.t3 GNDA.t91 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X85 GNDA.t117 VDDA.t222 VCO_FD_magic_0.vco2_3_0.V3.t2 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X86 GNDA.t215 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t3 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X87 pfd_8_0.opamp_out.t12 a_9360_6440.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X88 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t0 VCO_FD_magic_0.div120_2_0.div8.t4 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X89 GNDA.t219 a_6220_5810.t10 a_6320_5840.t12 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X90 a_1390_640.t1 pfd_8_0.F.t3 pfd_8_0.F_b.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X91 GNDA.t192 GNDA.t189 GNDA.t191 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X92 GNDA.t30 F_VCO.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t1 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X93 VDDA.t147 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t1 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X94 a_2350_1400.t1 pfd_8_0.before_Reset.t4 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X95 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t1 F_VCO.t5 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X96 GNDA.t261 a_6220_5810.t4 a_6220_5810.t5 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X97 GNDA.t188 GNDA.t185 GNDA.t187 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X98 VDDA.t23 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t3 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X99 GNDA.t184 GNDA.t182 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X100 a_5970_4630.t12 a_5970_4630.t11 a_5970_4630.t12 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X101 VDDA.t88 pfd_8_0.UP_input.t6 V_CONT.t3 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X102 pfd_8_0.F_b.t2 pfd_8_0.F.t4 GNDA.t263 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X103 VDDA.t102 pfd_8_0.F.t5 a_490_640.t1 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X104 GNDA.t271 loop_filter_2_0.R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X105 VDDA.t177 VDDA.t175 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X106 pfd_8_0.QA_b.t0 pfd_8_0.QA.t4 a_n30_1400.t1 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X107 GNDA.t181 GNDA.t179 GNDA.t181 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X108 GNDA.t99 VCO_FD_magic_0.div120_2_0.div8.t5 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t0 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X109 GNDA.t121 VCO_FD_magic_0.div120_2_0.div24.t6 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t1 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X110 GNDA.t14 pfd_8_0.F.t6 pfd_8_0.QB.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X111 GNDA.t8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t5 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X112 pfd_8_0.before_Reset.t0 pfd_8_0.QB.t4 VDDA.t43 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X113 GNDA.t36 V_CONT.t11 VCO_FD_magic_0.vco2_3_0.V7.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X114 GNDA.t24 VDDA.t223 VCO_FD_magic_0.vco2_3_0.V5.t1 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X115 VDDA.t220 VCO_FD_magic_0.vco2_3_0.V1.t4 VCO_FD_magic_0.vco2_3_0.V2.t1 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X116 VDDA.t137 VCO_FD_magic_0.div120_2_0.div24.t7 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t0 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X117 VDDA.t15 VCO_FD_magic_0.div120_2_0.div24.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t0 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X118 GNDA.t124 a_6490_4630.t6 pfd_8_0.opamp_out.t6 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X119 VDDA.t17 opamp_cell_4_0.n_right.t6 pfd_8_0.opamp_out.t0 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X120 opamp_cell_4_0.VIN+.t2 pfd_8_0.opamp_out.t13 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X121 VDDA.t25 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t6 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t0 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X122 a_490_1400.t0 pfd_8_0.QA_b.t5 pfd_8_0.QA.t1 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X123 pfd_8_0.UP_input.t2 pfd_8_0.UP_b.t3 pfd_8_0.opamp_out.t2 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X124 V_CONT.t0 pfd_8_0.UP_input.t7 VDDA.t61 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X125 VDDA.t151 GNDA.t272 VCO_FD_magic_0.vco2_3_0.V2.t2 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X126 GNDA.t18 pfd_8_0.Reset.t2 pfd_8_0.E_b.t0 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X127 GNDA.t101 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t4 VCO_FD_magic_0.div120_2_0.div2.t0 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X128 GNDA.t32 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 VCO_FD_magic_0.div120_2_0.div24.t0 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X129 VCO_FD_magic_0.vco2_3_0.V9.t0 V_OSC.t4 VCO_FD_magic_0.vco2_3_0.V7.t0 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X130 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t3 a_6330_n1440.t3 GNDA.t269 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X131 a_2530_190.t0 a_2350_1400.t2 GNDA.t227 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X132 VDDA.t80 opamp_cell_4_0.n_left.t4 opamp_cell_4_0.n_left.t5 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X133 VCO_FD_magic_0.div120_2_0.div24.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t5 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X134 a_6320_5840.t11 V_CONT.t12 opamp_cell_4_0.n_left.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X135 a_7630_n1440.t2 VCO_FD_magic_0.div120_2_0.div2.t3 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X136 VDDA.t143 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t6 VCO_FD_magic_0.div120_2_0.div24.t2 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X137 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t7 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X138 GNDA.t119 VCO_FD_magic_0.div120_2_0.div24.t9 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t0 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X139 pfd_8_0.E.t0 pfd_8_0.E_b.t4 a_870_1400.t0 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X140 pfd_8_0.UP_b.t2 pfd_8_0.UP.t4 VDDA.t196 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X141 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t0 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X142 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN.t2 sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X143 VDDA.t34 V_OSC.t5 a_8930_n1440.t1 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X144 VDDA.t76 VCO_FD_magic_0.div120_2_0.div8.t6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t1 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X145 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t0 VCO_FD_magic_0.div120_2_0.div24.t10 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t0 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X146 a_5970_4630.t10 a_5970_4630.t8 a_5970_4630.t9 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X147 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t2 a_6330_n1440.t4 GNDA.t217 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X148 GNDA.t178 GNDA.t175 GNDA.t177 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X149 VDDA.t28 a_1870_190.t2 pfd_8_0.Reset.t0 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X150 pfd_8_0.opamp_out.t1 a_6490_4630.t7 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X151 pfd_8_0.opamp_out.t7 opamp_cell_4_0.n_right.t7 VDDA.t149 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X152 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X153 GNDA.t267 VCO_FD_magic_0.div120_2_0.div4.t3 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t1 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X154 VDDA.t86 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t3 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X155 VDDA.t41 a_7630_n1440.t5 VCO_FD_magic_0.div120_2_0.div4.t0 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X156 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t1 a_6330_n1440.t5 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t1 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X157 GNDA.t40 a_1870_190.t3 pfd_8_0.Reset.t1 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X158 V_OSC.t1 VCO_FD_magic_0.vco2_3_0.V8.t3 VCO_FD_magic_0.vco2_3_0.V2.t0 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X159 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t1 VCO_FD_magic_0.div120_2_0.div2.t4 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X160 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t0 VCO_FD_magic_0.div120_2_0.div24.t11 VDDA.t74 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X161 VDDA.t174 VDDA.t171 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X162 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t1 VCO_FD_magic_0.div120_2_0.div24.t12 GNDA.t237 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X163 opamp_cell_4_0.p_bias.t3 opamp_cell_4_0.p_bias.t2 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X164 opamp_cell_4_0.p_bias.t8 a_6220_5810.t8 GNDA.t38 sky130_fd_pr__res_xhigh_po_5p73 l=1
X165 VDDA.t145 VCO_FD_magic_0.vco2_3_0.V1.t5 VCO_FD_magic_0.vco2_3_0.V6.t1 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X166 GNDA.t221 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t4 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t1 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X167 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t8 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t0 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X168 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.t2 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X169 GNDA.t16 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t4 F_VCO.t0 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X170 GNDA.t273 V_CONT.t5 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X171 opamp_cell_4_0.n_left.t0 V_CONT.t13 a_6320_5840.t10 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X172 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t7 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t0 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X173 VDDA.t57 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t0 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X174 a_5970_4630.t0 opamp_cell_4_0.p_bias.t11 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X175 pfd_8_0.before_Reset.t1 pfd_8_0.QA.t5 a_1910_2020.t0 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X176 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t6 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X177 VDDA.t150 GNDA.t274 VCO_FD_magic_0.vco2_3_0.V6.t2 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X178 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t1 a_7630_n1440.t6 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X179 GNDA.t66 pfd_8_0.E.t4 pfd_8_0.QA.t0 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X180 VDDA.t13 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X181 a_9360_6440.t1 a_6490_4630.t2 GNDA.t154 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X182 VDDA.t170 VDDA.t168 VDDA.t170 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X183 VDDA.t106 pfd_8_0.Reset.t3 a_1390_1400.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X184 pfd_8_0.F.t0 pfd_8_0.F_b.t3 a_870_640.t0 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X185 a_2530_190.t1 a_2350_1400.t3 VDDA.t64 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X186 GNDA.t174 GNDA.t172 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X187 GNDA.t150 a_6220_5810.t2 a_6220_5810.t3 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X188 GNDA.t156 a_6490_4630.t8 pfd_8_0.opamp_out.t8 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X189 VDDA.t70 opamp_cell_4_0.n_right.t8 pfd_8_0.opamp_out.t3 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X190 VDDA.t167 VDDA.t164 VDDA.t166 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X191 GNDA.t10 a_8930_n1440.t6 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t2 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X192 GNDA.t134 pfd_8_0.F_b.t4 pfd_8_0.F.t2 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X193 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t3 VCO_FD_magic_0.div120_2_0.div24.t13 GNDA.t259 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X194 GNDA.t12 a_6220_5810.t11 a_6320_5840.t0 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X195 pfd_8_0.QB_b.t0 pfd_8_0.QB.t5 a_n30_640.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X196 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t0 a_7630_n1440.t7 GNDA.t103 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X197 GNDA.t164 a_6200_5250.t6 a_6490_4630.t4 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X198 a_5970_4630.t2 opamp_cell_4_0.VIN+.t7 a_6490_4630.t1 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X199 VDDA.t98 opamp_cell_4_0.p_bias.t12 a_5970_4630.t4 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X200 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t9 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X201 GNDA.t63 VCO_FD_magic_0.div120_2_0.div2.t5 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t1 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X202 VDDA.t5 pfd_8_0.Reset.t4 a_1390_640.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X203 VDDA.t30 opamp_cell_4_0.p_bias.t0 opamp_cell_4_0.p_bias.t1 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X204 opamp_cell_4_0.n_right.t3 a_9360_3514.t1 GNDA.t154 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X205 pfd_8_0.UP_input.t0 pfd_8_0.UP.t5 VDDA.t47 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X206 VDDA.t163 VDDA.t160 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X207 a_6320_5840.t8 a_6320_5840.t6 a_6320_5840.t7 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X208 GNDA.t97 pfd_8_0.QB.t6 pfd_8_0.QB_b.t1 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X209 a_6320_5840.t1 a_6220_5810.t12 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X210 GNDA.t54 pfd_8_0.Reset.t5 pfd_8_0.F_b.t0 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X211 a_6330_n1440.t1 VCO_FD_magic_0.div120_2_0.div4.t4 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X212 VCO_FD_magic_0.vco2_3_0.V9.t1 V_OSC.t6 VCO_FD_magic_0.vco2_3_0.V6.t0 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X213 GNDA.t231 pfd_8_0.DOWN_input.t4 V_CONT.t6 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X214 a_6320_5840.t5 a_6320_5840.t4 a_6320_5840.t5 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X215 VDDA.t159 VDDA.t157 VDDA.t159 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X216 a_6220_5810.t1 a_6220_5810.t0 GNDA.t58 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X217 GNDA.t75 V_CONT.t14 VCO_FD_magic_0.vco2_3_0.V3.t1 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X218 VDDA.t127 VCO_FD_magic_0.div120_2_0.div2.t6 a_7630_n1440.t1 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X219 pfd_8_0.E.t1 pfd_8_0.QA_b.t6 GNDA.t255 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X220 GNDA.t34 I_IN.t6 opamp_cell_4_0.VIN+.t4 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X221 GNDA.t148 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t10 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t0 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X222 a_6330_n1440.t0 VCO_FD_magic_0.div120_2_0.div4.t5 GNDA.t244 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X223 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t11 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t1 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X224 GNDA.t142 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t0 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X225 VDDA.t125 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t2 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X226 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t8 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X227 a_n30_640.t1 F_VCO.t6 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X228 GNDA.t26 VDDA.t224 VCO_FD_magic_0.vco2_3_0.V7.t2 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X229 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 GNDA.t233 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X230 a_6490_4630.t3 a_6200_5250.t7 GNDA.t162 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X231 a_6490_4630.t0 opamp_cell_4_0.VIN+.t8 a_5970_4630.t1 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X232 VDDA.t198 a_6330_n1440.t6 VCO_FD_magic_0.div120_2_0.div8.t1 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X233 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 VDDA.t115 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X234 VDDA.t103 pfd_8_0.E.t5 a_490_1400.t1 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X235 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t1 VCO_FD_magic_0.div120_2_0.div4.t6 VDDA.t208 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X236 VDDA.t213 a_2200_190.t2 a_1870_190.t1 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X237 VDDA.t32 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t0 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X238 pfd_8_0.QA_b.t1 F_REF.t1 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X239 VDDA.t218 pfd_8_0.opamp_out.t14 opamp_cell_4_0.VIN+.t1 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X240 a_490_640.t0 pfd_8_0.QB_b.t5 pfd_8_0.QB.t2 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X241 V_CONT.t4 pfd_8_0.DOWN_input.t5 GNDA.t130 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X242 pfd_8_0.QB_b.t2 F_VCO.t7 GNDA.t111 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X243 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t10 GNDA.t257 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X244 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t1 a_8930_n1440.t7 GNDA.t95 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X245 VDDA.t7 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X246 VDDA.t131 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t3 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X247 VCO_FD_magic_0.vco2_3_0.V8.t0 VCO_FD_magic_0.vco2_3_0.V9.t3 VCO_FD_magic_0.vco2_3_0.V5.t2 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X248 GNDA.t72 a_2200_190.t3 a_1870_190.t0 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X249 GNDA.t61 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t4 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t1 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X250 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t0 VCO_FD_magic_0.div120_2_0.div24.t14 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X251 opamp_cell_4_0.VIN+.t5 I_IN.t7 GNDA.t160 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X252 a_6320_5840.t2 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t1 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X253 VDDA.t216 opamp_cell_4_0.n_left.t7 opamp_cell_4_0.n_right.t4 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X254 pfd_8_0.DOWN_PFD_b.t3 pfd_8_0.QB.t7 VDDA.t209 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X255 pfd_8_0.QB.t1 pfd_8_0.QB_b.t6 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X256 GNDA.t35 V_CONT.t15 VCO_FD_magic_0.vco2_3_0.V5.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X257 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t1 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X258 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t12 GNDA.t146 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X259 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t11 GNDA.t93 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X260 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t3 GNDA.t77 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X261 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t3 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X262 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t3 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X263 GNDA.t171 GNDA.t169 GNDA.t171 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X264 pfd_8_0.E_b.t2 pfd_8_0.E.t6 GNDA.t253 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X265 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t8 GNDA.t70 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X266 VCO_FD_magic_0.vco2_3_0.V1.t1 VCO_FD_magic_0.vco2_3_0.V1.t0 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X267 opamp_cell_4_0.VIN+.t0 pfd_8_0.opamp_out.t15 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X268 pfd_8_0.DOWN_b.t0 GNDA.t275 pfd_8_0.DOWN_PFD_b.t1 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X269 GNDA.t132 a_6330_n1440.t7 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t1 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
R0 a_6200_5250.n4 a_6200_5250.n0 427.647
R1 a_6200_5250.n1 a_6200_5250.t6 321.334
R2 a_6200_5250.n5 a_6200_5250.n4 210.601
R3 a_6200_5250.n2 a_6200_5250.n1 208.868
R4 a_6200_5250.n3 a_6200_5250.t2 174.056
R5 a_6200_5250.n4 a_6200_5250.n3 152
R6 a_6200_5250.n1 a_6200_5250.t7 112.468
R7 a_6200_5250.n2 a_6200_5250.t4 112.468
R8 a_6200_5250.n3 a_6200_5250.n2 61.5894
R9 a_6200_5250.t5 a_6200_5250.n5 60.0005
R10 a_6200_5250.n5 a_6200_5250.t3 60.0005
R11 a_6200_5250.n0 a_6200_5250.t0 49.2505
R12 a_6200_5250.n0 a_6200_5250.t1 49.2505
R13 GNDA.n724 GNDA.n723 337993
R14 GNDA.n723 GNDA.n722 309276
R15 GNDA.n724 GNDA.n23 164874
R16 GNDA.n494 GNDA.n493 36300
R17 GNDA.n492 GNDA.t78 10524.4
R18 GNDA.n131 GNDA.t67 2045.88
R19 GNDA.n206 GNDA.n24 1946.93
R20 GNDA.n557 GNDA.n60 1204.13
R21 GNDA.n532 GNDA.n531 1204.13
R22 GNDA.n425 GNDA.n424 1204.13
R23 GNDA.n252 GNDA.n251 1186
R24 GNDA.n205 GNDA.n204 1186
R25 GNDA.n198 GNDA.n197 1186
R26 GNDA.n259 GNDA.n258 1186
R27 GNDA.n688 GNDA.n687 1182.8
R28 GNDA.n50 GNDA.n25 1182.8
R29 GNDA.n497 GNDA.n496 1173.78
R30 GNDA.n168 GNDA.n112 1173.78
R31 GNDA.n123 GNDA.n122 1173.78
R32 GNDA.n132 GNDA.n131 1170
R33 GNDA.n131 GNDA.n23 811.765
R34 GNDA.t141 GNDA.t116 800
R35 GNDA.n298 GNDA.t127 783.001
R36 GNDA.t222 GNDA.t106 776.471
R37 GNDA.n123 GNDA.t272 728.524
R38 GNDA.n496 GNDA.t274 728.524
R39 GNDA.n112 GNDA.t270 728.524
R40 GNDA.n126 GNDA.n120 686.717
R41 GNDA.n499 GNDA.n498 686.717
R42 GNDA.n167 GNDA.n166 686.717
R43 GNDA.n167 GNDA.n114 686.717
R44 GNDA.n498 GNDA.n111 686.717
R45 GNDA.n125 GNDA.n120 686.717
R46 GNDA.n529 GNDA.n528 669.307
R47 GNDA.n526 GNDA.n73 669.307
R48 GNDA.n463 GNDA.n462 669.307
R49 GNDA.n466 GNDA.n465 669.307
R50 GNDA.n490 GNDA.n489 669.307
R51 GNDA.n484 GNDA.n368 669.307
R52 GNDA.t220 GNDA.t114 613.048
R53 GNDA.t224 GNDA.t252 601.333
R54 GNDA.t245 GNDA.t234 601.333
R55 GNDA.n727 GNDA.n726 585.003
R56 GNDA.n297 GNDA.n296 585.003
R57 GNDA.n294 GNDA.n293 585.001
R58 GNDA.n292 GNDA.n278 585.001
R59 GNDA.n291 GNDA.n275 585.001
R60 GNDA.n272 GNDA.n271 585.001
R61 GNDA.n250 GNDA.n249 585.001
R62 GNDA.n207 GNDA.n206 585.001
R63 GNDA.n367 GNDA.n366 585.001
R64 GNDA.n269 GNDA.n263 585.001
R65 GNDA.n270 GNDA.n266 585.001
R66 GNDA.n721 GNDA.n720 585.001
R67 GNDA.n36 GNDA.n31 585.001
R68 GNDA.n690 GNDA.n689 585.001
R69 GNDA.n732 GNDA.n731 585.001
R70 GNDA.n730 GNDA.n19 585.001
R71 GNDA.n729 GNDA.n16 585.001
R72 GNDA.n728 GNDA.n13 585.001
R73 GNDA.n725 GNDA.n2 585.001
R74 GNDA.n488 GNDA.n426 585
R75 GNDA.n486 GNDA.n485 585
R76 GNDA.n441 GNDA.n437 585
R77 GNDA.n439 GNDA.n436 585
R78 GNDA.n77 GNDA.n74 585
R79 GNDA.n80 GNDA.n79 585
R80 GNDA.n99 GNDA.n98 585
R81 GNDA.n100 GNDA.n99 585
R82 GNDA.n97 GNDA.n95 585
R83 GNDA.n93 GNDA.n91 585
R84 GNDA.n102 GNDA.n101 585
R85 GNDA.n101 GNDA.n100 585
R86 GNDA.n703 GNDA.t275 566.966
R87 GNDA.n100 GNDA.t45 522.179
R88 GNDA.t39 GNDA.t2 517.648
R89 GNDA.t31 GNDA.n36 482.353
R90 GNDA.t15 GNDA.n724 482.353
R91 GNDA.t81 GNDA.n730 458.825
R92 GNDA.t78 GNDA.t90 425.334
R93 GNDA.t226 GNDA.n270 418
R94 GNDA.n689 GNDA.t69 388.236
R95 GNDA.t198 GNDA.t129 376.654
R96 GNDA.t52 GNDA.t96 376.471
R97 GNDA.t190 GNDA.n530 359.534
R98 GNDA.n367 GNDA.t76 344.668
R99 GNDA.t228 GNDA.n269 344.668
R100 GNDA.n75 GNDA.t208 336.329
R101 GNDA.n75 GNDA.t189 336.329
R102 GNDA.n438 GNDA.t169 336.329
R103 GNDA.n438 GNDA.t197 336.329
R104 GNDA.t79 GNDA.t29 329.413
R105 GNDA.n103 GNDA.t185 320.7
R106 GNDA.n483 GNDA.t172 320.7
R107 GNDA.n688 GNDA.t73 317.647
R108 GNDA.t264 GNDA.t173 316.733
R109 GNDA.t33 GNDA.t243 316.733
R110 GNDA.t152 GNDA.t125 316.733
R111 GNDA.n531 GNDA.t170 308.171
R112 GNDA.t135 GNDA.n60 308.171
R113 GNDA.t60 GNDA.t39 305.882
R114 GNDA.n169 GNDA.t179 304.634
R115 GNDA.n253 GNDA.t201 304.634
R116 GNDA.n203 GNDA.t175 304.634
R117 GNDA.n199 GNDA.t182 304.634
R118 GNDA.n634 GNDA.t30 295.933
R119 GNDA.n606 GNDA.t142 295.933
R120 GNDA.n42 GNDA.t32 295.933
R121 GNDA.n248 GNDA.t205 292.584
R122 GNDA.n208 GNDA.t193 292.584
R123 GNDA.n491 GNDA.n425 291.051
R124 GNDA.t86 GNDA.n291 286
R125 GNDA.t68 GNDA.n25 270.589
R126 GNDA.n126 GNDA.t75 260
R127 GNDA.t75 GNDA.n125 260
R128 GNDA.t249 GNDA.t137 258.825
R129 GNDA.n721 GNDA.n25 258.825
R130 GNDA.t7 GNDA.t145 258.825
R131 GNDA.t84 GNDA.t108 258.825
R132 GNDA.t104 GNDA.t143 258.825
R133 GNDA.t13 GNDA.t79 258.825
R134 GNDA.t29 GNDA.t52 258.825
R135 GNDA.t92 GNDA.t15 258.825
R136 GNDA.n639 GNDA.n636 256.207
R137 GNDA.n491 GNDA.n490 250.349
R138 GNDA.n491 GNDA.n368 250.349
R139 GNDA.n464 GNDA.n463 250.349
R140 GNDA.n465 GNDA.n464 250.349
R141 GNDA.n530 GNDA.n529 250.349
R142 GNDA.n530 GNDA.n73 250.349
R143 GNDA.n100 GNDA.n94 250.349
R144 GNDA.n638 GNDA.n637 247.934
R145 GNDA.n630 GNDA.n629 247.934
R146 GNDA.n655 GNDA.n628 247.934
R147 GNDA.n662 GNDA.n625 247.934
R148 GNDA.n674 GNDA.n620 247.934
R149 GNDA.n618 GNDA.n617 247.934
R150 GNDA.n45 GNDA.n44 247.934
R151 GNDA.n594 GNDA.n47 247.934
R152 GNDA.n575 GNDA.n574 247.934
R153 GNDA.n572 GNDA.n55 247.934
R154 GNDA.t236 GNDA.n729 247.06
R155 GNDA.n560 GNDA.n559 246.714
R156 GNDA.n258 GNDA.t181 245
R157 GNDA.n252 GNDA.t204 245
R158 GNDA.n204 GNDA.t178 245
R159 GNDA.n198 GNDA.t184 245
R160 GNDA.n168 GNDA.n167 241.643
R161 GNDA.n498 GNDA.n497 241.643
R162 GNDA.n122 GNDA.n120 241.643
R163 GNDA.t42 GNDA.t7 235.294
R164 GNDA.n689 GNDA.n688 235.294
R165 GNDA.n124 GNDA.t117 233
R166 GNDA.n687 GNDA.t74 233
R167 GNDA.n50 GNDA.t138 233
R168 GNDA.n495 GNDA.t26 233
R169 GNDA.n113 GNDA.t24 233
R170 GNDA.t90 GNDA.n367 227.333
R171 GNDA.n269 GNDA.t76 227.333
R172 GNDA.n270 GNDA.t228 227.333
R173 GNDA.n551 GNDA.n63 219.133
R174 GNDA.n65 GNDA.n64 219.133
R175 GNDA.n539 GNDA.n69 219.133
R176 GNDA.n404 GNDA.n403 219.133
R177 GNDA.n410 GNDA.n401 219.133
R178 GNDA.n418 GNDA.n398 219.133
R179 GNDA.n392 GNDA.n372 219.133
R180 GNDA.n386 GNDA.n385 219.133
R181 GNDA.n378 GNDA.n377 219.133
R182 GNDA.t5 GNDA.n23 216.788
R183 GNDA.t71 GNDA.t236 211.766
R184 GNDA.t240 GNDA.t13 211.766
R185 GNDA.t96 GNDA.t256 211.766
R186 GNDA.t110 GNDA.t214 211.766
R187 GNDA.n294 GNDA.n292 205.333
R188 GNDA.n255 GNDA.n171 204.201
R189 GNDA.n201 GNDA.n195 204.201
R190 GNDA.n202 GNDA.n194 204.201
R191 GNDA.n200 GNDA.n196 204.201
R192 GNDA.n254 GNDA.n172 204.201
R193 GNDA.n257 GNDA.n256 204.201
R194 GNDA.n731 GNDA.t64 200
R195 GNDA.n3 GNDA.t97 198.058
R196 GNDA.n773 GNDA.t80 198.058
R197 GNDA.n761 GNDA.t134 198.058
R198 GNDA.n11 GNDA.t263 198.058
R199 GNDA.n323 GNDA.t253 198.058
R200 GNDA.n318 GNDA.t225 198.058
R201 GNDA.n288 GNDA.t235 198.058
R202 GNDA.n304 GNDA.t246 198.058
R203 GNDA.n271 GNDA.t226 198
R204 GNDA.n291 GNDA.t238 198
R205 GNDA.n292 GNDA.t47 198
R206 GNDA.t17 GNDA.n294 198
R207 GNDA.n297 GNDA.t254 198
R208 GNDA.t65 GNDA.n297 198
R209 GNDA.n79 GNDA.n74 197
R210 GNDA.n437 GNDA.n436 197
R211 GNDA.n485 GNDA.n426 197
R212 GNDA.n99 GNDA.n95 197
R213 GNDA.n101 GNDA.n93 197
R214 GNDA.t83 GNDA.t266 188.327
R215 GNDA.t19 GNDA.t112 188.327
R216 GNDA.t102 GNDA.t49 188.327
R217 GNDA.t98 GNDA.t87 188.327
R218 GNDA.t268 GNDA.t131 188.327
R219 GNDA.t216 GNDA.t55 188.327
R220 GNDA.t115 GNDA.t118 188.327
R221 GNDA.t147 GNDA.t211 188.327
R222 GNDA.t211 GNDA.t220 188.327
R223 GNDA.t114 GNDA.t0 188.236
R224 GNDA.t145 GNDA.t68 188.236
R225 GNDA.n528 GNDA.n527 185
R226 GNDA.n527 GNDA.n526 185
R227 GNDA.n462 GNDA.n435 185
R228 GNDA.n466 GNDA.n435 185
R229 GNDA.n489 GNDA.n427 185
R230 GNDA.n484 GNDA.n427 185
R231 GNDA.n98 GNDA.n92 185
R232 GNDA.n102 GNDA.n92 185
R233 GNDA.n528 GNDA.n75 166.63
R234 GNDA.n462 GNDA.n438 166.63
R235 GNDA.t44 GNDA.t53 164.707
R236 GNDA.t232 GNDA.t262 164.707
R237 GNDA.t133 GNDA.t120 164.707
R238 GNDA.t3 GNDA.t258 164.707
R239 GNDA.t209 GNDA.t216 162.647
R240 GNDA.t47 GNDA.t86 161.333
R241 GNDA.t252 GNDA.t17 161.333
R242 GNDA.t254 GNDA.t224 161.333
R243 GNDA.t234 GNDA.t65 161.333
R244 GNDA.t127 GNDA.t245 161.333
R245 GNDA.n728 GNDA.t44 152.941
R246 GNDA.t258 GNDA.n727 152.941
R247 GNDA.n725 GNDA.t92 152.941
R248 GNDA.n168 GNDA.t59 149.344
R249 GNDA.n497 GNDA.t23 149.344
R250 GNDA.t25 GNDA.t139 147.738
R251 GNDA.n464 GNDA.t102 145.525
R252 GNDA.n530 GNDA.t268 145.525
R253 GNDA.n722 GNDA.t45 145.525
R254 GNDA.n133 GNDA.n132 142.694
R255 GNDA.n723 GNDA.t238 139.333
R256 GNDA.n249 GNDA.t207 134.501
R257 GNDA.n207 GNDA.t196 134.501
R258 GNDA.n7 GNDA.t14 130.713
R259 GNDA.n2 GNDA.t111 130.001
R260 GNDA.n13 GNDA.t54 130.001
R261 GNDA.n16 GNDA.t40 130.001
R262 GNDA.n19 GNDA.t72 130.001
R263 GNDA.n732 GNDA.t82 130.001
R264 GNDA.n298 GNDA.t128 130.001
R265 GNDA.n293 GNDA.t18 130.001
R266 GNDA.n278 GNDA.t48 130.001
R267 GNDA.n275 GNDA.t239 130.001
R268 GNDA.n272 GNDA.t227 130.001
R269 GNDA.n8 GNDA.t4 130.001
R270 GNDA.n295 GNDA.t255 130.001
R271 GNDA.n287 GNDA.t66 130.001
R272 GNDA.n121 GNDA.t6 128.562
R273 GNDA.t266 GNDA.t230 128.405
R274 GNDA.t112 GNDA.t198 128.405
R275 GNDA.t159 GNDA.t98 128.405
R276 GNDA.t118 GNDA.t186 128.405
R277 GNDA.n165 GNDA.t35 127.754
R278 GNDA.n110 GNDA.t36 127.754
R279 GNDA.n690 GNDA.t70 122.501
R280 GNDA.n31 GNDA.t43 122.501
R281 GNDA.n720 GNDA.t1 122.501
R282 GNDA.n266 GNDA.t229 122.501
R283 GNDA.n263 GNDA.t77 122.501
R284 GNDA.n366 GNDA.t91 122.501
R285 GNDA.t69 GNDA.t141 117.647
R286 GNDA.t64 GNDA.t81 117.647
R287 GNDA.n250 GNDA.t37 112.451
R288 GNDA.n492 GNDA.t100 111.284
R289 GNDA.n36 GNDA.t84 105.882
R290 GNDA.t2 GNDA.n728 105.882
R291 GNDA.n727 GNDA.t240 105.882
R292 GNDA.t214 GNDA.n725 105.882
R293 GNDA.t247 GNDA.t9 100.001
R294 GNDA.t9 GNDA.t94 100.001
R295 GNDA.n176 GNDA.n175 97.8707
R296 GNDA.n180 GNDA.n179 97.8707
R297 GNDA.n184 GNDA.n183 97.8707
R298 GNDA.n188 GNDA.n187 97.8707
R299 GNDA.n193 GNDA.n192 97.8707
R300 GNDA.n197 GNDA.t250 97.7783
R301 GNDA.n251 GNDA.t202 95.1512
R302 GNDA.n259 GNDA.t180 94.9025
R303 GNDA.t53 GNDA.t232 94.1181
R304 GNDA.t262 GNDA.t222 94.1181
R305 GNDA.t106 GNDA.t133 94.1181
R306 GNDA.t120 GNDA.t3 94.1181
R307 GNDA.n473 GNDA.n472 92.2612
R308 GNDA.n481 GNDA.n480 92.2612
R309 GNDA.n459 GNDA.n458 92.2612
R310 GNDA.n452 GNDA.n447 92.2612
R311 GNDA.n520 GNDA.n87 92.2612
R312 GNDA.n514 GNDA.n90 92.2612
R313 GNDA.n527 GNDA.n78 91.3721
R314 GNDA.n86 GNDA.n76 91.3721
R315 GNDA.n86 GNDA.n81 91.3721
R316 GNDA.n440 GNDA.n435 91.3721
R317 GNDA.n461 GNDA.n460 91.3721
R318 GNDA.n460 GNDA.n434 91.3721
R319 GNDA.n487 GNDA.n427 90.7567
R320 GNDA.n96 GNDA.n92 90.7567
R321 GNDA.t250 GNDA.t242 89.1508
R322 GNDA.n205 GNDA.t194 86.275
R323 GNDA.n132 GNDA.t273 86.0829
R324 GNDA.n490 GNDA.n426 84.306
R325 GNDA.n485 GNDA.n368 84.306
R326 GNDA.n463 GNDA.n437 84.306
R327 GNDA.n465 GNDA.n436 84.306
R328 GNDA.n529 GNDA.n74 84.306
R329 GNDA.n79 GNDA.n73 84.306
R330 GNDA.n95 GNDA.n94 84.306
R331 GNDA.n94 GNDA.n93 84.306
R332 GNDA.n201 GNDA.n200 83.2005
R333 GNDA.n202 GNDA.n201 83.2005
R334 GNDA.n132 GNDA.t271 82.8829
R335 GNDA.n723 GNDA.n24 80.6672
R336 GNDA.t260 GNDA.t183 77.6476
R337 GNDA.n251 GNDA.n250 74.9677
R338 GNDA.t202 GNDA.t157 74.8697
R339 GNDA.t123 GNDA.t180 74.7717
R340 GNDA.t21 GNDA.t123 74.7717
R341 GNDA.t155 GNDA.t21 74.7717
R342 GNDA.t157 GNDA.t155 74.7717
R343 GNDA.t51 GNDA.t41 74.7717
R344 GNDA.t163 GNDA.t161 74.7717
R345 GNDA.t165 GNDA.t176 74.7717
R346 GNDA.t122 GNDA.t206 72.0844
R347 GNDA.t218 GNDA.t167 71.8959
R348 GNDA.t0 GNDA.t249 70.5887
R349 GNDA.t173 GNDA.n425 68.483
R350 GNDA.n531 GNDA.t33 68.483
R351 GNDA.t125 GNDA.n60 68.483
R352 GNDA.n256 GNDA.n255 66.5605
R353 GNDA.n255 GNDA.n254 66.5605
R354 GNDA.t151 GNDA.t88 66.1443
R355 GNDA.n271 GNDA.n24 66.0005
R356 GNDA.n255 GNDA.n170 65.9634
R357 GNDA.n733 GNDA.n732 60.29
R358 GNDA.n740 GNDA.n19 60.29
R359 GNDA.n746 GNDA.n16 60.29
R360 GNDA.n753 GNDA.n13 60.29
R361 GNDA.n781 GNDA.n2 60.29
R362 GNDA.n299 GNDA.n298 60.29
R363 GNDA.n293 GNDA.n281 60.29
R364 GNDA.n331 GNDA.n278 60.29
R365 GNDA.n338 GNDA.n275 60.29
R366 GNDA.n344 GNDA.n272 60.29
R367 GNDA.n171 GNDA.t22 60.0005
R368 GNDA.n171 GNDA.t156 60.0005
R369 GNDA.n195 GNDA.t162 60.0005
R370 GNDA.n195 GNDA.t168 60.0005
R371 GNDA.n194 GNDA.t166 60.0005
R372 GNDA.n194 GNDA.t177 60.0005
R373 GNDA.t184 GNDA.n196 60.0005
R374 GNDA.n196 GNDA.t164 60.0005
R375 GNDA.n172 GNDA.t158 60.0005
R376 GNDA.n172 GNDA.t203 60.0005
R377 GNDA.t181 GNDA.n257 60.0005
R378 GNDA.n257 GNDA.t124 60.0005
R379 GNDA.t230 GNDA.t264 59.9227
R380 GNDA.t129 GNDA.t83 59.9227
R381 GNDA.t243 GNDA.t159 59.9227
R382 GNDA.t87 GNDA.t190 59.9227
R383 GNDA.t186 GNDA.t152 59.9227
R384 GNDA.n352 GNDA.n266 59.5478
R385 GNDA.n359 GNDA.n263 59.5478
R386 GNDA.n366 GNDA.n365 59.5478
R387 GNDA.n493 GNDA.t247 59.0914
R388 GNDA.n708 GNDA.n31 58.9809
R389 GNDA.n691 GNDA.n690 58.9809
R390 GNDA.n720 GNDA.n719 58.9809
R391 GNDA.t137 GNDA.n721 58.824
R392 GNDA.n731 GNDA.t73 58.824
R393 GNDA.n766 GNDA.n8 54.4005
R394 GNDA.n768 GNDA.n7 54.4005
R395 GNDA.n687 GNDA.n686 54.4005
R396 GNDA.n588 GNDA.n50 54.4005
R397 GNDA.n312 GNDA.n287 54.4005
R398 GNDA.n295 GNDA.n286 54.4005
R399 GNDA.n493 GNDA.n259 51.7652
R400 GNDA.t149 GNDA.t151 48.8894
R401 GNDA.n636 GNDA.t93 48.0005
R402 GNDA.n636 GNDA.t16 48.0005
R403 GNDA.n637 GNDA.t257 48.0005
R404 GNDA.n637 GNDA.t215 48.0005
R405 GNDA.n629 GNDA.t259 48.0005
R406 GNDA.n629 GNDA.t241 48.0005
R407 GNDA.n628 GNDA.t107 48.0005
R408 GNDA.n628 GNDA.t121 48.0005
R409 GNDA.n625 GNDA.t233 48.0005
R410 GNDA.n625 GNDA.t223 48.0005
R411 GNDA.n620 GNDA.t237 48.0005
R412 GNDA.n620 GNDA.t61 48.0005
R413 GNDA.n617 GNDA.t105 48.0005
R414 GNDA.n617 GNDA.t144 48.0005
R415 GNDA.n44 GNDA.t109 48.0005
R416 GNDA.n44 GNDA.t85 48.0005
R417 GNDA.n47 GNDA.t146 48.0005
R418 GNDA.n47 GNDA.t8 48.0005
R419 GNDA.n574 GNDA.t212 48.0005
R420 GNDA.n574 GNDA.t221 48.0005
R421 GNDA.n55 GNDA.t46 48.0005
R422 GNDA.n55 GNDA.t148 48.0005
R423 GNDA.n559 GNDA.t153 48.0005
R424 GNDA.n559 GNDA.t119 48.0005
R425 GNDA.n63 GNDA.t217 48.0005
R426 GNDA.n63 GNDA.t56 48.0005
R427 GNDA.n64 GNDA.t269 48.0005
R428 GNDA.n64 GNDA.t132 48.0005
R429 GNDA.n69 GNDA.t244 48.0005
R430 GNDA.n69 GNDA.t99 48.0005
R431 GNDA.n403 GNDA.t103 48.0005
R432 GNDA.n403 GNDA.t50 48.0005
R433 GNDA.n401 GNDA.t113 48.0005
R434 GNDA.n401 GNDA.t20 48.0005
R435 GNDA.n398 GNDA.t265 48.0005
R436 GNDA.n398 GNDA.t267 48.0005
R437 GNDA.n372 GNDA.t95 48.0005
R438 GNDA.n372 GNDA.t101 48.0005
R439 GNDA.n385 GNDA.t248 48.0005
R440 GNDA.n385 GNDA.t10 48.0005
R441 GNDA.n377 GNDA.t140 48.0005
R442 GNDA.n377 GNDA.t63 48.0005
R443 GNDA.t116 GNDA.t31 47.0593
R444 GNDA.t143 GNDA.t71 47.0593
R445 GNDA.t256 GNDA.t110 47.0593
R446 GNDA.t213 GNDA.t154 44.964
R447 GNDA.n122 GNDA.t5 43.3582
R448 GNDA.n122 GNDA.t59 43.3582
R449 GNDA.t23 GNDA.n168 43.3582
R450 GNDA.n497 GNDA.t25 43.3582
R451 GNDA.t167 GNDA.t27 43.1378
R452 GNDA.t100 GNDA.n491 42.8021
R453 GNDA.n464 GNDA.t19 42.8021
R454 GNDA.n100 GNDA.t115 42.8021
R455 GNDA.n722 GNDA.t147 42.8021
R456 GNDA.n201 GNDA.n190 41.6005
R457 GNDA.n509 GNDA.n508 41.3005
R458 GNDA.t94 GNDA.n492 40.9096
R459 GNDA.t11 GNDA.t122 40.3637
R460 GNDA.t154 GNDA.n493 40.1465
R461 GNDA.n134 GNDA.n133 39.4989
R462 GNDA.n245 GNDA.n170 39.4985
R463 GNDA.t183 GNDA.t57 37.3861
R464 GNDA.t57 GNDA.t163 37.3861
R465 GNDA.n495 GNDA.n111 35.6576
R466 GNDA.n500 GNDA.n499 35.6576
R467 GNDA.n166 GNDA.n164 35.6576
R468 GNDA.n114 GNDA.n113 35.6576
R469 GNDA.t62 GNDA.t213 35.329
R470 GNDA.n125 GNDA.n124 34.3278
R471 GNDA.n146 GNDA.n126 34.3278
R472 GNDA.n782 GNDA.n781 33.0991
R473 GNDA.n299 GNDA.n0 33.0991
R474 GNDA.n473 GNDA.n471 32.0005
R475 GNDA.n471 GNDA.n431 32.0005
R476 GNDA.n479 GNDA.n478 32.0005
R477 GNDA.n478 GNDA.n429 32.0005
R478 GNDA.n474 GNDA.n429 32.0005
R479 GNDA.n442 GNDA.n433 32.0005
R480 GNDA.n457 GNDA.n445 32.0005
R481 GNDA.n453 GNDA.n445 32.0005
R482 GNDA.n453 GNDA.n452 32.0005
R483 GNDA.n451 GNDA.n448 32.0005
R484 GNDA.n448 GNDA.n82 32.0005
R485 GNDA.n525 GNDA.n83 32.0005
R486 GNDA.n521 GNDA.n83 32.0005
R487 GNDA.n519 GNDA.n88 32.0005
R488 GNDA.n515 GNDA.n88 32.0005
R489 GNDA.n513 GNDA.n104 32.0005
R490 GNDA.n718 GNDA.n27 32.0005
R491 GNDA.n714 GNDA.n27 32.0005
R492 GNDA.n714 GNDA.n713 32.0005
R493 GNDA.n713 GNDA.n712 32.0005
R494 GNDA.n712 GNDA.n29 32.0005
R495 GNDA.n708 GNDA.n29 32.0005
R496 GNDA.n708 GNDA.n707 32.0005
R497 GNDA.n707 GNDA.n706 32.0005
R498 GNDA.n706 GNDA.n32 32.0005
R499 GNDA.n701 GNDA.n32 32.0005
R500 GNDA.n701 GNDA.n700 32.0005
R501 GNDA.n700 GNDA.n699 32.0005
R502 GNDA.n699 GNDA.n34 32.0005
R503 GNDA.n695 GNDA.n694 32.0005
R504 GNDA.n694 GNDA.n693 32.0005
R505 GNDA.n693 GNDA.n22 32.0005
R506 GNDA.n734 GNDA.n22 32.0005
R507 GNDA.n738 GNDA.n20 32.0005
R508 GNDA.n739 GNDA.n738 32.0005
R509 GNDA.n741 GNDA.n17 32.0005
R510 GNDA.n745 GNDA.n17 32.0005
R511 GNDA.n748 GNDA.n747 32.0005
R512 GNDA.n748 GNDA.n14 32.0005
R513 GNDA.n752 GNDA.n14 32.0005
R514 GNDA.n755 GNDA.n754 32.0005
R515 GNDA.n755 GNDA.n11 32.0005
R516 GNDA.n759 GNDA.n11 32.0005
R517 GNDA.n760 GNDA.n759 32.0005
R518 GNDA.n761 GNDA.n760 32.0005
R519 GNDA.n761 GNDA.n9 32.0005
R520 GNDA.n765 GNDA.n9 32.0005
R521 GNDA.n769 GNDA.n5 32.0005
R522 GNDA.n773 GNDA.n5 32.0005
R523 GNDA.n774 GNDA.n773 32.0005
R524 GNDA.n775 GNDA.n774 32.0005
R525 GNDA.n775 GNDA.n3 32.0005
R526 GNDA.n779 GNDA.n3 32.0005
R527 GNDA.n780 GNDA.n779 32.0005
R528 GNDA.n147 GNDA.n118 32.0005
R529 GNDA.n151 GNDA.n118 32.0005
R530 GNDA.n152 GNDA.n151 32.0005
R531 GNDA.n153 GNDA.n152 32.0005
R532 GNDA.n153 GNDA.n115 32.0005
R533 GNDA.n379 GNDA.n375 32.0005
R534 GNDA.n383 GNDA.n375 32.0005
R535 GNDA.n384 GNDA.n383 32.0005
R536 GNDA.n387 GNDA.n384 32.0005
R537 GNDA.n391 GNDA.n373 32.0005
R538 GNDA.n394 GNDA.n393 32.0005
R539 GNDA.n394 GNDA.n369 32.0005
R540 GNDA.n423 GNDA.n370 32.0005
R541 GNDA.n419 GNDA.n370 32.0005
R542 GNDA.n417 GNDA.n416 32.0005
R543 GNDA.n416 GNDA.n399 32.0005
R544 GNDA.n412 GNDA.n399 32.0005
R545 GNDA.n412 GNDA.n411 32.0005
R546 GNDA.n409 GNDA.n402 32.0005
R547 GNDA.n405 GNDA.n72 32.0005
R548 GNDA.n533 GNDA.n72 32.0005
R549 GNDA.n537 GNDA.n70 32.0005
R550 GNDA.n538 GNDA.n537 32.0005
R551 GNDA.n540 GNDA.n67 32.0005
R552 GNDA.n544 GNDA.n67 32.0005
R553 GNDA.n545 GNDA.n544 32.0005
R554 GNDA.n546 GNDA.n545 32.0005
R555 GNDA.n550 GNDA.n549 32.0005
R556 GNDA.n552 GNDA.n61 32.0005
R557 GNDA.n556 GNDA.n61 32.0005
R558 GNDA.n561 GNDA.n558 32.0005
R559 GNDA.n565 GNDA.n58 32.0005
R560 GNDA.n566 GNDA.n565 32.0005
R561 GNDA.n567 GNDA.n566 32.0005
R562 GNDA.n567 GNDA.n56 32.0005
R563 GNDA.n571 GNDA.n56 32.0005
R564 GNDA.n576 GNDA.n573 32.0005
R565 GNDA.n580 GNDA.n53 32.0005
R566 GNDA.n581 GNDA.n580 32.0005
R567 GNDA.n582 GNDA.n581 32.0005
R568 GNDA.n582 GNDA.n51 32.0005
R569 GNDA.n586 GNDA.n51 32.0005
R570 GNDA.n587 GNDA.n586 32.0005
R571 GNDA.n589 GNDA.n48 32.0005
R572 GNDA.n593 GNDA.n48 32.0005
R573 GNDA.n596 GNDA.n595 32.0005
R574 GNDA.n600 GNDA.n599 32.0005
R575 GNDA.n601 GNDA.n600 32.0005
R576 GNDA.n605 GNDA.n604 32.0005
R577 GNDA.n607 GNDA.n605 32.0005
R578 GNDA.n611 GNDA.n40 32.0005
R579 GNDA.n612 GNDA.n611 32.0005
R580 GNDA.n613 GNDA.n612 32.0005
R581 GNDA.n613 GNDA.n37 32.0005
R582 GNDA.n685 GNDA.n38 32.0005
R583 GNDA.n681 GNDA.n38 32.0005
R584 GNDA.n681 GNDA.n680 32.0005
R585 GNDA.n680 GNDA.n679 32.0005
R586 GNDA.n676 GNDA.n675 32.0005
R587 GNDA.n673 GNDA.n621 32.0005
R588 GNDA.n669 GNDA.n621 32.0005
R589 GNDA.n669 GNDA.n668 32.0005
R590 GNDA.n668 GNDA.n667 32.0005
R591 GNDA.n667 GNDA.n623 32.0005
R592 GNDA.n663 GNDA.n623 32.0005
R593 GNDA.n661 GNDA.n660 32.0005
R594 GNDA.n660 GNDA.n626 32.0005
R595 GNDA.n656 GNDA.n626 32.0005
R596 GNDA.n654 GNDA.n653 32.0005
R597 GNDA.n650 GNDA.n649 32.0005
R598 GNDA.n649 GNDA.n648 32.0005
R599 GNDA.n648 GNDA.n632 32.0005
R600 GNDA.n644 GNDA.n643 32.0005
R601 GNDA.n643 GNDA.n642 32.0005
R602 GNDA.n642 GNDA.n635 32.0005
R603 GNDA.n164 GNDA.n116 32.0005
R604 GNDA.n160 GNDA.n116 32.0005
R605 GNDA.n160 GNDA.n159 32.0005
R606 GNDA.n159 GNDA.n158 32.0005
R607 GNDA.n158 GNDA.n109 32.0005
R608 GNDA.n500 GNDA.n107 32.0005
R609 GNDA.n504 GNDA.n107 32.0005
R610 GNDA.n365 GNDA.n364 32.0005
R611 GNDA.n364 GNDA.n261 32.0005
R612 GNDA.n360 GNDA.n261 32.0005
R613 GNDA.n358 GNDA.n357 32.0005
R614 GNDA.n357 GNDA.n264 32.0005
R615 GNDA.n353 GNDA.n264 32.0005
R616 GNDA.n351 GNDA.n350 32.0005
R617 GNDA.n350 GNDA.n267 32.0005
R618 GNDA.n346 GNDA.n267 32.0005
R619 GNDA.n346 GNDA.n345 32.0005
R620 GNDA.n343 GNDA.n273 32.0005
R621 GNDA.n339 GNDA.n273 32.0005
R622 GNDA.n337 GNDA.n336 32.0005
R623 GNDA.n336 GNDA.n276 32.0005
R624 GNDA.n332 GNDA.n276 32.0005
R625 GNDA.n330 GNDA.n329 32.0005
R626 GNDA.n329 GNDA.n279 32.0005
R627 GNDA.n325 GNDA.n324 32.0005
R628 GNDA.n324 GNDA.n323 32.0005
R629 GNDA.n323 GNDA.n282 32.0005
R630 GNDA.n319 GNDA.n282 32.0005
R631 GNDA.n319 GNDA.n318 32.0005
R632 GNDA.n318 GNDA.n317 32.0005
R633 GNDA.n317 GNDA.n284 32.0005
R634 GNDA.n311 GNDA.n310 32.0005
R635 GNDA.n310 GNDA.n288 32.0005
R636 GNDA.n306 GNDA.n288 32.0005
R637 GNDA.n306 GNDA.n305 32.0005
R638 GNDA.n305 GNDA.n304 32.0005
R639 GNDA.n304 GNDA.n290 32.0005
R640 GNDA.n300 GNDA.n290 32.0005
R641 GNDA.n245 GNDA.n244 32.0005
R642 GNDA.n244 GNDA.n243 32.0005
R643 GNDA.n243 GNDA.n174 32.0005
R644 GNDA.n239 GNDA.n174 32.0005
R645 GNDA.n239 GNDA.n238 32.0005
R646 GNDA.n238 GNDA.n237 32.0005
R647 GNDA.n237 GNDA.n178 32.0005
R648 GNDA.n233 GNDA.n178 32.0005
R649 GNDA.n233 GNDA.n232 32.0005
R650 GNDA.n232 GNDA.n231 32.0005
R651 GNDA.n231 GNDA.n182 32.0005
R652 GNDA.n227 GNDA.n182 32.0005
R653 GNDA.n227 GNDA.n226 32.0005
R654 GNDA.n226 GNDA.n225 32.0005
R655 GNDA.n225 GNDA.n186 32.0005
R656 GNDA.n221 GNDA.n220 32.0005
R657 GNDA.n220 GNDA.n219 32.0005
R658 GNDA.n219 GNDA.n191 32.0005
R659 GNDA.n214 GNDA.n191 32.0005
R660 GNDA.n214 GNDA.n213 32.0005
R661 GNDA.n213 GNDA.n212 32.0005
R662 GNDA.n135 GNDA.n134 32.0005
R663 GNDA.n135 GNDA.n129 32.0005
R664 GNDA.n139 GNDA.n129 32.0005
R665 GNDA.n140 GNDA.n139 32.0005
R666 GNDA.n141 GNDA.n140 32.0005
R667 GNDA.n141 GNDA.n127 32.0005
R668 GNDA.n145 GNDA.n127 32.0005
R669 GNDA.t41 GNDA.t11 31.6345
R670 GNDA.n505 GNDA.n504 29.4625
R671 GNDA.n526 GNDA.n525 29.0291
R672 GNDA.n467 GNDA.n466 29.0291
R673 GNDA.n379 GNDA.n378 28.8005
R674 GNDA.n418 GNDA.n417 28.8005
R675 GNDA.n540 GNDA.n539 28.8005
R676 GNDA.n561 GNDA.n560 28.8005
R677 GNDA.n596 GNDA.n45 28.8005
R678 GNDA.n607 GNDA.n606 28.8005
R679 GNDA.n638 GNDA.n635 28.8005
R680 GNDA.n360 GNDA.n359 28.8005
R681 GNDA.n344 GNDA.n343 28.8005
R682 GNDA.n206 GNDA.n205 28.7587
R683 GNDA.n253 GNDA.n252 27.2005
R684 GNDA.n258 GNDA.n169 27.2005
R685 GNDA.t242 GNDA.t149 25.8829
R686 GNDA.t139 GNDA.n494 25.6939
R687 GNDA.t49 GNDA.t170 25.6814
R688 GNDA.t131 GNDA.t209 25.6814
R689 GNDA.t55 GNDA.t135 25.6814
R690 GNDA.n467 GNDA.n433 25.6005
R691 GNDA.n520 GNDA.n519 25.6005
R692 GNDA.n515 GNDA.n514 25.6005
R693 GNDA.n719 GNDA.n718 25.6005
R694 GNDA.n691 GNDA.n34 25.6005
R695 GNDA.n733 GNDA.n20 25.6005
R696 GNDA.n746 GNDA.n745 25.6005
R697 GNDA.n753 GNDA.n752 25.6005
R698 GNDA.n767 GNDA.n766 25.6005
R699 GNDA.n147 GNDA.n146 25.6005
R700 GNDA.n392 GNDA.n391 25.6005
R701 GNDA.n404 GNDA.n402 25.6005
R702 GNDA.n551 GNDA.n550 25.6005
R703 GNDA.n576 GNDA.n575 25.6005
R704 GNDA.n676 GNDA.n618 25.6005
R705 GNDA.n662 GNDA.n661 25.6005
R706 GNDA.n653 GNDA.n630 25.6005
R707 GNDA.n644 GNDA.n634 25.6005
R708 GNDA.n353 GNDA.n352 25.6005
R709 GNDA.n332 GNDA.n331 25.6005
R710 GNDA.n281 GNDA.n279 25.6005
R711 GNDA.n313 GNDA.n286 25.6005
R712 GNDA.n313 GNDA.n312 25.6005
R713 GNDA.n204 GNDA.n203 25.6005
R714 GNDA.n199 GNDA.n198 25.6005
R715 GNDA.n221 GNDA.n190 25.6005
R716 GNDA.n212 GNDA 25.6005
R717 GNDA.n249 GNDA.n248 24.8279
R718 GNDA.n208 GNDA.n207 24.8279
R719 GNDA.n175 GNDA.t207 24.0005
R720 GNDA.n175 GNDA.t12 24.0005
R721 GNDA.n179 GNDA.t89 24.0005
R722 GNDA.n179 GNDA.t150 24.0005
R723 GNDA.n183 GNDA.t251 24.0005
R724 GNDA.n183 GNDA.t261 24.0005
R725 GNDA.n187 GNDA.t58 24.0005
R726 GNDA.n187 GNDA.t219 24.0005
R727 GNDA.n192 GNDA.t28 24.0005
R728 GNDA.n192 GNDA.t195 24.0005
R729 GNDA.t108 GNDA.t42 23.5299
R730 GNDA.n376 GNDA.n106 23.1831
R731 GNDA.n768 GNDA.n767 22.4005
R732 GNDA.n424 GNDA.n423 22.4005
R733 GNDA.n532 GNDA.n70 22.4005
R734 GNDA.n558 GNDA.n557 22.4005
R735 GNDA.n594 GNDA.n593 22.4005
R736 GNDA.n483 GNDA.n482 20.9665
R737 GNDA.n506 GNDA.n505 19.4202
R738 GNDA.n458 GNDA.n442 19.2005
R739 GNDA.n458 GNDA.n457 19.2005
R740 GNDA.n387 GNDA.n386 19.2005
R741 GNDA.n411 GNDA.n410 19.2005
R742 GNDA.n546 GNDA.n65 19.2005
R743 GNDA.n572 GNDA.n571 19.2005
R744 GNDA.n589 GNDA.n588 19.2005
R745 GNDA.n604 GNDA.n42 19.2005
R746 GNDA.n674 GNDA.n673 19.2005
R747 GNDA.n656 GNDA.n655 19.2005
R748 GNDA.n338 GNDA.n337 19.2005
R749 GNDA.n146 GNDA.n145 19.2005
R750 GNDA.t38 GNDA.t165 17.8306
R751 GNDA.n197 GNDA.t260 17.2554
R752 GNDA.n740 GNDA.n739 16.0005
R753 GNDA.n741 GNDA.n740 16.0005
R754 GNDA.n686 GNDA.n37 16.0005
R755 GNDA.n686 GNDA.n685 16.0005
R756 GNDA.n210 GNDA 15.7005
R757 GNDA.n484 GNDA.n483 15.6449
R758 GNDA.n103 GNDA.n102 15.6449
R759 GNDA.n472 GNDA.t130 15.0005
R760 GNDA.n472 GNDA.t199 15.0005
R761 GNDA.n480 GNDA.t174 15.0005
R762 GNDA.n480 GNDA.t231 15.0005
R763 GNDA.t171 GNDA.n459 15.0005
R764 GNDA.n459 GNDA.t34 15.0005
R765 GNDA.n447 GNDA.t160 15.0005
R766 GNDA.n447 GNDA.t191 15.0005
R767 GNDA.n87 GNDA.t210 15.0005
R768 GNDA.n87 GNDA.t136 15.0005
R769 GNDA.n90 GNDA.t126 15.0005
R770 GNDA.n90 GNDA.t187 15.0005
R771 GNDA.t210 GNDA.n86 15.0005
R772 GNDA.n527 GNDA.t192 15.0005
R773 GNDA.n460 GNDA.t171 15.0005
R774 GNDA.n435 GNDA.t200 15.0005
R775 GNDA.t174 GNDA.n427 15.0005
R776 GNDA.n92 GNDA.t188 15.0005
R777 GNDA.n104 GNDA.n103 14.4005
R778 GNDA.n254 GNDA.n253 14.0805
R779 GNDA.n256 GNDA.n169 14.0805
R780 GNDA.n719 GNDA.n26 13.9181
R781 GNDA.t27 GNDA.t38 13.8044
R782 GNDA.n210 GNDA.n105 13.1958
R783 GNDA.n260 GNDA.n105 12.8163
R784 GNDA.n467 GNDA.n431 12.8005
R785 GNDA.n481 GNDA.n479 12.8005
R786 GNDA.n521 GNDA.n520 12.8005
R787 GNDA.n514 GNDA.n513 12.8005
R788 GNDA.n164 GNDA.n115 12.8005
R789 GNDA.n386 GNDA.n373 12.8005
R790 GNDA.n410 GNDA.n409 12.8005
R791 GNDA.n549 GNDA.n65 12.8005
R792 GNDA.n573 GNDA.n572 12.8005
R793 GNDA.n588 GNDA.n587 12.8005
R794 GNDA.n601 GNDA.n42 12.8005
R795 GNDA.n675 GNDA.n674 12.8005
R796 GNDA.n655 GNDA.n654 12.8005
R797 GNDA.n500 GNDA.n109 12.8005
R798 GNDA.n339 GNDA.n338 12.8005
R799 GNDA.n203 GNDA.n202 12.8005
R800 GNDA.n200 GNDA.n199 12.8005
R801 GNDA GNDA.n0 12.7806
R802 GNDA GNDA.n782 11.8829
R803 GNDA.n730 GNDA.t104 11.7652
R804 GNDA.n729 GNDA.t60 11.7652
R805 GNDA.n506 GNDA.n26 11.7212
R806 GNDA.n508 GNDA.n507 11.6542
R807 GNDA.n378 GNDA.n376 10.7016
R808 GNDA.n639 GNDA.n638 10.4505
R809 GNDA.n494 GNDA.t62 9.63554
R810 GNDA.n769 GNDA.n768 9.6005
R811 GNDA.n424 GNDA.n369 9.6005
R812 GNDA.n533 GNDA.n532 9.6005
R813 GNDA.n557 GNDA.n556 9.6005
R814 GNDA.n595 GNDA.n594 9.6005
R815 GNDA.n248 GNDA.n247 9.58175
R816 GNDA.n216 GNDA.n208 9.58175
R817 GNDA.n640 GNDA.n635 9.3005
R818 GNDA.n642 GNDA.n641 9.3005
R819 GNDA.n643 GNDA.n633 9.3005
R820 GNDA.n645 GNDA.n644 9.3005
R821 GNDA.n646 GNDA.n632 9.3005
R822 GNDA.n648 GNDA.n647 9.3005
R823 GNDA.n649 GNDA.n631 9.3005
R824 GNDA.n651 GNDA.n650 9.3005
R825 GNDA.n653 GNDA.n652 9.3005
R826 GNDA.n654 GNDA.n627 9.3005
R827 GNDA.n657 GNDA.n656 9.3005
R828 GNDA.n658 GNDA.n626 9.3005
R829 GNDA.n660 GNDA.n659 9.3005
R830 GNDA.n661 GNDA.n624 9.3005
R831 GNDA.n664 GNDA.n663 9.3005
R832 GNDA.n665 GNDA.n623 9.3005
R833 GNDA.n667 GNDA.n666 9.3005
R834 GNDA.n668 GNDA.n622 9.3005
R835 GNDA.n670 GNDA.n669 9.3005
R836 GNDA.n671 GNDA.n621 9.3005
R837 GNDA.n673 GNDA.n672 9.3005
R838 GNDA.n675 GNDA.n619 9.3005
R839 GNDA.n677 GNDA.n676 9.3005
R840 GNDA.n679 GNDA.n678 9.3005
R841 GNDA.n680 GNDA.n616 9.3005
R842 GNDA.n682 GNDA.n681 9.3005
R843 GNDA.n683 GNDA.n38 9.3005
R844 GNDA.n685 GNDA.n684 9.3005
R845 GNDA.n615 GNDA.n37 9.3005
R846 GNDA.n614 GNDA.n613 9.3005
R847 GNDA.n612 GNDA.n39 9.3005
R848 GNDA.n611 GNDA.n610 9.3005
R849 GNDA.n609 GNDA.n40 9.3005
R850 GNDA.n608 GNDA.n607 9.3005
R851 GNDA.n605 GNDA.n41 9.3005
R852 GNDA.n604 GNDA.n603 9.3005
R853 GNDA.n602 GNDA.n601 9.3005
R854 GNDA.n600 GNDA.n43 9.3005
R855 GNDA.n599 GNDA.n598 9.3005
R856 GNDA.n597 GNDA.n596 9.3005
R857 GNDA.n595 GNDA.n46 9.3005
R858 GNDA.n593 GNDA.n592 9.3005
R859 GNDA.n591 GNDA.n48 9.3005
R860 GNDA.n590 GNDA.n589 9.3005
R861 GNDA.n587 GNDA.n49 9.3005
R862 GNDA.n586 GNDA.n585 9.3005
R863 GNDA.n584 GNDA.n51 9.3005
R864 GNDA.n583 GNDA.n582 9.3005
R865 GNDA.n581 GNDA.n52 9.3005
R866 GNDA.n580 GNDA.n579 9.3005
R867 GNDA.n578 GNDA.n53 9.3005
R868 GNDA.n577 GNDA.n576 9.3005
R869 GNDA.n573 GNDA.n54 9.3005
R870 GNDA.n571 GNDA.n570 9.3005
R871 GNDA.n569 GNDA.n56 9.3005
R872 GNDA.n568 GNDA.n567 9.3005
R873 GNDA.n566 GNDA.n57 9.3005
R874 GNDA.n565 GNDA.n564 9.3005
R875 GNDA.n563 GNDA.n58 9.3005
R876 GNDA.n562 GNDA.n561 9.3005
R877 GNDA.n558 GNDA.n59 9.3005
R878 GNDA.n556 GNDA.n555 9.3005
R879 GNDA.n554 GNDA.n61 9.3005
R880 GNDA.n553 GNDA.n552 9.3005
R881 GNDA.n550 GNDA.n62 9.3005
R882 GNDA.n549 GNDA.n548 9.3005
R883 GNDA.n547 GNDA.n546 9.3005
R884 GNDA.n545 GNDA.n66 9.3005
R885 GNDA.n544 GNDA.n543 9.3005
R886 GNDA.n542 GNDA.n67 9.3005
R887 GNDA.n541 GNDA.n540 9.3005
R888 GNDA.n538 GNDA.n68 9.3005
R889 GNDA.n537 GNDA.n536 9.3005
R890 GNDA.n535 GNDA.n70 9.3005
R891 GNDA.n534 GNDA.n533 9.3005
R892 GNDA.n72 GNDA.n71 9.3005
R893 GNDA.n406 GNDA.n405 9.3005
R894 GNDA.n407 GNDA.n402 9.3005
R895 GNDA.n409 GNDA.n408 9.3005
R896 GNDA.n411 GNDA.n400 9.3005
R897 GNDA.n413 GNDA.n412 9.3005
R898 GNDA.n414 GNDA.n399 9.3005
R899 GNDA.n416 GNDA.n415 9.3005
R900 GNDA.n417 GNDA.n397 9.3005
R901 GNDA.n420 GNDA.n419 9.3005
R902 GNDA.n421 GNDA.n370 9.3005
R903 GNDA.n423 GNDA.n422 9.3005
R904 GNDA.n396 GNDA.n369 9.3005
R905 GNDA.n395 GNDA.n394 9.3005
R906 GNDA.n393 GNDA.n371 9.3005
R907 GNDA.n391 GNDA.n390 9.3005
R908 GNDA.n389 GNDA.n373 9.3005
R909 GNDA.n388 GNDA.n387 9.3005
R910 GNDA.n384 GNDA.n374 9.3005
R911 GNDA.n383 GNDA.n382 9.3005
R912 GNDA.n381 GNDA.n375 9.3005
R913 GNDA.n380 GNDA.n379 9.3005
R914 GNDA.n148 GNDA.n147 9.3005
R915 GNDA.n149 GNDA.n118 9.3005
R916 GNDA.n151 GNDA.n150 9.3005
R917 GNDA.n152 GNDA.n117 9.3005
R918 GNDA.n154 GNDA.n153 9.3005
R919 GNDA.n155 GNDA.n115 9.3005
R920 GNDA.n162 GNDA.n116 9.3005
R921 GNDA.n161 GNDA.n160 9.3005
R922 GNDA.n159 GNDA.n156 9.3005
R923 GNDA.n158 GNDA.n157 9.3005
R924 GNDA.n109 GNDA.n108 9.3005
R925 GNDA.n504 GNDA.n503 9.3005
R926 GNDA.n502 GNDA.n107 9.3005
R927 GNDA.n501 GNDA.n500 9.3005
R928 GNDA.n164 GNDA.n163 9.3005
R929 GNDA.n314 GNDA.n313 9.3005
R930 GNDA.n301 GNDA.n300 9.3005
R931 GNDA.n302 GNDA.n290 9.3005
R932 GNDA.n304 GNDA.n303 9.3005
R933 GNDA.n305 GNDA.n289 9.3005
R934 GNDA.n307 GNDA.n306 9.3005
R935 GNDA.n308 GNDA.n288 9.3005
R936 GNDA.n310 GNDA.n309 9.3005
R937 GNDA.n311 GNDA.n285 9.3005
R938 GNDA.n315 GNDA.n284 9.3005
R939 GNDA.n317 GNDA.n316 9.3005
R940 GNDA.n318 GNDA.n283 9.3005
R941 GNDA.n320 GNDA.n319 9.3005
R942 GNDA.n321 GNDA.n282 9.3005
R943 GNDA.n323 GNDA.n322 9.3005
R944 GNDA.n324 GNDA.n280 9.3005
R945 GNDA.n326 GNDA.n325 9.3005
R946 GNDA.n327 GNDA.n279 9.3005
R947 GNDA.n329 GNDA.n328 9.3005
R948 GNDA.n330 GNDA.n277 9.3005
R949 GNDA.n333 GNDA.n332 9.3005
R950 GNDA.n334 GNDA.n276 9.3005
R951 GNDA.n336 GNDA.n335 9.3005
R952 GNDA.n337 GNDA.n274 9.3005
R953 GNDA.n340 GNDA.n339 9.3005
R954 GNDA.n341 GNDA.n273 9.3005
R955 GNDA.n343 GNDA.n342 9.3005
R956 GNDA.n345 GNDA.n268 9.3005
R957 GNDA.n347 GNDA.n346 9.3005
R958 GNDA.n348 GNDA.n267 9.3005
R959 GNDA.n350 GNDA.n349 9.3005
R960 GNDA.n351 GNDA.n265 9.3005
R961 GNDA.n354 GNDA.n353 9.3005
R962 GNDA.n355 GNDA.n264 9.3005
R963 GNDA.n357 GNDA.n356 9.3005
R964 GNDA.n358 GNDA.n262 9.3005
R965 GNDA.n361 GNDA.n360 9.3005
R966 GNDA.n362 GNDA.n261 9.3005
R967 GNDA.n364 GNDA.n363 9.3005
R968 GNDA.n246 GNDA.n245 9.3005
R969 GNDA.n244 GNDA.n173 9.3005
R970 GNDA.n243 GNDA.n242 9.3005
R971 GNDA.n241 GNDA.n174 9.3005
R972 GNDA.n240 GNDA.n239 9.3005
R973 GNDA.n238 GNDA.n177 9.3005
R974 GNDA.n237 GNDA.n236 9.3005
R975 GNDA.n235 GNDA.n178 9.3005
R976 GNDA.n234 GNDA.n233 9.3005
R977 GNDA.n232 GNDA.n181 9.3005
R978 GNDA.n231 GNDA.n230 9.3005
R979 GNDA.n229 GNDA.n182 9.3005
R980 GNDA.n228 GNDA.n227 9.3005
R981 GNDA.n226 GNDA.n185 9.3005
R982 GNDA.n225 GNDA.n224 9.3005
R983 GNDA.n223 GNDA.n186 9.3005
R984 GNDA.n222 GNDA.n221 9.3005
R985 GNDA.n220 GNDA.n189 9.3005
R986 GNDA.n219 GNDA.n218 9.3005
R987 GNDA.n217 GNDA.n191 9.3005
R988 GNDA.n215 GNDA.n214 9.3005
R989 GNDA.n213 GNDA.n209 9.3005
R990 GNDA.n212 GNDA.n211 9.3005
R991 GNDA.n146 GNDA.n119 9.3005
R992 GNDA.n134 GNDA.n130 9.3005
R993 GNDA.n136 GNDA.n135 9.3005
R994 GNDA.n137 GNDA.n129 9.3005
R995 GNDA.n139 GNDA.n138 9.3005
R996 GNDA.n140 GNDA.n128 9.3005
R997 GNDA.n142 GNDA.n141 9.3005
R998 GNDA.n143 GNDA.n127 9.3005
R999 GNDA.n145 GNDA.n144 9.3005
R1000 GNDA.n510 GNDA.n509 9.3005
R1001 GNDA.n511 GNDA.n104 9.3005
R1002 GNDA.n513 GNDA.n512 9.3005
R1003 GNDA.n514 GNDA.n89 9.3005
R1004 GNDA.n516 GNDA.n515 9.3005
R1005 GNDA.n517 GNDA.n88 9.3005
R1006 GNDA.n519 GNDA.n518 9.3005
R1007 GNDA.n520 GNDA.n85 9.3005
R1008 GNDA.n522 GNDA.n521 9.3005
R1009 GNDA.n523 GNDA.n83 9.3005
R1010 GNDA.n525 GNDA.n524 9.3005
R1011 GNDA.n479 GNDA.n428 9.3005
R1012 GNDA.n478 GNDA.n477 9.3005
R1013 GNDA.n476 GNDA.n429 9.3005
R1014 GNDA.n475 GNDA.n474 9.3005
R1015 GNDA.n473 GNDA.n430 9.3005
R1016 GNDA.n471 GNDA.n470 9.3005
R1017 GNDA.n469 GNDA.n431 9.3005
R1018 GNDA.n468 GNDA.n467 9.3005
R1019 GNDA.n433 GNDA.n432 9.3005
R1020 GNDA.n443 GNDA.n442 9.3005
R1021 GNDA.n458 GNDA.n444 9.3005
R1022 GNDA.n457 GNDA.n456 9.3005
R1023 GNDA.n455 GNDA.n445 9.3005
R1024 GNDA.n454 GNDA.n453 9.3005
R1025 GNDA.n452 GNDA.n446 9.3005
R1026 GNDA.n451 GNDA.n450 9.3005
R1027 GNDA.n449 GNDA.n448 9.3005
R1028 GNDA.n84 GNDA.n82 9.3005
R1029 GNDA.n718 GNDA.n717 9.3005
R1030 GNDA.n716 GNDA.n27 9.3005
R1031 GNDA.n715 GNDA.n714 9.3005
R1032 GNDA.n713 GNDA.n28 9.3005
R1033 GNDA.n712 GNDA.n711 9.3005
R1034 GNDA.n710 GNDA.n29 9.3005
R1035 GNDA.n709 GNDA.n708 9.3005
R1036 GNDA.n707 GNDA.n30 9.3005
R1037 GNDA.n706 GNDA.n705 9.3005
R1038 GNDA.n704 GNDA.n32 9.3005
R1039 GNDA.n702 GNDA.n701 9.3005
R1040 GNDA.n700 GNDA.n33 9.3005
R1041 GNDA.n699 GNDA.n698 9.3005
R1042 GNDA.n697 GNDA.n34 9.3005
R1043 GNDA.n696 GNDA.n695 9.3005
R1044 GNDA.n694 GNDA.n35 9.3005
R1045 GNDA.n693 GNDA.n692 9.3005
R1046 GNDA.n22 GNDA.n21 9.3005
R1047 GNDA.n735 GNDA.n734 9.3005
R1048 GNDA.n736 GNDA.n20 9.3005
R1049 GNDA.n738 GNDA.n737 9.3005
R1050 GNDA.n739 GNDA.n18 9.3005
R1051 GNDA.n742 GNDA.n741 9.3005
R1052 GNDA.n743 GNDA.n17 9.3005
R1053 GNDA.n745 GNDA.n744 9.3005
R1054 GNDA.n747 GNDA.n15 9.3005
R1055 GNDA.n749 GNDA.n748 9.3005
R1056 GNDA.n750 GNDA.n14 9.3005
R1057 GNDA.n752 GNDA.n751 9.3005
R1058 GNDA.n754 GNDA.n12 9.3005
R1059 GNDA.n756 GNDA.n755 9.3005
R1060 GNDA.n757 GNDA.n11 9.3005
R1061 GNDA.n759 GNDA.n758 9.3005
R1062 GNDA.n760 GNDA.n10 9.3005
R1063 GNDA.n762 GNDA.n761 9.3005
R1064 GNDA.n763 GNDA.n9 9.3005
R1065 GNDA.n765 GNDA.n764 9.3005
R1066 GNDA.n767 GNDA.n6 9.3005
R1067 GNDA.n770 GNDA.n769 9.3005
R1068 GNDA.n771 GNDA.n5 9.3005
R1069 GNDA.n773 GNDA.n772 9.3005
R1070 GNDA.n774 GNDA.n4 9.3005
R1071 GNDA.n776 GNDA.n775 9.3005
R1072 GNDA.n777 GNDA.n3 9.3005
R1073 GNDA.n779 GNDA.n778 9.3005
R1074 GNDA.n780 GNDA.n1 9.3005
R1075 GNDA.t88 GNDA.t51 8.62795
R1076 GNDA.t176 GNDA.t194 8.62795
R1077 GNDA.n365 GNDA.n260 7.49888
R1078 GNDA.n489 GNDA.n488 7.11161
R1079 GNDA.n486 GNDA.n484 7.11161
R1080 GNDA.n98 GNDA.n97 7.11161
R1081 GNDA.n102 GNDA.n91 7.11161
R1082 GNDA.n482 GNDA.n481 6.69883
R1083 GNDA.n474 GNDA.n473 6.4005
R1084 GNDA.n452 GNDA.n451 6.4005
R1085 GNDA.n525 GNDA.n82 6.4005
R1086 GNDA.n695 GNDA.n691 6.4005
R1087 GNDA.n734 GNDA.n733 6.4005
R1088 GNDA.n747 GNDA.n746 6.4005
R1089 GNDA.n754 GNDA.n753 6.4005
R1090 GNDA.n766 GNDA.n765 6.4005
R1091 GNDA.n781 GNDA.n780 6.4005
R1092 GNDA.n393 GNDA.n392 6.4005
R1093 GNDA.n405 GNDA.n404 6.4005
R1094 GNDA.n552 GNDA.n551 6.4005
R1095 GNDA.n575 GNDA.n53 6.4005
R1096 GNDA.n679 GNDA.n618 6.4005
R1097 GNDA.n663 GNDA.n662 6.4005
R1098 GNDA.n650 GNDA.n630 6.4005
R1099 GNDA.n634 GNDA.n632 6.4005
R1100 GNDA.n352 GNDA.n351 6.4005
R1101 GNDA.n331 GNDA.n330 6.4005
R1102 GNDA.n325 GNDA.n281 6.4005
R1103 GNDA.n286 GNDA.n284 6.4005
R1104 GNDA.n312 GNDA.n311 6.4005
R1105 GNDA.n300 GNDA.n299 6.4005
R1106 GNDA.n190 GNDA.n186 6.4005
R1107 GNDA.n509 GNDA.n104 6.4005
R1108 GNDA.n726 GNDA.n8 5.68939
R1109 GNDA.n296 GNDA.n295 5.68939
R1110 GNDA.n296 GNDA.n287 5.68939
R1111 GNDA.n726 GNDA.n7 4.97828
R1112 GNDA.n165 GNDA.n114 4.49344
R1113 GNDA.n111 GNDA.n110 4.49344
R1114 GNDA.n499 GNDA.n110 4.49344
R1115 GNDA.n166 GNDA.n165 4.49344
R1116 GNDA.n496 GNDA.n495 3.8278
R1117 GNDA.n113 GNDA.n112 3.8278
R1118 GNDA.n124 GNDA.n123 3.8278
R1119 GNDA.n488 GNDA.n487 3.48951
R1120 GNDA.n487 GNDA.n486 3.48951
R1121 GNDA.n97 GNDA.n96 3.48951
R1122 GNDA.n96 GNDA.n91 3.48951
R1123 GNDA.n419 GNDA.n418 3.2005
R1124 GNDA.n539 GNDA.n538 3.2005
R1125 GNDA.n560 GNDA.n58 3.2005
R1126 GNDA.n599 GNDA.n45 3.2005
R1127 GNDA.n606 GNDA.n40 3.2005
R1128 GNDA.n359 GNDA.n358 3.2005
R1129 GNDA.n345 GNDA.n344 3.2005
R1130 GNDA.t206 GNDA.t37 2.88386
R1131 GNDA.n125 GNDA.n121 2.8779
R1132 GNDA.n126 GNDA.n121 2.8779
R1133 GNDA.t161 GNDA.t218 2.87632
R1134 GNDA.n77 GNDA.n76 2.25882
R1135 GNDA.n78 GNDA.n77 2.25882
R1136 GNDA.n526 GNDA.n81 2.25882
R1137 GNDA.n80 GNDA.n78 2.25882
R1138 GNDA.n528 GNDA.n76 2.25882
R1139 GNDA.n81 GNDA.n80 2.25882
R1140 GNDA.n461 GNDA.n441 2.25882
R1141 GNDA.n441 GNDA.n440 2.25882
R1142 GNDA.n466 GNDA.n434 2.25882
R1143 GNDA.n440 GNDA.n439 2.25882
R1144 GNDA.n462 GNDA.n461 2.25882
R1145 GNDA.n439 GNDA.n434 2.25882
R1146 GNDA.n507 GNDA.n105 0.9875
R1147 GNDA.n482 GNDA.n428 0.703977
R1148 GNDA.n640 GNDA.n639 0.442364
R1149 GNDA.n363 GNDA.n260 0.193977
R1150 GNDA.n301 GNDA.n0 0.193881
R1151 GNDA.n782 GNDA.n1 0.193881
R1152 GNDA.n717 GNDA.n26 0.193695
R1153 GNDA.n380 GNDA.n376 0.193477
R1154 GNDA.n211 GNDA.n210 0.188
R1155 GNDA.n133 GNDA 0.162727
R1156 GNDA.n381 GNDA.n380 0.15675
R1157 GNDA.n382 GNDA.n381 0.15675
R1158 GNDA.n382 GNDA.n374 0.15675
R1159 GNDA.n388 GNDA.n374 0.15675
R1160 GNDA.n389 GNDA.n388 0.15675
R1161 GNDA.n390 GNDA.n389 0.15675
R1162 GNDA.n390 GNDA.n371 0.15675
R1163 GNDA.n395 GNDA.n371 0.15675
R1164 GNDA.n396 GNDA.n395 0.15675
R1165 GNDA.n422 GNDA.n396 0.15675
R1166 GNDA.n422 GNDA.n421 0.15675
R1167 GNDA.n421 GNDA.n420 0.15675
R1168 GNDA.n420 GNDA.n397 0.15675
R1169 GNDA.n415 GNDA.n397 0.15675
R1170 GNDA.n415 GNDA.n414 0.15675
R1171 GNDA.n414 GNDA.n413 0.15675
R1172 GNDA.n413 GNDA.n400 0.15675
R1173 GNDA.n408 GNDA.n400 0.15675
R1174 GNDA.n408 GNDA.n407 0.15675
R1175 GNDA.n407 GNDA.n406 0.15675
R1176 GNDA.n406 GNDA.n71 0.15675
R1177 GNDA.n534 GNDA.n71 0.15675
R1178 GNDA.n535 GNDA.n534 0.15675
R1179 GNDA.n536 GNDA.n535 0.15675
R1180 GNDA.n536 GNDA.n68 0.15675
R1181 GNDA.n541 GNDA.n68 0.15675
R1182 GNDA.n542 GNDA.n541 0.15675
R1183 GNDA.n543 GNDA.n542 0.15675
R1184 GNDA.n543 GNDA.n66 0.15675
R1185 GNDA.n547 GNDA.n66 0.15675
R1186 GNDA.n548 GNDA.n547 0.15675
R1187 GNDA.n548 GNDA.n62 0.15675
R1188 GNDA.n553 GNDA.n62 0.15675
R1189 GNDA.n554 GNDA.n553 0.15675
R1190 GNDA.n555 GNDA.n554 0.15675
R1191 GNDA.n555 GNDA.n59 0.15675
R1192 GNDA.n562 GNDA.n59 0.15675
R1193 GNDA.n563 GNDA.n562 0.15675
R1194 GNDA.n564 GNDA.n563 0.15675
R1195 GNDA.n564 GNDA.n57 0.15675
R1196 GNDA.n568 GNDA.n57 0.15675
R1197 GNDA.n569 GNDA.n568 0.15675
R1198 GNDA.n570 GNDA.n569 0.15675
R1199 GNDA.n570 GNDA.n54 0.15675
R1200 GNDA.n577 GNDA.n54 0.15675
R1201 GNDA.n578 GNDA.n577 0.15675
R1202 GNDA.n579 GNDA.n578 0.15675
R1203 GNDA.n579 GNDA.n52 0.15675
R1204 GNDA.n583 GNDA.n52 0.15675
R1205 GNDA.n584 GNDA.n583 0.15675
R1206 GNDA.n585 GNDA.n584 0.15675
R1207 GNDA.n585 GNDA.n49 0.15675
R1208 GNDA.n590 GNDA.n49 0.15675
R1209 GNDA.n591 GNDA.n590 0.15675
R1210 GNDA.n592 GNDA.n591 0.15675
R1211 GNDA.n592 GNDA.n46 0.15675
R1212 GNDA.n597 GNDA.n46 0.15675
R1213 GNDA.n598 GNDA.n597 0.15675
R1214 GNDA.n598 GNDA.n43 0.15675
R1215 GNDA.n602 GNDA.n43 0.15675
R1216 GNDA.n603 GNDA.n602 0.15675
R1217 GNDA.n603 GNDA.n41 0.15675
R1218 GNDA.n608 GNDA.n41 0.15675
R1219 GNDA.n609 GNDA.n608 0.15675
R1220 GNDA.n610 GNDA.n609 0.15675
R1221 GNDA.n610 GNDA.n39 0.15675
R1222 GNDA.n614 GNDA.n39 0.15675
R1223 GNDA.n615 GNDA.n614 0.15675
R1224 GNDA.n684 GNDA.n615 0.15675
R1225 GNDA.n684 GNDA.n683 0.15675
R1226 GNDA.n683 GNDA.n682 0.15675
R1227 GNDA.n682 GNDA.n616 0.15675
R1228 GNDA.n678 GNDA.n616 0.15675
R1229 GNDA.n678 GNDA.n677 0.15675
R1230 GNDA.n677 GNDA.n619 0.15675
R1231 GNDA.n672 GNDA.n619 0.15675
R1232 GNDA.n672 GNDA.n671 0.15675
R1233 GNDA.n671 GNDA.n670 0.15675
R1234 GNDA.n670 GNDA.n622 0.15675
R1235 GNDA.n666 GNDA.n622 0.15675
R1236 GNDA.n666 GNDA.n665 0.15675
R1237 GNDA.n665 GNDA.n664 0.15675
R1238 GNDA.n664 GNDA.n624 0.15675
R1239 GNDA.n659 GNDA.n624 0.15675
R1240 GNDA.n659 GNDA.n658 0.15675
R1241 GNDA.n658 GNDA.n657 0.15675
R1242 GNDA.n657 GNDA.n627 0.15675
R1243 GNDA.n652 GNDA.n627 0.15675
R1244 GNDA.n652 GNDA.n651 0.15675
R1245 GNDA.n651 GNDA.n631 0.15675
R1246 GNDA.n647 GNDA.n631 0.15675
R1247 GNDA.n647 GNDA.n646 0.15675
R1248 GNDA.n646 GNDA.n645 0.15675
R1249 GNDA.n645 GNDA.n633 0.15675
R1250 GNDA.n641 GNDA.n633 0.15675
R1251 GNDA.n641 GNDA.n640 0.15675
R1252 GNDA.n136 GNDA.n130 0.15675
R1253 GNDA.n137 GNDA.n136 0.15675
R1254 GNDA.n138 GNDA.n137 0.15675
R1255 GNDA.n138 GNDA.n128 0.15675
R1256 GNDA.n142 GNDA.n128 0.15675
R1257 GNDA.n143 GNDA.n142 0.15675
R1258 GNDA.n144 GNDA.n143 0.15675
R1259 GNDA.n144 GNDA.n119 0.15675
R1260 GNDA.n148 GNDA.n119 0.15675
R1261 GNDA.n149 GNDA.n148 0.15675
R1262 GNDA.n150 GNDA.n149 0.15675
R1263 GNDA.n150 GNDA.n117 0.15675
R1264 GNDA.n154 GNDA.n117 0.15675
R1265 GNDA.n155 GNDA.n154 0.15675
R1266 GNDA.n163 GNDA.n155 0.15675
R1267 GNDA.n163 GNDA.n162 0.15675
R1268 GNDA.n162 GNDA.n161 0.15675
R1269 GNDA.n161 GNDA.n156 0.15675
R1270 GNDA.n157 GNDA.n156 0.15675
R1271 GNDA.n157 GNDA.n108 0.15675
R1272 GNDA.n501 GNDA.n108 0.15675
R1273 GNDA.n502 GNDA.n501 0.15675
R1274 GNDA.n503 GNDA.n502 0.15675
R1275 GNDA.n363 GNDA.n362 0.15675
R1276 GNDA.n362 GNDA.n361 0.15675
R1277 GNDA.n361 GNDA.n262 0.15675
R1278 GNDA.n356 GNDA.n262 0.15675
R1279 GNDA.n356 GNDA.n355 0.15675
R1280 GNDA.n355 GNDA.n354 0.15675
R1281 GNDA.n354 GNDA.n265 0.15675
R1282 GNDA.n349 GNDA.n265 0.15675
R1283 GNDA.n349 GNDA.n348 0.15675
R1284 GNDA.n348 GNDA.n347 0.15675
R1285 GNDA.n347 GNDA.n268 0.15675
R1286 GNDA.n342 GNDA.n268 0.15675
R1287 GNDA.n342 GNDA.n341 0.15675
R1288 GNDA.n341 GNDA.n340 0.15675
R1289 GNDA.n340 GNDA.n274 0.15675
R1290 GNDA.n335 GNDA.n274 0.15675
R1291 GNDA.n335 GNDA.n334 0.15675
R1292 GNDA.n334 GNDA.n333 0.15675
R1293 GNDA.n333 GNDA.n277 0.15675
R1294 GNDA.n328 GNDA.n277 0.15675
R1295 GNDA.n328 GNDA.n327 0.15675
R1296 GNDA.n327 GNDA.n326 0.15675
R1297 GNDA.n326 GNDA.n280 0.15675
R1298 GNDA.n322 GNDA.n280 0.15675
R1299 GNDA.n322 GNDA.n321 0.15675
R1300 GNDA.n321 GNDA.n320 0.15675
R1301 GNDA.n320 GNDA.n283 0.15675
R1302 GNDA.n316 GNDA.n283 0.15675
R1303 GNDA.n316 GNDA.n315 0.15675
R1304 GNDA.n315 GNDA.n314 0.15675
R1305 GNDA.n314 GNDA.n285 0.15675
R1306 GNDA.n309 GNDA.n285 0.15675
R1307 GNDA.n309 GNDA.n308 0.15675
R1308 GNDA.n308 GNDA.n307 0.15675
R1309 GNDA.n307 GNDA.n289 0.15675
R1310 GNDA.n303 GNDA.n289 0.15675
R1311 GNDA.n303 GNDA.n302 0.15675
R1312 GNDA.n302 GNDA.n301 0.15675
R1313 GNDA.n246 GNDA.n173 0.15675
R1314 GNDA.n242 GNDA.n241 0.15675
R1315 GNDA.n241 GNDA.n240 0.15675
R1316 GNDA.n240 GNDA.n177 0.15675
R1317 GNDA.n236 GNDA.n235 0.15675
R1318 GNDA.n235 GNDA.n234 0.15675
R1319 GNDA.n234 GNDA.n181 0.15675
R1320 GNDA.n230 GNDA.n229 0.15675
R1321 GNDA.n229 GNDA.n228 0.15675
R1322 GNDA.n228 GNDA.n185 0.15675
R1323 GNDA.n224 GNDA.n223 0.15675
R1324 GNDA.n223 GNDA.n222 0.15675
R1325 GNDA.n222 GNDA.n189 0.15675
R1326 GNDA.n218 GNDA.n217 0.15675
R1327 GNDA.n215 GNDA.n209 0.15675
R1328 GNDA.n211 GNDA.n209 0.15675
R1329 GNDA.n477 GNDA.n428 0.15675
R1330 GNDA.n477 GNDA.n476 0.15675
R1331 GNDA.n476 GNDA.n475 0.15675
R1332 GNDA.n475 GNDA.n430 0.15675
R1333 GNDA.n470 GNDA.n430 0.15675
R1334 GNDA.n470 GNDA.n469 0.15675
R1335 GNDA.n469 GNDA.n468 0.15675
R1336 GNDA.n468 GNDA.n432 0.15675
R1337 GNDA.n443 GNDA.n432 0.15675
R1338 GNDA.n444 GNDA.n443 0.15675
R1339 GNDA.n456 GNDA.n444 0.15675
R1340 GNDA.n456 GNDA.n455 0.15675
R1341 GNDA.n455 GNDA.n454 0.15675
R1342 GNDA.n454 GNDA.n446 0.15675
R1343 GNDA.n450 GNDA.n446 0.15675
R1344 GNDA.n450 GNDA.n449 0.15675
R1345 GNDA.n449 GNDA.n84 0.15675
R1346 GNDA.n524 GNDA.n84 0.15675
R1347 GNDA.n524 GNDA.n523 0.15675
R1348 GNDA.n523 GNDA.n522 0.15675
R1349 GNDA.n522 GNDA.n85 0.15675
R1350 GNDA.n518 GNDA.n85 0.15675
R1351 GNDA.n518 GNDA.n517 0.15675
R1352 GNDA.n517 GNDA.n516 0.15675
R1353 GNDA.n516 GNDA.n89 0.15675
R1354 GNDA.n512 GNDA.n89 0.15675
R1355 GNDA.n512 GNDA.n511 0.15675
R1356 GNDA.n511 GNDA.n510 0.15675
R1357 GNDA.n717 GNDA.n716 0.15675
R1358 GNDA.n716 GNDA.n715 0.15675
R1359 GNDA.n715 GNDA.n28 0.15675
R1360 GNDA.n711 GNDA.n28 0.15675
R1361 GNDA.n711 GNDA.n710 0.15675
R1362 GNDA.n710 GNDA.n709 0.15675
R1363 GNDA.n709 GNDA.n30 0.15675
R1364 GNDA.n705 GNDA.n30 0.15675
R1365 GNDA.n705 GNDA.n704 0.15675
R1366 GNDA.n702 GNDA.n33 0.15675
R1367 GNDA.n698 GNDA.n33 0.15675
R1368 GNDA.n698 GNDA.n697 0.15675
R1369 GNDA.n697 GNDA.n696 0.15675
R1370 GNDA.n696 GNDA.n35 0.15675
R1371 GNDA.n692 GNDA.n35 0.15675
R1372 GNDA.n692 GNDA.n21 0.15675
R1373 GNDA.n735 GNDA.n21 0.15675
R1374 GNDA.n736 GNDA.n735 0.15675
R1375 GNDA.n737 GNDA.n736 0.15675
R1376 GNDA.n737 GNDA.n18 0.15675
R1377 GNDA.n742 GNDA.n18 0.15675
R1378 GNDA.n743 GNDA.n742 0.15675
R1379 GNDA.n744 GNDA.n743 0.15675
R1380 GNDA.n744 GNDA.n15 0.15675
R1381 GNDA.n749 GNDA.n15 0.15675
R1382 GNDA.n750 GNDA.n749 0.15675
R1383 GNDA.n751 GNDA.n750 0.15675
R1384 GNDA.n751 GNDA.n12 0.15675
R1385 GNDA.n756 GNDA.n12 0.15675
R1386 GNDA.n757 GNDA.n756 0.15675
R1387 GNDA.n758 GNDA.n757 0.15675
R1388 GNDA.n758 GNDA.n10 0.15675
R1389 GNDA.n762 GNDA.n10 0.15675
R1390 GNDA.n763 GNDA.n762 0.15675
R1391 GNDA.n764 GNDA.n763 0.15675
R1392 GNDA.n764 GNDA.n6 0.15675
R1393 GNDA.n770 GNDA.n6 0.15675
R1394 GNDA.n771 GNDA.n770 0.15675
R1395 GNDA.n772 GNDA.n771 0.15675
R1396 GNDA.n772 GNDA.n4 0.15675
R1397 GNDA.n776 GNDA.n4 0.15675
R1398 GNDA.n777 GNDA.n776 0.15675
R1399 GNDA.n778 GNDA.n777 0.15675
R1400 GNDA.n778 GNDA.n1 0.15675
R1401 GNDA.n503 GNDA.n106 0.141125
R1402 GNDA.n507 GNDA.n506 0.1321
R1403 GNDA.n247 GNDA.n170 0.131895
R1404 GNDA.n510 GNDA 0.1255
R1405 GNDA.n704 GNDA.n703 0.109875
R1406 GNDA.n176 GNDA.n173 0.09425
R1407 GNDA.n180 GNDA.n177 0.09425
R1408 GNDA.n184 GNDA.n181 0.09425
R1409 GNDA.n188 GNDA.n185 0.09425
R1410 GNDA.n193 GNDA.n189 0.09425
R1411 GNDA.n217 GNDA.n216 0.09425
R1412 GNDA.n247 GNDA.n246 0.063
R1413 GNDA.n242 GNDA.n176 0.063
R1414 GNDA.n236 GNDA.n180 0.063
R1415 GNDA.n230 GNDA.n184 0.063
R1416 GNDA.n224 GNDA.n188 0.063
R1417 GNDA.n218 GNDA.n193 0.063
R1418 GNDA.n216 GNDA.n215 0.063
R1419 GNDA.n508 GNDA 0.063
R1420 GNDA.n703 GNDA.n702 0.047375
R1421 GNDA.n505 GNDA.n106 0.0430057
R1422 GNDA GNDA.n130 0.03175
R1423 V_CONT.n10 V_CONT.t11 1156.8
R1424 V_CONT.n11 V_CONT.n10 964
R1425 VCO_FD_magic_0.V_CONT V_CONT.n12 562.333
R1426 V_CONT.n12 V_CONT.n11 433.8
R1427 V_CONT.n1 V_CONT.t8 377.567
R1428 V_CONT.n0 V_CONT.t12 297.233
R1429 V_CONT.n5 V_CONT.n4 242.903
R1430 V_CONT.n2 V_CONT.n0 237.851
R1431 V_CONT.n2 V_CONT.n1 232.809
R1432 V_CONT.n1 V_CONT.t9 216.9
R1433 V_CONT.n12 V_CONT.t10 192.8
R1434 V_CONT.n11 V_CONT.t14 192.8
R1435 V_CONT.n10 V_CONT.t15 192.8
R1436 V_CONT.n5 V_CONT.n3 172.502
R1437 V_CONT.n13 VCO_FD_magic_0.V_CONT 168.037
R1438 V_CONT.n8 V_CONT.t1 164.118
R1439 V_CONT.n0 V_CONT.t13 136.567
R1440 V_CONT.n15 V_CONT.n7 118.35
R1441 V_CONT.n7 V_CONT.n6 106.662
R1442 opamp_cell_4_0.VIN- V_CONT.n15 50.938
R1443 V_CONT.n3 V_CONT.t3 24.6255
R1444 V_CONT.n3 V_CONT.t0 24.6255
R1445 V_CONT.n4 V_CONT.t7 24.6255
R1446 V_CONT.n4 V_CONT.t2 24.6255
R1447 V_CONT.n7 V_CONT.n5 22.4005
R1448 V_CONT.n6 V_CONT.t6 15.0005
R1449 V_CONT.n6 V_CONT.t4 15.0005
R1450 V_CONT.n15 V_CONT.n14 9.45883
R1451 V_CONT.n14 V_CONT.n13 4.5005
R1452 V_CONT.n9 V_CONT.n8 4.5005
R1453 V_CONT.n9 V_CONT.t5 3.746
R1454 opamp_cell_4_0.VIN- V_CONT.n2 1.39633
R1455 V_CONT.n13 V_CONT.n9 0.172375
R1456 V_CONT.n14 V_CONT.n8 0.172375
R1457 a_5970_4630.n8 a_5970_4630.n6 522.322
R1458 a_5970_4630.n3 a_5970_4630.t8 384.967
R1459 a_5970_4630.n0 a_5970_4630.t11 384.967
R1460 a_5970_4630.n3 a_5970_4630.t10 379.166
R1461 a_5970_4630.t12 a_5970_4630.n0 376.56
R1462 a_5970_4630.n5 a_5970_4630.n1 315.647
R1463 a_5970_4630.n4 a_5970_4630.n2 315.647
R1464 a_5970_4630.n11 a_5970_4630.n10 314.502
R1465 a_5970_4630.n8 a_5970_4630.n7 160.721
R1466 a_5970_4630.n5 a_5970_4630.n4 83.2005
R1467 a_5970_4630.n1 a_5970_4630.t1 49.2505
R1468 a_5970_4630.n1 a_5970_4630.t7 49.2505
R1469 a_5970_4630.n2 a_5970_4630.t6 49.2505
R1470 a_5970_4630.n2 a_5970_4630.t9 49.2505
R1471 a_5970_4630.t12 a_5970_4630.n11 49.2505
R1472 a_5970_4630.n11 a_5970_4630.t2 49.2505
R1473 a_5970_4630.n10 a_5970_4630.n9 42.6672
R1474 a_5970_4630.n9 a_5970_4630.n8 37.763
R1475 a_5970_4630.n9 a_5970_4630.n5 23.4672
R1476 a_5970_4630.n6 a_5970_4630.t5 19.7005
R1477 a_5970_4630.n6 a_5970_4630.t0 19.7005
R1478 a_5970_4630.n7 a_5970_4630.t4 19.7005
R1479 a_5970_4630.n7 a_5970_4630.t3 19.7005
R1480 a_5970_4630.n4 a_5970_4630.n3 16.0005
R1481 a_5970_4630.n10 a_5970_4630.n0 16.0005
R1482 VDDA.t136 VDDA.t58 2804.76
R1483 VDDA.t14 VDDA.t44 2533.33
R1484 VDDA.t194 VDDA.t199 2307.14
R1485 VDDA.t210 VDDA.t0 2216.67
R1486 VDDA.t40 VDDA.t54 2216.67
R1487 VDDA.t197 VDDA.t95 2216.67
R1488 VDDA.t24 VDDA.t142 2126.19
R1489 VDDA.t116 VDDA.t201 1538.1
R1490 VDDA.t146 VDDA.t10 1492.86
R1491 VDDA.t8 VDDA.t120 1492.86
R1492 VDDA.t48 VDDA.t2 1317.78
R1493 VDDA.t85 VDDA.n91 1289.29
R1494 VDDA.t12 VDDA.n90 1289.29
R1495 VDDA.t33 VDDA.t112 1130.95
R1496 VDDA.t126 VDDA.t207 1130.95
R1497 VDDA.t65 VDDA.t38 1130.95
R1498 VDDA.t75 VDDA.t73 1130.95
R1499 VDDA.t93 VDDA.t114 1130.95
R1500 VDDA.t6 VDDA.n97 927.381
R1501 VDDA.t22 VDDA.n95 927.381
R1502 VDDA.t56 VDDA.n94 927.381
R1503 VDDA.t130 VDDA.n92 927.381
R1504 VDDA.n86 VDDA.n75 831.25
R1505 VDDA.n80 VDDA.n78 831.25
R1506 VDDA.n768 VDDA.n760 831.25
R1507 VDDA.n763 VDDA.n762 831.25
R1508 VDDA.n757 VDDA.n749 831.25
R1509 VDDA.n752 VDDA.n751 831.25
R1510 VDDA.n236 VDDA.t143 726.734
R1511 VDDA.n238 VDDA.t94 726.734
R1512 VDDA.n96 VDDA.t211 663.801
R1513 VDDA.n53 VDDA.t41 663.801
R1514 VDDA.n93 VDDA.t198 663.801
R1515 VDDA.n35 VDDA.t195 663.801
R1516 VDDA.n17 VDDA.t137 663.801
R1517 VDDA.n89 VDDA.t82 663.801
R1518 VDDA.n67 VDDA.n66 647.933
R1519 VDDA.n134 VDDA.n133 647.933
R1520 VDDA.n152 VDDA.n59 647.933
R1521 VDDA.n158 VDDA.n56 647.933
R1522 VDDA.n49 VDDA.n48 647.933
R1523 VDDA.n179 VDDA.n178 647.933
R1524 VDDA.n197 VDDA.n41 647.933
R1525 VDDA.n203 VDDA.n38 647.933
R1526 VDDA.n219 VDDA.n218 647.933
R1527 VDDA.n29 VDDA.n28 647.933
R1528 VDDA.n245 VDDA.n23 647.933
R1529 VDDA.n252 VDDA.n20 647.933
R1530 VDDA.n8 VDDA.n7 647.933
R1531 VDDA.n291 VDDA.n290 647.933
R1532 VDDA.n271 VDDA.n12 646.715
R1533 VDDA.n97 VDDA.t210 610.715
R1534 VDDA.n95 VDDA.t40 610.715
R1535 VDDA.n94 VDDA.t197 610.715
R1536 VDDA.n92 VDDA.t194 610.715
R1537 VDDA.n91 VDDA.t136 610.715
R1538 VDDA.n90 VDDA.t81 610.715
R1539 VDDA.n83 VDDA.n75 585
R1540 VDDA.n82 VDDA.n78 585
R1541 VDDA.n761 VDDA.n760 585
R1542 VDDA.n765 VDDA.n763 585
R1543 VDDA.n661 VDDA.n655 585
R1544 VDDA.n656 VDDA.n655 585
R1545 VDDA.n667 VDDA.n344 585
R1546 VDDA.n671 VDDA.n344 585
R1547 VDDA.n612 VDDA.n350 585
R1548 VDDA.n607 VDDA.n350 585
R1549 VDDA.n588 VDDA.n583 585
R1550 VDDA.n592 VDDA.n583 585
R1551 VDDA.n750 VDDA.n749 585
R1552 VDDA.n754 VDDA.n752 585
R1553 VDDA.n652 VDDA.n646 585
R1554 VDDA.n647 VDDA.n646 585
R1555 VDDA.n358 VDDA.n351 585
R1556 VDDA.n353 VDDA.n351 585
R1557 VDDA.n423 VDDA.n416 585
R1558 VDDA.n405 VDDA.n397 585
R1559 VDDA.n571 VDDA.n475 585
R1560 VDDA.n564 VDDA.n475 585
R1561 VDDA.n561 VDDA.n560 585
R1562 VDDA.n560 VDDA.n559 585
R1563 VDDA.n530 VDDA.n529 585
R1564 VDDA.n530 VDDA.n519 585
R1565 VDDA.n99 VDDA.t224 537.492
R1566 VDDA.n110 VDDA.t223 537.491
R1567 VDDA.n87 VDDA.t222 537.491
R1568 VDDA.t2 VDDA.t33 497.62
R1569 VDDA.t112 VDDA.t6 497.62
R1570 VDDA.t0 VDDA.t126 497.62
R1571 VDDA.t207 VDDA.t22 497.62
R1572 VDDA.t54 VDDA.t65 497.62
R1573 VDDA.t38 VDDA.t56 497.62
R1574 VDDA.t95 VDDA.t75 497.62
R1575 VDDA.t73 VDDA.t130 497.62
R1576 VDDA.t199 VDDA.t146 497.62
R1577 VDDA.t10 VDDA.t24 497.62
R1578 VDDA.t142 VDDA.t93 497.62
R1579 VDDA.t114 VDDA.t116 497.62
R1580 VDDA.t201 VDDA.t85 497.62
R1581 VDDA.t58 VDDA.t31 497.62
R1582 VDDA.t31 VDDA.t8 497.62
R1583 VDDA.t120 VDDA.t14 497.62
R1584 VDDA.t44 VDDA.t12 497.62
R1585 VDDA.t37 VDDA.n76 465.079
R1586 VDDA.n81 VDDA.t37 465.079
R1587 VDDA.n767 VDDA.t214 465.079
R1588 VDDA.t214 VDDA.n766 465.079
R1589 VDDA.n756 VDDA.t134 465.079
R1590 VDDA.t134 VDDA.n755 465.079
R1591 VDDA.n105 VDDA.t145 464.281
R1592 VDDA.n102 VDDA.t145 464.281
R1593 VDDA.n113 VDDA.t100 464.281
R1594 VDDA.t100 VDDA.n72 464.281
R1595 VDDA.t84 VDDA.n636 464.281
R1596 VDDA.n638 VDDA.t84 464.281
R1597 VDDA.n744 VDDA.t132 464.281
R1598 VDDA.t132 VDDA.n743 464.281
R1599 VDDA.n781 VDDA.t106 464.281
R1600 VDDA.t106 VDDA.n780 464.281
R1601 VDDA.n725 VDDA.t43 464.281
R1602 VDDA.t43 VDDA.n724 464.281
R1603 VDDA.n703 VDDA.t206 464.281
R1604 VDDA.t206 VDDA.n702 464.281
R1605 VDDA.n633 VDDA.t64 464.281
R1606 VDDA.t64 VDDA.n632 464.281
R1607 VDDA.t111 VDDA.n733 464.281
R1608 VDDA.n734 VDDA.t111 464.281
R1609 VDDA.t5 VDDA.n317 464.281
R1610 VDDA.n771 VDDA.t5 464.281
R1611 VDDA.t28 VDDA.n325 464.281
R1612 VDDA.n706 VDDA.t28 464.281
R1613 VDDA.t213 VDDA.n621 464.281
R1614 VDDA.n622 VDDA.t213 464.281
R1615 VDDA.n341 VDDA.t221 415.336
R1616 VDDA.n386 VDDA.t175 384.967
R1617 VDDA.n428 VDDA.t181 384.967
R1618 VDDA.n391 VDDA.t160 384.967
R1619 VDDA.n411 VDDA.t157 384.967
R1620 VDDA.n95 VDDA.n53 382.8
R1621 VDDA.n94 VDDA.n93 382.8
R1622 VDDA.n92 VDDA.n35 382.8
R1623 VDDA.n91 VDDA.n17 382.8
R1624 VDDA.n90 VDDA.n89 382.8
R1625 VDDA.n97 VDDA.n96 382.8
R1626 VDDA.n423 VDDA.t168 374.878
R1627 VDDA.t179 VDDA.t87 360.346
R1628 VDDA.t87 VDDA.t60 360.346
R1629 VDDA.t60 VDDA.t203 360.346
R1630 VDDA.t203 VDDA.t77 360.346
R1631 VDDA.t77 VDDA.t172 360.346
R1632 VDDA.t217 VDDA.t186 360.346
R1633 VDDA.t89 VDDA.t217 360.346
R1634 VDDA.t91 VDDA.t89 360.346
R1635 VDDA.t118 VDDA.t91 360.346
R1636 VDDA.t189 VDDA.t118 360.346
R1637 VDDA.n110 VDDA.t152 359.752
R1638 VDDA.n87 VDDA.t151 359.752
R1639 VDDA.n99 VDDA.t150 359.752
R1640 VDDA.n396 VDDA.t164 352.834
R1641 VDDA.n525 VDDA.t179 343.966
R1642 VDDA.n563 VDDA.t172 343.966
R1643 VDDA.t186 VDDA.n563 343.966
R1644 VDDA.n569 VDDA.t189 343.966
R1645 VDDA.n412 VDDA.t159 341.752
R1646 VDDA.n427 VDDA.t184 341.752
R1647 VDDA.n387 VDDA.t177 341.752
R1648 VDDA.n392 VDDA.t163 341.752
R1649 VDDA.n558 VDDA.t185 336.329
R1650 VDDA.n558 VDDA.t171 336.329
R1651 VDDA.n520 VDDA.t178 320.7
R1652 VDDA.n572 VDDA.t188 320.7
R1653 VDDA.n385 VDDA.n383 315.647
R1654 VDDA.n379 VDDA.n378 315.647
R1655 VDDA.n410 VDDA.n409 315.647
R1656 VDDA.n390 VDDA.n389 315.647
R1657 VDDA.n430 VDDA.n382 315.647
R1658 VDDA.n429 VDDA.n384 315.647
R1659 VDDA.n324 VDDA.t125 315.25
R1660 VDDA.t35 VDDA.t9 314.113
R1661 VDDA.t128 VDDA.t26 314.113
R1662 VDDA.t176 VDDA.n387 304.659
R1663 VDDA.n560 VDDA.n483 291.363
R1664 VDDA.n556 VDDA.n481 291.363
R1665 VDDA.n557 VDDA.n556 291.363
R1666 VDDA.n659 VDDA.n655 290.733
R1667 VDDA.n665 VDDA.n344 290.733
R1668 VDDA.n610 VDDA.n350 290.733
R1669 VDDA.n586 VDDA.n583 290.733
R1670 VDDA.n650 VDDA.n646 290.733
R1671 VDDA.n352 VDDA.n351 290.733
R1672 VDDA.n421 VDDA.n416 290.733
R1673 VDDA.n417 VDDA.n416 290.733
R1674 VDDA.n403 VDDA.n397 290.733
R1675 VDDA.n398 VDDA.n397 290.733
R1676 VDDA.n565 VDDA.n475 290.733
R1677 VDDA.n530 VDDA.n518 290.733
R1678 VDDA.n745 VDDA.n744 243.698
R1679 VDDA.n782 VDDA.n781 243.698
R1680 VDDA.n726 VDDA.n725 243.698
R1681 VDDA.n704 VDDA.n703 243.698
R1682 VDDA.n634 VDDA.n633 243.698
R1683 VDDA.n734 VDDA.n731 243.698
R1684 VDDA.n775 VDDA.n771 243.698
R1685 VDDA.n710 VDDA.n706 243.698
R1686 VDDA.n622 VDDA.n619 243.698
R1687 VDDA.n107 VDDA.n106 238.367
R1688 VDDA.n101 VDDA.n88 238.367
R1689 VDDA.n115 VDDA.n114 238.367
R1690 VDDA.n118 VDDA.n117 238.367
R1691 VDDA.n86 VDDA.n85 238.367
R1692 VDDA.n80 VDDA.n79 238.367
R1693 VDDA.n730 VDDA.n301 238.367
R1694 VDDA.n769 VDDA.n768 238.367
R1695 VDDA.n762 VDDA.n729 238.367
R1696 VDDA.n728 VDDA.n316 238.367
R1697 VDDA.n721 VDDA.n319 238.367
R1698 VDDA.n699 VDDA.n327 238.367
R1699 VDDA.n618 VDDA.n335 238.367
R1700 VDDA.n738 VDDA.n302 238.367
R1701 VDDA.n758 VDDA.n757 238.367
R1702 VDDA.n785 VDDA.n784 238.367
R1703 VDDA.n713 VDDA.n712 238.367
R1704 VDDA.n626 VDDA.n331 238.367
R1705 VDDA.n751 VDDA.n747 238.367
R1706 VDDA.n417 VDDA.n388 233.841
R1707 VDDA.n398 VDDA.n394 233.841
R1708 VDDA.n662 VDDA.n661 230.308
R1709 VDDA.n656 VDDA.n615 230.308
R1710 VDDA.n668 VDDA.n667 230.308
R1711 VDDA.n671 VDDA.n670 230.308
R1712 VDDA.n613 VDDA.n612 230.308
R1713 VDDA.n607 VDDA.n346 230.308
R1714 VDDA.n589 VDDA.n588 230.308
R1715 VDDA.n592 VDDA.n591 230.308
R1716 VDDA.n653 VDDA.n652 230.308
R1717 VDDA.n358 VDDA.n348 230.308
R1718 VDDA.n353 VDDA.n347 230.308
R1719 VDDA.n647 VDDA.n644 230.308
R1720 VDDA.n424 VDDA.n423 230.308
R1721 VDDA.n571 VDDA.n570 230.308
R1722 VDDA.n568 VDDA.n564 230.308
R1723 VDDA.n562 VDDA.n561 230.308
R1724 VDDA.n559 VDDA.n478 230.308
R1725 VDDA.t107 VDDA.t192 222.178
R1726 VDDA.n74 VDDA.t36 219.232
R1727 VDDA.t219 VDDA.n74 219.232
R1728 VDDA.n116 VDDA.t99 219.232
R1729 VDDA.n108 VDDA.t144 219.232
R1730 VDDA.n663 VDDA.n643 199.195
R1731 VDDA.n492 VDDA.n491 196.502
R1732 VDDA.n489 VDDA.n488 196.502
R1733 VDDA.n555 VDDA.n554 196.502
R1734 VDDA.n546 VDDA.n511 196.502
R1735 VDDA.n539 VDDA.n514 196.502
R1736 VDDA.n532 VDDA.n531 196.502
R1737 VDDA.n638 VDDA.n617 190.333
R1738 VDDA.n110 VDDA.t99 185.002
R1739 VDDA.t219 VDDA.n87 185.002
R1740 VDDA.n99 VDDA.t144 185.002
R1741 VDDA.n427 VDDA.n426 185.001
R1742 VDDA.n413 VDDA.n412 185.001
R1743 VDDA.n408 VDDA.n392 185.001
R1744 VDDA.n84 VDDA.n83 185
R1745 VDDA.n82 VDDA.n77 185
R1746 VDDA.n112 VDDA.n109 185
R1747 VDDA.n111 VDDA.n73 185
R1748 VDDA.n104 VDDA.n98 185
R1749 VDDA.n103 VDDA.n100 185
R1750 VDDA.n357 VDDA.n356 185
R1751 VDDA.n355 VDDA.n354 185
R1752 VDDA.n651 VDDA.n645 185
R1753 VDDA.n649 VDDA.n648 185
R1754 VDDA.n625 VDDA.n624 185
R1755 VDDA.n623 VDDA.n620 185
R1756 VDDA.n707 VDDA.n326 185
R1757 VDDA.n709 VDDA.n708 185
R1758 VDDA.n772 VDDA.n318 185
R1759 VDDA.n774 VDDA.n773 185
R1760 VDDA.n750 VDDA.n748 185
R1761 VDDA.n754 VDDA.n753 185
R1762 VDDA.n737 VDDA.n736 185
R1763 VDDA.n735 VDDA.n732 185
R1764 VDDA.n587 VDDA.n585 185
R1765 VDDA.n584 VDDA.n582 185
R1766 VDDA.n611 VDDA.n349 185
R1767 VDDA.n609 VDDA.n608 185
R1768 VDDA.n666 VDDA.n664 185
R1769 VDDA.n345 VDDA.n343 185
R1770 VDDA.n660 VDDA.n654 185
R1771 VDDA.n658 VDDA.n657 185
R1772 VDDA.n629 VDDA.n628 185
R1773 VDDA.n631 VDDA.n630 185
R1774 VDDA.n329 VDDA.n328 185
R1775 VDDA.n701 VDDA.n700 185
R1776 VDDA.n321 VDDA.n320 185
R1777 VDDA.n723 VDDA.n722 185
R1778 VDDA.n777 VDDA.n776 185
R1779 VDDA.n779 VDDA.n778 185
R1780 VDDA.n761 VDDA.n759 185
R1781 VDDA.n765 VDDA.n764 185
R1782 VDDA.n740 VDDA.n739 185
R1783 VDDA.n742 VDDA.n741 185
R1784 VDDA.n642 VDDA.n334 185
R1785 VDDA.n643 VDDA.n642 185
R1786 VDDA.n641 VDDA.n640 185
R1787 VDDA.n639 VDDA.n637 185
R1788 VDDA.n643 VDDA.n617 185
R1789 VDDA.n422 VDDA.n415 185
R1790 VDDA.n420 VDDA.n414 185
R1791 VDDA.n425 VDDA.n414 185
R1792 VDDA.n419 VDDA.n418 185
R1793 VDDA.n406 VDDA.n405 185
R1794 VDDA.n407 VDDA.n406 185
R1795 VDDA.n404 VDDA.n395 185
R1796 VDDA.n402 VDDA.n401 185
R1797 VDDA.n400 VDDA.n399 185
R1798 VDDA.n482 VDDA.n479 185
R1799 VDDA.n485 VDDA.n484 185
R1800 VDDA.n477 VDDA.n476 185
R1801 VDDA.n567 VDDA.n566 185
R1802 VDDA.n529 VDDA.n521 185
R1803 VDDA.n525 VDDA.n521 185
R1804 VDDA.n528 VDDA.n527 185
R1805 VDDA.n523 VDDA.n522 185
R1806 VDDA.n524 VDDA.n519 185
R1807 VDDA.n525 VDDA.n524 185
R1808 VDDA.n590 VDDA.t107 172.38
R1809 VDDA.t104 VDDA.n614 172.38
R1810 VDDA.n669 VDDA.t67 172.38
R1811 VDDA.n559 VDDA.n558 166.63
R1812 VDDA.n116 VDDA.t129 158.333
R1813 VDDA.t135 VDDA.n108 158.333
R1814 VDDA.n100 VDDA.n98 150
R1815 VDDA.n109 VDDA.n73 150
R1816 VDDA.n84 VDDA.n77 150
R1817 VDDA.n741 VDDA.n739 150
R1818 VDDA.n764 VDDA.n759 150
R1819 VDDA.n778 VDDA.n776 150
R1820 VDDA.n722 VDDA.n320 150
R1821 VDDA.n700 VDDA.n328 150
R1822 VDDA.n630 VDDA.n628 150
R1823 VDDA.n737 VDDA.n732 150
R1824 VDDA.n753 VDDA.n748 150
R1825 VDDA.n774 VDDA.n318 150
R1826 VDDA.n709 VDDA.n326 150
R1827 VDDA.n625 VDDA.n620 150
R1828 VDDA.n642 VDDA.n641 150
R1829 VDDA.n637 VDDA.n617 150
R1830 VDDA.t29 VDDA.t108 145.038
R1831 VDDA.n635 VDDA.n627 137.904
R1832 VDDA.n711 VDDA.n705 137.904
R1833 VDDA.n590 VDDA.t46 126.412
R1834 VDDA.n614 VDDA.t192 126.412
R1835 VDDA.n669 VDDA.t104 126.412
R1836 VDDA.t67 VDDA.n663 126.412
R1837 VDDA.t220 VDDA.n75 123.126
R1838 VDDA.n78 VDDA.t220 123.126
R1839 VDDA.t103 VDDA.n760 123.126
R1840 VDDA.n763 VDDA.t103 123.126
R1841 VDDA.t102 VDDA.n749 123.126
R1842 VDDA.n752 VDDA.t102 123.126
R1843 VDDA.n657 VDDA.n654 120.001
R1844 VDDA.n664 VDDA.n345 120.001
R1845 VDDA.n608 VDDA.n349 120.001
R1846 VDDA.n585 VDDA.n584 120.001
R1847 VDDA.n648 VDDA.n645 120.001
R1848 VDDA.n356 VDDA.n355 120.001
R1849 VDDA.n415 VDDA.n414 120.001
R1850 VDDA.n418 VDDA.n414 120.001
R1851 VDDA.n406 VDDA.n395 120.001
R1852 VDDA.n401 VDDA.n400 120.001
R1853 VDDA.n567 VDDA.n477 120.001
R1854 VDDA.n484 VDDA.n479 120.001
R1855 VDDA.n527 VDDA.n521 120.001
R1856 VDDA.n524 VDDA.n523 120.001
R1857 VDDA.n461 VDDA.n367 119.737
R1858 VDDA.n454 VDDA.n370 119.737
R1859 VDDA.n447 VDDA.n373 119.737
R1860 VDDA.n440 VDDA.n376 119.737
R1861 VDDA.n432 VDDA.n381 119.737
R1862 VDDA.n426 VDDA.t182 119.656
R1863 VDDA.t129 VDDA.t219 109.615
R1864 VDDA.t99 VDDA.t135 109.615
R1865 VDDA.t144 VDDA.t48 109.615
R1866 VDDA.n425 VDDA.n413 108.779
R1867 VDDA.n783 VDDA.n727 107.258
R1868 VDDA.n783 VDDA.t4 103.427
R1869 VDDA.t133 VDDA.n770 103.427
R1870 VDDA.n770 VDDA.t101 103.427
R1871 VDDA.t110 VDDA.n746 103.427
R1872 VDDA.n727 VDDA.t27 95.7666
R1873 VDDA.t16 VDDA.t176 94.2753
R1874 VDDA.t148 VDDA.t16 94.2753
R1875 VDDA.t69 VDDA.t148 94.2753
R1876 VDDA.t122 VDDA.t69 94.2753
R1877 VDDA.t182 VDDA.t122 94.2753
R1878 VDDA.t215 VDDA.t50 94.2753
R1879 VDDA.t52 VDDA.t161 94.2753
R1880 VDDA.t20 VDDA.n408 94.2753
R1881 VDDA.t156 VDDA.t62 94.2753
R1882 VDDA.t154 VDDA.t153 94.2753
R1883 VDDA.t63 VDDA.t83 91.936
R1884 VDDA.t205 VDDA.t212 91.936
R1885 VDDA.n87 VDDA.n86 90.5056
R1886 VDDA.t124 VDDA.t42 84.2747
R1887 VDDA.t4 VDDA.t35 84.2747
R1888 VDDA.t9 VDDA.t133 84.2747
R1889 VDDA.t101 VDDA.t128 84.2747
R1890 VDDA.t26 VDDA.t110 84.2747
R1891 VDDA.t169 VDDA.t158 83.3974
R1892 VDDA.t97 VDDA.t49 83.3974
R1893 VDDA.n410 VDDA.n379 83.2005
R1894 VDDA.n390 VDDA.n379 83.2005
R1895 VDDA.n430 VDDA.n383 83.2005
R1896 VDDA.n430 VDDA.n429 83.2005
R1897 VDDA.n66 VDDA.t3 78.8005
R1898 VDDA.n66 VDDA.t34 78.8005
R1899 VDDA.n133 VDDA.t113 78.8005
R1900 VDDA.n133 VDDA.t7 78.8005
R1901 VDDA.n59 VDDA.t1 78.8005
R1902 VDDA.n59 VDDA.t127 78.8005
R1903 VDDA.n56 VDDA.t208 78.8005
R1904 VDDA.n56 VDDA.t23 78.8005
R1905 VDDA.n48 VDDA.t55 78.8005
R1906 VDDA.n48 VDDA.t66 78.8005
R1907 VDDA.n178 VDDA.t39 78.8005
R1908 VDDA.n178 VDDA.t57 78.8005
R1909 VDDA.n41 VDDA.t96 78.8005
R1910 VDDA.n41 VDDA.t76 78.8005
R1911 VDDA.n38 VDDA.t74 78.8005
R1912 VDDA.n38 VDDA.t131 78.8005
R1913 VDDA.n218 VDDA.t200 78.8005
R1914 VDDA.n218 VDDA.t147 78.8005
R1915 VDDA.n28 VDDA.t11 78.8005
R1916 VDDA.n28 VDDA.t25 78.8005
R1917 VDDA.n23 VDDA.t115 78.8005
R1918 VDDA.n23 VDDA.t117 78.8005
R1919 VDDA.n20 VDDA.t202 78.8005
R1920 VDDA.n20 VDDA.t86 78.8005
R1921 VDDA.n12 VDDA.t59 78.8005
R1922 VDDA.n12 VDDA.t32 78.8005
R1923 VDDA.n7 VDDA.t121 78.8005
R1924 VDDA.n7 VDDA.t15 78.8005
R1925 VDDA.n290 VDDA.t45 78.8005
R1926 VDDA.n290 VDDA.t13 78.8005
R1927 VDDA.t18 VDDA.t79 76.1455
R1928 VDDA.t165 VDDA.t155 76.1455
R1929 VDDA.n114 VDDA.n110 74.7688
R1930 VDDA.n106 VDDA.n99 74.7688
R1931 VDDA.n614 VDDA.n348 69.8479
R1932 VDDA.n614 VDDA.n347 69.8479
R1933 VDDA.n663 VDDA.n653 69.8479
R1934 VDDA.n663 VDDA.n644 69.8479
R1935 VDDA.n590 VDDA.n589 69.8479
R1936 VDDA.n591 VDDA.n590 69.8479
R1937 VDDA.n614 VDDA.n613 69.8479
R1938 VDDA.n614 VDDA.n346 69.8479
R1939 VDDA.n669 VDDA.n668 69.8479
R1940 VDDA.n670 VDDA.n669 69.8479
R1941 VDDA.n663 VDDA.n662 69.8479
R1942 VDDA.n663 VDDA.n615 69.8479
R1943 VDDA.n425 VDDA.n424 69.8479
R1944 VDDA.n425 VDDA.n388 69.8479
R1945 VDDA.n407 VDDA.n393 69.8479
R1946 VDDA.n407 VDDA.n394 69.8479
R1947 VDDA.n563 VDDA.n562 69.8479
R1948 VDDA.n563 VDDA.n478 69.8479
R1949 VDDA.n570 VDDA.n569 69.8479
R1950 VDDA.n569 VDDA.n568 69.8479
R1951 VDDA.n526 VDDA.n525 69.8479
R1952 VDDA.n431 VDDA.n430 69.3203
R1953 VDDA.t79 VDDA.t140 68.8936
R1954 VDDA.t155 VDDA.n407 68.8936
R1955 VDDA.n85 VDDA.n74 65.8183
R1956 VDDA.n79 VDDA.n74 65.8183
R1957 VDDA.n116 VDDA.n115 65.8183
R1958 VDDA.n117 VDDA.n116 65.8183
R1959 VDDA.n108 VDDA.n107 65.8183
R1960 VDDA.n108 VDDA.n88 65.8183
R1961 VDDA.n627 VDDA.n626 65.8183
R1962 VDDA.n627 VDDA.n619 65.8183
R1963 VDDA.n712 VDDA.n711 65.8183
R1964 VDDA.n711 VDDA.n710 65.8183
R1965 VDDA.n784 VDDA.n783 65.8183
R1966 VDDA.n783 VDDA.n775 65.8183
R1967 VDDA.n770 VDDA.n758 65.8183
R1968 VDDA.n770 VDDA.n747 65.8183
R1969 VDDA.n746 VDDA.n738 65.8183
R1970 VDDA.n746 VDDA.n731 65.8183
R1971 VDDA.n635 VDDA.n634 65.8183
R1972 VDDA.n635 VDDA.n618 65.8183
R1973 VDDA.n705 VDDA.n704 65.8183
R1974 VDDA.n705 VDDA.n327 65.8183
R1975 VDDA.n727 VDDA.n726 65.8183
R1976 VDDA.n727 VDDA.n319 65.8183
R1977 VDDA.n783 VDDA.n782 65.8183
R1978 VDDA.n783 VDDA.n728 65.8183
R1979 VDDA.n770 VDDA.n769 65.8183
R1980 VDDA.n770 VDDA.n729 65.8183
R1981 VDDA.n746 VDDA.n745 65.8183
R1982 VDDA.n746 VDDA.n730 65.8183
R1983 VDDA.n643 VDDA.n616 65.8183
R1984 VDDA.t158 VDDA.t138 61.6417
R1985 VDDA.t49 VDDA.t71 61.6417
R1986 VDDA.n816 VDDA.n301 58.0576
R1987 VDDA.n786 VDDA.n316 58.0576
R1988 VDDA.n721 VDDA.n720 58.0576
R1989 VDDA.n699 VDDA.n698 58.0576
R1990 VDDA.n689 VDDA.n335 58.0576
R1991 VDDA.n816 VDDA.n302 58.0576
R1992 VDDA.n786 VDDA.n785 58.0576
R1993 VDDA.n714 VDDA.n713 58.0576
R1994 VDDA.n697 VDDA.n331 58.0576
R1995 VDDA.n690 VDDA.n334 58.0576
R1996 VDDA.n656 VDDA.n338 57.2449
R1997 VDDA.n672 VDDA.n671 57.2449
R1998 VDDA.n607 VDDA.n606 57.2449
R1999 VDDA.n593 VDDA.n592 57.2449
R2000 VDDA.n652 VDDA.n338 57.2449
R2001 VDDA.n606 VDDA.n358 57.2449
R2002 VDDA.n165 VDDA.n53 54.4005
R2003 VDDA.n93 VDDA.n44 54.4005
R2004 VDDA.n210 VDDA.n35 54.4005
R2005 VDDA.n259 VDDA.n17 54.4005
R2006 VDDA.n89 VDDA.n1 54.4005
R2007 VDDA.n96 VDDA.n62 54.4005
R2008 VDDA.n803 VDDA.n307 54.4005
R2009 VDDA.n309 VDDA.n307 54.4005
R2010 VDDA.n309 VDDA.n308 54.4005
R2011 VDDA.n803 VDDA.n308 54.4005
R2012 VDDA.n85 VDDA.n84 53.3664
R2013 VDDA.n79 VDDA.n77 53.3664
R2014 VDDA.n115 VDDA.n109 53.3664
R2015 VDDA.n117 VDDA.n73 53.3664
R2016 VDDA.n107 VDDA.n98 53.3664
R2017 VDDA.n100 VDDA.n88 53.3664
R2018 VDDA.n732 VDDA.n731 53.3664
R2019 VDDA.n753 VDDA.n747 53.3664
R2020 VDDA.n775 VDDA.n774 53.3664
R2021 VDDA.n626 VDDA.n625 53.3664
R2022 VDDA.n620 VDDA.n619 53.3664
R2023 VDDA.n712 VDDA.n326 53.3664
R2024 VDDA.n710 VDDA.n709 53.3664
R2025 VDDA.n784 VDDA.n318 53.3664
R2026 VDDA.n758 VDDA.n748 53.3664
R2027 VDDA.n738 VDDA.n737 53.3664
R2028 VDDA.n634 VDDA.n628 53.3664
R2029 VDDA.n630 VDDA.n618 53.3664
R2030 VDDA.n704 VDDA.n328 53.3664
R2031 VDDA.n700 VDDA.n327 53.3664
R2032 VDDA.n726 VDDA.n320 53.3664
R2033 VDDA.n722 VDDA.n319 53.3664
R2034 VDDA.n782 VDDA.n776 53.3664
R2035 VDDA.n778 VDDA.n728 53.3664
R2036 VDDA.n769 VDDA.n759 53.3664
R2037 VDDA.n764 VDDA.n729 53.3664
R2038 VDDA.n745 VDDA.n739 53.3664
R2039 VDDA.n741 VDDA.n730 53.3664
R2040 VDDA.n641 VDDA.n616 53.3664
R2041 VDDA.n637 VDDA.n616 53.3664
R2042 VDDA.n408 VDDA.t29 50.7639
R2043 VDDA.t177 VDDA.n385 49.2505
R2044 VDDA.n385 VDDA.t17 49.2505
R2045 VDDA.n378 VDDA.t51 49.2505
R2046 VDDA.n378 VDDA.t80 49.2505
R2047 VDDA.n409 VDDA.t159 49.2505
R2048 VDDA.n409 VDDA.t216 49.2505
R2049 VDDA.n389 VDDA.t53 49.2505
R2050 VDDA.n389 VDDA.t162 49.2505
R2051 VDDA.n382 VDDA.t149 49.2505
R2052 VDDA.n382 VDDA.t70 49.2505
R2053 VDDA.n384 VDDA.t123 49.2505
R2054 VDDA.n384 VDDA.t183 49.2505
R2055 VDDA.n818 VDDA.n817 47.7005
R2056 VDDA.n648 VDDA.n644 45.3071
R2057 VDDA.n355 VDDA.n347 45.3071
R2058 VDDA.n356 VDDA.n348 45.3071
R2059 VDDA.n653 VDDA.n645 45.3071
R2060 VDDA.n589 VDDA.n585 45.3071
R2061 VDDA.n591 VDDA.n584 45.3071
R2062 VDDA.n613 VDDA.n349 45.3071
R2063 VDDA.n608 VDDA.n346 45.3071
R2064 VDDA.n668 VDDA.n664 45.3071
R2065 VDDA.n670 VDDA.n345 45.3071
R2066 VDDA.n662 VDDA.n654 45.3071
R2067 VDDA.n657 VDDA.n615 45.3071
R2068 VDDA.n418 VDDA.n388 45.3071
R2069 VDDA.n424 VDDA.n415 45.3071
R2070 VDDA.n395 VDDA.n393 45.3071
R2071 VDDA.n400 VDDA.n394 45.3071
R2072 VDDA.n401 VDDA.n393 45.3071
R2073 VDDA.n562 VDDA.n479 45.3071
R2074 VDDA.n484 VDDA.n478 45.3071
R2075 VDDA.n570 VDDA.n477 45.3071
R2076 VDDA.n568 VDDA.n567 45.3071
R2077 VDDA.n527 VDDA.n526 45.3071
R2078 VDDA.n526 VDDA.n523 45.3071
R2079 VDDA.n437 VDDA.n379 41.6005
R2080 VDDA.t108 VDDA.t156 39.886
R2081 VDDA.n431 VDDA.n380 39.4988
R2082 VDDA.n579 VDDA.n578 38.1005
R2083 VDDA.n413 VDDA.t169 36.26
R2084 VDDA.t138 VDDA.t215 32.6341
R2085 VDDA.t71 VDDA.t154 32.6341
R2086 VDDA.n561 VDDA.n480 32.2291
R2087 VDDA.n120 VDDA.n70 32.0005
R2088 VDDA.n124 VDDA.n70 32.0005
R2089 VDDA.n125 VDDA.n124 32.0005
R2090 VDDA.n126 VDDA.n125 32.0005
R2091 VDDA.n132 VDDA.n131 32.0005
R2092 VDDA.n135 VDDA.n132 32.0005
R2093 VDDA.n139 VDDA.n64 32.0005
R2094 VDDA.n140 VDDA.n139 32.0005
R2095 VDDA.n141 VDDA.n140 32.0005
R2096 VDDA.n145 VDDA.n144 32.0005
R2097 VDDA.n146 VDDA.n145 32.0005
R2098 VDDA.n146 VDDA.n60 32.0005
R2099 VDDA.n150 VDDA.n60 32.0005
R2100 VDDA.n151 VDDA.n150 32.0005
R2101 VDDA.n153 VDDA.n57 32.0005
R2102 VDDA.n157 VDDA.n57 32.0005
R2103 VDDA.n160 VDDA.n159 32.0005
R2104 VDDA.n160 VDDA.n54 32.0005
R2105 VDDA.n164 VDDA.n54 32.0005
R2106 VDDA.n167 VDDA.n166 32.0005
R2107 VDDA.n167 VDDA.n51 32.0005
R2108 VDDA.n171 VDDA.n51 32.0005
R2109 VDDA.n172 VDDA.n171 32.0005
R2110 VDDA.n173 VDDA.n172 32.0005
R2111 VDDA.n177 VDDA.n176 32.0005
R2112 VDDA.n180 VDDA.n177 32.0005
R2113 VDDA.n184 VDDA.n46 32.0005
R2114 VDDA.n185 VDDA.n184 32.0005
R2115 VDDA.n186 VDDA.n185 32.0005
R2116 VDDA.n190 VDDA.n189 32.0005
R2117 VDDA.n191 VDDA.n190 32.0005
R2118 VDDA.n191 VDDA.n42 32.0005
R2119 VDDA.n195 VDDA.n42 32.0005
R2120 VDDA.n196 VDDA.n195 32.0005
R2121 VDDA.n198 VDDA.n39 32.0005
R2122 VDDA.n202 VDDA.n39 32.0005
R2123 VDDA.n205 VDDA.n204 32.0005
R2124 VDDA.n205 VDDA.n36 32.0005
R2125 VDDA.n209 VDDA.n36 32.0005
R2126 VDDA.n212 VDDA.n211 32.0005
R2127 VDDA.n212 VDDA.n33 32.0005
R2128 VDDA.n216 VDDA.n33 32.0005
R2129 VDDA.n217 VDDA.n216 32.0005
R2130 VDDA.n220 VDDA.n217 32.0005
R2131 VDDA.n224 VDDA.n31 32.0005
R2132 VDDA.n225 VDDA.n224 32.0005
R2133 VDDA.n226 VDDA.n225 32.0005
R2134 VDDA.n230 VDDA.n229 32.0005
R2135 VDDA.n231 VDDA.n230 32.0005
R2136 VDDA.n231 VDDA.n26 32.0005
R2137 VDDA.n235 VDDA.n26 32.0005
R2138 VDDA.n239 VDDA.n237 32.0005
R2139 VDDA.n243 VDDA.n24 32.0005
R2140 VDDA.n244 VDDA.n243 32.0005
R2141 VDDA.n246 VDDA.n21 32.0005
R2142 VDDA.n250 VDDA.n21 32.0005
R2143 VDDA.n251 VDDA.n250 32.0005
R2144 VDDA.n253 VDDA.n18 32.0005
R2145 VDDA.n257 VDDA.n18 32.0005
R2146 VDDA.n258 VDDA.n257 32.0005
R2147 VDDA.n260 VDDA.n15 32.0005
R2148 VDDA.n264 VDDA.n15 32.0005
R2149 VDDA.n265 VDDA.n264 32.0005
R2150 VDDA.n266 VDDA.n265 32.0005
R2151 VDDA.n266 VDDA.n13 32.0005
R2152 VDDA.n270 VDDA.n13 32.0005
R2153 VDDA.n273 VDDA.n272 32.0005
R2154 VDDA.n273 VDDA.n10 32.0005
R2155 VDDA.n277 VDDA.n10 32.0005
R2156 VDDA.n278 VDDA.n277 32.0005
R2157 VDDA.n279 VDDA.n278 32.0005
R2158 VDDA.n283 VDDA.n282 32.0005
R2159 VDDA.n284 VDDA.n283 32.0005
R2160 VDDA.n284 VDDA.n5 32.0005
R2161 VDDA.n288 VDDA.n5 32.0005
R2162 VDDA.n289 VDDA.n288 32.0005
R2163 VDDA.n292 VDDA.n289 32.0005
R2164 VDDA.n296 VDDA.n3 32.0005
R2165 VDDA.n297 VDDA.n296 32.0005
R2166 VDDA.n298 VDDA.n297 32.0005
R2167 VDDA.n594 VDDA.n362 32.0005
R2168 VDDA.n598 VDDA.n362 32.0005
R2169 VDDA.n599 VDDA.n598 32.0005
R2170 VDDA.n600 VDDA.n599 32.0005
R2171 VDDA.n600 VDDA.n359 32.0005
R2172 VDDA.n606 VDDA.n359 32.0005
R2173 VDDA.n606 VDDA.n360 32.0005
R2174 VDDA.n360 VDDA.n342 32.0005
R2175 VDDA.n673 VDDA.n342 32.0005
R2176 VDDA.n677 VDDA.n340 32.0005
R2177 VDDA.n678 VDDA.n677 32.0005
R2178 VDDA.n679 VDDA.n678 32.0005
R2179 VDDA.n683 VDDA.n682 32.0005
R2180 VDDA.n684 VDDA.n683 32.0005
R2181 VDDA.n684 VDDA.n336 32.0005
R2182 VDDA.n688 VDDA.n336 32.0005
R2183 VDDA.n692 VDDA.n691 32.0005
R2184 VDDA.n692 VDDA.n330 32.0005
R2185 VDDA.n696 VDDA.n332 32.0005
R2186 VDDA.n719 VDDA.n322 32.0005
R2187 VDDA.n787 VDDA.n315 32.0005
R2188 VDDA.n791 VDDA.n313 32.0005
R2189 VDDA.n792 VDDA.n791 32.0005
R2190 VDDA.n793 VDDA.n792 32.0005
R2191 VDDA.n793 VDDA.n311 32.0005
R2192 VDDA.n797 VDDA.n311 32.0005
R2193 VDDA.n798 VDDA.n797 32.0005
R2194 VDDA.n799 VDDA.n798 32.0005
R2195 VDDA.n805 VDDA.n804 32.0005
R2196 VDDA.n805 VDDA.n305 32.0005
R2197 VDDA.n809 VDDA.n305 32.0005
R2198 VDDA.n810 VDDA.n809 32.0005
R2199 VDDA.n811 VDDA.n810 32.0005
R2200 VDDA.n811 VDDA.n303 32.0005
R2201 VDDA.n815 VDDA.n303 32.0005
R2202 VDDA.n435 VDDA.n380 32.0005
R2203 VDDA.n436 VDDA.n435 32.0005
R2204 VDDA.n438 VDDA.n375 32.0005
R2205 VDDA.n443 VDDA.n375 32.0005
R2206 VDDA.n444 VDDA.n443 32.0005
R2207 VDDA.n445 VDDA.n444 32.0005
R2208 VDDA.n445 VDDA.n372 32.0005
R2209 VDDA.n450 VDDA.n372 32.0005
R2210 VDDA.n451 VDDA.n450 32.0005
R2211 VDDA.n452 VDDA.n451 32.0005
R2212 VDDA.n452 VDDA.n369 32.0005
R2213 VDDA.n457 VDDA.n369 32.0005
R2214 VDDA.n458 VDDA.n457 32.0005
R2215 VDDA.n459 VDDA.n458 32.0005
R2216 VDDA.n459 VDDA.n366 32.0005
R2217 VDDA.n464 VDDA.n366 32.0005
R2218 VDDA.n465 VDDA.n464 32.0005
R2219 VDDA.n465 VDDA.n364 32.0005
R2220 VDDA.n469 VDDA.n364 32.0005
R2221 VDDA.n470 VDDA.n469 32.0005
R2222 VDDA.n574 VDDA.n472 32.0005
R2223 VDDA.n578 VDDA.n472 32.0005
R2224 VDDA.n498 VDDA.n497 32.0005
R2225 VDDA.n497 VDDA.n496 32.0005
R2226 VDDA.n504 VDDA.n486 32.0005
R2227 VDDA.n504 VDDA.n503 32.0005
R2228 VDDA.n503 VDDA.n502 32.0005
R2229 VDDA.n553 VDDA.n508 32.0005
R2230 VDDA.n548 VDDA.n547 32.0005
R2231 VDDA.n541 VDDA.n540 32.0005
R2232 VDDA.n541 VDDA.n512 32.0005
R2233 VDDA.n545 VDDA.n512 32.0005
R2234 VDDA.n534 VDDA.n533 32.0005
R2235 VDDA.n534 VDDA.n515 32.0005
R2236 VDDA.n538 VDDA.n515 32.0005
R2237 VDDA.n428 VDDA.n427 30.754
R2238 VDDA.n392 VDDA.n391 30.754
R2239 VDDA.n80 VDDA.n71 30.2632
R2240 VDDA.n412 VDDA.n411 30.186
R2241 VDDA.n387 VDDA.n386 30.186
R2242 VDDA.n131 VDDA.n67 28.8005
R2243 VDDA.n144 VDDA.n62 28.8005
R2244 VDDA.n153 VDDA.n152 28.8005
R2245 VDDA.n166 VDDA.n165 28.8005
R2246 VDDA.n176 VDDA.n49 28.8005
R2247 VDDA.n189 VDDA.n44 28.8005
R2248 VDDA.n198 VDDA.n197 28.8005
R2249 VDDA.n211 VDDA.n210 28.8005
R2250 VDDA.n246 VDDA.n245 28.8005
R2251 VDDA.n271 VDDA.n270 28.8005
R2252 VDDA.n673 VDDA.n672 28.8005
R2253 VDDA.n573 VDDA.n474 28.8005
R2254 VDDA.n498 VDDA.n489 28.8005
R2255 VDDA.n554 VDDA.n553 28.8005
R2256 VDDA.n259 VDDA.n258 25.6005
R2257 VDDA.n594 VDDA.n593 25.6005
R2258 VDDA.n679 VDDA.n338 25.6005
R2259 VDDA.n691 VDDA.n690 25.6005
R2260 VDDA.n715 VDDA.n714 25.6005
R2261 VDDA.n720 VDDA.n315 25.6005
R2262 VDDA.n787 VDDA.n786 25.6005
R2263 VDDA.n802 VDDA.n309 25.6005
R2264 VDDA.n803 VDDA.n802 25.6005
R2265 VDDA.n817 VDDA.n816 25.6005
R2266 VDDA.n437 VDDA.n436 25.6005
R2267 VDDA VDDA.n470 25.6005
R2268 VDDA.t140 VDDA.t52 25.3822
R2269 VDDA.t161 VDDA.t20 25.3822
R2270 VDDA.n119 VDDA.n118 24.991
R2271 VDDA.n101 VDDA.n68 24.991
R2272 VDDA.n818 VDDA.n300 24.8806
R2273 VDDA.n655 VDDA.t68 24.6255
R2274 VDDA.n344 VDDA.t105 24.6255
R2275 VDDA.n350 VDDA.t196 24.6255
R2276 VDDA.n583 VDDA.t47 24.6255
R2277 VDDA.n646 VDDA.t209 24.6255
R2278 VDDA.n351 VDDA.t193 24.6255
R2279 VDDA.n491 VDDA.t119 24.6255
R2280 VDDA.n491 VDDA.t190 24.6255
R2281 VDDA.n488 VDDA.t90 24.6255
R2282 VDDA.n488 VDDA.t92 24.6255
R2283 VDDA.t187 VDDA.n555 24.6255
R2284 VDDA.n555 VDDA.t218 24.6255
R2285 VDDA.n511 VDDA.t78 24.6255
R2286 VDDA.n511 VDDA.t173 24.6255
R2287 VDDA.n514 VDDA.t61 24.6255
R2288 VDDA.n514 VDDA.t204 24.6255
R2289 VDDA.n531 VDDA.t180 24.6255
R2290 VDDA.n531 VDDA.t88 24.6255
R2291 VDDA.t180 VDDA.n530 24.6255
R2292 VDDA.n475 VDDA.t191 24.6255
R2293 VDDA.n556 VDDA.t187 24.6255
R2294 VDDA.n560 VDDA.t174 24.6255
R2295 VDDA.n520 VDDA.n517 24.361
R2296 VDDA.n129 VDDA.n128 24.1919
R2297 VDDA.n300 VDDA.n1 23.4989
R2298 VDDA.n120 VDDA.n119 22.4005
R2299 VDDA.n126 VDDA.n68 22.4005
R2300 VDDA.n135 VDDA.n134 22.4005
R2301 VDDA.n158 VDDA.n157 22.4005
R2302 VDDA.n180 VDDA.n179 22.4005
R2303 VDDA.n203 VDDA.n202 22.4005
R2304 VDDA.n219 VDDA.n31 22.4005
R2305 VDDA.n226 VDDA.n29 22.4005
R2306 VDDA.n291 VDDA.n3 22.4005
R2307 VDDA.n496 VDDA.n492 22.4005
R2308 VDDA.n547 VDDA.n546 22.4005
R2309 VDDA.n548 VDDA.n480 22.4005
R2310 VDDA.n405 VDDA.n396 22.0449
R2311 VDDA.n416 VDDA.t170 19.7005
R2312 VDDA.n397 VDDA.t167 19.7005
R2313 VDDA.n367 VDDA.t72 19.7005
R2314 VDDA.n367 VDDA.t166 19.7005
R2315 VDDA.n370 VDDA.t109 19.7005
R2316 VDDA.n370 VDDA.t98 19.7005
R2317 VDDA.n373 VDDA.t21 19.7005
R2318 VDDA.n373 VDDA.t30 19.7005
R2319 VDDA.n376 VDDA.t19 19.7005
R2320 VDDA.n376 VDDA.t141 19.7005
R2321 VDDA.t170 VDDA.n381 19.7005
R2322 VDDA.n381 VDDA.t139 19.7005
R2323 VDDA.n237 VDDA.n236 19.2005
R2324 VDDA.n239 VDDA.n238 19.2005
R2325 VDDA.n279 VDDA.n8 19.2005
R2326 VDDA.n332 VDDA.n324 19.2005
R2327 VDDA.t50 VDDA.t18 18.1303
R2328 VDDA.t153 VDDA.t165 18.1303
R2329 VDDA.n573 VDDA.n572 17.6005
R2330 VDDA.n252 VDDA.n251 16.0005
R2331 VDDA.n253 VDDA.n252 16.0005
R2332 VDDA.n298 VDDA.n1 16.0005
R2333 VDDA.n697 VDDA.n696 16.0005
R2334 VDDA.n429 VDDA.n428 16.0005
R2335 VDDA.n391 VDDA.n390 16.0005
R2336 VDDA.n411 VDDA.n410 16.0005
R2337 VDDA.n386 VDDA.n383 16.0005
R2338 VDDA.n492 VDDA.n474 16.0005
R2339 VDDA.n508 VDDA.n480 16.0005
R2340 VDDA.n546 VDDA.n545 16.0005
R2341 VDDA.n533 VDDA.n532 16.0005
R2342 VDDA.n471 VDDA 15.7005
R2343 VDDA.n572 VDDA.n571 15.6449
R2344 VDDA.n529 VDDA.n520 15.6449
R2345 VDDA.n593 VDDA.n581 13.8989
R2346 VDDA.n236 VDDA.n235 12.8005
R2347 VDDA.n238 VDDA.n24 12.8005
R2348 VDDA.n282 VDDA.n8 12.8005
R2349 VDDA.n698 VDDA.n330 12.8005
R2350 VDDA.n715 VDDA.n324 12.8005
R2351 VDDA.n580 VDDA.n471 12.7493
R2352 VDDA.n581 VDDA.n580 12.3383
R2353 VDDA.n580 VDDA.n579 11.579
R2354 VDDA.n643 VDDA.t63 11.4924
R2355 VDDA.t83 VDDA.n635 11.4924
R2356 VDDA.n627 VDDA.t205 11.4924
R2357 VDDA.n705 VDDA.t212 11.4924
R2358 VDDA.n711 VDDA.t124 11.4924
R2359 VDDA.t62 VDDA.t97 10.8784
R2360 VDDA.n129 VDDA.n67 10.7016
R2361 VDDA.n396 VDDA.n365 9.613
R2362 VDDA.n134 VDDA.n64 9.6005
R2363 VDDA.n159 VDDA.n158 9.6005
R2364 VDDA.n179 VDDA.n46 9.6005
R2365 VDDA.n204 VDDA.n203 9.6005
R2366 VDDA.n220 VDDA.n219 9.6005
R2367 VDDA.n229 VDDA.n29 9.6005
R2368 VDDA.n292 VDDA.n291 9.6005
R2369 VDDA.n574 VDDA.n573 9.6005
R2370 VDDA.n554 VDDA.n486 9.6005
R2371 VDDA.n502 VDDA.n489 9.6005
R2372 VDDA.n121 VDDA.n120 9.3005
R2373 VDDA.n122 VDDA.n70 9.3005
R2374 VDDA.n124 VDDA.n123 9.3005
R2375 VDDA.n125 VDDA.n69 9.3005
R2376 VDDA.n127 VDDA.n126 9.3005
R2377 VDDA.n131 VDDA.n130 9.3005
R2378 VDDA.n132 VDDA.n65 9.3005
R2379 VDDA.n136 VDDA.n135 9.3005
R2380 VDDA.n137 VDDA.n64 9.3005
R2381 VDDA.n139 VDDA.n138 9.3005
R2382 VDDA.n140 VDDA.n63 9.3005
R2383 VDDA.n142 VDDA.n141 9.3005
R2384 VDDA.n144 VDDA.n143 9.3005
R2385 VDDA.n145 VDDA.n61 9.3005
R2386 VDDA.n147 VDDA.n146 9.3005
R2387 VDDA.n148 VDDA.n60 9.3005
R2388 VDDA.n150 VDDA.n149 9.3005
R2389 VDDA.n151 VDDA.n58 9.3005
R2390 VDDA.n154 VDDA.n153 9.3005
R2391 VDDA.n155 VDDA.n57 9.3005
R2392 VDDA.n157 VDDA.n156 9.3005
R2393 VDDA.n159 VDDA.n55 9.3005
R2394 VDDA.n161 VDDA.n160 9.3005
R2395 VDDA.n162 VDDA.n54 9.3005
R2396 VDDA.n164 VDDA.n163 9.3005
R2397 VDDA.n166 VDDA.n52 9.3005
R2398 VDDA.n168 VDDA.n167 9.3005
R2399 VDDA.n169 VDDA.n51 9.3005
R2400 VDDA.n171 VDDA.n170 9.3005
R2401 VDDA.n172 VDDA.n50 9.3005
R2402 VDDA.n174 VDDA.n173 9.3005
R2403 VDDA.n176 VDDA.n175 9.3005
R2404 VDDA.n177 VDDA.n47 9.3005
R2405 VDDA.n181 VDDA.n180 9.3005
R2406 VDDA.n182 VDDA.n46 9.3005
R2407 VDDA.n184 VDDA.n183 9.3005
R2408 VDDA.n185 VDDA.n45 9.3005
R2409 VDDA.n187 VDDA.n186 9.3005
R2410 VDDA.n189 VDDA.n188 9.3005
R2411 VDDA.n190 VDDA.n43 9.3005
R2412 VDDA.n192 VDDA.n191 9.3005
R2413 VDDA.n193 VDDA.n42 9.3005
R2414 VDDA.n195 VDDA.n194 9.3005
R2415 VDDA.n196 VDDA.n40 9.3005
R2416 VDDA.n199 VDDA.n198 9.3005
R2417 VDDA.n200 VDDA.n39 9.3005
R2418 VDDA.n202 VDDA.n201 9.3005
R2419 VDDA.n204 VDDA.n37 9.3005
R2420 VDDA.n206 VDDA.n205 9.3005
R2421 VDDA.n207 VDDA.n36 9.3005
R2422 VDDA.n209 VDDA.n208 9.3005
R2423 VDDA.n211 VDDA.n34 9.3005
R2424 VDDA.n213 VDDA.n212 9.3005
R2425 VDDA.n214 VDDA.n33 9.3005
R2426 VDDA.n216 VDDA.n215 9.3005
R2427 VDDA.n217 VDDA.n32 9.3005
R2428 VDDA.n221 VDDA.n220 9.3005
R2429 VDDA.n222 VDDA.n31 9.3005
R2430 VDDA.n224 VDDA.n223 9.3005
R2431 VDDA.n225 VDDA.n30 9.3005
R2432 VDDA.n227 VDDA.n226 9.3005
R2433 VDDA.n229 VDDA.n228 9.3005
R2434 VDDA.n230 VDDA.n27 9.3005
R2435 VDDA.n232 VDDA.n231 9.3005
R2436 VDDA.n233 VDDA.n26 9.3005
R2437 VDDA.n235 VDDA.n234 9.3005
R2438 VDDA.n237 VDDA.n25 9.3005
R2439 VDDA.n240 VDDA.n239 9.3005
R2440 VDDA.n241 VDDA.n24 9.3005
R2441 VDDA.n243 VDDA.n242 9.3005
R2442 VDDA.n244 VDDA.n22 9.3005
R2443 VDDA.n247 VDDA.n246 9.3005
R2444 VDDA.n248 VDDA.n21 9.3005
R2445 VDDA.n250 VDDA.n249 9.3005
R2446 VDDA.n251 VDDA.n19 9.3005
R2447 VDDA.n254 VDDA.n253 9.3005
R2448 VDDA.n255 VDDA.n18 9.3005
R2449 VDDA.n257 VDDA.n256 9.3005
R2450 VDDA.n258 VDDA.n16 9.3005
R2451 VDDA.n261 VDDA.n260 9.3005
R2452 VDDA.n262 VDDA.n15 9.3005
R2453 VDDA.n264 VDDA.n263 9.3005
R2454 VDDA.n265 VDDA.n14 9.3005
R2455 VDDA.n267 VDDA.n266 9.3005
R2456 VDDA.n268 VDDA.n13 9.3005
R2457 VDDA.n270 VDDA.n269 9.3005
R2458 VDDA.n272 VDDA.n11 9.3005
R2459 VDDA.n274 VDDA.n273 9.3005
R2460 VDDA.n275 VDDA.n10 9.3005
R2461 VDDA.n277 VDDA.n276 9.3005
R2462 VDDA.n278 VDDA.n9 9.3005
R2463 VDDA.n280 VDDA.n279 9.3005
R2464 VDDA.n282 VDDA.n281 9.3005
R2465 VDDA.n283 VDDA.n6 9.3005
R2466 VDDA.n285 VDDA.n284 9.3005
R2467 VDDA.n286 VDDA.n5 9.3005
R2468 VDDA.n288 VDDA.n287 9.3005
R2469 VDDA.n289 VDDA.n4 9.3005
R2470 VDDA.n293 VDDA.n292 9.3005
R2471 VDDA.n294 VDDA.n3 9.3005
R2472 VDDA.n296 VDDA.n295 9.3005
R2473 VDDA.n297 VDDA.n2 9.3005
R2474 VDDA.n299 VDDA.n298 9.3005
R2475 VDDA.n470 VDDA.n363 9.3005
R2476 VDDA.n469 VDDA.n468 9.3005
R2477 VDDA.n467 VDDA.n364 9.3005
R2478 VDDA.n466 VDDA.n465 9.3005
R2479 VDDA.n464 VDDA.n463 9.3005
R2480 VDDA.n462 VDDA.n366 9.3005
R2481 VDDA.n460 VDDA.n459 9.3005
R2482 VDDA.n458 VDDA.n368 9.3005
R2483 VDDA.n457 VDDA.n456 9.3005
R2484 VDDA.n455 VDDA.n369 9.3005
R2485 VDDA.n453 VDDA.n452 9.3005
R2486 VDDA.n451 VDDA.n371 9.3005
R2487 VDDA.n450 VDDA.n449 9.3005
R2488 VDDA.n448 VDDA.n372 9.3005
R2489 VDDA.n446 VDDA.n445 9.3005
R2490 VDDA.n444 VDDA.n374 9.3005
R2491 VDDA.n443 VDDA.n442 9.3005
R2492 VDDA.n441 VDDA.n375 9.3005
R2493 VDDA.n439 VDDA.n438 9.3005
R2494 VDDA.n433 VDDA.n380 9.3005
R2495 VDDA.n435 VDDA.n434 9.3005
R2496 VDDA.n436 VDDA.n377 9.3005
R2497 VDDA.n533 VDDA.n516 9.3005
R2498 VDDA.n535 VDDA.n534 9.3005
R2499 VDDA.n536 VDDA.n515 9.3005
R2500 VDDA.n538 VDDA.n537 9.3005
R2501 VDDA.n540 VDDA.n513 9.3005
R2502 VDDA.n542 VDDA.n541 9.3005
R2503 VDDA.n543 VDDA.n512 9.3005
R2504 VDDA.n545 VDDA.n544 9.3005
R2505 VDDA.n546 VDDA.n510 9.3005
R2506 VDDA.n547 VDDA.n509 9.3005
R2507 VDDA.n549 VDDA.n548 9.3005
R2508 VDDA.n550 VDDA.n480 9.3005
R2509 VDDA.n551 VDDA.n508 9.3005
R2510 VDDA.n553 VDDA.n552 9.3005
R2511 VDDA.n554 VDDA.n507 9.3005
R2512 VDDA.n506 VDDA.n486 9.3005
R2513 VDDA.n505 VDDA.n504 9.3005
R2514 VDDA.n503 VDDA.n487 9.3005
R2515 VDDA.n502 VDDA.n501 9.3005
R2516 VDDA.n500 VDDA.n489 9.3005
R2517 VDDA.n499 VDDA.n498 9.3005
R2518 VDDA.n497 VDDA.n490 9.3005
R2519 VDDA.n496 VDDA.n495 9.3005
R2520 VDDA.n494 VDDA.n492 9.3005
R2521 VDDA.n493 VDDA.n474 9.3005
R2522 VDDA.n573 VDDA.n473 9.3005
R2523 VDDA.n575 VDDA.n574 9.3005
R2524 VDDA.n576 VDDA.n472 9.3005
R2525 VDDA.n578 VDDA.n577 9.3005
R2526 VDDA.n817 VDDA.n0 9.3005
R2527 VDDA.n595 VDDA.n594 9.3005
R2528 VDDA.n596 VDDA.n362 9.3005
R2529 VDDA.n598 VDDA.n597 9.3005
R2530 VDDA.n599 VDDA.n361 9.3005
R2531 VDDA.n601 VDDA.n600 9.3005
R2532 VDDA.n602 VDDA.n359 9.3005
R2533 VDDA.n606 VDDA.n605 9.3005
R2534 VDDA.n604 VDDA.n360 9.3005
R2535 VDDA.n603 VDDA.n342 9.3005
R2536 VDDA.n674 VDDA.n673 9.3005
R2537 VDDA.n675 VDDA.n340 9.3005
R2538 VDDA.n677 VDDA.n676 9.3005
R2539 VDDA.n678 VDDA.n339 9.3005
R2540 VDDA.n680 VDDA.n679 9.3005
R2541 VDDA.n682 VDDA.n681 9.3005
R2542 VDDA.n683 VDDA.n337 9.3005
R2543 VDDA.n685 VDDA.n684 9.3005
R2544 VDDA.n686 VDDA.n336 9.3005
R2545 VDDA.n688 VDDA.n687 9.3005
R2546 VDDA.n691 VDDA.n333 9.3005
R2547 VDDA.n693 VDDA.n692 9.3005
R2548 VDDA.n694 VDDA.n330 9.3005
R2549 VDDA.n696 VDDA.n695 9.3005
R2550 VDDA.n332 VDDA.n323 9.3005
R2551 VDDA.n716 VDDA.n715 9.3005
R2552 VDDA.n717 VDDA.n322 9.3005
R2553 VDDA.n719 VDDA.n718 9.3005
R2554 VDDA.n315 VDDA.n314 9.3005
R2555 VDDA.n788 VDDA.n787 9.3005
R2556 VDDA.n789 VDDA.n313 9.3005
R2557 VDDA.n791 VDDA.n790 9.3005
R2558 VDDA.n792 VDDA.n312 9.3005
R2559 VDDA.n794 VDDA.n793 9.3005
R2560 VDDA.n795 VDDA.n311 9.3005
R2561 VDDA.n797 VDDA.n796 9.3005
R2562 VDDA.n798 VDDA.n310 9.3005
R2563 VDDA.n800 VDDA.n799 9.3005
R2564 VDDA.n802 VDDA.n801 9.3005
R2565 VDDA.n804 VDDA.n306 9.3005
R2566 VDDA.n806 VDDA.n805 9.3005
R2567 VDDA.n807 VDDA.n305 9.3005
R2568 VDDA.n809 VDDA.n808 9.3005
R2569 VDDA.n810 VDDA.n304 9.3005
R2570 VDDA.n812 VDDA.n811 9.3005
R2571 VDDA.n813 VDDA.n303 9.3005
R2572 VDDA.n815 VDDA.n814 9.3005
R2573 VDDA.n112 VDDA.n111 9.14336
R2574 VDDA.n104 VDDA.n103 9.14336
R2575 VDDA.n742 VDDA.n740 9.14336
R2576 VDDA.n779 VDDA.n777 9.14336
R2577 VDDA.n723 VDDA.n321 9.14336
R2578 VDDA.n701 VDDA.n329 9.14336
R2579 VDDA.n631 VDDA.n629 9.14336
R2580 VDDA.n736 VDDA.n735 9.14336
R2581 VDDA.n773 VDDA.n772 9.14336
R2582 VDDA.n708 VDDA.n707 9.14336
R2583 VDDA.n624 VDDA.n623 9.14336
R2584 VDDA.n640 VDDA.n639 9.14336
R2585 VDDA.t42 VDDA.t27 7.66179
R2586 VDDA.n426 VDDA.n425 7.25241
R2587 VDDA.n661 VDDA.n660 7.11161
R2588 VDDA.n658 VDDA.n656 7.11161
R2589 VDDA.n667 VDDA.n666 7.11161
R2590 VDDA.n671 VDDA.n343 7.11161
R2591 VDDA.n612 VDDA.n611 7.11161
R2592 VDDA.n609 VDDA.n607 7.11161
R2593 VDDA.n588 VDDA.n587 7.11161
R2594 VDDA.n592 VDDA.n582 7.11161
R2595 VDDA.n652 VDDA.n651 7.11161
R2596 VDDA.n649 VDDA.n647 7.11161
R2597 VDDA.n358 VDDA.n357 7.11161
R2598 VDDA.n354 VDDA.n353 7.11161
R2599 VDDA.n423 VDDA.n422 7.11161
R2600 VDDA.n420 VDDA.n419 7.11161
R2601 VDDA.n405 VDDA.n404 7.11161
R2602 VDDA.n402 VDDA.n399 7.11161
R2603 VDDA.n571 VDDA.n476 7.11161
R2604 VDDA.n566 VDDA.n564 7.11161
R2605 VDDA.n529 VDDA.n528 7.11161
R2606 VDDA.n522 VDDA.n519 7.11161
R2607 VDDA.n128 VDDA.n68 7.05969
R2608 VDDA.n119 VDDA.n71 7.05957
R2609 VDDA.n532 VDDA.n517 6.54033
R2610 VDDA.n260 VDDA.n259 6.4005
R2611 VDDA.n682 VDDA.n338 6.4005
R2612 VDDA.n714 VDDA.n322 6.4005
R2613 VDDA.n720 VDDA.n719 6.4005
R2614 VDDA.n786 VDDA.n313 6.4005
R2615 VDDA.n799 VDDA.n309 6.4005
R2616 VDDA.n804 VDDA.n803 6.4005
R2617 VDDA.n816 VDDA.n815 6.4005
R2618 VDDA.n438 VDDA.n437 6.4005
R2619 VDDA.n83 VDDA.n82 5.81868
R2620 VDDA.n765 VDDA.n761 5.81868
R2621 VDDA.n754 VDDA.n750 5.81868
R2622 VDDA.n106 VDDA.n105 5.33286
R2623 VDDA.n114 VDDA.n113 5.33286
R2624 VDDA.n118 VDDA.n72 5.33286
R2625 VDDA.n102 VDDA.n101 5.33286
R2626 VDDA.n636 VDDA.n334 5.33286
R2627 VDDA.n743 VDDA.n301 5.33286
R2628 VDDA.n780 VDDA.n316 5.33286
R2629 VDDA.n724 VDDA.n721 5.33286
R2630 VDDA.n702 VDDA.n699 5.33286
R2631 VDDA.n632 VDDA.n335 5.33286
R2632 VDDA.n733 VDDA.n302 5.33286
R2633 VDDA.n785 VDDA.n317 5.33286
R2634 VDDA.n713 VDDA.n325 5.33286
R2635 VDDA.n621 VDDA.n331 5.33286
R2636 VDDA.n113 VDDA.n112 3.75335
R2637 VDDA.n111 VDDA.n72 3.75335
R2638 VDDA.n105 VDDA.n104 3.75335
R2639 VDDA.n103 VDDA.n102 3.75335
R2640 VDDA.n744 VDDA.n740 3.75335
R2641 VDDA.n743 VDDA.n742 3.75335
R2642 VDDA.n781 VDDA.n777 3.75335
R2643 VDDA.n780 VDDA.n779 3.75335
R2644 VDDA.n725 VDDA.n321 3.75335
R2645 VDDA.n724 VDDA.n723 3.75335
R2646 VDDA.n703 VDDA.n329 3.75335
R2647 VDDA.n702 VDDA.n701 3.75335
R2648 VDDA.n633 VDDA.n629 3.75335
R2649 VDDA.n632 VDDA.n631 3.75335
R2650 VDDA.n736 VDDA.n733 3.75335
R2651 VDDA.n735 VDDA.n734 3.75335
R2652 VDDA.n772 VDDA.n317 3.75335
R2653 VDDA.n773 VDDA.n771 3.75335
R2654 VDDA.n707 VDDA.n325 3.75335
R2655 VDDA.n708 VDDA.n706 3.75335
R2656 VDDA.n624 VDDA.n621 3.75335
R2657 VDDA.n623 VDDA.n622 3.75335
R2658 VDDA.n640 VDDA.n636 3.75335
R2659 VDDA.n639 VDDA.n638 3.75335
R2660 VDDA.n660 VDDA.n659 3.53508
R2661 VDDA.n659 VDDA.n658 3.53508
R2662 VDDA.n666 VDDA.n665 3.53508
R2663 VDDA.n665 VDDA.n343 3.53508
R2664 VDDA.n611 VDDA.n610 3.53508
R2665 VDDA.n610 VDDA.n609 3.53508
R2666 VDDA.n587 VDDA.n586 3.53508
R2667 VDDA.n586 VDDA.n582 3.53508
R2668 VDDA.n651 VDDA.n650 3.53508
R2669 VDDA.n650 VDDA.n649 3.53508
R2670 VDDA.n357 VDDA.n352 3.53508
R2671 VDDA.n354 VDDA.n352 3.53508
R2672 VDDA.n422 VDDA.n421 3.53508
R2673 VDDA.n419 VDDA.n417 3.53508
R2674 VDDA.n421 VDDA.n420 3.53508
R2675 VDDA.n404 VDDA.n403 3.53508
R2676 VDDA.n399 VDDA.n398 3.53508
R2677 VDDA.n403 VDDA.n402 3.53508
R2678 VDDA.n565 VDDA.n476 3.53508
R2679 VDDA.n566 VDDA.n565 3.53508
R2680 VDDA.n528 VDDA.n518 3.53508
R2681 VDDA.n522 VDDA.n518 3.53508
R2682 VDDA.n86 VDDA.n76 3.40194
R2683 VDDA.n81 VDDA.n80 3.40194
R2684 VDDA.n768 VDDA.n767 3.40194
R2685 VDDA.n766 VDDA.n762 3.40194
R2686 VDDA.n757 VDDA.n756 3.40194
R2687 VDDA.n755 VDDA.n751 3.40194
R2688 VDDA.n141 VDDA.n62 3.2005
R2689 VDDA.n152 VDDA.n151 3.2005
R2690 VDDA.n165 VDDA.n164 3.2005
R2691 VDDA.n173 VDDA.n49 3.2005
R2692 VDDA.n186 VDDA.n44 3.2005
R2693 VDDA.n197 VDDA.n196 3.2005
R2694 VDDA.n210 VDDA.n209 3.2005
R2695 VDDA.n245 VDDA.n244 3.2005
R2696 VDDA.n272 VDDA.n271 3.2005
R2697 VDDA.n672 VDDA.n340 3.2005
R2698 VDDA.n689 VDDA.n688 3.2005
R2699 VDDA.n690 VDDA.n689 3.2005
R2700 VDDA.n698 VDDA.n697 3.2005
R2701 VDDA.n540 VDDA.n539 3.2005
R2702 VDDA.n539 VDDA.n538 3.2005
R2703 VDDA.n83 VDDA.n76 2.39444
R2704 VDDA.n82 VDDA.n81 2.39444
R2705 VDDA.n767 VDDA.n761 2.39444
R2706 VDDA.n766 VDDA.n765 2.39444
R2707 VDDA.n756 VDDA.n750 2.39444
R2708 VDDA.n755 VDDA.n754 2.39444
R2709 VDDA.n762 VDDA.n307 2.32777
R2710 VDDA.n757 VDDA.n308 2.32777
R2711 VDDA.n482 VDDA.n481 2.27782
R2712 VDDA.n483 VDDA.n482 2.27782
R2713 VDDA.n559 VDDA.n557 2.27782
R2714 VDDA.n485 VDDA.n483 2.27782
R2715 VDDA.n561 VDDA.n481 2.27782
R2716 VDDA.n557 VDDA.n485 2.27782
R2717 VDDA.n517 VDDA.n516 0.703395
R2718 VDDA.n121 VDDA.n71 0.203053
R2719 VDDA.n128 VDDA.n127 0.202927
R2720 VDDA.n595 VDDA.n581 0.193961
R2721 VDDA.n300 VDDA.n299 0.193958
R2722 VDDA.n130 VDDA.n129 0.193477
R2723 VDDA.n471 VDDA.n363 0.188
R2724 VDDA.n122 VDDA.n121 0.15675
R2725 VDDA.n123 VDDA.n122 0.15675
R2726 VDDA.n123 VDDA.n69 0.15675
R2727 VDDA.n127 VDDA.n69 0.15675
R2728 VDDA.n130 VDDA.n65 0.15675
R2729 VDDA.n136 VDDA.n65 0.15675
R2730 VDDA.n137 VDDA.n136 0.15675
R2731 VDDA.n138 VDDA.n137 0.15675
R2732 VDDA.n138 VDDA.n63 0.15675
R2733 VDDA.n142 VDDA.n63 0.15675
R2734 VDDA.n143 VDDA.n142 0.15675
R2735 VDDA.n143 VDDA.n61 0.15675
R2736 VDDA.n147 VDDA.n61 0.15675
R2737 VDDA.n148 VDDA.n147 0.15675
R2738 VDDA.n149 VDDA.n148 0.15675
R2739 VDDA.n149 VDDA.n58 0.15675
R2740 VDDA.n154 VDDA.n58 0.15675
R2741 VDDA.n155 VDDA.n154 0.15675
R2742 VDDA.n156 VDDA.n155 0.15675
R2743 VDDA.n156 VDDA.n55 0.15675
R2744 VDDA.n161 VDDA.n55 0.15675
R2745 VDDA.n162 VDDA.n161 0.15675
R2746 VDDA.n163 VDDA.n162 0.15675
R2747 VDDA.n163 VDDA.n52 0.15675
R2748 VDDA.n168 VDDA.n52 0.15675
R2749 VDDA.n169 VDDA.n168 0.15675
R2750 VDDA.n170 VDDA.n169 0.15675
R2751 VDDA.n170 VDDA.n50 0.15675
R2752 VDDA.n174 VDDA.n50 0.15675
R2753 VDDA.n175 VDDA.n174 0.15675
R2754 VDDA.n175 VDDA.n47 0.15675
R2755 VDDA.n181 VDDA.n47 0.15675
R2756 VDDA.n182 VDDA.n181 0.15675
R2757 VDDA.n183 VDDA.n182 0.15675
R2758 VDDA.n183 VDDA.n45 0.15675
R2759 VDDA.n187 VDDA.n45 0.15675
R2760 VDDA.n188 VDDA.n187 0.15675
R2761 VDDA.n188 VDDA.n43 0.15675
R2762 VDDA.n192 VDDA.n43 0.15675
R2763 VDDA.n193 VDDA.n192 0.15675
R2764 VDDA.n194 VDDA.n193 0.15675
R2765 VDDA.n194 VDDA.n40 0.15675
R2766 VDDA.n199 VDDA.n40 0.15675
R2767 VDDA.n200 VDDA.n199 0.15675
R2768 VDDA.n201 VDDA.n200 0.15675
R2769 VDDA.n201 VDDA.n37 0.15675
R2770 VDDA.n206 VDDA.n37 0.15675
R2771 VDDA.n207 VDDA.n206 0.15675
R2772 VDDA.n208 VDDA.n207 0.15675
R2773 VDDA.n208 VDDA.n34 0.15675
R2774 VDDA.n213 VDDA.n34 0.15675
R2775 VDDA.n214 VDDA.n213 0.15675
R2776 VDDA.n215 VDDA.n214 0.15675
R2777 VDDA.n215 VDDA.n32 0.15675
R2778 VDDA.n221 VDDA.n32 0.15675
R2779 VDDA.n222 VDDA.n221 0.15675
R2780 VDDA.n223 VDDA.n222 0.15675
R2781 VDDA.n223 VDDA.n30 0.15675
R2782 VDDA.n227 VDDA.n30 0.15675
R2783 VDDA.n228 VDDA.n227 0.15675
R2784 VDDA.n228 VDDA.n27 0.15675
R2785 VDDA.n232 VDDA.n27 0.15675
R2786 VDDA.n233 VDDA.n232 0.15675
R2787 VDDA.n234 VDDA.n233 0.15675
R2788 VDDA.n234 VDDA.n25 0.15675
R2789 VDDA.n240 VDDA.n25 0.15675
R2790 VDDA.n241 VDDA.n240 0.15675
R2791 VDDA.n242 VDDA.n241 0.15675
R2792 VDDA.n242 VDDA.n22 0.15675
R2793 VDDA.n247 VDDA.n22 0.15675
R2794 VDDA.n248 VDDA.n247 0.15675
R2795 VDDA.n249 VDDA.n248 0.15675
R2796 VDDA.n249 VDDA.n19 0.15675
R2797 VDDA.n254 VDDA.n19 0.15675
R2798 VDDA.n255 VDDA.n254 0.15675
R2799 VDDA.n256 VDDA.n255 0.15675
R2800 VDDA.n256 VDDA.n16 0.15675
R2801 VDDA.n261 VDDA.n16 0.15675
R2802 VDDA.n262 VDDA.n261 0.15675
R2803 VDDA.n263 VDDA.n262 0.15675
R2804 VDDA.n263 VDDA.n14 0.15675
R2805 VDDA.n267 VDDA.n14 0.15675
R2806 VDDA.n268 VDDA.n267 0.15675
R2807 VDDA.n269 VDDA.n268 0.15675
R2808 VDDA.n269 VDDA.n11 0.15675
R2809 VDDA.n274 VDDA.n11 0.15675
R2810 VDDA.n275 VDDA.n274 0.15675
R2811 VDDA.n276 VDDA.n275 0.15675
R2812 VDDA.n276 VDDA.n9 0.15675
R2813 VDDA.n280 VDDA.n9 0.15675
R2814 VDDA.n281 VDDA.n280 0.15675
R2815 VDDA.n281 VDDA.n6 0.15675
R2816 VDDA.n285 VDDA.n6 0.15675
R2817 VDDA.n286 VDDA.n285 0.15675
R2818 VDDA.n287 VDDA.n286 0.15675
R2819 VDDA.n287 VDDA.n4 0.15675
R2820 VDDA.n293 VDDA.n4 0.15675
R2821 VDDA.n294 VDDA.n293 0.15675
R2822 VDDA.n295 VDDA.n294 0.15675
R2823 VDDA.n295 VDDA.n2 0.15675
R2824 VDDA.n299 VDDA.n2 0.15675
R2825 VDDA.n434 VDDA.n433 0.15675
R2826 VDDA.n434 VDDA.n377 0.15675
R2827 VDDA.n439 VDDA.n377 0.15675
R2828 VDDA.n442 VDDA.n441 0.15675
R2829 VDDA.n442 VDDA.n374 0.15675
R2830 VDDA.n446 VDDA.n374 0.15675
R2831 VDDA.n449 VDDA.n448 0.15675
R2832 VDDA.n449 VDDA.n371 0.15675
R2833 VDDA.n453 VDDA.n371 0.15675
R2834 VDDA.n456 VDDA.n455 0.15675
R2835 VDDA.n456 VDDA.n368 0.15675
R2836 VDDA.n460 VDDA.n368 0.15675
R2837 VDDA.n463 VDDA.n462 0.15675
R2838 VDDA.n467 VDDA.n466 0.15675
R2839 VDDA.n468 VDDA.n467 0.15675
R2840 VDDA.n468 VDDA.n363 0.15675
R2841 VDDA.n535 VDDA.n516 0.15675
R2842 VDDA.n536 VDDA.n535 0.15675
R2843 VDDA.n537 VDDA.n536 0.15675
R2844 VDDA.n537 VDDA.n513 0.15675
R2845 VDDA.n542 VDDA.n513 0.15675
R2846 VDDA.n543 VDDA.n542 0.15675
R2847 VDDA.n544 VDDA.n543 0.15675
R2848 VDDA.n544 VDDA.n510 0.15675
R2849 VDDA.n510 VDDA.n509 0.15675
R2850 VDDA.n549 VDDA.n509 0.15675
R2851 VDDA.n550 VDDA.n549 0.15675
R2852 VDDA.n551 VDDA.n550 0.15675
R2853 VDDA.n552 VDDA.n551 0.15675
R2854 VDDA.n552 VDDA.n507 0.15675
R2855 VDDA.n507 VDDA.n506 0.15675
R2856 VDDA.n506 VDDA.n505 0.15675
R2857 VDDA.n505 VDDA.n487 0.15675
R2858 VDDA.n501 VDDA.n487 0.15675
R2859 VDDA.n501 VDDA.n500 0.15675
R2860 VDDA.n500 VDDA.n499 0.15675
R2861 VDDA.n499 VDDA.n490 0.15675
R2862 VDDA.n495 VDDA.n490 0.15675
R2863 VDDA.n495 VDDA.n494 0.15675
R2864 VDDA.n494 VDDA.n493 0.15675
R2865 VDDA.n493 VDDA.n473 0.15675
R2866 VDDA.n575 VDDA.n473 0.15675
R2867 VDDA.n576 VDDA.n575 0.15675
R2868 VDDA.n577 VDDA.n576 0.15675
R2869 VDDA.n596 VDDA.n595 0.15675
R2870 VDDA.n597 VDDA.n596 0.15675
R2871 VDDA.n597 VDDA.n361 0.15675
R2872 VDDA.n601 VDDA.n361 0.15675
R2873 VDDA.n602 VDDA.n601 0.15675
R2874 VDDA.n605 VDDA.n602 0.15675
R2875 VDDA.n605 VDDA.n604 0.15675
R2876 VDDA.n604 VDDA.n603 0.15675
R2877 VDDA.n675 VDDA.n674 0.15675
R2878 VDDA.n676 VDDA.n675 0.15675
R2879 VDDA.n676 VDDA.n339 0.15675
R2880 VDDA.n680 VDDA.n339 0.15675
R2881 VDDA.n681 VDDA.n680 0.15675
R2882 VDDA.n681 VDDA.n337 0.15675
R2883 VDDA.n685 VDDA.n337 0.15675
R2884 VDDA.n686 VDDA.n685 0.15675
R2885 VDDA.n687 VDDA.n686 0.15675
R2886 VDDA.n687 VDDA.n333 0.15675
R2887 VDDA.n693 VDDA.n333 0.15675
R2888 VDDA.n694 VDDA.n693 0.15675
R2889 VDDA.n695 VDDA.n694 0.15675
R2890 VDDA.n695 VDDA.n323 0.15675
R2891 VDDA.n716 VDDA.n323 0.15675
R2892 VDDA.n717 VDDA.n716 0.15675
R2893 VDDA.n718 VDDA.n717 0.15675
R2894 VDDA.n718 VDDA.n314 0.15675
R2895 VDDA.n788 VDDA.n314 0.15675
R2896 VDDA.n789 VDDA.n788 0.15675
R2897 VDDA.n790 VDDA.n789 0.15675
R2898 VDDA.n790 VDDA.n312 0.15675
R2899 VDDA.n794 VDDA.n312 0.15675
R2900 VDDA.n795 VDDA.n794 0.15675
R2901 VDDA.n796 VDDA.n795 0.15675
R2902 VDDA.n796 VDDA.n310 0.15675
R2903 VDDA.n800 VDDA.n310 0.15675
R2904 VDDA.n801 VDDA.n800 0.15675
R2905 VDDA.n801 VDDA.n306 0.15675
R2906 VDDA.n806 VDDA.n306 0.15675
R2907 VDDA.n807 VDDA.n806 0.15675
R2908 VDDA.n808 VDDA.n807 0.15675
R2909 VDDA.n808 VDDA.n304 0.15675
R2910 VDDA.n812 VDDA.n304 0.15675
R2911 VDDA.n813 VDDA.n812 0.15675
R2912 VDDA.n814 VDDA.n813 0.15675
R2913 VDDA.n814 VDDA.n0 0.15675
R2914 VDDA VDDA.n0 0.1255
R2915 VDDA.n577 VDDA 0.122375
R2916 VDDA.n432 VDDA.n431 0.100307
R2917 VDDA.n433 VDDA.n432 0.09425
R2918 VDDA.n441 VDDA.n440 0.09425
R2919 VDDA.n448 VDDA.n447 0.09425
R2920 VDDA.n455 VDDA.n454 0.09425
R2921 VDDA.n462 VDDA.n461 0.09425
R2922 VDDA.n466 VDDA.n365 0.09425
R2923 VDDA.n603 VDDA.n341 0.078625
R2924 VDDA.n674 VDDA.n341 0.078625
R2925 VDDA VDDA.n818 0.063
R2926 VDDA.n440 VDDA.n439 0.063
R2927 VDDA.n447 VDDA.n446 0.063
R2928 VDDA.n454 VDDA.n453 0.063
R2929 VDDA.n461 VDDA.n460 0.063
R2930 VDDA.n463 VDDA.n365 0.063
R2931 VDDA.n579 VDDA 0.0505
R2932 VCO_FD_magic_0.div120_2_0.div2.t4 VCO_FD_magic_0.div120_2_0.div2.t5 1012.2
R2933 VCO_FD_magic_0.div120_2_0.div2.n0 VCO_FD_magic_0.div120_2_0.div2.t1 663.801
R2934 VCO_FD_magic_0.div120_2_0.div2.n2 VCO_FD_magic_0.div120_2_0.div2.n1 431.401
R2935 VCO_FD_magic_0.div120_2_0.div2.t3 VCO_FD_magic_0.div120_2_0.div2.t6 401.668
R2936 VCO_FD_magic_0.div120_2_0.div2.n0 VCO_FD_magic_0.div120_2_0.div2.t4 361.692
R2937 VCO_FD_magic_0.div120_2_0.div2.n1 VCO_FD_magic_0.div120_2_0.div2.t2 353.467
R2938 VCO_FD_magic_0.div120_2_0.div2.t0 VCO_FD_magic_0.div120_2_0.div2.n2 298.921
R2939 VCO_FD_magic_0.div120_2_0.div2.n1 VCO_FD_magic_0.div120_2_0.div2.t3 257.067
R2940 VCO_FD_magic_0.div120_2_0.div2.n2 VCO_FD_magic_0.div120_2_0.div2.n0 67.2005
R2941 a_7630_n1440.n4 a_7630_n1440.t1 752.333
R2942 a_7630_n1440.t2 a_7630_n1440.n5 752.333
R2943 a_7630_n1440.n0 a_7630_n1440.t5 514.134
R2944 a_7630_n1440.n3 a_7630_n1440.n2 366.856
R2945 a_7630_n1440.n5 a_7630_n1440.t0 254.333
R2946 a_7630_n1440.n3 a_7630_n1440.t3 190.123
R2947 a_7630_n1440.n4 a_7630_n1440.n3 187.201
R2948 a_7630_n1440.n2 a_7630_n1440.n1 176.733
R2949 a_7630_n1440.n1 a_7630_n1440.n0 176.733
R2950 a_7630_n1440.n2 a_7630_n1440.t6 112.468
R2951 a_7630_n1440.n1 a_7630_n1440.t4 112.468
R2952 a_7630_n1440.n0 a_7630_n1440.t7 112.468
R2953 a_7630_n1440.n5 a_7630_n1440.n4 70.4005
R2954 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R2955 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R2956 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R2957 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R2958 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R2959 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R2960 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R2961 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t0 221.411
R2962 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t2 24.0005
R2963 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t1 24.0005
R2964 a_870_1400.t0 a_870_1400.t1 39.4005
R2965 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 203.528
R2966 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.DOWN_PFD_b.n1 203.528
R2967 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t2 183.935
R2968 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t0 183.935
R2969 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R2970 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R2971 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R2972 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R2973 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R2974 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R2975 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R2976 pfd_8_0.DOWN_b.t0 pfd_8_0.DOWN_b.n2 211.847
R2977 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t1 173.055
R2978 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.J.t2 710.734
R2979 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t4 553.534
R2980 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t0 254.333
R2981 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 206.333
R2982 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n1 70.4005
R2983 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t1 48.0005
R2984 VCO_FD_magic_0.div120_2_0.div5_2_0.J.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.J.t3 48.0005
R2985 VCO_FD_magic_0.div120_2_0.div5_2_0.J VCO_FD_magic_0.div120_2_0.div5_2_0.J.n2 12.8005
R2986 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t0 777.4
R2987 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t6 514.134
R2988 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 364.178
R2989 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 353.467
R2990 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t2 353.467
R2991 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t8 318.702
R2992 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t5 307.909
R2993 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t3 289.2
R2994 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 257.079
R2995 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t1 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 233
R2996 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t11 192.8
R2997 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 176.733
R2998 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t9 112.468
R2999 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n4 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t10 112.468
R3000 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t4 112.468
R3001 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n5 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.t7 112.468
R3002 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n3 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n2 96.4005
R3003 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n1 38.2642
R3004 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n7 VCO_FD_magic_0.div120_2_0.div5_2_0.Q2_b.n6 21.3338
R3005 VCO_FD_magic_0.div120_2_0.div24.n3 VCO_FD_magic_0.div120_2_0.div24.n2 919.244
R3006 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div24.n7 912.303
R3007 VCO_FD_magic_0.div120_2_0.div24.t9 VCO_FD_magic_0.div120_2_0.div24.t11 819.4
R3008 VCO_FD_magic_0.div120_2_0.div24.n9 VCO_FD_magic_0.div120_2_0.div24.n8 628.734
R3009 VCO_FD_magic_0.div120_2_0.div24.n2 VCO_FD_magic_0.div120_2_0.div24.n1 520.361
R3010 VCO_FD_magic_0.div120_2_0.div24.n7 VCO_FD_magic_0.div120_2_0.div24.n6 364.178
R3011 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t8 337.401
R3012 VCO_FD_magic_0.div120_2_0.div24.n10 VCO_FD_magic_0.div120_2_0.div24.t9 336.25
R3013 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t13 305.267
R3014 VCO_FD_magic_0.div120_2_0.div24.n9 VCO_FD_magic_0.div120_2_0.div24.t0 257.534
R3015 VCO_FD_magic_0.div120_2_0.div24.n4 VCO_FD_magic_0.div120_2_0.div24.t12 192.8
R3016 VCO_FD_magic_0.div120_2_0.div24.n1 VCO_FD_magic_0.div120_2_0.div24.n0 176.733
R3017 VCO_FD_magic_0.div120_2_0.div24.n6 VCO_FD_magic_0.div120_2_0.div24.n5 176.733
R3018 VCO_FD_magic_0.div120_2_0.div24.n4 VCO_FD_magic_0.div120_2_0.div24.n3 160.667
R3019 VCO_FD_magic_0.div120_2_0.div24.n3 VCO_FD_magic_0.div120_2_0.div24.t7 144.601
R3020 VCO_FD_magic_0.div120_2_0.div24.n2 VCO_FD_magic_0.div120_2_0.div24.t4 131.976
R3021 VCO_FD_magic_0.div120_2_0.div24.n1 VCO_FD_magic_0.div120_2_0.div24.t3 128.534
R3022 VCO_FD_magic_0.div120_2_0.div24.n0 VCO_FD_magic_0.div120_2_0.div24.t6 128.534
R3023 VCO_FD_magic_0.div120_2_0.div24.n6 VCO_FD_magic_0.div120_2_0.div24.t14 112.468
R3024 VCO_FD_magic_0.div120_2_0.div24.n5 VCO_FD_magic_0.div120_2_0.div24.t5 112.468
R3025 VCO_FD_magic_0.div120_2_0.div24.n7 VCO_FD_magic_0.div120_2_0.div24.t10 112.468
R3026 VCO_FD_magic_0.div120_2_0.div24.n5 VCO_FD_magic_0.div120_2_0.div24.n4 96.4005
R3027 VCO_FD_magic_0.div120_2_0.div24.n8 VCO_FD_magic_0.div120_2_0.div24.t2 78.8005
R3028 VCO_FD_magic_0.div120_2_0.div24.n8 VCO_FD_magic_0.div120_2_0.div24.t1 78.8005
R3029 VCO_FD_magic_0.div120_2_0.div24.n10 VCO_FD_magic_0.div120_2_0.div24.n9 11.2005
R3030 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div24.n10 6.4005
R3031 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div3_3_0.H.t1 710.734
R3032 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t4 553.534
R3033 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t3 254.333
R3034 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 206.333
R3035 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n1 70.4005
R3036 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t0 48.0005
R3037 VCO_FD_magic_0.div120_2_0.div3_3_0.H.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.H.t2 48.0005
R3038 VCO_FD_magic_0.div120_2_0.div3_3_0.H VCO_FD_magic_0.div120_2_0.div3_3_0.H.n2 12.8005
R3039 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t0 663.801
R3040 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t2 514.134
R3041 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t3 479.284
R3042 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 344.8
R3043 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t5 289.2
R3044 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 275.454
R3045 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t4 241
R3046 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.I.t6 112.468
R3047 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n0 97.9205
R3048 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.I.n1 64.2672
R3049 pfd_8_0.DOWN.t3 pfd_8_0.DOWN.n0 605.311
R3050 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t3 399.497
R3051 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 240.327
R3052 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t0 148.736
R3053 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t2 24.487
R3054 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t3 326.658
R3055 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t6 297.233
R3056 pfd_8_0.UP_input.t5 pfd_8_0.UP_input.n5 297.233
R3057 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n1 257.067
R3058 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 246.275
R3059 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t2 241.928
R3060 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n1 226.942
R3061 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n2 226.942
R3062 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.n4 216.9
R3063 pfd_8_0.UP_input.t0 pfd_8_0.UP_input.n7 209.928
R3064 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t1 145.536
R3065 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n0 144
R3066 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t6 92.3838
R3067 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t5 92.3838
R3068 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t7 80.3338
R3069 pfd_8_0.UP_input.t7 pfd_8_0.UP_input.n3 80.3338
R3070 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t4 80.3338
R3071 pfd_8_0.UP_input.t4 pfd_8_0.UP_input.n1 80.3338
R3072 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.n1 507.072
R3073 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.n0 409.067
R3074 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.t3 369.534
R3075 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 209.928
R3076 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t0 177.536
R3077 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.t1 24.0223
R3078 VCO_FD_magic_0.vco2_3_0.V1.n1 VCO_FD_magic_0.vco2_3_0.V1.t5 600.206
R3079 VCO_FD_magic_0.vco2_3_0.V1.t2 VCO_FD_magic_0.vco2_3_0.V1.n5 576.192
R3080 VCO_FD_magic_0.vco2_3_0.V1.n2 VCO_FD_magic_0.vco2_3_0.V1.n1 568.072
R3081 VCO_FD_magic_0.vco2_3_0.V1.n4 VCO_FD_magic_0.vco2_3_0.V1.n2 392.486
R3082 VCO_FD_magic_0.vco2_3_0.V1.n0 VCO_FD_magic_0.vco2_3_0.V1.t1 289.791
R3083 VCO_FD_magic_0.vco2_3_0.V1.n5 VCO_FD_magic_0.vco2_3_0.V1.n4 168.067
R3084 VCO_FD_magic_0.vco2_3_0.V1.n3 VCO_FD_magic_0.vco2_3_0.V1.n0 97.9242
R3085 VCO_FD_magic_0.vco2_3_0.V1.n4 VCO_FD_magic_0.vco2_3_0.V1.n3 37.7572
R3086 VCO_FD_magic_0.vco2_3_0.V1.n1 VCO_FD_magic_0.vco2_3_0.V1.t3 32.1338
R3087 VCO_FD_magic_0.vco2_3_0.V1.n2 VCO_FD_magic_0.vco2_3_0.V1.t4 32.1338
R3088 VCO_FD_magic_0.vco2_3_0.V1.n3 VCO_FD_magic_0.vco2_3_0.V1.t0 32.1338
R3089 VCO_FD_magic_0.vco2_3_0.V1.n5 VCO_FD_magic_0.vco2_3_0.V1.n0 28.3357
R3090 VCO_FD_magic_0.vco2_3_0.V4.n0 VCO_FD_magic_0.vco2_3_0.V4.t1 421.027
R3091 VCO_FD_magic_0.vco2_3_0.V4.n0 VCO_FD_magic_0.vco2_3_0.V4.t2 348.81
R3092 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V4.t0 280.05
R3093 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V4.n0 36.1094
R3094 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t1 685.134
R3095 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.G.t0 663.801
R3096 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t3 534.268
R3097 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.G.t2 340.521
R3098 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.G.n0 105.6
R3099 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.G.n1 21.3338
R3100 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n5 424.447
R3101 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n4 354.048
R3102 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n1 313
R3103 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.t14 297.233
R3104 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t14 297.233
R3105 pfd_8_0.opamp_out.t13 pfd_8_0.opamp_out.n11 297.233
R3106 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t2 281.596
R3107 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n0 242.601
R3108 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.n2 220.8
R3109 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.n6 220.8
R3110 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.n10 216.9
R3111 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n8 216.9
R3112 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n12 215.107
R3113 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.n8 184.768
R3114 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t4 118.666
R3115 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t15 80.3338
R3116 pfd_8_0.opamp_out.t15 pfd_8_0.opamp_out.n9 80.3338
R3117 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t10 80.3338
R3118 pfd_8_0.opamp_out.t10 pfd_8_0.opamp_out.n8 80.3338
R3119 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t13 80.3338
R3120 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n14 78.9255
R3121 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.t12 70.0829
R3122 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t11 63.6829
R3123 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n3 62.4005
R3124 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n7 60.8005
R3125 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n13 60.2361
R3126 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t6 60.0005
R3127 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t1 60.0005
R3128 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t8 60.0005
R3129 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t9 60.0005
R3130 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t3 49.2505
R3131 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t5 49.2505
R3132 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t0 49.2505
R3133 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t7 49.2505
R3134 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n15 1.6005
R3135 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t8 377.567
R3136 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t6 321.334
R3137 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 233.476
R3138 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t7 216.9
R3139 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n4 199.462
R3140 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 189.898
R3141 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n3 172.502
R3142 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 172.5
R3143 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t9 112.468
R3144 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n5 70.4005
R3145 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 50.088
R3146 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t1 24.6255
R3147 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t0 24.6255
R3148 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t3 24.6255
R3149 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t2 24.6255
R3150 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t4 15.0005
R3151 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t5 15.0005
R3152 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.313
R3153 a_6320_5840.n7 a_6320_5840.n5 482.582
R3154 a_6320_5840.n10 a_6320_5840.t6 304.634
R3155 a_6320_5840.n3 a_6320_5840.t4 304.634
R3156 a_6320_5840.t8 a_6320_5840.n10 277.914
R3157 a_6320_5840.n3 a_6320_5840.t5 276.289
R3158 a_6320_5840.n8 a_6320_5840.n1 204.201
R3159 a_6320_5840.n4 a_6320_5840.n2 204.201
R3160 a_6320_5840.n9 a_6320_5840.n0 204.201
R3161 a_6320_5840.n7 a_6320_5840.n6 120.981
R3162 a_6320_5840.n8 a_6320_5840.n4 74.6672
R3163 a_6320_5840.n9 a_6320_5840.n8 74.6672
R3164 a_6320_5840.n1 a_6320_5840.t3 60.0005
R3165 a_6320_5840.n1 a_6320_5840.t11 60.0005
R3166 a_6320_5840.t5 a_6320_5840.n2 60.0005
R3167 a_6320_5840.n2 a_6320_5840.t2 60.0005
R3168 a_6320_5840.n0 a_6320_5840.t10 60.0005
R3169 a_6320_5840.n0 a_6320_5840.t7 60.0005
R3170 a_6320_5840.n8 a_6320_5840.n7 37.763
R3171 a_6320_5840.n5 a_6320_5840.t12 24.0005
R3172 a_6320_5840.n5 a_6320_5840.t1 24.0005
R3173 a_6320_5840.n6 a_6320_5840.t0 24.0005
R3174 a_6320_5840.n6 a_6320_5840.t9 24.0005
R3175 a_6320_5840.n4 a_6320_5840.n3 16.0005
R3176 a_6320_5840.n10 a_6320_5840.n9 16.0005
R3177 opamp_cell_4_0.n_right.t3 opamp_cell_4_0.n_right.n6 1010.36
R3178 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 404.8
R3179 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 322.048
R3180 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 316.2
R3181 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t8 289.2
R3182 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R3183 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t6 289.2
R3184 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t5 232.968
R3185 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R3186 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R3187 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 199.829
R3188 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R3189 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t2 60.0005
R3190 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t4 49.2505
R3191 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t0 49.2505
R3192 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 359.894
R3193 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R3194 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R3195 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t2 252.248
R3196 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R3197 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t4 192.8
R3198 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 192.8
R3199 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R3200 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t1 60.0005
R3201 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t0 60.0005
R3202 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R3203 opamp_cell_4_0.n_left.t5 opamp_cell_4_0.n_left.n5 49.2505
R3204 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t3 49.2505
R3205 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.C.t0 702.201
R3206 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t4 349.433
R3207 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t3 276.733
R3208 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 206.333
R3209 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 48.0005
R3210 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n1 48.0005
R3211 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t1 48.0005
R3212 VCO_FD_magic_0.div120_2_0.div2_4_0.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.C.t2 48.0005
R3213 VCO_FD_magic_0.div120_2_0.div8.t4 VCO_FD_magic_0.div120_2_0.div8.t5 1012.2
R3214 VCO_FD_magic_0.div120_2_0.div8.n0 VCO_FD_magic_0.div120_2_0.div8.t1 663.801
R3215 VCO_FD_magic_0.div120_2_0.div8.n2 VCO_FD_magic_0.div120_2_0.div8.n1 431.401
R3216 VCO_FD_magic_0.div120_2_0.div8.t3 VCO_FD_magic_0.div120_2_0.div8.t6 401.668
R3217 VCO_FD_magic_0.div120_2_0.div8.n0 VCO_FD_magic_0.div120_2_0.div8.t4 361.692
R3218 VCO_FD_magic_0.div120_2_0.div8.t0 VCO_FD_magic_0.div120_2_0.div8.n2 298.921
R3219 VCO_FD_magic_0.div120_2_0.div8.n1 VCO_FD_magic_0.div120_2_0.div8.t3 257.067
R3220 VCO_FD_magic_0.div120_2_0.div8.n1 VCO_FD_magic_0.div120_2_0.div8.t2 208.868
R3221 VCO_FD_magic_0.div120_2_0.div8.n2 VCO_FD_magic_0.div120_2_0.div8.n0 67.2005
R3222 a_6490_4630.t2 a_6490_4630.n6 1112.76
R3223 a_6490_4630.n3 a_6490_4630.n2 441.433
R3224 a_6490_4630.n2 a_6490_4630.n1 379.647
R3225 a_6490_4630.n2 a_6490_4630.n0 258.601
R3226 a_6490_4630.n6 a_6490_4630.t6 208.868
R3227 a_6490_4630.n5 a_6490_4630.t7 208.868
R3228 a_6490_4630.n4 a_6490_4630.t8 208.868
R3229 a_6490_4630.n3 a_6490_4630.t5 208.868
R3230 a_6490_4630.n6 a_6490_4630.n5 208.868
R3231 a_6490_4630.n5 a_6490_4630.n4 208.868
R3232 a_6490_4630.n4 a_6490_4630.n3 208.868
R3233 a_6490_4630.n0 a_6490_4630.t4 60.0005
R3234 a_6490_4630.n0 a_6490_4630.t3 60.0005
R3235 a_6490_4630.n1 a_6490_4630.t1 49.2505
R3236 a_6490_4630.n1 a_6490_4630.t0 49.2505
R3237 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R3238 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R3239 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R3240 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R3241 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t1 172.458
R3242 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R3243 pfd_8_0.before_Reset.t0 pfd_8_0.before_Reset.n2 19.7005
R3244 a_2350_1400.t1 a_2350_1400.n2 500.086
R3245 a_2350_1400.n1 a_2350_1400.n0 473.334
R3246 a_2350_1400.n0 a_2350_1400.t3 465.933
R3247 a_2350_1400.t1 a_2350_1400.n2 461.389
R3248 a_2350_1400.n0 a_2350_1400.t2 321.334
R3249 a_2350_1400.n1 a_2350_1400.t0 177.577
R3250 a_2350_1400.n2 a_2350_1400.n1 48.3899
R3251 VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t1 713.933
R3252 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.A.t0 327.401
R3253 VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.A.t2 314.233
R3254 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.A.n0 9.6005
R3255 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_2.B.t1 96.0005
R3256 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t8 918.318
R3257 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R3258 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t10 377.567
R3259 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t9 377.567
R3260 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R3261 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R3262 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R3263 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R3264 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R3265 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R3266 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R3267 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t12 120.501
R3268 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t4 120.501
R3269 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t0 120.501
R3270 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t2 120.501
R3271 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t11 120.501
R3272 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t6 120.501
R3273 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R3274 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R3275 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R3276 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R3277 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R3278 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t1 19.7005
R3279 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t5 19.7005
R3280 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t7 19.7005
R3281 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t3 19.7005
R3282 F_REF.n0 F_REF.t0 514.134
R3283 F_REF.n0 F_REF.t1 273.134
R3284 F_REF F_REF.n0 216.9
R3285 a_n30_1400.t0 a_n30_1400.t1 39.4005
R3286 I_IN.n1 I_IN.n0 1269.42
R3287 I_IN.n1 I_IN.t0 275.325
R3288 I_IN.n6 I_IN.n2 248.4
R3289 I_IN.n4 I_IN.t4 238.892
R3290 I_IN.n4 I_IN.t5 161.371
R3291 I_IN.n0 I_IN.t6 151.792
R3292 I_IN.n5 I_IN.n4 151.34
R3293 I_IN.n2 I_IN.t2 140.583
R3294 I_IN.n2 I_IN.t0 140.583
R3295 I_IN.n6 I_IN.n3 98.6614
R3296 I_IN.t2 I_IN.n1 80.3338
R3297 I_IN.n0 I_IN.t7 44.2902
R3298 I_IN.n3 I_IN.t3 15.0005
R3299 I_IN.n3 I_IN.t1 15.0005
R3300 I_IN.n6 I_IN.n5 9.3005
R3301 I_IN I_IN.n6 3.2005
R3302 I_IN.n5 I_IN 0.063
R3303 VCO_FD_magic_0.div120_2_0.div4.t6 VCO_FD_magic_0.div120_2_0.div4.t3 1012.2
R3304 VCO_FD_magic_0.div120_2_0.div4.n0 VCO_FD_magic_0.div120_2_0.div4.t0 663.801
R3305 VCO_FD_magic_0.div120_2_0.div4.n2 VCO_FD_magic_0.div120_2_0.div4.n1 431.401
R3306 VCO_FD_magic_0.div120_2_0.div4.t4 VCO_FD_magic_0.div120_2_0.div4.t2 401.668
R3307 VCO_FD_magic_0.div120_2_0.div4.n0 VCO_FD_magic_0.div120_2_0.div4.t6 361.692
R3308 VCO_FD_magic_0.div120_2_0.div4.n1 VCO_FD_magic_0.div120_2_0.div4.t5 353.467
R3309 VCO_FD_magic_0.div120_2_0.div4.t1 VCO_FD_magic_0.div120_2_0.div4.n2 298.921
R3310 VCO_FD_magic_0.div120_2_0.div4.n1 VCO_FD_magic_0.div120_2_0.div4.t4 257.067
R3311 VCO_FD_magic_0.div120_2_0.div4.n2 VCO_FD_magic_0.div120_2_0.div4.n0 67.2005
R3312 a_6330_n1440.n0 a_6330_n1440.t1 752.333
R3313 a_6330_n1440.t2 a_6330_n1440.n5 752.333
R3314 a_6330_n1440.n1 a_6330_n1440.t6 514.134
R3315 a_6330_n1440.n4 a_6330_n1440.n3 366.856
R3316 a_6330_n1440.n0 a_6330_n1440.t0 254.333
R3317 a_6330_n1440.n4 a_6330_n1440.t5 190.123
R3318 a_6330_n1440.n5 a_6330_n1440.n4 187.201
R3319 a_6330_n1440.n3 a_6330_n1440.n2 176.733
R3320 a_6330_n1440.n2 a_6330_n1440.n1 176.733
R3321 a_6330_n1440.n3 a_6330_n1440.t3 112.468
R3322 a_6330_n1440.n2 a_6330_n1440.t7 112.468
R3323 a_6330_n1440.n1 a_6330_n1440.t4 112.468
R3324 a_6330_n1440.n5 a_6330_n1440.n0 70.4005
R3325 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R3326 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R3327 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R3328 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R3329 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R3330 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R3331 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R3332 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R3333 pfd_8_0.QA.n4 pfd_8_0.QA.t1 221.411
R3334 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R3335 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R3336 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R3337 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R3338 pfd_8_0.QA.n3 pfd_8_0.QA.t0 24.0005
R3339 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R3340 a_8930_n1440.n5 a_8930_n1440.t0 752.333
R3341 a_8930_n1440.n4 a_8930_n1440.t1 752.333
R3342 a_8930_n1440.n0 a_8930_n1440.t4 514.134
R3343 a_8930_n1440.n3 a_8930_n1440.n2 366.856
R3344 a_8930_n1440.t2 a_8930_n1440.n5 254.333
R3345 a_8930_n1440.n3 a_8930_n1440.t5 190.123
R3346 a_8930_n1440.n4 a_8930_n1440.n3 187.201
R3347 a_8930_n1440.n2 a_8930_n1440.n1 176.733
R3348 a_8930_n1440.n1 a_8930_n1440.n0 176.733
R3349 a_8930_n1440.n2 a_8930_n1440.t3 112.468
R3350 a_8930_n1440.n1 a_8930_n1440.t6 112.468
R3351 a_8930_n1440.n0 a_8930_n1440.t7 112.468
R3352 a_8930_n1440.n5 a_8930_n1440.n4 70.4005
R3353 VCO_FD_magic_0.div120_2_0.div2_4_1.C VCO_FD_magic_0.div120_2_0.div2_4_1.C.t0 702.201
R3354 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t4 349.433
R3355 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t3 276.733
R3356 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 206.333
R3357 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t2 48.0005
R3358 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.C.t1 48.0005
R3359 VCO_FD_magic_0.div120_2_0.div2_4_1.C VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 48.0005
R3360 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_1.C.n1 48.0005
R3361 pfd_8_0.DOWN_input.t5 pfd_8_0.DOWN_input.t4 377.567
R3362 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t3 326.658
R3363 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 237.65
R3364 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t1 229.127
R3365 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 196.817
R3366 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t0 158.335
R3367 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t2 158.335
R3368 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 121.6
R3369 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.n2 92.3838
R3370 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t5 92.3838
R3371 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 3.2005
R3372 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 742.51
R3373 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t1 723.534
R3374 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 723.534
R3375 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 684.806
R3376 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 366.856
R3377 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t6 337.401
R3378 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t9 305.267
R3379 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t0 254.333
R3380 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 224.934
R3381 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t11 190.123
R3382 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n7 187.201
R3383 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 176.733
R3384 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 176.733
R3385 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 176.733
R3386 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n3 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t3 144.601
R3387 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t8 131.976
R3388 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t12 128.534
R3389 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t5 128.534
R3390 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n6 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t7 112.468
R3391 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n5 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t10 112.468
R3392 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n4 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.t4 112.468
R3393 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n9 VCO_FD_magic_0.div120_2_0.div3_3_0.CLK.n8 70.4005
R3394 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 701.467
R3395 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t0 694.201
R3396 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t2 321.334
R3397 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.D.t1 260.521
R3398 VCO_FD_magic_0.div120_2_0.div3_3_0.D.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.D.t3 144.601
R3399 VCO_FD_magic_0.div120_2_0.div3_3_0.D VCO_FD_magic_0.div120_2_0.div3_3_0.D.n1 54.4005
R3400 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.C.t3 702.201
R3401 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t4 350.349
R3402 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t1 276.733
R3403 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 206.333
R3404 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n1 48.0005
R3405 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t0 48.0005
R3406 VCO_FD_magic_0.div120_2_0.div3_3_0.C.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.C.t2 48.0005
R3407 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.C.n2 19.2005
R3408 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R3409 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R3410 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R3411 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R3412 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R3413 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R3414 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R3415 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R3416 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R3417 pfd_8_0.QB.n4 pfd_8_0.QB.t2 221.411
R3418 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R3419 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R3420 pfd_8_0.QB.n3 pfd_8_0.QB.t0 24.0005
R3421 pfd_8_0.QB.n3 pfd_8_0.QB.t1 24.0005
R3422 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R3423 a_1910_2020.t0 a_1910_2020.t1 48.0005
R3424 a_6220_5810.n4 a_6220_5810.t12 317.317
R3425 a_6220_5810.n2 a_6220_5810.t11 317.317
R3426 a_6220_5810.n5 a_6220_5810.n4 257.067
R3427 a_6220_5810.n3 a_6220_5810.n2 257.067
R3428 a_6220_5810.n10 a_6220_5810.n9 257.067
R3429 a_6220_5810.t8 a_6220_5810.n12 194.478
R3430 a_6220_5810.n8 a_6220_5810.n7 152
R3431 a_6220_5810.n12 a_6220_5810.n11 152
R3432 a_6220_5810.n1 a_6220_5810.n0 120.981
R3433 a_6220_5810.n7 a_6220_5810.n6 117.781
R3434 a_6220_5810.n7 a_6220_5810.n1 108.8
R3435 a_6220_5810.n8 a_6220_5810.n5 85.6894
R3436 a_6220_5810.n11 a_6220_5810.n3 85.6894
R3437 a_6220_5810.n11 a_6220_5810.n10 85.6894
R3438 a_6220_5810.n9 a_6220_5810.n8 85.6894
R3439 a_6220_5810.n4 a_6220_5810.t10 60.2505
R3440 a_6220_5810.n5 a_6220_5810.t0 60.2505
R3441 a_6220_5810.n2 a_6220_5810.t9 60.2505
R3442 a_6220_5810.n3 a_6220_5810.t2 60.2505
R3443 a_6220_5810.n10 a_6220_5810.t6 60.2505
R3444 a_6220_5810.n9 a_6220_5810.t4 60.2505
R3445 a_6220_5810.n6 a_6220_5810.t5 24.0005
R3446 a_6220_5810.n6 a_6220_5810.t1 24.0005
R3447 a_6220_5810.n0 a_6220_5810.t3 24.0005
R3448 a_6220_5810.n0 a_6220_5810.t7 24.0005
R3449 a_6220_5810.n12 a_6220_5810.n1 3.2005
R3450 VCO_FD_magic_0.div120_2_0.div2_4_2.C VCO_FD_magic_0.div120_2_0.div2_4_2.C.t3 702.201
R3451 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t4 349.433
R3452 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t1 276.733
R3453 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 206.333
R3454 VCO_FD_magic_0.div120_2_0.div2_4_2.C VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 48.0005
R3455 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n2 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n1 48.0005
R3456 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t2 48.0005
R3457 VCO_FD_magic_0.div120_2_0.div2_4_2.C.n0 VCO_FD_magic_0.div120_2_0.div2_4_2.C.t0 48.0005
R3458 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R3459 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R3460 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R3461 pfd_8_0.UP_PFD_b.t1 pfd_8_0.UP_PFD_b.n1 219.528
R3462 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t0 167.935
R3463 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R3464 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R3465 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R3466 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R3467 pfd_8_0.UP.t1 pfd_8_0.UP.n3 229.127
R3468 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R3469 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R3470 pfd_8_0.UP.n3 pfd_8_0.UP.t0 158.335
R3471 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R3472 F_VCO.n3 F_VCO.t3 772.196
R3473 F_VCO.n5 F_VCO.t1 751.801
R3474 F_VCO.n4 F_VCO.n3 607.465
R3475 F_VCO.t3 F_VCO.t2 514.134
R3476 F_VCO.n0 F_VCO.t6 514.134
R3477 F_VCO.n2 F_VCO.t4 289.2
R3478 F_VCO.n0 F_VCO.t7 273.134
R3479 F_VCO.n4 F_VCO.t0 233
R3480 F_VCO F_VCO.n0 216.9
R3481 F_VCO.n3 F_VCO.n2 208.868
R3482 F_VCO F_VCO.n1 194.333
R3483 F_VCO.n2 F_VCO.t5 176.733
R3484 F_VCO.n5 F_VCO.n4 40.3205
R3485 F_VCO F_VCO.n5 38.4005
R3486 F_VCO.n1 F_VCO 24.1005
R3487 F_VCO.n1 F_VCO 24.1005
R3488 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 279.933
R3489 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.I.t1 251.133
R3490 VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t0 48.0005
R3491 VCO_FD_magic_0.div120_2_0.div5_2_0.I.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.I.t2 48.0005
R3492 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.H.t1 96.0005
R3493 V_OSC.t2 V_OSC.t5 401.668
R3494 V_OSC.n1 V_OSC.t1 372.118
R3495 V_OSC.n3 V_OSC.t3 353.467
R3496 V_OSC V_OSC.n3 313.3
R3497 V_OSC.n3 V_OSC.t2 257.067
R3498 V_OSC.n1 V_OSC.t0 247.934
R3499 V_OSC.n2 V_OSC.n1 236.756
R3500 V_OSC.n0 V_OSC.t6 224.934
R3501 V_OSC.n2 V_OSC.n0 224.934
R3502 V_OSC.n0 V_OSC.t4 144.601
R3503 V_OSC V_OSC.n2 120.501
R3504 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t1 755.534
R3505 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 685.134
R3506 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 389.733
R3507 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t0 340.2
R3508 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t3 321.334
R3509 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.A.t4 144.601
R3510 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.A.n1 19.2005
R3511 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.C.t1 96.0005
R3512 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R3513 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R3514 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R3515 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R3516 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R3517 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R3518 pfd_8_0.E.t0 pfd_8_0.E.n4 221.411
R3519 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R3520 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R3521 pfd_8_0.E.n1 pfd_8_0.E.t2 24.0005
R3522 pfd_8_0.E.n1 pfd_8_0.E.t1 24.0005
R3523 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R3524 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R3525 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R3526 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R3527 pfd_8_0.E_b.t1 pfd_8_0.E_b.n2 221.411
R3528 pfd_8_0.E_b.n1 pfd_8_0.E_b.t0 24.0005
R3529 pfd_8_0.E_b.n1 pfd_8_0.E_b.t2 24.0005
R3530 a_1390_1400.t0 a_1390_1400.t1 39.4005
R3531 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R3532 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R3533 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R3534 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R3535 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R3536 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R3537 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R3538 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t0 221.411
R3539 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t1 24.0005
R3540 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R3541 a_870_640.t0 a_870_640.t1 39.4005
R3542 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.F.t1 157.601
R3543 a_2530_190.t1 a_2530_190.n2 500.086
R3544 a_2530_190.n0 a_2530_190.t2 465.933
R3545 a_2530_190.t1 a_2530_190.n2 461.389
R3546 a_2530_190.n1 a_2530_190.n0 392.623
R3547 a_2530_190.n0 a_2530_190.t3 321.334
R3548 a_2530_190.n1 a_2530_190.t0 177.577
R3549 a_2530_190.n2 a_2530_190.n1 48.3899
R3550 a_2200_190.t1 a_2200_190.n2 500.086
R3551 a_2200_190.n1 a_2200_190.n0 473.334
R3552 a_2200_190.n0 a_2200_190.t2 465.933
R3553 a_2200_190.t1 a_2200_190.n2 461.389
R3554 a_2200_190.n0 a_2200_190.t3 321.334
R3555 a_2200_190.n1 a_2200_190.t0 177.577
R3556 a_2200_190.n2 a_2200_190.n1 48.3898
R3557 loop_filter_2_0.R1_C1.t0 loop_filter_2_0.R1_C1.t1 167.429
R3558 a_9360_3514.t1 a_9360_3514.t0 323.964
R3559 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t1 663.801
R3560 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 397.053
R3561 VCO_FD_magic_0.div120_2_0.div5_2_0.B.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.B.t2 348.851
R3562 VCO_FD_magic_0.vco2_3_0.V9.n1 VCO_FD_magic_0.vco2_3_0.V9.n0 437.733
R3563 VCO_FD_magic_0.vco2_3_0.V9.t1 VCO_FD_magic_0.vco2_3_0.V9.n1 372.118
R3564 VCO_FD_magic_0.vco2_3_0.V9.n1 VCO_FD_magic_0.vco2_3_0.V9.t0 247.934
R3565 VCO_FD_magic_0.vco2_3_0.V9.n0 VCO_FD_magic_0.vco2_3_0.V9.t2 224.934
R3566 VCO_FD_magic_0.vco2_3_0.V9.n0 VCO_FD_magic_0.vco2_3_0.V9.t3 144.601
R3567 VCO_FD_magic_0.vco2_3_0.V8.n1 VCO_FD_magic_0.vco2_3_0.V8.n0 437.733
R3568 VCO_FD_magic_0.vco2_3_0.V8.t1 VCO_FD_magic_0.vco2_3_0.V8.n1 372.118
R3569 VCO_FD_magic_0.vco2_3_0.V8.n1 VCO_FD_magic_0.vco2_3_0.V8.t0 247.934
R3570 VCO_FD_magic_0.vco2_3_0.V8.n0 VCO_FD_magic_0.vco2_3_0.V8.t3 224.934
R3571 VCO_FD_magic_0.vco2_3_0.V8.n0 VCO_FD_magic_0.vco2_3_0.V8.t2 144.601
R3572 VCO_FD_magic_0.vco2_3_0.V3.n0 VCO_FD_magic_0.vco2_3_0.V3.t0 284.2
R3573 VCO_FD_magic_0.vco2_3_0.V3.n0 VCO_FD_magic_0.vco2_3_0.V3.t2 233
R3574 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V3.t1 162.857
R3575 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V3.n0 21.3338
R3576 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R3577 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R3578 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R3579 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R3580 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R3581 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R3582 pfd_8_0.F.t0 pfd_8_0.F.n4 221.411
R3583 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R3584 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R3585 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R3586 pfd_8_0.F.n1 pfd_8_0.F.t1 24.0005
R3587 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.D.t3 742.201
R3588 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t4 350.349
R3589 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t0 254.333
R3590 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 206.333
R3591 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n1 70.4005
R3592 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t2 48.0005
R3593 VCO_FD_magic_0.div120_2_0.div5_2_0.D.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.D.t1 48.0005
R3594 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.D.n2 19.2005
R3595 VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t1 713.933
R3596 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.A.t0 327.401
R3597 VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_1.A.t2 314.233
R3598 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.A.n0 9.6005
R3599 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_1.B.t1 96.0005
R3600 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.G.t1 96.0005
R3601 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.M.t0 739
R3602 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t4 349.433
R3603 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t2 254.333
R3604 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 206.333
R3605 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n1 70.4005
R3606 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t3 48.0005
R3607 VCO_FD_magic_0.div120_2_0.div5_2_0.M.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.M.t1 48.0005
R3608 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.M.n2 22.4005
R3609 a_9360_6440.t1 a_9360_6440.t0 245.883
R3610 VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t0 713.933
R3611 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.A.t1 327.401
R3612 VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 VCO_FD_magic_0.div120_2_0.div2_4_0.A.t2 314.233
R3613 VCO_FD_magic_0.div120_2_0.div2_4_0.A VCO_FD_magic_0.div120_2_0.div2_4_0.A.n0 9.6005
R3614 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R3615 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R3616 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R3617 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R3618 pfd_8_0.F_b.t1 pfd_8_0.F_b.n2 221.411
R3619 pfd_8_0.F_b.n1 pfd_8_0.F_b.t0 24.0005
R3620 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R3621 a_1390_640.t0 a_1390_640.t1 39.4005
R3622 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t0 VCO_FD_magic_0.div120_2_0.div5_2_0.L.t1 96.0005
R3623 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t1 685.134
R3624 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t2 663.801
R3625 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t3 534.268
R3626 VCO_FD_magic_0.div120_2_0.div3_3_0.E.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 362.921
R3627 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n1 VCO_FD_magic_0.div120_2_0.div3_3_0.E.n0 91.7338
R3628 VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t1 663.801
R3629 VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.K.t2 355.378
R3630 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.K.t0 276.521
R3631 VCO_FD_magic_0.div120_2_0.div5_2_0.K VCO_FD_magic_0.div120_2_0.div5_2_0.K.n0 120.534
R3632 a_490_640.t0 a_490_640.t1 39.4005
R3633 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t0 VCO_FD_magic_0.div120_2_0.div2_4_0.B.t1 96.0005
R3634 VCO_FD_magic_0.vco2_3_0.V7.n0 VCO_FD_magic_0.vco2_3_0.V7.t0 284.2
R3635 VCO_FD_magic_0.vco2_3_0.V7.n0 VCO_FD_magic_0.vco2_3_0.V7.t2 233
R3636 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V7.t1 162.857
R3637 VCO_FD_magic_0.vco2_3_0.V7 VCO_FD_magic_0.vco2_3_0.V7.n0 21.3338
R3638 VCO_FD_magic_0.vco2_3_0.V5.n0 VCO_FD_magic_0.vco2_3_0.V5.t2 284.2
R3639 VCO_FD_magic_0.vco2_3_0.V5.n0 VCO_FD_magic_0.vco2_3_0.V5.t1 233
R3640 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V5.t0 162.857
R3641 VCO_FD_magic_0.vco2_3_0.V5 VCO_FD_magic_0.vco2_3_0.V5.n0 21.3338
R3642 VCO_FD_magic_0.vco2_3_0.V2.n0 VCO_FD_magic_0.vco2_3_0.V2.t0 421.027
R3643 VCO_FD_magic_0.vco2_3_0.V2.n0 VCO_FD_magic_0.vco2_3_0.V2.t2 348.81
R3644 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V2.t1 284.317
R3645 VCO_FD_magic_0.vco2_3_0.V2 VCO_FD_magic_0.vco2_3_0.V2.n0 31.8427
R3646 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t0 723
R3647 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t2 514.134
R3648 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t3 332.783
R3649 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 VCO_FD_magic_0.div120_2_0.div5_2_0.E.t1 314.921
R3650 VCO_FD_magic_0.div120_2_0.div5_2_0.E VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 6.4005
R3651 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n1 VCO_FD_magic_0.div120_2_0.div5_2_0.E.n0 3.2005
R3652 a_490_1400.t0 a_490_1400.t1 39.4005
R3653 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R3654 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R3655 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R3656 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R3657 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R3658 pfd_8_0.Reset.t0 pfd_8_0.Reset.n3 288.37
R3659 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R3660 pfd_8_0.Reset.n3 pfd_8_0.Reset.t1 177.577
R3661 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R3662 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.B.t1 96.0005
R3663 a_1870_190.t1 a_1870_190.n2 500.086
R3664 a_1870_190.n1 a_1870_190.n0 473.334
R3665 a_1870_190.n0 a_1870_190.t2 465.933
R3666 a_1870_190.t1 a_1870_190.n2 461.389
R3667 a_1870_190.n0 a_1870_190.t3 321.334
R3668 a_1870_190.n1 a_1870_190.t0 177.577
R3669 a_1870_190.n2 a_1870_190.n1 48.3898
R3670 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t0 713.933
R3671 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t2 314.233
R3672 VCO_FD_magic_0.div120_2_0.div3_3_0.A.t1 VCO_FD_magic_0.div120_2_0.div3_3_0.A.n0 308.2
R3673 VCO_FD_magic_0.vco2_3_0.V6.n0 VCO_FD_magic_0.vco2_3_0.V6.t0 421.027
R3674 VCO_FD_magic_0.vco2_3_0.V6.n0 VCO_FD_magic_0.vco2_3_0.V6.t2 348.81
R3675 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V6.t1 280.05
R3676 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V6.n0 36.1094
R3677 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t0 VCO_FD_magic_0.div120_2_0.div3_3_0.F.t1 96.0005
R3678 a_n30_640.t0 a_n30_640.t1 39.4005
C0 VDDA VCO_FD_magic_0.div120_2_0.div2_4_1.A 0.126015f
C1 VCO_FD_magic_0.div120_2_0.div2_4_0.C VDDA 0.111144f
C2 VCO_FD_magic_0.vco2_3_0.V4 VDDA 0.413959f
C3 pfd_8_0.QA_b F_REF 0.027208f
C4 VCO_FD_magic_0.div120_2_0.div2_4_2.A VCO_FD_magic_0.div120_2_0.div2_4_2.C 0.122602f
C5 VDDA VCO_FD_magic_0.vco2_3_0.V7 0.033517f
C6 VDDA F_REF 0.098433f
C7 VCO_FD_magic_0.vco2_3_0.V3 V_OSC 0.046941f
C8 VCO_FD_magic_0.div120_2_0.div2_4_0.C VCO_FD_magic_0.div120_2_0.div2_4_0.A 0.122602f
C9 VCO_FD_magic_0.vco2_3_0.V3 VCO_FD_magic_0.vco2_3_0.V2 0.010316f
C10 VCO_FD_magic_0.div120_2_0.div5_2_0.G F_VCO 0.081976f
C11 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN+ 0.100967f
C12 VCO_FD_magic_0.div120_2_0.div5_2_0.D VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.070599f
C13 I_IN pfd_8_0.DOWN_input 0.928029f
C14 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.H 0.106696f
C15 VCO_FD_magic_0.div120_2_0.div5_2_0.D VDDA 0.144695f
C16 VCO_FD_magic_0.vco2_3_0.V6 VDDA 0.281338f
C17 opamp_cell_4_0.VIN+ pfd_8_0.DOWN_input 0.080549f
C18 pfd_8_0.QB_b F_VCO 0.044529f
C19 VDDA opamp_cell_4_0.p_bias 2.86573f
C20 V_OSC VCO_FD_magic_0.vco2_3_0.V2 0.063469f
C21 VDDA VCO_FD_magic_0.div120_2_0.div2_4_1.C 0.111409f
C22 V_OSC VCO_FD_magic_0.vco2_3_0.V5 0.017652f
C23 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.I 0.069172f
C24 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.112235f
C25 VDDA pfd_8_0.DOWN_input 0.221484f
C26 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.061186f
C27 VCO_FD_magic_0.vco2_3_0.V3 VDDA 0.040599f
C28 VCO_FD_magic_0.div120_2_0.div5_2_0.G VDDA 0.25905f
C29 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.D 0.163145f
C30 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div3_3_0.H 0.038583f
C31 VDDA VCO_FD_magic_0.div120_2_0.div2_4_2.C 0.111144f
C32 VCO_FD_magic_0.div120_2_0.div3_3_0.C VCO_FD_magic_0.div120_2_0.div3_3_0.D 0.060684f
C33 VDDA VCO_FD_magic_0.div120_2_0.div3_3_0.D 0.311052f
C34 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.K 0.174679f
C35 VCO_FD_magic_0.div120_2_0.div2_4_2.A VDDA 0.125335f
C36 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.M 0.119081f
C37 pfd_8_0.QB_b VDDA 0.512673f
C38 VCO_FD_magic_0.div120_2_0.div5_2_0.M VCO_FD_magic_0.div120_2_0.div5_2_0.K 0.169071f
C39 V_OSC VDDA 0.627267f
C40 VCO_FD_magic_0.div120_2_0.div5_2_0.G VCO_FD_magic_0.div120_2_0.div24 0.240642f
C41 pfd_8_0.QB_b pfd_8_0.QB 0.388258f
C42 VCO_FD_magic_0.vco2_3_0.V6 VCO_FD_magic_0.vco2_3_0.V7 0.010316f
C43 VCO_FD_magic_0.div120_2_0.div2_4_1.A VCO_FD_magic_0.div120_2_0.div2_4_1.C 0.122602f
C44 VCO_FD_magic_0.div120_2_0.div5_2_0.I F_VCO 0.021863f
C45 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.139506f
C46 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div3_3_0.D 0.024014f
C47 VCO_FD_magic_0.vco2_3_0.V2 VDDA 0.410554f
C48 I_IN opamp_cell_4_0.VIN+ 0.166322f
C49 F_VCO VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.036046f
C50 F_VCO VDDA 1.25401f
C51 VDDA VCO_FD_magic_0.vco2_3_0.V5 0.040599f
C52 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C53 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.K 0.482256f
C54 F_VCO pfd_8_0.QB 0.060952f
C55 VDDA pfd_8_0.QA 0.550605f
C56 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.M 0.157966f
C57 I_IN VDDA 0.541032f
C58 pfd_8_0.QA pfd_8_0.QB 0.074487f
C59 VDDA opamp_cell_4_0.VIN+ 0.832915f
C60 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.021344f
C61 VCO_FD_magic_0.div120_2_0.div24 F_VCO 0.067501f
C62 VCO_FD_magic_0.div120_2_0.div5_2_0.I VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.016448f
C63 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.53342f
C64 pfd_8_0.QA_b VDDA 0.52066f
C65 VCO_FD_magic_0.div120_2_0.div3_3_0.C VDDA 0.125686f
C66 VDDA VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.104998f
C67 V_OSC VCO_FD_magic_0.vco2_3_0.V7 0.108092f
C68 VDDA pfd_8_0.QB 2.75013f
C69 VCO_FD_magic_0.vco2_3_0.V4 VCO_FD_magic_0.vco2_3_0.V5 0.010316f
C70 VCO_FD_magic_0.div120_2_0.div2_4_0.A VDDA 0.125335f
C71 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.I 0.076865f
C72 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.E 0.108607f
C73 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div3_3_0.C 0.03648f
C74 VCO_FD_magic_0.div120_2_0.div24 VCO_FD_magic_0.div120_2_0.div5_2_0.J 0.176046f
C75 VCO_FD_magic_0.div120_2_0.div24 VDDA 0.654009f
C76 F_REF pfd_8_0.QA 0.056f
C77 VCO_FD_magic_0.vco2_3_0.V6 V_OSC 0.019495f
C78 V_OSC GNDA 2.90637f
C79 I_IN GNDA 2.82399f
C80 F_REF GNDA 0.277742f
C81 VDDA GNDA 71.3612f
C82 VCO_FD_magic_0.vco2_3_0.V2 GNDA 0.045471f
C83 VCO_FD_magic_0.vco2_3_0.V4 GNDA 0.045471f
C84 VCO_FD_magic_0.vco2_3_0.V6 GNDA 0.157087f
C85 VCO_FD_magic_0.div120_2_0.div2_4_1.A GNDA 0.200071f
C86 VCO_FD_magic_0.div120_2_0.div2_4_2.A GNDA 0.200074f
C87 VCO_FD_magic_0.div120_2_0.div2_4_0.A GNDA 0.200071f
C88 VCO_FD_magic_0.div120_2_0.div5_2_0.G GNDA 0.195152f
C89 VCO_FD_magic_0.div120_2_0.div5_2_0.I GNDA 0.152847f
C90 VCO_FD_magic_0.div120_2_0.div3_3_0.C GNDA 0.36191f
C91 VCO_FD_magic_0.div120_2_0.div3_3_0.D GNDA 0.301961f
C92 VCO_FD_magic_0.div120_2_0.div3_3_0.H GNDA 0.423425f
C93 VCO_FD_magic_0.div120_2_0.div5_2_0.D GNDA 0.366928f
C94 VCO_FD_magic_0.div120_2_0.div5_2_0.E GNDA 0.297109f
C95 VCO_FD_magic_0.div120_2_0.div5_2_0.J GNDA 0.398061f
C96 VCO_FD_magic_0.div120_2_0.div5_2_0.K GNDA 0.180033f
C97 VCO_FD_magic_0.div120_2_0.div5_2_0.M GNDA 0.397035f
C98 VCO_FD_magic_0.div120_2_0.div2_4_1.C GNDA 0.45763f
C99 VCO_FD_magic_0.div120_2_0.div2_4_2.C GNDA 0.457627f
C100 VCO_FD_magic_0.div120_2_0.div2_4_0.C GNDA 0.46146f
C101 VCO_FD_magic_0.div120_2_0.div24 GNDA 3.78529f
C102 VCO_FD_magic_0.vco2_3_0.V3 GNDA 0.300759f
C103 VCO_FD_magic_0.vco2_3_0.V5 GNDA 0.302737f
C104 VCO_FD_magic_0.vco2_3_0.V7 GNDA 0.314921f
C105 pfd_8_0.DOWN_input GNDA 3.02729f
C106 pfd_8_0.QB_b GNDA 1.04775f
C107 F_VCO GNDA 3.25572f
C108 pfd_8_0.QB GNDA 1.307779f
C109 pfd_8_0.QA GNDA 3.10102f
C110 pfd_8_0.QA_b GNDA 1.05138f
C111 opamp_cell_4_0.VIN+ GNDA 2.37749f
C112 opamp_cell_4_0.p_bias GNDA 3.954681f
C113 loop_filter_2_0.R1_C1.t1 GNDA 2.39887f
C114 pfd_8_0.QB.t7 GNDA 0.069179f
C115 pfd_8_0.QB.t8 GNDA 0.032493f
C116 pfd_8_0.QB.n0 GNDA 0.099932f
C117 pfd_8_0.QB.t3 GNDA 0.069179f
C118 pfd_8_0.QB.t4 GNDA 0.104293f
C119 pfd_8_0.QB.n1 GNDA 1.25065f
C120 pfd_8_0.QB.t5 GNDA 0.069862f
C121 pfd_8_0.QB.t6 GNDA 0.030633f
C122 pfd_8_0.QB.n2 GNDA 0.176466f
C123 pfd_8_0.QB.t2 GNDA 0.147114f
C124 pfd_8_0.QB.t0 GNDA 0.027951f
C125 pfd_8_0.QB.t1 GNDA 0.027951f
C126 pfd_8_0.QB.n3 GNDA 0.149246f
C127 pfd_8_0.QB.n4 GNDA 0.265156f
C128 pfd_8_0.QB.n5 GNDA 0.226459f
C129 opamp_cell_4_0.p_bias.t8 GNDA 1.66267f
C130 opamp_cell_4_0.p_bias.t1 GNDA 0.019693f
C131 opamp_cell_4_0.p_bias.t5 GNDA 0.019693f
C132 opamp_cell_4_0.p_bias.n0 GNDA 0.054067f
C133 opamp_cell_4_0.p_bias.t7 GNDA 0.019693f
C134 opamp_cell_4_0.p_bias.t3 GNDA 0.019693f
C135 opamp_cell_4_0.p_bias.n1 GNDA 0.054067f
C136 opamp_cell_4_0.p_bias.n2 GNDA 0.068502f
C137 opamp_cell_4_0.p_bias.t0 GNDA 0.054353f
C138 opamp_cell_4_0.p_bias.t2 GNDA 0.054353f
C139 opamp_cell_4_0.p_bias.t6 GNDA 0.054353f
C140 opamp_cell_4_0.p_bias.t11 GNDA 0.054353f
C141 opamp_cell_4_0.p_bias.t9 GNDA 0.074733f
C142 opamp_cell_4_0.p_bias.n3 GNDA 0.04185f
C143 opamp_cell_4_0.p_bias.n4 GNDA 0.029697f
C144 opamp_cell_4_0.p_bias.n5 GNDA 0.012761f
C145 opamp_cell_4_0.p_bias.n6 GNDA 0.029697f
C146 opamp_cell_4_0.p_bias.n7 GNDA 0.029697f
C147 opamp_cell_4_0.p_bias.t4 GNDA 0.054353f
C148 opamp_cell_4_0.p_bias.t12 GNDA 0.054353f
C149 opamp_cell_4_0.p_bias.t10 GNDA 0.074733f
C150 opamp_cell_4_0.p_bias.n8 GNDA 0.04185f
C151 opamp_cell_4_0.p_bias.n9 GNDA 0.029697f
C152 opamp_cell_4_0.p_bias.n10 GNDA 0.012761f
C153 opamp_cell_4_0.p_bias.n11 GNDA 0.120625f
C154 pfd_8_0.opamp_out.t12 GNDA 0.957954f
C155 pfd_8_0.opamp_out.t11 GNDA 0.957546f
C156 pfd_8_0.opamp_out.n6 GNDA 0.012958f
C157 pfd_8_0.opamp_out.t14 GNDA 0.012873f
C158 pfd_8_0.opamp_out.t2 GNDA 0.012026f
C159 pfd_8_0.opamp_out.n13 GNDA 0.015342f
C160 pfd_8_0.opamp_out.n14 GNDA 0.081091f
C161 pfd_8_0.opamp_out.n15 GNDA 0.047633f
C162 VCO_FD_magic_0.vco2_3_0.V1.t1 GNDA 0.104706f
C163 VCO_FD_magic_0.vco2_3_0.V1.n0 GNDA 0.184398f
C164 VCO_FD_magic_0.vco2_3_0.V1.t4 GNDA 0.298444f
C165 VCO_FD_magic_0.vco2_3_0.V1.t3 GNDA 0.298444f
C166 VCO_FD_magic_0.vco2_3_0.V1.t5 GNDA 0.497217f
C167 VCO_FD_magic_0.vco2_3_0.V1.n1 GNDA 0.243367f
C168 VCO_FD_magic_0.vco2_3_0.V1.n2 GNDA 0.217957f
C169 VCO_FD_magic_0.vco2_3_0.V1.t0 GNDA 0.298444f
C170 VCO_FD_magic_0.vco2_3_0.V1.n3 GNDA 0.169192f
C171 VCO_FD_magic_0.vco2_3_0.V1.n4 GNDA 0.045341f
C172 VCO_FD_magic_0.vco2_3_0.V1.n5 GNDA 0.177452f
C173 VCO_FD_magic_0.vco2_3_0.V1.t2 GNDA 0.165036f
C174 VDDA.n71 GNDA 0.051784f
C175 VDDA.t36 GNDA 0.173447f
C176 VDDA.n74 GNDA 0.115632f
C177 VDDA.n80 GNDA 0.01246f
C178 VDDA.n86 GNDA 0.014434f
C179 VDDA.n87 GNDA 0.03888f
C180 VDDA.t219 GNDA 0.089652f
C181 VDDA.t129 GNDA 0.070664f
C182 VDDA.t81 GNDA 0.033245f
C183 VDDA.n90 GNDA 0.014698f
C184 VDDA.t12 GNDA 0.015182f
C185 VDDA.t44 GNDA 0.025751f
C186 VDDA.t14 GNDA 0.025751f
C187 VDDA.t120 GNDA 0.016911f
C188 VDDA.t8 GNDA 0.016911f
C189 VDDA.t58 GNDA 0.028057f
C190 VDDA.t136 GNDA 0.029018f
C191 VDDA.n91 GNDA 0.014698f
C192 VDDA.t85 GNDA 0.015182f
C193 VDDA.t201 GNDA 0.017295f
C194 VDDA.t116 GNDA 0.017295f
C195 VDDA.t114 GNDA 0.013836f
C196 VDDA.t93 GNDA 0.013836f
C197 VDDA.t142 GNDA 0.022292f
C198 VDDA.t24 GNDA 0.022292f
C199 VDDA.t10 GNDA 0.016911f
C200 VDDA.t146 GNDA 0.016911f
C201 VDDA.t199 GNDA 0.023829f
C202 VDDA.t194 GNDA 0.02479f
C203 VDDA.n92 GNDA 0.011623f
C204 VDDA.t130 GNDA 0.012107f
C205 VDDA.t73 GNDA 0.013836f
C206 VDDA.t75 GNDA 0.013836f
C207 VDDA.t95 GNDA 0.02306f
C208 VDDA.t197 GNDA 0.024021f
C209 VDDA.n94 GNDA 0.011623f
C210 VDDA.t56 GNDA 0.012107f
C211 VDDA.t38 GNDA 0.013836f
C212 VDDA.t65 GNDA 0.013836f
C213 VDDA.t54 GNDA 0.02306f
C214 VDDA.t40 GNDA 0.024021f
C215 VDDA.n95 GNDA 0.011623f
C216 VDDA.t22 GNDA 0.012107f
C217 VDDA.t207 GNDA 0.013836f
C218 VDDA.t126 GNDA 0.013836f
C219 VDDA.t0 GNDA 0.02306f
C220 VDDA.t210 GNDA 0.024021f
C221 VDDA.n97 GNDA 0.011623f
C222 VDDA.t6 GNDA 0.012107f
C223 VDDA.t112 GNDA 0.013836f
C224 VDDA.t33 GNDA 0.013836f
C225 VDDA.t2 GNDA 0.0214f
C226 VDDA.t48 GNDA 0.100683f
C227 VDDA.t144 GNDA 0.089652f
C228 VDDA.n99 GNDA 0.038136f
C229 VDDA.n108 GNDA 0.099572f
C230 VDDA.t135 GNDA 0.070664f
C231 VDDA.t99 GNDA 0.089652f
C232 VDDA.n110 GNDA 0.038136f
C233 VDDA.n116 GNDA 0.099572f
C234 VDDA.n128 GNDA 0.05312f
C235 VDDA.n129 GNDA 0.039691f
C236 VDDA.n300 GNDA 0.093595f
C237 VDDA.t27 GNDA 0.030637f
C238 VDDA.t125 GNDA 0.011111f
C239 VDDA.n324 GNDA 0.012169f
C240 VDDA.t212 GNDA 0.030637f
C241 VDDA.n341 GNDA 0.028191f
C242 VDDA.n344 GNDA 0.010981f
C243 VDDA.t192 GNDA 0.10326f
C244 VDDA.n350 GNDA 0.010981f
C245 VDDA.n351 GNDA 0.010981f
C246 VDDA.n379 GNDA 0.010229f
C247 VDDA.n387 GNDA 0.050308f
C248 VDDA.t176 GNDA 0.123217f
C249 VDDA.t16 GNDA 0.062336f
C250 VDDA.t148 GNDA 0.062336f
C251 VDDA.t69 GNDA 0.062336f
C252 VDDA.t122 GNDA 0.062336f
C253 VDDA.t182 GNDA 0.070728f
C254 VDDA.n392 GNDA 0.013768f
C255 VDDA.t164 GNDA 0.018131f
C256 VDDA.n397 GNDA 0.013726f
C257 VDDA.n407 GNDA 0.099498f
C258 VDDA.t155 GNDA 0.047951f
C259 VDDA.t165 GNDA 0.031168f
C260 VDDA.t153 GNDA 0.037162f
C261 VDDA.t154 GNDA 0.041957f
C262 VDDA.t71 GNDA 0.031168f
C263 VDDA.t49 GNDA 0.047951f
C264 VDDA.t97 GNDA 0.031168f
C265 VDDA.t62 GNDA 0.034764f
C266 VDDA.t156 GNDA 0.044355f
C267 VDDA.t108 GNDA 0.061138f
C268 VDDA.t29 GNDA 0.064734f
C269 VDDA.n408 GNDA 0.051668f
C270 VDDA.t20 GNDA 0.03956f
C271 VDDA.t161 GNDA 0.03956f
C272 VDDA.t52 GNDA 0.03956f
C273 VDDA.t140 GNDA 0.031168f
C274 VDDA.t79 GNDA 0.047951f
C275 VDDA.t18 GNDA 0.031168f
C276 VDDA.t50 GNDA 0.037162f
C277 VDDA.t215 GNDA 0.041957f
C278 VDDA.t138 GNDA 0.031168f
C279 VDDA.t158 GNDA 0.047951f
C280 VDDA.t169 GNDA 0.03956f
C281 VDDA.n412 GNDA 0.016359f
C282 VDDA.n413 GNDA 0.046733f
C283 VDDA.t168 GNDA 0.018502f
C284 VDDA.n416 GNDA 0.013726f
C285 VDDA.n423 GNDA 0.012928f
C286 VDDA.n425 GNDA 0.037812f
C287 VDDA.n426 GNDA 0.045674f
C288 VDDA.n427 GNDA 0.013768f
C289 VDDA.n430 GNDA 0.011329f
C290 VDDA.n431 GNDA 0.032916f
C291 VDDA.n432 GNDA 0.033073f
C292 VDDA.n440 GNDA 0.032073f
C293 VDDA.n447 GNDA 0.032073f
C294 VDDA.n454 GNDA 0.032073f
C295 VDDA.n461 GNDA 0.032073f
C296 VDDA.n471 GNDA 0.021537f
C297 VDDA.n475 GNDA 0.010981f
C298 VDDA.t172 GNDA 0.045645f
C299 VDDA.n482 GNDA 0.010249f
C300 VDDA.n485 GNDA 0.010249f
C301 VDDA.n488 GNDA 0.010584f
C302 VDDA.n489 GNDA 0.014893f
C303 VDDA.n491 GNDA 0.010584f
C304 VDDA.n492 GNDA 0.014893f
C305 VDDA.n511 GNDA 0.010584f
C306 VDDA.n514 GNDA 0.010584f
C307 VDDA.t178 GNDA 0.018245f
C308 VDDA.t77 GNDA 0.046707f
C309 VDDA.t203 GNDA 0.046707f
C310 VDDA.t60 GNDA 0.046707f
C311 VDDA.t87 GNDA 0.046707f
C312 VDDA.t179 GNDA 0.045645f
C313 VDDA.n525 GNDA 0.041399f
C314 VDDA.n530 GNDA 0.010981f
C315 VDDA.n531 GNDA 0.010584f
C316 VDDA.n532 GNDA 0.015082f
C317 VDDA.n539 GNDA 0.014161f
C318 VDDA.n546 GNDA 0.014893f
C319 VDDA.n554 GNDA 0.014893f
C320 VDDA.n555 GNDA 0.010584f
C321 VDDA.n556 GNDA 0.010981f
C322 VDDA.t171 GNDA 0.017216f
C323 VDDA.t185 GNDA 0.017216f
C324 VDDA.n559 GNDA 0.013217f
C325 VDDA.n560 GNDA 0.010981f
C326 VDDA.n561 GNDA 0.012452f
C327 VDDA.n563 GNDA 0.044583f
C328 VDDA.t186 GNDA 0.045645f
C329 VDDA.t217 GNDA 0.046707f
C330 VDDA.t89 GNDA 0.046707f
C331 VDDA.t91 GNDA 0.046707f
C332 VDDA.t118 GNDA 0.046707f
C333 VDDA.t189 GNDA 0.045645f
C334 VDDA.n569 GNDA 0.041399f
C335 VDDA.t188 GNDA 0.018245f
C336 VDDA.n579 GNDA 0.014987f
C337 VDDA.n580 GNDA 0.156827f
C338 VDDA.n581 GNDA 0.028105f
C339 VDDA.n583 GNDA 0.010981f
C340 VDDA.t46 GNDA 0.107798f
C341 VDDA.t107 GNDA 0.116876f
C342 VDDA.n590 GNDA 0.088508f
C343 VDDA.n614 GNDA 0.088508f
C344 VDDA.t104 GNDA 0.088508f
C345 VDDA.t205 GNDA 0.030637f
C346 VDDA.n627 GNDA 0.044254f
C347 VDDA.n635 GNDA 0.044254f
C348 VDDA.t83 GNDA 0.030637f
C349 VDDA.t63 GNDA 0.030637f
C350 VDDA.n643 GNDA 0.06241f
C351 VDDA.n646 GNDA 0.010981f
C352 VDDA.n655 GNDA 0.010981f
C353 VDDA.n663 GNDA 0.096451f
C354 VDDA.t67 GNDA 0.088508f
C355 VDDA.n669 GNDA 0.088508f
C356 VDDA.n705 GNDA 0.044254f
C357 VDDA.t42 GNDA 0.027233f
C358 VDDA.t124 GNDA 0.028368f
C359 VDDA.n711 GNDA 0.044254f
C360 VDDA.n727 GNDA 0.06014f
C361 VDDA.n746 GNDA 0.066949f
C362 VDDA.t110 GNDA 0.055601f
C363 VDDA.t26 GNDA 0.118011f
C364 VDDA.t128 GNDA 0.118011f
C365 VDDA.t101 GNDA 0.055601f
C366 VDDA.n770 GNDA 0.061275f
C367 VDDA.t133 GNDA 0.055601f
C368 VDDA.t9 GNDA 0.118011f
C369 VDDA.t35 GNDA 0.118011f
C370 VDDA.t4 GNDA 0.055601f
C371 VDDA.n783 GNDA 0.06241f
C372 VDDA.n818 GNDA 0.082395f
C373 a_5970_4630.t11 GNDA 0.030769f
C374 a_5970_4630.n0 GNDA 0.124795f
C375 a_5970_4630.t2 GNDA 0.020325f
C376 a_5970_4630.t1 GNDA 0.020325f
C377 a_5970_4630.t7 GNDA 0.020325f
C378 a_5970_4630.n1 GNDA 0.044943f
C379 a_5970_4630.t6 GNDA 0.020325f
C380 a_5970_4630.t9 GNDA 0.020325f
C381 a_5970_4630.n2 GNDA 0.044943f
C382 a_5970_4630.t10 GNDA 0.077457f
C383 a_5970_4630.t8 GNDA 0.030769f
C384 a_5970_4630.n3 GNDA 0.097952f
C385 a_5970_4630.n4 GNDA 0.087903f
C386 a_5970_4630.n5 GNDA 0.089425f
C387 a_5970_4630.t5 GNDA 0.050813f
C388 a_5970_4630.t0 GNDA 0.050813f
C389 a_5970_4630.n6 GNDA 0.295522f
C390 a_5970_4630.t4 GNDA 0.050813f
C391 a_5970_4630.t3 GNDA 0.050813f
C392 a_5970_4630.n7 GNDA 0.144587f
C393 a_5970_4630.n8 GNDA 0.360746f
C394 a_5970_4630.n9 GNDA 0.13437f
C395 a_5970_4630.n10 GNDA 0.085474f
C396 a_5970_4630.n11 GNDA 0.045257f
C397 a_5970_4630.t12 GNDA 0.100208f
C398 V_CONT.n2 GNDA 0.013537f
C399 V_CONT.n5 GNDA 0.01164f
C400 V_CONT.n8 GNDA 0.078062f
C401 V_CONT.t5 GNDA 4.34239f
C402 V_CONT.n9 GNDA 0.031107f
C403 V_CONT.n15 GNDA 0.037822f
C404 opamp_cell_4_0.VIN- GNDA 0.020154f
.ends

