magic
tech sky130A
timestamp 1739895002
<< nwell >>
rect 605 150 1145 255
<< nmos >>
rect 665 -35 680 15
rect 720 -35 735 15
rect 775 -35 790 15
rect 940 -35 955 15
rect 995 -35 1010 15
rect 1050 -35 1065 15
rect 1105 -35 1120 15
<< pmos >>
rect 665 170 680 220
rect 720 170 735 220
rect 845 170 860 220
rect 900 170 915 220
rect 1070 170 1085 220
<< ndiff >>
rect 625 0 665 15
rect 625 -20 635 0
rect 655 -20 665 0
rect 625 -35 665 -20
rect 680 0 720 15
rect 680 -20 690 0
rect 710 -20 720 0
rect 680 -35 720 -20
rect 735 0 775 15
rect 735 -20 745 0
rect 765 -20 775 0
rect 735 -35 775 -20
rect 790 0 830 15
rect 790 -20 800 0
rect 820 -20 830 0
rect 790 -35 830 -20
rect 900 0 940 15
rect 900 -20 910 0
rect 930 -20 940 0
rect 900 -35 940 -20
rect 955 0 995 15
rect 955 -20 965 0
rect 985 -20 995 0
rect 955 -35 995 -20
rect 1010 0 1050 15
rect 1010 -20 1020 0
rect 1040 -20 1050 0
rect 1010 -35 1050 -20
rect 1065 0 1105 15
rect 1065 -20 1075 0
rect 1095 -20 1105 0
rect 1065 -35 1105 -20
rect 1120 0 1160 15
rect 1120 -20 1130 0
rect 1150 -20 1160 0
rect 1120 -35 1160 -20
<< pdiff >>
rect 625 205 665 220
rect 625 185 635 205
rect 655 185 665 205
rect 625 170 665 185
rect 680 205 720 220
rect 680 185 690 205
rect 710 185 720 205
rect 680 170 720 185
rect 735 205 775 220
rect 735 185 745 205
rect 765 185 775 205
rect 735 170 775 185
rect 805 205 845 220
rect 805 185 815 205
rect 835 185 845 205
rect 805 170 845 185
rect 860 205 900 220
rect 860 185 870 205
rect 890 185 900 205
rect 860 170 900 185
rect 915 205 955 220
rect 915 185 925 205
rect 945 185 955 205
rect 915 170 955 185
rect 1030 205 1070 220
rect 1030 185 1040 205
rect 1060 185 1070 205
rect 1030 170 1070 185
rect 1085 205 1125 220
rect 1085 185 1095 205
rect 1115 185 1125 205
rect 1085 170 1125 185
<< ndiffc >>
rect 635 -20 655 0
rect 690 -20 710 0
rect 745 -20 765 0
rect 800 -20 820 0
rect 910 -20 930 0
rect 965 -20 985 0
rect 1020 -20 1040 0
rect 1075 -20 1095 0
rect 1130 -20 1150 0
<< pdiffc >>
rect 635 185 655 205
rect 690 185 710 205
rect 745 185 765 205
rect 815 185 835 205
rect 870 185 890 205
rect 925 185 945 205
rect 1040 185 1060 205
rect 1095 185 1115 205
<< psubdiff >>
rect 1190 0 1230 15
rect 1190 -20 1200 0
rect 1220 -20 1230 0
rect 1190 -35 1230 -20
<< nsubdiff >>
rect 990 205 1030 220
rect 990 185 1000 205
rect 1020 185 1030 205
rect 990 170 1030 185
<< psubdiffcont >>
rect 1200 -20 1220 0
<< nsubdiffcont >>
rect 1000 185 1020 205
<< poly >>
rect 805 265 860 275
rect 805 245 815 265
rect 835 245 860 265
rect 665 230 735 245
rect 805 235 860 245
rect 665 220 680 230
rect 720 220 735 230
rect 845 220 860 235
rect 900 220 915 235
rect 1070 220 1085 235
rect 665 115 680 170
rect 720 155 735 170
rect 845 115 860 170
rect 900 155 915 170
rect 1070 155 1085 170
rect 885 145 925 155
rect 885 125 895 145
rect 915 125 925 145
rect 885 115 925 125
rect 1050 140 1085 155
rect 605 100 680 115
rect 665 15 680 100
rect 720 100 860 115
rect 720 15 735 100
rect 800 60 840 70
rect 800 40 810 60
rect 830 40 840 60
rect 1050 40 1065 140
rect 775 25 1065 40
rect 1090 60 1130 70
rect 1090 40 1100 60
rect 1120 40 1130 60
rect 1090 30 1130 40
rect 775 15 790 25
rect 940 15 955 25
rect 995 15 1010 25
rect 1050 15 1065 25
rect 1105 15 1120 30
rect 665 -50 680 -35
rect 720 -50 735 -35
rect 775 -50 790 -35
rect 940 -50 955 -35
rect 995 -50 1010 -35
rect 1050 -50 1065 -35
rect 1105 -50 1120 -35
<< polycont >>
rect 815 245 835 265
rect 895 125 915 145
rect 810 40 830 60
rect 1100 40 1120 60
<< locali >>
rect 605 300 635 320
rect 655 300 685 320
rect 705 300 735 320
rect 755 300 785 320
rect 805 300 835 320
rect 855 300 885 320
rect 905 300 935 320
rect 955 300 985 320
rect 1005 300 1035 320
rect 1055 300 1085 320
rect 1105 300 1135 320
rect 1155 300 1185 320
rect 1205 300 1235 320
rect 1255 300 1265 320
rect 690 215 710 300
rect 805 265 845 275
rect 805 245 815 265
rect 835 245 845 265
rect 805 235 845 245
rect 870 215 890 300
rect 1040 215 1060 300
rect 1095 265 1135 275
rect 1095 245 1105 265
rect 1125 245 1135 265
rect 1095 235 1135 245
rect 1095 215 1115 235
rect 630 205 660 215
rect 630 185 635 205
rect 655 185 660 205
rect 630 175 660 185
rect 685 205 715 215
rect 685 185 690 205
rect 710 185 715 205
rect 685 175 715 185
rect 740 205 770 215
rect 740 185 745 205
rect 765 185 770 205
rect 740 175 770 185
rect 810 205 840 215
rect 810 185 815 205
rect 835 185 840 205
rect 810 175 840 185
rect 865 205 895 215
rect 865 185 870 205
rect 890 185 895 205
rect 865 175 895 185
rect 920 205 965 215
rect 920 185 925 205
rect 945 185 965 205
rect 920 175 965 185
rect 995 205 1065 215
rect 995 185 1000 205
rect 1020 185 1040 205
rect 1060 185 1065 205
rect 995 175 1065 185
rect 1090 205 1120 215
rect 1090 185 1095 205
rect 1115 185 1175 205
rect 1090 175 1120 185
rect 635 50 655 175
rect 745 50 765 175
rect 815 155 835 175
rect 815 145 925 155
rect 815 135 895 145
rect 865 125 895 135
rect 915 125 925 145
rect 865 115 925 125
rect 800 60 840 70
rect 800 50 810 60
rect 635 40 810 50
rect 830 40 840 60
rect 635 30 840 40
rect 635 10 655 30
rect 865 10 885 115
rect 945 50 965 175
rect 1155 125 1175 185
rect 1155 105 1230 125
rect 1090 60 1130 70
rect 1090 50 1100 60
rect 910 40 1100 50
rect 1120 40 1130 60
rect 910 30 1130 40
rect 910 10 930 30
rect 1020 10 1040 30
rect 1155 10 1175 105
rect 630 0 660 10
rect 630 -20 635 0
rect 655 -20 660 0
rect 630 -30 660 -20
rect 685 0 715 10
rect 685 -20 690 0
rect 710 -20 715 0
rect 685 -30 715 -20
rect 740 0 770 10
rect 740 -20 745 0
rect 765 -20 770 0
rect 740 -30 770 -20
rect 795 0 885 10
rect 795 -20 800 0
rect 820 -10 885 0
rect 905 0 935 10
rect 820 -20 825 -10
rect 795 -30 825 -20
rect 905 -20 910 0
rect 930 -20 935 0
rect 905 -30 935 -20
rect 960 0 990 10
rect 960 -20 965 0
rect 985 -20 990 0
rect 960 -30 990 -20
rect 1015 0 1045 10
rect 1015 -20 1020 0
rect 1040 -20 1045 0
rect 1015 -30 1045 -20
rect 1070 0 1100 10
rect 1070 -20 1075 0
rect 1095 -20 1100 0
rect 1070 -30 1100 -20
rect 1125 0 1175 10
rect 1125 -20 1130 0
rect 1150 -20 1175 0
rect 1195 0 1225 10
rect 1195 -20 1200 0
rect 1220 -20 1225 0
rect 1125 -30 1155 -20
rect 1195 -30 1225 -20
rect 690 -70 710 -30
rect 965 -70 985 -30
rect 1075 -70 1095 -30
rect 1200 -70 1220 -30
rect 605 -90 635 -70
rect 655 -90 685 -70
rect 705 -90 735 -70
rect 755 -90 785 -70
rect 805 -90 835 -70
rect 855 -90 885 -70
rect 905 -90 935 -70
rect 955 -90 985 -70
rect 1005 -90 1035 -70
rect 1055 -90 1085 -70
rect 1105 -90 1135 -70
rect 1155 -90 1185 -70
rect 1205 -90 1235 -70
rect 1255 -90 1265 -70
<< viali >>
rect 635 300 655 320
rect 685 300 705 320
rect 735 300 755 320
rect 785 300 805 320
rect 835 300 855 320
rect 885 300 905 320
rect 935 300 955 320
rect 985 300 1005 320
rect 1035 300 1055 320
rect 1085 300 1105 320
rect 1135 300 1155 320
rect 1185 300 1205 320
rect 1235 300 1255 320
rect 815 245 835 265
rect 1105 245 1125 265
rect 635 -90 655 -70
rect 685 -90 705 -70
rect 735 -90 755 -70
rect 785 -90 805 -70
rect 835 -90 855 -70
rect 885 -90 905 -70
rect 935 -90 955 -70
rect 985 -90 1005 -70
rect 1035 -90 1055 -70
rect 1085 -90 1105 -70
rect 1135 -90 1155 -70
rect 1185 -90 1205 -70
rect 1235 -90 1255 -70
<< metal1 >>
rect 605 320 1265 330
rect 605 300 635 320
rect 655 300 685 320
rect 705 300 735 320
rect 755 300 785 320
rect 805 300 835 320
rect 855 300 885 320
rect 905 300 935 320
rect 955 300 985 320
rect 1005 300 1035 320
rect 1055 300 1085 320
rect 1105 300 1135 320
rect 1155 300 1185 320
rect 1205 300 1235 320
rect 1255 300 1265 320
rect 605 290 1265 300
rect 805 265 845 275
rect 805 245 815 265
rect 835 255 845 265
rect 1095 265 1135 275
rect 1095 255 1105 265
rect 835 245 1105 255
rect 1125 245 1135 265
rect 805 235 1135 245
rect 1095 215 1115 235
rect 605 -70 1265 -60
rect 605 -90 635 -70
rect 655 -90 685 -70
rect 705 -90 735 -70
rect 755 -90 785 -70
rect 805 -90 835 -70
rect 855 -90 885 -70
rect 905 -90 935 -70
rect 955 -90 985 -70
rect 1005 -90 1035 -70
rect 1055 -90 1085 -70
rect 1105 -90 1135 -70
rect 1155 -90 1185 -70
rect 1205 -90 1235 -70
rect 1255 -90 1265 -70
rect 605 -100 1265 -90
<< labels >>
flabel locali 755 -30 755 -30 5 FreeSans 160 0 0 -80 B
flabel metal1 605 -80 605 -80 7 FreeSans 160 0 -80 0 GNDA
port 4 w
flabel metal1 605 310 605 310 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel poly 605 105 605 105 7 FreeSans 160 0 -80 0 VIN
port 2 w
flabel locali 965 125 965 125 3 FreeSans 160 0 80 0 C
flabel locali 1230 115 1230 115 3 FreeSans 160 0 80 0 VOUT
port 1 e
flabel space 700 95 700 95 1 FreeSans 160 0 0 80 CLK
flabel locali 885 100 885 100 3 FreeSans 160 0 80 0 A
<< end >>
