* PEX produced on Mon Feb  3 12:34:26 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from phase_frequency_detector_magic.ext - technology: sky130A

.subckt phase_frequency_detector_magic F_REF F_VCO VDDA QA QB GNDA
X0 GNDA.t32 Reset.t2 F_b.t0 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1 a_1430_320.t1 E.t3 E_b.t1 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X2 QB_b.t2 QB.t3 a_1790_320.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X3 a_3930_0.t1 before_Reset.t3 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X4 F.t2 QB_b.t3 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X5 F.t0 F_b.t3 a_2690_320.t0 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 a_550_320.t1 QA_b.t3 QA.t1 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X7 E.t0 E_b.t3 a_910_320.t0 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X8 QA_b.t0 F_REF.t0 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X9 GNDA.t21 QA.t3 QA_b.t1 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X10 E.t2 QA_b.t4 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X11 E_b.t2 E.t4 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X12 GNDA.t34 F_b.t4 F.t1 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 VDDA.t16 QA.t4 before_Reset.t0 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X14 GNDA.t26 E_b.t4 E.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X15 QB.t0 QB_b.t4 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 a_4430_0.t1 a_4180_0.t2 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X17 GNDA.t30 Reset.t3 E_b.t0 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X18 Reset.t0 a_4680_0.t2 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X19 a_2310_320.t1 QB_b.t5 QB.t1 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X20 a_3210_320.t1 F.t3 F_b.t2 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X21 a_4430_0.t0 a_4180_0.t3 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X22 a_4680_0.t1 a_4430_0.t2 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X23 GNDA.t40 F.t4 QB.t2 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X24 VDDA.t24 Reset.t4 a_1430_320.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X25 QB_b.t0 F_VCO.t0 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X26 a_3930_0.t0 before_Reset.t4 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X27 QA_b.t2 QA.t5 a_30_320.t0 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 VDDA.t27 E.t5 a_550_320.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X29 a_4680_0.t0 a_4430_0.t3 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X30 a_1790_320.t0 F_VCO.t1 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X31 GNDA.t24 QB.t4 QB_b.t1 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X32 a_2690_320.t1 QB_b.t6 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X33 before_Reset.t1 QB.t5 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X34 a_4180_0.t0 a_3930_0.t2 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X35 a_910_320.t1 QA_b.t5 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X36 a_3570_0.t0 QA.t6 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X37 a_30_320.t1 F_REF.t1 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X38 VDDA.t33 F.t5 a_2310_320.t0 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X39 QA.t2 QA_b.t6 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X40 Reset.t1 a_4680_0.t3 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X41 F_b.t1 F.t6 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X42 before_Reset.t2 QB.t6 a_3570_0.t1 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X43 VDDA.t22 Reset.t5 a_3210_320.t0 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X44 a_4180_0.t1 a_3930_0.t3 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X45 GNDA.t17 E.t6 QA.t0 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
R0 Reset.n1 Reset.n0 3646.5
R1 Reset.n0 Reset.t4 3277.6
R2 Reset.t4 Reset.t3 594.467
R3 Reset.t5 Reset.t2 594.467
R4 Reset.n0 Reset.t5 417.733
R5 Reset.t1 Reset.n1 378.62
R6 Reset.n1 Reset.t0 275.454
R7 F_b.n0 F_b.t3 356.68
R8 F_b.n2 F_b.n0 333.334
R9 F_b.t2 F_b.n2 331.901
R10 F_b.n2 F_b.n1 311.933
R11 F_b.n0 F_b.t4 147.814
R12 F_b.n1 F_b.t0 48.0005
R13 F_b.n1 F_b.t1 48.0005
R14 GNDA.t33 GNDA.t37 3838.3
R15 GNDA.t6 GNDA.t23 3838.3
R16 GNDA.t0 GNDA.t25 3838.3
R17 GNDA.t43 GNDA.t20 3838.3
R18 GNDA.t12 GNDA.t14 2340.43
R19 GNDA.t8 GNDA.t12 2340.43
R20 GNDA.t27 GNDA.t8 2340.43
R21 GNDA.t35 GNDA.t27 2340.43
R22 GNDA.t22 GNDA.t35 2340.43
R23 GNDA.t31 GNDA.t18 2340.43
R24 GNDA.t4 GNDA.t29 2340.43
R25 GNDA.t41 GNDA.t16 2340.43
R26 GNDA.n11 GNDA.t2 1263.83
R27 GNDA.n11 GNDA.t39 1263.83
R28 GNDA.n12 GNDA.n11 1170
R29 GNDA.t18 GNDA.t22 1029.79
R30 GNDA.t37 GNDA.t31 1029.79
R31 GNDA.t2 GNDA.t33 1029.79
R32 GNDA.t39 GNDA.t6 1029.79
R33 GNDA.t23 GNDA.t4 1029.79
R34 GNDA.t29 GNDA.t0 1029.79
R35 GNDA.t25 GNDA.t41 1029.79
R36 GNDA.t16 GNDA.t43 1029.79
R37 GNDA.t20 GNDA.t10 1029.79
R38 GNDA.n1 GNDA.t15 242.613
R39 GNDA.n25 GNDA.t11 242.3
R40 GNDA.n24 GNDA.t21 242.3
R41 GNDA.n23 GNDA.t44 242.3
R42 GNDA.n22 GNDA.t17 242.3
R43 GNDA.n21 GNDA.t42 242.3
R44 GNDA.n20 GNDA.t26 242.3
R45 GNDA.n19 GNDA.t1 242.3
R46 GNDA.n18 GNDA.t30 242.3
R47 GNDA.n17 GNDA.t5 242.3
R48 GNDA.n16 GNDA.t24 242.3
R49 GNDA.n15 GNDA.t7 242.3
R50 GNDA.n8 GNDA.t34 242.3
R51 GNDA.n7 GNDA.t38 242.3
R52 GNDA.n6 GNDA.t32 242.3
R53 GNDA.n5 GNDA.t19 242.3
R54 GNDA.n4 GNDA.t36 242.3
R55 GNDA.n3 GNDA.t28 242.3
R56 GNDA.n2 GNDA.t9 242.3
R57 GNDA.n1 GNDA.t13 242.3
R58 GNDA.n13 GNDA.t40 233
R59 GNDA.n10 GNDA.t3 233
R60 GNDA.n12 GNDA.n10 12.8005
R61 GNDA.n13 GNDA.n12 12.8005
R62 GNDA.n10 GNDA.n9 9.3005
R63 GNDA.n12 GNDA.n0 9.3005
R64 GNDA.n14 GNDA.n13 9.3005
R65 GNDA.n5 GNDA.n4 0.4505
R66 GNDA.n8 GNDA.n7 0.3755
R67 GNDA.n16 GNDA.n15 0.3755
R68 GNDA.n20 GNDA.n19 0.3755
R69 GNDA.n24 GNDA.n23 0.3755
R70 GNDA.n2 GNDA.n1 0.313
R71 GNDA.n3 GNDA.n2 0.313
R72 GNDA.n4 GNDA.n3 0.313
R73 GNDA.n7 GNDA.n6 0.2755
R74 GNDA.n9 GNDA.n8 0.2755
R75 GNDA.n15 GNDA.n14 0.2755
R76 GNDA.n17 GNDA.n16 0.2755
R77 GNDA.n19 GNDA.n18 0.2755
R78 GNDA.n21 GNDA.n20 0.2755
R79 GNDA.n23 GNDA.n22 0.2755
R80 GNDA.n25 GNDA.n24 0.2755
R81 GNDA.n6 GNDA.n5 0.1755
R82 GNDA.n18 GNDA.n17 0.1755
R83 GNDA.n22 GNDA.n21 0.1755
R84 GNDA.n9 GNDA.n0 0.1005
R85 GNDA.n14 GNDA.n0 0.1005
R86 GNDA GNDA.n25 0.0505
R87 E.n4 E.n0 977.808
R88 E.n0 E.t3 401.668
R89 E.t0 E.n4 331.901
R90 E.n2 E.t6 276.348
R91 E.n3 E.n1 244.733
R92 E.n2 E.t5 228.148
R93 E.n3 E.n2 225.601
R94 E.n0 E.t4 144.601
R95 E.n4 E.n3 70.4005
R96 E.n1 E.t1 48.0005
R97 E.n1 E.t2 48.0005
R98 E_b.n0 E_b.t3 356.68
R99 E_b.n2 E_b.n0 333.334
R100 E_b.t1 E_b.n2 331.901
R101 E_b.n2 E_b.n1 311.933
R102 E_b.n0 E_b.t4 147.814
R103 E_b.n1 E_b.t0 48.0005
R104 E_b.n1 E_b.t2 48.0005
R105 a_1430_320.t0 a_1430_320.t1 78.8005
R106 VDDA.t25 VDDA.t35 1391.07
R107 VDDA.t8 VDDA.t13 1391.07
R108 VDDA.t28 VDDA.t34 1391.07
R109 VDDA.t14 VDDA.t31 1391.07
R110 VDDA.t9 VDDA.t17 848.215
R111 VDDA.t6 VDDA.t9 848.215
R112 VDDA.t29 VDDA.t6 848.215
R113 VDDA.t19 VDDA.t29 848.215
R114 VDDA.t4 VDDA.t19 848.215
R115 VDDA.t21 VDDA.t15 848.215
R116 VDDA.t2 VDDA.t23 848.215
R117 VDDA.t36 VDDA.t26 848.215
R118 VDDA.n10 VDDA.t11 458.036
R119 VDDA.n10 VDDA.t32 458.036
R120 VDDA.t15 VDDA.t4 373.214
R121 VDDA.t35 VDDA.t21 373.214
R122 VDDA.t11 VDDA.t25 373.214
R123 VDDA.t32 VDDA.t8 373.214
R124 VDDA.t13 VDDA.t2 373.214
R125 VDDA.t23 VDDA.t28 373.214
R126 VDDA.t34 VDDA.t36 373.214
R127 VDDA.t26 VDDA.t14 373.214
R128 VDDA.t31 VDDA.t0 373.214
R129 VDDA.n1 VDDA.t18 336.707
R130 VDDA.n18 VDDA.t1 336.55
R131 VDDA.n17 VDDA.t27 336.55
R132 VDDA.n16 VDDA.t37 336.55
R133 VDDA.n15 VDDA.t24 336.55
R134 VDDA.n14 VDDA.t3 336.55
R135 VDDA.n7 VDDA.t22 336.55
R136 VDDA.n4 VDDA.t20 336.55
R137 VDDA.n3 VDDA.t30 336.55
R138 VDDA.n2 VDDA.t7 336.55
R139 VDDA.n1 VDDA.t10 336.55
R140 VDDA.n12 VDDA.t33 331.901
R141 VDDA.n9 VDDA.t12 331.901
R142 VDDA.n6 VDDA.n5 297.151
R143 VDDA.n11 VDDA.n10 185
R144 VDDA.n5 VDDA.t5 39.4005
R145 VDDA.n5 VDDA.t16 39.4005
R146 VDDA.n11 VDDA.n9 5.68939
R147 VDDA.n12 VDDA.n11 5.68939
R148 VDDA.n9 VDDA.n8 4.6505
R149 VDDA.n11 VDDA.n0 4.6505
R150 VDDA.n13 VDDA.n12 4.6505
R151 VDDA.n8 VDDA.n7 0.463
R152 VDDA.n14 VDDA.n13 0.463
R153 VDDA.n16 VDDA.n15 0.463
R154 VDDA.n18 VDDA.n17 0.463
R155 VDDA.n2 VDDA.n1 0.15675
R156 VDDA.n3 VDDA.n2 0.15675
R157 VDDA.n4 VDDA.n3 0.15675
R158 VDDA.n6 VDDA.n4 0.15675
R159 VDDA.n7 VDDA.n6 0.15675
R160 VDDA.n15 VDDA.n14 0.088
R161 VDDA.n17 VDDA.n16 0.088
R162 VDDA.n8 VDDA.n0 0.0505
R163 VDDA.n13 VDDA.n0 0.0505
R164 VDDA VDDA.n18 0.0255
R165 QB.t6 QB.t5 594.467
R166 QB.n4 QB.n3 443.733
R167 QB QB.n4 432
R168 QB.n0 QB.t3 356.68
R169 QB.n1 QB.n0 333.334
R170 QB.n1 QB.t1 331.901
R171 QB.n4 QB.t6 304.634
R172 QB.n3 QB.n2 185
R173 QB.n0 QB.t4 147.814
R174 QB.n3 QB.n1 126.933
R175 QB.n2 QB.t2 48.0005
R176 QB.n2 QB.t0 48.0005
R177 a_1790_320.t0 a_1790_320.t1 78.8005
R178 QB_b.t4 QB_b.t3 1028.27
R179 QB_b.t3 QB_b.t6 594.467
R180 QB_b QB_b.n2 514.134
R181 QB_b QB_b.n1 463.673
R182 QB_b.n2 QB_b.t5 401.668
R183 QB_b.n1 QB_b.t2 331.901
R184 QB_b.n1 QB_b.n0 315.134
R185 QB_b.n2 QB_b.t4 144.601
R186 QB_b.n0 QB_b.t1 48.0005
R187 QB_b.n0 QB_b.t0 48.0005
R188 before_Reset.t0 before_Reset.n2 427.901
R189 before_Reset.n2 before_Reset.t1 370.3
R190 before_Reset.n1 before_Reset.n0 349.601
R191 before_Reset.n0 before_Reset.t3 305.267
R192 before_Reset.n1 before_Reset.t2 284.841
R193 before_Reset.n0 before_Reset.t4 241
R194 before_Reset.n2 before_Reset.n1 16.0005
R195 a_3930_0.t1 a_3930_0.n1 378.62
R196 a_3930_0.n1 a_3930_0.n0 344.8
R197 a_3930_0.n0 a_3930_0.t3 305.267
R198 a_3930_0.n1 a_3930_0.t0 275.454
R199 a_3930_0.n0 a_3930_0.t2 241
R200 F.n4 F.n0 977.808
R201 F.n0 F.t3 401.668
R202 F.t0 F.n4 331.901
R203 F.n2 F.t4 276.348
R204 F.n3 F.n1 244.733
R205 F.n3 F.n2 232
R206 F.n2 F.t5 228.148
R207 F.n0 F.t6 144.601
R208 F.n4 F.n3 70.4005
R209 F.n1 F.t1 48.0005
R210 F.n1 F.t2 48.0005
R211 a_2690_320.t0 a_2690_320.t1 78.8005
R212 QA_b.t6 QA_b.t4 996.134
R213 QA_b.t4 QA_b.t5 594.467
R214 QA_b QA_b.n1 495.808
R215 QA_b QA_b.n2 482
R216 QA_b.n2 QA_b.t3 401.668
R217 QA_b.n1 QA_b.t2 331.901
R218 QA_b.n1 QA_b.n0 315.134
R219 QA_b.n2 QA_b.t6 144.601
R220 QA_b.n0 QA_b.t1 48.0005
R221 QA_b.n0 QA_b.t0 48.0005
R222 QA.n4 QA.n3 1001.6
R223 QA.t4 QA.t6 594.467
R224 QA QA.n4 483.2
R225 QA.n4 QA.t4 384.967
R226 QA.n0 QA.t5 356.68
R227 QA.n2 QA.t1 331.901
R228 QA.n2 QA.n1 311.933
R229 QA.n3 QA.n0 299.2
R230 QA.n0 QA.t3 147.814
R231 QA.n1 QA.t0 48.0005
R232 QA.n1 QA.t2 48.0005
R233 QA.n3 QA.n2 34.1338
R234 a_550_320.t0 a_550_320.t1 78.8005
R235 a_910_320.t0 a_910_320.t1 78.8005
R236 F_REF.n0 F_REF.t1 353.467
R237 F_REF F_REF.n0 216.9
R238 F_REF.n0 F_REF.t0 192.8
R239 a_4180_0.t1 a_4180_0.n1 378.62
R240 a_4180_0.n1 a_4180_0.n0 344.8
R241 a_4180_0.n0 a_4180_0.t2 305.267
R242 a_4180_0.n1 a_4180_0.t0 275.454
R243 a_4180_0.n0 a_4180_0.t3 241
R244 a_4430_0.t1 a_4430_0.n1 378.62
R245 a_4430_0.n1 a_4430_0.n0 344.8
R246 a_4430_0.n0 a_4430_0.t2 305.267
R247 a_4430_0.n1 a_4430_0.t0 275.454
R248 a_4430_0.n0 a_4430_0.t3 241
R249 a_4680_0.t1 a_4680_0.n1 378.62
R250 a_4680_0.n1 a_4680_0.n0 344.8
R251 a_4680_0.n0 a_4680_0.t3 305.267
R252 a_4680_0.n1 a_4680_0.t0 275.454
R253 a_4680_0.n0 a_4680_0.t2 241
R254 a_2310_320.t0 a_2310_320.t1 78.8005
R255 a_3210_320.t0 a_3210_320.t1 78.8005
R256 F_VCO F_VCO.t0 3382.03
R257 F_VCO.t0 F_VCO.t1 594.467
R258 a_30_320.t0 a_30_320.t1 78.8005
R259 a_3570_0.t0 a_3570_0.t1 96.0005
C0 F_VCO QA_b 0.141561f
C1 VDDA QB 0.312516f
C2 QA QA_b 0.321451f
C3 VDDA F_VCO 0.058995f
C4 VDDA QA 1.39534f
C5 VDDA QB_b 0.451913f
C6 F_VCO QB 0.056132f
C7 QA QB 0.159324f
C8 QA F_VCO 0.017952f
C9 QB_b QB 0.354572f
C10 F_REF QA_b 0.021974f
C11 F_VCO QB_b 0.021493f
C12 QA QB_b 0.08944f
C13 VDDA F_REF 0.062052f
C14 VDDA QA_b 0.44408f
C15 QA F_REF 0.056153f
C16 QB GNDA 2.0664f
C17 F_VCO GNDA 1.33173f
C18 F_REF GNDA 0.228052f
C19 QA GNDA 1.85881f
C20 VDDA GNDA 6.31463f
C21 QB_b GNDA 0.914709f
C22 QA_b GNDA 0.906621f
.ends

