magic
tech sky130A
timestamp 1751481783
<< metal1 >>
rect 6370 5475 6410 5480
rect 6370 5445 6375 5475
rect 6405 5445 6410 5475
rect 6370 5440 6410 5445
rect 9975 5475 10015 5480
rect 9975 5445 9980 5475
rect 10010 5445 10015 5475
rect 9975 5440 10015 5445
rect 6270 5430 6310 5435
rect 6270 5400 6275 5430
rect 6305 5400 6310 5430
rect 6270 5395 6310 5400
rect 6280 5290 6300 5395
rect 6270 5285 6310 5290
rect 6270 5255 6275 5285
rect 6305 5255 6310 5285
rect 6270 5250 6310 5255
rect 6380 5140 6400 5440
rect 6370 5135 6410 5140
rect 6370 5105 6375 5135
rect 6405 5105 6410 5135
rect 6370 5100 6410 5105
rect 2935 5090 2975 5095
rect 2935 5060 2940 5090
rect 2970 5060 2975 5090
rect 2935 5055 2975 5060
rect 9875 5065 9915 5070
rect 2365 3215 2405 3220
rect 2365 3185 2370 3215
rect 2400 3185 2405 3215
rect 2365 3180 2405 3185
rect 2375 940 2395 3180
rect 2945 3045 2965 5055
rect 9875 5035 9880 5065
rect 9910 5035 9915 5065
rect 9875 5030 9915 5035
rect 9885 5010 9905 5030
rect 7120 4760 7160 4765
rect 7120 4730 7125 4760
rect 7155 4730 7160 4760
rect 7120 4725 7160 4730
rect 5025 4715 5065 4720
rect 5025 4685 5030 4715
rect 5060 4685 5065 4715
rect 5025 4680 5065 4685
rect 5035 4410 5055 4680
rect 6295 4465 6335 4470
rect 6295 4435 6300 4465
rect 6330 4435 6335 4465
rect 6295 4430 6335 4435
rect 6305 4410 6325 4430
rect 5025 4405 5065 4410
rect 5025 4375 5030 4405
rect 5060 4375 5065 4405
rect 5025 4370 5065 4375
rect 6295 4405 6335 4410
rect 6295 4375 6300 4405
rect 6330 4375 6335 4405
rect 6295 4370 6335 4375
rect 2980 3215 3020 3220
rect 2980 3185 2985 3215
rect 3015 3185 3020 3215
rect 2980 3180 3020 3185
rect 7075 3215 7115 3220
rect 7075 3185 7080 3215
rect 7110 3185 7115 3215
rect 7075 3180 7115 3185
rect 2990 2850 3010 3180
rect 7085 2855 7105 3180
rect 7130 3045 7150 4725
rect 9855 4515 9895 4520
rect 9855 4485 9860 4515
rect 9890 4485 9895 4515
rect 9855 4480 9895 4485
rect 9620 4415 9660 4420
rect 9620 4385 9625 4415
rect 9655 4385 9660 4415
rect 9620 4380 9660 4385
rect 7790 4370 7830 4375
rect 7790 4340 7795 4370
rect 7825 4340 7830 4370
rect 7790 4335 7830 4340
rect 7685 3215 7725 3220
rect 7685 3185 7690 3215
rect 7720 3185 7725 3215
rect 7685 3180 7725 3185
rect 5960 2405 6000 2410
rect 5960 2375 5965 2405
rect 5995 2375 6000 2405
rect 5960 2370 6000 2375
rect 2365 935 2405 940
rect 2365 905 2370 935
rect 2400 905 2405 935
rect 2365 900 2405 905
rect 3985 895 4005 1260
rect 5970 1155 5990 2370
rect 7695 1960 7715 3180
rect 7685 1955 7725 1960
rect 7685 1925 7690 1955
rect 7720 1925 7725 1955
rect 7685 1920 7725 1925
rect 7800 1155 7820 4335
rect 9630 3450 9650 4380
rect 9865 4375 9885 4480
rect 9855 4370 9895 4375
rect 9855 4340 9860 4370
rect 9890 4340 9895 4370
rect 9855 4335 9895 4340
rect 9855 4195 9895 4200
rect 9855 4165 9860 4195
rect 9890 4165 9895 4195
rect 9855 4160 9895 4165
rect 9620 3445 9660 3450
rect 9620 3415 9625 3445
rect 9655 3415 9660 3445
rect 9620 3410 9660 3415
rect 5960 1150 6000 1155
rect 5960 1120 5965 1150
rect 5995 1120 6000 1150
rect 5960 1115 6000 1120
rect 7790 1150 7830 1155
rect 7790 1120 7795 1150
rect 7825 1120 7830 1150
rect 7790 1115 7830 1120
rect 9865 895 9885 4160
rect 9985 1915 10005 5440
rect 10030 5430 10070 5435
rect 10030 5400 10035 5430
rect 10065 5400 10070 5430
rect 10030 5395 10070 5400
rect 9975 1910 10015 1915
rect 9975 1880 9980 1910
rect 10010 1880 10015 1910
rect 9975 1875 10015 1880
rect 10045 1870 10065 5395
rect 10090 4715 10130 4720
rect 10090 4685 10095 4715
rect 10125 4685 10130 4715
rect 10090 4680 10130 4685
rect 10035 1865 10075 1870
rect 10035 1835 10040 1865
rect 10070 1835 10075 1865
rect 10035 1830 10075 1835
rect 10100 1825 10120 4680
rect 11160 1955 11200 1960
rect 11160 1925 11165 1955
rect 11195 1925 11200 1955
rect 11160 1920 11200 1925
rect 11785 1870 11805 1950
rect 11895 1915 11915 1950
rect 11885 1910 11925 1915
rect 11885 1880 11890 1910
rect 11920 1880 11925 1910
rect 11885 1875 11925 1880
rect 11775 1865 11815 1870
rect 11775 1835 11780 1865
rect 11810 1835 11815 1865
rect 11775 1830 11815 1835
rect 12005 1825 12025 1950
rect 10090 1820 10130 1825
rect 10090 1790 10095 1820
rect 10125 1790 10130 1820
rect 10090 1785 10130 1790
rect 11995 1820 12035 1825
rect 11995 1790 12000 1820
rect 12030 1790 12035 1820
rect 11995 1785 12035 1790
rect 12620 940 12640 1950
rect 12610 935 12650 940
rect 12610 905 12615 935
rect 12645 905 12650 935
rect 12610 900 12650 905
rect 3975 890 4015 895
rect 3975 860 3980 890
rect 4010 860 4015 890
rect 3975 855 4015 860
rect 9855 890 9895 895
rect 9855 860 9860 890
rect 9890 860 9895 890
rect 9855 855 9895 860
<< via1 >>
rect 6375 5445 6405 5475
rect 9980 5445 10010 5475
rect 6275 5400 6305 5430
rect 6275 5255 6305 5285
rect 6375 5105 6405 5135
rect 2940 5060 2970 5090
rect 2370 3185 2400 3215
rect 9880 5035 9910 5065
rect 7125 4730 7155 4760
rect 5030 4685 5060 4715
rect 6300 4435 6330 4465
rect 5030 4375 5060 4405
rect 6300 4375 6330 4405
rect 2985 3185 3015 3215
rect 7080 3185 7110 3215
rect 9860 4485 9890 4515
rect 9625 4385 9655 4415
rect 7795 4340 7825 4370
rect 7690 3185 7720 3215
rect 5965 2375 5995 2405
rect 2370 905 2400 935
rect 7690 1925 7720 1955
rect 9860 4340 9890 4370
rect 9860 4165 9890 4195
rect 9625 3415 9655 3445
rect 5965 1120 5995 1150
rect 7795 1120 7825 1150
rect 10035 5400 10065 5430
rect 9980 1880 10010 1910
rect 10095 4685 10125 4715
rect 10040 1835 10070 1865
rect 11165 1925 11195 1955
rect 11890 1880 11920 1910
rect 11780 1835 11810 1865
rect 10095 1790 10125 1820
rect 12000 1790 12030 1820
rect 12615 905 12645 935
rect 3980 860 4010 890
rect 9860 860 9890 890
<< metal2 >>
rect 6370 5475 6410 5480
rect 6370 5445 6375 5475
rect 6405 5470 6410 5475
rect 9975 5475 10015 5480
rect 9975 5470 9980 5475
rect 6405 5450 9980 5470
rect 6405 5445 6410 5450
rect 6370 5440 6410 5445
rect 9975 5445 9980 5450
rect 10010 5445 10015 5475
rect 9975 5440 10015 5445
rect 6270 5430 6310 5435
rect 6270 5400 6275 5430
rect 6305 5425 6310 5430
rect 10030 5430 10070 5435
rect 10030 5425 10035 5430
rect 6305 5405 10035 5425
rect 6305 5400 6310 5405
rect 6270 5395 6310 5400
rect 10030 5400 10035 5405
rect 10065 5400 10070 5430
rect 10030 5395 10070 5400
rect 6270 5285 6310 5290
rect 6270 5280 6275 5285
rect 5630 5260 6275 5280
rect 6270 5255 6275 5260
rect 6305 5255 6310 5285
rect 6270 5250 6310 5255
rect 6370 5135 6410 5140
rect 6370 5130 6375 5135
rect 5580 5110 6375 5130
rect 6370 5105 6375 5110
rect 6405 5105 6410 5135
rect 6370 5100 6410 5105
rect 2935 5090 2975 5095
rect 2935 5060 2940 5090
rect 2970 5085 2975 5090
rect 2970 5065 9915 5085
rect 2970 5060 2975 5065
rect 2935 5055 2975 5060
rect 9875 5035 9880 5065
rect 9910 5035 9915 5065
rect 9875 5030 9915 5035
rect 7120 4760 7160 4765
rect 7120 4730 7125 4760
rect 7155 4755 7160 4760
rect 7155 4735 9885 4755
rect 7155 4730 7160 4735
rect 7120 4725 7160 4730
rect 5025 4715 5065 4720
rect 5025 4685 5030 4715
rect 5060 4710 5065 4715
rect 10090 4715 10130 4720
rect 10090 4710 10095 4715
rect 5060 4690 10095 4710
rect 5060 4685 5065 4690
rect 5025 4680 5065 4685
rect 10090 4685 10095 4690
rect 10125 4685 10130 4715
rect 10090 4680 10130 4685
rect 9855 4515 9895 4520
rect 9855 4485 9860 4515
rect 9890 4485 9895 4515
rect 9855 4480 9895 4485
rect 6295 4465 6335 4470
rect 6295 4460 6300 4465
rect 5785 4440 6300 4460
rect 6295 4435 6300 4440
rect 6330 4435 6335 4465
rect 6295 4430 6335 4435
rect 9620 4415 9660 4420
rect 9620 4410 9625 4415
rect 5025 4405 5065 4410
rect 5025 4400 5030 4405
rect 4860 4380 5030 4400
rect 5025 4375 5030 4380
rect 5060 4375 5065 4405
rect 5025 4370 5065 4375
rect 6295 4405 9625 4410
rect 6295 4375 6300 4405
rect 6330 4390 9625 4405
rect 6330 4375 6335 4390
rect 9620 4385 9625 4390
rect 9655 4385 9660 4415
rect 9620 4380 9660 4385
rect 6295 4370 6335 4375
rect 7790 4370 7830 4375
rect 7790 4340 7795 4370
rect 7825 4365 7830 4370
rect 9855 4370 9895 4375
rect 9855 4365 9860 4370
rect 7825 4345 9860 4365
rect 7825 4340 7830 4345
rect 7790 4335 7830 4340
rect 9855 4340 9860 4345
rect 9890 4340 9895 4370
rect 9855 4335 9895 4340
rect 9855 4195 9895 4200
rect 9855 4165 9860 4195
rect 9890 4165 9895 4195
rect 9855 4160 9895 4165
rect 9620 3445 9660 3450
rect 9620 3415 9625 3445
rect 9655 3440 9660 3445
rect 9655 3420 9885 3440
rect 9655 3415 9660 3420
rect 9620 3410 9660 3415
rect 2365 3215 2405 3220
rect 2365 3185 2370 3215
rect 2400 3210 2405 3215
rect 2980 3215 3020 3220
rect 2980 3210 2985 3215
rect 2400 3190 2985 3210
rect 2400 3185 2405 3190
rect 2365 3180 2405 3185
rect 2980 3185 2985 3190
rect 3015 3185 3020 3215
rect 2980 3180 3020 3185
rect 7075 3215 7115 3220
rect 7075 3185 7080 3215
rect 7110 3210 7115 3215
rect 7685 3215 7725 3220
rect 7685 3210 7690 3215
rect 7110 3190 7690 3210
rect 7110 3185 7115 3190
rect 7075 3180 7115 3185
rect 7685 3185 7690 3190
rect 7720 3185 7725 3215
rect 7685 3180 7725 3185
rect 5960 2405 6000 2410
rect 5960 2400 5965 2405
rect 5125 2380 5965 2400
rect 5960 2375 5965 2380
rect 5995 2375 6000 2405
rect 5960 2370 6000 2375
rect 7685 1955 7725 1960
rect 7685 1925 7690 1955
rect 7720 1950 7725 1955
rect 11160 1955 11200 1960
rect 11160 1950 11165 1955
rect 7720 1930 11165 1950
rect 7720 1925 7725 1930
rect 7685 1920 7725 1925
rect 11160 1925 11165 1930
rect 11195 1925 11200 1955
rect 11160 1920 11200 1925
rect 9975 1910 10015 1915
rect 9975 1880 9980 1910
rect 10010 1905 10015 1910
rect 11885 1910 11925 1915
rect 11885 1905 11890 1910
rect 10010 1885 11890 1905
rect 10010 1880 10015 1885
rect 9975 1875 10015 1880
rect 11885 1880 11890 1885
rect 11920 1880 11925 1910
rect 11885 1875 11925 1880
rect 10035 1865 10075 1870
rect 10035 1835 10040 1865
rect 10070 1860 10075 1865
rect 11775 1865 11815 1870
rect 11775 1860 11780 1865
rect 10070 1840 11780 1860
rect 10070 1835 10075 1840
rect 10035 1830 10075 1835
rect 11775 1835 11780 1840
rect 11810 1835 11815 1865
rect 11775 1830 11815 1835
rect 10090 1820 10130 1825
rect 10090 1790 10095 1820
rect 10125 1815 10130 1820
rect 11995 1820 12035 1825
rect 11995 1815 12000 1820
rect 10125 1795 12000 1815
rect 10125 1790 10130 1795
rect 10090 1785 10130 1790
rect 11995 1790 12000 1795
rect 12030 1790 12035 1820
rect 11995 1785 12035 1790
rect 5960 1150 6000 1155
rect 5960 1120 5965 1150
rect 5995 1145 6000 1150
rect 7790 1150 7830 1155
rect 7790 1145 7795 1150
rect 5995 1125 7795 1145
rect 5995 1120 6000 1125
rect 5960 1115 6000 1120
rect 7790 1120 7795 1125
rect 7825 1120 7830 1150
rect 7790 1115 7830 1120
rect 2365 935 2405 940
rect 2365 905 2370 935
rect 2400 930 2405 935
rect 12610 935 12650 940
rect 12610 930 12615 935
rect 2400 910 12615 930
rect 2400 905 2405 910
rect 2365 900 2405 905
rect 12610 905 12615 910
rect 12645 905 12650 935
rect 12610 900 12650 905
rect 3975 890 4015 895
rect 3975 860 3980 890
rect 4010 885 4015 890
rect 9855 890 9895 895
rect 9855 885 9860 890
rect 4010 865 9860 885
rect 4010 860 4015 865
rect 3975 855 4015 860
rect 9855 860 9860 865
rect 9890 860 9895 890
rect 9855 855 9895 860
<< metal3 >>
rect 10280 50 10320 2015
rect 10275 45 10325 50
rect 10275 5 10280 45
rect 10320 5 10325 45
rect 10275 0 10325 5
<< via3 >>
rect 10280 5 10320 45
<< metal4 >>
rect 9690 6700 10190 6750
rect 9690 45 10325 50
rect 9690 5 10280 45
rect 10320 5 10325 45
rect 9690 0 10325 5
use bgr  bgr_0
timestamp 1751468312
transform -1 0 15985 0 1 1400
box -200 535 6100 5350
use two_stage_opamp_dummy_magic  two_stage_opamp_dummy_magic_0
timestamp 1751466479
transform 1 0 -26855 0 1 555
box 26855 -555 36545 6195
<< labels >>
flabel metal4 10000 0 10000 0 5 FreeSans 800 0 0 -400 GNDA
port 2 s
flabel metal4 9965 6750 9965 6750 1 FreeSans 800 0 0 400 VDDA
port 1 n
<< end >>
