** sch_path: /foss/designs/my_design/projects/montecarlo/xschem_ngspice/inverter/common_source_mc.sch
**.subckt common_source_mc
XM1 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdd VDD GND 1.8
Vin Vin GND sin(1.2 0.01 1k)
XR1 VDD Vout GND sky130_fd_pr__res_xhigh_po_0p35 L=0.70 mult=1 m=1
**** begin user architecture code



.option wnflag=1
.option savecurrents
.save
+@m.xm1.msky130_fd_pr__nfet_01v8[gm]
+@m.xm1.msky130_fd_pr__nfet_01v8[vth]
+@m.xm2.msky130_fd_pr__pfet_01v8[gm]
+@m.xm2.msky130_fd_pr__pfet_01v8[vth]

.control

  let runs=100
  let run=1

  dowhile run <= runs
    save all
    * dc vin 0 1.8 0.01
    tran 1u 3m
    write common_source_mc.raw
    set appendwrite
    reset
    let run = run + 1
  end

.endc



.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice mc
**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
