magic
tech sky130A
timestamp 1739204916
<< nwell >>
rect 9230 2165 10840 2455
<< nmos >>
rect 9250 1805 9310 2005
rect 9360 1805 9420 2005
rect 9470 1805 9530 2005
rect 9580 1805 9640 2005
rect 9790 1805 9850 2005
rect 9900 1805 9960 2005
rect 10010 1805 10070 2005
rect 10120 1805 10180 2005
rect 10330 1805 10390 2005
rect 10440 1805 10500 2005
rect 10550 1805 10610 2005
rect 10660 1805 10720 2005
<< pmos >>
rect 9350 2235 9410 2435
rect 9460 2235 9520 2435
rect 9570 2235 9630 2435
rect 9680 2235 9740 2435
rect 9790 2235 9850 2435
rect 9900 2235 9960 2435
rect 10110 2235 10170 2435
rect 10220 2235 10280 2435
rect 10330 2235 10390 2435
rect 10440 2235 10500 2435
rect 10550 2235 10610 2435
rect 10660 2235 10720 2435
<< ndiff >>
rect 9200 1990 9250 2005
rect 9200 1970 9215 1990
rect 9235 1970 9250 1990
rect 9200 1940 9250 1970
rect 9200 1920 9215 1940
rect 9235 1920 9250 1940
rect 9200 1890 9250 1920
rect 9200 1870 9215 1890
rect 9235 1870 9250 1890
rect 9200 1840 9250 1870
rect 9200 1820 9215 1840
rect 9235 1820 9250 1840
rect 9200 1805 9250 1820
rect 9310 1990 9360 2005
rect 9310 1970 9325 1990
rect 9345 1970 9360 1990
rect 9310 1940 9360 1970
rect 9310 1920 9325 1940
rect 9345 1920 9360 1940
rect 9310 1890 9360 1920
rect 9310 1870 9325 1890
rect 9345 1870 9360 1890
rect 9310 1840 9360 1870
rect 9310 1820 9325 1840
rect 9345 1820 9360 1840
rect 9310 1805 9360 1820
rect 9420 1990 9470 2005
rect 9420 1970 9435 1990
rect 9455 1970 9470 1990
rect 9420 1940 9470 1970
rect 9420 1920 9435 1940
rect 9455 1920 9470 1940
rect 9420 1890 9470 1920
rect 9420 1870 9435 1890
rect 9455 1870 9470 1890
rect 9420 1840 9470 1870
rect 9420 1820 9435 1840
rect 9455 1820 9470 1840
rect 9420 1805 9470 1820
rect 9530 1990 9580 2005
rect 9530 1970 9545 1990
rect 9565 1970 9580 1990
rect 9530 1940 9580 1970
rect 9530 1920 9545 1940
rect 9565 1920 9580 1940
rect 9530 1890 9580 1920
rect 9530 1870 9545 1890
rect 9565 1870 9580 1890
rect 9530 1840 9580 1870
rect 9530 1820 9545 1840
rect 9565 1820 9580 1840
rect 9530 1805 9580 1820
rect 9640 1990 9690 2005
rect 9740 1990 9790 2005
rect 9640 1970 9655 1990
rect 9675 1970 9690 1990
rect 9740 1970 9755 1990
rect 9775 1970 9790 1990
rect 9640 1940 9690 1970
rect 9740 1940 9790 1970
rect 9640 1920 9655 1940
rect 9675 1920 9690 1940
rect 9740 1920 9755 1940
rect 9775 1920 9790 1940
rect 9640 1890 9690 1920
rect 9740 1890 9790 1920
rect 9640 1870 9655 1890
rect 9675 1870 9690 1890
rect 9740 1870 9755 1890
rect 9775 1870 9790 1890
rect 9640 1840 9690 1870
rect 9740 1840 9790 1870
rect 9640 1820 9655 1840
rect 9675 1820 9690 1840
rect 9740 1820 9755 1840
rect 9775 1820 9790 1840
rect 9640 1805 9690 1820
rect 9740 1805 9790 1820
rect 9850 1990 9900 2005
rect 9850 1970 9865 1990
rect 9885 1970 9900 1990
rect 9850 1940 9900 1970
rect 9850 1920 9865 1940
rect 9885 1920 9900 1940
rect 9850 1890 9900 1920
rect 9850 1870 9865 1890
rect 9885 1870 9900 1890
rect 9850 1840 9900 1870
rect 9850 1820 9865 1840
rect 9885 1820 9900 1840
rect 9850 1805 9900 1820
rect 9960 1990 10010 2005
rect 9960 1970 9975 1990
rect 9995 1970 10010 1990
rect 9960 1940 10010 1970
rect 9960 1920 9975 1940
rect 9995 1920 10010 1940
rect 9960 1890 10010 1920
rect 9960 1870 9975 1890
rect 9995 1870 10010 1890
rect 9960 1840 10010 1870
rect 9960 1820 9975 1840
rect 9995 1820 10010 1840
rect 9960 1805 10010 1820
rect 10070 1990 10120 2005
rect 10070 1970 10085 1990
rect 10105 1970 10120 1990
rect 10070 1940 10120 1970
rect 10070 1920 10085 1940
rect 10105 1920 10120 1940
rect 10070 1890 10120 1920
rect 10070 1870 10085 1890
rect 10105 1870 10120 1890
rect 10070 1840 10120 1870
rect 10070 1820 10085 1840
rect 10105 1820 10120 1840
rect 10070 1805 10120 1820
rect 10180 1990 10230 2005
rect 10280 1990 10330 2005
rect 10180 1970 10195 1990
rect 10215 1970 10230 1990
rect 10280 1970 10295 1990
rect 10315 1970 10330 1990
rect 10180 1940 10230 1970
rect 10280 1940 10330 1970
rect 10180 1920 10195 1940
rect 10215 1920 10230 1940
rect 10280 1920 10295 1940
rect 10315 1920 10330 1940
rect 10180 1890 10230 1920
rect 10280 1890 10330 1920
rect 10180 1870 10195 1890
rect 10215 1870 10230 1890
rect 10280 1870 10295 1890
rect 10315 1870 10330 1890
rect 10180 1840 10230 1870
rect 10280 1840 10330 1870
rect 10180 1820 10195 1840
rect 10215 1820 10230 1840
rect 10280 1820 10295 1840
rect 10315 1820 10330 1840
rect 10180 1805 10230 1820
rect 10280 1805 10330 1820
rect 10390 1990 10440 2005
rect 10390 1970 10405 1990
rect 10425 1970 10440 1990
rect 10390 1940 10440 1970
rect 10390 1920 10405 1940
rect 10425 1920 10440 1940
rect 10390 1890 10440 1920
rect 10390 1870 10405 1890
rect 10425 1870 10440 1890
rect 10390 1840 10440 1870
rect 10390 1820 10405 1840
rect 10425 1820 10440 1840
rect 10390 1805 10440 1820
rect 10500 1990 10550 2005
rect 10500 1970 10515 1990
rect 10535 1970 10550 1990
rect 10500 1940 10550 1970
rect 10500 1920 10515 1940
rect 10535 1920 10550 1940
rect 10500 1890 10550 1920
rect 10500 1870 10515 1890
rect 10535 1870 10550 1890
rect 10500 1840 10550 1870
rect 10500 1820 10515 1840
rect 10535 1820 10550 1840
rect 10500 1805 10550 1820
rect 10610 1990 10660 2005
rect 10610 1970 10625 1990
rect 10645 1970 10660 1990
rect 10610 1940 10660 1970
rect 10610 1920 10625 1940
rect 10645 1920 10660 1940
rect 10610 1890 10660 1920
rect 10610 1870 10625 1890
rect 10645 1870 10660 1890
rect 10610 1840 10660 1870
rect 10610 1820 10625 1840
rect 10645 1820 10660 1840
rect 10610 1805 10660 1820
rect 10720 1990 10770 2005
rect 10720 1970 10735 1990
rect 10755 1970 10770 1990
rect 10720 1940 10770 1970
rect 10720 1920 10735 1940
rect 10755 1920 10770 1940
rect 10720 1890 10770 1920
rect 10720 1870 10735 1890
rect 10755 1870 10770 1890
rect 10720 1840 10770 1870
rect 10720 1820 10735 1840
rect 10755 1820 10770 1840
rect 10720 1805 10770 1820
<< pdiff >>
rect 9300 2420 9350 2435
rect 9300 2400 9315 2420
rect 9335 2400 9350 2420
rect 9300 2370 9350 2400
rect 9300 2350 9315 2370
rect 9335 2350 9350 2370
rect 9300 2320 9350 2350
rect 9300 2300 9315 2320
rect 9335 2300 9350 2320
rect 9300 2270 9350 2300
rect 9300 2250 9315 2270
rect 9335 2250 9350 2270
rect 9300 2235 9350 2250
rect 9410 2420 9460 2435
rect 9410 2400 9425 2420
rect 9445 2400 9460 2420
rect 9410 2370 9460 2400
rect 9410 2350 9425 2370
rect 9445 2350 9460 2370
rect 9410 2320 9460 2350
rect 9410 2300 9425 2320
rect 9445 2300 9460 2320
rect 9410 2270 9460 2300
rect 9410 2250 9425 2270
rect 9445 2250 9460 2270
rect 9410 2235 9460 2250
rect 9520 2420 9570 2435
rect 9520 2400 9535 2420
rect 9555 2400 9570 2420
rect 9520 2370 9570 2400
rect 9520 2350 9535 2370
rect 9555 2350 9570 2370
rect 9520 2320 9570 2350
rect 9520 2300 9535 2320
rect 9555 2300 9570 2320
rect 9520 2270 9570 2300
rect 9520 2250 9535 2270
rect 9555 2250 9570 2270
rect 9520 2235 9570 2250
rect 9630 2420 9680 2435
rect 9630 2400 9645 2420
rect 9665 2400 9680 2420
rect 9630 2370 9680 2400
rect 9630 2350 9645 2370
rect 9665 2350 9680 2370
rect 9630 2320 9680 2350
rect 9630 2300 9645 2320
rect 9665 2300 9680 2320
rect 9630 2270 9680 2300
rect 9630 2250 9645 2270
rect 9665 2250 9680 2270
rect 9630 2235 9680 2250
rect 9740 2420 9790 2435
rect 9740 2400 9755 2420
rect 9775 2400 9790 2420
rect 9740 2370 9790 2400
rect 9740 2350 9755 2370
rect 9775 2350 9790 2370
rect 9740 2320 9790 2350
rect 9740 2300 9755 2320
rect 9775 2300 9790 2320
rect 9740 2270 9790 2300
rect 9740 2250 9755 2270
rect 9775 2250 9790 2270
rect 9740 2235 9790 2250
rect 9850 2420 9900 2435
rect 9850 2400 9865 2420
rect 9885 2400 9900 2420
rect 9850 2370 9900 2400
rect 9850 2350 9865 2370
rect 9885 2350 9900 2370
rect 9850 2320 9900 2350
rect 9850 2300 9865 2320
rect 9885 2300 9900 2320
rect 9850 2270 9900 2300
rect 9850 2250 9865 2270
rect 9885 2250 9900 2270
rect 9850 2235 9900 2250
rect 9960 2420 10010 2435
rect 10060 2420 10110 2435
rect 9960 2400 9975 2420
rect 9995 2400 10010 2420
rect 10060 2400 10075 2420
rect 10095 2400 10110 2420
rect 9960 2370 10010 2400
rect 10060 2370 10110 2400
rect 9960 2350 9975 2370
rect 9995 2350 10010 2370
rect 10060 2350 10075 2370
rect 10095 2350 10110 2370
rect 9960 2320 10010 2350
rect 10060 2320 10110 2350
rect 9960 2300 9975 2320
rect 9995 2300 10010 2320
rect 10060 2300 10075 2320
rect 10095 2300 10110 2320
rect 9960 2270 10010 2300
rect 10060 2270 10110 2300
rect 9960 2250 9975 2270
rect 9995 2250 10010 2270
rect 10060 2250 10075 2270
rect 10095 2250 10110 2270
rect 9960 2235 10010 2250
rect 10060 2235 10110 2250
rect 10170 2420 10220 2435
rect 10170 2400 10185 2420
rect 10205 2400 10220 2420
rect 10170 2370 10220 2400
rect 10170 2350 10185 2370
rect 10205 2350 10220 2370
rect 10170 2320 10220 2350
rect 10170 2300 10185 2320
rect 10205 2300 10220 2320
rect 10170 2270 10220 2300
rect 10170 2250 10185 2270
rect 10205 2250 10220 2270
rect 10170 2235 10220 2250
rect 10280 2420 10330 2435
rect 10280 2400 10295 2420
rect 10315 2400 10330 2420
rect 10280 2370 10330 2400
rect 10280 2350 10295 2370
rect 10315 2350 10330 2370
rect 10280 2320 10330 2350
rect 10280 2300 10295 2320
rect 10315 2300 10330 2320
rect 10280 2270 10330 2300
rect 10280 2250 10295 2270
rect 10315 2250 10330 2270
rect 10280 2235 10330 2250
rect 10390 2420 10440 2435
rect 10390 2400 10405 2420
rect 10425 2400 10440 2420
rect 10390 2370 10440 2400
rect 10390 2350 10405 2370
rect 10425 2350 10440 2370
rect 10390 2320 10440 2350
rect 10390 2300 10405 2320
rect 10425 2300 10440 2320
rect 10390 2270 10440 2300
rect 10390 2250 10405 2270
rect 10425 2250 10440 2270
rect 10390 2235 10440 2250
rect 10500 2420 10550 2435
rect 10500 2400 10515 2420
rect 10535 2400 10550 2420
rect 10500 2370 10550 2400
rect 10500 2350 10515 2370
rect 10535 2350 10550 2370
rect 10500 2320 10550 2350
rect 10500 2300 10515 2320
rect 10535 2300 10550 2320
rect 10500 2270 10550 2300
rect 10500 2250 10515 2270
rect 10535 2250 10550 2270
rect 10500 2235 10550 2250
rect 10610 2420 10660 2435
rect 10610 2400 10625 2420
rect 10645 2400 10660 2420
rect 10610 2370 10660 2400
rect 10610 2350 10625 2370
rect 10645 2350 10660 2370
rect 10610 2320 10660 2350
rect 10610 2300 10625 2320
rect 10645 2300 10660 2320
rect 10610 2270 10660 2300
rect 10610 2250 10625 2270
rect 10645 2250 10660 2270
rect 10610 2235 10660 2250
rect 10720 2420 10770 2435
rect 10720 2400 10735 2420
rect 10755 2400 10770 2420
rect 10720 2370 10770 2400
rect 10720 2350 10735 2370
rect 10755 2350 10770 2370
rect 10720 2320 10770 2350
rect 10720 2300 10735 2320
rect 10755 2300 10770 2320
rect 10720 2270 10770 2300
rect 10720 2250 10735 2270
rect 10755 2250 10770 2270
rect 10720 2235 10770 2250
<< ndiffc >>
rect 9215 1970 9235 1990
rect 9215 1920 9235 1940
rect 9215 1870 9235 1890
rect 9215 1820 9235 1840
rect 9325 1970 9345 1990
rect 9325 1920 9345 1940
rect 9325 1870 9345 1890
rect 9325 1820 9345 1840
rect 9435 1970 9455 1990
rect 9435 1920 9455 1940
rect 9435 1870 9455 1890
rect 9435 1820 9455 1840
rect 9545 1970 9565 1990
rect 9545 1920 9565 1940
rect 9545 1870 9565 1890
rect 9545 1820 9565 1840
rect 9655 1970 9675 1990
rect 9755 1970 9775 1990
rect 9655 1920 9675 1940
rect 9755 1920 9775 1940
rect 9655 1870 9675 1890
rect 9755 1870 9775 1890
rect 9655 1820 9675 1840
rect 9755 1820 9775 1840
rect 9865 1970 9885 1990
rect 9865 1920 9885 1940
rect 9865 1870 9885 1890
rect 9865 1820 9885 1840
rect 9975 1970 9995 1990
rect 9975 1920 9995 1940
rect 9975 1870 9995 1890
rect 9975 1820 9995 1840
rect 10085 1970 10105 1990
rect 10085 1920 10105 1940
rect 10085 1870 10105 1890
rect 10085 1820 10105 1840
rect 10195 1970 10215 1990
rect 10295 1970 10315 1990
rect 10195 1920 10215 1940
rect 10295 1920 10315 1940
rect 10195 1870 10215 1890
rect 10295 1870 10315 1890
rect 10195 1820 10215 1840
rect 10295 1820 10315 1840
rect 10405 1970 10425 1990
rect 10405 1920 10425 1940
rect 10405 1870 10425 1890
rect 10405 1820 10425 1840
rect 10515 1970 10535 1990
rect 10515 1920 10535 1940
rect 10515 1870 10535 1890
rect 10515 1820 10535 1840
rect 10625 1970 10645 1990
rect 10625 1920 10645 1940
rect 10625 1870 10645 1890
rect 10625 1820 10645 1840
rect 10735 1970 10755 1990
rect 10735 1920 10755 1940
rect 10735 1870 10755 1890
rect 10735 1820 10755 1840
<< pdiffc >>
rect 9315 2400 9335 2420
rect 9315 2350 9335 2370
rect 9315 2300 9335 2320
rect 9315 2250 9335 2270
rect 9425 2400 9445 2420
rect 9425 2350 9445 2370
rect 9425 2300 9445 2320
rect 9425 2250 9445 2270
rect 9535 2400 9555 2420
rect 9535 2350 9555 2370
rect 9535 2300 9555 2320
rect 9535 2250 9555 2270
rect 9645 2400 9665 2420
rect 9645 2350 9665 2370
rect 9645 2300 9665 2320
rect 9645 2250 9665 2270
rect 9755 2400 9775 2420
rect 9755 2350 9775 2370
rect 9755 2300 9775 2320
rect 9755 2250 9775 2270
rect 9865 2400 9885 2420
rect 9865 2350 9885 2370
rect 9865 2300 9885 2320
rect 9865 2250 9885 2270
rect 9975 2400 9995 2420
rect 10075 2400 10095 2420
rect 9975 2350 9995 2370
rect 10075 2350 10095 2370
rect 9975 2300 9995 2320
rect 10075 2300 10095 2320
rect 9975 2250 9995 2270
rect 10075 2250 10095 2270
rect 10185 2400 10205 2420
rect 10185 2350 10205 2370
rect 10185 2300 10205 2320
rect 10185 2250 10205 2270
rect 10295 2400 10315 2420
rect 10295 2350 10315 2370
rect 10295 2300 10315 2320
rect 10295 2250 10315 2270
rect 10405 2400 10425 2420
rect 10405 2350 10425 2370
rect 10405 2300 10425 2320
rect 10405 2250 10425 2270
rect 10515 2400 10535 2420
rect 10515 2350 10535 2370
rect 10515 2300 10535 2320
rect 10515 2250 10535 2270
rect 10625 2400 10645 2420
rect 10625 2350 10645 2370
rect 10625 2300 10645 2320
rect 10625 2250 10645 2270
rect 10735 2400 10755 2420
rect 10735 2350 10755 2370
rect 10735 2300 10755 2320
rect 10735 2250 10755 2270
<< psubdiff >>
rect 9150 1990 9200 2005
rect 9150 1970 9165 1990
rect 9185 1970 9200 1990
rect 9150 1940 9200 1970
rect 9150 1920 9165 1940
rect 9185 1920 9200 1940
rect 9150 1890 9200 1920
rect 9150 1870 9165 1890
rect 9185 1870 9200 1890
rect 9150 1840 9200 1870
rect 9150 1820 9165 1840
rect 9185 1820 9200 1840
rect 9150 1805 9200 1820
rect 9690 1990 9740 2005
rect 9690 1970 9705 1990
rect 9725 1970 9740 1990
rect 9690 1940 9740 1970
rect 9690 1920 9705 1940
rect 9725 1920 9740 1940
rect 9690 1890 9740 1920
rect 9690 1870 9705 1890
rect 9725 1870 9740 1890
rect 9690 1840 9740 1870
rect 9690 1820 9705 1840
rect 9725 1820 9740 1840
rect 9690 1805 9740 1820
rect 10230 1990 10280 2005
rect 10230 1970 10245 1990
rect 10265 1970 10280 1990
rect 10230 1940 10280 1970
rect 10230 1920 10245 1940
rect 10265 1920 10280 1940
rect 10230 1890 10280 1920
rect 10230 1870 10245 1890
rect 10265 1870 10280 1890
rect 10230 1840 10280 1870
rect 10230 1820 10245 1840
rect 10265 1820 10280 1840
rect 10230 1805 10280 1820
rect 10770 1990 10820 2005
rect 10770 1970 10785 1990
rect 10805 1970 10820 1990
rect 10770 1940 10820 1970
rect 10770 1920 10785 1940
rect 10805 1920 10820 1940
rect 10770 1890 10820 1920
rect 10770 1870 10785 1890
rect 10805 1870 10820 1890
rect 10770 1840 10820 1870
rect 10770 1820 10785 1840
rect 10805 1820 10820 1840
rect 10770 1805 10820 1820
<< nsubdiff >>
rect 9250 2420 9300 2435
rect 9250 2400 9265 2420
rect 9285 2400 9300 2420
rect 9250 2370 9300 2400
rect 9250 2350 9265 2370
rect 9285 2350 9300 2370
rect 9250 2320 9300 2350
rect 9250 2300 9265 2320
rect 9285 2300 9300 2320
rect 9250 2270 9300 2300
rect 9250 2250 9265 2270
rect 9285 2250 9300 2270
rect 9250 2235 9300 2250
rect 10010 2420 10060 2435
rect 10010 2400 10025 2420
rect 10045 2400 10060 2420
rect 10010 2370 10060 2400
rect 10010 2350 10025 2370
rect 10045 2350 10060 2370
rect 10010 2320 10060 2350
rect 10010 2300 10025 2320
rect 10045 2300 10060 2320
rect 10010 2270 10060 2300
rect 10010 2250 10025 2270
rect 10045 2250 10060 2270
rect 10010 2235 10060 2250
rect 10770 2420 10820 2435
rect 10770 2400 10785 2420
rect 10805 2400 10820 2420
rect 10770 2370 10820 2400
rect 10770 2350 10785 2370
rect 10805 2350 10820 2370
rect 10770 2320 10820 2350
rect 10770 2300 10785 2320
rect 10805 2300 10820 2320
rect 10770 2270 10820 2300
rect 10770 2250 10785 2270
rect 10805 2250 10820 2270
rect 10770 2235 10820 2250
<< psubdiffcont >>
rect 9165 1970 9185 1990
rect 9165 1920 9185 1940
rect 9165 1870 9185 1890
rect 9165 1820 9185 1840
rect 9705 1970 9725 1990
rect 9705 1920 9725 1940
rect 9705 1870 9725 1890
rect 9705 1820 9725 1840
rect 10245 1970 10265 1990
rect 10245 1920 10265 1940
rect 10245 1870 10265 1890
rect 10245 1820 10265 1840
rect 10785 1970 10805 1990
rect 10785 1920 10805 1940
rect 10785 1870 10805 1890
rect 10785 1820 10805 1840
<< nsubdiffcont >>
rect 9265 2400 9285 2420
rect 9265 2350 9285 2370
rect 9265 2300 9285 2320
rect 9265 2250 9285 2270
rect 10025 2400 10045 2420
rect 10025 2350 10045 2370
rect 10025 2300 10045 2320
rect 10025 2250 10045 2270
rect 10785 2400 10805 2420
rect 10785 2350 10805 2370
rect 10785 2300 10805 2320
rect 10785 2250 10805 2270
<< poly >>
rect 10505 2500 10560 2515
rect 10505 2475 10520 2500
rect 10545 2475 10560 2500
rect 10505 2460 10560 2475
rect 9350 2435 9410 2450
rect 9460 2435 9520 2450
rect 9570 2435 9630 2450
rect 9680 2435 9740 2450
rect 9790 2435 9850 2450
rect 9900 2435 9960 2450
rect 10110 2435 10170 2450
rect 10220 2445 10610 2460
rect 10220 2435 10280 2445
rect 10330 2435 10390 2445
rect 10440 2435 10500 2445
rect 10550 2435 10610 2445
rect 10660 2435 10720 2450
rect 9350 2225 9410 2235
rect 9305 2210 9410 2225
rect 9305 2190 9315 2210
rect 9335 2205 9410 2210
rect 9460 2225 9520 2235
rect 9570 2225 9630 2235
rect 9680 2225 9740 2235
rect 9790 2225 9850 2235
rect 9460 2205 9850 2225
rect 9900 2225 9960 2235
rect 10110 2225 10170 2235
rect 9900 2210 10170 2225
rect 10220 2220 10280 2235
rect 10330 2220 10390 2235
rect 10440 2220 10500 2235
rect 10550 2220 10610 2235
rect 10660 2225 10720 2235
rect 10660 2210 10765 2225
rect 9335 2190 9345 2205
rect 9305 2180 9345 2190
rect 10015 2190 10025 2210
rect 10045 2190 10055 2210
rect 10015 2180 10055 2190
rect 10725 2190 10735 2210
rect 10755 2190 10765 2210
rect 10725 2180 10765 2190
rect 9205 2050 9245 2060
rect 9205 2030 9215 2050
rect 9235 2030 9245 2050
rect 9370 2050 9410 2060
rect 9370 2030 9380 2050
rect 9400 2030 9410 2050
rect 9480 2050 9520 2060
rect 9480 2030 9490 2050
rect 9510 2030 9520 2050
rect 9695 2050 9735 2060
rect 9695 2030 9705 2050
rect 9725 2030 9735 2050
rect 10235 2050 10275 2060
rect 10235 2030 10245 2050
rect 10265 2030 10275 2050
rect 10725 2050 10765 2060
rect 10725 2030 10735 2050
rect 10755 2030 10765 2050
rect 9205 2015 9310 2030
rect 9250 2005 9310 2015
rect 9360 2015 9530 2030
rect 9360 2005 9420 2015
rect 9470 2005 9530 2015
rect 9580 2015 9850 2030
rect 9580 2005 9640 2015
rect 9790 2005 9850 2015
rect 9900 2015 10070 2030
rect 9900 2005 9960 2015
rect 10010 2005 10070 2015
rect 10120 2015 10390 2030
rect 10120 2005 10180 2015
rect 10330 2005 10390 2015
rect 10440 2005 10500 2020
rect 10550 2005 10610 2020
rect 10660 2015 10765 2030
rect 10660 2005 10720 2015
rect 9250 1790 9310 1805
rect 9360 1790 9420 1805
rect 9470 1765 9530 1805
rect 9580 1790 9640 1805
rect 9790 1790 9850 1805
rect 9900 1765 9960 1805
rect 10010 1790 10070 1805
rect 10120 1790 10180 1805
rect 10330 1790 10390 1805
rect 10440 1795 10500 1805
rect 10550 1795 10610 1805
rect 10440 1780 10610 1795
rect 10660 1790 10720 1805
rect 9470 1750 9960 1765
rect 10505 1765 10560 1780
rect 10505 1740 10520 1765
rect 10545 1740 10560 1765
rect 10505 1725 10560 1740
<< polycont >>
rect 10520 2475 10545 2500
rect 9315 2190 9335 2210
rect 10025 2190 10045 2210
rect 10735 2190 10755 2210
rect 9215 2030 9235 2050
rect 9380 2030 9400 2050
rect 9490 2030 9510 2050
rect 9705 2030 9725 2050
rect 10245 2030 10265 2050
rect 10735 2030 10755 2050
rect 10520 1740 10545 1765
<< locali >>
rect 10850 2885 10905 2895
rect 10850 2850 10860 2885
rect 10895 2850 10905 2885
rect 10850 2840 10905 2850
rect 9150 2575 9180 2595
rect 9200 2575 9230 2595
rect 9250 2575 9280 2595
rect 9300 2575 9330 2595
rect 9350 2575 9380 2595
rect 9400 2575 9430 2595
rect 9450 2575 9480 2595
rect 9500 2575 9530 2595
rect 9550 2575 9580 2595
rect 9600 2575 9630 2595
rect 9650 2575 9680 2595
rect 9700 2575 9730 2595
rect 9750 2575 9780 2595
rect 9800 2575 9830 2595
rect 9850 2575 9880 2595
rect 9900 2575 9930 2595
rect 9950 2575 9980 2595
rect 10000 2575 10030 2595
rect 10050 2575 10080 2595
rect 10100 2575 10130 2595
rect 10150 2575 10180 2595
rect 10200 2575 10230 2595
rect 10250 2575 10280 2595
rect 10300 2575 10330 2595
rect 10350 2575 10380 2595
rect 10400 2575 10430 2595
rect 10450 2575 10480 2595
rect 10500 2575 10530 2595
rect 10550 2575 10580 2595
rect 10600 2575 10630 2595
rect 10650 2575 10680 2595
rect 10700 2575 10730 2595
rect 10750 2575 10780 2595
rect 10800 2575 10835 2595
rect 9305 2430 9345 2575
rect 9255 2420 9345 2430
rect 9255 2400 9265 2420
rect 9285 2400 9315 2420
rect 9335 2400 9345 2420
rect 9255 2370 9345 2400
rect 9255 2350 9265 2370
rect 9285 2350 9315 2370
rect 9335 2350 9345 2370
rect 9255 2320 9345 2350
rect 9255 2300 9265 2320
rect 9285 2300 9315 2320
rect 9335 2300 9345 2320
rect 9255 2270 9345 2300
rect 9255 2250 9265 2270
rect 9285 2250 9315 2270
rect 9335 2250 9345 2270
rect 9255 2240 9345 2250
rect 9415 2420 9455 2575
rect 9415 2400 9425 2420
rect 9445 2400 9455 2420
rect 9415 2370 9455 2400
rect 9415 2350 9425 2370
rect 9445 2350 9455 2370
rect 9415 2320 9455 2350
rect 9415 2300 9425 2320
rect 9445 2300 9455 2320
rect 9415 2270 9455 2300
rect 9415 2250 9425 2270
rect 9445 2250 9455 2270
rect 9415 2240 9455 2250
rect 9525 2420 9565 2430
rect 9525 2400 9535 2420
rect 9555 2400 9565 2420
rect 9525 2370 9565 2400
rect 9525 2350 9535 2370
rect 9555 2350 9565 2370
rect 9525 2320 9565 2350
rect 9525 2300 9535 2320
rect 9555 2300 9565 2320
rect 9525 2270 9565 2300
rect 9525 2250 9535 2270
rect 9555 2250 9565 2270
rect 9305 2210 9345 2240
rect 9305 2190 9315 2210
rect 9335 2190 9345 2210
rect 9305 2180 9345 2190
rect 9525 2220 9565 2250
rect 9635 2420 9675 2575
rect 9635 2400 9645 2420
rect 9665 2400 9675 2420
rect 9635 2370 9675 2400
rect 9635 2350 9645 2370
rect 9665 2350 9675 2370
rect 9635 2320 9675 2350
rect 9635 2300 9645 2320
rect 9665 2300 9675 2320
rect 9635 2270 9675 2300
rect 9635 2250 9645 2270
rect 9665 2250 9675 2270
rect 9635 2240 9675 2250
rect 9745 2420 9785 2430
rect 9745 2400 9755 2420
rect 9775 2400 9785 2420
rect 9745 2370 9785 2400
rect 9745 2350 9755 2370
rect 9775 2350 9785 2370
rect 9745 2320 9785 2350
rect 9745 2300 9755 2320
rect 9775 2300 9785 2320
rect 9745 2270 9785 2300
rect 9745 2250 9755 2270
rect 9775 2250 9785 2270
rect 9745 2220 9785 2250
rect 9855 2420 9895 2575
rect 10015 2430 10055 2575
rect 9855 2400 9865 2420
rect 9885 2400 9895 2420
rect 9855 2370 9895 2400
rect 9855 2350 9865 2370
rect 9885 2350 9895 2370
rect 9855 2320 9895 2350
rect 9855 2300 9865 2320
rect 9885 2300 9895 2320
rect 9855 2270 9895 2300
rect 9855 2250 9865 2270
rect 9885 2250 9895 2270
rect 9855 2240 9895 2250
rect 9965 2420 10105 2430
rect 9965 2400 9975 2420
rect 9995 2400 10025 2420
rect 10045 2400 10075 2420
rect 10095 2400 10105 2420
rect 9965 2370 10105 2400
rect 9965 2350 9975 2370
rect 9995 2350 10025 2370
rect 10045 2350 10075 2370
rect 10095 2350 10105 2370
rect 9965 2320 10105 2350
rect 9965 2300 9975 2320
rect 9995 2300 10025 2320
rect 10045 2300 10075 2320
rect 10095 2300 10105 2320
rect 9965 2270 10105 2300
rect 9965 2250 9975 2270
rect 9995 2250 10025 2270
rect 10045 2250 10075 2270
rect 10095 2250 10105 2270
rect 9965 2240 10105 2250
rect 10175 2420 10215 2575
rect 10175 2400 10185 2420
rect 10205 2400 10215 2420
rect 10175 2370 10215 2400
rect 10175 2350 10185 2370
rect 10205 2350 10215 2370
rect 10175 2320 10215 2350
rect 10175 2300 10185 2320
rect 10205 2300 10215 2320
rect 10175 2270 10215 2300
rect 10175 2250 10185 2270
rect 10205 2250 10215 2270
rect 10175 2240 10215 2250
rect 10285 2420 10325 2430
rect 10285 2400 10295 2420
rect 10315 2400 10325 2420
rect 10285 2370 10325 2400
rect 10285 2350 10295 2370
rect 10315 2350 10325 2370
rect 10285 2320 10325 2350
rect 10285 2300 10295 2320
rect 10315 2300 10325 2320
rect 10285 2270 10325 2300
rect 10285 2250 10295 2270
rect 10315 2250 10325 2270
rect 9525 2180 9785 2220
rect 10015 2210 10055 2240
rect 10015 2190 10025 2210
rect 10045 2190 10055 2210
rect 10015 2180 10055 2190
rect 10285 2220 10325 2250
rect 10395 2420 10435 2575
rect 10505 2500 10560 2515
rect 10505 2475 10520 2500
rect 10545 2475 10560 2500
rect 10505 2460 10560 2475
rect 10395 2400 10405 2420
rect 10425 2400 10435 2420
rect 10395 2370 10435 2400
rect 10395 2350 10405 2370
rect 10425 2350 10435 2370
rect 10395 2320 10435 2350
rect 10395 2300 10405 2320
rect 10425 2300 10435 2320
rect 10395 2270 10435 2300
rect 10395 2250 10405 2270
rect 10425 2250 10435 2270
rect 10395 2240 10435 2250
rect 10505 2420 10545 2430
rect 10505 2400 10515 2420
rect 10535 2400 10545 2420
rect 10505 2370 10545 2400
rect 10505 2350 10515 2370
rect 10535 2350 10545 2370
rect 10505 2320 10545 2350
rect 10505 2300 10515 2320
rect 10535 2300 10545 2320
rect 10505 2270 10545 2300
rect 10505 2250 10515 2270
rect 10535 2250 10545 2270
rect 10505 2220 10545 2250
rect 10615 2420 10655 2575
rect 10615 2400 10625 2420
rect 10645 2400 10655 2420
rect 10615 2370 10655 2400
rect 10615 2350 10625 2370
rect 10645 2350 10655 2370
rect 10615 2320 10655 2350
rect 10615 2300 10625 2320
rect 10645 2300 10655 2320
rect 10615 2270 10655 2300
rect 10615 2250 10625 2270
rect 10645 2250 10655 2270
rect 10615 2240 10655 2250
rect 10725 2430 10765 2575
rect 10850 2505 10905 2515
rect 10850 2470 10860 2505
rect 10895 2470 10905 2505
rect 10850 2460 10905 2470
rect 10725 2420 10815 2430
rect 10725 2400 10735 2420
rect 10755 2400 10785 2420
rect 10805 2400 10815 2420
rect 10725 2370 10815 2400
rect 10725 2350 10735 2370
rect 10755 2350 10785 2370
rect 10805 2350 10815 2370
rect 10725 2320 10815 2350
rect 10725 2300 10735 2320
rect 10755 2300 10785 2320
rect 10805 2300 10815 2320
rect 10725 2270 10815 2300
rect 10725 2250 10735 2270
rect 10755 2250 10785 2270
rect 10805 2250 10815 2270
rect 10725 2240 10815 2250
rect 10285 2180 10545 2220
rect 10725 2210 10765 2240
rect 10725 2190 10735 2210
rect 10755 2190 10765 2210
rect 10725 2180 10765 2190
rect 9745 2135 9785 2180
rect 8815 2080 9410 2100
rect 9745 2095 10005 2135
rect 9370 2060 9410 2080
rect 9205 2050 9245 2060
rect 9205 2030 9215 2050
rect 9235 2030 9245 2050
rect 9205 2000 9245 2030
rect 9370 2050 9520 2060
rect 9370 2030 9380 2050
rect 9400 2030 9490 2050
rect 9510 2030 9520 2050
rect 9370 2020 9520 2030
rect 9695 2050 9735 2060
rect 9695 2030 9705 2050
rect 9725 2030 9735 2050
rect 9155 1990 9245 2000
rect 9155 1970 9165 1990
rect 9185 1970 9215 1990
rect 9235 1970 9245 1990
rect 9155 1940 9245 1970
rect 9155 1920 9165 1940
rect 9185 1920 9215 1940
rect 9235 1920 9245 1940
rect 9155 1890 9245 1920
rect 9155 1870 9165 1890
rect 9185 1870 9215 1890
rect 9235 1870 9245 1890
rect 9155 1840 9245 1870
rect 9155 1820 9165 1840
rect 9185 1820 9215 1840
rect 9235 1820 9245 1840
rect 9155 1810 9245 1820
rect 9205 1665 9245 1810
rect 9315 1990 9355 2000
rect 9315 1970 9325 1990
rect 9345 1970 9355 1990
rect 9315 1940 9355 1970
rect 9315 1920 9325 1940
rect 9345 1920 9355 1940
rect 9315 1890 9355 1920
rect 9315 1870 9325 1890
rect 9345 1870 9355 1890
rect 9315 1840 9355 1870
rect 9315 1820 9325 1840
rect 9345 1820 9355 1840
rect 9315 1665 9355 1820
rect 9425 1990 9465 2020
rect 9695 2000 9735 2030
rect 9425 1970 9435 1990
rect 9455 1970 9465 1990
rect 9425 1940 9465 1970
rect 9425 1920 9435 1940
rect 9455 1920 9465 1940
rect 9425 1890 9465 1920
rect 9425 1870 9435 1890
rect 9455 1870 9465 1890
rect 9425 1840 9465 1870
rect 9425 1820 9435 1840
rect 9455 1820 9465 1840
rect 9425 1810 9465 1820
rect 9535 1990 9575 2000
rect 9535 1970 9545 1990
rect 9565 1970 9575 1990
rect 9535 1940 9575 1970
rect 9535 1920 9545 1940
rect 9565 1920 9575 1940
rect 9535 1890 9575 1920
rect 9535 1870 9545 1890
rect 9565 1870 9575 1890
rect 9535 1840 9575 1870
rect 9535 1820 9545 1840
rect 9565 1820 9575 1840
rect 9535 1665 9575 1820
rect 9645 1990 9785 2000
rect 9645 1970 9655 1990
rect 9675 1970 9705 1990
rect 9725 1970 9755 1990
rect 9775 1970 9785 1990
rect 9645 1940 9785 1970
rect 9645 1920 9655 1940
rect 9675 1920 9705 1940
rect 9725 1920 9755 1940
rect 9775 1920 9785 1940
rect 9645 1890 9785 1920
rect 9645 1870 9655 1890
rect 9675 1870 9705 1890
rect 9725 1870 9755 1890
rect 9775 1870 9785 1890
rect 9645 1840 9785 1870
rect 9645 1820 9655 1840
rect 9675 1820 9705 1840
rect 9725 1820 9755 1840
rect 9775 1820 9785 1840
rect 9645 1810 9785 1820
rect 9855 1990 9895 2000
rect 9855 1970 9865 1990
rect 9885 1970 9895 1990
rect 9855 1940 9895 1970
rect 9855 1920 9865 1940
rect 9885 1920 9895 1940
rect 9855 1890 9895 1920
rect 9855 1870 9865 1890
rect 9885 1870 9895 1890
rect 9855 1840 9895 1870
rect 9855 1820 9865 1840
rect 9885 1820 9895 1840
rect 9695 1665 9735 1810
rect 9855 1665 9895 1820
rect 9965 1990 10005 2095
rect 10235 2050 10275 2060
rect 10235 2030 10245 2050
rect 10265 2030 10275 2050
rect 10235 2000 10275 2030
rect 9965 1970 9975 1990
rect 9995 1970 10005 1990
rect 9965 1940 10005 1970
rect 9965 1920 9975 1940
rect 9995 1920 10005 1940
rect 9965 1890 10005 1920
rect 9965 1870 9975 1890
rect 9995 1870 10005 1890
rect 9965 1840 10005 1870
rect 9965 1820 9975 1840
rect 9995 1820 10005 1840
rect 9965 1810 10005 1820
rect 10075 1990 10115 2000
rect 10075 1970 10085 1990
rect 10105 1970 10115 1990
rect 10075 1940 10115 1970
rect 10075 1920 10085 1940
rect 10105 1920 10115 1940
rect 10075 1890 10115 1920
rect 10075 1870 10085 1890
rect 10105 1870 10115 1890
rect 10075 1840 10115 1870
rect 10075 1820 10085 1840
rect 10105 1820 10115 1840
rect 10075 1665 10115 1820
rect 10185 1990 10325 2000
rect 10185 1970 10195 1990
rect 10215 1970 10245 1990
rect 10265 1970 10295 1990
rect 10315 1970 10325 1990
rect 10185 1940 10325 1970
rect 10185 1920 10195 1940
rect 10215 1920 10245 1940
rect 10265 1920 10295 1940
rect 10315 1920 10325 1940
rect 10185 1890 10325 1920
rect 10185 1870 10195 1890
rect 10215 1870 10245 1890
rect 10265 1870 10295 1890
rect 10315 1870 10325 1890
rect 10185 1840 10325 1870
rect 10185 1820 10195 1840
rect 10215 1820 10245 1840
rect 10265 1820 10295 1840
rect 10315 1820 10325 1840
rect 10185 1810 10325 1820
rect 10395 1990 10435 2000
rect 10395 1970 10405 1990
rect 10425 1970 10435 1990
rect 10395 1940 10435 1970
rect 10395 1920 10405 1940
rect 10425 1920 10435 1940
rect 10395 1890 10435 1920
rect 10395 1870 10405 1890
rect 10425 1870 10435 1890
rect 10395 1840 10435 1870
rect 10395 1820 10405 1840
rect 10425 1820 10435 1840
rect 10235 1665 10275 1810
rect 10395 1665 10435 1820
rect 10505 1990 10545 2180
rect 10725 2050 10765 2060
rect 10725 2030 10735 2050
rect 10755 2030 10765 2050
rect 10725 2000 10765 2030
rect 10505 1970 10515 1990
rect 10535 1970 10545 1990
rect 10505 1940 10545 1970
rect 10505 1920 10515 1940
rect 10535 1920 10545 1940
rect 10505 1890 10545 1920
rect 10505 1870 10515 1890
rect 10535 1870 10545 1890
rect 10505 1840 10545 1870
rect 10505 1820 10515 1840
rect 10535 1820 10545 1840
rect 10505 1810 10545 1820
rect 10615 1990 10655 2000
rect 10615 1970 10625 1990
rect 10645 1970 10655 1990
rect 10615 1940 10655 1970
rect 10615 1920 10625 1940
rect 10645 1920 10655 1940
rect 10615 1890 10655 1920
rect 10615 1870 10625 1890
rect 10645 1870 10655 1890
rect 10615 1840 10655 1870
rect 10615 1820 10625 1840
rect 10645 1820 10655 1840
rect 10505 1765 10560 1780
rect 10505 1740 10520 1765
rect 10545 1740 10560 1765
rect 10505 1725 10560 1740
rect 10615 1665 10655 1820
rect 10725 1990 10815 2000
rect 10725 1970 10735 1990
rect 10755 1970 10785 1990
rect 10805 1970 10815 1990
rect 10725 1940 10815 1970
rect 10725 1920 10735 1940
rect 10755 1920 10785 1940
rect 10805 1920 10815 1940
rect 10725 1890 10815 1920
rect 10725 1870 10735 1890
rect 10755 1870 10785 1890
rect 10805 1870 10815 1890
rect 10725 1840 10815 1870
rect 10725 1820 10735 1840
rect 10755 1820 10785 1840
rect 10805 1820 10815 1840
rect 10725 1810 10815 1820
rect 10725 1665 10765 1810
rect 10890 1770 10945 1780
rect 10890 1735 10900 1770
rect 10935 1735 10945 1770
rect 10890 1725 10945 1735
rect 9155 1645 9185 1665
rect 9205 1645 9235 1665
rect 9255 1645 9285 1665
rect 9305 1645 9335 1665
rect 9355 1645 9385 1665
rect 9405 1645 9435 1665
rect 9455 1645 9485 1665
rect 9505 1645 9535 1665
rect 9555 1645 9585 1665
rect 9605 1645 9635 1665
rect 9655 1645 9685 1665
rect 9705 1645 9735 1665
rect 9755 1645 9785 1665
rect 9805 1645 9835 1665
rect 9855 1645 9885 1665
rect 9905 1645 9935 1665
rect 9955 1645 9985 1665
rect 10005 1645 10035 1665
rect 10055 1645 10085 1665
rect 10105 1645 10135 1665
rect 10155 1645 10185 1665
rect 10205 1645 10235 1665
rect 10255 1645 10285 1665
rect 10305 1645 10335 1665
rect 10355 1645 10385 1665
rect 10405 1645 10435 1665
rect 10455 1645 10485 1665
rect 10505 1645 10535 1665
rect 10555 1645 10585 1665
rect 10605 1645 10635 1665
rect 10655 1645 10685 1665
rect 10705 1645 10735 1665
rect 10755 1645 10785 1665
rect 10805 1645 10840 1665
rect 10890 1550 10945 1560
rect 10890 1515 10900 1550
rect 10935 1515 10945 1550
rect 10890 1505 10945 1515
<< viali >>
rect 10860 2850 10895 2885
rect 9180 2575 9200 2595
rect 9230 2575 9250 2595
rect 9280 2575 9300 2595
rect 9330 2575 9350 2595
rect 9380 2575 9400 2595
rect 9430 2575 9450 2595
rect 9480 2575 9500 2595
rect 9530 2575 9550 2595
rect 9580 2575 9600 2595
rect 9630 2575 9650 2595
rect 9680 2575 9700 2595
rect 9730 2575 9750 2595
rect 9780 2575 9800 2595
rect 9830 2575 9850 2595
rect 9880 2575 9900 2595
rect 9930 2575 9950 2595
rect 9980 2575 10000 2595
rect 10030 2575 10050 2595
rect 10080 2575 10100 2595
rect 10130 2575 10150 2595
rect 10180 2575 10200 2595
rect 10230 2575 10250 2595
rect 10280 2575 10300 2595
rect 10330 2575 10350 2595
rect 10380 2575 10400 2595
rect 10430 2575 10450 2595
rect 10480 2575 10500 2595
rect 10530 2575 10550 2595
rect 10580 2575 10600 2595
rect 10630 2575 10650 2595
rect 10680 2575 10700 2595
rect 10730 2575 10750 2595
rect 10780 2575 10800 2595
rect 10520 2475 10545 2500
rect 10860 2470 10895 2505
rect 10520 1740 10545 1765
rect 10900 1735 10935 1770
rect 9185 1645 9205 1665
rect 9235 1645 9255 1665
rect 9285 1645 9305 1665
rect 9335 1645 9355 1665
rect 9385 1645 9405 1665
rect 9435 1645 9455 1665
rect 9485 1645 9505 1665
rect 9535 1645 9555 1665
rect 9585 1645 9605 1665
rect 9635 1645 9655 1665
rect 9685 1645 9705 1665
rect 9735 1645 9755 1665
rect 9785 1645 9805 1665
rect 9835 1645 9855 1665
rect 9885 1645 9905 1665
rect 9935 1645 9955 1665
rect 9985 1645 10005 1665
rect 10035 1645 10055 1665
rect 10085 1645 10105 1665
rect 10135 1645 10155 1665
rect 10185 1645 10205 1665
rect 10235 1645 10255 1665
rect 10285 1645 10305 1665
rect 10335 1645 10355 1665
rect 10385 1645 10405 1665
rect 10435 1645 10455 1665
rect 10485 1645 10505 1665
rect 10535 1645 10555 1665
rect 10585 1645 10605 1665
rect 10635 1645 10655 1665
rect 10685 1645 10705 1665
rect 10735 1645 10755 1665
rect 10785 1645 10805 1665
rect 10900 1515 10935 1550
<< metal1 >>
rect 8205 2885 10905 2895
rect 8205 2850 10860 2885
rect 10895 2850 10905 2885
rect 8205 2840 10905 2850
rect 9150 2595 10835 2605
rect 9150 2575 9180 2595
rect 9200 2575 9230 2595
rect 9250 2575 9280 2595
rect 9300 2575 9330 2595
rect 9350 2575 9380 2595
rect 9400 2575 9430 2595
rect 9450 2575 9480 2595
rect 9500 2575 9530 2595
rect 9550 2575 9580 2595
rect 9600 2575 9630 2595
rect 9650 2575 9680 2595
rect 9700 2575 9730 2595
rect 9750 2575 9780 2595
rect 9800 2575 9830 2595
rect 9850 2575 9880 2595
rect 9900 2575 9930 2595
rect 9950 2575 9980 2595
rect 10000 2575 10030 2595
rect 10050 2575 10080 2595
rect 10100 2575 10130 2595
rect 10150 2575 10180 2595
rect 10200 2575 10230 2595
rect 10250 2575 10280 2595
rect 10300 2575 10330 2595
rect 10350 2575 10380 2595
rect 10400 2575 10430 2595
rect 10450 2575 10480 2595
rect 10500 2575 10530 2595
rect 10550 2575 10580 2595
rect 10600 2575 10630 2595
rect 10650 2575 10680 2595
rect 10700 2575 10730 2595
rect 10750 2575 10780 2595
rect 10800 2575 10835 2595
rect 9150 2565 10835 2575
rect 10505 2505 10905 2515
rect 10505 2500 10860 2505
rect 10505 2475 10520 2500
rect 10545 2475 10860 2500
rect 10505 2470 10860 2475
rect 10895 2470 10905 2505
rect 10505 2460 10905 2470
rect 10505 1770 10945 1780
rect 10505 1765 10900 1770
rect 10505 1740 10520 1765
rect 10545 1740 10900 1765
rect 10505 1735 10900 1740
rect 10935 1735 10945 1770
rect 10505 1725 10945 1735
rect 9155 1665 10840 1675
rect 9155 1645 9185 1665
rect 9205 1645 9235 1665
rect 9255 1645 9285 1665
rect 9305 1645 9335 1665
rect 9355 1645 9385 1665
rect 9405 1645 9435 1665
rect 9455 1645 9485 1665
rect 9505 1645 9535 1665
rect 9555 1645 9585 1665
rect 9605 1645 9635 1665
rect 9655 1645 9685 1665
rect 9705 1645 9735 1665
rect 9755 1645 9785 1665
rect 9805 1645 9835 1665
rect 9855 1645 9885 1665
rect 9905 1645 9935 1665
rect 9955 1645 9985 1665
rect 10005 1645 10035 1665
rect 10055 1645 10085 1665
rect 10105 1645 10135 1665
rect 10155 1645 10185 1665
rect 10205 1645 10235 1665
rect 10255 1645 10285 1665
rect 10305 1645 10335 1665
rect 10355 1645 10385 1665
rect 10405 1645 10435 1665
rect 10455 1645 10485 1665
rect 10505 1645 10535 1665
rect 10555 1645 10585 1665
rect 10605 1645 10635 1665
rect 10655 1645 10685 1665
rect 10705 1645 10735 1665
rect 10755 1645 10785 1665
rect 10805 1645 10840 1665
rect 9155 1635 10840 1645
rect 8250 1550 10945 1560
rect 8250 1515 10900 1550
rect 10935 1515 10945 1550
rect 8250 1505 10945 1515
<< via1 >>
rect 10860 2850 10895 2885
rect 10860 2470 10895 2505
rect 10900 1735 10935 1770
rect 10900 1515 10935 1550
<< metal2 >>
rect 10850 2885 10905 2895
rect 10850 2850 10860 2885
rect 10895 2850 10905 2885
rect 10850 2840 10905 2850
rect 10850 2505 10905 2515
rect 10850 2470 10860 2505
rect 10895 2470 10905 2505
rect 10850 2460 10905 2470
rect 10890 1770 10945 1780
rect 10890 1735 10900 1770
rect 10935 1735 10945 1770
rect 10890 1725 10945 1735
rect 10890 1550 10945 1560
rect 10890 1515 10900 1550
rect 10935 1515 10945 1550
rect 10890 1505 10945 1515
<< via2 >>
rect 10860 2850 10895 2885
rect 10860 2470 10895 2505
rect 10900 1735 10935 1770
rect 10900 1515 10935 1550
<< metal3 >>
rect 10850 2885 11655 2895
rect 10850 2850 10860 2885
rect 10895 2850 11655 2885
rect 10850 2840 11655 2850
rect 10850 2505 10905 2515
rect 10850 2470 10860 2505
rect 10895 2470 10905 2505
rect 10850 2460 10905 2470
rect 11025 2445 11655 2840
rect 10890 1770 10945 1780
rect 10890 1735 10900 1770
rect 10935 1735 10945 1770
rect 10890 1725 10945 1735
rect 11065 1560 11355 1795
rect 10890 1550 11355 1560
rect 10890 1515 10900 1550
rect 10935 1515 11355 1550
rect 10890 1505 11355 1515
<< via3 >>
rect 10860 2470 10895 2505
rect 10900 1735 10935 1770
<< mimcap >>
rect 11040 2505 11640 2880
rect 11040 2470 11050 2505
rect 11085 2470 11640 2505
rect 11040 2460 11640 2470
rect 11080 1770 11340 1780
rect 11080 1735 11090 1770
rect 11125 1735 11340 1770
rect 11080 1520 11340 1735
<< mimcapcontact >>
rect 11050 2470 11085 2505
rect 11090 1735 11125 1770
<< metal4 >>
rect 10850 2505 11095 2515
rect 10850 2470 10860 2505
rect 10895 2470 11050 2505
rect 11085 2470 11095 2505
rect 10850 2460 11095 2470
rect 10890 1770 11135 1780
rect 10890 1735 10900 1770
rect 10935 1735 11090 1770
rect 11125 1735 11135 1770
rect 10890 1725 11135 1735
<< labels >>
flabel locali 8815 2090 8815 2090 7 FreeSans 400 0 -200 0 I_IN
port 3 w
flabel locali 10545 2105 10545 2105 3 FreeSans 400 0 160 0 vout
port 6 e
flabel locali 10005 2120 10005 2120 3 FreeSans 400 0 200 0 x
flabel metal1 9150 2585 9150 2585 7 FreeSans 400 0 -200 0 VDDA
port 1 w
flabel metal1 9155 1655 9155 1655 7 FreeSans 400 0 -200 0 GNDA
port 2 w
flabel poly 9460 2205 9460 2205 5 FreeSans 400 0 0 -200 opamp_out
flabel metal1 10530 1725 10530 1725 5 FreeSans 400 0 0 -200 DOWN_input
port 8 s
flabel metal1 8250 1530 8250 1530 7 FreeSans 400 0 -200 0 DOWN
port 5 w
flabel metal1 10530 2515 10530 2515 1 FreeSans 400 0 0 200 UP_input
port 7 n
flabel metal1 8205 2865 8205 2865 7 FreeSans 400 0 -200 0 UP_b
port 4 w
<< end >>
