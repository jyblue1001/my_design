magic
tech sky130A
timestamp 1738582453
<< nwell >>
rect -60 140 2525 280
<< nmos >>
rect 0 0 15 50
rect 55 0 70 50
rect 260 0 275 50
rect 315 0 330 50
rect 440 0 455 50
rect 495 0 510 50
rect 700 0 715 50
rect 755 0 770 50
rect 880 0 895 50
rect 935 0 950 50
rect 1140 0 1155 50
rect 1195 0 1210 50
rect 1330 0 1345 50
rect 1385 0 1400 50
rect 1590 0 1605 50
rect 1645 0 1660 50
rect 1770 0 1785 50
rect 1825 0 1840 50
rect 1950 0 1965 50
rect 2075 0 2090 50
rect 2200 0 2215 50
rect 2325 0 2340 50
rect 2450 0 2465 50
<< pmos >>
rect 0 160 15 260
rect 55 160 70 260
rect 260 160 275 260
rect 315 160 330 260
rect 440 160 455 260
rect 495 160 510 260
rect 700 160 715 260
rect 755 160 770 260
rect 880 160 895 260
rect 935 160 950 260
rect 1140 160 1155 260
rect 1195 160 1210 260
rect 1330 160 1345 260
rect 1385 160 1400 260
rect 1590 160 1605 260
rect 1645 160 1660 260
rect 1770 160 1785 260
rect 1825 160 1840 260
rect 1950 160 1965 260
rect 2075 160 2090 260
rect 2200 160 2215 260
rect 2325 160 2340 260
rect 2450 160 2465 260
<< ndiff >>
rect -40 35 0 50
rect -40 15 -30 35
rect -10 15 0 35
rect -40 0 0 15
rect 15 35 55 50
rect 15 15 25 35
rect 45 15 55 35
rect 15 0 55 15
rect 70 35 110 50
rect 70 15 80 35
rect 100 15 110 35
rect 70 0 110 15
rect 220 35 260 50
rect 220 15 230 35
rect 250 15 260 35
rect 220 0 260 15
rect 275 35 315 50
rect 275 15 285 35
rect 305 15 315 35
rect 275 0 315 15
rect 330 35 370 50
rect 330 15 340 35
rect 360 15 370 35
rect 330 0 370 15
rect 400 35 440 50
rect 400 15 410 35
rect 430 15 440 35
rect 400 0 440 15
rect 455 35 495 50
rect 455 15 465 35
rect 485 15 495 35
rect 455 0 495 15
rect 510 35 550 50
rect 510 15 520 35
rect 540 15 550 35
rect 510 0 550 15
rect 660 35 700 50
rect 660 15 670 35
rect 690 15 700 35
rect 660 0 700 15
rect 715 35 755 50
rect 715 15 725 35
rect 745 15 755 35
rect 715 0 755 15
rect 770 35 810 50
rect 770 15 780 35
rect 800 15 810 35
rect 770 0 810 15
rect 840 35 880 50
rect 840 15 850 35
rect 870 15 880 35
rect 840 0 880 15
rect 895 35 935 50
rect 895 15 905 35
rect 925 15 935 35
rect 895 0 935 15
rect 950 35 990 50
rect 950 15 960 35
rect 980 15 990 35
rect 950 0 990 15
rect 1100 35 1140 50
rect 1100 15 1110 35
rect 1130 15 1140 35
rect 1100 0 1140 15
rect 1155 35 1195 50
rect 1155 15 1165 35
rect 1185 15 1195 35
rect 1155 0 1195 15
rect 1210 35 1250 50
rect 1290 35 1330 50
rect 1210 15 1220 35
rect 1240 15 1250 35
rect 1290 15 1300 35
rect 1320 15 1330 35
rect 1210 0 1250 15
rect 1290 0 1330 15
rect 1345 35 1385 50
rect 1345 15 1355 35
rect 1375 15 1385 35
rect 1345 0 1385 15
rect 1400 35 1440 50
rect 1400 15 1410 35
rect 1430 15 1440 35
rect 1400 0 1440 15
rect 1550 35 1590 50
rect 1550 15 1560 35
rect 1580 15 1590 35
rect 1550 0 1590 15
rect 1605 35 1645 50
rect 1605 15 1615 35
rect 1635 15 1645 35
rect 1605 0 1645 15
rect 1660 35 1700 50
rect 1660 15 1670 35
rect 1690 15 1700 35
rect 1660 0 1700 15
rect 1730 35 1770 50
rect 1730 15 1740 35
rect 1760 15 1770 35
rect 1730 0 1770 15
rect 1785 35 1825 50
rect 1785 15 1795 35
rect 1815 15 1825 35
rect 1785 0 1825 15
rect 1840 35 1880 50
rect 1840 15 1850 35
rect 1870 15 1880 35
rect 1840 0 1880 15
rect 1910 35 1950 50
rect 1910 15 1920 35
rect 1940 15 1950 35
rect 1910 0 1950 15
rect 1965 35 2005 50
rect 1965 15 1975 35
rect 1995 15 2005 35
rect 1965 0 2005 15
rect 2035 35 2075 50
rect 2035 15 2045 35
rect 2065 15 2075 35
rect 2035 0 2075 15
rect 2090 35 2130 50
rect 2090 15 2100 35
rect 2120 15 2130 35
rect 2090 0 2130 15
rect 2160 35 2200 50
rect 2160 15 2170 35
rect 2190 15 2200 35
rect 2160 0 2200 15
rect 2215 35 2255 50
rect 2215 15 2225 35
rect 2245 15 2255 35
rect 2215 0 2255 15
rect 2285 35 2325 50
rect 2285 15 2295 35
rect 2315 15 2325 35
rect 2285 0 2325 15
rect 2340 35 2380 50
rect 2340 15 2350 35
rect 2370 15 2380 35
rect 2340 0 2380 15
rect 2410 35 2450 50
rect 2410 15 2420 35
rect 2440 15 2450 35
rect 2410 0 2450 15
rect 2465 35 2505 50
rect 2465 15 2475 35
rect 2495 15 2505 35
rect 2465 0 2505 15
<< pdiff >>
rect -40 245 0 260
rect -40 175 -30 245
rect -10 175 0 245
rect -40 160 0 175
rect 15 245 55 260
rect 15 175 25 245
rect 45 175 55 245
rect 15 160 55 175
rect 70 245 110 260
rect 70 175 80 245
rect 100 175 110 245
rect 70 160 110 175
rect 220 245 260 260
rect 220 175 230 245
rect 250 175 260 245
rect 220 160 260 175
rect 275 245 315 260
rect 275 175 285 245
rect 305 175 315 245
rect 275 160 315 175
rect 330 245 370 260
rect 330 175 340 245
rect 360 175 370 245
rect 330 160 370 175
rect 400 245 440 260
rect 400 175 410 245
rect 430 175 440 245
rect 400 160 440 175
rect 455 245 495 260
rect 455 175 465 245
rect 485 175 495 245
rect 455 160 495 175
rect 510 245 550 260
rect 510 175 520 245
rect 540 175 550 245
rect 510 160 550 175
rect 660 245 700 260
rect 660 175 670 245
rect 690 175 700 245
rect 660 160 700 175
rect 715 245 755 260
rect 715 175 725 245
rect 745 175 755 245
rect 715 160 755 175
rect 770 245 810 260
rect 770 175 780 245
rect 800 175 810 245
rect 770 160 810 175
rect 840 245 880 260
rect 840 175 850 245
rect 870 175 880 245
rect 840 160 880 175
rect 895 245 935 260
rect 895 175 905 245
rect 925 175 935 245
rect 895 160 935 175
rect 950 245 990 260
rect 950 175 960 245
rect 980 175 990 245
rect 950 160 990 175
rect 1100 245 1140 260
rect 1100 175 1110 245
rect 1130 175 1140 245
rect 1100 160 1140 175
rect 1155 245 1195 260
rect 1155 175 1165 245
rect 1185 175 1195 245
rect 1155 160 1195 175
rect 1210 245 1250 260
rect 1290 245 1330 260
rect 1210 175 1220 245
rect 1240 175 1250 245
rect 1290 175 1300 245
rect 1320 175 1330 245
rect 1210 160 1250 175
rect 1290 160 1330 175
rect 1345 245 1385 260
rect 1345 175 1355 245
rect 1375 175 1385 245
rect 1345 160 1385 175
rect 1400 245 1440 260
rect 1400 175 1410 245
rect 1430 175 1440 245
rect 1400 160 1440 175
rect 1550 245 1590 260
rect 1550 175 1560 245
rect 1580 175 1590 245
rect 1550 160 1590 175
rect 1605 245 1645 260
rect 1605 175 1615 245
rect 1635 175 1645 245
rect 1605 160 1645 175
rect 1660 245 1700 260
rect 1660 175 1670 245
rect 1690 175 1700 245
rect 1660 160 1700 175
rect 1730 245 1770 260
rect 1730 175 1740 245
rect 1760 175 1770 245
rect 1730 160 1770 175
rect 1785 245 1825 260
rect 1785 175 1795 245
rect 1815 175 1825 245
rect 1785 160 1825 175
rect 1840 245 1880 260
rect 1840 175 1850 245
rect 1870 175 1880 245
rect 1840 160 1880 175
rect 1910 245 1950 260
rect 1910 175 1920 245
rect 1940 175 1950 245
rect 1910 160 1950 175
rect 1965 245 2005 260
rect 1965 175 1975 245
rect 1995 175 2005 245
rect 1965 160 2005 175
rect 2035 245 2075 260
rect 2035 175 2045 245
rect 2065 175 2075 245
rect 2035 160 2075 175
rect 2090 245 2130 260
rect 2090 175 2100 245
rect 2120 175 2130 245
rect 2090 160 2130 175
rect 2160 245 2200 260
rect 2160 175 2170 245
rect 2190 175 2200 245
rect 2160 160 2200 175
rect 2215 245 2255 260
rect 2215 175 2225 245
rect 2245 175 2255 245
rect 2215 160 2255 175
rect 2285 245 2325 260
rect 2285 175 2295 245
rect 2315 175 2325 245
rect 2285 160 2325 175
rect 2340 245 2380 260
rect 2340 175 2350 245
rect 2370 175 2380 245
rect 2340 160 2380 175
rect 2410 245 2450 260
rect 2410 175 2420 245
rect 2440 175 2450 245
rect 2410 160 2450 175
rect 2465 245 2505 260
rect 2465 175 2475 245
rect 2495 175 2505 245
rect 2465 160 2505 175
<< ndiffc >>
rect -30 15 -10 35
rect 25 15 45 35
rect 80 15 100 35
rect 230 15 250 35
rect 285 15 305 35
rect 340 15 360 35
rect 410 15 430 35
rect 465 15 485 35
rect 520 15 540 35
rect 670 15 690 35
rect 725 15 745 35
rect 780 15 800 35
rect 850 15 870 35
rect 905 15 925 35
rect 960 15 980 35
rect 1110 15 1130 35
rect 1165 15 1185 35
rect 1220 15 1240 35
rect 1300 15 1320 35
rect 1355 15 1375 35
rect 1410 15 1430 35
rect 1560 15 1580 35
rect 1615 15 1635 35
rect 1670 15 1690 35
rect 1740 15 1760 35
rect 1795 15 1815 35
rect 1850 15 1870 35
rect 1920 15 1940 35
rect 1975 15 1995 35
rect 2045 15 2065 35
rect 2100 15 2120 35
rect 2170 15 2190 35
rect 2225 15 2245 35
rect 2295 15 2315 35
rect 2350 15 2370 35
rect 2420 15 2440 35
rect 2475 15 2495 35
<< pdiffc >>
rect -30 175 -10 245
rect 25 175 45 245
rect 80 175 100 245
rect 230 175 250 245
rect 285 175 305 245
rect 340 175 360 245
rect 410 175 430 245
rect 465 175 485 245
rect 520 175 540 245
rect 670 175 690 245
rect 725 175 745 245
rect 780 175 800 245
rect 850 175 870 245
rect 905 175 925 245
rect 960 175 980 245
rect 1110 175 1130 245
rect 1165 175 1185 245
rect 1220 175 1240 245
rect 1300 175 1320 245
rect 1355 175 1375 245
rect 1410 175 1430 245
rect 1560 175 1580 245
rect 1615 175 1635 245
rect 1670 175 1690 245
rect 1740 175 1760 245
rect 1795 175 1815 245
rect 1850 175 1870 245
rect 1920 175 1940 245
rect 1975 175 1995 245
rect 2045 175 2065 245
rect 2100 175 2120 245
rect 2170 175 2190 245
rect 2225 175 2245 245
rect 2295 175 2315 245
rect 2350 175 2370 245
rect 2420 175 2440 245
rect 2475 175 2495 245
<< psubdiff >>
rect 1250 35 1290 50
rect 1250 15 1260 35
rect 1280 15 1290 35
rect 1250 0 1290 15
<< nsubdiff >>
rect 1250 245 1290 260
rect 1250 175 1260 245
rect 1280 175 1290 245
rect 1250 160 1290 175
<< psubdiffcont >>
rect 1260 15 1280 35
<< nsubdiffcont >>
rect 1260 175 1280 245
<< poly >>
rect 755 340 2530 355
rect 185 305 225 315
rect 185 285 195 305
rect 215 285 225 305
rect 185 275 225 285
rect 0 260 15 275
rect 55 260 70 275
rect 260 260 275 275
rect 315 260 330 275
rect 440 260 455 275
rect 495 260 510 275
rect 700 260 715 275
rect 755 260 770 340
rect 880 260 895 275
rect 935 260 950 275
rect 1140 260 1155 275
rect 1195 260 1210 275
rect 1330 260 1345 275
rect 1385 260 1400 275
rect 1590 260 1605 275
rect 1645 260 1660 340
rect 1745 305 1785 315
rect 1745 285 1755 305
rect 1775 285 1785 305
rect 1745 275 1785 285
rect 1770 260 1785 275
rect 1825 260 1840 275
rect 1950 260 1965 275
rect 2075 260 2090 275
rect 2200 260 2215 275
rect 2325 260 2340 275
rect 2450 260 2465 275
rect 125 245 165 255
rect 125 225 135 245
rect 155 225 165 245
rect 125 215 165 225
rect 0 100 15 160
rect -60 85 15 100
rect 0 50 15 85
rect 55 105 70 160
rect 55 95 105 105
rect 55 75 75 95
rect 95 75 105 95
rect 55 65 105 75
rect 150 85 165 215
rect 565 245 605 255
rect 565 225 575 245
rect 595 225 605 245
rect 565 215 605 225
rect 260 85 275 160
rect 150 70 275 85
rect 55 50 70 65
rect 260 50 275 70
rect 315 145 330 160
rect 315 135 365 145
rect 315 115 335 135
rect 355 115 365 135
rect 315 105 365 115
rect 315 50 330 105
rect 440 50 455 160
rect 495 105 510 160
rect 495 95 545 105
rect 495 75 515 95
rect 535 75 545 95
rect 495 65 545 75
rect 590 85 605 215
rect 1005 245 1045 255
rect 1005 225 1015 245
rect 1035 225 1045 245
rect 1005 215 1045 225
rect 700 85 715 160
rect 590 70 715 85
rect 495 50 510 65
rect 700 50 715 70
rect 755 50 770 160
rect 880 50 895 160
rect 935 105 950 160
rect 935 95 985 105
rect 935 75 955 95
rect 975 75 985 95
rect 935 65 985 75
rect 1030 85 1045 215
rect 1455 245 1495 255
rect 1455 225 1465 245
rect 1485 225 1495 245
rect 1455 215 1495 225
rect 1140 85 1155 160
rect 1030 70 1155 85
rect 935 50 950 65
rect 1140 50 1155 70
rect 1195 145 1210 160
rect 1195 135 1245 145
rect 1195 115 1215 135
rect 1235 115 1245 135
rect 1195 105 1245 115
rect 1195 50 1210 105
rect 1330 50 1345 160
rect 1385 105 1400 160
rect 1385 95 1435 105
rect 1385 75 1405 95
rect 1425 75 1435 95
rect 1385 65 1435 75
rect 1480 85 1495 215
rect 1590 85 1605 160
rect 1480 70 1605 85
rect 1385 50 1400 65
rect 1590 50 1605 70
rect 1645 50 1660 160
rect 1770 50 1785 160
rect 1825 50 1840 160
rect 1865 120 1905 130
rect 1865 100 1875 120
rect 1895 115 1905 120
rect 1950 115 1965 160
rect 1895 100 1965 115
rect 1865 90 1905 100
rect 1950 50 1965 100
rect 1990 120 2030 130
rect 1990 100 2000 120
rect 2020 115 2030 120
rect 2075 115 2090 160
rect 2020 100 2090 115
rect 1990 90 2030 100
rect 2075 50 2090 100
rect 2115 120 2155 130
rect 2115 100 2125 120
rect 2145 115 2155 120
rect 2200 115 2215 160
rect 2145 100 2215 115
rect 2115 90 2155 100
rect 2200 50 2215 100
rect 2240 120 2280 130
rect 2240 100 2250 120
rect 2270 115 2280 120
rect 2325 115 2340 160
rect 2270 100 2340 115
rect 2240 90 2280 100
rect 2325 50 2340 100
rect 2365 120 2405 130
rect 2365 100 2375 120
rect 2395 115 2405 120
rect 2450 115 2465 160
rect 2515 130 2530 340
rect 2395 100 2465 115
rect 2365 90 2405 100
rect 2450 50 2465 100
rect 2490 120 2530 130
rect 2490 100 2500 120
rect 2520 100 2530 120
rect 2490 90 2530 100
rect 0 -15 15 0
rect 55 -15 70 0
rect 260 -40 275 0
rect 315 -15 330 0
rect 440 -40 455 0
rect 495 -15 510 0
rect 700 -15 715 0
rect 755 -15 770 0
rect 260 -55 455 -40
rect 880 -80 895 0
rect 935 -15 950 0
rect 1140 -40 1155 0
rect 1195 -15 1210 0
rect 1330 -40 1345 0
rect 1385 -15 1400 0
rect 1590 -15 1605 0
rect 1645 -15 1660 0
rect 1770 -15 1785 0
rect 1825 -15 1840 0
rect 1950 -15 1965 0
rect 2075 -15 2090 0
rect 2200 -15 2215 0
rect 2325 -15 2340 0
rect 2450 -15 2465 0
rect 1140 -55 1345 -40
rect 1825 -25 1865 -15
rect 1825 -45 1835 -25
rect 1855 -45 1865 -25
rect 1825 -55 1865 -45
rect -60 -95 895 -80
<< polycont >>
rect 195 285 215 305
rect 1755 285 1775 305
rect 135 225 155 245
rect 75 75 95 95
rect 575 225 595 245
rect 335 115 355 135
rect 515 75 535 95
rect 1015 225 1035 245
rect 955 75 975 95
rect 1465 225 1485 245
rect 1215 115 1235 135
rect 1405 75 1425 95
rect 1875 100 1895 120
rect 2000 100 2020 120
rect 2125 100 2145 120
rect 2250 100 2270 120
rect 2375 100 2395 120
rect 2500 100 2520 120
rect 1835 -45 1855 -25
<< locali >>
rect 185 305 225 315
rect 185 285 195 305
rect 215 295 225 305
rect 1745 305 1785 315
rect 1745 295 1755 305
rect 215 285 1755 295
rect 1775 295 1785 305
rect 1775 285 2530 295
rect 185 275 2530 285
rect 185 255 205 275
rect -35 245 -5 255
rect -35 175 -30 245
rect -10 175 -5 245
rect -35 165 -5 175
rect 20 245 50 255
rect 20 175 25 245
rect 45 175 50 245
rect 20 165 50 175
rect 75 245 165 255
rect 75 175 80 245
rect 100 230 135 245
rect 100 175 105 230
rect 125 225 135 230
rect 155 225 165 245
rect 125 215 165 225
rect 185 245 255 255
rect 185 235 230 245
rect 75 165 105 175
rect 80 145 100 165
rect 20 125 100 145
rect 20 45 40 125
rect 185 105 205 235
rect 225 175 230 235
rect 250 175 255 245
rect 225 165 255 175
rect 280 245 310 255
rect 280 175 285 245
rect 305 175 310 245
rect 280 165 310 175
rect 335 245 365 255
rect 335 175 340 245
rect 360 175 365 245
rect 335 165 365 175
rect 405 245 435 255
rect 405 175 410 245
rect 430 175 435 245
rect 405 165 435 175
rect 460 245 490 255
rect 460 175 465 245
rect 485 175 490 245
rect 460 165 490 175
rect 515 245 605 255
rect 515 175 520 245
rect 540 230 575 245
rect 540 175 545 230
rect 565 225 575 230
rect 595 225 605 245
rect 565 215 605 225
rect 625 245 695 255
rect 625 235 670 245
rect 515 165 545 175
rect 230 145 250 165
rect 520 145 540 165
rect 230 125 305 145
rect 65 95 205 105
rect 65 75 75 95
rect 95 85 205 95
rect 95 75 105 85
rect 65 65 105 75
rect 285 45 305 125
rect 325 135 540 145
rect 325 115 335 135
rect 355 125 540 135
rect 355 115 365 125
rect 325 105 365 115
rect 460 45 480 125
rect 625 105 645 235
rect 665 175 670 235
rect 690 175 695 245
rect 665 165 695 175
rect 720 245 750 255
rect 720 175 725 245
rect 745 175 750 245
rect 720 165 750 175
rect 775 245 805 255
rect 775 175 780 245
rect 800 175 805 245
rect 775 165 805 175
rect 845 245 875 255
rect 845 175 850 245
rect 870 175 875 245
rect 845 165 875 175
rect 900 245 930 255
rect 900 175 905 245
rect 925 175 930 245
rect 900 165 930 175
rect 955 245 1045 255
rect 955 175 960 245
rect 980 230 1015 245
rect 980 175 985 230
rect 1005 225 1015 230
rect 1035 225 1045 245
rect 1005 215 1045 225
rect 1065 245 1135 255
rect 1065 235 1110 245
rect 955 165 985 175
rect 670 145 690 165
rect 960 145 980 165
rect 670 125 745 145
rect 505 95 645 105
rect 505 75 515 95
rect 535 85 645 95
rect 535 75 545 85
rect 505 65 545 75
rect 725 45 745 125
rect 900 125 980 145
rect 900 45 920 125
rect 1065 105 1085 235
rect 1105 175 1110 235
rect 1130 175 1135 245
rect 1105 165 1135 175
rect 1160 245 1190 255
rect 1160 175 1165 245
rect 1185 175 1190 245
rect 1160 165 1190 175
rect 1215 245 1325 255
rect 1215 175 1220 245
rect 1240 175 1260 245
rect 1280 175 1300 245
rect 1320 175 1325 245
rect 1215 165 1325 175
rect 1350 245 1380 255
rect 1350 175 1355 245
rect 1375 175 1380 245
rect 1350 165 1380 175
rect 1405 245 1495 255
rect 1405 175 1410 245
rect 1430 230 1465 245
rect 1430 175 1435 230
rect 1455 225 1465 230
rect 1485 225 1495 245
rect 1455 215 1495 225
rect 1515 245 1585 255
rect 1515 235 1560 245
rect 1405 165 1435 175
rect 1110 145 1130 165
rect 1410 145 1430 165
rect 1110 125 1185 145
rect 945 95 1085 105
rect 945 75 955 95
rect 975 85 1085 95
rect 975 75 985 85
rect 945 65 985 75
rect 1165 45 1185 125
rect 1205 135 1430 145
rect 1205 115 1215 135
rect 1235 125 1430 135
rect 1235 115 1245 125
rect 1205 105 1245 115
rect 1350 45 1370 125
rect 1515 105 1535 235
rect 1555 175 1560 235
rect 1580 175 1585 245
rect 1555 165 1585 175
rect 1610 245 1640 255
rect 1610 175 1615 245
rect 1635 175 1640 245
rect 1610 165 1640 175
rect 1665 245 1695 255
rect 1665 175 1670 245
rect 1690 175 1695 245
rect 1665 165 1695 175
rect 1735 245 1765 255
rect 1735 175 1740 245
rect 1760 175 1765 245
rect 1735 165 1765 175
rect 1790 245 1820 255
rect 1790 175 1795 245
rect 1815 175 1820 245
rect 1790 165 1820 175
rect 1845 245 1875 255
rect 1845 175 1850 245
rect 1870 175 1875 245
rect 1845 165 1875 175
rect 1915 245 1945 255
rect 1915 175 1920 245
rect 1940 175 1945 245
rect 1915 165 1945 175
rect 1970 245 2000 255
rect 1970 175 1975 245
rect 1995 175 2000 245
rect 1970 165 2000 175
rect 2040 245 2070 255
rect 2040 175 2045 245
rect 2065 175 2070 245
rect 2040 165 2070 175
rect 2095 245 2125 255
rect 2095 175 2100 245
rect 2120 175 2125 245
rect 2095 165 2125 175
rect 2165 245 2195 255
rect 2165 175 2170 245
rect 2190 175 2195 245
rect 2165 165 2195 175
rect 2220 245 2250 255
rect 2220 175 2225 245
rect 2245 175 2250 245
rect 2220 165 2250 175
rect 2290 245 2320 255
rect 2290 175 2295 245
rect 2315 175 2320 245
rect 2290 165 2320 175
rect 2345 245 2375 255
rect 2345 175 2350 245
rect 2370 175 2375 245
rect 2345 165 2375 175
rect 2415 245 2445 255
rect 2415 175 2420 245
rect 2440 175 2445 245
rect 2415 165 2445 175
rect 2470 245 2500 255
rect 2470 175 2475 245
rect 2495 175 2500 245
rect 2470 165 2500 175
rect 1560 145 1580 165
rect 1740 145 1760 165
rect 1850 145 1870 165
rect 1560 125 1635 145
rect 1740 130 1870 145
rect 1980 130 2000 165
rect 2105 130 2125 165
rect 2230 130 2250 165
rect 2355 130 2375 165
rect 2480 130 2500 165
rect 1740 125 1905 130
rect 1395 95 1535 105
rect 1395 75 1405 95
rect 1425 85 1535 95
rect 1425 75 1435 85
rect 1395 65 1435 75
rect 1615 45 1635 125
rect 1850 120 1905 125
rect 1850 100 1875 120
rect 1895 100 1905 120
rect 1850 90 1905 100
rect 1980 120 2030 130
rect 1980 100 2000 120
rect 2020 100 2030 120
rect 1980 90 2030 100
rect 2105 120 2155 130
rect 2105 100 2125 120
rect 2145 100 2155 120
rect 2105 90 2155 100
rect 2230 120 2280 130
rect 2230 100 2250 120
rect 2270 100 2280 120
rect 2230 90 2280 100
rect 2355 120 2405 130
rect 2355 100 2375 120
rect 2395 100 2405 120
rect 2355 90 2405 100
rect 2480 120 2530 130
rect 2480 100 2500 120
rect 2520 100 2530 120
rect 2480 90 2530 100
rect 1850 45 1870 90
rect 1980 45 2000 90
rect 2105 45 2125 90
rect 2230 45 2250 90
rect 2355 45 2375 90
rect 2480 45 2500 90
rect -35 35 -5 45
rect -35 15 -30 35
rect -10 15 -5 35
rect -35 5 -5 15
rect 20 35 50 45
rect 20 15 25 35
rect 45 15 50 35
rect 20 5 50 15
rect 75 35 105 45
rect 75 15 80 35
rect 100 15 105 35
rect 75 5 105 15
rect 225 35 255 45
rect 225 15 230 35
rect 250 15 255 35
rect 225 5 255 15
rect 280 35 310 45
rect 280 15 285 35
rect 305 15 310 35
rect 280 5 310 15
rect 335 35 365 45
rect 335 15 340 35
rect 360 15 365 35
rect 335 5 365 15
rect 405 35 435 45
rect 405 15 410 35
rect 430 15 435 35
rect 405 5 435 15
rect 460 35 490 45
rect 460 15 465 35
rect 485 15 490 35
rect 460 5 490 15
rect 515 35 545 45
rect 515 15 520 35
rect 540 15 545 35
rect 515 5 545 15
rect 665 35 695 45
rect 665 15 670 35
rect 690 15 695 35
rect 665 5 695 15
rect 720 35 750 45
rect 720 15 725 35
rect 745 15 750 35
rect 720 5 750 15
rect 775 35 805 45
rect 775 15 780 35
rect 800 15 805 35
rect 775 5 805 15
rect 845 35 875 45
rect 845 15 850 35
rect 870 15 875 35
rect 845 5 875 15
rect 900 35 930 45
rect 900 15 905 35
rect 925 15 930 35
rect 900 5 930 15
rect 955 35 985 45
rect 955 15 960 35
rect 980 15 985 35
rect 955 5 985 15
rect 1105 35 1135 45
rect 1105 15 1110 35
rect 1130 15 1135 35
rect 1105 5 1135 15
rect 1160 35 1190 45
rect 1160 15 1165 35
rect 1185 15 1190 35
rect 1160 5 1190 15
rect 1215 35 1325 45
rect 1215 15 1220 35
rect 1240 15 1260 35
rect 1280 15 1300 35
rect 1320 15 1325 35
rect 1215 5 1325 15
rect 1350 35 1380 45
rect 1350 15 1355 35
rect 1375 15 1380 35
rect 1350 5 1380 15
rect 1405 35 1435 45
rect 1405 15 1410 35
rect 1430 15 1435 35
rect 1405 5 1435 15
rect 1555 35 1585 45
rect 1555 15 1560 35
rect 1580 15 1585 35
rect 1555 5 1585 15
rect 1610 35 1640 45
rect 1610 15 1615 35
rect 1635 15 1640 35
rect 1610 5 1640 15
rect 1665 35 1695 45
rect 1665 15 1670 35
rect 1690 15 1695 35
rect 1665 5 1695 15
rect 1735 35 1765 45
rect 1735 15 1740 35
rect 1760 15 1765 35
rect 1735 5 1765 15
rect 1790 35 1820 45
rect 1790 15 1795 35
rect 1815 15 1820 35
rect 1790 5 1820 15
rect 1845 35 1875 45
rect 1845 15 1850 35
rect 1870 15 1875 35
rect 1845 5 1875 15
rect 1915 35 1945 45
rect 1915 15 1920 35
rect 1940 15 1945 35
rect 1915 5 1945 15
rect 1970 35 2000 45
rect 1970 15 1975 35
rect 1995 15 2000 35
rect 1970 5 2000 15
rect 2040 35 2070 45
rect 2040 15 2045 35
rect 2065 15 2070 35
rect 2040 5 2070 15
rect 2095 35 2125 45
rect 2095 15 2100 35
rect 2120 15 2125 35
rect 2095 5 2125 15
rect 2165 35 2195 45
rect 2165 15 2170 35
rect 2190 15 2195 35
rect 2165 5 2195 15
rect 2220 35 2250 45
rect 2220 15 2225 35
rect 2245 15 2250 35
rect 2220 5 2250 15
rect 2290 35 2320 45
rect 2290 15 2295 35
rect 2315 15 2320 35
rect 2290 5 2320 15
rect 2345 35 2375 45
rect 2345 15 2350 35
rect 2370 15 2375 35
rect 2345 5 2375 15
rect 2415 35 2445 45
rect 2415 15 2420 35
rect 2440 15 2445 35
rect 2415 5 2445 15
rect 2470 35 2500 45
rect 2470 15 2475 35
rect 2495 15 2500 35
rect 2470 5 2500 15
rect 1165 -15 1185 5
rect 1165 -25 2530 -15
rect 1165 -35 1835 -25
rect 1825 -45 1835 -35
rect 1855 -35 2530 -25
rect 1855 -45 1865 -35
rect 1825 -55 1865 -45
<< viali >>
rect -30 175 -10 245
rect 340 175 360 245
rect 410 175 430 245
rect 780 175 800 245
rect 850 175 870 245
rect 1220 175 1240 245
rect 1260 175 1280 245
rect 1300 175 1320 245
rect 1670 175 1690 245
rect 1795 175 1815 245
rect 1920 175 1940 245
rect 2045 175 2065 245
rect 2170 175 2190 245
rect 2295 175 2315 245
rect 2420 175 2440 245
rect -30 15 -10 35
rect 80 15 100 35
rect 230 15 250 35
rect 340 15 360 35
rect 410 15 430 35
rect 520 15 540 35
rect 670 15 690 35
rect 780 15 800 35
rect 850 15 870 35
rect 960 15 980 35
rect 1110 15 1130 35
rect 1220 15 1240 35
rect 1260 15 1280 35
rect 1300 15 1320 35
rect 1410 15 1430 35
rect 1560 15 1580 35
rect 1670 15 1690 35
rect 1740 15 1760 35
rect 1920 15 1940 35
rect 2045 15 2065 35
rect 2170 15 2190 35
rect 2295 15 2315 35
rect 2420 15 2440 35
<< metal1 >>
rect -40 245 2505 260
rect -40 175 -30 245
rect -10 175 340 245
rect 360 175 410 245
rect 430 175 780 245
rect 800 175 850 245
rect 870 175 1220 245
rect 1240 175 1260 245
rect 1280 175 1300 245
rect 1320 175 1670 245
rect 1690 175 1795 245
rect 1815 175 1920 245
rect 1940 175 2045 245
rect 2065 175 2170 245
rect 2190 175 2295 245
rect 2315 175 2420 245
rect 2440 175 2505 245
rect -40 160 2505 175
rect -40 35 2505 50
rect -40 15 -30 35
rect -10 15 80 35
rect 100 15 230 35
rect 250 15 340 35
rect 360 15 410 35
rect 430 15 520 35
rect 540 15 670 35
rect 690 15 780 35
rect 800 15 850 35
rect 870 15 960 35
rect 980 15 1110 35
rect 1130 15 1220 35
rect 1240 15 1260 35
rect 1280 15 1300 35
rect 1320 15 1410 35
rect 1430 15 1560 35
rect 1580 15 1670 35
rect 1690 15 1740 35
rect 1760 15 1920 35
rect 1940 15 2045 35
rect 2065 15 2170 35
rect 2190 15 2295 35
rect 2315 15 2420 35
rect 2440 15 2505 35
rect -40 0 2505 15
<< labels >>
flabel poly -60 95 -60 95 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel poly 150 125 150 125 7 FreeSans 160 0 -80 0 QA_b
flabel locali 540 125 540 125 3 FreeSans 160 0 80 0 E
flabel locali 745 125 745 125 3 FreeSans 160 0 80 0 E_b
flabel poly 770 325 770 325 3 FreeSans 160 0 80 0 Reset
flabel locali 1905 130 1905 130 3 FreeSans 160 0 80 0 before_Reset
flabel poly -60 -85 -60 -85 7 FreeSans 160 0 -80 0 F_VCO
port 2 w
flabel poly 1030 135 1030 135 7 FreeSans 160 0 -80 0 QB_b
flabel locali 1430 125 1430 125 3 FreeSans 160 0 80 0 F
flabel locali 1635 110 1635 110 3 FreeSans 160 0 80 0 F_b
flabel metal1 -40 25 -40 25 7 FreeSans 160 0 -80 0 GNDA
port 6 w
flabel metal1 -40 210 -40 210 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel locali 2530 285 2530 285 3 FreeSans 160 0 80 0 QA
port 4 e
flabel locali 2530 -25 2530 -25 3 FreeSans 160 0 80 0 QB
port 5 e
<< end >>
