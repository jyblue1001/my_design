magic
tech sky130A
timestamp 1723040855
<< nwell >>
rect -270 630 -65 985
<< nmos >>
rect -200 425 -185 525
<< pmos >>
rect -200 650 -185 750
<< ndiff >>
rect -250 510 -200 525
rect -250 440 -235 510
rect -215 440 -200 510
rect -250 425 -200 440
rect -185 510 -135 525
rect -185 440 -170 510
rect -150 440 -135 510
rect -185 425 -135 440
<< pdiff >>
rect -250 735 -200 750
rect -250 665 -235 735
rect -215 665 -200 735
rect -250 650 -200 665
rect -185 735 -135 750
rect -185 665 -170 735
rect -150 665 -135 735
rect -185 650 -135 665
<< ndiffc >>
rect -235 440 -215 510
rect -170 440 -150 510
<< pdiffc >>
rect -235 665 -215 735
rect -170 665 -150 735
<< psubdiff >>
rect -135 510 -85 525
rect -135 440 -120 510
rect -100 440 -85 510
rect -135 425 -85 440
<< nsubdiff >>
rect -135 735 -85 750
rect -135 665 -120 735
rect -100 665 -85 735
rect -135 650 -85 665
<< psubdiffcont >>
rect -120 440 -100 510
<< nsubdiffcont >>
rect -120 665 -100 735
<< poly >>
rect -130 845 -65 855
rect -130 825 -120 845
rect -100 840 -65 845
rect -100 825 -90 840
rect -130 815 -90 825
rect -200 750 -185 765
rect -200 605 -185 650
rect -200 595 -160 605
rect -200 575 -190 595
rect -170 575 -160 595
rect -200 565 -160 575
rect -200 525 -185 565
rect -200 410 -185 425
rect -130 350 -90 360
rect -130 330 -120 350
rect -100 335 -90 350
rect -100 330 -65 335
rect -130 320 -65 330
<< polycont >>
rect -120 825 -100 845
rect -190 575 -170 595
rect -120 330 -100 350
<< locali >>
rect -130 845 -90 855
rect -130 835 -120 845
rect -225 825 -120 835
rect -100 825 -90 845
rect -225 815 -90 825
rect -225 745 -205 815
rect -245 735 -205 745
rect -245 665 -235 735
rect -215 665 -205 735
rect -245 655 -205 665
rect -180 735 -90 745
rect -180 665 -170 735
rect -150 665 -120 735
rect -100 665 -90 735
rect -180 655 -90 665
rect -245 520 -225 655
rect -200 595 -160 605
rect -200 575 -190 595
rect -170 585 -160 595
rect -170 575 -65 585
rect -200 565 -65 575
rect -245 510 -205 520
rect -245 440 -235 510
rect -215 440 -205 510
rect -245 430 -205 440
rect -180 510 -90 520
rect -180 440 -170 510
rect -150 440 -120 510
rect -100 440 -90 510
rect -180 430 -90 440
rect -225 360 -205 430
rect -225 350 -90 360
rect -225 340 -120 350
rect -130 330 -120 340
rect -100 330 -90 350
rect -130 320 -90 330
<< viali >>
rect -170 665 -150 735
rect -120 665 -100 735
rect -190 575 -170 595
rect -170 440 -150 510
rect -120 440 -100 510
<< metal1 >>
rect -270 735 -65 965
rect -270 665 -170 735
rect -150 665 -120 735
rect -100 665 -65 735
rect -270 650 -65 665
rect -260 595 -160 605
rect -260 575 -190 595
rect -170 575 -160 595
rect -260 565 -160 575
rect -260 510 -65 525
rect -260 440 -170 510
rect -150 440 -120 510
rect -100 440 -65 510
rect -260 210 -65 440
<< end >>
