* PEX produced on Sat Feb  1 02:34:58 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from TSPC_FF_ratioed_divide5_magic.ext - technology: sky130A

.subckt TSPC_FF_ratioed_divide5_magic VOUT VIN VDDA GNDA
X0 M.t3 Q2_b.t2 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1 E.t0 VIN.t0 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X2 D.t2 VIN.t1 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 I.t0 VOUT.t2 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 Q2_b.t1 VIN.t2 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X5 F.t1 E.t2 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X6 GNDA.t31 VIN.t3 J.t2 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 A.t2 Q2_b.t3 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 B.t1 VIN.t4 C.t1 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 I.t1 Q2_b.t4 H.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X10 A.t0 Q2_b.t5 GNDA.t24 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X11 GNDA.t16 VIN.t5 D.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X12 VDDA.t12 A.t3 B.t0 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X13 K.t1 Q2_b.t6 L.t1 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X14 GNDA.t29 VIN.t6 J.t1 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 GNDA.t21 Q2_b.t7 M.t2 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X16 VDDA.t1 VOUT.t3 K.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 GNDA.t19 Q2_b.t8 M.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 G.t1 VOUT.t4 F.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X19 GNDA.t14 VIN.t7 D.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X20 GNDA.t33 E.t3 I.t2 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X21 J.t0 VIN.t8 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X22 E.t1 D.t4 GNDA.t35 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 VDDA.t10 G.t3 J.t3 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X24 D.t3 B.t2 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X25 VDDA.t20 Q2_b.t9 G.t2 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X26 VDDA.t18 Q2_b.t10 A.t1 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 C.t0 A.t4 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X28 H.t0 VIN.t9 G.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X29 Q2_b.t0 J.t4 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X30 VOUT.t1 M.t4 GNDA.t6 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X31 M.t0 K.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X32 VOUT.t0 Q2_b.t11 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X33 L.t0 VOUT.t5 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
R0 Q2_b.n6 Q2_b.t5 2779.53
R1 Q2_b.n7 Q2_b.n6 1206
R2 Q2_b.n4 Q2_b.t1 777.4
R3 Q2_b.t4 Q2_b.t9 514.134
R4 Q2_b.n3 Q2_b.n2 364.178
R5 Q2_b.n0 Q2_b.t11 353.467
R6 Q2_b.t5 Q2_b.n5 353.467
R7 Q2_b.n5 Q2_b.t3 289.2
R8 Q2_b.n4 Q2_b.n3 257.079
R9 Q2_b.t0 Q2_b.n7 233
R10 Q2_b.n6 Q2_b.t4 208.868
R11 Q2_b.n0 Q2_b.t7 192.8
R12 Q2_b.n2 Q2_b.n1 176.733
R13 Q2_b.n2 Q2_b.t8 112.468
R14 Q2_b.n1 Q2_b.t2 112.468
R15 Q2_b.n3 Q2_b.t6 112.468
R16 Q2_b.n5 Q2_b.t10 112.468
R17 Q2_b.n1 Q2_b.n0 96.4005
R18 Q2_b.n7 Q2_b.n4 21.3338
R19 GNDA.t34 GNDA.t2 3500
R20 GNDA.t3 GNDA.t7 3400
R21 GNDA.t0 GNDA.t30 3300
R22 GNDA.n16 GNDA.t23 3150
R23 GNDA.t22 GNDA.t18 2500
R24 GNDA.t17 GNDA.t13 2500
R25 GNDA.n16 GNDA.t9 1350
R26 GNDA.n17 GNDA.n16 1170
R27 GNDA.t20 GNDA.t5 1100
R28 GNDA.t26 GNDA.t20 1100
R29 GNDA.t18 GNDA.t26 1100
R30 GNDA.t7 GNDA.t22 1100
R31 GNDA.t28 GNDA.t3 1100
R32 GNDA.t11 GNDA.t28 1100
R33 GNDA.t30 GNDA.t11 1100
R34 GNDA.t32 GNDA.t0 1100
R35 GNDA.t25 GNDA.t32 1100
R36 GNDA.t2 GNDA.t25 1100
R37 GNDA.t15 GNDA.t34 1100
R38 GNDA.t36 GNDA.t15 1100
R39 GNDA.t13 GNDA.t36 1100
R40 GNDA.t9 GNDA.t17 1100
R41 GNDA.n19 GNDA.t24 242.3
R42 GNDA.n3 GNDA.t8 242.3
R43 GNDA.n15 GNDA.t10 233
R44 GNDA.n2 GNDA.n0 194.576
R45 GNDA.n13 GNDA.n12 194.3
R46 GNDA.n11 GNDA.n10 194.3
R47 GNDA.n9 GNDA.n8 194.3
R48 GNDA.n7 GNDA.n6 194.3
R49 GNDA.n5 GNDA.n4 194.3
R50 GNDA.n2 GNDA.n1 194.3
R51 GNDA.n12 GNDA.t37 48.0005
R52 GNDA.n12 GNDA.t14 48.0005
R53 GNDA.n10 GNDA.t35 48.0005
R54 GNDA.n10 GNDA.t16 48.0005
R55 GNDA.n8 GNDA.t1 48.0005
R56 GNDA.n8 GNDA.t33 48.0005
R57 GNDA.n6 GNDA.t12 48.0005
R58 GNDA.n6 GNDA.t31 48.0005
R59 GNDA.n4 GNDA.t4 48.0005
R60 GNDA.n4 GNDA.t29 48.0005
R61 GNDA.n1 GNDA.t27 48.0005
R62 GNDA.n1 GNDA.t19 48.0005
R63 GNDA.n0 GNDA.t6 48.0005
R64 GNDA.n0 GNDA.t21 48.0005
R65 GNDA.n17 GNDA.n15 12.8005
R66 GNDA.n15 GNDA.n14 9.3005
R67 GNDA.n18 GNDA.n17 9.3005
R68 GNDA.n11 GNDA.n9 0.8505
R69 GNDA.n3 GNDA.n2 0.588
R70 GNDA.n14 GNDA.n13 0.588
R71 GNDA.n9 GNDA.n7 0.5505
R72 GNDA.n19 GNDA.n18 0.463
R73 GNDA.n5 GNDA.n3 0.4255
R74 GNDA.n7 GNDA.n5 0.2755
R75 GNDA.n13 GNDA.n11 0.2755
R76 GNDA.n18 GNDA.n14 0.1005
R77 GNDA GNDA.n19 0.1005
R78 M.n0 M.t0 761.4
R79 M.n1 M.t4 349.433
R80 M.n0 M.t1 254.333
R81 M.n2 M.n1 206.333
R82 M.n1 M.n0 70.4005
R83 M.n2 M.t2 48.0005
R84 M.t3 M.n2 48.0005
R85 VIN.n3 VIN.n2 919.244
R86 VIN VIN.n7 893.102
R87 VIN.n2 VIN.n1 758.606
R88 VIN.n7 VIN.n6 364.178
R89 VIN.n0 VIN.t2 337.401
R90 VIN.n0 VIN.t6 305.267
R91 VIN.n4 VIN.t5 192.8
R92 VIN.n1 VIN.n0 176.733
R93 VIN.n6 VIN.n5 176.733
R94 VIN.n4 VIN.n3 160.667
R95 VIN.n3 VIN.t0 144.601
R96 VIN.n2 VIN.t9 131.976
R97 VIN.n0 VIN.t8 128.534
R98 VIN.n1 VIN.t3 128.534
R99 VIN.n6 VIN.t7 112.468
R100 VIN.n5 VIN.t1 112.468
R101 VIN.n7 VIN.t4 112.468
R102 VIN.n5 VIN.n4 96.4005
R103 VDDA.t7 VDDA.t19 2804.76
R104 VDDA.t5 VDDA.t0 2533.33
R105 VDDA.t11 VDDA.t21 1538.1
R106 VDDA.t4 VDDA.t9 1492.86
R107 VDDA.t2 VDDA.n9 1289.29
R108 VDDA.n10 VDDA.t23 1289.29
R109 VDDA.n8 VDDA.t16 667.62
R110 VDDA.n1 VDDA.t8 663.801
R111 VDDA.n9 VDDA.t15 610.715
R112 VDDA.n10 VDDA.t7 610.715
R113 VDDA.n16 VDDA.n15 594.301
R114 VDDA.n14 VDDA.n13 594.301
R115 VDDA.n3 VDDA.n2 594.301
R116 VDDA.n5 VDDA.n4 594.301
R117 VDDA.n7 VDDA.n6 594.301
R118 VDDA.t0 VDDA.t2 497.62
R119 VDDA.t9 VDDA.t5 497.62
R120 VDDA.t13 VDDA.t4 497.62
R121 VDDA.t19 VDDA.t13 497.62
R122 VDDA.t23 VDDA.t11 497.62
R123 VDDA.t21 VDDA.t17 497.62
R124 VDDA.n9 VDDA.n8 373.781
R125 VDDA.n11 VDDA.n10 370
R126 VDDA.n15 VDDA.t22 78.8005
R127 VDDA.n15 VDDA.t18 78.8005
R128 VDDA.n13 VDDA.t24 78.8005
R129 VDDA.n13 VDDA.t12 78.8005
R130 VDDA.n2 VDDA.t14 78.8005
R131 VDDA.n2 VDDA.t20 78.8005
R132 VDDA.n4 VDDA.t6 78.8005
R133 VDDA.n4 VDDA.t10 78.8005
R134 VDDA.n6 VDDA.t3 78.8005
R135 VDDA.n6 VDDA.t1 78.8005
R136 VDDA.n11 VDDA.n1 12.8005
R137 VDDA.n1 VDDA.n0 9.3005
R138 VDDA.n12 VDDA.n11 9.3005
R139 VDDA.n8 VDDA.n7 3.20124
R140 VDDA.n3 VDDA.n0 0.913
R141 VDDA.n7 VDDA.n5 0.838
R142 VDDA.n5 VDDA.n3 0.688
R143 VDDA.n16 VDDA.n14 0.563
R144 VDDA.n14 VDDA.n12 0.4255
R145 VDDA VDDA.n16 0.238
R146 VDDA.n12 VDDA.n0 0.1005
R147 E.n0 E.t2 1207.57
R148 E.n0 E.t0 723
R149 E.t2 E.t3 514.134
R150 E.t1 E.n0 314.921
R151 D.n0 D.t3 761.4
R152 D.n1 D.t4 350.349
R153 D.n0 D.t0 254.333
R154 D.n2 D.n1 206.333
R155 D.n1 D.n0 70.4005
R156 D.n2 D.t1 48.0005
R157 D.t2 D.n2 48.0005
R158 VOUT.n2 VOUT.n1 2120.39
R159 VOUT.n1 VOUT.t4 1992.27
R160 VOUT.n3 VOUT.t0 751.801
R161 VOUT.t4 VOUT.t2 514.134
R162 VOUT.n0 VOUT.t5 289.2
R163 VOUT.n2 VOUT.t1 233
R164 VOUT.n1 VOUT.n0 208.868
R165 VOUT.n0 VOUT.t3 176.733
R166 VOUT.n3 VOUT.n2 40.3205
R167 VOUT VOUT.n3 32.0005
R168 I.t0 I.n0 531.067
R169 I.n0 I.t2 48.0005
R170 I.n0 I.t1 48.0005
R171 F.t0 F.t1 157.601
R172 J.n2 J.t3 723.534
R173 J.n1 J.t4 553.534
R174 J.t2 J.n2 254.333
R175 J.n1 J.n0 206.333
R176 J.n2 J.n1 70.4005
R177 J.n0 J.t1 48.0005
R178 J.n0 J.t0 48.0005
R179 A.n2 A.t1 755.534
R180 A.t2 A.n2 685.134
R181 A.n1 A.n0 389.733
R182 A.n1 A.t0 340.2
R183 A.n0 A.t4 321.334
R184 A.n0 A.t3 144.601
R185 A.n2 A.n1 19.2005
R186 C.t0 C.t1 96.0005
R187 B.n0 B.t0 663.801
R188 B.n0 B.t2 380.368
R189 B B.t1 282.921
R190 B B.n0 114.133
R191 H.t0 H.t1 96.0005
R192 L.t0 L.t1 96.0005
R193 K.n0 K.t0 663.801
R194 K.t1 K.n0 397.053
R195 K.n0 K.t2 380.368
R196 G.n0 G.t1 685.134
R197 G.n1 G.t2 685.134
R198 G.n0 G.t3 534.268
R199 G.t0 G.n1 340.521
R200 G.n1 G.n0 105.6
C0 VIN B 0.143413f
C1 VDDA VIN 0.290147f
C2 VOUT VDDA 0.659192f
C3 VOUT VIN 0.065488f
C4 VDDA B 0.305296f
C5 VOUT GNDA 1.86297f
C6 VIN GNDA 1.85246f
C7 VDDA GNDA 3.92947f
C8 B GNDA 0.256727f
.ends

