magic
tech sky130A
timestamp 1739198281
<< nwell >>
rect -190 -3460 2265 -2840
<< nmos >>
rect -90 -2750 -75 -2650
rect -35 -2750 -20 -2650
rect 170 -2750 185 -2650
rect 225 -2750 240 -2650
rect 360 -2750 375 -2650
rect 415 -2750 430 -2650
rect 620 -2750 635 -2650
rect 675 -2750 690 -2650
rect 840 -2750 855 -2650
rect 895 -2750 910 -2650
rect 1060 -2750 1075 -2650
rect 1225 -2750 1240 -2650
rect 1450 -2750 1465 -2650
rect 1645 -2750 1660 -2650
rect 1840 -2750 1855 -2650
rect 1985 -2750 2000 -2650
rect -90 -3650 -75 -3550
rect -35 -3650 -20 -3550
rect 170 -3650 185 -3550
rect 225 -3650 240 -3550
rect 360 -3650 375 -3550
rect 415 -3650 430 -3550
rect 620 -3650 635 -3550
rect 675 -3650 690 -3550
rect 875 -3650 890 -3550
rect 1040 -3650 1055 -3550
rect 1205 -3650 1220 -3550
rect 1450 -3650 1465 -3550
rect 1645 -3650 1660 -3550
rect 1840 -3650 1855 -3550
rect 1985 -3650 2000 -3550
rect 2180 -3650 2195 -3550
<< pmos >>
rect -90 -3060 -75 -2860
rect -35 -3060 -20 -2860
rect 170 -3060 185 -2860
rect 225 -3060 240 -2860
rect 360 -3060 375 -2860
rect 415 -3060 430 -2860
rect 620 -3060 635 -2860
rect 675 -3060 690 -2860
rect 840 -3060 855 -2860
rect 895 -3060 910 -2860
rect 1060 -3060 1075 -2860
rect 1225 -3060 1240 -2860
rect 1450 -3060 1465 -2860
rect 1645 -3060 1660 -2860
rect 1840 -3060 1855 -2860
rect 1985 -3060 2000 -2860
rect 2180 -3060 2195 -2860
rect -90 -3440 -75 -3240
rect -35 -3440 -20 -3240
rect 170 -3440 185 -3240
rect 225 -3440 240 -3240
rect 360 -3440 375 -3240
rect 415 -3440 430 -3240
rect 620 -3440 635 -3240
rect 675 -3440 690 -3240
rect 875 -3440 890 -3240
rect 1040 -3440 1055 -3240
rect 1205 -3440 1220 -3240
rect 1450 -3440 1465 -3240
rect 1645 -3440 1660 -3240
rect 1840 -3440 1855 -3240
rect 1985 -3440 2000 -3240
<< ndiff >>
rect -130 -2665 -90 -2650
rect -130 -2685 -120 -2665
rect -100 -2685 -90 -2665
rect -130 -2715 -90 -2685
rect -130 -2735 -120 -2715
rect -100 -2735 -90 -2715
rect -130 -2750 -90 -2735
rect -75 -2665 -35 -2650
rect -75 -2685 -65 -2665
rect -45 -2685 -35 -2665
rect -75 -2715 -35 -2685
rect -75 -2735 -65 -2715
rect -45 -2735 -35 -2715
rect -75 -2750 -35 -2735
rect -20 -2665 20 -2650
rect -20 -2685 -10 -2665
rect 10 -2685 20 -2665
rect -20 -2715 20 -2685
rect -20 -2735 -10 -2715
rect 10 -2735 20 -2715
rect -20 -2750 20 -2735
rect 130 -2665 170 -2650
rect 130 -2685 140 -2665
rect 160 -2685 170 -2665
rect 130 -2715 170 -2685
rect 130 -2735 140 -2715
rect 160 -2735 170 -2715
rect 130 -2750 170 -2735
rect 185 -2665 225 -2650
rect 185 -2685 195 -2665
rect 215 -2685 225 -2665
rect 185 -2715 225 -2685
rect 185 -2735 195 -2715
rect 215 -2735 225 -2715
rect 185 -2750 225 -2735
rect 240 -2665 280 -2650
rect 320 -2665 360 -2650
rect 240 -2685 250 -2665
rect 270 -2685 280 -2665
rect 320 -2685 330 -2665
rect 350 -2685 360 -2665
rect 240 -2715 280 -2685
rect 320 -2715 360 -2685
rect 240 -2735 250 -2715
rect 270 -2735 280 -2715
rect 320 -2735 330 -2715
rect 350 -2735 360 -2715
rect 240 -2750 280 -2735
rect 320 -2750 360 -2735
rect 375 -2665 415 -2650
rect 375 -2685 385 -2665
rect 405 -2685 415 -2665
rect 375 -2715 415 -2685
rect 375 -2735 385 -2715
rect 405 -2735 415 -2715
rect 375 -2750 415 -2735
rect 430 -2665 470 -2650
rect 430 -2685 440 -2665
rect 460 -2685 470 -2665
rect 430 -2715 470 -2685
rect 430 -2735 440 -2715
rect 460 -2735 470 -2715
rect 430 -2750 470 -2735
rect 580 -2665 620 -2650
rect 580 -2685 590 -2665
rect 610 -2685 620 -2665
rect 580 -2715 620 -2685
rect 580 -2735 590 -2715
rect 610 -2735 620 -2715
rect 580 -2750 620 -2735
rect 635 -2665 675 -2650
rect 635 -2685 645 -2665
rect 665 -2685 675 -2665
rect 635 -2715 675 -2685
rect 635 -2735 645 -2715
rect 665 -2735 675 -2715
rect 635 -2750 675 -2735
rect 690 -2665 730 -2650
rect 690 -2685 700 -2665
rect 720 -2685 730 -2665
rect 690 -2715 730 -2685
rect 690 -2735 700 -2715
rect 720 -2735 730 -2715
rect 690 -2750 730 -2735
rect 800 -2665 840 -2650
rect 800 -2685 810 -2665
rect 830 -2685 840 -2665
rect 800 -2715 840 -2685
rect 800 -2735 810 -2715
rect 830 -2735 840 -2715
rect 800 -2750 840 -2735
rect 855 -2665 895 -2650
rect 855 -2685 865 -2665
rect 885 -2685 895 -2665
rect 855 -2715 895 -2685
rect 855 -2735 865 -2715
rect 885 -2735 895 -2715
rect 855 -2750 895 -2735
rect 910 -2665 950 -2650
rect 910 -2685 920 -2665
rect 940 -2685 950 -2665
rect 910 -2715 950 -2685
rect 910 -2735 920 -2715
rect 940 -2735 950 -2715
rect 910 -2750 950 -2735
rect 1020 -2665 1060 -2650
rect 1020 -2685 1030 -2665
rect 1050 -2685 1060 -2665
rect 1020 -2715 1060 -2685
rect 1020 -2735 1030 -2715
rect 1050 -2735 1060 -2715
rect 1020 -2750 1060 -2735
rect 1075 -2665 1115 -2650
rect 1075 -2685 1085 -2665
rect 1105 -2685 1115 -2665
rect 1075 -2715 1115 -2685
rect 1075 -2735 1085 -2715
rect 1105 -2735 1115 -2715
rect 1075 -2750 1115 -2735
rect 1185 -2665 1225 -2650
rect 1185 -2685 1195 -2665
rect 1215 -2685 1225 -2665
rect 1185 -2715 1225 -2685
rect 1185 -2735 1195 -2715
rect 1215 -2735 1225 -2715
rect 1185 -2750 1225 -2735
rect 1240 -2665 1280 -2650
rect 1240 -2685 1250 -2665
rect 1270 -2685 1280 -2665
rect 1240 -2715 1280 -2685
rect 1240 -2735 1250 -2715
rect 1270 -2735 1280 -2715
rect 1240 -2750 1280 -2735
rect 1400 -2665 1450 -2650
rect 1400 -2685 1415 -2665
rect 1435 -2685 1450 -2665
rect 1400 -2715 1450 -2685
rect 1400 -2735 1415 -2715
rect 1435 -2735 1450 -2715
rect 1400 -2750 1450 -2735
rect 1465 -2665 1515 -2650
rect 1465 -2685 1480 -2665
rect 1500 -2685 1515 -2665
rect 1465 -2715 1515 -2685
rect 1465 -2735 1480 -2715
rect 1500 -2735 1515 -2715
rect 1465 -2750 1515 -2735
rect 1595 -2665 1645 -2650
rect 1595 -2685 1610 -2665
rect 1630 -2685 1645 -2665
rect 1595 -2715 1645 -2685
rect 1595 -2735 1610 -2715
rect 1630 -2735 1645 -2715
rect 1595 -2750 1645 -2735
rect 1660 -2665 1710 -2650
rect 1660 -2685 1675 -2665
rect 1695 -2685 1710 -2665
rect 1660 -2715 1710 -2685
rect 1660 -2735 1675 -2715
rect 1695 -2735 1710 -2715
rect 1660 -2750 1710 -2735
rect 1790 -2665 1840 -2650
rect 1790 -2685 1805 -2665
rect 1825 -2685 1840 -2665
rect 1790 -2715 1840 -2685
rect 1790 -2735 1805 -2715
rect 1825 -2735 1840 -2715
rect 1790 -2750 1840 -2735
rect 1855 -2665 1905 -2650
rect 1855 -2685 1870 -2665
rect 1890 -2685 1905 -2665
rect 1855 -2715 1905 -2685
rect 1855 -2735 1870 -2715
rect 1890 -2735 1905 -2715
rect 1855 -2750 1905 -2735
rect 1935 -2665 1985 -2650
rect 1935 -2685 1950 -2665
rect 1970 -2685 1985 -2665
rect 1935 -2715 1985 -2685
rect 1935 -2735 1950 -2715
rect 1970 -2735 1985 -2715
rect 1935 -2750 1985 -2735
rect 2000 -2665 2050 -2650
rect 2000 -2685 2015 -2665
rect 2035 -2685 2050 -2665
rect 2000 -2715 2050 -2685
rect 2000 -2735 2015 -2715
rect 2035 -2735 2050 -2715
rect 2000 -2750 2050 -2735
rect -130 -3565 -90 -3550
rect -130 -3585 -120 -3565
rect -100 -3585 -90 -3565
rect -130 -3615 -90 -3585
rect -130 -3635 -120 -3615
rect -100 -3635 -90 -3615
rect -130 -3650 -90 -3635
rect -75 -3565 -35 -3550
rect -75 -3585 -65 -3565
rect -45 -3585 -35 -3565
rect -75 -3615 -35 -3585
rect -75 -3635 -65 -3615
rect -45 -3635 -35 -3615
rect -75 -3650 -35 -3635
rect -20 -3565 20 -3550
rect -20 -3585 -10 -3565
rect 10 -3585 20 -3565
rect -20 -3615 20 -3585
rect -20 -3635 -10 -3615
rect 10 -3635 20 -3615
rect -20 -3650 20 -3635
rect 130 -3565 170 -3550
rect 130 -3585 140 -3565
rect 160 -3585 170 -3565
rect 130 -3615 170 -3585
rect 130 -3635 140 -3615
rect 160 -3635 170 -3615
rect 130 -3650 170 -3635
rect 185 -3565 225 -3550
rect 185 -3585 195 -3565
rect 215 -3585 225 -3565
rect 185 -3615 225 -3585
rect 185 -3635 195 -3615
rect 215 -3635 225 -3615
rect 185 -3650 225 -3635
rect 240 -3565 280 -3550
rect 320 -3565 360 -3550
rect 240 -3585 250 -3565
rect 270 -3585 280 -3565
rect 320 -3585 330 -3565
rect 350 -3585 360 -3565
rect 240 -3615 280 -3585
rect 320 -3615 360 -3585
rect 240 -3635 250 -3615
rect 270 -3635 280 -3615
rect 320 -3635 330 -3615
rect 350 -3635 360 -3615
rect 240 -3650 280 -3635
rect 320 -3650 360 -3635
rect 375 -3565 415 -3550
rect 375 -3585 385 -3565
rect 405 -3585 415 -3565
rect 375 -3615 415 -3585
rect 375 -3635 385 -3615
rect 405 -3635 415 -3615
rect 375 -3650 415 -3635
rect 430 -3565 470 -3550
rect 430 -3585 440 -3565
rect 460 -3585 470 -3565
rect 430 -3615 470 -3585
rect 430 -3635 440 -3615
rect 460 -3635 470 -3615
rect 430 -3650 470 -3635
rect 580 -3565 620 -3550
rect 580 -3585 590 -3565
rect 610 -3585 620 -3565
rect 580 -3615 620 -3585
rect 580 -3635 590 -3615
rect 610 -3635 620 -3615
rect 580 -3650 620 -3635
rect 635 -3565 675 -3550
rect 635 -3585 645 -3565
rect 665 -3585 675 -3565
rect 635 -3615 675 -3585
rect 635 -3635 645 -3615
rect 665 -3635 675 -3615
rect 635 -3650 675 -3635
rect 690 -3565 730 -3550
rect 690 -3585 700 -3565
rect 720 -3585 730 -3565
rect 690 -3615 730 -3585
rect 690 -3635 700 -3615
rect 720 -3635 730 -3615
rect 690 -3650 730 -3635
rect 835 -3565 875 -3550
rect 835 -3585 845 -3565
rect 865 -3585 875 -3565
rect 835 -3615 875 -3585
rect 835 -3635 845 -3615
rect 865 -3635 875 -3615
rect 835 -3650 875 -3635
rect 890 -3565 930 -3550
rect 890 -3585 900 -3565
rect 920 -3585 930 -3565
rect 890 -3615 930 -3585
rect 890 -3635 900 -3615
rect 920 -3635 930 -3615
rect 890 -3650 930 -3635
rect 1000 -3565 1040 -3550
rect 1000 -3585 1010 -3565
rect 1030 -3585 1040 -3565
rect 1000 -3615 1040 -3585
rect 1000 -3635 1010 -3615
rect 1030 -3635 1040 -3615
rect 1000 -3650 1040 -3635
rect 1055 -3565 1095 -3550
rect 1055 -3585 1065 -3565
rect 1085 -3585 1095 -3565
rect 1055 -3615 1095 -3585
rect 1055 -3635 1065 -3615
rect 1085 -3635 1095 -3615
rect 1055 -3650 1095 -3635
rect 1165 -3565 1205 -3550
rect 1165 -3585 1175 -3565
rect 1195 -3585 1205 -3565
rect 1165 -3615 1205 -3585
rect 1165 -3635 1175 -3615
rect 1195 -3635 1205 -3615
rect 1165 -3650 1205 -3635
rect 1220 -3565 1260 -3550
rect 1220 -3585 1230 -3565
rect 1250 -3585 1260 -3565
rect 1220 -3615 1260 -3585
rect 1220 -3635 1230 -3615
rect 1250 -3635 1260 -3615
rect 1220 -3650 1260 -3635
rect 1400 -3565 1450 -3550
rect 1400 -3585 1415 -3565
rect 1435 -3585 1450 -3565
rect 1400 -3615 1450 -3585
rect 1400 -3635 1415 -3615
rect 1435 -3635 1450 -3615
rect 1400 -3650 1450 -3635
rect 1465 -3565 1515 -3550
rect 1465 -3585 1480 -3565
rect 1500 -3585 1515 -3565
rect 1465 -3615 1515 -3585
rect 1465 -3635 1480 -3615
rect 1500 -3635 1515 -3615
rect 1465 -3650 1515 -3635
rect 1595 -3565 1645 -3550
rect 1595 -3585 1610 -3565
rect 1630 -3585 1645 -3565
rect 1595 -3615 1645 -3585
rect 1595 -3635 1610 -3615
rect 1630 -3635 1645 -3615
rect 1595 -3650 1645 -3635
rect 1660 -3565 1710 -3550
rect 1660 -3585 1675 -3565
rect 1695 -3585 1710 -3565
rect 1660 -3615 1710 -3585
rect 1660 -3635 1675 -3615
rect 1695 -3635 1710 -3615
rect 1660 -3650 1710 -3635
rect 1790 -3565 1840 -3550
rect 1790 -3585 1805 -3565
rect 1825 -3585 1840 -3565
rect 1790 -3615 1840 -3585
rect 1790 -3635 1805 -3615
rect 1825 -3635 1840 -3615
rect 1790 -3650 1840 -3635
rect 1855 -3565 1905 -3550
rect 1855 -3585 1870 -3565
rect 1890 -3585 1905 -3565
rect 1855 -3615 1905 -3585
rect 1855 -3635 1870 -3615
rect 1890 -3635 1905 -3615
rect 1855 -3650 1905 -3635
rect 1935 -3565 1985 -3550
rect 1935 -3585 1950 -3565
rect 1970 -3585 1985 -3565
rect 1935 -3615 1985 -3585
rect 1935 -3635 1950 -3615
rect 1970 -3635 1985 -3615
rect 1935 -3650 1985 -3635
rect 2000 -3565 2050 -3550
rect 2000 -3585 2015 -3565
rect 2035 -3585 2050 -3565
rect 2000 -3615 2050 -3585
rect 2000 -3635 2015 -3615
rect 2035 -3635 2050 -3615
rect 2000 -3650 2050 -3635
rect 2130 -3565 2180 -3550
rect 2130 -3585 2145 -3565
rect 2165 -3585 2180 -3565
rect 2130 -3615 2180 -3585
rect 2130 -3635 2145 -3615
rect 2165 -3635 2180 -3615
rect 2130 -3650 2180 -3635
rect 2195 -3565 2245 -3550
rect 2195 -3585 2210 -3565
rect 2230 -3585 2245 -3565
rect 2195 -3615 2245 -3585
rect 2195 -3635 2210 -3615
rect 2230 -3635 2245 -3615
rect 2195 -3650 2245 -3635
<< pdiff >>
rect -130 -2875 -90 -2860
rect -130 -2895 -120 -2875
rect -100 -2895 -90 -2875
rect -130 -2925 -90 -2895
rect -130 -2945 -120 -2925
rect -100 -2945 -90 -2925
rect -130 -2975 -90 -2945
rect -130 -2995 -120 -2975
rect -100 -2995 -90 -2975
rect -130 -3025 -90 -2995
rect -130 -3045 -120 -3025
rect -100 -3045 -90 -3025
rect -130 -3060 -90 -3045
rect -75 -2875 -35 -2860
rect -75 -2895 -65 -2875
rect -45 -2895 -35 -2875
rect -75 -2925 -35 -2895
rect -75 -2945 -65 -2925
rect -45 -2945 -35 -2925
rect -75 -2975 -35 -2945
rect -75 -2995 -65 -2975
rect -45 -2995 -35 -2975
rect -75 -3025 -35 -2995
rect -75 -3045 -65 -3025
rect -45 -3045 -35 -3025
rect -75 -3060 -35 -3045
rect -20 -2875 20 -2860
rect -20 -2895 -10 -2875
rect 10 -2895 20 -2875
rect -20 -2925 20 -2895
rect -20 -2945 -10 -2925
rect 10 -2945 20 -2925
rect -20 -2975 20 -2945
rect -20 -2995 -10 -2975
rect 10 -2995 20 -2975
rect -20 -3025 20 -2995
rect -20 -3045 -10 -3025
rect 10 -3045 20 -3025
rect -20 -3060 20 -3045
rect 130 -2875 170 -2860
rect 130 -2895 140 -2875
rect 160 -2895 170 -2875
rect 130 -2925 170 -2895
rect 130 -2945 140 -2925
rect 160 -2945 170 -2925
rect 130 -2975 170 -2945
rect 130 -2995 140 -2975
rect 160 -2995 170 -2975
rect 130 -3025 170 -2995
rect 130 -3045 140 -3025
rect 160 -3045 170 -3025
rect 130 -3060 170 -3045
rect 185 -2875 225 -2860
rect 185 -2895 195 -2875
rect 215 -2895 225 -2875
rect 185 -2925 225 -2895
rect 185 -2945 195 -2925
rect 215 -2945 225 -2925
rect 185 -2975 225 -2945
rect 185 -2995 195 -2975
rect 215 -2995 225 -2975
rect 185 -3025 225 -2995
rect 185 -3045 195 -3025
rect 215 -3045 225 -3025
rect 185 -3060 225 -3045
rect 240 -2875 280 -2860
rect 320 -2875 360 -2860
rect 240 -2895 250 -2875
rect 270 -2895 280 -2875
rect 320 -2895 330 -2875
rect 350 -2895 360 -2875
rect 240 -2925 280 -2895
rect 320 -2925 360 -2895
rect 240 -2945 250 -2925
rect 270 -2945 280 -2925
rect 320 -2945 330 -2925
rect 350 -2945 360 -2925
rect 240 -2975 280 -2945
rect 320 -2975 360 -2945
rect 240 -2995 250 -2975
rect 270 -2995 280 -2975
rect 320 -2995 330 -2975
rect 350 -2995 360 -2975
rect 240 -3025 280 -2995
rect 320 -3025 360 -2995
rect 240 -3045 250 -3025
rect 270 -3045 280 -3025
rect 320 -3045 330 -3025
rect 350 -3045 360 -3025
rect 240 -3060 280 -3045
rect 320 -3060 360 -3045
rect 375 -2875 415 -2860
rect 375 -2895 385 -2875
rect 405 -2895 415 -2875
rect 375 -2925 415 -2895
rect 375 -2945 385 -2925
rect 405 -2945 415 -2925
rect 375 -2975 415 -2945
rect 375 -2995 385 -2975
rect 405 -2995 415 -2975
rect 375 -3025 415 -2995
rect 375 -3045 385 -3025
rect 405 -3045 415 -3025
rect 375 -3060 415 -3045
rect 430 -2875 470 -2860
rect 430 -2895 440 -2875
rect 460 -2895 470 -2875
rect 430 -2925 470 -2895
rect 430 -2945 440 -2925
rect 460 -2945 470 -2925
rect 430 -2975 470 -2945
rect 430 -2995 440 -2975
rect 460 -2995 470 -2975
rect 430 -3025 470 -2995
rect 430 -3045 440 -3025
rect 460 -3045 470 -3025
rect 430 -3060 470 -3045
rect 580 -2875 620 -2860
rect 580 -2895 590 -2875
rect 610 -2895 620 -2875
rect 580 -2925 620 -2895
rect 580 -2945 590 -2925
rect 610 -2945 620 -2925
rect 580 -2975 620 -2945
rect 580 -2995 590 -2975
rect 610 -2995 620 -2975
rect 580 -3025 620 -2995
rect 580 -3045 590 -3025
rect 610 -3045 620 -3025
rect 580 -3060 620 -3045
rect 635 -2875 675 -2860
rect 635 -2895 645 -2875
rect 665 -2895 675 -2875
rect 635 -2925 675 -2895
rect 635 -2945 645 -2925
rect 665 -2945 675 -2925
rect 635 -2975 675 -2945
rect 635 -2995 645 -2975
rect 665 -2995 675 -2975
rect 635 -3025 675 -2995
rect 635 -3045 645 -3025
rect 665 -3045 675 -3025
rect 635 -3060 675 -3045
rect 690 -2875 730 -2860
rect 690 -2895 700 -2875
rect 720 -2895 730 -2875
rect 690 -2925 730 -2895
rect 690 -2945 700 -2925
rect 720 -2945 730 -2925
rect 690 -2975 730 -2945
rect 690 -2995 700 -2975
rect 720 -2995 730 -2975
rect 690 -3025 730 -2995
rect 690 -3045 700 -3025
rect 720 -3045 730 -3025
rect 690 -3060 730 -3045
rect 800 -2875 840 -2860
rect 800 -2895 810 -2875
rect 830 -2895 840 -2875
rect 800 -2925 840 -2895
rect 800 -2945 810 -2925
rect 830 -2945 840 -2925
rect 800 -2975 840 -2945
rect 800 -2995 810 -2975
rect 830 -2995 840 -2975
rect 800 -3025 840 -2995
rect 800 -3045 810 -3025
rect 830 -3045 840 -3025
rect 800 -3060 840 -3045
rect 855 -2875 895 -2860
rect 855 -2895 865 -2875
rect 885 -2895 895 -2875
rect 855 -2925 895 -2895
rect 855 -2945 865 -2925
rect 885 -2945 895 -2925
rect 855 -2975 895 -2945
rect 855 -2995 865 -2975
rect 885 -2995 895 -2975
rect 855 -3025 895 -2995
rect 855 -3045 865 -3025
rect 885 -3045 895 -3025
rect 855 -3060 895 -3045
rect 910 -2875 950 -2860
rect 910 -2895 920 -2875
rect 940 -2895 950 -2875
rect 910 -2925 950 -2895
rect 910 -2945 920 -2925
rect 940 -2945 950 -2925
rect 910 -2975 950 -2945
rect 910 -2995 920 -2975
rect 940 -2995 950 -2975
rect 910 -3025 950 -2995
rect 910 -3045 920 -3025
rect 940 -3045 950 -3025
rect 910 -3060 950 -3045
rect 1020 -2875 1060 -2860
rect 1020 -2895 1030 -2875
rect 1050 -2895 1060 -2875
rect 1020 -2925 1060 -2895
rect 1020 -2945 1030 -2925
rect 1050 -2945 1060 -2925
rect 1020 -2975 1060 -2945
rect 1020 -2995 1030 -2975
rect 1050 -2995 1060 -2975
rect 1020 -3025 1060 -2995
rect 1020 -3045 1030 -3025
rect 1050 -3045 1060 -3025
rect 1020 -3060 1060 -3045
rect 1075 -2875 1115 -2860
rect 1075 -2895 1085 -2875
rect 1105 -2895 1115 -2875
rect 1075 -2925 1115 -2895
rect 1075 -2945 1085 -2925
rect 1105 -2945 1115 -2925
rect 1075 -2975 1115 -2945
rect 1075 -2995 1085 -2975
rect 1105 -2995 1115 -2975
rect 1075 -3025 1115 -2995
rect 1075 -3045 1085 -3025
rect 1105 -3045 1115 -3025
rect 1075 -3060 1115 -3045
rect 1185 -2875 1225 -2860
rect 1185 -2895 1195 -2875
rect 1215 -2895 1225 -2875
rect 1185 -2925 1225 -2895
rect 1185 -2945 1195 -2925
rect 1215 -2945 1225 -2925
rect 1185 -2975 1225 -2945
rect 1185 -2995 1195 -2975
rect 1215 -2995 1225 -2975
rect 1185 -3025 1225 -2995
rect 1185 -3045 1195 -3025
rect 1215 -3045 1225 -3025
rect 1185 -3060 1225 -3045
rect 1240 -2875 1280 -2860
rect 1240 -2895 1250 -2875
rect 1270 -2895 1280 -2875
rect 1240 -2925 1280 -2895
rect 1240 -2945 1250 -2925
rect 1270 -2945 1280 -2925
rect 1240 -2975 1280 -2945
rect 1240 -2995 1250 -2975
rect 1270 -2995 1280 -2975
rect 1240 -3025 1280 -2995
rect 1240 -3045 1250 -3025
rect 1270 -3045 1280 -3025
rect 1240 -3060 1280 -3045
rect 1400 -2875 1450 -2860
rect 1400 -2895 1415 -2875
rect 1435 -2895 1450 -2875
rect 1400 -2925 1450 -2895
rect 1400 -2945 1415 -2925
rect 1435 -2945 1450 -2925
rect 1400 -2975 1450 -2945
rect 1400 -2995 1415 -2975
rect 1435 -2995 1450 -2975
rect 1400 -3025 1450 -2995
rect 1400 -3045 1415 -3025
rect 1435 -3045 1450 -3025
rect 1400 -3060 1450 -3045
rect 1465 -2875 1515 -2860
rect 1465 -2895 1480 -2875
rect 1500 -2895 1515 -2875
rect 1465 -2925 1515 -2895
rect 1465 -2945 1480 -2925
rect 1500 -2945 1515 -2925
rect 1465 -2975 1515 -2945
rect 1465 -2995 1480 -2975
rect 1500 -2995 1515 -2975
rect 1465 -3025 1515 -2995
rect 1465 -3045 1480 -3025
rect 1500 -3045 1515 -3025
rect 1465 -3060 1515 -3045
rect 1595 -2875 1645 -2860
rect 1595 -2895 1610 -2875
rect 1630 -2895 1645 -2875
rect 1595 -2925 1645 -2895
rect 1595 -2945 1610 -2925
rect 1630 -2945 1645 -2925
rect 1595 -2975 1645 -2945
rect 1595 -2995 1610 -2975
rect 1630 -2995 1645 -2975
rect 1595 -3025 1645 -2995
rect 1595 -3045 1610 -3025
rect 1630 -3045 1645 -3025
rect 1595 -3060 1645 -3045
rect 1660 -2875 1710 -2860
rect 1660 -2895 1675 -2875
rect 1695 -2895 1710 -2875
rect 1660 -2925 1710 -2895
rect 1660 -2945 1675 -2925
rect 1695 -2945 1710 -2925
rect 1660 -2975 1710 -2945
rect 1660 -2995 1675 -2975
rect 1695 -2995 1710 -2975
rect 1660 -3025 1710 -2995
rect 1660 -3045 1675 -3025
rect 1695 -3045 1710 -3025
rect 1660 -3060 1710 -3045
rect 1790 -2875 1840 -2860
rect 1790 -2895 1805 -2875
rect 1825 -2895 1840 -2875
rect 1790 -2925 1840 -2895
rect 1790 -2945 1805 -2925
rect 1825 -2945 1840 -2925
rect 1790 -2975 1840 -2945
rect 1790 -2995 1805 -2975
rect 1825 -2995 1840 -2975
rect 1790 -3025 1840 -2995
rect 1790 -3045 1805 -3025
rect 1825 -3045 1840 -3025
rect 1790 -3060 1840 -3045
rect 1855 -2875 1905 -2860
rect 1855 -2895 1870 -2875
rect 1890 -2895 1905 -2875
rect 1855 -2925 1905 -2895
rect 1855 -2945 1870 -2925
rect 1890 -2945 1905 -2925
rect 1855 -2975 1905 -2945
rect 1855 -2995 1870 -2975
rect 1890 -2995 1905 -2975
rect 1855 -3025 1905 -2995
rect 1855 -3045 1870 -3025
rect 1890 -3045 1905 -3025
rect 1855 -3060 1905 -3045
rect 1935 -2875 1985 -2860
rect 1935 -2895 1950 -2875
rect 1970 -2895 1985 -2875
rect 1935 -2925 1985 -2895
rect 1935 -2945 1950 -2925
rect 1970 -2945 1985 -2925
rect 1935 -2975 1985 -2945
rect 1935 -2995 1950 -2975
rect 1970 -2995 1985 -2975
rect 1935 -3025 1985 -2995
rect 1935 -3045 1950 -3025
rect 1970 -3045 1985 -3025
rect 1935 -3060 1985 -3045
rect 2000 -2875 2050 -2860
rect 2000 -2895 2015 -2875
rect 2035 -2895 2050 -2875
rect 2000 -2925 2050 -2895
rect 2000 -2945 2015 -2925
rect 2035 -2945 2050 -2925
rect 2000 -2975 2050 -2945
rect 2000 -2995 2015 -2975
rect 2035 -2995 2050 -2975
rect 2000 -3025 2050 -2995
rect 2000 -3045 2015 -3025
rect 2035 -3045 2050 -3025
rect 2000 -3060 2050 -3045
rect 2130 -2875 2180 -2860
rect 2130 -2895 2145 -2875
rect 2165 -2895 2180 -2875
rect 2130 -2925 2180 -2895
rect 2130 -2945 2145 -2925
rect 2165 -2945 2180 -2925
rect 2130 -2975 2180 -2945
rect 2130 -2995 2145 -2975
rect 2165 -2995 2180 -2975
rect 2130 -3025 2180 -2995
rect 2130 -3045 2145 -3025
rect 2165 -3045 2180 -3025
rect 2130 -3060 2180 -3045
rect 2195 -2875 2245 -2860
rect 2195 -2895 2210 -2875
rect 2230 -2895 2245 -2875
rect 2195 -2925 2245 -2895
rect 2195 -2945 2210 -2925
rect 2230 -2945 2245 -2925
rect 2195 -2975 2245 -2945
rect 2195 -2995 2210 -2975
rect 2230 -2995 2245 -2975
rect 2195 -3025 2245 -2995
rect 2195 -3045 2210 -3025
rect 2230 -3045 2245 -3025
rect 2195 -3060 2245 -3045
rect -130 -3255 -90 -3240
rect -130 -3275 -120 -3255
rect -100 -3275 -90 -3255
rect -130 -3305 -90 -3275
rect -130 -3325 -120 -3305
rect -100 -3325 -90 -3305
rect -130 -3355 -90 -3325
rect -130 -3375 -120 -3355
rect -100 -3375 -90 -3355
rect -130 -3405 -90 -3375
rect -130 -3425 -120 -3405
rect -100 -3425 -90 -3405
rect -130 -3440 -90 -3425
rect -75 -3255 -35 -3240
rect -75 -3275 -65 -3255
rect -45 -3275 -35 -3255
rect -75 -3305 -35 -3275
rect -75 -3325 -65 -3305
rect -45 -3325 -35 -3305
rect -75 -3355 -35 -3325
rect -75 -3375 -65 -3355
rect -45 -3375 -35 -3355
rect -75 -3405 -35 -3375
rect -75 -3425 -65 -3405
rect -45 -3425 -35 -3405
rect -75 -3440 -35 -3425
rect -20 -3255 20 -3240
rect -20 -3275 -10 -3255
rect 10 -3275 20 -3255
rect -20 -3305 20 -3275
rect -20 -3325 -10 -3305
rect 10 -3325 20 -3305
rect -20 -3355 20 -3325
rect -20 -3375 -10 -3355
rect 10 -3375 20 -3355
rect -20 -3405 20 -3375
rect -20 -3425 -10 -3405
rect 10 -3425 20 -3405
rect -20 -3440 20 -3425
rect 130 -3255 170 -3240
rect 130 -3275 140 -3255
rect 160 -3275 170 -3255
rect 130 -3305 170 -3275
rect 130 -3325 140 -3305
rect 160 -3325 170 -3305
rect 130 -3355 170 -3325
rect 130 -3375 140 -3355
rect 160 -3375 170 -3355
rect 130 -3405 170 -3375
rect 130 -3425 140 -3405
rect 160 -3425 170 -3405
rect 130 -3440 170 -3425
rect 185 -3255 225 -3240
rect 185 -3275 195 -3255
rect 215 -3275 225 -3255
rect 185 -3305 225 -3275
rect 185 -3325 195 -3305
rect 215 -3325 225 -3305
rect 185 -3355 225 -3325
rect 185 -3375 195 -3355
rect 215 -3375 225 -3355
rect 185 -3405 225 -3375
rect 185 -3425 195 -3405
rect 215 -3425 225 -3405
rect 185 -3440 225 -3425
rect 240 -3255 280 -3240
rect 320 -3255 360 -3240
rect 240 -3275 250 -3255
rect 270 -3275 280 -3255
rect 320 -3275 330 -3255
rect 350 -3275 360 -3255
rect 240 -3305 280 -3275
rect 320 -3305 360 -3275
rect 240 -3325 250 -3305
rect 270 -3325 280 -3305
rect 320 -3325 330 -3305
rect 350 -3325 360 -3305
rect 240 -3355 280 -3325
rect 320 -3355 360 -3325
rect 240 -3375 250 -3355
rect 270 -3375 280 -3355
rect 320 -3375 330 -3355
rect 350 -3375 360 -3355
rect 240 -3405 280 -3375
rect 320 -3405 360 -3375
rect 240 -3425 250 -3405
rect 270 -3425 280 -3405
rect 320 -3425 330 -3405
rect 350 -3425 360 -3405
rect 240 -3440 280 -3425
rect 320 -3440 360 -3425
rect 375 -3255 415 -3240
rect 375 -3275 385 -3255
rect 405 -3275 415 -3255
rect 375 -3305 415 -3275
rect 375 -3325 385 -3305
rect 405 -3325 415 -3305
rect 375 -3355 415 -3325
rect 375 -3375 385 -3355
rect 405 -3375 415 -3355
rect 375 -3405 415 -3375
rect 375 -3425 385 -3405
rect 405 -3425 415 -3405
rect 375 -3440 415 -3425
rect 430 -3255 470 -3240
rect 430 -3275 440 -3255
rect 460 -3275 470 -3255
rect 430 -3305 470 -3275
rect 430 -3325 440 -3305
rect 460 -3325 470 -3305
rect 430 -3355 470 -3325
rect 430 -3375 440 -3355
rect 460 -3375 470 -3355
rect 430 -3405 470 -3375
rect 430 -3425 440 -3405
rect 460 -3425 470 -3405
rect 430 -3440 470 -3425
rect 580 -3255 620 -3240
rect 580 -3275 590 -3255
rect 610 -3275 620 -3255
rect 580 -3305 620 -3275
rect 580 -3325 590 -3305
rect 610 -3325 620 -3305
rect 580 -3355 620 -3325
rect 580 -3375 590 -3355
rect 610 -3375 620 -3355
rect 580 -3405 620 -3375
rect 580 -3425 590 -3405
rect 610 -3425 620 -3405
rect 580 -3440 620 -3425
rect 635 -3255 675 -3240
rect 635 -3275 645 -3255
rect 665 -3275 675 -3255
rect 635 -3305 675 -3275
rect 635 -3325 645 -3305
rect 665 -3325 675 -3305
rect 635 -3355 675 -3325
rect 635 -3375 645 -3355
rect 665 -3375 675 -3355
rect 635 -3405 675 -3375
rect 635 -3425 645 -3405
rect 665 -3425 675 -3405
rect 635 -3440 675 -3425
rect 690 -3255 730 -3240
rect 690 -3275 700 -3255
rect 720 -3275 730 -3255
rect 690 -3305 730 -3275
rect 690 -3325 700 -3305
rect 720 -3325 730 -3305
rect 690 -3355 730 -3325
rect 690 -3375 700 -3355
rect 720 -3375 730 -3355
rect 690 -3405 730 -3375
rect 690 -3425 700 -3405
rect 720 -3425 730 -3405
rect 690 -3440 730 -3425
rect 835 -3255 875 -3240
rect 835 -3275 845 -3255
rect 865 -3275 875 -3255
rect 835 -3305 875 -3275
rect 835 -3325 845 -3305
rect 865 -3325 875 -3305
rect 835 -3355 875 -3325
rect 835 -3375 845 -3355
rect 865 -3375 875 -3355
rect 835 -3405 875 -3375
rect 835 -3425 845 -3405
rect 865 -3425 875 -3405
rect 835 -3440 875 -3425
rect 890 -3255 930 -3240
rect 890 -3275 900 -3255
rect 920 -3275 930 -3255
rect 890 -3305 930 -3275
rect 890 -3325 900 -3305
rect 920 -3325 930 -3305
rect 890 -3355 930 -3325
rect 890 -3375 900 -3355
rect 920 -3375 930 -3355
rect 890 -3405 930 -3375
rect 890 -3425 900 -3405
rect 920 -3425 930 -3405
rect 890 -3440 930 -3425
rect 1000 -3255 1040 -3240
rect 1000 -3275 1010 -3255
rect 1030 -3275 1040 -3255
rect 1000 -3305 1040 -3275
rect 1000 -3325 1010 -3305
rect 1030 -3325 1040 -3305
rect 1000 -3355 1040 -3325
rect 1000 -3375 1010 -3355
rect 1030 -3375 1040 -3355
rect 1000 -3405 1040 -3375
rect 1000 -3425 1010 -3405
rect 1030 -3425 1040 -3405
rect 1000 -3440 1040 -3425
rect 1055 -3255 1095 -3240
rect 1055 -3275 1065 -3255
rect 1085 -3275 1095 -3255
rect 1055 -3305 1095 -3275
rect 1055 -3325 1065 -3305
rect 1085 -3325 1095 -3305
rect 1055 -3355 1095 -3325
rect 1055 -3375 1065 -3355
rect 1085 -3375 1095 -3355
rect 1055 -3405 1095 -3375
rect 1055 -3425 1065 -3405
rect 1085 -3425 1095 -3405
rect 1055 -3440 1095 -3425
rect 1165 -3255 1205 -3240
rect 1165 -3275 1175 -3255
rect 1195 -3275 1205 -3255
rect 1165 -3305 1205 -3275
rect 1165 -3325 1175 -3305
rect 1195 -3325 1205 -3305
rect 1165 -3355 1205 -3325
rect 1165 -3375 1175 -3355
rect 1195 -3375 1205 -3355
rect 1165 -3405 1205 -3375
rect 1165 -3425 1175 -3405
rect 1195 -3425 1205 -3405
rect 1165 -3440 1205 -3425
rect 1220 -3255 1260 -3240
rect 1220 -3275 1230 -3255
rect 1250 -3275 1260 -3255
rect 1220 -3305 1260 -3275
rect 1220 -3325 1230 -3305
rect 1250 -3325 1260 -3305
rect 1220 -3355 1260 -3325
rect 1220 -3375 1230 -3355
rect 1250 -3375 1260 -3355
rect 1220 -3405 1260 -3375
rect 1220 -3425 1230 -3405
rect 1250 -3425 1260 -3405
rect 1220 -3440 1260 -3425
rect 1400 -3255 1450 -3240
rect 1400 -3275 1415 -3255
rect 1435 -3275 1450 -3255
rect 1400 -3305 1450 -3275
rect 1400 -3325 1415 -3305
rect 1435 -3325 1450 -3305
rect 1400 -3355 1450 -3325
rect 1400 -3375 1415 -3355
rect 1435 -3375 1450 -3355
rect 1400 -3405 1450 -3375
rect 1400 -3425 1415 -3405
rect 1435 -3425 1450 -3405
rect 1400 -3440 1450 -3425
rect 1465 -3255 1515 -3240
rect 1465 -3275 1480 -3255
rect 1500 -3275 1515 -3255
rect 1465 -3305 1515 -3275
rect 1465 -3325 1480 -3305
rect 1500 -3325 1515 -3305
rect 1465 -3355 1515 -3325
rect 1465 -3375 1480 -3355
rect 1500 -3375 1515 -3355
rect 1465 -3405 1515 -3375
rect 1465 -3425 1480 -3405
rect 1500 -3425 1515 -3405
rect 1465 -3440 1515 -3425
rect 1595 -3255 1645 -3240
rect 1595 -3275 1610 -3255
rect 1630 -3275 1645 -3255
rect 1595 -3305 1645 -3275
rect 1595 -3325 1610 -3305
rect 1630 -3325 1645 -3305
rect 1595 -3355 1645 -3325
rect 1595 -3375 1610 -3355
rect 1630 -3375 1645 -3355
rect 1595 -3405 1645 -3375
rect 1595 -3425 1610 -3405
rect 1630 -3425 1645 -3405
rect 1595 -3440 1645 -3425
rect 1660 -3255 1710 -3240
rect 1660 -3275 1675 -3255
rect 1695 -3275 1710 -3255
rect 1660 -3305 1710 -3275
rect 1660 -3325 1675 -3305
rect 1695 -3325 1710 -3305
rect 1660 -3355 1710 -3325
rect 1660 -3375 1675 -3355
rect 1695 -3375 1710 -3355
rect 1660 -3405 1710 -3375
rect 1660 -3425 1675 -3405
rect 1695 -3425 1710 -3405
rect 1660 -3440 1710 -3425
rect 1790 -3255 1840 -3240
rect 1790 -3275 1805 -3255
rect 1825 -3275 1840 -3255
rect 1790 -3305 1840 -3275
rect 1790 -3325 1805 -3305
rect 1825 -3325 1840 -3305
rect 1790 -3355 1840 -3325
rect 1790 -3375 1805 -3355
rect 1825 -3375 1840 -3355
rect 1790 -3405 1840 -3375
rect 1790 -3425 1805 -3405
rect 1825 -3425 1840 -3405
rect 1790 -3440 1840 -3425
rect 1855 -3255 1905 -3240
rect 1855 -3275 1870 -3255
rect 1890 -3275 1905 -3255
rect 1855 -3305 1905 -3275
rect 1855 -3325 1870 -3305
rect 1890 -3325 1905 -3305
rect 1855 -3355 1905 -3325
rect 1855 -3375 1870 -3355
rect 1890 -3375 1905 -3355
rect 1855 -3405 1905 -3375
rect 1855 -3425 1870 -3405
rect 1890 -3425 1905 -3405
rect 1855 -3440 1905 -3425
rect 1935 -3255 1985 -3240
rect 1935 -3275 1950 -3255
rect 1970 -3275 1985 -3255
rect 1935 -3305 1985 -3275
rect 1935 -3325 1950 -3305
rect 1970 -3325 1985 -3305
rect 1935 -3355 1985 -3325
rect 1935 -3375 1950 -3355
rect 1970 -3375 1985 -3355
rect 1935 -3405 1985 -3375
rect 1935 -3425 1950 -3405
rect 1970 -3425 1985 -3405
rect 1935 -3440 1985 -3425
rect 2000 -3255 2050 -3240
rect 2000 -3275 2015 -3255
rect 2035 -3275 2050 -3255
rect 2000 -3305 2050 -3275
rect 2000 -3325 2015 -3305
rect 2035 -3325 2050 -3305
rect 2000 -3355 2050 -3325
rect 2000 -3375 2015 -3355
rect 2035 -3375 2050 -3355
rect 2000 -3405 2050 -3375
rect 2000 -3425 2015 -3405
rect 2035 -3425 2050 -3405
rect 2000 -3440 2050 -3425
<< ndiffc >>
rect -120 -2685 -100 -2665
rect -120 -2735 -100 -2715
rect -65 -2685 -45 -2665
rect -65 -2735 -45 -2715
rect -10 -2685 10 -2665
rect -10 -2735 10 -2715
rect 140 -2685 160 -2665
rect 140 -2735 160 -2715
rect 195 -2685 215 -2665
rect 195 -2735 215 -2715
rect 250 -2685 270 -2665
rect 330 -2685 350 -2665
rect 250 -2735 270 -2715
rect 330 -2735 350 -2715
rect 385 -2685 405 -2665
rect 385 -2735 405 -2715
rect 440 -2685 460 -2665
rect 440 -2735 460 -2715
rect 590 -2685 610 -2665
rect 590 -2735 610 -2715
rect 645 -2685 665 -2665
rect 645 -2735 665 -2715
rect 700 -2685 720 -2665
rect 700 -2735 720 -2715
rect 810 -2685 830 -2665
rect 810 -2735 830 -2715
rect 865 -2685 885 -2665
rect 865 -2735 885 -2715
rect 920 -2685 940 -2665
rect 920 -2735 940 -2715
rect 1030 -2685 1050 -2665
rect 1030 -2735 1050 -2715
rect 1085 -2685 1105 -2665
rect 1085 -2735 1105 -2715
rect 1195 -2685 1215 -2665
rect 1195 -2735 1215 -2715
rect 1250 -2685 1270 -2665
rect 1250 -2735 1270 -2715
rect 1415 -2685 1435 -2665
rect 1415 -2735 1435 -2715
rect 1480 -2685 1500 -2665
rect 1480 -2735 1500 -2715
rect 1610 -2685 1630 -2665
rect 1610 -2735 1630 -2715
rect 1675 -2685 1695 -2665
rect 1675 -2735 1695 -2715
rect 1805 -2685 1825 -2665
rect 1805 -2735 1825 -2715
rect 1870 -2685 1890 -2665
rect 1870 -2735 1890 -2715
rect 1950 -2685 1970 -2665
rect 1950 -2735 1970 -2715
rect 2015 -2685 2035 -2665
rect 2015 -2735 2035 -2715
rect -120 -3585 -100 -3565
rect -120 -3635 -100 -3615
rect -65 -3585 -45 -3565
rect -65 -3635 -45 -3615
rect -10 -3585 10 -3565
rect -10 -3635 10 -3615
rect 140 -3585 160 -3565
rect 140 -3635 160 -3615
rect 195 -3585 215 -3565
rect 195 -3635 215 -3615
rect 250 -3585 270 -3565
rect 330 -3585 350 -3565
rect 250 -3635 270 -3615
rect 330 -3635 350 -3615
rect 385 -3585 405 -3565
rect 385 -3635 405 -3615
rect 440 -3585 460 -3565
rect 440 -3635 460 -3615
rect 590 -3585 610 -3565
rect 590 -3635 610 -3615
rect 645 -3585 665 -3565
rect 645 -3635 665 -3615
rect 700 -3585 720 -3565
rect 700 -3635 720 -3615
rect 845 -3585 865 -3565
rect 845 -3635 865 -3615
rect 900 -3585 920 -3565
rect 900 -3635 920 -3615
rect 1010 -3585 1030 -3565
rect 1010 -3635 1030 -3615
rect 1065 -3585 1085 -3565
rect 1065 -3635 1085 -3615
rect 1175 -3585 1195 -3565
rect 1175 -3635 1195 -3615
rect 1230 -3585 1250 -3565
rect 1230 -3635 1250 -3615
rect 1415 -3585 1435 -3565
rect 1415 -3635 1435 -3615
rect 1480 -3585 1500 -3565
rect 1480 -3635 1500 -3615
rect 1610 -3585 1630 -3565
rect 1610 -3635 1630 -3615
rect 1675 -3585 1695 -3565
rect 1675 -3635 1695 -3615
rect 1805 -3585 1825 -3565
rect 1805 -3635 1825 -3615
rect 1870 -3585 1890 -3565
rect 1870 -3635 1890 -3615
rect 1950 -3585 1970 -3565
rect 1950 -3635 1970 -3615
rect 2015 -3585 2035 -3565
rect 2015 -3635 2035 -3615
rect 2145 -3585 2165 -3565
rect 2145 -3635 2165 -3615
rect 2210 -3585 2230 -3565
rect 2210 -3635 2230 -3615
<< pdiffc >>
rect -120 -2895 -100 -2875
rect -120 -2945 -100 -2925
rect -120 -2995 -100 -2975
rect -120 -3045 -100 -3025
rect -65 -2895 -45 -2875
rect -65 -2945 -45 -2925
rect -65 -2995 -45 -2975
rect -65 -3045 -45 -3025
rect -10 -2895 10 -2875
rect -10 -2945 10 -2925
rect -10 -2995 10 -2975
rect -10 -3045 10 -3025
rect 140 -2895 160 -2875
rect 140 -2945 160 -2925
rect 140 -2995 160 -2975
rect 140 -3045 160 -3025
rect 195 -2895 215 -2875
rect 195 -2945 215 -2925
rect 195 -2995 215 -2975
rect 195 -3045 215 -3025
rect 250 -2895 270 -2875
rect 330 -2895 350 -2875
rect 250 -2945 270 -2925
rect 330 -2945 350 -2925
rect 250 -2995 270 -2975
rect 330 -2995 350 -2975
rect 250 -3045 270 -3025
rect 330 -3045 350 -3025
rect 385 -2895 405 -2875
rect 385 -2945 405 -2925
rect 385 -2995 405 -2975
rect 385 -3045 405 -3025
rect 440 -2895 460 -2875
rect 440 -2945 460 -2925
rect 440 -2995 460 -2975
rect 440 -3045 460 -3025
rect 590 -2895 610 -2875
rect 590 -2945 610 -2925
rect 590 -2995 610 -2975
rect 590 -3045 610 -3025
rect 645 -2895 665 -2875
rect 645 -2945 665 -2925
rect 645 -2995 665 -2975
rect 645 -3045 665 -3025
rect 700 -2895 720 -2875
rect 700 -2945 720 -2925
rect 700 -2995 720 -2975
rect 700 -3045 720 -3025
rect 810 -2895 830 -2875
rect 810 -2945 830 -2925
rect 810 -2995 830 -2975
rect 810 -3045 830 -3025
rect 865 -2895 885 -2875
rect 865 -2945 885 -2925
rect 865 -2995 885 -2975
rect 865 -3045 885 -3025
rect 920 -2895 940 -2875
rect 920 -2945 940 -2925
rect 920 -2995 940 -2975
rect 920 -3045 940 -3025
rect 1030 -2895 1050 -2875
rect 1030 -2945 1050 -2925
rect 1030 -2995 1050 -2975
rect 1030 -3045 1050 -3025
rect 1085 -2895 1105 -2875
rect 1085 -2945 1105 -2925
rect 1085 -2995 1105 -2975
rect 1085 -3045 1105 -3025
rect 1195 -2895 1215 -2875
rect 1195 -2945 1215 -2925
rect 1195 -2995 1215 -2975
rect 1195 -3045 1215 -3025
rect 1250 -2895 1270 -2875
rect 1250 -2945 1270 -2925
rect 1250 -2995 1270 -2975
rect 1250 -3045 1270 -3025
rect 1415 -2895 1435 -2875
rect 1415 -2945 1435 -2925
rect 1415 -2995 1435 -2975
rect 1415 -3045 1435 -3025
rect 1480 -2895 1500 -2875
rect 1480 -2945 1500 -2925
rect 1480 -2995 1500 -2975
rect 1480 -3045 1500 -3025
rect 1610 -2895 1630 -2875
rect 1610 -2945 1630 -2925
rect 1610 -2995 1630 -2975
rect 1610 -3045 1630 -3025
rect 1675 -2895 1695 -2875
rect 1675 -2945 1695 -2925
rect 1675 -2995 1695 -2975
rect 1675 -3045 1695 -3025
rect 1805 -2895 1825 -2875
rect 1805 -2945 1825 -2925
rect 1805 -2995 1825 -2975
rect 1805 -3045 1825 -3025
rect 1870 -2895 1890 -2875
rect 1870 -2945 1890 -2925
rect 1870 -2995 1890 -2975
rect 1870 -3045 1890 -3025
rect 1950 -2895 1970 -2875
rect 1950 -2945 1970 -2925
rect 1950 -2995 1970 -2975
rect 1950 -3045 1970 -3025
rect 2015 -2895 2035 -2875
rect 2015 -2945 2035 -2925
rect 2015 -2995 2035 -2975
rect 2015 -3045 2035 -3025
rect 2145 -2895 2165 -2875
rect 2145 -2945 2165 -2925
rect 2145 -2995 2165 -2975
rect 2145 -3045 2165 -3025
rect 2210 -2895 2230 -2875
rect 2210 -2945 2230 -2925
rect 2210 -2995 2230 -2975
rect 2210 -3045 2230 -3025
rect -120 -3275 -100 -3255
rect -120 -3325 -100 -3305
rect -120 -3375 -100 -3355
rect -120 -3425 -100 -3405
rect -65 -3275 -45 -3255
rect -65 -3325 -45 -3305
rect -65 -3375 -45 -3355
rect -65 -3425 -45 -3405
rect -10 -3275 10 -3255
rect -10 -3325 10 -3305
rect -10 -3375 10 -3355
rect -10 -3425 10 -3405
rect 140 -3275 160 -3255
rect 140 -3325 160 -3305
rect 140 -3375 160 -3355
rect 140 -3425 160 -3405
rect 195 -3275 215 -3255
rect 195 -3325 215 -3305
rect 195 -3375 215 -3355
rect 195 -3425 215 -3405
rect 250 -3275 270 -3255
rect 330 -3275 350 -3255
rect 250 -3325 270 -3305
rect 330 -3325 350 -3305
rect 250 -3375 270 -3355
rect 330 -3375 350 -3355
rect 250 -3425 270 -3405
rect 330 -3425 350 -3405
rect 385 -3275 405 -3255
rect 385 -3325 405 -3305
rect 385 -3375 405 -3355
rect 385 -3425 405 -3405
rect 440 -3275 460 -3255
rect 440 -3325 460 -3305
rect 440 -3375 460 -3355
rect 440 -3425 460 -3405
rect 590 -3275 610 -3255
rect 590 -3325 610 -3305
rect 590 -3375 610 -3355
rect 590 -3425 610 -3405
rect 645 -3275 665 -3255
rect 645 -3325 665 -3305
rect 645 -3375 665 -3355
rect 645 -3425 665 -3405
rect 700 -3275 720 -3255
rect 700 -3325 720 -3305
rect 700 -3375 720 -3355
rect 700 -3425 720 -3405
rect 845 -3275 865 -3255
rect 845 -3325 865 -3305
rect 845 -3375 865 -3355
rect 845 -3425 865 -3405
rect 900 -3275 920 -3255
rect 900 -3325 920 -3305
rect 900 -3375 920 -3355
rect 900 -3425 920 -3405
rect 1010 -3275 1030 -3255
rect 1010 -3325 1030 -3305
rect 1010 -3375 1030 -3355
rect 1010 -3425 1030 -3405
rect 1065 -3275 1085 -3255
rect 1065 -3325 1085 -3305
rect 1065 -3375 1085 -3355
rect 1065 -3425 1085 -3405
rect 1175 -3275 1195 -3255
rect 1175 -3325 1195 -3305
rect 1175 -3375 1195 -3355
rect 1175 -3425 1195 -3405
rect 1230 -3275 1250 -3255
rect 1230 -3325 1250 -3305
rect 1230 -3375 1250 -3355
rect 1230 -3425 1250 -3405
rect 1415 -3275 1435 -3255
rect 1415 -3325 1435 -3305
rect 1415 -3375 1435 -3355
rect 1415 -3425 1435 -3405
rect 1480 -3275 1500 -3255
rect 1480 -3325 1500 -3305
rect 1480 -3375 1500 -3355
rect 1480 -3425 1500 -3405
rect 1610 -3275 1630 -3255
rect 1610 -3325 1630 -3305
rect 1610 -3375 1630 -3355
rect 1610 -3425 1630 -3405
rect 1675 -3275 1695 -3255
rect 1675 -3325 1695 -3305
rect 1675 -3375 1695 -3355
rect 1675 -3425 1695 -3405
rect 1805 -3275 1825 -3255
rect 1805 -3325 1825 -3305
rect 1805 -3375 1825 -3355
rect 1805 -3425 1825 -3405
rect 1870 -3275 1890 -3255
rect 1870 -3325 1890 -3305
rect 1870 -3375 1890 -3355
rect 1870 -3425 1890 -3405
rect 1950 -3275 1970 -3255
rect 1950 -3325 1970 -3305
rect 1950 -3375 1970 -3355
rect 1950 -3425 1970 -3405
rect 2015 -3275 2035 -3255
rect 2015 -3325 2035 -3305
rect 2015 -3375 2035 -3355
rect 2015 -3425 2035 -3405
<< psubdiff >>
rect -170 -2665 -130 -2650
rect -170 -2685 -160 -2665
rect -140 -2685 -130 -2665
rect -170 -2715 -130 -2685
rect -170 -2735 -160 -2715
rect -140 -2735 -130 -2715
rect -170 -2750 -130 -2735
rect 280 -2665 320 -2650
rect 280 -2685 290 -2665
rect 310 -2685 320 -2665
rect 280 -2715 320 -2685
rect 280 -2735 290 -2715
rect 310 -2735 320 -2715
rect 280 -2750 320 -2735
rect 730 -2665 770 -2650
rect 730 -2685 740 -2665
rect 760 -2685 770 -2665
rect 730 -2715 770 -2685
rect 730 -2735 740 -2715
rect 760 -2735 770 -2715
rect 730 -2750 770 -2735
rect 980 -2665 1020 -2650
rect 980 -2685 990 -2665
rect 1010 -2685 1020 -2665
rect 980 -2715 1020 -2685
rect 980 -2735 990 -2715
rect 1010 -2735 1020 -2715
rect 980 -2750 1020 -2735
rect 1145 -2665 1185 -2650
rect 1145 -2685 1155 -2665
rect 1175 -2685 1185 -2665
rect 1145 -2715 1185 -2685
rect 1145 -2735 1155 -2715
rect 1175 -2735 1185 -2715
rect 1145 -2750 1185 -2735
rect 1360 -2665 1400 -2650
rect 1360 -2685 1370 -2665
rect 1390 -2685 1400 -2665
rect 1360 -2715 1400 -2685
rect 1360 -2735 1370 -2715
rect 1390 -2735 1400 -2715
rect 1360 -2750 1400 -2735
rect 1555 -2665 1595 -2650
rect 1555 -2685 1565 -2665
rect 1585 -2685 1595 -2665
rect 1555 -2715 1595 -2685
rect 1555 -2735 1565 -2715
rect 1585 -2735 1595 -2715
rect 1555 -2750 1595 -2735
rect 1750 -2665 1790 -2650
rect 1750 -2685 1760 -2665
rect 1780 -2685 1790 -2665
rect 1750 -2715 1790 -2685
rect 1750 -2735 1760 -2715
rect 1780 -2735 1790 -2715
rect 1750 -2750 1790 -2735
rect -170 -3565 -130 -3550
rect -170 -3585 -160 -3565
rect -140 -3585 -130 -3565
rect -170 -3615 -130 -3585
rect -170 -3635 -160 -3615
rect -140 -3635 -130 -3615
rect -170 -3650 -130 -3635
rect 280 -3565 320 -3550
rect 280 -3585 290 -3565
rect 310 -3585 320 -3565
rect 280 -3615 320 -3585
rect 280 -3635 290 -3615
rect 310 -3635 320 -3615
rect 280 -3650 320 -3635
rect 730 -3565 770 -3550
rect 730 -3585 740 -3565
rect 760 -3585 770 -3565
rect 730 -3615 770 -3585
rect 730 -3635 740 -3615
rect 760 -3635 770 -3615
rect 730 -3650 770 -3635
rect 930 -3565 970 -3550
rect 930 -3585 940 -3565
rect 960 -3585 970 -3565
rect 930 -3615 970 -3585
rect 930 -3635 940 -3615
rect 960 -3635 970 -3615
rect 930 -3650 970 -3635
rect 1095 -3565 1135 -3550
rect 1095 -3585 1105 -3565
rect 1125 -3585 1135 -3565
rect 1095 -3615 1135 -3585
rect 1095 -3635 1105 -3615
rect 1125 -3635 1135 -3615
rect 1095 -3650 1135 -3635
rect 1260 -3565 1300 -3550
rect 1260 -3585 1270 -3565
rect 1290 -3585 1300 -3565
rect 1260 -3615 1300 -3585
rect 1260 -3635 1270 -3615
rect 1290 -3635 1300 -3615
rect 1260 -3650 1300 -3635
rect 1350 -3565 1400 -3550
rect 1350 -3585 1365 -3565
rect 1385 -3585 1400 -3565
rect 1350 -3615 1400 -3585
rect 1350 -3635 1365 -3615
rect 1385 -3635 1400 -3615
rect 1350 -3650 1400 -3635
rect 1740 -3565 1790 -3550
rect 1740 -3585 1755 -3565
rect 1775 -3585 1790 -3565
rect 1740 -3615 1790 -3585
rect 1740 -3635 1755 -3615
rect 1775 -3635 1790 -3615
rect 1740 -3650 1790 -3635
rect 2080 -3565 2130 -3550
rect 2080 -3585 2095 -3565
rect 2115 -3585 2130 -3565
rect 2080 -3615 2130 -3585
rect 2080 -3635 2095 -3615
rect 2115 -3635 2130 -3615
rect 2080 -3650 2130 -3635
<< nsubdiff >>
rect -170 -2875 -130 -2860
rect -170 -2895 -160 -2875
rect -140 -2895 -130 -2875
rect -170 -2925 -130 -2895
rect -170 -2945 -160 -2925
rect -140 -2945 -130 -2925
rect -170 -2975 -130 -2945
rect -170 -2995 -160 -2975
rect -140 -2995 -130 -2975
rect -170 -3025 -130 -2995
rect -170 -3045 -160 -3025
rect -140 -3045 -130 -3025
rect -170 -3060 -130 -3045
rect 280 -2875 320 -2860
rect 280 -2895 290 -2875
rect 310 -2895 320 -2875
rect 280 -2925 320 -2895
rect 280 -2945 290 -2925
rect 310 -2945 320 -2925
rect 280 -2975 320 -2945
rect 280 -2995 290 -2975
rect 310 -2995 320 -2975
rect 280 -3025 320 -2995
rect 280 -3045 290 -3025
rect 310 -3045 320 -3025
rect 280 -3060 320 -3045
rect 730 -2875 770 -2860
rect 730 -2895 740 -2875
rect 760 -2895 770 -2875
rect 730 -2925 770 -2895
rect 730 -2945 740 -2925
rect 760 -2945 770 -2925
rect 730 -2975 770 -2945
rect 730 -2995 740 -2975
rect 760 -2995 770 -2975
rect 730 -3025 770 -2995
rect 730 -3045 740 -3025
rect 760 -3045 770 -3025
rect 730 -3060 770 -3045
rect 980 -2875 1020 -2860
rect 980 -2895 990 -2875
rect 1010 -2895 1020 -2875
rect 980 -2925 1020 -2895
rect 980 -2945 990 -2925
rect 1010 -2945 1020 -2925
rect 980 -2975 1020 -2945
rect 980 -2995 990 -2975
rect 1010 -2995 1020 -2975
rect 980 -3025 1020 -2995
rect 980 -3045 990 -3025
rect 1010 -3045 1020 -3025
rect 980 -3060 1020 -3045
rect 1145 -2875 1185 -2860
rect 1145 -2895 1155 -2875
rect 1175 -2895 1185 -2875
rect 1145 -2925 1185 -2895
rect 1145 -2945 1155 -2925
rect 1175 -2945 1185 -2925
rect 1145 -2975 1185 -2945
rect 1145 -2995 1155 -2975
rect 1175 -2995 1185 -2975
rect 1145 -3025 1185 -2995
rect 1145 -3045 1155 -3025
rect 1175 -3045 1185 -3025
rect 1145 -3060 1185 -3045
rect 1350 -2875 1400 -2860
rect 1350 -2895 1365 -2875
rect 1385 -2895 1400 -2875
rect 1350 -2925 1400 -2895
rect 1350 -2945 1365 -2925
rect 1385 -2945 1400 -2925
rect 1350 -2975 1400 -2945
rect 1350 -2995 1365 -2975
rect 1385 -2995 1400 -2975
rect 1350 -3025 1400 -2995
rect 1350 -3045 1365 -3025
rect 1385 -3045 1400 -3025
rect 1350 -3060 1400 -3045
rect 1545 -2875 1595 -2860
rect 1545 -2895 1560 -2875
rect 1580 -2895 1595 -2875
rect 1545 -2925 1595 -2895
rect 1545 -2945 1560 -2925
rect 1580 -2945 1595 -2925
rect 1545 -2975 1595 -2945
rect 1545 -2995 1560 -2975
rect 1580 -2995 1595 -2975
rect 1545 -3025 1595 -2995
rect 1545 -3045 1560 -3025
rect 1580 -3045 1595 -3025
rect 1545 -3060 1595 -3045
rect 1740 -2875 1790 -2860
rect 1740 -2895 1755 -2875
rect 1775 -2895 1790 -2875
rect 1740 -2925 1790 -2895
rect 1740 -2945 1755 -2925
rect 1775 -2945 1790 -2925
rect 1740 -2975 1790 -2945
rect 1740 -2995 1755 -2975
rect 1775 -2995 1790 -2975
rect 1740 -3025 1790 -2995
rect 1740 -3045 1755 -3025
rect 1775 -3045 1790 -3025
rect 1740 -3060 1790 -3045
rect 2080 -2875 2130 -2860
rect 2080 -2895 2095 -2875
rect 2115 -2895 2130 -2875
rect 2080 -2925 2130 -2895
rect 2080 -2945 2095 -2925
rect 2115 -2945 2130 -2925
rect 2080 -2975 2130 -2945
rect 2080 -2995 2095 -2975
rect 2115 -2995 2130 -2975
rect 2080 -3025 2130 -2995
rect 2080 -3045 2095 -3025
rect 2115 -3045 2130 -3025
rect 2080 -3060 2130 -3045
rect -170 -3255 -130 -3240
rect -170 -3275 -160 -3255
rect -140 -3275 -130 -3255
rect -170 -3305 -130 -3275
rect -170 -3325 -160 -3305
rect -140 -3325 -130 -3305
rect -170 -3355 -130 -3325
rect -170 -3375 -160 -3355
rect -140 -3375 -130 -3355
rect -170 -3405 -130 -3375
rect -170 -3425 -160 -3405
rect -140 -3425 -130 -3405
rect -170 -3440 -130 -3425
rect 280 -3255 320 -3240
rect 280 -3275 290 -3255
rect 310 -3275 320 -3255
rect 280 -3305 320 -3275
rect 280 -3325 290 -3305
rect 310 -3325 320 -3305
rect 280 -3355 320 -3325
rect 280 -3375 290 -3355
rect 310 -3375 320 -3355
rect 280 -3405 320 -3375
rect 280 -3425 290 -3405
rect 310 -3425 320 -3405
rect 280 -3440 320 -3425
rect 730 -3255 770 -3240
rect 730 -3275 740 -3255
rect 760 -3275 770 -3255
rect 730 -3305 770 -3275
rect 730 -3325 740 -3305
rect 760 -3325 770 -3305
rect 730 -3355 770 -3325
rect 730 -3375 740 -3355
rect 760 -3375 770 -3355
rect 730 -3405 770 -3375
rect 730 -3425 740 -3405
rect 760 -3425 770 -3405
rect 730 -3440 770 -3425
rect 930 -3255 970 -3240
rect 930 -3275 940 -3255
rect 960 -3275 970 -3255
rect 930 -3305 970 -3275
rect 930 -3325 940 -3305
rect 960 -3325 970 -3305
rect 930 -3355 970 -3325
rect 930 -3375 940 -3355
rect 960 -3375 970 -3355
rect 930 -3405 970 -3375
rect 930 -3425 940 -3405
rect 960 -3425 970 -3405
rect 930 -3440 970 -3425
rect 1095 -3255 1135 -3240
rect 1095 -3275 1105 -3255
rect 1125 -3275 1135 -3255
rect 1095 -3305 1135 -3275
rect 1095 -3325 1105 -3305
rect 1125 -3325 1135 -3305
rect 1095 -3355 1135 -3325
rect 1095 -3375 1105 -3355
rect 1125 -3375 1135 -3355
rect 1095 -3405 1135 -3375
rect 1095 -3425 1105 -3405
rect 1125 -3425 1135 -3405
rect 1095 -3440 1135 -3425
rect 1260 -3255 1300 -3240
rect 1260 -3275 1270 -3255
rect 1290 -3275 1300 -3255
rect 1260 -3305 1300 -3275
rect 1260 -3325 1270 -3305
rect 1290 -3325 1300 -3305
rect 1260 -3355 1300 -3325
rect 1260 -3375 1270 -3355
rect 1290 -3375 1300 -3355
rect 1260 -3405 1300 -3375
rect 1260 -3425 1270 -3405
rect 1290 -3425 1300 -3405
rect 1260 -3440 1300 -3425
rect 1350 -3255 1400 -3240
rect 1350 -3275 1365 -3255
rect 1385 -3275 1400 -3255
rect 1350 -3305 1400 -3275
rect 1350 -3325 1365 -3305
rect 1385 -3325 1400 -3305
rect 1350 -3355 1400 -3325
rect 1350 -3375 1365 -3355
rect 1385 -3375 1400 -3355
rect 1350 -3405 1400 -3375
rect 1350 -3425 1365 -3405
rect 1385 -3425 1400 -3405
rect 1350 -3440 1400 -3425
rect 1740 -3255 1790 -3240
rect 1740 -3275 1755 -3255
rect 1775 -3275 1790 -3255
rect 1740 -3305 1790 -3275
rect 1740 -3325 1755 -3305
rect 1775 -3325 1790 -3305
rect 1740 -3355 1790 -3325
rect 1740 -3375 1755 -3355
rect 1775 -3375 1790 -3355
rect 1740 -3405 1790 -3375
rect 1740 -3425 1755 -3405
rect 1775 -3425 1790 -3405
rect 1740 -3440 1790 -3425
<< psubdiffcont >>
rect -160 -2685 -140 -2665
rect -160 -2735 -140 -2715
rect 290 -2685 310 -2665
rect 290 -2735 310 -2715
rect 740 -2685 760 -2665
rect 740 -2735 760 -2715
rect 990 -2685 1010 -2665
rect 990 -2735 1010 -2715
rect 1155 -2685 1175 -2665
rect 1155 -2735 1175 -2715
rect 1370 -2685 1390 -2665
rect 1370 -2735 1390 -2715
rect 1565 -2685 1585 -2665
rect 1565 -2735 1585 -2715
rect 1760 -2685 1780 -2665
rect 1760 -2735 1780 -2715
rect -160 -3585 -140 -3565
rect -160 -3635 -140 -3615
rect 290 -3585 310 -3565
rect 290 -3635 310 -3615
rect 740 -3585 760 -3565
rect 740 -3635 760 -3615
rect 940 -3585 960 -3565
rect 940 -3635 960 -3615
rect 1105 -3585 1125 -3565
rect 1105 -3635 1125 -3615
rect 1270 -3585 1290 -3565
rect 1270 -3635 1290 -3615
rect 1365 -3585 1385 -3565
rect 1365 -3635 1385 -3615
rect 1755 -3585 1775 -3565
rect 1755 -3635 1775 -3615
rect 2095 -3585 2115 -3565
rect 2095 -3635 2115 -3615
<< nsubdiffcont >>
rect -160 -2895 -140 -2875
rect -160 -2945 -140 -2925
rect -160 -2995 -140 -2975
rect -160 -3045 -140 -3025
rect 290 -2895 310 -2875
rect 290 -2945 310 -2925
rect 290 -2995 310 -2975
rect 290 -3045 310 -3025
rect 740 -2895 760 -2875
rect 740 -2945 760 -2925
rect 740 -2995 760 -2975
rect 740 -3045 760 -3025
rect 990 -2895 1010 -2875
rect 990 -2945 1010 -2925
rect 990 -2995 1010 -2975
rect 990 -3045 1010 -3025
rect 1155 -2895 1175 -2875
rect 1155 -2945 1175 -2925
rect 1155 -2995 1175 -2975
rect 1155 -3045 1175 -3025
rect 1365 -2895 1385 -2875
rect 1365 -2945 1385 -2925
rect 1365 -2995 1385 -2975
rect 1365 -3045 1385 -3025
rect 1560 -2895 1580 -2875
rect 1560 -2945 1580 -2925
rect 1560 -2995 1580 -2975
rect 1560 -3045 1580 -3025
rect 1755 -2895 1775 -2875
rect 1755 -2945 1775 -2925
rect 1755 -2995 1775 -2975
rect 1755 -3045 1775 -3025
rect 2095 -2895 2115 -2875
rect 2095 -2945 2115 -2925
rect 2095 -2995 2115 -2975
rect 2095 -3045 2115 -3025
rect -160 -3275 -140 -3255
rect -160 -3325 -140 -3305
rect -160 -3375 -140 -3355
rect -160 -3425 -140 -3405
rect 290 -3275 310 -3255
rect 290 -3325 310 -3305
rect 290 -3375 310 -3355
rect 290 -3425 310 -3405
rect 740 -3275 760 -3255
rect 740 -3325 760 -3305
rect 740 -3375 760 -3355
rect 740 -3425 760 -3405
rect 940 -3275 960 -3255
rect 940 -3325 960 -3305
rect 940 -3375 960 -3355
rect 940 -3425 960 -3405
rect 1105 -3275 1125 -3255
rect 1105 -3325 1125 -3305
rect 1105 -3375 1125 -3355
rect 1105 -3425 1125 -3405
rect 1270 -3275 1290 -3255
rect 1270 -3325 1290 -3305
rect 1270 -3375 1290 -3355
rect 1270 -3425 1290 -3405
rect 1365 -3275 1385 -3255
rect 1365 -3325 1385 -3305
rect 1365 -3375 1385 -3355
rect 1365 -3425 1385 -3405
rect 1755 -3275 1775 -3255
rect 1755 -3325 1775 -3305
rect 1755 -3375 1775 -3355
rect 1755 -3425 1775 -3405
<< poly >>
rect 170 -2610 375 -2595
rect -90 -2650 -75 -2635
rect -35 -2650 -20 -2635
rect 170 -2650 185 -2610
rect 225 -2650 240 -2635
rect 360 -2650 375 -2610
rect 895 -2605 935 -2595
rect 895 -2625 905 -2605
rect 925 -2625 935 -2605
rect 895 -2635 935 -2625
rect 415 -2650 430 -2635
rect 620 -2650 635 -2635
rect 675 -2650 690 -2635
rect 840 -2650 855 -2635
rect 895 -2650 910 -2635
rect 1060 -2650 1075 -2635
rect 1225 -2650 1240 -2635
rect 1450 -2650 1465 -2635
rect 1645 -2650 1660 -2635
rect 1840 -2650 1855 -2635
rect 1985 -2650 2000 -2635
rect -90 -2785 -75 -2750
rect -150 -2800 -75 -2785
rect -90 -2860 -75 -2800
rect -35 -2765 -20 -2750
rect -35 -2775 15 -2765
rect 170 -2770 185 -2750
rect -35 -2795 -15 -2775
rect 5 -2795 15 -2775
rect -35 -2805 15 -2795
rect 60 -2785 185 -2770
rect -35 -2860 -20 -2805
rect 60 -3015 75 -2785
rect 170 -2860 185 -2785
rect 225 -2805 240 -2750
rect 225 -2815 275 -2805
rect 225 -2835 245 -2815
rect 265 -2835 275 -2815
rect 225 -2845 275 -2835
rect 225 -2860 240 -2845
rect 360 -2860 375 -2750
rect 415 -2765 430 -2750
rect 415 -2775 465 -2765
rect 620 -2770 635 -2750
rect 415 -2795 435 -2775
rect 455 -2795 465 -2775
rect 415 -2805 465 -2795
rect 510 -2785 635 -2770
rect 415 -2860 430 -2805
rect 35 -3025 75 -3015
rect 35 -3045 45 -3025
rect 65 -3045 75 -3025
rect 35 -3055 75 -3045
rect 510 -3015 525 -2785
rect 620 -2860 635 -2785
rect 675 -2770 690 -2750
rect 675 -2780 760 -2770
rect 675 -2785 730 -2780
rect 675 -2860 690 -2785
rect 720 -2800 730 -2785
rect 750 -2800 760 -2780
rect 720 -2810 760 -2800
rect 840 -2860 855 -2750
rect 895 -2860 910 -2750
rect 935 -2800 975 -2790
rect 1060 -2800 1075 -2750
rect 935 -2820 945 -2800
rect 965 -2815 1075 -2800
rect 965 -2820 975 -2815
rect 935 -2830 975 -2820
rect 1060 -2860 1075 -2815
rect 1100 -2800 1140 -2790
rect 1225 -2800 1240 -2750
rect 1335 -2785 1375 -2775
rect 1100 -2820 1110 -2800
rect 1130 -2815 1240 -2800
rect 1130 -2820 1140 -2815
rect 1100 -2830 1140 -2820
rect 1225 -2860 1240 -2815
rect 1265 -2800 1305 -2790
rect 1265 -2820 1275 -2800
rect 1295 -2820 1305 -2800
rect 1335 -2805 1345 -2785
rect 1365 -2800 1375 -2785
rect 1450 -2800 1465 -2750
rect 1645 -2790 1660 -2750
rect 1840 -2765 1855 -2750
rect 1985 -2765 2000 -2750
rect 1365 -2805 1465 -2800
rect 1335 -2815 1465 -2805
rect 1265 -2830 1305 -2820
rect 1450 -2860 1465 -2815
rect 1620 -2800 1660 -2790
rect 1620 -2820 1630 -2800
rect 1650 -2820 1660 -2800
rect 1815 -2775 2195 -2765
rect 1815 -2795 1825 -2775
rect 1845 -2780 2195 -2775
rect 1845 -2795 1855 -2780
rect 1815 -2805 1855 -2795
rect 1620 -2830 1660 -2820
rect 1645 -2860 1660 -2830
rect 1840 -2860 1855 -2805
rect 1880 -2815 1920 -2805
rect 1880 -2835 1890 -2815
rect 1910 -2830 1920 -2815
rect 1910 -2835 2000 -2830
rect 1880 -2845 2000 -2835
rect 1985 -2860 2000 -2845
rect 2180 -2860 2195 -2780
rect 485 -3025 525 -3015
rect 485 -3045 495 -3025
rect 515 -3045 525 -3025
rect 485 -3055 525 -3045
rect -90 -3075 -75 -3060
rect -35 -3075 -20 -3060
rect 170 -3075 185 -3060
rect 225 -3075 240 -3060
rect 360 -3075 375 -3060
rect 415 -3075 430 -3060
rect 620 -3075 635 -3060
rect 675 -3075 690 -3060
rect 840 -3075 855 -3060
rect 895 -3075 910 -3060
rect 1060 -3075 1075 -3060
rect 1225 -3075 1240 -3060
rect 1450 -3075 1465 -3060
rect 1645 -3075 1660 -3060
rect 1840 -3075 1855 -3060
rect 1985 -3075 2000 -3060
rect 2180 -3075 2195 -3060
rect 810 -3085 855 -3075
rect 810 -3105 820 -3085
rect 840 -3105 855 -3085
rect 810 -3115 855 -3105
rect 1620 -3195 1660 -3185
rect 1620 -3215 1630 -3195
rect 1650 -3215 1660 -3195
rect 1620 -3225 1660 -3215
rect -90 -3240 -75 -3225
rect -35 -3240 -20 -3225
rect 170 -3240 185 -3225
rect 225 -3240 240 -3225
rect 360 -3240 375 -3225
rect 415 -3240 430 -3225
rect 620 -3240 635 -3225
rect 675 -3240 690 -3225
rect 875 -3240 890 -3225
rect 1040 -3240 1055 -3225
rect 1205 -3240 1220 -3225
rect 1450 -3240 1465 -3225
rect 1645 -3240 1660 -3225
rect 1840 -3240 1855 -3225
rect 1985 -3240 2000 -3225
rect 35 -3255 75 -3245
rect 35 -3275 45 -3255
rect 65 -3275 75 -3255
rect 35 -3285 75 -3275
rect -90 -3500 -75 -3440
rect -150 -3515 -75 -3500
rect -90 -3550 -75 -3515
rect -35 -3495 -20 -3440
rect -35 -3505 15 -3495
rect -35 -3525 -15 -3505
rect 5 -3525 15 -3505
rect -35 -3535 15 -3525
rect 60 -3515 75 -3285
rect 485 -3255 525 -3245
rect 485 -3275 495 -3255
rect 515 -3275 525 -3255
rect 485 -3285 525 -3275
rect 170 -3515 185 -3440
rect 60 -3530 185 -3515
rect -35 -3550 -20 -3535
rect 170 -3550 185 -3530
rect 225 -3455 240 -3440
rect 225 -3465 275 -3455
rect 225 -3485 245 -3465
rect 265 -3485 275 -3465
rect 225 -3495 275 -3485
rect 225 -3550 240 -3495
rect 360 -3550 375 -3440
rect 415 -3495 430 -3440
rect 415 -3505 465 -3495
rect 415 -3525 435 -3505
rect 455 -3525 465 -3505
rect 415 -3535 465 -3525
rect 510 -3515 525 -3285
rect 620 -3515 635 -3440
rect 510 -3530 635 -3515
rect 415 -3550 430 -3535
rect 620 -3550 635 -3530
rect 675 -3470 690 -3440
rect 675 -3480 850 -3470
rect 675 -3485 740 -3480
rect 675 -3550 690 -3485
rect 730 -3500 740 -3485
rect 760 -3485 820 -3480
rect 760 -3500 770 -3485
rect 730 -3510 770 -3500
rect 810 -3500 820 -3485
rect 840 -3500 850 -3480
rect 810 -3510 850 -3500
rect 875 -3485 890 -3440
rect 975 -3480 1015 -3470
rect 975 -3485 985 -3480
rect 875 -3500 985 -3485
rect 1005 -3500 1015 -3480
rect 875 -3550 890 -3500
rect 975 -3510 1015 -3500
rect 1040 -3485 1055 -3440
rect 1140 -3480 1180 -3470
rect 1140 -3485 1150 -3480
rect 1040 -3500 1150 -3485
rect 1170 -3500 1180 -3480
rect 1040 -3550 1055 -3500
rect 1140 -3510 1180 -3500
rect 1205 -3485 1220 -3440
rect 1270 -3480 1310 -3470
rect 1270 -3485 1280 -3480
rect 1205 -3500 1280 -3485
rect 1300 -3500 1310 -3480
rect 1205 -3550 1220 -3500
rect 1270 -3510 1310 -3500
rect 1335 -3485 1375 -3475
rect 1335 -3505 1345 -3485
rect 1365 -3500 1375 -3485
rect 1450 -3500 1465 -3440
rect 1645 -3455 1660 -3440
rect 1685 -3465 1725 -3455
rect 1840 -3465 1855 -3440
rect 1985 -3465 2000 -3440
rect 1685 -3485 1695 -3465
rect 1715 -3480 2195 -3465
rect 1715 -3485 1725 -3480
rect 1685 -3495 1725 -3485
rect 1365 -3505 1465 -3500
rect 1335 -3515 1465 -3505
rect 1450 -3550 1465 -3515
rect 1645 -3550 1660 -3535
rect 1840 -3550 1855 -3480
rect 1880 -3510 1920 -3505
rect 1880 -3530 1890 -3510
rect 1910 -3525 1920 -3510
rect 1910 -3530 2000 -3525
rect 1880 -3540 2000 -3530
rect 1985 -3550 2000 -3540
rect 2180 -3550 2195 -3480
rect -90 -3665 -75 -3650
rect -35 -3665 -20 -3650
rect 170 -3690 185 -3650
rect 225 -3665 240 -3650
rect 360 -3690 375 -3650
rect 415 -3665 430 -3650
rect 620 -3665 635 -3650
rect 675 -3665 690 -3650
rect 875 -3665 890 -3650
rect 1040 -3665 1055 -3650
rect 1205 -3665 1220 -3650
rect 1450 -3665 1465 -3650
rect 1645 -3665 1660 -3650
rect 1840 -3665 1855 -3650
rect 1985 -3665 2000 -3650
rect 2180 -3665 2195 -3650
rect 170 -3705 375 -3690
rect 1645 -3675 1700 -3665
rect 1645 -3695 1670 -3675
rect 1690 -3695 1700 -3675
rect 1645 -3705 1700 -3695
<< polycont >>
rect 905 -2625 925 -2605
rect -15 -2795 5 -2775
rect 245 -2835 265 -2815
rect 435 -2795 455 -2775
rect 45 -3045 65 -3025
rect 730 -2800 750 -2780
rect 945 -2820 965 -2800
rect 1110 -2820 1130 -2800
rect 1275 -2820 1295 -2800
rect 1345 -2805 1365 -2785
rect 1630 -2820 1650 -2800
rect 1825 -2795 1845 -2775
rect 1890 -2835 1910 -2815
rect 495 -3045 515 -3025
rect 820 -3105 840 -3085
rect 1630 -3215 1650 -3195
rect 45 -3275 65 -3255
rect -15 -3525 5 -3505
rect 495 -3275 515 -3255
rect 245 -3485 265 -3465
rect 435 -3525 455 -3505
rect 740 -3500 760 -3480
rect 820 -3500 840 -3480
rect 985 -3500 1005 -3480
rect 1150 -3500 1170 -3480
rect 1280 -3500 1300 -3480
rect 1345 -3505 1365 -3485
rect 1695 -3485 1715 -3465
rect 1890 -3530 1910 -3510
rect 1670 -3695 1690 -3675
<< locali >>
rect -340 -2550 -290 -2540
rect -340 -2555 -260 -2550
rect -340 -2575 -325 -2555
rect -305 -2570 -260 -2555
rect -240 -2570 -210 -2550
rect -190 -2570 -160 -2550
rect -140 -2570 -110 -2550
rect -90 -2570 -60 -2550
rect -40 -2570 -10 -2550
rect 10 -2570 40 -2550
rect 60 -2570 90 -2550
rect 110 -2570 140 -2550
rect 160 -2570 190 -2550
rect 210 -2570 240 -2550
rect 260 -2570 290 -2550
rect 310 -2570 340 -2550
rect 360 -2570 390 -2550
rect 410 -2570 440 -2550
rect 460 -2570 490 -2550
rect 510 -2570 540 -2550
rect 560 -2570 590 -2550
rect 610 -2570 640 -2550
rect 660 -2570 690 -2550
rect 710 -2570 740 -2550
rect 760 -2570 790 -2550
rect 810 -2570 840 -2550
rect 860 -2570 890 -2550
rect 910 -2570 940 -2550
rect 960 -2570 990 -2550
rect 1010 -2570 1040 -2550
rect 1060 -2570 1090 -2550
rect 1110 -2570 1140 -2550
rect 1160 -2570 1190 -2550
rect 1210 -2570 1240 -2550
rect 1260 -2570 1290 -2550
rect 1310 -2570 1340 -2550
rect 1360 -2570 1390 -2550
rect 1410 -2570 1440 -2550
rect 1460 -2570 1490 -2550
rect 1510 -2570 1540 -2550
rect 1560 -2570 1590 -2550
rect 1610 -2570 1640 -2550
rect 1660 -2570 1690 -2550
rect 1710 -2570 1740 -2550
rect 1760 -2570 1790 -2550
rect 1810 -2570 1840 -2550
rect 1860 -2570 1890 -2550
rect 1910 -2570 1940 -2550
rect 1960 -2570 1990 -2550
rect 2010 -2570 2040 -2550
rect 2060 -2570 2090 -2550
rect 2110 -2570 2140 -2550
rect 2160 -2570 2190 -2550
rect 2210 -2570 2240 -2550
rect 2260 -2570 2305 -2550
rect -305 -2575 -290 -2570
rect -340 -2590 -290 -2575
rect -120 -2655 -100 -2570
rect -10 -2655 10 -2570
rect 75 -2605 115 -2595
rect 75 -2625 85 -2605
rect 105 -2625 115 -2605
rect 75 -2635 115 -2625
rect -165 -2665 -95 -2655
rect -165 -2685 -160 -2665
rect -140 -2685 -120 -2665
rect -100 -2685 -95 -2665
rect -165 -2715 -95 -2685
rect -165 -2735 -160 -2715
rect -140 -2735 -120 -2715
rect -100 -2735 -95 -2715
rect -165 -2745 -95 -2735
rect -70 -2665 -40 -2655
rect -70 -2685 -65 -2665
rect -45 -2685 -40 -2665
rect -70 -2715 -40 -2685
rect -70 -2735 -65 -2715
rect -45 -2735 -40 -2715
rect -70 -2745 -40 -2735
rect -15 -2665 15 -2655
rect -15 -2685 -10 -2665
rect 10 -2685 15 -2665
rect -15 -2715 15 -2685
rect -15 -2735 -10 -2715
rect 10 -2735 15 -2715
rect -15 -2745 15 -2735
rect -70 -2825 -50 -2745
rect -25 -2775 15 -2765
rect -25 -2795 -15 -2775
rect 5 -2785 15 -2775
rect 95 -2785 115 -2635
rect 140 -2655 160 -2570
rect 250 -2655 270 -2570
rect 330 -2655 350 -2570
rect 440 -2655 460 -2570
rect 590 -2655 610 -2570
rect 700 -2655 720 -2570
rect 810 -2655 830 -2570
rect 895 -2605 935 -2595
rect 895 -2625 905 -2605
rect 925 -2625 935 -2605
rect 895 -2635 935 -2625
rect 1195 -2655 1215 -2570
rect 1415 -2655 1435 -2570
rect 1610 -2655 1630 -2570
rect 1805 -2655 1825 -2570
rect 135 -2665 165 -2655
rect 135 -2685 140 -2665
rect 160 -2685 165 -2665
rect 135 -2715 165 -2685
rect 135 -2735 140 -2715
rect 160 -2735 165 -2715
rect 135 -2745 165 -2735
rect 190 -2665 220 -2655
rect 190 -2685 195 -2665
rect 215 -2685 220 -2665
rect 190 -2715 220 -2685
rect 190 -2735 195 -2715
rect 215 -2735 220 -2715
rect 190 -2745 220 -2735
rect 245 -2665 355 -2655
rect 245 -2685 250 -2665
rect 270 -2685 290 -2665
rect 310 -2685 330 -2665
rect 350 -2685 355 -2665
rect 245 -2715 355 -2685
rect 245 -2735 250 -2715
rect 270 -2735 290 -2715
rect 310 -2735 330 -2715
rect 350 -2735 355 -2715
rect 245 -2745 355 -2735
rect 380 -2665 410 -2655
rect 380 -2685 385 -2665
rect 405 -2685 410 -2665
rect 380 -2715 410 -2685
rect 380 -2735 385 -2715
rect 405 -2735 410 -2715
rect 380 -2745 410 -2735
rect 435 -2665 465 -2655
rect 435 -2685 440 -2665
rect 460 -2685 465 -2665
rect 435 -2715 465 -2685
rect 435 -2735 440 -2715
rect 460 -2735 465 -2715
rect 435 -2745 465 -2735
rect 585 -2665 615 -2655
rect 585 -2685 590 -2665
rect 610 -2685 615 -2665
rect 585 -2715 615 -2685
rect 585 -2735 590 -2715
rect 610 -2735 615 -2715
rect 585 -2745 615 -2735
rect 640 -2665 670 -2655
rect 640 -2685 645 -2665
rect 665 -2685 670 -2665
rect 640 -2715 670 -2685
rect 640 -2735 645 -2715
rect 665 -2735 670 -2715
rect 640 -2745 670 -2735
rect 695 -2665 765 -2655
rect 695 -2685 700 -2665
rect 720 -2685 740 -2665
rect 760 -2685 765 -2665
rect 695 -2715 765 -2685
rect 695 -2735 700 -2715
rect 720 -2735 740 -2715
rect 760 -2735 765 -2715
rect 695 -2745 765 -2735
rect 805 -2665 835 -2655
rect 805 -2685 810 -2665
rect 830 -2685 835 -2665
rect 805 -2715 835 -2685
rect 805 -2735 810 -2715
rect 830 -2735 835 -2715
rect 805 -2745 835 -2735
rect 860 -2665 890 -2655
rect 860 -2685 865 -2665
rect 885 -2685 890 -2665
rect 860 -2715 890 -2685
rect 860 -2735 865 -2715
rect 885 -2735 890 -2715
rect 860 -2745 890 -2735
rect 915 -2665 945 -2655
rect 915 -2685 920 -2665
rect 940 -2685 945 -2665
rect 915 -2715 945 -2685
rect 915 -2735 920 -2715
rect 940 -2735 945 -2715
rect 915 -2745 945 -2735
rect 985 -2665 1055 -2655
rect 985 -2685 990 -2665
rect 1010 -2685 1030 -2665
rect 1050 -2685 1055 -2665
rect 985 -2715 1055 -2685
rect 985 -2735 990 -2715
rect 1010 -2735 1030 -2715
rect 1050 -2735 1055 -2715
rect 985 -2745 1055 -2735
rect 1080 -2665 1110 -2655
rect 1080 -2685 1085 -2665
rect 1105 -2685 1110 -2665
rect 1080 -2715 1110 -2685
rect 1080 -2735 1085 -2715
rect 1105 -2735 1110 -2715
rect 1080 -2745 1110 -2735
rect 1150 -2665 1220 -2655
rect 1150 -2685 1155 -2665
rect 1175 -2685 1195 -2665
rect 1215 -2685 1220 -2665
rect 1150 -2715 1220 -2685
rect 1150 -2735 1155 -2715
rect 1175 -2735 1195 -2715
rect 1215 -2735 1220 -2715
rect 1150 -2745 1220 -2735
rect 1245 -2665 1275 -2655
rect 1245 -2685 1250 -2665
rect 1270 -2685 1275 -2665
rect 1245 -2715 1275 -2685
rect 1245 -2735 1250 -2715
rect 1270 -2735 1275 -2715
rect 1245 -2745 1275 -2735
rect 1365 -2665 1445 -2655
rect 1365 -2685 1370 -2665
rect 1390 -2685 1415 -2665
rect 1435 -2685 1445 -2665
rect 1365 -2715 1445 -2685
rect 1365 -2735 1370 -2715
rect 1390 -2735 1415 -2715
rect 1435 -2735 1445 -2715
rect 1365 -2745 1445 -2735
rect 1470 -2665 1510 -2655
rect 1470 -2685 1480 -2665
rect 1500 -2685 1510 -2665
rect 1470 -2715 1510 -2685
rect 1470 -2735 1480 -2715
rect 1500 -2735 1510 -2715
rect 1470 -2745 1510 -2735
rect 1560 -2665 1640 -2655
rect 1560 -2685 1565 -2665
rect 1585 -2685 1610 -2665
rect 1630 -2685 1640 -2665
rect 1560 -2715 1640 -2685
rect 1560 -2735 1565 -2715
rect 1585 -2735 1610 -2715
rect 1630 -2735 1640 -2715
rect 1560 -2745 1640 -2735
rect 1665 -2665 1705 -2655
rect 1665 -2685 1675 -2665
rect 1695 -2685 1705 -2665
rect 1665 -2715 1705 -2685
rect 1665 -2735 1675 -2715
rect 1695 -2735 1705 -2715
rect 1665 -2745 1705 -2735
rect 1755 -2665 1835 -2655
rect 1755 -2685 1760 -2665
rect 1780 -2685 1805 -2665
rect 1825 -2685 1835 -2665
rect 1755 -2715 1835 -2685
rect 1755 -2735 1760 -2715
rect 1780 -2735 1805 -2715
rect 1825 -2735 1835 -2715
rect 1755 -2745 1835 -2735
rect 1860 -2665 1900 -2655
rect 1860 -2685 1870 -2665
rect 1890 -2685 1900 -2665
rect 1860 -2715 1900 -2685
rect 1860 -2735 1870 -2715
rect 1890 -2735 1900 -2715
rect 1860 -2745 1900 -2735
rect 1940 -2665 1980 -2655
rect 1940 -2685 1950 -2665
rect 1970 -2685 1980 -2665
rect 1940 -2715 1980 -2685
rect 1940 -2735 1950 -2715
rect 1970 -2735 1980 -2715
rect 1940 -2745 1980 -2735
rect 2005 -2665 2045 -2655
rect 2005 -2685 2015 -2665
rect 2035 -2685 2045 -2665
rect 2005 -2715 2045 -2685
rect 2005 -2735 2015 -2715
rect 2035 -2735 2045 -2715
rect 2005 -2745 2045 -2735
rect 5 -2795 115 -2785
rect -25 -2805 115 -2795
rect -70 -2845 10 -2825
rect -10 -2865 10 -2845
rect -165 -2875 -95 -2865
rect -165 -2895 -160 -2875
rect -140 -2895 -120 -2875
rect -100 -2895 -95 -2875
rect -165 -2925 -95 -2895
rect -165 -2945 -160 -2925
rect -140 -2945 -120 -2925
rect -100 -2945 -95 -2925
rect -165 -2975 -95 -2945
rect -165 -2995 -160 -2975
rect -140 -2995 -120 -2975
rect -100 -2995 -95 -2975
rect -165 -3025 -95 -2995
rect -165 -3045 -160 -3025
rect -140 -3045 -120 -3025
rect -100 -3045 -95 -3025
rect -165 -3055 -95 -3045
rect -70 -2875 -40 -2865
rect -70 -2895 -65 -2875
rect -45 -2895 -40 -2875
rect -70 -2925 -40 -2895
rect -70 -2945 -65 -2925
rect -45 -2945 -40 -2925
rect -70 -2975 -40 -2945
rect -70 -2995 -65 -2975
rect -45 -2995 -40 -2975
rect -70 -3025 -40 -2995
rect -70 -3045 -65 -3025
rect -45 -3045 -40 -3025
rect -70 -3055 -40 -3045
rect -15 -2875 15 -2865
rect -15 -2895 -10 -2875
rect 10 -2895 15 -2875
rect -15 -2925 15 -2895
rect -15 -2945 -10 -2925
rect 10 -2945 15 -2925
rect -15 -2975 15 -2945
rect -15 -2995 -10 -2975
rect 10 -2995 15 -2975
rect -15 -3025 15 -2995
rect -15 -3045 -10 -3025
rect 10 -3030 15 -3025
rect 35 -3025 75 -3015
rect 35 -3030 45 -3025
rect 10 -3045 45 -3030
rect 65 -3045 75 -3025
rect -15 -3055 75 -3045
rect 95 -3035 115 -2805
rect 195 -2825 215 -2745
rect 140 -2845 215 -2825
rect 235 -2815 275 -2805
rect 235 -2835 245 -2815
rect 265 -2825 275 -2815
rect 380 -2825 400 -2745
rect 425 -2775 465 -2765
rect 425 -2795 435 -2775
rect 455 -2785 465 -2775
rect 455 -2795 565 -2785
rect 425 -2805 565 -2795
rect 265 -2835 460 -2825
rect 235 -2845 460 -2835
rect 140 -2865 160 -2845
rect 440 -2865 460 -2845
rect 135 -2875 165 -2865
rect 135 -2895 140 -2875
rect 160 -2895 165 -2875
rect 135 -2925 165 -2895
rect 135 -2945 140 -2925
rect 160 -2945 165 -2925
rect 135 -2975 165 -2945
rect 135 -2995 140 -2975
rect 160 -2995 165 -2975
rect 135 -3025 165 -2995
rect 135 -3035 140 -3025
rect 95 -3045 140 -3035
rect 160 -3045 165 -3025
rect 95 -3055 165 -3045
rect 190 -2875 220 -2865
rect 190 -2895 195 -2875
rect 215 -2895 220 -2875
rect 190 -2925 220 -2895
rect 190 -2945 195 -2925
rect 215 -2945 220 -2925
rect 190 -2975 220 -2945
rect 190 -2995 195 -2975
rect 215 -2995 220 -2975
rect 190 -3025 220 -2995
rect 190 -3045 195 -3025
rect 215 -3045 220 -3025
rect 190 -3055 220 -3045
rect 245 -2875 355 -2865
rect 245 -2895 250 -2875
rect 270 -2895 290 -2875
rect 310 -2895 330 -2875
rect 350 -2895 355 -2875
rect 245 -2925 355 -2895
rect 245 -2945 250 -2925
rect 270 -2945 290 -2925
rect 310 -2945 330 -2925
rect 350 -2945 355 -2925
rect 245 -2975 355 -2945
rect 245 -2995 250 -2975
rect 270 -2995 290 -2975
rect 310 -2995 330 -2975
rect 350 -2995 355 -2975
rect 245 -3025 355 -2995
rect 245 -3045 250 -3025
rect 270 -3045 290 -3025
rect 310 -3045 330 -3025
rect 350 -3045 355 -3025
rect 245 -3055 355 -3045
rect 380 -2875 410 -2865
rect 380 -2895 385 -2875
rect 405 -2895 410 -2875
rect 380 -2925 410 -2895
rect 380 -2945 385 -2925
rect 405 -2945 410 -2925
rect 380 -2975 410 -2945
rect 380 -2995 385 -2975
rect 405 -2995 410 -2975
rect 380 -3025 410 -2995
rect 380 -3045 385 -3025
rect 405 -3045 410 -3025
rect 380 -3055 410 -3045
rect 435 -2875 465 -2865
rect 435 -2895 440 -2875
rect 460 -2895 465 -2875
rect 435 -2925 465 -2895
rect 435 -2945 440 -2925
rect 460 -2945 465 -2925
rect 435 -2975 465 -2945
rect 435 -2995 440 -2975
rect 460 -2995 465 -2975
rect 435 -3025 465 -2995
rect 435 -3045 440 -3025
rect 460 -3030 465 -3025
rect 485 -3025 525 -3015
rect 485 -3030 495 -3025
rect 460 -3045 495 -3030
rect 515 -3045 525 -3025
rect 435 -3055 525 -3045
rect 545 -3035 565 -2805
rect 645 -2825 665 -2745
rect 720 -2780 760 -2770
rect 720 -2800 730 -2780
rect 750 -2800 760 -2780
rect 720 -2810 760 -2800
rect 920 -2790 940 -2745
rect 1090 -2790 1110 -2745
rect 1255 -2790 1275 -2745
rect 1335 -2785 1375 -2775
rect 920 -2800 975 -2790
rect 920 -2820 945 -2800
rect 965 -2820 975 -2800
rect 920 -2825 975 -2820
rect 590 -2845 665 -2825
rect 810 -2830 975 -2825
rect 1090 -2800 1140 -2790
rect 1090 -2820 1110 -2800
rect 1130 -2820 1140 -2800
rect 1090 -2830 1140 -2820
rect 1255 -2800 1305 -2790
rect 1255 -2820 1275 -2800
rect 1295 -2820 1305 -2800
rect 1335 -2805 1345 -2785
rect 1365 -2805 1375 -2785
rect 1335 -2815 1375 -2805
rect 1490 -2800 1510 -2745
rect 1685 -2785 1705 -2745
rect 1815 -2775 1855 -2765
rect 1815 -2785 1825 -2775
rect 1620 -2800 1660 -2790
rect 1255 -2830 1305 -2820
rect 1490 -2820 1630 -2800
rect 1650 -2820 1660 -2800
rect 810 -2845 940 -2830
rect 590 -2865 610 -2845
rect 810 -2865 830 -2845
rect 920 -2865 940 -2845
rect 1090 -2865 1110 -2830
rect 1255 -2865 1275 -2830
rect 1490 -2865 1510 -2820
rect 1620 -2830 1660 -2820
rect 1685 -2795 1825 -2785
rect 1845 -2795 1855 -2775
rect 1685 -2805 1855 -2795
rect 1880 -2805 1900 -2745
rect 1685 -2865 1705 -2805
rect 1880 -2815 1920 -2805
rect 1880 -2835 1890 -2815
rect 1910 -2835 1920 -2815
rect 1880 -2845 1920 -2835
rect 1880 -2865 1900 -2845
rect 1950 -2865 1970 -2745
rect 2015 -2800 2035 -2745
rect 2015 -2820 2325 -2800
rect 2015 -2865 2035 -2820
rect 2210 -2865 2230 -2820
rect 585 -2875 615 -2865
rect 585 -2895 590 -2875
rect 610 -2895 615 -2875
rect 585 -2925 615 -2895
rect 585 -2945 590 -2925
rect 610 -2945 615 -2925
rect 585 -2975 615 -2945
rect 585 -2995 590 -2975
rect 610 -2995 615 -2975
rect 585 -3025 615 -2995
rect 585 -3035 590 -3025
rect 545 -3045 590 -3035
rect 610 -3045 615 -3025
rect 545 -3055 615 -3045
rect 640 -2875 670 -2865
rect 640 -2895 645 -2875
rect 665 -2895 670 -2875
rect 640 -2925 670 -2895
rect 640 -2945 645 -2925
rect 665 -2945 670 -2925
rect 640 -2975 670 -2945
rect 640 -2995 645 -2975
rect 665 -2995 670 -2975
rect 640 -3025 670 -2995
rect 640 -3045 645 -3025
rect 665 -3045 670 -3025
rect 640 -3055 670 -3045
rect 695 -2875 765 -2865
rect 695 -2895 700 -2875
rect 720 -2895 740 -2875
rect 760 -2895 765 -2875
rect 695 -2925 765 -2895
rect 695 -2945 700 -2925
rect 720 -2945 740 -2925
rect 760 -2945 765 -2925
rect 695 -2975 765 -2945
rect 695 -2995 700 -2975
rect 720 -2995 740 -2975
rect 760 -2995 765 -2975
rect 695 -3025 765 -2995
rect 695 -3045 700 -3025
rect 720 -3045 740 -3025
rect 760 -3045 765 -3025
rect 695 -3055 765 -3045
rect 805 -2875 835 -2865
rect 805 -2895 810 -2875
rect 830 -2895 835 -2875
rect 805 -2925 835 -2895
rect 805 -2945 810 -2925
rect 830 -2945 835 -2925
rect 805 -2975 835 -2945
rect 805 -2995 810 -2975
rect 830 -2995 835 -2975
rect 805 -3025 835 -2995
rect 805 -3045 810 -3025
rect 830 -3045 835 -3025
rect 805 -3055 835 -3045
rect 860 -2875 890 -2865
rect 860 -2895 865 -2875
rect 885 -2895 890 -2875
rect 860 -2925 890 -2895
rect 860 -2945 865 -2925
rect 885 -2945 890 -2925
rect 860 -2975 890 -2945
rect 860 -2995 865 -2975
rect 885 -2995 890 -2975
rect 860 -3025 890 -2995
rect 860 -3045 865 -3025
rect 885 -3045 890 -3025
rect 860 -3055 890 -3045
rect 915 -2875 945 -2865
rect 915 -2895 920 -2875
rect 940 -2895 945 -2875
rect 915 -2925 945 -2895
rect 915 -2945 920 -2925
rect 940 -2945 945 -2925
rect 915 -2975 945 -2945
rect 915 -2995 920 -2975
rect 940 -2995 945 -2975
rect 915 -3025 945 -2995
rect 915 -3045 920 -3025
rect 940 -3045 945 -3025
rect 915 -3055 945 -3045
rect 985 -2875 1055 -2865
rect 985 -2895 990 -2875
rect 1010 -2895 1030 -2875
rect 1050 -2895 1055 -2875
rect 985 -2925 1055 -2895
rect 985 -2945 990 -2925
rect 1010 -2945 1030 -2925
rect 1050 -2945 1055 -2925
rect 985 -2975 1055 -2945
rect 985 -2995 990 -2975
rect 1010 -2995 1030 -2975
rect 1050 -2995 1055 -2975
rect 985 -3025 1055 -2995
rect 985 -3045 990 -3025
rect 1010 -3045 1030 -3025
rect 1050 -3045 1055 -3025
rect 985 -3055 1055 -3045
rect 1080 -2875 1110 -2865
rect 1080 -2895 1085 -2875
rect 1105 -2895 1110 -2875
rect 1080 -2925 1110 -2895
rect 1080 -2945 1085 -2925
rect 1105 -2945 1110 -2925
rect 1080 -2975 1110 -2945
rect 1080 -2995 1085 -2975
rect 1105 -2995 1110 -2975
rect 1080 -3025 1110 -2995
rect 1080 -3045 1085 -3025
rect 1105 -3045 1110 -3025
rect 1080 -3055 1110 -3045
rect 1150 -2875 1220 -2865
rect 1150 -2895 1155 -2875
rect 1175 -2895 1195 -2875
rect 1215 -2895 1220 -2875
rect 1150 -2925 1220 -2895
rect 1150 -2945 1155 -2925
rect 1175 -2945 1195 -2925
rect 1215 -2945 1220 -2925
rect 1150 -2975 1220 -2945
rect 1150 -2995 1155 -2975
rect 1175 -2995 1195 -2975
rect 1215 -2995 1220 -2975
rect 1150 -3025 1220 -2995
rect 1150 -3045 1155 -3025
rect 1175 -3045 1195 -3025
rect 1215 -3045 1220 -3025
rect 1150 -3055 1220 -3045
rect 1245 -2875 1275 -2865
rect 1245 -2895 1250 -2875
rect 1270 -2895 1275 -2875
rect 1245 -2925 1275 -2895
rect 1245 -2945 1250 -2925
rect 1270 -2945 1275 -2925
rect 1245 -2975 1275 -2945
rect 1245 -2995 1250 -2975
rect 1270 -2995 1275 -2975
rect 1245 -3025 1275 -2995
rect 1245 -3045 1250 -3025
rect 1270 -3045 1275 -3025
rect 1245 -3055 1275 -3045
rect 1355 -2875 1445 -2865
rect 1355 -2895 1365 -2875
rect 1385 -2895 1415 -2875
rect 1435 -2895 1445 -2875
rect 1355 -2925 1445 -2895
rect 1355 -2945 1365 -2925
rect 1385 -2945 1415 -2925
rect 1435 -2945 1445 -2925
rect 1355 -2975 1445 -2945
rect 1355 -2995 1365 -2975
rect 1385 -2995 1415 -2975
rect 1435 -2995 1445 -2975
rect 1355 -3025 1445 -2995
rect 1355 -3045 1365 -3025
rect 1385 -3045 1415 -3025
rect 1435 -3045 1445 -3025
rect 1355 -3055 1445 -3045
rect 1470 -2875 1510 -2865
rect 1470 -2895 1480 -2875
rect 1500 -2895 1510 -2875
rect 1470 -2925 1510 -2895
rect 1470 -2945 1480 -2925
rect 1500 -2945 1510 -2925
rect 1470 -2975 1510 -2945
rect 1470 -2995 1480 -2975
rect 1500 -2995 1510 -2975
rect 1470 -3025 1510 -2995
rect 1470 -3045 1480 -3025
rect 1500 -3045 1510 -3025
rect 1470 -3055 1510 -3045
rect 1550 -2875 1640 -2865
rect 1550 -2895 1560 -2875
rect 1580 -2895 1610 -2875
rect 1630 -2895 1640 -2875
rect 1550 -2925 1640 -2895
rect 1550 -2945 1560 -2925
rect 1580 -2945 1610 -2925
rect 1630 -2945 1640 -2925
rect 1550 -2975 1640 -2945
rect 1550 -2995 1560 -2975
rect 1580 -2995 1610 -2975
rect 1630 -2995 1640 -2975
rect 1550 -3025 1640 -2995
rect 1550 -3045 1560 -3025
rect 1580 -3045 1610 -3025
rect 1630 -3045 1640 -3025
rect 1550 -3055 1640 -3045
rect 1665 -2875 1705 -2865
rect 1665 -2895 1675 -2875
rect 1695 -2895 1705 -2875
rect 1665 -2925 1705 -2895
rect 1665 -2945 1675 -2925
rect 1695 -2945 1705 -2925
rect 1665 -2975 1705 -2945
rect 1665 -2995 1675 -2975
rect 1695 -2995 1705 -2975
rect 1665 -3025 1705 -2995
rect 1665 -3045 1675 -3025
rect 1695 -3045 1705 -3025
rect 1665 -3055 1705 -3045
rect 1745 -2875 1835 -2865
rect 1745 -2895 1755 -2875
rect 1775 -2895 1805 -2875
rect 1825 -2895 1835 -2875
rect 1745 -2925 1835 -2895
rect 1745 -2945 1755 -2925
rect 1775 -2945 1805 -2925
rect 1825 -2945 1835 -2925
rect 1745 -2975 1835 -2945
rect 1745 -2995 1755 -2975
rect 1775 -2995 1805 -2975
rect 1825 -2995 1835 -2975
rect 1745 -3025 1835 -2995
rect 1745 -3045 1755 -3025
rect 1775 -3045 1805 -3025
rect 1825 -3045 1835 -3025
rect 1745 -3055 1835 -3045
rect 1860 -2875 1900 -2865
rect 1860 -2895 1870 -2875
rect 1890 -2895 1900 -2875
rect 1860 -2925 1900 -2895
rect 1860 -2945 1870 -2925
rect 1890 -2945 1900 -2925
rect 1860 -2975 1900 -2945
rect 1860 -2995 1870 -2975
rect 1890 -2995 1900 -2975
rect 1860 -3025 1900 -2995
rect 1860 -3045 1870 -3025
rect 1890 -3045 1900 -3025
rect 1860 -3055 1900 -3045
rect 1940 -2875 1980 -2865
rect 1940 -2895 1950 -2875
rect 1970 -2895 1980 -2875
rect 1940 -2925 1980 -2895
rect 1940 -2945 1950 -2925
rect 1970 -2945 1980 -2925
rect 1940 -2975 1980 -2945
rect 1940 -2995 1950 -2975
rect 1970 -2995 1980 -2975
rect 1940 -3025 1980 -2995
rect 1940 -3045 1950 -3025
rect 1970 -3045 1980 -3025
rect 1940 -3055 1980 -3045
rect 2005 -2875 2045 -2865
rect 2005 -2895 2015 -2875
rect 2035 -2895 2045 -2875
rect 2005 -2925 2045 -2895
rect 2005 -2945 2015 -2925
rect 2035 -2945 2045 -2925
rect 2005 -2975 2045 -2945
rect 2005 -2995 2015 -2975
rect 2035 -2995 2045 -2975
rect 2005 -3025 2045 -2995
rect 2005 -3045 2015 -3025
rect 2035 -3045 2045 -3025
rect 2005 -3055 2045 -3045
rect 2085 -2875 2175 -2865
rect 2085 -2895 2095 -2875
rect 2115 -2895 2145 -2875
rect 2165 -2895 2175 -2875
rect 2085 -2925 2175 -2895
rect 2085 -2945 2095 -2925
rect 2115 -2945 2145 -2925
rect 2165 -2945 2175 -2925
rect 2085 -2975 2175 -2945
rect 2085 -2995 2095 -2975
rect 2115 -2995 2145 -2975
rect 2165 -2995 2175 -2975
rect 2085 -3025 2175 -2995
rect 2085 -3045 2095 -3025
rect 2115 -3045 2145 -3025
rect 2165 -3045 2175 -3025
rect 2085 -3055 2175 -3045
rect 2200 -2875 2240 -2865
rect 2200 -2895 2210 -2875
rect 2230 -2895 2240 -2875
rect 2200 -2925 2240 -2895
rect 2200 -2945 2210 -2925
rect 2230 -2945 2240 -2925
rect 2200 -2975 2240 -2945
rect 2200 -2995 2210 -2975
rect 2230 -2995 2240 -2975
rect 2200 -3025 2240 -2995
rect 2200 -3045 2210 -3025
rect 2230 -3045 2240 -3025
rect 2200 -3055 2240 -3045
rect -120 -3140 -100 -3055
rect 250 -3140 270 -3055
rect 330 -3140 350 -3055
rect 700 -3140 720 -3055
rect 810 -3085 850 -3075
rect 810 -3105 820 -3085
rect 840 -3105 850 -3085
rect 810 -3115 850 -3105
rect 870 -3140 890 -3055
rect 1030 -3140 1050 -3055
rect 1195 -3140 1215 -3055
rect 1415 -3140 1435 -3055
rect 1610 -3140 1630 -3055
rect 1805 -3140 1825 -3055
rect 2145 -3140 2165 -3055
rect -190 -3160 -160 -3140
rect -140 -3160 -110 -3140
rect -90 -3160 -60 -3140
rect -40 -3160 -10 -3140
rect 10 -3160 40 -3140
rect 60 -3160 90 -3140
rect 110 -3160 140 -3140
rect 160 -3160 190 -3140
rect 210 -3160 240 -3140
rect 260 -3160 290 -3140
rect 310 -3160 340 -3140
rect 360 -3160 390 -3140
rect 410 -3160 440 -3140
rect 460 -3160 490 -3140
rect 510 -3160 540 -3140
rect 560 -3160 590 -3140
rect 610 -3160 640 -3140
rect 660 -3160 690 -3140
rect 710 -3160 740 -3140
rect 760 -3160 790 -3140
rect 810 -3160 840 -3140
rect 860 -3160 890 -3140
rect 910 -3160 940 -3140
rect 960 -3160 990 -3140
rect 1010 -3160 1040 -3140
rect 1060 -3160 1090 -3140
rect 1110 -3160 1140 -3140
rect 1160 -3160 1190 -3140
rect 1210 -3160 1240 -3140
rect 1260 -3160 1290 -3140
rect 1310 -3160 1340 -3140
rect 1360 -3160 1390 -3140
rect 1410 -3160 1440 -3140
rect 1460 -3160 1490 -3140
rect 1510 -3160 1540 -3140
rect 1560 -3160 1590 -3140
rect 1610 -3160 1640 -3140
rect 1660 -3160 1690 -3140
rect 1710 -3160 1740 -3140
rect 1760 -3160 1790 -3140
rect 1810 -3160 1840 -3140
rect 1860 -3160 1890 -3140
rect 1910 -3160 1940 -3140
rect 1960 -3160 1990 -3140
rect 2010 -3160 2040 -3140
rect 2060 -3160 2090 -3140
rect 2110 -3160 2140 -3140
rect 2160 -3160 2190 -3140
rect 2210 -3160 2240 -3140
rect 2260 -3160 2305 -3140
rect -120 -3245 -100 -3160
rect 95 -3195 135 -3185
rect 95 -3215 105 -3195
rect 125 -3215 135 -3195
rect 95 -3225 135 -3215
rect 95 -3245 115 -3225
rect 250 -3245 270 -3160
rect 330 -3245 350 -3160
rect 700 -3245 720 -3160
rect 900 -3245 920 -3160
rect 1065 -3245 1085 -3160
rect 1230 -3245 1250 -3160
rect 1415 -3245 1435 -3160
rect 1620 -3195 1660 -3185
rect 1620 -3215 1630 -3195
rect 1650 -3215 1660 -3195
rect 1620 -3225 1660 -3215
rect 1805 -3245 1825 -3160
rect -165 -3255 -95 -3245
rect -165 -3275 -160 -3255
rect -140 -3275 -120 -3255
rect -100 -3275 -95 -3255
rect -165 -3305 -95 -3275
rect -165 -3325 -160 -3305
rect -140 -3325 -120 -3305
rect -100 -3325 -95 -3305
rect -165 -3355 -95 -3325
rect -165 -3375 -160 -3355
rect -140 -3375 -120 -3355
rect -100 -3375 -95 -3355
rect -165 -3405 -95 -3375
rect -165 -3425 -160 -3405
rect -140 -3425 -120 -3405
rect -100 -3425 -95 -3405
rect -165 -3435 -95 -3425
rect -70 -3255 -40 -3245
rect -70 -3275 -65 -3255
rect -45 -3275 -40 -3255
rect -70 -3305 -40 -3275
rect -70 -3325 -65 -3305
rect -45 -3325 -40 -3305
rect -70 -3355 -40 -3325
rect -70 -3375 -65 -3355
rect -45 -3375 -40 -3355
rect -70 -3405 -40 -3375
rect -70 -3425 -65 -3405
rect -45 -3425 -40 -3405
rect -70 -3435 -40 -3425
rect -15 -3255 75 -3245
rect -15 -3275 -10 -3255
rect 10 -3270 45 -3255
rect 10 -3275 15 -3270
rect -15 -3305 15 -3275
rect 35 -3275 45 -3270
rect 65 -3275 75 -3255
rect 35 -3285 75 -3275
rect 95 -3255 165 -3245
rect 95 -3265 140 -3255
rect -15 -3325 -10 -3305
rect 10 -3325 15 -3305
rect -15 -3355 15 -3325
rect -15 -3375 -10 -3355
rect 10 -3375 15 -3355
rect -15 -3405 15 -3375
rect -15 -3425 -10 -3405
rect 10 -3425 15 -3405
rect -15 -3435 15 -3425
rect -10 -3455 10 -3435
rect -70 -3475 10 -3455
rect -70 -3555 -50 -3475
rect 95 -3495 115 -3265
rect 135 -3275 140 -3265
rect 160 -3275 165 -3255
rect 135 -3305 165 -3275
rect 135 -3325 140 -3305
rect 160 -3325 165 -3305
rect 135 -3355 165 -3325
rect 135 -3375 140 -3355
rect 160 -3375 165 -3355
rect 135 -3405 165 -3375
rect 135 -3425 140 -3405
rect 160 -3425 165 -3405
rect 135 -3435 165 -3425
rect 190 -3255 220 -3245
rect 190 -3275 195 -3255
rect 215 -3275 220 -3255
rect 190 -3305 220 -3275
rect 190 -3325 195 -3305
rect 215 -3325 220 -3305
rect 190 -3355 220 -3325
rect 190 -3375 195 -3355
rect 215 -3375 220 -3355
rect 190 -3405 220 -3375
rect 190 -3425 195 -3405
rect 215 -3425 220 -3405
rect 190 -3435 220 -3425
rect 245 -3255 355 -3245
rect 245 -3275 250 -3255
rect 270 -3275 290 -3255
rect 310 -3275 330 -3255
rect 350 -3275 355 -3255
rect 245 -3305 355 -3275
rect 245 -3325 250 -3305
rect 270 -3325 290 -3305
rect 310 -3325 330 -3305
rect 350 -3325 355 -3305
rect 245 -3355 355 -3325
rect 245 -3375 250 -3355
rect 270 -3375 290 -3355
rect 310 -3375 330 -3355
rect 350 -3375 355 -3355
rect 245 -3405 355 -3375
rect 245 -3425 250 -3405
rect 270 -3425 290 -3405
rect 310 -3425 330 -3405
rect 350 -3425 355 -3405
rect 245 -3435 355 -3425
rect 380 -3255 410 -3245
rect 380 -3275 385 -3255
rect 405 -3275 410 -3255
rect 380 -3305 410 -3275
rect 380 -3325 385 -3305
rect 405 -3325 410 -3305
rect 380 -3355 410 -3325
rect 380 -3375 385 -3355
rect 405 -3375 410 -3355
rect 380 -3405 410 -3375
rect 380 -3425 385 -3405
rect 405 -3425 410 -3405
rect 380 -3435 410 -3425
rect 435 -3255 525 -3245
rect 435 -3275 440 -3255
rect 460 -3270 495 -3255
rect 460 -3275 465 -3270
rect 435 -3305 465 -3275
rect 485 -3275 495 -3270
rect 515 -3275 525 -3255
rect 485 -3285 525 -3275
rect 545 -3255 615 -3245
rect 545 -3265 590 -3255
rect 435 -3325 440 -3305
rect 460 -3325 465 -3305
rect 435 -3355 465 -3325
rect 435 -3375 440 -3355
rect 460 -3375 465 -3355
rect 435 -3405 465 -3375
rect 435 -3425 440 -3405
rect 460 -3425 465 -3405
rect 435 -3435 465 -3425
rect 140 -3455 160 -3435
rect 440 -3455 460 -3435
rect 140 -3475 215 -3455
rect -25 -3505 115 -3495
rect -25 -3525 -15 -3505
rect 5 -3515 115 -3505
rect 5 -3525 15 -3515
rect -25 -3535 15 -3525
rect 195 -3555 215 -3475
rect 235 -3465 460 -3455
rect 235 -3485 245 -3465
rect 265 -3475 460 -3465
rect 265 -3485 275 -3475
rect 235 -3495 275 -3485
rect 380 -3555 400 -3475
rect 545 -3495 565 -3265
rect 585 -3275 590 -3265
rect 610 -3275 615 -3255
rect 585 -3305 615 -3275
rect 585 -3325 590 -3305
rect 610 -3325 615 -3305
rect 585 -3355 615 -3325
rect 585 -3375 590 -3355
rect 610 -3375 615 -3355
rect 585 -3405 615 -3375
rect 585 -3425 590 -3405
rect 610 -3425 615 -3405
rect 585 -3435 615 -3425
rect 640 -3255 670 -3245
rect 640 -3275 645 -3255
rect 665 -3275 670 -3255
rect 640 -3305 670 -3275
rect 640 -3325 645 -3305
rect 665 -3325 670 -3305
rect 640 -3355 670 -3325
rect 640 -3375 645 -3355
rect 665 -3375 670 -3355
rect 640 -3405 670 -3375
rect 640 -3425 645 -3405
rect 665 -3425 670 -3405
rect 640 -3435 670 -3425
rect 695 -3255 765 -3245
rect 695 -3275 700 -3255
rect 720 -3275 740 -3255
rect 760 -3275 765 -3255
rect 695 -3305 765 -3275
rect 695 -3325 700 -3305
rect 720 -3325 740 -3305
rect 760 -3325 765 -3305
rect 695 -3355 765 -3325
rect 695 -3375 700 -3355
rect 720 -3375 740 -3355
rect 760 -3375 765 -3355
rect 695 -3405 765 -3375
rect 695 -3425 700 -3405
rect 720 -3425 740 -3405
rect 760 -3425 765 -3405
rect 695 -3435 765 -3425
rect 840 -3255 870 -3245
rect 840 -3275 845 -3255
rect 865 -3275 870 -3255
rect 840 -3305 870 -3275
rect 840 -3325 845 -3305
rect 865 -3325 870 -3305
rect 840 -3355 870 -3325
rect 840 -3375 845 -3355
rect 865 -3375 870 -3355
rect 840 -3405 870 -3375
rect 840 -3425 845 -3405
rect 865 -3425 870 -3405
rect 840 -3435 870 -3425
rect 895 -3255 965 -3245
rect 895 -3275 900 -3255
rect 920 -3275 940 -3255
rect 960 -3275 965 -3255
rect 895 -3305 965 -3275
rect 895 -3325 900 -3305
rect 920 -3325 940 -3305
rect 960 -3325 965 -3305
rect 895 -3355 965 -3325
rect 895 -3375 900 -3355
rect 920 -3375 940 -3355
rect 960 -3375 965 -3355
rect 895 -3405 965 -3375
rect 895 -3425 900 -3405
rect 920 -3425 940 -3405
rect 960 -3425 965 -3405
rect 895 -3435 965 -3425
rect 1005 -3255 1035 -3245
rect 1005 -3275 1010 -3255
rect 1030 -3275 1035 -3255
rect 1005 -3305 1035 -3275
rect 1005 -3325 1010 -3305
rect 1030 -3325 1035 -3305
rect 1005 -3355 1035 -3325
rect 1005 -3375 1010 -3355
rect 1030 -3375 1035 -3355
rect 1005 -3405 1035 -3375
rect 1005 -3425 1010 -3405
rect 1030 -3425 1035 -3405
rect 1005 -3435 1035 -3425
rect 1060 -3255 1130 -3245
rect 1060 -3275 1065 -3255
rect 1085 -3275 1105 -3255
rect 1125 -3275 1130 -3255
rect 1060 -3305 1130 -3275
rect 1060 -3325 1065 -3305
rect 1085 -3325 1105 -3305
rect 1125 -3325 1130 -3305
rect 1060 -3355 1130 -3325
rect 1060 -3375 1065 -3355
rect 1085 -3375 1105 -3355
rect 1125 -3375 1130 -3355
rect 1060 -3405 1130 -3375
rect 1060 -3425 1065 -3405
rect 1085 -3425 1105 -3405
rect 1125 -3425 1130 -3405
rect 1060 -3435 1130 -3425
rect 1170 -3255 1200 -3245
rect 1170 -3275 1175 -3255
rect 1195 -3275 1200 -3255
rect 1170 -3305 1200 -3275
rect 1170 -3325 1175 -3305
rect 1195 -3325 1200 -3305
rect 1170 -3355 1200 -3325
rect 1170 -3375 1175 -3355
rect 1195 -3375 1200 -3355
rect 1170 -3405 1200 -3375
rect 1170 -3425 1175 -3405
rect 1195 -3425 1200 -3405
rect 1170 -3435 1200 -3425
rect 1225 -3255 1295 -3245
rect 1225 -3275 1230 -3255
rect 1250 -3275 1270 -3255
rect 1290 -3275 1295 -3255
rect 1225 -3305 1295 -3275
rect 1225 -3325 1230 -3305
rect 1250 -3325 1270 -3305
rect 1290 -3325 1295 -3305
rect 1225 -3355 1295 -3325
rect 1225 -3375 1230 -3355
rect 1250 -3375 1270 -3355
rect 1290 -3375 1295 -3355
rect 1225 -3405 1295 -3375
rect 1225 -3425 1230 -3405
rect 1250 -3425 1270 -3405
rect 1290 -3425 1295 -3405
rect 1225 -3435 1295 -3425
rect 1355 -3255 1445 -3245
rect 1355 -3275 1365 -3255
rect 1385 -3275 1415 -3255
rect 1435 -3275 1445 -3255
rect 1355 -3305 1445 -3275
rect 1355 -3325 1365 -3305
rect 1385 -3325 1415 -3305
rect 1435 -3325 1445 -3305
rect 1355 -3355 1445 -3325
rect 1355 -3375 1365 -3355
rect 1385 -3375 1415 -3355
rect 1435 -3375 1445 -3355
rect 1355 -3405 1445 -3375
rect 1355 -3425 1365 -3405
rect 1385 -3425 1415 -3405
rect 1435 -3425 1445 -3405
rect 1355 -3435 1445 -3425
rect 1470 -3255 1510 -3245
rect 1470 -3275 1480 -3255
rect 1500 -3275 1510 -3255
rect 1470 -3305 1510 -3275
rect 1470 -3325 1480 -3305
rect 1500 -3325 1510 -3305
rect 1470 -3355 1510 -3325
rect 1470 -3375 1480 -3355
rect 1500 -3375 1510 -3355
rect 1470 -3405 1510 -3375
rect 1470 -3425 1480 -3405
rect 1500 -3425 1510 -3405
rect 1470 -3435 1510 -3425
rect 1600 -3255 1640 -3245
rect 1600 -3275 1610 -3255
rect 1630 -3275 1640 -3255
rect 1600 -3305 1640 -3275
rect 1600 -3325 1610 -3305
rect 1630 -3325 1640 -3305
rect 1600 -3355 1640 -3325
rect 1600 -3375 1610 -3355
rect 1630 -3375 1640 -3355
rect 1600 -3405 1640 -3375
rect 1600 -3425 1610 -3405
rect 1630 -3425 1640 -3405
rect 1600 -3435 1640 -3425
rect 1665 -3255 1705 -3245
rect 1665 -3275 1675 -3255
rect 1695 -3275 1705 -3255
rect 1665 -3305 1705 -3275
rect 1665 -3325 1675 -3305
rect 1695 -3325 1705 -3305
rect 1665 -3355 1705 -3325
rect 1665 -3375 1675 -3355
rect 1695 -3375 1705 -3355
rect 1665 -3405 1705 -3375
rect 1665 -3425 1675 -3405
rect 1695 -3425 1705 -3405
rect 1665 -3435 1705 -3425
rect 1745 -3255 1835 -3245
rect 1745 -3275 1755 -3255
rect 1775 -3275 1805 -3255
rect 1825 -3275 1835 -3255
rect 1745 -3305 1835 -3275
rect 1745 -3325 1755 -3305
rect 1775 -3325 1805 -3305
rect 1825 -3325 1835 -3305
rect 1745 -3355 1835 -3325
rect 1745 -3375 1755 -3355
rect 1775 -3375 1805 -3355
rect 1825 -3375 1835 -3355
rect 1745 -3405 1835 -3375
rect 1745 -3425 1755 -3405
rect 1775 -3425 1805 -3405
rect 1825 -3425 1835 -3405
rect 1745 -3435 1835 -3425
rect 1860 -3255 1900 -3245
rect 1860 -3275 1870 -3255
rect 1890 -3275 1900 -3255
rect 1860 -3305 1900 -3275
rect 1860 -3325 1870 -3305
rect 1890 -3325 1900 -3305
rect 1860 -3355 1900 -3325
rect 1860 -3375 1870 -3355
rect 1890 -3375 1900 -3355
rect 1860 -3405 1900 -3375
rect 1860 -3425 1870 -3405
rect 1890 -3425 1900 -3405
rect 1860 -3435 1900 -3425
rect 1940 -3255 1980 -3245
rect 1940 -3275 1950 -3255
rect 1970 -3275 1980 -3255
rect 1940 -3305 1980 -3275
rect 1940 -3325 1950 -3305
rect 1970 -3325 1980 -3305
rect 1940 -3355 1980 -3325
rect 1940 -3375 1950 -3355
rect 1970 -3375 1980 -3355
rect 1940 -3405 1980 -3375
rect 1940 -3425 1950 -3405
rect 1970 -3425 1980 -3405
rect 1940 -3435 1980 -3425
rect 2005 -3255 2045 -3245
rect 2005 -3275 2015 -3255
rect 2035 -3275 2045 -3255
rect 2005 -3305 2045 -3275
rect 2005 -3325 2015 -3305
rect 2035 -3325 2045 -3305
rect 2005 -3355 2045 -3325
rect 2005 -3375 2015 -3355
rect 2035 -3375 2045 -3355
rect 2005 -3405 2045 -3375
rect 2005 -3425 2015 -3405
rect 2035 -3425 2045 -3405
rect 2005 -3435 2045 -3425
rect 590 -3455 610 -3435
rect 590 -3475 665 -3455
rect 840 -3470 860 -3435
rect 1005 -3470 1025 -3435
rect 1170 -3470 1190 -3435
rect 1480 -3455 1500 -3435
rect 1610 -3455 1630 -3435
rect 425 -3505 565 -3495
rect 425 -3525 435 -3505
rect 455 -3515 565 -3505
rect 455 -3525 465 -3515
rect 425 -3535 465 -3525
rect 645 -3555 665 -3475
rect 730 -3480 770 -3470
rect 730 -3500 740 -3480
rect 760 -3500 770 -3480
rect 730 -3510 770 -3500
rect 810 -3480 860 -3470
rect 810 -3500 820 -3480
rect 840 -3500 860 -3480
rect 810 -3510 860 -3500
rect 975 -3480 1025 -3470
rect 975 -3500 985 -3480
rect 1005 -3500 1025 -3480
rect 975 -3510 1025 -3500
rect 1140 -3480 1190 -3470
rect 1140 -3500 1150 -3480
rect 1170 -3500 1190 -3480
rect 1140 -3510 1190 -3500
rect 1270 -3480 1310 -3470
rect 1480 -3475 1630 -3455
rect 1270 -3500 1280 -3480
rect 1300 -3500 1310 -3480
rect 1270 -3510 1310 -3500
rect 1335 -3485 1375 -3475
rect 1335 -3505 1345 -3485
rect 1365 -3505 1375 -3485
rect 840 -3555 860 -3510
rect 1005 -3555 1025 -3510
rect 1170 -3555 1190 -3510
rect 1335 -3515 1375 -3505
rect 1480 -3555 1500 -3475
rect 1610 -3555 1630 -3475
rect 1675 -3455 1695 -3435
rect 1675 -3465 1725 -3455
rect 1675 -3485 1695 -3465
rect 1715 -3485 1725 -3465
rect 1675 -3495 1725 -3485
rect 1675 -3555 1695 -3495
rect 1880 -3505 1900 -3435
rect 1880 -3510 1920 -3505
rect 1880 -3530 1890 -3510
rect 1910 -3530 1920 -3510
rect 1880 -3540 1920 -3530
rect 1880 -3555 1900 -3540
rect 1950 -3555 1970 -3435
rect 2015 -3495 2035 -3435
rect 2015 -3515 2325 -3495
rect 2015 -3555 2035 -3515
rect 2210 -3555 2230 -3515
rect -165 -3565 -95 -3555
rect -165 -3585 -160 -3565
rect -140 -3585 -120 -3565
rect -100 -3585 -95 -3565
rect -165 -3615 -95 -3585
rect -165 -3635 -160 -3615
rect -140 -3635 -120 -3615
rect -100 -3635 -95 -3615
rect -165 -3645 -95 -3635
rect -70 -3565 -40 -3555
rect -70 -3585 -65 -3565
rect -45 -3585 -40 -3565
rect -70 -3615 -40 -3585
rect -70 -3635 -65 -3615
rect -45 -3635 -40 -3615
rect -70 -3645 -40 -3635
rect -15 -3565 15 -3555
rect -15 -3585 -10 -3565
rect 10 -3585 15 -3565
rect -15 -3615 15 -3585
rect -15 -3635 -10 -3615
rect 10 -3635 15 -3615
rect -15 -3645 15 -3635
rect 135 -3565 165 -3555
rect 135 -3585 140 -3565
rect 160 -3585 165 -3565
rect 135 -3615 165 -3585
rect 135 -3635 140 -3615
rect 160 -3635 165 -3615
rect 135 -3645 165 -3635
rect 190 -3565 220 -3555
rect 190 -3585 195 -3565
rect 215 -3585 220 -3565
rect 190 -3615 220 -3585
rect 190 -3635 195 -3615
rect 215 -3635 220 -3615
rect 190 -3645 220 -3635
rect 245 -3565 355 -3555
rect 245 -3585 250 -3565
rect 270 -3585 290 -3565
rect 310 -3585 330 -3565
rect 350 -3585 355 -3565
rect 245 -3615 355 -3585
rect 245 -3635 250 -3615
rect 270 -3635 290 -3615
rect 310 -3635 330 -3615
rect 350 -3635 355 -3615
rect 245 -3645 355 -3635
rect 380 -3565 410 -3555
rect 380 -3585 385 -3565
rect 405 -3585 410 -3565
rect 380 -3615 410 -3585
rect 380 -3635 385 -3615
rect 405 -3635 410 -3615
rect 380 -3645 410 -3635
rect 435 -3565 465 -3555
rect 435 -3585 440 -3565
rect 460 -3585 465 -3565
rect 435 -3615 465 -3585
rect 435 -3635 440 -3615
rect 460 -3635 465 -3615
rect 435 -3645 465 -3635
rect 585 -3565 615 -3555
rect 585 -3585 590 -3565
rect 610 -3585 615 -3565
rect 585 -3615 615 -3585
rect 585 -3635 590 -3615
rect 610 -3635 615 -3615
rect 585 -3645 615 -3635
rect 640 -3565 670 -3555
rect 640 -3585 645 -3565
rect 665 -3585 670 -3565
rect 640 -3615 670 -3585
rect 640 -3635 645 -3615
rect 665 -3635 670 -3615
rect 640 -3645 670 -3635
rect 695 -3565 765 -3555
rect 695 -3585 700 -3565
rect 720 -3585 740 -3565
rect 760 -3585 765 -3565
rect 695 -3615 765 -3585
rect 695 -3635 700 -3615
rect 720 -3635 740 -3615
rect 760 -3635 765 -3615
rect 695 -3645 765 -3635
rect 840 -3565 870 -3555
rect 840 -3585 845 -3565
rect 865 -3585 870 -3565
rect 840 -3615 870 -3585
rect 840 -3635 845 -3615
rect 865 -3635 870 -3615
rect 840 -3645 870 -3635
rect 895 -3565 965 -3555
rect 895 -3585 900 -3565
rect 920 -3585 940 -3565
rect 960 -3585 965 -3565
rect 895 -3615 965 -3585
rect 895 -3635 900 -3615
rect 920 -3635 940 -3615
rect 960 -3635 965 -3615
rect 895 -3645 965 -3635
rect 1005 -3565 1035 -3555
rect 1005 -3585 1010 -3565
rect 1030 -3585 1035 -3565
rect 1005 -3615 1035 -3585
rect 1005 -3635 1010 -3615
rect 1030 -3635 1035 -3615
rect 1005 -3645 1035 -3635
rect 1060 -3565 1130 -3555
rect 1060 -3585 1065 -3565
rect 1085 -3585 1105 -3565
rect 1125 -3585 1130 -3565
rect 1060 -3615 1130 -3585
rect 1060 -3635 1065 -3615
rect 1085 -3635 1105 -3615
rect 1125 -3635 1130 -3615
rect 1060 -3645 1130 -3635
rect 1170 -3565 1200 -3555
rect 1170 -3585 1175 -3565
rect 1195 -3585 1200 -3565
rect 1170 -3615 1200 -3585
rect 1170 -3635 1175 -3615
rect 1195 -3635 1200 -3615
rect 1170 -3645 1200 -3635
rect 1225 -3565 1295 -3555
rect 1225 -3585 1230 -3565
rect 1250 -3585 1270 -3565
rect 1290 -3585 1295 -3565
rect 1225 -3615 1295 -3585
rect 1225 -3635 1230 -3615
rect 1250 -3635 1270 -3615
rect 1290 -3635 1295 -3615
rect 1225 -3645 1295 -3635
rect 1355 -3565 1445 -3555
rect 1355 -3585 1365 -3565
rect 1385 -3585 1415 -3565
rect 1435 -3585 1445 -3565
rect 1355 -3615 1445 -3585
rect 1355 -3635 1365 -3615
rect 1385 -3635 1415 -3615
rect 1435 -3635 1445 -3615
rect 1355 -3645 1445 -3635
rect 1470 -3565 1510 -3555
rect 1470 -3585 1480 -3565
rect 1500 -3585 1510 -3565
rect 1470 -3615 1510 -3585
rect 1470 -3635 1480 -3615
rect 1500 -3635 1510 -3615
rect 1470 -3645 1510 -3635
rect 1600 -3565 1640 -3555
rect 1600 -3585 1610 -3565
rect 1630 -3585 1640 -3565
rect 1600 -3615 1640 -3585
rect 1600 -3635 1610 -3615
rect 1630 -3635 1640 -3615
rect 1600 -3645 1640 -3635
rect 1665 -3565 1705 -3555
rect 1665 -3585 1675 -3565
rect 1695 -3585 1705 -3565
rect 1665 -3615 1705 -3585
rect 1665 -3635 1675 -3615
rect 1695 -3635 1705 -3615
rect 1665 -3645 1705 -3635
rect 1745 -3565 1835 -3555
rect 1745 -3585 1755 -3565
rect 1775 -3585 1805 -3565
rect 1825 -3585 1835 -3565
rect 1745 -3615 1835 -3585
rect 1745 -3635 1755 -3615
rect 1775 -3635 1805 -3615
rect 1825 -3635 1835 -3615
rect 1745 -3645 1835 -3635
rect 1860 -3565 1900 -3555
rect 1860 -3585 1870 -3565
rect 1890 -3585 1900 -3565
rect 1860 -3615 1900 -3585
rect 1860 -3635 1870 -3615
rect 1890 -3635 1900 -3615
rect 1860 -3645 1900 -3635
rect 1940 -3565 1980 -3555
rect 1940 -3585 1950 -3565
rect 1970 -3585 1980 -3565
rect 1940 -3615 1980 -3585
rect 1940 -3635 1950 -3615
rect 1970 -3635 1980 -3615
rect 1940 -3645 1980 -3635
rect 2005 -3565 2045 -3555
rect 2005 -3585 2015 -3565
rect 2035 -3585 2045 -3565
rect 2005 -3615 2045 -3585
rect 2005 -3635 2015 -3615
rect 2035 -3635 2045 -3615
rect 2005 -3645 2045 -3635
rect 2085 -3565 2175 -3555
rect 2085 -3585 2095 -3565
rect 2115 -3585 2145 -3565
rect 2165 -3585 2175 -3565
rect 2085 -3615 2175 -3585
rect 2085 -3635 2095 -3615
rect 2115 -3635 2145 -3615
rect 2165 -3635 2175 -3615
rect 2085 -3645 2175 -3635
rect 2200 -3565 2240 -3555
rect 2200 -3585 2210 -3565
rect 2230 -3585 2240 -3565
rect 2200 -3615 2240 -3585
rect 2200 -3635 2210 -3615
rect 2230 -3635 2240 -3615
rect 2200 -3645 2240 -3635
rect -340 -3725 -290 -3710
rect -340 -3745 -325 -3725
rect -305 -3730 -290 -3725
rect -120 -3730 -100 -3645
rect -10 -3730 10 -3645
rect 140 -3730 160 -3645
rect 255 -3730 275 -3645
rect 330 -3730 350 -3645
rect 440 -3730 460 -3645
rect 590 -3730 610 -3645
rect 700 -3730 720 -3645
rect 900 -3730 920 -3645
rect 1065 -3730 1085 -3645
rect 1230 -3730 1250 -3645
rect 1415 -3730 1435 -3645
rect 1660 -3675 1700 -3665
rect 1660 -3695 1670 -3675
rect 1690 -3695 1700 -3675
rect 1660 -3705 1700 -3695
rect 1805 -3730 1825 -3645
rect 2145 -3730 2165 -3645
rect -305 -3745 -260 -3730
rect -340 -3750 -260 -3745
rect -240 -3750 -210 -3730
rect -190 -3750 -160 -3730
rect -140 -3750 -110 -3730
rect -90 -3750 -60 -3730
rect -40 -3750 -10 -3730
rect 10 -3750 40 -3730
rect 60 -3750 90 -3730
rect 110 -3750 140 -3730
rect 160 -3750 190 -3730
rect 210 -3750 240 -3730
rect 260 -3750 290 -3730
rect 310 -3750 340 -3730
rect 360 -3750 390 -3730
rect 410 -3750 440 -3730
rect 460 -3750 490 -3730
rect 510 -3750 540 -3730
rect 560 -3750 590 -3730
rect 610 -3750 640 -3730
rect 660 -3750 690 -3730
rect 710 -3750 740 -3730
rect 760 -3750 790 -3730
rect 810 -3750 840 -3730
rect 860 -3750 890 -3730
rect 910 -3750 940 -3730
rect 960 -3750 990 -3730
rect 1010 -3750 1040 -3730
rect 1060 -3750 1090 -3730
rect 1110 -3750 1140 -3730
rect 1160 -3750 1190 -3730
rect 1210 -3750 1240 -3730
rect 1260 -3750 1290 -3730
rect 1310 -3750 1340 -3730
rect 1360 -3750 1390 -3730
rect 1410 -3750 1440 -3730
rect 1460 -3750 1490 -3730
rect 1510 -3750 1540 -3730
rect 1560 -3750 1590 -3730
rect 1610 -3750 1640 -3730
rect 1660 -3750 1690 -3730
rect 1710 -3750 1740 -3730
rect 1760 -3750 1790 -3730
rect 1810 -3750 1840 -3730
rect 1860 -3750 1890 -3730
rect 1910 -3750 1940 -3730
rect 1960 -3750 1990 -3730
rect 2010 -3750 2040 -3730
rect 2060 -3750 2090 -3730
rect 2110 -3750 2140 -3730
rect 2160 -3750 2190 -3730
rect 2210 -3750 2240 -3730
rect 2260 -3750 2305 -3730
rect -340 -3760 -290 -3750
<< viali >>
rect -325 -2575 -305 -2555
rect -260 -2570 -240 -2550
rect -210 -2570 -190 -2550
rect -160 -2570 -140 -2550
rect -110 -2570 -90 -2550
rect -60 -2570 -40 -2550
rect -10 -2570 10 -2550
rect 40 -2570 60 -2550
rect 90 -2570 110 -2550
rect 140 -2570 160 -2550
rect 190 -2570 210 -2550
rect 240 -2570 260 -2550
rect 290 -2570 310 -2550
rect 340 -2570 360 -2550
rect 390 -2570 410 -2550
rect 440 -2570 460 -2550
rect 490 -2570 510 -2550
rect 540 -2570 560 -2550
rect 590 -2570 610 -2550
rect 640 -2570 660 -2550
rect 690 -2570 710 -2550
rect 740 -2570 760 -2550
rect 790 -2570 810 -2550
rect 840 -2570 860 -2550
rect 890 -2570 910 -2550
rect 940 -2570 960 -2550
rect 990 -2570 1010 -2550
rect 1040 -2570 1060 -2550
rect 1090 -2570 1110 -2550
rect 1140 -2570 1160 -2550
rect 1190 -2570 1210 -2550
rect 1240 -2570 1260 -2550
rect 1290 -2570 1310 -2550
rect 1340 -2570 1360 -2550
rect 1390 -2570 1410 -2550
rect 1440 -2570 1460 -2550
rect 1490 -2570 1510 -2550
rect 1540 -2570 1560 -2550
rect 1590 -2570 1610 -2550
rect 1640 -2570 1660 -2550
rect 1690 -2570 1710 -2550
rect 1740 -2570 1760 -2550
rect 1790 -2570 1810 -2550
rect 1840 -2570 1860 -2550
rect 1890 -2570 1910 -2550
rect 1940 -2570 1960 -2550
rect 1990 -2570 2010 -2550
rect 2040 -2570 2060 -2550
rect 2090 -2570 2110 -2550
rect 2140 -2570 2160 -2550
rect 2190 -2570 2210 -2550
rect 2240 -2570 2260 -2550
rect 85 -2625 105 -2605
rect 905 -2625 925 -2605
rect 730 -2800 750 -2780
rect 1275 -2820 1295 -2800
rect 1345 -2805 1365 -2785
rect 820 -3105 840 -3085
rect -160 -3160 -140 -3140
rect -110 -3160 -90 -3140
rect -60 -3160 -40 -3140
rect -10 -3160 10 -3140
rect 40 -3160 60 -3140
rect 90 -3160 110 -3140
rect 140 -3160 160 -3140
rect 190 -3160 210 -3140
rect 240 -3160 260 -3140
rect 290 -3160 310 -3140
rect 340 -3160 360 -3140
rect 390 -3160 410 -3140
rect 440 -3160 460 -3140
rect 490 -3160 510 -3140
rect 540 -3160 560 -3140
rect 590 -3160 610 -3140
rect 640 -3160 660 -3140
rect 690 -3160 710 -3140
rect 740 -3160 760 -3140
rect 790 -3160 810 -3140
rect 840 -3160 860 -3140
rect 890 -3160 910 -3140
rect 940 -3160 960 -3140
rect 990 -3160 1010 -3140
rect 1040 -3160 1060 -3140
rect 1090 -3160 1110 -3140
rect 1140 -3160 1160 -3140
rect 1190 -3160 1210 -3140
rect 1240 -3160 1260 -3140
rect 1290 -3160 1310 -3140
rect 1340 -3160 1360 -3140
rect 1390 -3160 1410 -3140
rect 1440 -3160 1460 -3140
rect 1490 -3160 1510 -3140
rect 1540 -3160 1560 -3140
rect 1590 -3160 1610 -3140
rect 1640 -3160 1660 -3140
rect 1690 -3160 1710 -3140
rect 1740 -3160 1760 -3140
rect 1790 -3160 1810 -3140
rect 1840 -3160 1860 -3140
rect 1890 -3160 1910 -3140
rect 1940 -3160 1960 -3140
rect 1990 -3160 2010 -3140
rect 2040 -3160 2060 -3140
rect 2090 -3160 2110 -3140
rect 2140 -3160 2160 -3140
rect 2190 -3160 2210 -3140
rect 2240 -3160 2260 -3140
rect 105 -3215 125 -3195
rect 1630 -3215 1650 -3195
rect 740 -3500 760 -3480
rect 1280 -3500 1300 -3480
rect 1345 -3505 1365 -3485
rect -325 -3745 -305 -3725
rect 1670 -3695 1690 -3675
rect -260 -3750 -240 -3730
rect -210 -3750 -190 -3730
rect -160 -3750 -140 -3730
rect -110 -3750 -90 -3730
rect -60 -3750 -40 -3730
rect -10 -3750 10 -3730
rect 40 -3750 60 -3730
rect 90 -3750 110 -3730
rect 140 -3750 160 -3730
rect 190 -3750 210 -3730
rect 240 -3750 260 -3730
rect 290 -3750 310 -3730
rect 340 -3750 360 -3730
rect 390 -3750 410 -3730
rect 440 -3750 460 -3730
rect 490 -3750 510 -3730
rect 540 -3750 560 -3730
rect 590 -3750 610 -3730
rect 640 -3750 660 -3730
rect 690 -3750 710 -3730
rect 740 -3750 760 -3730
rect 790 -3750 810 -3730
rect 840 -3750 860 -3730
rect 890 -3750 910 -3730
rect 940 -3750 960 -3730
rect 990 -3750 1010 -3730
rect 1040 -3750 1060 -3730
rect 1090 -3750 1110 -3730
rect 1140 -3750 1160 -3730
rect 1190 -3750 1210 -3730
rect 1240 -3750 1260 -3730
rect 1290 -3750 1310 -3730
rect 1340 -3750 1360 -3730
rect 1390 -3750 1410 -3730
rect 1440 -3750 1460 -3730
rect 1490 -3750 1510 -3730
rect 1540 -3750 1560 -3730
rect 1590 -3750 1610 -3730
rect 1640 -3750 1660 -3730
rect 1690 -3750 1710 -3730
rect 1740 -3750 1760 -3730
rect 1790 -3750 1810 -3730
rect 1840 -3750 1860 -3730
rect 1890 -3750 1910 -3730
rect 1940 -3750 1960 -3730
rect 1990 -3750 2010 -3730
rect 2040 -3750 2060 -3730
rect 2090 -3750 2110 -3730
rect 2140 -3750 2160 -3730
rect 2190 -3750 2210 -3730
rect 2240 -3750 2260 -3730
<< metal1 >>
rect -340 -2545 2255 -2540
rect -340 -2550 2305 -2545
rect -340 -2580 -330 -2550
rect -300 -2570 -260 -2550
rect -240 -2570 -210 -2550
rect -190 -2570 -160 -2550
rect -140 -2570 -110 -2550
rect -90 -2570 -60 -2550
rect -40 -2570 -10 -2550
rect 10 -2570 40 -2550
rect 60 -2570 90 -2550
rect 110 -2570 140 -2550
rect 160 -2570 190 -2550
rect 210 -2570 240 -2550
rect 260 -2570 290 -2550
rect 310 -2570 340 -2550
rect 360 -2570 390 -2550
rect 410 -2570 440 -2550
rect 460 -2570 490 -2550
rect 510 -2570 540 -2550
rect 560 -2570 590 -2550
rect 610 -2570 640 -2550
rect 660 -2570 690 -2550
rect 710 -2570 740 -2550
rect 760 -2570 790 -2550
rect 810 -2570 840 -2550
rect 860 -2570 890 -2550
rect 910 -2570 940 -2550
rect 960 -2570 990 -2550
rect 1010 -2570 1040 -2550
rect 1060 -2570 1090 -2550
rect 1110 -2570 1140 -2550
rect 1160 -2570 1190 -2550
rect 1210 -2570 1240 -2550
rect 1260 -2570 1290 -2550
rect 1310 -2570 1340 -2550
rect 1360 -2570 1390 -2550
rect 1410 -2570 1440 -2550
rect 1460 -2570 1490 -2550
rect 1510 -2570 1540 -2550
rect 1560 -2570 1590 -2550
rect 1610 -2570 1640 -2550
rect 1660 -2570 1690 -2550
rect 1710 -2570 1740 -2550
rect 1760 -2570 1790 -2550
rect 1810 -2570 1840 -2550
rect 1860 -2570 1890 -2550
rect 1910 -2570 1940 -2550
rect 1960 -2570 1990 -2550
rect 2010 -2570 2040 -2550
rect 2060 -2570 2090 -2550
rect 2110 -2570 2140 -2550
rect 2160 -2570 2190 -2550
rect 2210 -2570 2240 -2550
rect 2260 -2570 2305 -2550
rect -300 -2580 2305 -2570
rect -340 -2590 -290 -2580
rect 75 -2605 115 -2595
rect 75 -2625 85 -2605
rect 105 -2615 115 -2605
rect 895 -2605 935 -2595
rect 895 -2615 905 -2605
rect 105 -2625 905 -2615
rect 925 -2615 935 -2605
rect 925 -2625 1355 -2615
rect 75 -2635 1355 -2625
rect 720 -2775 760 -2770
rect 720 -2805 725 -2775
rect 755 -2805 760 -2775
rect 1335 -2775 1355 -2635
rect 1335 -2785 1375 -2775
rect 720 -2810 760 -2805
rect 1265 -2795 1305 -2790
rect 1265 -2825 1270 -2795
rect 1300 -2825 1305 -2795
rect 1335 -2805 1345 -2785
rect 1365 -2805 1375 -2785
rect 1335 -2815 1375 -2805
rect 1265 -2830 1305 -2825
rect 810 -3080 850 -3075
rect 810 -3110 815 -3080
rect 845 -3110 850 -3080
rect 810 -3115 850 -3110
rect -190 -3140 2305 -3130
rect -190 -3160 -160 -3140
rect -140 -3160 -110 -3140
rect -90 -3160 -60 -3140
rect -40 -3160 -10 -3140
rect 10 -3160 40 -3140
rect 60 -3160 90 -3140
rect 110 -3160 140 -3140
rect 160 -3160 190 -3140
rect 210 -3160 240 -3140
rect 260 -3160 290 -3140
rect 310 -3160 340 -3140
rect 360 -3160 390 -3140
rect 410 -3160 440 -3140
rect 460 -3160 490 -3140
rect 510 -3160 540 -3140
rect 560 -3160 590 -3140
rect 610 -3160 640 -3140
rect 660 -3160 690 -3140
rect 710 -3160 740 -3140
rect 760 -3160 790 -3140
rect 810 -3160 840 -3140
rect 860 -3160 890 -3140
rect 910 -3160 940 -3140
rect 960 -3160 990 -3140
rect 1010 -3160 1040 -3140
rect 1060 -3160 1090 -3140
rect 1110 -3160 1140 -3140
rect 1160 -3160 1190 -3140
rect 1210 -3160 1240 -3140
rect 1260 -3160 1290 -3140
rect 1310 -3160 1340 -3140
rect 1360 -3160 1390 -3140
rect 1410 -3160 1440 -3140
rect 1460 -3160 1490 -3140
rect 1510 -3160 1540 -3140
rect 1560 -3160 1590 -3140
rect 1610 -3160 1640 -3140
rect 1660 -3160 1690 -3140
rect 1710 -3160 1740 -3140
rect 1760 -3160 1790 -3140
rect 1810 -3160 1840 -3140
rect 1860 -3160 1890 -3140
rect 1910 -3160 1940 -3140
rect 1960 -3160 1990 -3140
rect 2010 -3160 2040 -3140
rect 2060 -3160 2090 -3140
rect 2110 -3160 2140 -3140
rect 2160 -3160 2190 -3140
rect 2210 -3160 2240 -3140
rect 2260 -3160 2305 -3140
rect -190 -3170 2305 -3160
rect 1680 -3185 1700 -3170
rect 95 -3195 135 -3185
rect 95 -3215 105 -3195
rect 125 -3200 135 -3195
rect 1620 -3190 1660 -3185
rect 125 -3205 1355 -3200
rect 125 -3215 785 -3205
rect 95 -3220 785 -3215
rect 95 -3225 135 -3220
rect 780 -3235 785 -3220
rect 815 -3220 1355 -3205
rect 815 -3235 820 -3220
rect 780 -3240 820 -3235
rect 730 -3475 770 -3470
rect 730 -3505 735 -3475
rect 765 -3505 770 -3475
rect 730 -3510 770 -3505
rect 1270 -3475 1310 -3470
rect 1270 -3505 1275 -3475
rect 1305 -3505 1310 -3475
rect 1270 -3510 1310 -3505
rect 1335 -3475 1355 -3220
rect 1620 -3220 1625 -3190
rect 1655 -3220 1660 -3190
rect 1620 -3225 1660 -3220
rect 1680 -3190 1720 -3185
rect 1680 -3220 1685 -3190
rect 1715 -3220 1720 -3190
rect 1680 -3225 1720 -3220
rect 1335 -3485 1375 -3475
rect 1335 -3505 1345 -3485
rect 1365 -3505 1375 -3485
rect 1335 -3515 1375 -3505
rect 1600 -3670 1640 -3665
rect 1600 -3700 1605 -3670
rect 1635 -3700 1640 -3670
rect 1600 -3705 1640 -3700
rect 1660 -3670 1700 -3665
rect 1660 -3700 1665 -3670
rect 1695 -3700 1700 -3670
rect 1660 -3705 1700 -3700
rect -340 -3720 -290 -3710
rect 1620 -3720 1640 -3705
rect -340 -3750 -330 -3720
rect -300 -3730 2305 -3720
rect -300 -3750 -260 -3730
rect -240 -3750 -210 -3730
rect -190 -3750 -160 -3730
rect -140 -3750 -110 -3730
rect -90 -3750 -60 -3730
rect -40 -3750 -10 -3730
rect 10 -3750 40 -3730
rect 60 -3750 90 -3730
rect 110 -3750 140 -3730
rect 160 -3750 190 -3730
rect 210 -3750 240 -3730
rect 260 -3750 290 -3730
rect 310 -3750 340 -3730
rect 360 -3750 390 -3730
rect 410 -3750 440 -3730
rect 460 -3750 490 -3730
rect 510 -3750 540 -3730
rect 560 -3750 590 -3730
rect 610 -3750 640 -3730
rect 660 -3750 690 -3730
rect 710 -3750 740 -3730
rect 760 -3750 790 -3730
rect 810 -3750 840 -3730
rect 860 -3750 890 -3730
rect 910 -3750 940 -3730
rect 960 -3750 990 -3730
rect 1010 -3750 1040 -3730
rect 1060 -3750 1090 -3730
rect 1110 -3750 1140 -3730
rect 1160 -3750 1190 -3730
rect 1210 -3750 1240 -3730
rect 1260 -3750 1290 -3730
rect 1310 -3750 1340 -3730
rect 1360 -3750 1390 -3730
rect 1410 -3750 1440 -3730
rect 1460 -3750 1490 -3730
rect 1510 -3750 1540 -3730
rect 1560 -3750 1590 -3730
rect 1610 -3750 1640 -3730
rect 1660 -3750 1690 -3730
rect 1710 -3750 1740 -3730
rect 1760 -3750 1790 -3730
rect 1810 -3750 1840 -3730
rect 1860 -3750 1890 -3730
rect 1910 -3750 1940 -3730
rect 1960 -3750 1990 -3730
rect 2010 -3750 2040 -3730
rect 2060 -3750 2090 -3730
rect 2110 -3750 2140 -3730
rect 2160 -3750 2190 -3730
rect 2210 -3750 2240 -3730
rect 2260 -3750 2305 -3730
rect -340 -3760 2305 -3750
<< via1 >>
rect -330 -2555 -300 -2550
rect -330 -2575 -325 -2555
rect -325 -2575 -305 -2555
rect -305 -2575 -300 -2555
rect -330 -2580 -300 -2575
rect 725 -2780 755 -2775
rect 725 -2800 730 -2780
rect 730 -2800 750 -2780
rect 750 -2800 755 -2780
rect 725 -2805 755 -2800
rect 1270 -2800 1300 -2795
rect 1270 -2820 1275 -2800
rect 1275 -2820 1295 -2800
rect 1295 -2820 1300 -2800
rect 1270 -2825 1300 -2820
rect 815 -3085 845 -3080
rect 815 -3105 820 -3085
rect 820 -3105 840 -3085
rect 840 -3105 845 -3085
rect 815 -3110 845 -3105
rect 785 -3235 815 -3205
rect 735 -3480 765 -3475
rect 735 -3500 740 -3480
rect 740 -3500 760 -3480
rect 760 -3500 765 -3480
rect 735 -3505 765 -3500
rect 1275 -3480 1305 -3475
rect 1275 -3500 1280 -3480
rect 1280 -3500 1300 -3480
rect 1300 -3500 1305 -3480
rect 1275 -3505 1305 -3500
rect 1625 -3195 1655 -3190
rect 1625 -3215 1630 -3195
rect 1630 -3215 1650 -3195
rect 1650 -3215 1655 -3195
rect 1625 -3220 1655 -3215
rect 1685 -3220 1715 -3190
rect 1605 -3700 1635 -3670
rect 1665 -3675 1695 -3670
rect 1665 -3695 1670 -3675
rect 1670 -3695 1690 -3675
rect 1690 -3695 1695 -3675
rect 1665 -3700 1695 -3695
rect -330 -3725 -300 -3720
rect -330 -3745 -325 -3725
rect -325 -3745 -305 -3725
rect -305 -3745 -300 -3725
rect -330 -3750 -300 -3745
<< metal2 >>
rect -340 -2550 -290 -2540
rect -340 -2580 -330 -2550
rect -300 -2580 -290 -2550
rect -340 -2590 -290 -2580
rect 720 -2775 760 -2770
rect 720 -2805 725 -2775
rect 755 -2805 760 -2775
rect 720 -2810 760 -2805
rect 740 -3470 760 -2810
rect 1265 -2795 1310 -2790
rect 1265 -2825 1270 -2795
rect 1300 -2825 1310 -2795
rect 1265 -2830 1310 -2825
rect 800 -3080 850 -3075
rect 800 -3110 815 -3080
rect 845 -3110 850 -3080
rect 800 -3115 850 -3110
rect 800 -3200 820 -3115
rect 780 -3205 820 -3200
rect 780 -3235 785 -3205
rect 815 -3235 820 -3205
rect 780 -3240 820 -3235
rect 1290 -3470 1310 -2830
rect 730 -3475 770 -3470
rect 730 -3505 735 -3475
rect 765 -3505 770 -3475
rect 730 -3510 770 -3505
rect 1270 -3475 1310 -3470
rect 1270 -3505 1275 -3475
rect 1305 -3505 1310 -3475
rect 1270 -3510 1310 -3505
rect 1620 -3190 1660 -3185
rect 1620 -3220 1625 -3190
rect 1655 -3220 1660 -3190
rect 1620 -3225 1660 -3220
rect 1680 -3190 1720 -3185
rect 1680 -3220 1685 -3190
rect 1715 -3220 1720 -3190
rect 1680 -3225 1720 -3220
rect 1620 -3665 1640 -3225
rect 1680 -3665 1700 -3225
rect 1600 -3670 1640 -3665
rect 1600 -3700 1605 -3670
rect 1635 -3700 1640 -3670
rect 1600 -3705 1640 -3700
rect 1660 -3670 1700 -3665
rect 1660 -3700 1665 -3670
rect 1695 -3700 1700 -3670
rect 1660 -3705 1700 -3700
rect -340 -3720 -290 -3710
rect -340 -3750 -330 -3720
rect -300 -3750 -290 -3720
rect -340 -3760 -290 -3750
<< via2 >>
rect -330 -2580 -300 -2550
rect -330 -3750 -300 -3720
<< metal3 >>
rect -340 -2545 -290 -2540
rect -340 -2585 -335 -2545
rect -295 -2585 -290 -2545
rect -340 -2590 -290 -2585
rect -340 -3715 -290 -3710
rect -340 -3755 -335 -3715
rect -295 -3755 -290 -3715
rect -340 -3760 -290 -3755
<< via3 >>
rect -335 -2550 -295 -2545
rect -335 -2580 -330 -2550
rect -330 -2580 -300 -2550
rect -300 -2580 -295 -2550
rect -335 -2585 -295 -2580
rect -335 -3720 -295 -3715
rect -335 -3750 -330 -3720
rect -330 -3750 -300 -3720
rect -300 -3750 -295 -3720
rect -335 -3755 -295 -3750
<< metal4 >>
rect -340 -2545 -290 -2540
rect -340 -2585 -335 -2545
rect -295 -2585 -290 -2545
rect -340 -3715 -290 -2585
rect -340 -3755 -335 -3715
rect -295 -3755 -290 -3715
rect -340 -3760 -290 -3755
<< labels >>
flabel poly 60 -2825 60 -2825 7 FreeSans 160 0 -80 0 QA_b
flabel poly -150 -2795 -150 -2795 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel locali 665 -2825 665 -2825 3 FreeSans 160 0 80 0 E_b
flabel locali 460 -2825 460 -2825 3 FreeSans 160 0 80 0 E
flabel poly -150 -3510 -150 -3510 7 FreeSans 160 0 -80 0 F_VCO
port 2 w
flabel poly 60 -3345 60 -3345 7 FreeSans 160 0 -80 0 QB_b
flabel locali 460 -3475 460 -3475 3 FreeSans 160 0 80 0 F
flabel locali 665 -3475 665 -3475 3 FreeSans 160 0 80 0 F_b
flabel locali 975 -2790 975 -2790 3 FreeSans 160 0 80 0 before_Reset
flabel locali 810 -3510 810 -3510 5 FreeSans 160 0 0 -80 Reset
flabel locali 2325 -3505 2325 -3505 3 FreeSans 160 0 80 0 DOWN_input
port 6 e
flabel locali 1510 -2775 1510 -2775 3 FreeSans 160 0 80 0 UP_PFD_b
flabel locali 1705 -2775 1705 -2775 3 FreeSans 160 0 80 0 UP
flabel locali 2325 -2810 2325 -2810 3 FreeSans 160 0 80 0 UP_input
port 5 e
flabel locali 1500 -3495 1500 -3495 3 FreeSans 160 0 80 0 DOWN_PFD_b
flabel poly 1820 -3480 1820 -3480 5 FreeSans 160 0 0 -80 DOWN_b
flabel metal4 -340 -3625 -340 -3625 7 FreeSans 160 0 -80 0 GNDA
port 4 w
flabel metal1 -190 -3150 -190 -3150 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel poly 2195 -3465 2195 -3465 3 FreeSans 160 0 80 0 DOWN
port 8 e
flabel locali 1970 -3515 1970 -3515 3 FreeSans 160 0 80 0 I_IN
port 10 e
flabel locali 1970 -2810 1970 -2810 3 FreeSans 160 0 80 0 opamp_out
flabel locali 1900 -2790 1900 -2790 3 FreeSans 160 0 80 0 UP_b
flabel locali 95 -2690 95 -2690 7 FreeSans 160 0 -80 0 QA
flabel locali 95 -3225 95 -3225 7 FreeSans 160 0 -80 0 QB
<< end >>
