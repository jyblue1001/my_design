magic
tech sky130A
timestamp 1739762179
<< nwell >>
rect -60 140 2525 380
<< nmos >>
rect 0 -50 15 50
rect 55 -50 70 50
rect 260 -50 275 50
rect 315 -50 330 50
rect 440 -50 455 50
rect 495 -50 510 50
rect 700 -50 715 50
rect 755 -50 770 50
rect 880 -50 895 50
rect 935 -50 950 50
rect 1140 -50 1155 50
rect 1195 -50 1210 50
rect 1330 -50 1345 50
rect 1385 -50 1400 50
rect 1590 -50 1605 50
rect 1645 -50 1660 50
rect 1770 -50 1785 50
rect 1825 -50 1840 50
rect 1950 -50 1965 50
rect 2075 -50 2090 50
rect 2200 -50 2215 50
rect 2325 -50 2340 50
rect 2450 -50 2465 50
<< pmos >>
rect 0 160 15 360
rect 55 160 70 360
rect 260 160 275 360
rect 315 160 330 360
rect 440 160 455 360
rect 495 160 510 360
rect 700 160 715 360
rect 755 160 770 360
rect 880 160 895 360
rect 935 160 950 360
rect 1140 160 1155 360
rect 1195 160 1210 360
rect 1330 160 1345 360
rect 1385 160 1400 360
rect 1590 160 1605 360
rect 1645 160 1660 360
rect 1770 160 1785 360
rect 1825 160 1840 360
rect 1950 160 1965 360
rect 2075 160 2090 360
rect 2200 160 2215 360
rect 2325 160 2340 360
rect 2450 160 2465 360
<< ndiff >>
rect -40 35 0 50
rect -40 -35 -30 35
rect -10 -35 0 35
rect -40 -50 0 -35
rect 15 35 55 50
rect 15 -35 25 35
rect 45 -35 55 35
rect 15 -50 55 -35
rect 70 35 110 50
rect 70 -35 80 35
rect 100 -35 110 35
rect 70 -50 110 -35
rect 220 35 260 50
rect 220 -35 230 35
rect 250 -35 260 35
rect 220 -50 260 -35
rect 275 35 315 50
rect 275 -35 285 35
rect 305 -35 315 35
rect 275 -50 315 -35
rect 330 35 370 50
rect 330 -35 340 35
rect 360 -35 370 35
rect 330 -50 370 -35
rect 400 35 440 50
rect 400 -35 410 35
rect 430 -35 440 35
rect 400 -50 440 -35
rect 455 35 495 50
rect 455 -35 465 35
rect 485 -35 495 35
rect 455 -50 495 -35
rect 510 35 550 50
rect 510 -35 520 35
rect 540 -35 550 35
rect 510 -50 550 -35
rect 660 35 700 50
rect 660 -35 670 35
rect 690 -35 700 35
rect 660 -50 700 -35
rect 715 35 755 50
rect 715 -35 725 35
rect 745 -35 755 35
rect 715 -50 755 -35
rect 770 35 810 50
rect 770 -35 780 35
rect 800 -35 810 35
rect 770 -50 810 -35
rect 840 35 880 50
rect 840 -35 850 35
rect 870 -35 880 35
rect 840 -50 880 -35
rect 895 35 935 50
rect 895 -35 905 35
rect 925 -35 935 35
rect 895 -50 935 -35
rect 950 35 990 50
rect 950 -35 960 35
rect 980 -35 990 35
rect 950 -50 990 -35
rect 1100 35 1140 50
rect 1100 -35 1110 35
rect 1130 -35 1140 35
rect 1100 -50 1140 -35
rect 1155 35 1195 50
rect 1155 -35 1165 35
rect 1185 -35 1195 35
rect 1155 -50 1195 -35
rect 1210 35 1250 50
rect 1290 35 1330 50
rect 1210 -35 1220 35
rect 1240 -35 1250 35
rect 1290 -35 1300 35
rect 1320 -35 1330 35
rect 1210 -50 1250 -35
rect 1290 -50 1330 -35
rect 1345 35 1385 50
rect 1345 -35 1355 35
rect 1375 -35 1385 35
rect 1345 -50 1385 -35
rect 1400 35 1440 50
rect 1400 -35 1410 35
rect 1430 -35 1440 35
rect 1400 -50 1440 -35
rect 1550 35 1590 50
rect 1550 -35 1560 35
rect 1580 -35 1590 35
rect 1550 -50 1590 -35
rect 1605 35 1645 50
rect 1605 -35 1615 35
rect 1635 -35 1645 35
rect 1605 -50 1645 -35
rect 1660 35 1700 50
rect 1660 -35 1670 35
rect 1690 -35 1700 35
rect 1660 -50 1700 -35
rect 1730 35 1770 50
rect 1730 -35 1740 35
rect 1760 -35 1770 35
rect 1730 -50 1770 -35
rect 1785 35 1825 50
rect 1785 -35 1795 35
rect 1815 -35 1825 35
rect 1785 -50 1825 -35
rect 1840 35 1880 50
rect 1840 -35 1850 35
rect 1870 -35 1880 35
rect 1840 -50 1880 -35
rect 1910 35 1950 50
rect 1910 -35 1920 35
rect 1940 -35 1950 35
rect 1910 -50 1950 -35
rect 1965 35 2005 50
rect 1965 -35 1975 35
rect 1995 -35 2005 35
rect 1965 -50 2005 -35
rect 2035 35 2075 50
rect 2035 -35 2045 35
rect 2065 -35 2075 35
rect 2035 -50 2075 -35
rect 2090 35 2130 50
rect 2090 -35 2100 35
rect 2120 -35 2130 35
rect 2090 -50 2130 -35
rect 2160 35 2200 50
rect 2160 -35 2170 35
rect 2190 -35 2200 35
rect 2160 -50 2200 -35
rect 2215 35 2255 50
rect 2215 -35 2225 35
rect 2245 -35 2255 35
rect 2215 -50 2255 -35
rect 2285 35 2325 50
rect 2285 -35 2295 35
rect 2315 -35 2325 35
rect 2285 -50 2325 -35
rect 2340 35 2380 50
rect 2340 -35 2350 35
rect 2370 -35 2380 35
rect 2340 -50 2380 -35
rect 2410 35 2450 50
rect 2410 -35 2420 35
rect 2440 -35 2450 35
rect 2410 -50 2450 -35
rect 2465 35 2505 50
rect 2465 -35 2475 35
rect 2495 -35 2505 35
rect 2465 -50 2505 -35
<< pdiff >>
rect -40 345 0 360
rect -40 175 -30 345
rect -10 175 0 345
rect -40 160 0 175
rect 15 345 55 360
rect 15 175 25 345
rect 45 175 55 345
rect 15 160 55 175
rect 70 345 110 360
rect 70 175 80 345
rect 100 175 110 345
rect 70 160 110 175
rect 220 345 260 360
rect 220 175 230 345
rect 250 175 260 345
rect 220 160 260 175
rect 275 345 315 360
rect 275 175 285 345
rect 305 175 315 345
rect 275 160 315 175
rect 330 345 370 360
rect 330 175 340 345
rect 360 175 370 345
rect 330 160 370 175
rect 400 345 440 360
rect 400 175 410 345
rect 430 175 440 345
rect 400 160 440 175
rect 455 345 495 360
rect 455 175 465 345
rect 485 175 495 345
rect 455 160 495 175
rect 510 345 550 360
rect 510 175 520 345
rect 540 175 550 345
rect 510 160 550 175
rect 660 345 700 360
rect 660 175 670 345
rect 690 175 700 345
rect 660 160 700 175
rect 715 345 755 360
rect 715 175 725 345
rect 745 175 755 345
rect 715 160 755 175
rect 770 345 810 360
rect 770 175 780 345
rect 800 175 810 345
rect 770 160 810 175
rect 840 345 880 360
rect 840 175 850 345
rect 870 175 880 345
rect 840 160 880 175
rect 895 345 935 360
rect 895 175 905 345
rect 925 175 935 345
rect 895 160 935 175
rect 950 345 990 360
rect 950 175 960 345
rect 980 175 990 345
rect 950 160 990 175
rect 1100 345 1140 360
rect 1100 175 1110 345
rect 1130 175 1140 345
rect 1100 160 1140 175
rect 1155 345 1195 360
rect 1155 175 1165 345
rect 1185 175 1195 345
rect 1155 160 1195 175
rect 1210 345 1250 360
rect 1290 345 1330 360
rect 1210 175 1220 345
rect 1240 175 1250 345
rect 1290 175 1300 345
rect 1320 175 1330 345
rect 1210 160 1250 175
rect 1290 160 1330 175
rect 1345 345 1385 360
rect 1345 175 1355 345
rect 1375 175 1385 345
rect 1345 160 1385 175
rect 1400 345 1440 360
rect 1400 175 1410 345
rect 1430 175 1440 345
rect 1400 160 1440 175
rect 1550 345 1590 360
rect 1550 175 1560 345
rect 1580 175 1590 345
rect 1550 160 1590 175
rect 1605 345 1645 360
rect 1605 175 1615 345
rect 1635 175 1645 345
rect 1605 160 1645 175
rect 1660 345 1700 360
rect 1660 175 1670 345
rect 1690 175 1700 345
rect 1660 160 1700 175
rect 1730 345 1770 360
rect 1730 175 1740 345
rect 1760 175 1770 345
rect 1730 160 1770 175
rect 1785 345 1825 360
rect 1785 175 1795 345
rect 1815 175 1825 345
rect 1785 160 1825 175
rect 1840 345 1880 360
rect 1840 175 1850 345
rect 1870 175 1880 345
rect 1840 160 1880 175
rect 1910 345 1950 360
rect 1910 175 1920 345
rect 1940 175 1950 345
rect 1910 160 1950 175
rect 1965 345 2005 360
rect 1965 175 1975 345
rect 1995 175 2005 345
rect 1965 160 2005 175
rect 2035 345 2075 360
rect 2035 175 2045 345
rect 2065 175 2075 345
rect 2035 160 2075 175
rect 2090 345 2130 360
rect 2090 175 2100 345
rect 2120 175 2130 345
rect 2090 160 2130 175
rect 2160 345 2200 360
rect 2160 175 2170 345
rect 2190 175 2200 345
rect 2160 160 2200 175
rect 2215 345 2255 360
rect 2215 175 2225 345
rect 2245 175 2255 345
rect 2215 160 2255 175
rect 2285 345 2325 360
rect 2285 175 2295 345
rect 2315 175 2325 345
rect 2285 160 2325 175
rect 2340 345 2380 360
rect 2340 175 2350 345
rect 2370 175 2380 345
rect 2340 160 2380 175
rect 2410 345 2450 360
rect 2410 175 2420 345
rect 2440 175 2450 345
rect 2410 160 2450 175
rect 2465 345 2505 360
rect 2465 175 2475 345
rect 2495 175 2505 345
rect 2465 160 2505 175
<< ndiffc >>
rect -30 -35 -10 35
rect 25 -35 45 35
rect 80 -35 100 35
rect 230 -35 250 35
rect 285 -35 305 35
rect 340 -35 360 35
rect 410 -35 430 35
rect 465 -35 485 35
rect 520 -35 540 35
rect 670 -35 690 35
rect 725 -35 745 35
rect 780 -35 800 35
rect 850 -35 870 35
rect 905 -35 925 35
rect 960 -35 980 35
rect 1110 -35 1130 35
rect 1165 -35 1185 35
rect 1220 -35 1240 35
rect 1300 -35 1320 35
rect 1355 -35 1375 35
rect 1410 -35 1430 35
rect 1560 -35 1580 35
rect 1615 -35 1635 35
rect 1670 -35 1690 35
rect 1740 -35 1760 35
rect 1795 -35 1815 35
rect 1850 -35 1870 35
rect 1920 -35 1940 35
rect 1975 -35 1995 35
rect 2045 -35 2065 35
rect 2100 -35 2120 35
rect 2170 -35 2190 35
rect 2225 -35 2245 35
rect 2295 -35 2315 35
rect 2350 -35 2370 35
rect 2420 -35 2440 35
rect 2475 -35 2495 35
<< pdiffc >>
rect -30 175 -10 345
rect 25 175 45 345
rect 80 175 100 345
rect 230 175 250 345
rect 285 175 305 345
rect 340 175 360 345
rect 410 175 430 345
rect 465 175 485 345
rect 520 175 540 345
rect 670 175 690 345
rect 725 175 745 345
rect 780 175 800 345
rect 850 175 870 345
rect 905 175 925 345
rect 960 175 980 345
rect 1110 175 1130 345
rect 1165 175 1185 345
rect 1220 175 1240 345
rect 1300 175 1320 345
rect 1355 175 1375 345
rect 1410 175 1430 345
rect 1560 175 1580 345
rect 1615 175 1635 345
rect 1670 175 1690 345
rect 1740 175 1760 345
rect 1795 175 1815 345
rect 1850 175 1870 345
rect 1920 175 1940 345
rect 1975 175 1995 345
rect 2045 175 2065 345
rect 2100 175 2120 345
rect 2170 175 2190 345
rect 2225 175 2245 345
rect 2295 175 2315 345
rect 2350 175 2370 345
rect 2420 175 2440 345
rect 2475 175 2495 345
<< psubdiff >>
rect 1250 35 1290 50
rect 1250 -35 1260 35
rect 1280 -35 1290 35
rect 1250 -50 1290 -35
<< nsubdiff >>
rect 1250 345 1290 360
rect 1250 175 1260 345
rect 1280 175 1290 345
rect 1250 160 1290 175
<< psubdiffcont >>
rect 1260 -35 1280 35
<< nsubdiffcont >>
rect 1260 175 1280 345
<< poly >>
rect 755 440 2530 455
rect 185 405 225 415
rect 185 385 195 405
rect 215 385 225 405
rect 185 375 225 385
rect 0 360 15 375
rect 55 360 70 375
rect 260 360 275 375
rect 315 360 330 375
rect 440 360 455 375
rect 495 360 510 375
rect 700 360 715 375
rect 755 360 770 440
rect 880 360 895 375
rect 935 360 950 375
rect 1140 360 1155 375
rect 1195 360 1210 375
rect 1330 360 1345 375
rect 1385 360 1400 375
rect 1590 360 1605 375
rect 1645 360 1660 440
rect 1745 405 1785 415
rect 1745 385 1755 405
rect 1775 385 1785 405
rect 1745 375 1785 385
rect 1770 360 1785 375
rect 1825 360 1840 375
rect 1950 360 1965 375
rect 2075 360 2090 375
rect 2200 360 2215 375
rect 2325 360 2340 375
rect 2450 360 2465 375
rect 125 345 165 355
rect 125 225 135 345
rect 155 225 165 345
rect 125 215 165 225
rect 0 100 15 160
rect -60 85 15 100
rect 0 50 15 85
rect 55 105 70 160
rect 55 95 105 105
rect 55 75 75 95
rect 95 75 105 95
rect 55 65 105 75
rect 150 85 165 215
rect 565 345 605 355
rect 565 225 575 345
rect 595 225 605 345
rect 565 215 605 225
rect 260 85 275 160
rect 150 70 275 85
rect 55 50 70 65
rect 260 50 275 70
rect 315 145 330 160
rect 315 135 365 145
rect 315 115 335 135
rect 355 115 365 135
rect 315 105 365 115
rect 315 50 330 105
rect 440 50 455 160
rect 495 105 510 160
rect 495 95 545 105
rect 495 75 515 95
rect 535 75 545 95
rect 495 65 545 75
rect 590 85 605 215
rect 1005 345 1045 355
rect 1005 225 1015 345
rect 1035 225 1045 345
rect 1005 215 1045 225
rect 700 85 715 160
rect 590 70 715 85
rect 495 50 510 65
rect 700 50 715 70
rect 755 50 770 160
rect 880 50 895 160
rect 935 105 950 160
rect 935 95 985 105
rect 935 75 955 95
rect 975 75 985 95
rect 935 65 985 75
rect 1030 85 1045 215
rect 1455 345 1495 355
rect 1455 225 1465 345
rect 1485 225 1495 345
rect 1455 215 1495 225
rect 1140 85 1155 160
rect 1030 70 1155 85
rect 935 50 950 65
rect 1140 50 1155 70
rect 1195 145 1210 160
rect 1195 135 1245 145
rect 1195 115 1215 135
rect 1235 115 1245 135
rect 1195 105 1245 115
rect 1195 50 1210 105
rect 1330 50 1345 160
rect 1385 105 1400 160
rect 1385 95 1435 105
rect 1385 75 1405 95
rect 1425 75 1435 95
rect 1385 65 1435 75
rect 1480 85 1495 215
rect 1590 85 1605 160
rect 1480 70 1605 85
rect 1385 50 1400 65
rect 1590 50 1605 70
rect 1645 50 1660 160
rect 1770 50 1785 160
rect 1825 50 1840 160
rect 1865 120 1905 130
rect 1865 100 1875 120
rect 1895 115 1905 120
rect 1950 115 1965 160
rect 1895 100 1965 115
rect 1865 90 1905 100
rect 1950 50 1965 100
rect 1990 120 2030 130
rect 1990 100 2000 120
rect 2020 115 2030 120
rect 2075 115 2090 160
rect 2020 100 2090 115
rect 1990 90 2030 100
rect 2075 50 2090 100
rect 2115 120 2155 130
rect 2115 100 2125 120
rect 2145 115 2155 120
rect 2200 115 2215 160
rect 2145 100 2215 115
rect 2115 90 2155 100
rect 2200 50 2215 100
rect 2240 120 2280 130
rect 2240 100 2250 120
rect 2270 115 2280 120
rect 2325 115 2340 160
rect 2270 100 2340 115
rect 2240 90 2280 100
rect 2325 50 2340 100
rect 2365 120 2405 130
rect 2365 100 2375 120
rect 2395 115 2405 120
rect 2450 115 2465 160
rect 2515 130 2530 440
rect 2395 100 2465 115
rect 2365 90 2405 100
rect 2450 50 2465 100
rect 2490 120 2530 130
rect 2490 100 2500 120
rect 2520 100 2530 120
rect 2490 90 2530 100
rect 0 -65 15 -50
rect 55 -65 70 -50
rect 260 -90 275 -50
rect 315 -65 330 -50
rect 440 -90 455 -50
rect 495 -65 510 -50
rect 700 -65 715 -50
rect 755 -65 770 -50
rect 260 -105 455 -90
rect 880 -130 895 -50
rect 935 -65 950 -50
rect 1140 -90 1155 -50
rect 1195 -65 1210 -50
rect 1330 -90 1345 -50
rect 1385 -65 1400 -50
rect 1590 -65 1605 -50
rect 1645 -65 1660 -50
rect 1770 -65 1785 -50
rect 1825 -65 1840 -50
rect 1950 -65 1965 -50
rect 2075 -65 2090 -50
rect 2200 -65 2215 -50
rect 2325 -65 2340 -50
rect 2450 -65 2465 -50
rect 1140 -105 1345 -90
rect 1825 -75 1865 -65
rect 1825 -95 1835 -75
rect 1855 -95 1865 -75
rect 1825 -105 1865 -95
rect -60 -145 895 -130
<< polycont >>
rect 195 385 215 405
rect 1755 385 1775 405
rect 135 225 155 345
rect 75 75 95 95
rect 575 225 595 345
rect 335 115 355 135
rect 515 75 535 95
rect 1015 225 1035 345
rect 955 75 975 95
rect 1465 225 1485 345
rect 1215 115 1235 135
rect 1405 75 1425 95
rect 1875 100 1895 120
rect 2000 100 2020 120
rect 2125 100 2145 120
rect 2250 100 2270 120
rect 2375 100 2395 120
rect 2500 100 2520 120
rect 1835 -95 1855 -75
<< locali >>
rect 185 405 225 415
rect 185 385 195 405
rect 215 395 225 405
rect 1745 405 1785 415
rect 1745 395 1755 405
rect 215 385 1755 395
rect 1775 395 1785 405
rect 1775 385 2530 395
rect 185 375 2530 385
rect 185 355 205 375
rect -35 345 -5 355
rect -35 175 -30 345
rect -10 175 -5 345
rect -35 165 -5 175
rect 20 345 50 355
rect 20 175 25 345
rect 45 175 50 345
rect 20 165 50 175
rect 75 345 165 355
rect 75 175 80 345
rect 100 230 135 345
rect 100 175 105 230
rect 125 225 135 230
rect 155 225 165 345
rect 125 215 165 225
rect 185 345 255 355
rect 185 235 230 345
rect 75 165 105 175
rect 80 145 100 165
rect 20 125 100 145
rect 20 45 40 125
rect 185 105 205 235
rect 225 175 230 235
rect 250 175 255 345
rect 225 165 255 175
rect 280 345 310 355
rect 280 175 285 345
rect 305 175 310 345
rect 280 165 310 175
rect 335 345 365 355
rect 335 175 340 345
rect 360 175 365 345
rect 335 165 365 175
rect 405 345 435 355
rect 405 175 410 345
rect 430 175 435 345
rect 405 165 435 175
rect 460 345 490 355
rect 460 175 465 345
rect 485 175 490 345
rect 460 165 490 175
rect 515 345 605 355
rect 515 175 520 345
rect 540 230 575 345
rect 540 175 545 230
rect 565 225 575 230
rect 595 225 605 345
rect 565 215 605 225
rect 625 345 695 355
rect 625 235 670 345
rect 515 165 545 175
rect 230 145 250 165
rect 520 145 540 165
rect 230 125 305 145
rect 65 95 205 105
rect 65 75 75 95
rect 95 85 205 95
rect 95 75 105 85
rect 65 65 105 75
rect 285 45 305 125
rect 325 135 540 145
rect 325 115 335 135
rect 355 125 540 135
rect 355 115 365 125
rect 325 105 365 115
rect 460 45 480 125
rect 625 105 645 235
rect 665 175 670 235
rect 690 175 695 345
rect 665 165 695 175
rect 720 345 750 355
rect 720 175 725 345
rect 745 175 750 345
rect 720 165 750 175
rect 775 345 805 355
rect 775 175 780 345
rect 800 175 805 345
rect 775 165 805 175
rect 845 345 875 355
rect 845 175 850 345
rect 870 175 875 345
rect 845 165 875 175
rect 900 345 930 355
rect 900 175 905 345
rect 925 175 930 345
rect 900 165 930 175
rect 955 345 1045 355
rect 955 175 960 345
rect 980 230 1015 345
rect 980 175 985 230
rect 1005 225 1015 230
rect 1035 225 1045 345
rect 1005 215 1045 225
rect 1065 345 1135 355
rect 1065 235 1110 345
rect 955 165 985 175
rect 670 145 690 165
rect 960 145 980 165
rect 670 125 745 145
rect 505 95 645 105
rect 505 75 515 95
rect 535 85 645 95
rect 535 75 545 85
rect 505 65 545 75
rect 725 45 745 125
rect 900 125 980 145
rect 900 45 920 125
rect 1065 105 1085 235
rect 1105 175 1110 235
rect 1130 175 1135 345
rect 1105 165 1135 175
rect 1160 345 1190 355
rect 1160 175 1165 345
rect 1185 175 1190 345
rect 1160 165 1190 175
rect 1215 345 1325 355
rect 1215 175 1220 345
rect 1240 175 1260 345
rect 1280 175 1300 345
rect 1320 175 1325 345
rect 1215 165 1325 175
rect 1350 345 1380 355
rect 1350 175 1355 345
rect 1375 175 1380 345
rect 1350 165 1380 175
rect 1405 345 1495 355
rect 1405 175 1410 345
rect 1430 230 1465 345
rect 1430 175 1435 230
rect 1455 225 1465 230
rect 1485 225 1495 345
rect 1455 215 1495 225
rect 1515 345 1585 355
rect 1515 235 1560 345
rect 1405 165 1435 175
rect 1110 145 1130 165
rect 1410 145 1430 165
rect 1110 125 1185 145
rect 945 95 1085 105
rect 945 75 955 95
rect 975 85 1085 95
rect 975 75 985 85
rect 945 65 985 75
rect 1165 45 1185 125
rect 1205 135 1430 145
rect 1205 115 1215 135
rect 1235 125 1430 135
rect 1235 115 1245 125
rect 1205 105 1245 115
rect 1350 45 1370 125
rect 1515 105 1535 235
rect 1555 175 1560 235
rect 1580 175 1585 345
rect 1555 165 1585 175
rect 1610 345 1640 355
rect 1610 175 1615 345
rect 1635 175 1640 345
rect 1610 165 1640 175
rect 1665 345 1695 355
rect 1665 175 1670 345
rect 1690 175 1695 345
rect 1665 165 1695 175
rect 1735 345 1765 355
rect 1735 175 1740 345
rect 1760 175 1765 345
rect 1735 165 1765 175
rect 1790 345 1820 355
rect 1790 175 1795 345
rect 1815 175 1820 345
rect 1790 165 1820 175
rect 1845 345 1875 355
rect 1845 175 1850 345
rect 1870 175 1875 345
rect 1845 165 1875 175
rect 1915 345 1945 355
rect 1915 175 1920 345
rect 1940 175 1945 345
rect 1915 165 1945 175
rect 1970 345 2000 355
rect 1970 175 1975 345
rect 1995 175 2000 345
rect 1970 165 2000 175
rect 2040 345 2070 355
rect 2040 175 2045 345
rect 2065 175 2070 345
rect 2040 165 2070 175
rect 2095 345 2125 355
rect 2095 175 2100 345
rect 2120 175 2125 345
rect 2095 165 2125 175
rect 2165 345 2195 355
rect 2165 175 2170 345
rect 2190 175 2195 345
rect 2165 165 2195 175
rect 2220 345 2250 355
rect 2220 175 2225 345
rect 2245 175 2250 345
rect 2220 165 2250 175
rect 2290 345 2320 355
rect 2290 175 2295 345
rect 2315 175 2320 345
rect 2290 165 2320 175
rect 2345 345 2375 355
rect 2345 175 2350 345
rect 2370 175 2375 345
rect 2345 165 2375 175
rect 2415 345 2445 355
rect 2415 175 2420 345
rect 2440 175 2445 345
rect 2415 165 2445 175
rect 2470 345 2500 355
rect 2470 175 2475 345
rect 2495 175 2500 345
rect 2470 165 2500 175
rect 1560 145 1580 165
rect 1740 145 1760 165
rect 1850 145 1870 165
rect 1560 125 1635 145
rect 1740 130 1870 145
rect 1980 130 2000 165
rect 2105 130 2125 165
rect 2230 130 2250 165
rect 2355 130 2375 165
rect 2480 130 2500 165
rect 1740 125 1905 130
rect 1395 95 1535 105
rect 1395 75 1405 95
rect 1425 85 1535 95
rect 1425 75 1435 85
rect 1395 65 1435 75
rect 1615 45 1635 125
rect 1850 120 1905 125
rect 1850 100 1875 120
rect 1895 100 1905 120
rect 1850 90 1905 100
rect 1980 120 2030 130
rect 1980 100 2000 120
rect 2020 100 2030 120
rect 1980 90 2030 100
rect 2105 120 2155 130
rect 2105 100 2125 120
rect 2145 100 2155 120
rect 2105 90 2155 100
rect 2230 120 2280 130
rect 2230 100 2250 120
rect 2270 100 2280 120
rect 2230 90 2280 100
rect 2355 120 2405 130
rect 2355 100 2375 120
rect 2395 100 2405 120
rect 2355 90 2405 100
rect 2480 120 2530 130
rect 2480 100 2500 120
rect 2520 100 2530 120
rect 2480 90 2530 100
rect 1850 45 1870 90
rect 1980 45 2000 90
rect 2105 45 2125 90
rect 2230 45 2250 90
rect 2355 45 2375 90
rect 2480 45 2500 90
rect -35 35 -5 45
rect -35 -35 -30 35
rect -10 -35 -5 35
rect -35 -45 -5 -35
rect 20 35 50 45
rect 20 -35 25 35
rect 45 -35 50 35
rect 20 -45 50 -35
rect 75 35 105 45
rect 75 -35 80 35
rect 100 -35 105 35
rect 75 -45 105 -35
rect 225 35 255 45
rect 225 -35 230 35
rect 250 -35 255 35
rect 225 -45 255 -35
rect 280 35 310 45
rect 280 -35 285 35
rect 305 -35 310 35
rect 280 -45 310 -35
rect 335 35 365 45
rect 335 -35 340 35
rect 360 -35 365 35
rect 335 -45 365 -35
rect 405 35 435 45
rect 405 -35 410 35
rect 430 -35 435 35
rect 405 -45 435 -35
rect 460 35 490 45
rect 460 -35 465 35
rect 485 -35 490 35
rect 460 -45 490 -35
rect 515 35 545 45
rect 515 -35 520 35
rect 540 -35 545 35
rect 515 -45 545 -35
rect 665 35 695 45
rect 665 -35 670 35
rect 690 -35 695 35
rect 665 -45 695 -35
rect 720 35 750 45
rect 720 -35 725 35
rect 745 -35 750 35
rect 720 -45 750 -35
rect 775 35 805 45
rect 775 -35 780 35
rect 800 -35 805 35
rect 775 -45 805 -35
rect 845 35 875 45
rect 845 -35 850 35
rect 870 -35 875 35
rect 845 -45 875 -35
rect 900 35 930 45
rect 900 -35 905 35
rect 925 -35 930 35
rect 900 -45 930 -35
rect 955 35 985 45
rect 955 -35 960 35
rect 980 -35 985 35
rect 955 -45 985 -35
rect 1105 35 1135 45
rect 1105 -35 1110 35
rect 1130 -35 1135 35
rect 1105 -45 1135 -35
rect 1160 35 1190 45
rect 1160 -35 1165 35
rect 1185 -35 1190 35
rect 1160 -45 1190 -35
rect 1215 35 1325 45
rect 1215 -35 1220 35
rect 1240 -35 1260 35
rect 1280 -35 1300 35
rect 1320 -35 1325 35
rect 1215 -45 1325 -35
rect 1350 35 1380 45
rect 1350 -35 1355 35
rect 1375 -35 1380 35
rect 1350 -45 1380 -35
rect 1405 35 1435 45
rect 1405 -35 1410 35
rect 1430 -35 1435 35
rect 1405 -45 1435 -35
rect 1555 35 1585 45
rect 1555 -35 1560 35
rect 1580 -35 1585 35
rect 1555 -45 1585 -35
rect 1610 35 1640 45
rect 1610 -35 1615 35
rect 1635 -35 1640 35
rect 1610 -45 1640 -35
rect 1665 35 1695 45
rect 1665 -35 1670 35
rect 1690 -35 1695 35
rect 1665 -45 1695 -35
rect 1735 35 1765 45
rect 1735 -35 1740 35
rect 1760 -35 1765 35
rect 1735 -45 1765 -35
rect 1790 35 1820 45
rect 1790 -35 1795 35
rect 1815 -35 1820 35
rect 1790 -45 1820 -35
rect 1845 35 1875 45
rect 1845 -35 1850 35
rect 1870 -35 1875 35
rect 1845 -45 1875 -35
rect 1915 35 1945 45
rect 1915 -35 1920 35
rect 1940 -35 1945 35
rect 1915 -45 1945 -35
rect 1970 35 2000 45
rect 1970 -35 1975 35
rect 1995 -35 2000 35
rect 1970 -45 2000 -35
rect 2040 35 2070 45
rect 2040 -35 2045 35
rect 2065 -35 2070 35
rect 2040 -45 2070 -35
rect 2095 35 2125 45
rect 2095 -35 2100 35
rect 2120 -35 2125 35
rect 2095 -45 2125 -35
rect 2165 35 2195 45
rect 2165 -35 2170 35
rect 2190 -35 2195 35
rect 2165 -45 2195 -35
rect 2220 35 2250 45
rect 2220 -35 2225 35
rect 2245 -35 2250 35
rect 2220 -45 2250 -35
rect 2290 35 2320 45
rect 2290 -35 2295 35
rect 2315 -35 2320 35
rect 2290 -45 2320 -35
rect 2345 35 2375 45
rect 2345 -35 2350 35
rect 2370 -35 2375 35
rect 2345 -45 2375 -35
rect 2415 35 2445 45
rect 2415 -35 2420 35
rect 2440 -35 2445 35
rect 2415 -45 2445 -35
rect 2470 35 2500 45
rect 2470 -35 2475 35
rect 2495 -35 2500 35
rect 2470 -45 2500 -35
rect 1165 -65 1185 -45
rect 1165 -75 2530 -65
rect 1165 -85 1835 -75
rect 1825 -95 1835 -85
rect 1855 -85 2530 -75
rect 1855 -95 1865 -85
rect 1825 -105 1865 -95
<< viali >>
rect -30 175 -10 345
rect 340 175 360 345
rect 410 175 430 345
rect 780 175 800 345
rect 850 175 870 345
rect 1220 175 1240 345
rect 1260 175 1280 345
rect 1300 175 1320 345
rect 1670 175 1690 345
rect 1795 175 1815 345
rect 1920 175 1940 345
rect 2045 175 2065 345
rect 2170 175 2190 345
rect 2295 175 2315 345
rect 2420 175 2440 345
rect -30 -35 -10 35
rect 80 -35 100 35
rect 230 -35 250 35
rect 340 -35 360 35
rect 410 -35 430 35
rect 520 -35 540 35
rect 670 -35 690 35
rect 780 -35 800 35
rect 850 -35 870 35
rect 960 -35 980 35
rect 1110 -35 1130 35
rect 1220 -35 1240 35
rect 1260 -35 1280 35
rect 1300 -35 1320 35
rect 1410 -35 1430 35
rect 1560 -35 1580 35
rect 1670 -35 1690 35
rect 1740 -35 1760 35
rect 1920 -35 1940 35
rect 2045 -35 2065 35
rect 2170 -35 2190 35
rect 2295 -35 2315 35
rect 2420 -35 2440 35
<< metal1 >>
rect -40 345 2505 360
rect -40 175 -30 345
rect -10 175 340 345
rect 360 175 410 345
rect 430 175 780 345
rect 800 175 850 345
rect 870 175 1220 345
rect 1240 175 1260 345
rect 1280 175 1300 345
rect 1320 175 1670 345
rect 1690 175 1795 345
rect 1815 175 1920 345
rect 1940 175 2045 345
rect 2065 175 2170 345
rect 2190 175 2295 345
rect 2315 175 2420 345
rect 2440 175 2505 345
rect -40 160 2505 175
rect -40 35 2505 50
rect -40 -35 -30 35
rect -10 -35 80 35
rect 100 -35 230 35
rect 250 -35 340 35
rect 360 -35 410 35
rect 430 -35 520 35
rect 540 -35 670 35
rect 690 -35 780 35
rect 800 -35 850 35
rect 870 -35 960 35
rect 980 -35 1110 35
rect 1130 -35 1220 35
rect 1240 -35 1260 35
rect 1280 -35 1300 35
rect 1320 -35 1410 35
rect 1430 -35 1560 35
rect 1580 -35 1670 35
rect 1690 -35 1740 35
rect 1760 -35 1920 35
rect 1940 -35 2045 35
rect 2065 -35 2170 35
rect 2190 -35 2295 35
rect 2315 -35 2420 35
rect 2440 -35 2505 35
rect -40 -50 2505 -35
<< labels >>
flabel poly -60 95 -60 95 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel poly 150 125 150 125 7 FreeSans 160 0 -80 0 QA_b
flabel locali 540 125 540 125 3 FreeSans 160 0 80 0 E
flabel locali 745 125 745 125 3 FreeSans 160 0 80 0 E_b
flabel locali 1905 130 1905 130 3 FreeSans 160 0 80 0 before_Reset
flabel poly 1030 135 1030 135 7 FreeSans 160 0 -80 0 QB_b
flabel locali 1430 125 1430 125 3 FreeSans 160 0 80 0 F
flabel locali 1635 110 1635 110 3 FreeSans 160 0 80 0 F_b
flabel metal1 -40 25 -40 25 7 FreeSans 160 0 -80 0 GNDA
port 6 w
flabel metal1 -40 210 -40 210 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel poly -60 -135 -60 -135 7 FreeSans 160 0 -80 0 F_VCO
port 2 w
flabel locali 2530 -75 2530 -75 3 FreeSans 160 0 80 0 QB
port 5 e
flabel poly 770 425 770 425 3 FreeSans 160 0 80 0 Reset
flabel locali 2530 385 2530 385 3 FreeSans 160 0 80 0 QA
port 4 e
<< end >>
