magic
tech sky130A
timestamp 1754061271
<< nwell >>
rect 56025 4510 56365 4900
rect 56495 4510 56835 4730
rect 56965 4510 57305 4900
rect 57435 4510 57775 4900
rect 54610 3645 55490 4035
rect 55945 3645 56825 4035
rect 56975 3645 57855 4035
rect 58310 3645 59190 4035
rect 54640 2535 55460 3175
rect 56450 2890 57350 3180
rect 58340 2535 59160 3175
rect 58835 2530 58975 2535
rect 54640 1660 55460 1900
rect 58340 1660 59160 1900
<< nmos >>
rect 56810 2315 56825 2565
rect 56865 2315 56880 2565
rect 56920 2315 56935 2565
rect 56975 2315 56990 2565
rect 56070 1745 56085 1895
rect 56125 1745 56140 1895
rect 56180 1745 56195 1895
rect 56235 1745 56250 1895
rect 56290 1745 56305 1895
rect 56345 1745 56360 1895
rect 56400 1745 56415 1895
rect 56455 1745 56470 1895
rect 56510 1745 56525 1895
rect 56565 1745 56580 1895
rect 56620 1745 56635 1895
rect 56675 1745 56690 1895
rect 57110 1745 57125 1895
rect 57165 1745 57180 1895
rect 57220 1745 57235 1895
rect 57275 1745 57290 1895
rect 57330 1745 57345 1895
rect 57385 1745 57400 1895
rect 57440 1745 57455 1895
rect 57495 1745 57510 1895
rect 57550 1745 57565 1895
rect 57605 1745 57620 1895
rect 57660 1745 57675 1895
rect 57715 1745 57730 1895
rect 54740 1140 54755 1440
rect 54795 1140 54810 1440
rect 54850 1140 54865 1440
rect 54905 1140 54920 1440
rect 54960 1140 54975 1440
rect 55015 1140 55030 1440
rect 55070 1140 55085 1440
rect 55125 1140 55140 1440
rect 55180 1140 55195 1440
rect 55235 1140 55250 1440
rect 55290 1140 55305 1440
rect 55345 1140 55360 1440
rect 56070 1070 56085 1220
rect 56125 1070 56140 1220
rect 56180 1070 56195 1220
rect 56235 1070 56250 1220
rect 56290 1070 56305 1220
rect 56345 1070 56360 1220
rect 56400 1070 56415 1220
rect 56455 1070 56470 1220
rect 56510 1070 56525 1220
rect 56565 1070 56580 1220
rect 56620 1070 56635 1220
rect 56675 1070 56690 1220
rect 56810 1070 56825 1220
rect 56865 1070 56880 1220
rect 56920 1070 56935 1220
rect 56975 1070 56990 1220
rect 57110 1070 57125 1220
rect 57165 1070 57180 1220
rect 57220 1070 57235 1220
rect 57275 1070 57290 1220
rect 57330 1070 57345 1220
rect 57385 1070 57400 1220
rect 57440 1070 57455 1220
rect 57495 1070 57510 1220
rect 57550 1070 57565 1220
rect 57605 1070 57620 1220
rect 57660 1070 57675 1220
rect 57715 1070 57730 1220
rect 58440 1140 58455 1440
rect 58495 1140 58510 1440
rect 58550 1140 58565 1440
rect 58605 1140 58620 1440
rect 58660 1140 58675 1440
rect 58715 1140 58730 1440
rect 58770 1140 58785 1440
rect 58825 1140 58840 1440
rect 58880 1140 58895 1440
rect 58935 1140 58950 1440
rect 58990 1140 59005 1440
rect 59045 1140 59060 1440
rect 54770 -520 54830 180
rect 54870 -520 54930 180
rect 54970 -520 55030 180
rect 55070 -520 55130 180
rect 55170 -520 55230 180
rect 55270 -520 55330 180
rect 56260 80 56275 330
rect 56315 80 56330 330
rect 56370 80 56385 330
rect 56425 80 56440 330
rect 56480 80 56495 330
rect 56535 80 56550 330
rect 56590 80 56605 330
rect 56645 80 56660 330
rect 56700 80 56715 330
rect 56755 80 56770 330
rect 56810 80 56825 330
rect 56865 80 56880 330
rect 56920 80 56935 330
rect 56975 80 56990 330
rect 57030 80 57045 330
rect 57085 80 57100 330
rect 57140 80 57155 330
rect 57195 80 57210 330
rect 57250 80 57265 330
rect 57305 80 57320 330
rect 57360 80 57375 330
rect 57415 80 57430 330
rect 57470 80 57485 330
rect 56470 -475 56485 -325
rect 56525 -475 56540 -325
rect 56580 -475 56595 -325
rect 56635 -475 56650 -325
rect 56690 -475 56705 -325
rect 56745 -475 56760 -325
rect 56910 -475 57210 -325
rect 58470 -520 58530 180
rect 58570 -520 58630 180
rect 58670 -520 58730 180
rect 58770 -520 58830 180
rect 58870 -520 58930 180
rect 58970 -520 59030 180
<< pmos >>
rect 56125 4530 56145 4880
rect 56185 4530 56205 4880
rect 56245 4530 56265 4880
rect 56595 4530 56615 4710
rect 56655 4530 56675 4710
rect 56715 4530 56735 4710
rect 57065 4530 57085 4880
rect 57125 4530 57145 4880
rect 57185 4530 57205 4880
rect 57535 4530 57555 4880
rect 57595 4530 57615 4880
rect 57655 4530 57675 4880
rect 54710 3665 54730 4015
rect 54770 3665 54790 4015
rect 54830 3665 54850 4015
rect 54890 3665 54910 4015
rect 54950 3665 54970 4015
rect 55010 3665 55030 4015
rect 55070 3665 55090 4015
rect 55130 3665 55150 4015
rect 55190 3665 55210 4015
rect 55250 3665 55270 4015
rect 55310 3665 55330 4015
rect 55370 3665 55390 4015
rect 56045 3665 56065 4015
rect 56105 3665 56125 4015
rect 56165 3665 56185 4015
rect 56225 3665 56245 4015
rect 56285 3665 56305 4015
rect 56345 3665 56365 4015
rect 56405 3665 56425 4015
rect 56465 3665 56485 4015
rect 56525 3665 56545 4015
rect 56585 3665 56605 4015
rect 56645 3665 56665 4015
rect 56705 3665 56725 4015
rect 57075 3665 57095 4015
rect 57135 3665 57155 4015
rect 57195 3665 57215 4015
rect 57255 3665 57275 4015
rect 57315 3665 57335 4015
rect 57375 3665 57395 4015
rect 57435 3665 57455 4015
rect 57495 3665 57515 4015
rect 57555 3665 57575 4015
rect 57615 3665 57635 4015
rect 57675 3665 57695 4015
rect 57735 3665 57755 4015
rect 58410 3665 58430 4015
rect 58470 3665 58490 4015
rect 58530 3665 58550 4015
rect 58590 3665 58610 4015
rect 58650 3665 58670 4015
rect 58710 3665 58730 4015
rect 58770 3665 58790 4015
rect 58830 3665 58850 4015
rect 58890 3665 58910 4015
rect 58950 3665 58970 4015
rect 59010 3665 59030 4015
rect 59070 3665 59090 4015
rect 54740 2555 54755 3155
rect 54795 2555 54810 3155
rect 54850 2555 54865 3155
rect 54905 2555 54920 3155
rect 54960 2555 54975 3155
rect 55015 2555 55030 3155
rect 55070 2555 55085 3155
rect 55125 2555 55140 3155
rect 55180 2555 55195 3155
rect 55235 2555 55250 3155
rect 55290 2555 55305 3155
rect 55345 2555 55360 3155
rect 56550 2910 56565 3160
rect 56605 2910 56620 3160
rect 56660 2910 56675 3160
rect 56715 2910 56730 3160
rect 56770 2910 56785 3160
rect 56825 2910 56840 3160
rect 56960 2910 56975 3160
rect 57015 2910 57030 3160
rect 57070 2910 57085 3160
rect 57125 2910 57140 3160
rect 57180 2910 57195 3160
rect 57235 2910 57250 3160
rect 58440 2555 58455 3155
rect 58495 2555 58510 3155
rect 58550 2555 58565 3155
rect 58605 2555 58620 3155
rect 58660 2555 58675 3155
rect 58715 2555 58730 3155
rect 58770 2555 58785 3155
rect 58825 2555 58840 3155
rect 58880 2555 58895 3155
rect 58935 2555 58950 3155
rect 58990 2555 59005 3155
rect 59045 2555 59060 3155
rect 54740 1680 54755 1880
rect 54795 1680 54810 1880
rect 54850 1680 54865 1880
rect 54905 1680 54920 1880
rect 54960 1680 54975 1880
rect 55015 1680 55030 1880
rect 55070 1680 55085 1880
rect 55125 1680 55140 1880
rect 55180 1680 55195 1880
rect 55235 1680 55250 1880
rect 55290 1680 55305 1880
rect 55345 1680 55360 1880
rect 58440 1680 58455 1880
rect 58495 1680 58510 1880
rect 58550 1680 58565 1880
rect 58605 1680 58620 1880
rect 58660 1680 58675 1880
rect 58715 1680 58730 1880
rect 58770 1680 58785 1880
rect 58825 1680 58840 1880
rect 58880 1680 58895 1880
rect 58935 1680 58950 1880
rect 58990 1680 59005 1880
rect 59045 1680 59060 1880
<< ndiff >>
rect 56770 2550 56810 2565
rect 56770 2330 56780 2550
rect 56800 2330 56810 2550
rect 56770 2315 56810 2330
rect 56825 2550 56865 2565
rect 56825 2330 56835 2550
rect 56855 2330 56865 2550
rect 56825 2315 56865 2330
rect 56880 2550 56920 2565
rect 56880 2330 56890 2550
rect 56910 2330 56920 2550
rect 56880 2315 56920 2330
rect 56935 2550 56975 2565
rect 56935 2330 56945 2550
rect 56965 2330 56975 2550
rect 56935 2315 56975 2330
rect 56990 2550 57030 2565
rect 56990 2330 57000 2550
rect 57020 2330 57030 2550
rect 56990 2315 57030 2330
rect 56030 1880 56070 1895
rect 56030 1760 56040 1880
rect 56060 1760 56070 1880
rect 56030 1745 56070 1760
rect 56085 1880 56125 1895
rect 56085 1760 56095 1880
rect 56115 1760 56125 1880
rect 56085 1745 56125 1760
rect 56140 1880 56180 1895
rect 56140 1760 56150 1880
rect 56170 1760 56180 1880
rect 56140 1745 56180 1760
rect 56195 1880 56235 1895
rect 56195 1760 56205 1880
rect 56225 1760 56235 1880
rect 56195 1745 56235 1760
rect 56250 1880 56290 1895
rect 56250 1760 56260 1880
rect 56280 1760 56290 1880
rect 56250 1745 56290 1760
rect 56305 1880 56345 1895
rect 56305 1760 56315 1880
rect 56335 1760 56345 1880
rect 56305 1745 56345 1760
rect 56360 1880 56400 1895
rect 56360 1760 56370 1880
rect 56390 1760 56400 1880
rect 56360 1745 56400 1760
rect 56415 1880 56455 1895
rect 56415 1760 56425 1880
rect 56445 1760 56455 1880
rect 56415 1745 56455 1760
rect 56470 1880 56510 1895
rect 56470 1760 56480 1880
rect 56500 1760 56510 1880
rect 56470 1745 56510 1760
rect 56525 1880 56565 1895
rect 56525 1760 56535 1880
rect 56555 1760 56565 1880
rect 56525 1745 56565 1760
rect 56580 1880 56620 1895
rect 56580 1760 56590 1880
rect 56610 1760 56620 1880
rect 56580 1745 56620 1760
rect 56635 1880 56675 1895
rect 56635 1760 56645 1880
rect 56665 1760 56675 1880
rect 56635 1745 56675 1760
rect 56690 1880 56730 1895
rect 56690 1760 56700 1880
rect 56720 1760 56730 1880
rect 56690 1745 56730 1760
rect 57070 1880 57110 1895
rect 57070 1760 57080 1880
rect 57100 1760 57110 1880
rect 57070 1745 57110 1760
rect 57125 1880 57165 1895
rect 57125 1760 57135 1880
rect 57155 1760 57165 1880
rect 57125 1745 57165 1760
rect 57180 1880 57220 1895
rect 57180 1760 57190 1880
rect 57210 1760 57220 1880
rect 57180 1745 57220 1760
rect 57235 1880 57275 1895
rect 57235 1760 57245 1880
rect 57265 1760 57275 1880
rect 57235 1745 57275 1760
rect 57290 1880 57330 1895
rect 57290 1760 57300 1880
rect 57320 1760 57330 1880
rect 57290 1745 57330 1760
rect 57345 1880 57385 1895
rect 57345 1760 57355 1880
rect 57375 1760 57385 1880
rect 57345 1745 57385 1760
rect 57400 1880 57440 1895
rect 57400 1760 57410 1880
rect 57430 1760 57440 1880
rect 57400 1745 57440 1760
rect 57455 1880 57495 1895
rect 57455 1760 57465 1880
rect 57485 1760 57495 1880
rect 57455 1745 57495 1760
rect 57510 1880 57550 1895
rect 57510 1760 57520 1880
rect 57540 1760 57550 1880
rect 57510 1745 57550 1760
rect 57565 1880 57605 1895
rect 57565 1760 57575 1880
rect 57595 1760 57605 1880
rect 57565 1745 57605 1760
rect 57620 1880 57660 1895
rect 57620 1760 57630 1880
rect 57650 1760 57660 1880
rect 57620 1745 57660 1760
rect 57675 1880 57715 1895
rect 57675 1760 57685 1880
rect 57705 1760 57715 1880
rect 57675 1745 57715 1760
rect 57730 1880 57770 1895
rect 57730 1760 57740 1880
rect 57760 1760 57770 1880
rect 57730 1745 57770 1760
rect 54700 1425 54740 1440
rect 54700 1155 54710 1425
rect 54730 1155 54740 1425
rect 54700 1140 54740 1155
rect 54755 1425 54795 1440
rect 54755 1155 54765 1425
rect 54785 1155 54795 1425
rect 54755 1140 54795 1155
rect 54810 1425 54850 1440
rect 54810 1155 54820 1425
rect 54840 1155 54850 1425
rect 54810 1140 54850 1155
rect 54865 1425 54905 1440
rect 54865 1155 54875 1425
rect 54895 1155 54905 1425
rect 54865 1140 54905 1155
rect 54920 1425 54960 1440
rect 54920 1155 54930 1425
rect 54950 1155 54960 1425
rect 54920 1140 54960 1155
rect 54975 1425 55015 1440
rect 54975 1155 54985 1425
rect 55005 1155 55015 1425
rect 54975 1140 55015 1155
rect 55030 1425 55070 1440
rect 55030 1155 55040 1425
rect 55060 1155 55070 1425
rect 55030 1140 55070 1155
rect 55085 1425 55125 1440
rect 55085 1155 55095 1425
rect 55115 1155 55125 1425
rect 55085 1140 55125 1155
rect 55140 1425 55180 1440
rect 55140 1155 55150 1425
rect 55170 1155 55180 1425
rect 55140 1140 55180 1155
rect 55195 1425 55235 1440
rect 55195 1155 55205 1425
rect 55225 1155 55235 1425
rect 55195 1140 55235 1155
rect 55250 1425 55290 1440
rect 55250 1155 55260 1425
rect 55280 1155 55290 1425
rect 55250 1140 55290 1155
rect 55305 1425 55345 1440
rect 55305 1155 55315 1425
rect 55335 1155 55345 1425
rect 55305 1140 55345 1155
rect 55360 1425 55400 1440
rect 55360 1155 55370 1425
rect 55390 1155 55400 1425
rect 58400 1425 58440 1440
rect 55360 1140 55400 1155
rect 56030 1205 56070 1220
rect 56030 1085 56040 1205
rect 56060 1085 56070 1205
rect 56030 1070 56070 1085
rect 56085 1205 56125 1220
rect 56085 1085 56095 1205
rect 56115 1085 56125 1205
rect 56085 1070 56125 1085
rect 56140 1205 56180 1220
rect 56140 1085 56150 1205
rect 56170 1085 56180 1205
rect 56140 1070 56180 1085
rect 56195 1205 56235 1220
rect 56195 1085 56205 1205
rect 56225 1085 56235 1205
rect 56195 1070 56235 1085
rect 56250 1205 56290 1220
rect 56250 1085 56260 1205
rect 56280 1085 56290 1205
rect 56250 1070 56290 1085
rect 56305 1205 56345 1220
rect 56305 1085 56315 1205
rect 56335 1085 56345 1205
rect 56305 1070 56345 1085
rect 56360 1205 56400 1220
rect 56360 1085 56370 1205
rect 56390 1085 56400 1205
rect 56360 1070 56400 1085
rect 56415 1205 56455 1220
rect 56415 1085 56425 1205
rect 56445 1085 56455 1205
rect 56415 1070 56455 1085
rect 56470 1205 56510 1220
rect 56470 1085 56480 1205
rect 56500 1085 56510 1205
rect 56470 1070 56510 1085
rect 56525 1205 56565 1220
rect 56525 1085 56535 1205
rect 56555 1085 56565 1205
rect 56525 1070 56565 1085
rect 56580 1205 56620 1220
rect 56580 1085 56590 1205
rect 56610 1085 56620 1205
rect 56580 1070 56620 1085
rect 56635 1205 56675 1220
rect 56635 1085 56645 1205
rect 56665 1085 56675 1205
rect 56635 1070 56675 1085
rect 56690 1205 56730 1220
rect 56770 1205 56810 1220
rect 56690 1085 56700 1205
rect 56720 1085 56730 1205
rect 56770 1085 56780 1205
rect 56800 1085 56810 1205
rect 56690 1070 56730 1085
rect 56770 1070 56810 1085
rect 56825 1205 56865 1220
rect 56825 1085 56835 1205
rect 56855 1085 56865 1205
rect 56825 1070 56865 1085
rect 56880 1205 56920 1220
rect 56880 1085 56890 1205
rect 56910 1085 56920 1205
rect 56880 1070 56920 1085
rect 56935 1205 56975 1220
rect 56935 1085 56945 1205
rect 56965 1085 56975 1205
rect 56935 1070 56975 1085
rect 56990 1205 57030 1220
rect 57070 1205 57110 1220
rect 56990 1085 57000 1205
rect 57020 1085 57030 1205
rect 57070 1085 57080 1205
rect 57100 1085 57110 1205
rect 56990 1070 57030 1085
rect 57070 1070 57110 1085
rect 57125 1205 57165 1220
rect 57125 1085 57135 1205
rect 57155 1085 57165 1205
rect 57125 1070 57165 1085
rect 57180 1205 57220 1220
rect 57180 1085 57190 1205
rect 57210 1085 57220 1205
rect 57180 1070 57220 1085
rect 57235 1205 57275 1220
rect 57235 1085 57245 1205
rect 57265 1085 57275 1205
rect 57235 1070 57275 1085
rect 57290 1205 57330 1220
rect 57290 1085 57300 1205
rect 57320 1085 57330 1205
rect 57290 1070 57330 1085
rect 57345 1205 57385 1220
rect 57345 1085 57355 1205
rect 57375 1085 57385 1205
rect 57345 1070 57385 1085
rect 57400 1205 57440 1220
rect 57400 1085 57410 1205
rect 57430 1085 57440 1205
rect 57400 1070 57440 1085
rect 57455 1205 57495 1220
rect 57455 1085 57465 1205
rect 57485 1085 57495 1205
rect 57455 1070 57495 1085
rect 57510 1205 57550 1220
rect 57510 1085 57520 1205
rect 57540 1085 57550 1205
rect 57510 1070 57550 1085
rect 57565 1205 57605 1220
rect 57565 1085 57575 1205
rect 57595 1085 57605 1205
rect 57565 1070 57605 1085
rect 57620 1205 57660 1220
rect 57620 1085 57630 1205
rect 57650 1085 57660 1205
rect 57620 1070 57660 1085
rect 57675 1205 57715 1220
rect 57675 1085 57685 1205
rect 57705 1085 57715 1205
rect 57675 1070 57715 1085
rect 57730 1205 57770 1220
rect 57730 1085 57740 1205
rect 57760 1085 57770 1205
rect 58400 1155 58410 1425
rect 58430 1155 58440 1425
rect 58400 1140 58440 1155
rect 58455 1425 58495 1440
rect 58455 1155 58465 1425
rect 58485 1155 58495 1425
rect 58455 1140 58495 1155
rect 58510 1425 58550 1440
rect 58510 1155 58520 1425
rect 58540 1155 58550 1425
rect 58510 1140 58550 1155
rect 58565 1425 58605 1440
rect 58565 1155 58575 1425
rect 58595 1155 58605 1425
rect 58565 1140 58605 1155
rect 58620 1425 58660 1440
rect 58620 1155 58630 1425
rect 58650 1155 58660 1425
rect 58620 1140 58660 1155
rect 58675 1425 58715 1440
rect 58675 1155 58685 1425
rect 58705 1155 58715 1425
rect 58675 1140 58715 1155
rect 58730 1425 58770 1440
rect 58730 1155 58740 1425
rect 58760 1155 58770 1425
rect 58730 1140 58770 1155
rect 58785 1425 58825 1440
rect 58785 1155 58795 1425
rect 58815 1155 58825 1425
rect 58785 1140 58825 1155
rect 58840 1425 58880 1440
rect 58840 1155 58850 1425
rect 58870 1155 58880 1425
rect 58840 1140 58880 1155
rect 58895 1425 58935 1440
rect 58895 1155 58905 1425
rect 58925 1155 58935 1425
rect 58895 1140 58935 1155
rect 58950 1425 58990 1440
rect 58950 1155 58960 1425
rect 58980 1155 58990 1425
rect 58950 1140 58990 1155
rect 59005 1425 59045 1440
rect 59005 1155 59015 1425
rect 59035 1155 59045 1425
rect 59005 1140 59045 1155
rect 59060 1425 59100 1440
rect 59060 1155 59070 1425
rect 59090 1155 59100 1425
rect 59060 1140 59100 1155
rect 57730 1070 57770 1085
rect 56220 315 56260 330
rect 54730 165 54770 180
rect 54730 -505 54740 165
rect 54760 -505 54770 165
rect 54730 -520 54770 -505
rect 54830 165 54870 180
rect 54830 -505 54840 165
rect 54860 -505 54870 165
rect 54830 -520 54870 -505
rect 54930 165 54970 180
rect 54930 -505 54940 165
rect 54960 -505 54970 165
rect 54930 -520 54970 -505
rect 55030 165 55070 180
rect 55030 -505 55040 165
rect 55060 -505 55070 165
rect 55030 -520 55070 -505
rect 55130 165 55170 180
rect 55130 -505 55140 165
rect 55160 -505 55170 165
rect 55130 -520 55170 -505
rect 55230 165 55270 180
rect 55230 -505 55240 165
rect 55260 -505 55270 165
rect 55230 -520 55270 -505
rect 55330 165 55370 180
rect 55330 -505 55340 165
rect 55360 -505 55370 165
rect 56220 95 56230 315
rect 56250 95 56260 315
rect 56220 80 56260 95
rect 56275 315 56315 330
rect 56275 95 56285 315
rect 56305 95 56315 315
rect 56275 80 56315 95
rect 56330 315 56370 330
rect 56330 95 56340 315
rect 56360 95 56370 315
rect 56330 80 56370 95
rect 56385 315 56425 330
rect 56385 95 56395 315
rect 56415 95 56425 315
rect 56385 80 56425 95
rect 56440 315 56480 330
rect 56440 95 56450 315
rect 56470 95 56480 315
rect 56440 80 56480 95
rect 56495 315 56535 330
rect 56495 95 56505 315
rect 56525 95 56535 315
rect 56495 80 56535 95
rect 56550 315 56590 330
rect 56550 95 56560 315
rect 56580 95 56590 315
rect 56550 80 56590 95
rect 56605 315 56645 330
rect 56605 95 56615 315
rect 56635 95 56645 315
rect 56605 80 56645 95
rect 56660 315 56700 330
rect 56660 95 56670 315
rect 56690 95 56700 315
rect 56660 80 56700 95
rect 56715 315 56755 330
rect 56715 95 56725 315
rect 56745 95 56755 315
rect 56715 80 56755 95
rect 56770 315 56810 330
rect 56770 95 56780 315
rect 56800 95 56810 315
rect 56770 80 56810 95
rect 56825 315 56865 330
rect 56825 95 56835 315
rect 56855 95 56865 315
rect 56825 80 56865 95
rect 56880 315 56920 330
rect 56880 95 56890 315
rect 56910 95 56920 315
rect 56880 80 56920 95
rect 56935 315 56975 330
rect 56935 95 56945 315
rect 56965 95 56975 315
rect 56935 80 56975 95
rect 56990 315 57030 330
rect 56990 95 57000 315
rect 57020 95 57030 315
rect 56990 80 57030 95
rect 57045 315 57085 330
rect 57045 95 57055 315
rect 57075 95 57085 315
rect 57045 80 57085 95
rect 57100 315 57140 330
rect 57100 95 57110 315
rect 57130 95 57140 315
rect 57100 80 57140 95
rect 57155 315 57195 330
rect 57155 95 57165 315
rect 57185 95 57195 315
rect 57155 80 57195 95
rect 57210 315 57250 330
rect 57210 95 57220 315
rect 57240 95 57250 315
rect 57210 80 57250 95
rect 57265 315 57305 330
rect 57265 95 57275 315
rect 57295 95 57305 315
rect 57265 80 57305 95
rect 57320 315 57360 330
rect 57320 95 57330 315
rect 57350 95 57360 315
rect 57320 80 57360 95
rect 57375 315 57415 330
rect 57375 95 57385 315
rect 57405 95 57415 315
rect 57375 80 57415 95
rect 57430 315 57470 330
rect 57430 95 57440 315
rect 57460 95 57470 315
rect 57430 80 57470 95
rect 57485 315 57525 330
rect 57485 95 57495 315
rect 57515 95 57525 315
rect 57485 80 57525 95
rect 58430 165 58470 180
rect 56430 -340 56470 -325
rect 56430 -460 56440 -340
rect 56460 -460 56470 -340
rect 56430 -475 56470 -460
rect 56485 -340 56525 -325
rect 56485 -460 56495 -340
rect 56515 -460 56525 -340
rect 56485 -475 56525 -460
rect 56540 -340 56580 -325
rect 56540 -460 56550 -340
rect 56570 -460 56580 -340
rect 56540 -475 56580 -460
rect 56595 -340 56635 -325
rect 56595 -460 56605 -340
rect 56625 -460 56635 -340
rect 56595 -475 56635 -460
rect 56650 -340 56690 -325
rect 56650 -460 56660 -340
rect 56680 -460 56690 -340
rect 56650 -475 56690 -460
rect 56705 -340 56745 -325
rect 56705 -460 56715 -340
rect 56735 -460 56745 -340
rect 56705 -475 56745 -460
rect 56760 -340 56800 -325
rect 56760 -460 56770 -340
rect 56790 -460 56800 -340
rect 56760 -475 56800 -460
rect 56870 -340 56910 -325
rect 56870 -460 56880 -340
rect 56900 -460 56910 -340
rect 56870 -475 56910 -460
rect 57210 -340 57250 -325
rect 57210 -460 57220 -340
rect 57240 -460 57250 -340
rect 57210 -475 57250 -460
rect 55330 -520 55370 -505
rect 58430 -505 58440 165
rect 58460 -505 58470 165
rect 58430 -520 58470 -505
rect 58530 165 58570 180
rect 58530 -505 58540 165
rect 58560 -505 58570 165
rect 58530 -520 58570 -505
rect 58630 165 58670 180
rect 58630 -505 58640 165
rect 58660 -505 58670 165
rect 58630 -520 58670 -505
rect 58730 165 58770 180
rect 58730 -505 58740 165
rect 58760 -505 58770 165
rect 58730 -520 58770 -505
rect 58830 165 58870 180
rect 58830 -505 58840 165
rect 58860 -505 58870 165
rect 58830 -520 58870 -505
rect 58930 165 58970 180
rect 58930 -505 58940 165
rect 58960 -505 58970 165
rect 58930 -520 58970 -505
rect 59030 165 59070 180
rect 59030 -505 59040 165
rect 59060 -505 59070 165
rect 59030 -520 59070 -505
<< pdiff >>
rect 56085 4865 56125 4880
rect 56085 4545 56095 4865
rect 56115 4545 56125 4865
rect 56085 4530 56125 4545
rect 56145 4865 56185 4880
rect 56145 4545 56155 4865
rect 56175 4545 56185 4865
rect 56145 4530 56185 4545
rect 56205 4865 56245 4880
rect 56205 4545 56215 4865
rect 56235 4545 56245 4865
rect 56205 4530 56245 4545
rect 56265 4865 56305 4880
rect 56265 4545 56275 4865
rect 56295 4545 56305 4865
rect 57025 4865 57065 4880
rect 56265 4530 56305 4545
rect 56555 4695 56595 4710
rect 56555 4545 56565 4695
rect 56585 4545 56595 4695
rect 56555 4530 56595 4545
rect 56615 4695 56655 4710
rect 56615 4545 56625 4695
rect 56645 4545 56655 4695
rect 56615 4530 56655 4545
rect 56675 4695 56715 4710
rect 56675 4545 56685 4695
rect 56705 4545 56715 4695
rect 56675 4530 56715 4545
rect 56735 4695 56775 4710
rect 56735 4545 56745 4695
rect 56765 4545 56775 4695
rect 56735 4530 56775 4545
rect 57025 4545 57035 4865
rect 57055 4545 57065 4865
rect 57025 4530 57065 4545
rect 57085 4865 57125 4880
rect 57085 4545 57095 4865
rect 57115 4545 57125 4865
rect 57085 4530 57125 4545
rect 57145 4865 57185 4880
rect 57145 4545 57155 4865
rect 57175 4545 57185 4865
rect 57145 4530 57185 4545
rect 57205 4865 57245 4880
rect 57205 4545 57215 4865
rect 57235 4545 57245 4865
rect 57205 4530 57245 4545
rect 57495 4865 57535 4880
rect 57495 4545 57505 4865
rect 57525 4545 57535 4865
rect 57495 4530 57535 4545
rect 57555 4865 57595 4880
rect 57555 4545 57565 4865
rect 57585 4545 57595 4865
rect 57555 4530 57595 4545
rect 57615 4865 57655 4880
rect 57615 4545 57625 4865
rect 57645 4545 57655 4865
rect 57615 4530 57655 4545
rect 57675 4865 57715 4880
rect 57675 4545 57685 4865
rect 57705 4545 57715 4865
rect 57675 4530 57715 4545
rect 54670 4000 54710 4015
rect 54670 3680 54680 4000
rect 54700 3680 54710 4000
rect 54670 3665 54710 3680
rect 54730 4000 54770 4015
rect 54730 3680 54740 4000
rect 54760 3680 54770 4000
rect 54730 3665 54770 3680
rect 54790 4000 54830 4015
rect 54790 3680 54800 4000
rect 54820 3680 54830 4000
rect 54790 3665 54830 3680
rect 54850 4000 54890 4015
rect 54850 3680 54860 4000
rect 54880 3680 54890 4000
rect 54850 3665 54890 3680
rect 54910 4000 54950 4015
rect 54910 3680 54920 4000
rect 54940 3680 54950 4000
rect 54910 3665 54950 3680
rect 54970 4000 55010 4015
rect 54970 3680 54980 4000
rect 55000 3680 55010 4000
rect 54970 3665 55010 3680
rect 55030 4000 55070 4015
rect 55030 3680 55040 4000
rect 55060 3680 55070 4000
rect 55030 3665 55070 3680
rect 55090 4000 55130 4015
rect 55090 3680 55100 4000
rect 55120 3680 55130 4000
rect 55090 3665 55130 3680
rect 55150 4000 55190 4015
rect 55150 3680 55160 4000
rect 55180 3680 55190 4000
rect 55150 3665 55190 3680
rect 55210 4000 55250 4015
rect 55210 3680 55220 4000
rect 55240 3680 55250 4000
rect 55210 3665 55250 3680
rect 55270 4000 55310 4015
rect 55270 3680 55280 4000
rect 55300 3680 55310 4000
rect 55270 3665 55310 3680
rect 55330 4000 55370 4015
rect 55330 3680 55340 4000
rect 55360 3680 55370 4000
rect 55330 3665 55370 3680
rect 55390 4000 55430 4015
rect 55390 3680 55400 4000
rect 55420 3680 55430 4000
rect 55390 3665 55430 3680
rect 56005 4000 56045 4015
rect 56005 3680 56015 4000
rect 56035 3680 56045 4000
rect 56005 3665 56045 3680
rect 56065 4000 56105 4015
rect 56065 3680 56075 4000
rect 56095 3680 56105 4000
rect 56065 3665 56105 3680
rect 56125 4000 56165 4015
rect 56125 3680 56135 4000
rect 56155 3680 56165 4000
rect 56125 3665 56165 3680
rect 56185 4000 56225 4015
rect 56185 3680 56195 4000
rect 56215 3680 56225 4000
rect 56185 3665 56225 3680
rect 56245 4000 56285 4015
rect 56245 3680 56255 4000
rect 56275 3680 56285 4000
rect 56245 3665 56285 3680
rect 56305 4000 56345 4015
rect 56305 3680 56315 4000
rect 56335 3680 56345 4000
rect 56305 3665 56345 3680
rect 56365 4000 56405 4015
rect 56365 3680 56375 4000
rect 56395 3680 56405 4000
rect 56365 3665 56405 3680
rect 56425 4000 56465 4015
rect 56425 3680 56435 4000
rect 56455 3680 56465 4000
rect 56425 3665 56465 3680
rect 56485 4000 56525 4015
rect 56485 3680 56495 4000
rect 56515 3680 56525 4000
rect 56485 3665 56525 3680
rect 56545 4000 56585 4015
rect 56545 3680 56555 4000
rect 56575 3680 56585 4000
rect 56545 3665 56585 3680
rect 56605 4000 56645 4015
rect 56605 3680 56615 4000
rect 56635 3680 56645 4000
rect 56605 3665 56645 3680
rect 56665 4000 56705 4015
rect 56665 3680 56675 4000
rect 56695 3680 56705 4000
rect 56665 3665 56705 3680
rect 56725 4000 56765 4015
rect 56725 3680 56735 4000
rect 56755 3680 56765 4000
rect 56725 3665 56765 3680
rect 57035 4000 57075 4015
rect 57035 3680 57045 4000
rect 57065 3680 57075 4000
rect 57035 3665 57075 3680
rect 57095 4000 57135 4015
rect 57095 3680 57105 4000
rect 57125 3680 57135 4000
rect 57095 3665 57135 3680
rect 57155 4000 57195 4015
rect 57155 3680 57165 4000
rect 57185 3680 57195 4000
rect 57155 3665 57195 3680
rect 57215 4000 57255 4015
rect 57215 3680 57225 4000
rect 57245 3680 57255 4000
rect 57215 3665 57255 3680
rect 57275 4000 57315 4015
rect 57275 3680 57285 4000
rect 57305 3680 57315 4000
rect 57275 3665 57315 3680
rect 57335 4000 57375 4015
rect 57335 3680 57345 4000
rect 57365 3680 57375 4000
rect 57335 3665 57375 3680
rect 57395 4000 57435 4015
rect 57395 3680 57405 4000
rect 57425 3680 57435 4000
rect 57395 3665 57435 3680
rect 57455 4000 57495 4015
rect 57455 3680 57465 4000
rect 57485 3680 57495 4000
rect 57455 3665 57495 3680
rect 57515 4000 57555 4015
rect 57515 3680 57525 4000
rect 57545 3680 57555 4000
rect 57515 3665 57555 3680
rect 57575 4000 57615 4015
rect 57575 3680 57585 4000
rect 57605 3680 57615 4000
rect 57575 3665 57615 3680
rect 57635 4000 57675 4015
rect 57635 3680 57645 4000
rect 57665 3680 57675 4000
rect 57635 3665 57675 3680
rect 57695 4000 57735 4015
rect 57695 3680 57705 4000
rect 57725 3680 57735 4000
rect 57695 3665 57735 3680
rect 57755 4000 57795 4015
rect 57755 3680 57765 4000
rect 57785 3680 57795 4000
rect 57755 3665 57795 3680
rect 58370 4000 58410 4015
rect 58370 3680 58380 4000
rect 58400 3680 58410 4000
rect 58370 3665 58410 3680
rect 58430 4000 58470 4015
rect 58430 3680 58440 4000
rect 58460 3680 58470 4000
rect 58430 3665 58470 3680
rect 58490 4000 58530 4015
rect 58490 3680 58500 4000
rect 58520 3680 58530 4000
rect 58490 3665 58530 3680
rect 58550 4000 58590 4015
rect 58550 3680 58560 4000
rect 58580 3680 58590 4000
rect 58550 3665 58590 3680
rect 58610 4000 58650 4015
rect 58610 3680 58620 4000
rect 58640 3680 58650 4000
rect 58610 3665 58650 3680
rect 58670 4000 58710 4015
rect 58670 3680 58680 4000
rect 58700 3680 58710 4000
rect 58670 3665 58710 3680
rect 58730 4000 58770 4015
rect 58730 3680 58740 4000
rect 58760 3680 58770 4000
rect 58730 3665 58770 3680
rect 58790 4000 58830 4015
rect 58790 3680 58800 4000
rect 58820 3680 58830 4000
rect 58790 3665 58830 3680
rect 58850 4000 58890 4015
rect 58850 3680 58860 4000
rect 58880 3680 58890 4000
rect 58850 3665 58890 3680
rect 58910 4000 58950 4015
rect 58910 3680 58920 4000
rect 58940 3680 58950 4000
rect 58910 3665 58950 3680
rect 58970 4000 59010 4015
rect 58970 3680 58980 4000
rect 59000 3680 59010 4000
rect 58970 3665 59010 3680
rect 59030 4000 59070 4015
rect 59030 3680 59040 4000
rect 59060 3680 59070 4000
rect 59030 3665 59070 3680
rect 59090 4000 59130 4015
rect 59090 3680 59100 4000
rect 59120 3680 59130 4000
rect 59090 3665 59130 3680
rect 54700 3140 54740 3155
rect 54700 2570 54710 3140
rect 54730 2570 54740 3140
rect 54700 2555 54740 2570
rect 54755 3140 54795 3155
rect 54755 2570 54765 3140
rect 54785 2570 54795 3140
rect 54755 2555 54795 2570
rect 54810 3140 54850 3155
rect 54810 2570 54820 3140
rect 54840 2570 54850 3140
rect 54810 2555 54850 2570
rect 54865 3140 54905 3155
rect 54865 2570 54875 3140
rect 54895 2570 54905 3140
rect 54865 2555 54905 2570
rect 54920 3140 54960 3155
rect 54920 2570 54930 3140
rect 54950 2570 54960 3140
rect 54920 2555 54960 2570
rect 54975 3140 55015 3155
rect 54975 2570 54985 3140
rect 55005 2570 55015 3140
rect 54975 2555 55015 2570
rect 55030 3140 55070 3155
rect 55030 2570 55040 3140
rect 55060 2570 55070 3140
rect 55030 2555 55070 2570
rect 55085 3140 55125 3155
rect 55085 2570 55095 3140
rect 55115 2570 55125 3140
rect 55085 2555 55125 2570
rect 55140 3140 55180 3155
rect 55140 2570 55150 3140
rect 55170 2570 55180 3140
rect 55140 2555 55180 2570
rect 55195 3140 55235 3155
rect 55195 2570 55205 3140
rect 55225 2570 55235 3140
rect 55195 2555 55235 2570
rect 55250 3140 55290 3155
rect 55250 2570 55260 3140
rect 55280 2570 55290 3140
rect 55250 2555 55290 2570
rect 55305 3140 55345 3155
rect 55305 2570 55315 3140
rect 55335 2570 55345 3140
rect 55305 2555 55345 2570
rect 55360 3140 55400 3155
rect 55360 2570 55370 3140
rect 55390 2570 55400 3140
rect 56510 3145 56550 3160
rect 56510 3125 56520 3145
rect 56540 3125 56550 3145
rect 56510 3095 56550 3125
rect 56510 3075 56520 3095
rect 56540 3075 56550 3095
rect 56510 3045 56550 3075
rect 56510 3025 56520 3045
rect 56540 3025 56550 3045
rect 56510 2995 56550 3025
rect 56510 2975 56520 2995
rect 56540 2975 56550 2995
rect 56510 2945 56550 2975
rect 56510 2925 56520 2945
rect 56540 2925 56550 2945
rect 56510 2910 56550 2925
rect 56565 3145 56605 3160
rect 56565 3125 56575 3145
rect 56595 3125 56605 3145
rect 56565 3095 56605 3125
rect 56565 3075 56575 3095
rect 56595 3075 56605 3095
rect 56565 3045 56605 3075
rect 56565 3025 56575 3045
rect 56595 3025 56605 3045
rect 56565 2995 56605 3025
rect 56565 2975 56575 2995
rect 56595 2975 56605 2995
rect 56565 2945 56605 2975
rect 56565 2925 56575 2945
rect 56595 2925 56605 2945
rect 56565 2910 56605 2925
rect 56620 3145 56660 3160
rect 56620 3125 56630 3145
rect 56650 3125 56660 3145
rect 56620 3095 56660 3125
rect 56620 3075 56630 3095
rect 56650 3075 56660 3095
rect 56620 3045 56660 3075
rect 56620 3025 56630 3045
rect 56650 3025 56660 3045
rect 56620 2995 56660 3025
rect 56620 2975 56630 2995
rect 56650 2975 56660 2995
rect 56620 2945 56660 2975
rect 56620 2925 56630 2945
rect 56650 2925 56660 2945
rect 56620 2910 56660 2925
rect 56675 3145 56715 3160
rect 56675 3125 56685 3145
rect 56705 3125 56715 3145
rect 56675 3095 56715 3125
rect 56675 3075 56685 3095
rect 56705 3075 56715 3095
rect 56675 3045 56715 3075
rect 56675 3025 56685 3045
rect 56705 3025 56715 3045
rect 56675 2995 56715 3025
rect 56675 2975 56685 2995
rect 56705 2975 56715 2995
rect 56675 2945 56715 2975
rect 56675 2925 56685 2945
rect 56705 2925 56715 2945
rect 56675 2910 56715 2925
rect 56730 3145 56770 3160
rect 56730 3125 56740 3145
rect 56760 3125 56770 3145
rect 56730 3095 56770 3125
rect 56730 3075 56740 3095
rect 56760 3075 56770 3095
rect 56730 3045 56770 3075
rect 56730 3025 56740 3045
rect 56760 3025 56770 3045
rect 56730 2995 56770 3025
rect 56730 2975 56740 2995
rect 56760 2975 56770 2995
rect 56730 2945 56770 2975
rect 56730 2925 56740 2945
rect 56760 2925 56770 2945
rect 56730 2910 56770 2925
rect 56785 3145 56825 3160
rect 56785 3125 56795 3145
rect 56815 3125 56825 3145
rect 56785 3095 56825 3125
rect 56785 3075 56795 3095
rect 56815 3075 56825 3095
rect 56785 3045 56825 3075
rect 56785 3025 56795 3045
rect 56815 3025 56825 3045
rect 56785 2995 56825 3025
rect 56785 2975 56795 2995
rect 56815 2975 56825 2995
rect 56785 2945 56825 2975
rect 56785 2925 56795 2945
rect 56815 2925 56825 2945
rect 56785 2910 56825 2925
rect 56840 3145 56880 3160
rect 56920 3145 56960 3160
rect 56840 3125 56850 3145
rect 56870 3125 56880 3145
rect 56920 3125 56930 3145
rect 56950 3125 56960 3145
rect 56840 3095 56880 3125
rect 56920 3095 56960 3125
rect 56840 3075 56850 3095
rect 56870 3075 56880 3095
rect 56920 3075 56930 3095
rect 56950 3075 56960 3095
rect 56840 3045 56880 3075
rect 56920 3045 56960 3075
rect 56840 3025 56850 3045
rect 56870 3025 56880 3045
rect 56920 3025 56930 3045
rect 56950 3025 56960 3045
rect 56840 2995 56880 3025
rect 56920 2995 56960 3025
rect 56840 2975 56850 2995
rect 56870 2975 56880 2995
rect 56920 2975 56930 2995
rect 56950 2975 56960 2995
rect 56840 2945 56880 2975
rect 56920 2945 56960 2975
rect 56840 2925 56850 2945
rect 56870 2925 56880 2945
rect 56920 2925 56930 2945
rect 56950 2925 56960 2945
rect 56840 2910 56880 2925
rect 56920 2910 56960 2925
rect 56975 3145 57015 3160
rect 56975 3125 56985 3145
rect 57005 3125 57015 3145
rect 56975 3095 57015 3125
rect 56975 3075 56985 3095
rect 57005 3075 57015 3095
rect 56975 3045 57015 3075
rect 56975 3025 56985 3045
rect 57005 3025 57015 3045
rect 56975 2995 57015 3025
rect 56975 2975 56985 2995
rect 57005 2975 57015 2995
rect 56975 2945 57015 2975
rect 56975 2925 56985 2945
rect 57005 2925 57015 2945
rect 56975 2910 57015 2925
rect 57030 3145 57070 3160
rect 57030 3125 57040 3145
rect 57060 3125 57070 3145
rect 57030 3095 57070 3125
rect 57030 3075 57040 3095
rect 57060 3075 57070 3095
rect 57030 3045 57070 3075
rect 57030 3025 57040 3045
rect 57060 3025 57070 3045
rect 57030 2995 57070 3025
rect 57030 2975 57040 2995
rect 57060 2975 57070 2995
rect 57030 2945 57070 2975
rect 57030 2925 57040 2945
rect 57060 2925 57070 2945
rect 57030 2910 57070 2925
rect 57085 3145 57125 3160
rect 57085 3125 57095 3145
rect 57115 3125 57125 3145
rect 57085 3095 57125 3125
rect 57085 3075 57095 3095
rect 57115 3075 57125 3095
rect 57085 3045 57125 3075
rect 57085 3025 57095 3045
rect 57115 3025 57125 3045
rect 57085 2995 57125 3025
rect 57085 2975 57095 2995
rect 57115 2975 57125 2995
rect 57085 2945 57125 2975
rect 57085 2925 57095 2945
rect 57115 2925 57125 2945
rect 57085 2910 57125 2925
rect 57140 3145 57180 3160
rect 57140 3125 57150 3145
rect 57170 3125 57180 3145
rect 57140 3095 57180 3125
rect 57140 3075 57150 3095
rect 57170 3075 57180 3095
rect 57140 3045 57180 3075
rect 57140 3025 57150 3045
rect 57170 3025 57180 3045
rect 57140 2995 57180 3025
rect 57140 2975 57150 2995
rect 57170 2975 57180 2995
rect 57140 2945 57180 2975
rect 57140 2925 57150 2945
rect 57170 2925 57180 2945
rect 57140 2910 57180 2925
rect 57195 3145 57235 3160
rect 57195 3125 57205 3145
rect 57225 3125 57235 3145
rect 57195 3095 57235 3125
rect 57195 3075 57205 3095
rect 57225 3075 57235 3095
rect 57195 3045 57235 3075
rect 57195 3025 57205 3045
rect 57225 3025 57235 3045
rect 57195 2995 57235 3025
rect 57195 2975 57205 2995
rect 57225 2975 57235 2995
rect 57195 2945 57235 2975
rect 57195 2925 57205 2945
rect 57225 2925 57235 2945
rect 57195 2910 57235 2925
rect 57250 3145 57290 3160
rect 57250 3125 57260 3145
rect 57280 3125 57290 3145
rect 57250 3095 57290 3125
rect 57250 3075 57260 3095
rect 57280 3075 57290 3095
rect 57250 3045 57290 3075
rect 57250 3025 57260 3045
rect 57280 3025 57290 3045
rect 57250 2995 57290 3025
rect 57250 2975 57260 2995
rect 57280 2975 57290 2995
rect 57250 2945 57290 2975
rect 57250 2925 57260 2945
rect 57280 2925 57290 2945
rect 57250 2910 57290 2925
rect 58400 3140 58440 3155
rect 55360 2555 55400 2570
rect 58400 2570 58410 3140
rect 58430 2570 58440 3140
rect 58400 2555 58440 2570
rect 58455 3140 58495 3155
rect 58455 2570 58465 3140
rect 58485 2570 58495 3140
rect 58455 2555 58495 2570
rect 58510 3140 58550 3155
rect 58510 2570 58520 3140
rect 58540 2570 58550 3140
rect 58510 2555 58550 2570
rect 58565 3140 58605 3155
rect 58565 2570 58575 3140
rect 58595 2570 58605 3140
rect 58565 2555 58605 2570
rect 58620 3140 58660 3155
rect 58620 2570 58630 3140
rect 58650 2570 58660 3140
rect 58620 2555 58660 2570
rect 58675 3140 58715 3155
rect 58675 2570 58685 3140
rect 58705 2570 58715 3140
rect 58675 2555 58715 2570
rect 58730 3140 58770 3155
rect 58730 2570 58740 3140
rect 58760 2570 58770 3140
rect 58730 2555 58770 2570
rect 58785 3140 58825 3155
rect 58785 2570 58795 3140
rect 58815 2570 58825 3140
rect 58785 2555 58825 2570
rect 58840 3140 58880 3155
rect 58840 2570 58850 3140
rect 58870 2570 58880 3140
rect 58840 2555 58880 2570
rect 58895 3140 58935 3155
rect 58895 2570 58905 3140
rect 58925 2570 58935 3140
rect 58895 2555 58935 2570
rect 58950 3140 58990 3155
rect 58950 2570 58960 3140
rect 58980 2570 58990 3140
rect 58950 2555 58990 2570
rect 59005 3140 59045 3155
rect 59005 2570 59015 3140
rect 59035 2570 59045 3140
rect 59005 2555 59045 2570
rect 59060 3140 59100 3155
rect 59060 2570 59070 3140
rect 59090 2570 59100 3140
rect 59060 2555 59100 2570
rect 54700 1865 54740 1880
rect 54700 1695 54710 1865
rect 54730 1695 54740 1865
rect 54700 1680 54740 1695
rect 54755 1865 54795 1880
rect 54755 1695 54765 1865
rect 54785 1695 54795 1865
rect 54755 1680 54795 1695
rect 54810 1865 54850 1880
rect 54810 1695 54820 1865
rect 54840 1695 54850 1865
rect 54810 1680 54850 1695
rect 54865 1865 54905 1880
rect 54865 1695 54875 1865
rect 54895 1695 54905 1865
rect 54865 1680 54905 1695
rect 54920 1865 54960 1880
rect 54920 1695 54930 1865
rect 54950 1695 54960 1865
rect 54920 1680 54960 1695
rect 54975 1865 55015 1880
rect 54975 1695 54985 1865
rect 55005 1695 55015 1865
rect 54975 1680 55015 1695
rect 55030 1865 55070 1880
rect 55030 1695 55040 1865
rect 55060 1695 55070 1865
rect 55030 1680 55070 1695
rect 55085 1865 55125 1880
rect 55085 1695 55095 1865
rect 55115 1695 55125 1865
rect 55085 1680 55125 1695
rect 55140 1865 55180 1880
rect 55140 1695 55150 1865
rect 55170 1695 55180 1865
rect 55140 1680 55180 1695
rect 55195 1865 55235 1880
rect 55195 1695 55205 1865
rect 55225 1695 55235 1865
rect 55195 1680 55235 1695
rect 55250 1865 55290 1880
rect 55250 1695 55260 1865
rect 55280 1695 55290 1865
rect 55250 1680 55290 1695
rect 55305 1865 55345 1880
rect 55305 1695 55315 1865
rect 55335 1695 55345 1865
rect 55305 1680 55345 1695
rect 55360 1865 55400 1880
rect 55360 1695 55370 1865
rect 55390 1695 55400 1865
rect 58400 1865 58440 1880
rect 55360 1680 55400 1695
rect 58400 1695 58410 1865
rect 58430 1695 58440 1865
rect 58400 1680 58440 1695
rect 58455 1865 58495 1880
rect 58455 1695 58465 1865
rect 58485 1695 58495 1865
rect 58455 1680 58495 1695
rect 58510 1865 58550 1880
rect 58510 1695 58520 1865
rect 58540 1695 58550 1865
rect 58510 1680 58550 1695
rect 58565 1865 58605 1880
rect 58565 1695 58575 1865
rect 58595 1695 58605 1865
rect 58565 1680 58605 1695
rect 58620 1865 58660 1880
rect 58620 1695 58630 1865
rect 58650 1695 58660 1865
rect 58620 1680 58660 1695
rect 58675 1865 58715 1880
rect 58675 1695 58685 1865
rect 58705 1695 58715 1865
rect 58675 1680 58715 1695
rect 58730 1865 58770 1880
rect 58730 1695 58740 1865
rect 58760 1695 58770 1865
rect 58730 1680 58770 1695
rect 58785 1865 58825 1880
rect 58785 1695 58795 1865
rect 58815 1695 58825 1865
rect 58785 1680 58825 1695
rect 58840 1865 58880 1880
rect 58840 1695 58850 1865
rect 58870 1695 58880 1865
rect 58840 1680 58880 1695
rect 58895 1865 58935 1880
rect 58895 1695 58905 1865
rect 58925 1695 58935 1865
rect 58895 1680 58935 1695
rect 58950 1865 58990 1880
rect 58950 1695 58960 1865
rect 58980 1695 58990 1865
rect 58950 1680 58990 1695
rect 59005 1865 59045 1880
rect 59005 1695 59015 1865
rect 59035 1695 59045 1865
rect 59005 1680 59045 1695
rect 59060 1865 59100 1880
rect 59060 1695 59070 1865
rect 59090 1695 59100 1865
rect 59060 1680 59100 1695
<< ndiffc >>
rect 56780 2330 56800 2550
rect 56835 2330 56855 2550
rect 56890 2330 56910 2550
rect 56945 2330 56965 2550
rect 57000 2330 57020 2550
rect 56040 1760 56060 1880
rect 56095 1760 56115 1880
rect 56150 1760 56170 1880
rect 56205 1760 56225 1880
rect 56260 1760 56280 1880
rect 56315 1760 56335 1880
rect 56370 1760 56390 1880
rect 56425 1760 56445 1880
rect 56480 1760 56500 1880
rect 56535 1760 56555 1880
rect 56590 1760 56610 1880
rect 56645 1760 56665 1880
rect 56700 1760 56720 1880
rect 57080 1760 57100 1880
rect 57135 1760 57155 1880
rect 57190 1760 57210 1880
rect 57245 1760 57265 1880
rect 57300 1760 57320 1880
rect 57355 1760 57375 1880
rect 57410 1760 57430 1880
rect 57465 1760 57485 1880
rect 57520 1760 57540 1880
rect 57575 1760 57595 1880
rect 57630 1760 57650 1880
rect 57685 1760 57705 1880
rect 57740 1760 57760 1880
rect 54710 1155 54730 1425
rect 54765 1155 54785 1425
rect 54820 1155 54840 1425
rect 54875 1155 54895 1425
rect 54930 1155 54950 1425
rect 54985 1155 55005 1425
rect 55040 1155 55060 1425
rect 55095 1155 55115 1425
rect 55150 1155 55170 1425
rect 55205 1155 55225 1425
rect 55260 1155 55280 1425
rect 55315 1155 55335 1425
rect 55370 1155 55390 1425
rect 56040 1085 56060 1205
rect 56095 1085 56115 1205
rect 56150 1085 56170 1205
rect 56205 1085 56225 1205
rect 56260 1085 56280 1205
rect 56315 1085 56335 1205
rect 56370 1085 56390 1205
rect 56425 1085 56445 1205
rect 56480 1085 56500 1205
rect 56535 1085 56555 1205
rect 56590 1085 56610 1205
rect 56645 1085 56665 1205
rect 56700 1085 56720 1205
rect 56780 1085 56800 1205
rect 56835 1085 56855 1205
rect 56890 1085 56910 1205
rect 56945 1085 56965 1205
rect 57000 1085 57020 1205
rect 57080 1085 57100 1205
rect 57135 1085 57155 1205
rect 57190 1085 57210 1205
rect 57245 1085 57265 1205
rect 57300 1085 57320 1205
rect 57355 1085 57375 1205
rect 57410 1085 57430 1205
rect 57465 1085 57485 1205
rect 57520 1085 57540 1205
rect 57575 1085 57595 1205
rect 57630 1085 57650 1205
rect 57685 1085 57705 1205
rect 57740 1085 57760 1205
rect 58410 1155 58430 1425
rect 58465 1155 58485 1425
rect 58520 1155 58540 1425
rect 58575 1155 58595 1425
rect 58630 1155 58650 1425
rect 58685 1155 58705 1425
rect 58740 1155 58760 1425
rect 58795 1155 58815 1425
rect 58850 1155 58870 1425
rect 58905 1155 58925 1425
rect 58960 1155 58980 1425
rect 59015 1155 59035 1425
rect 59070 1155 59090 1425
rect 54740 -505 54760 165
rect 54840 -505 54860 165
rect 54940 -505 54960 165
rect 55040 -505 55060 165
rect 55140 -505 55160 165
rect 55240 -505 55260 165
rect 55340 -505 55360 165
rect 56230 95 56250 315
rect 56285 95 56305 315
rect 56340 95 56360 315
rect 56395 95 56415 315
rect 56450 95 56470 315
rect 56505 95 56525 315
rect 56560 95 56580 315
rect 56615 95 56635 315
rect 56670 95 56690 315
rect 56725 95 56745 315
rect 56780 95 56800 315
rect 56835 95 56855 315
rect 56890 95 56910 315
rect 56945 95 56965 315
rect 57000 95 57020 315
rect 57055 95 57075 315
rect 57110 95 57130 315
rect 57165 95 57185 315
rect 57220 95 57240 315
rect 57275 95 57295 315
rect 57330 95 57350 315
rect 57385 95 57405 315
rect 57440 95 57460 315
rect 57495 95 57515 315
rect 56440 -460 56460 -340
rect 56495 -460 56515 -340
rect 56550 -460 56570 -340
rect 56605 -460 56625 -340
rect 56660 -460 56680 -340
rect 56715 -460 56735 -340
rect 56770 -460 56790 -340
rect 56880 -460 56900 -340
rect 57220 -460 57240 -340
rect 58440 -505 58460 165
rect 58540 -505 58560 165
rect 58640 -505 58660 165
rect 58740 -505 58760 165
rect 58840 -505 58860 165
rect 58940 -505 58960 165
rect 59040 -505 59060 165
<< pdiffc >>
rect 56095 4545 56115 4865
rect 56155 4545 56175 4865
rect 56215 4545 56235 4865
rect 56275 4545 56295 4865
rect 56565 4545 56585 4695
rect 56625 4545 56645 4695
rect 56685 4545 56705 4695
rect 56745 4545 56765 4695
rect 57035 4545 57055 4865
rect 57095 4545 57115 4865
rect 57155 4545 57175 4865
rect 57215 4545 57235 4865
rect 57505 4545 57525 4865
rect 57565 4545 57585 4865
rect 57625 4545 57645 4865
rect 57685 4545 57705 4865
rect 54680 3680 54700 4000
rect 54740 3680 54760 4000
rect 54800 3680 54820 4000
rect 54860 3680 54880 4000
rect 54920 3680 54940 4000
rect 54980 3680 55000 4000
rect 55040 3680 55060 4000
rect 55100 3680 55120 4000
rect 55160 3680 55180 4000
rect 55220 3680 55240 4000
rect 55280 3680 55300 4000
rect 55340 3680 55360 4000
rect 55400 3680 55420 4000
rect 56015 3680 56035 4000
rect 56075 3680 56095 4000
rect 56135 3680 56155 4000
rect 56195 3680 56215 4000
rect 56255 3680 56275 4000
rect 56315 3680 56335 4000
rect 56375 3680 56395 4000
rect 56435 3680 56455 4000
rect 56495 3680 56515 4000
rect 56555 3680 56575 4000
rect 56615 3680 56635 4000
rect 56675 3680 56695 4000
rect 56735 3680 56755 4000
rect 57045 3680 57065 4000
rect 57105 3680 57125 4000
rect 57165 3680 57185 4000
rect 57225 3680 57245 4000
rect 57285 3680 57305 4000
rect 57345 3680 57365 4000
rect 57405 3680 57425 4000
rect 57465 3680 57485 4000
rect 57525 3680 57545 4000
rect 57585 3680 57605 4000
rect 57645 3680 57665 4000
rect 57705 3680 57725 4000
rect 57765 3680 57785 4000
rect 58380 3680 58400 4000
rect 58440 3680 58460 4000
rect 58500 3680 58520 4000
rect 58560 3680 58580 4000
rect 58620 3680 58640 4000
rect 58680 3680 58700 4000
rect 58740 3680 58760 4000
rect 58800 3680 58820 4000
rect 58860 3680 58880 4000
rect 58920 3680 58940 4000
rect 58980 3680 59000 4000
rect 59040 3680 59060 4000
rect 59100 3680 59120 4000
rect 54710 2570 54730 3140
rect 54765 2570 54785 3140
rect 54820 2570 54840 3140
rect 54875 2570 54895 3140
rect 54930 2570 54950 3140
rect 54985 2570 55005 3140
rect 55040 2570 55060 3140
rect 55095 2570 55115 3140
rect 55150 2570 55170 3140
rect 55205 2570 55225 3140
rect 55260 2570 55280 3140
rect 55315 2570 55335 3140
rect 55370 2570 55390 3140
rect 56520 3125 56540 3145
rect 56520 3075 56540 3095
rect 56520 3025 56540 3045
rect 56520 2975 56540 2995
rect 56520 2925 56540 2945
rect 56575 3125 56595 3145
rect 56575 3075 56595 3095
rect 56575 3025 56595 3045
rect 56575 2975 56595 2995
rect 56575 2925 56595 2945
rect 56630 3125 56650 3145
rect 56630 3075 56650 3095
rect 56630 3025 56650 3045
rect 56630 2975 56650 2995
rect 56630 2925 56650 2945
rect 56685 3125 56705 3145
rect 56685 3075 56705 3095
rect 56685 3025 56705 3045
rect 56685 2975 56705 2995
rect 56685 2925 56705 2945
rect 56740 3125 56760 3145
rect 56740 3075 56760 3095
rect 56740 3025 56760 3045
rect 56740 2975 56760 2995
rect 56740 2925 56760 2945
rect 56795 3125 56815 3145
rect 56795 3075 56815 3095
rect 56795 3025 56815 3045
rect 56795 2975 56815 2995
rect 56795 2925 56815 2945
rect 56850 3125 56870 3145
rect 56930 3125 56950 3145
rect 56850 3075 56870 3095
rect 56930 3075 56950 3095
rect 56850 3025 56870 3045
rect 56930 3025 56950 3045
rect 56850 2975 56870 2995
rect 56930 2975 56950 2995
rect 56850 2925 56870 2945
rect 56930 2925 56950 2945
rect 56985 3125 57005 3145
rect 56985 3075 57005 3095
rect 56985 3025 57005 3045
rect 56985 2975 57005 2995
rect 56985 2925 57005 2945
rect 57040 3125 57060 3145
rect 57040 3075 57060 3095
rect 57040 3025 57060 3045
rect 57040 2975 57060 2995
rect 57040 2925 57060 2945
rect 57095 3125 57115 3145
rect 57095 3075 57115 3095
rect 57095 3025 57115 3045
rect 57095 2975 57115 2995
rect 57095 2925 57115 2945
rect 57150 3125 57170 3145
rect 57150 3075 57170 3095
rect 57150 3025 57170 3045
rect 57150 2975 57170 2995
rect 57150 2925 57170 2945
rect 57205 3125 57225 3145
rect 57205 3075 57225 3095
rect 57205 3025 57225 3045
rect 57205 2975 57225 2995
rect 57205 2925 57225 2945
rect 57260 3125 57280 3145
rect 57260 3075 57280 3095
rect 57260 3025 57280 3045
rect 57260 2975 57280 2995
rect 57260 2925 57280 2945
rect 58410 2570 58430 3140
rect 58465 2570 58485 3140
rect 58520 2570 58540 3140
rect 58575 2570 58595 3140
rect 58630 2570 58650 3140
rect 58685 2570 58705 3140
rect 58740 2570 58760 3140
rect 58795 2570 58815 3140
rect 58850 2570 58870 3140
rect 58905 2570 58925 3140
rect 58960 2570 58980 3140
rect 59015 2570 59035 3140
rect 59070 2570 59090 3140
rect 54710 1695 54730 1865
rect 54765 1695 54785 1865
rect 54820 1695 54840 1865
rect 54875 1695 54895 1865
rect 54930 1695 54950 1865
rect 54985 1695 55005 1865
rect 55040 1695 55060 1865
rect 55095 1695 55115 1865
rect 55150 1695 55170 1865
rect 55205 1695 55225 1865
rect 55260 1695 55280 1865
rect 55315 1695 55335 1865
rect 55370 1695 55390 1865
rect 58410 1695 58430 1865
rect 58465 1695 58485 1865
rect 58520 1695 58540 1865
rect 58575 1695 58595 1865
rect 58630 1695 58650 1865
rect 58685 1695 58705 1865
rect 58740 1695 58760 1865
rect 58795 1695 58815 1865
rect 58850 1695 58870 1865
rect 58905 1695 58925 1865
rect 58960 1695 58980 1865
rect 59015 1695 59035 1865
rect 59070 1695 59090 1865
<< psubdiff >>
rect 56730 2550 56770 2565
rect 56730 2330 56740 2550
rect 56760 2330 56770 2550
rect 56730 2315 56770 2330
rect 57030 2550 57070 2565
rect 57030 2330 57040 2550
rect 57060 2330 57070 2550
rect 57030 2315 57070 2330
rect 55990 1880 56030 1895
rect 55990 1760 56000 1880
rect 56020 1760 56030 1880
rect 55990 1745 56030 1760
rect 56730 1880 56770 1895
rect 56730 1760 56740 1880
rect 56760 1760 56770 1880
rect 56730 1745 56770 1760
rect 57030 1880 57070 1895
rect 57030 1760 57040 1880
rect 57060 1760 57070 1880
rect 57030 1745 57070 1760
rect 57770 1880 57810 1895
rect 57770 1760 57780 1880
rect 57800 1760 57810 1880
rect 57770 1745 57810 1760
rect 54660 1425 54700 1440
rect 54660 1155 54670 1425
rect 54690 1155 54700 1425
rect 54660 1140 54700 1155
rect 55400 1425 55440 1440
rect 55400 1155 55410 1425
rect 55430 1155 55440 1425
rect 58360 1425 58400 1440
rect 55400 1140 55440 1155
rect 55990 1205 56030 1220
rect 55990 1085 56000 1205
rect 56020 1085 56030 1205
rect 55990 1070 56030 1085
rect 56730 1205 56770 1220
rect 56730 1085 56740 1205
rect 56760 1085 56770 1205
rect 56730 1070 56770 1085
rect 57030 1205 57070 1220
rect 57030 1085 57040 1205
rect 57060 1085 57070 1205
rect 57030 1070 57070 1085
rect 57770 1205 57810 1220
rect 57770 1085 57780 1205
rect 57800 1085 57810 1205
rect 58360 1155 58370 1425
rect 58390 1155 58400 1425
rect 58360 1140 58400 1155
rect 59100 1425 59140 1440
rect 59100 1155 59110 1425
rect 59130 1155 59140 1425
rect 59100 1140 59140 1155
rect 57770 1070 57810 1085
rect 56180 315 56220 330
rect 54690 165 54730 180
rect 54690 -505 54700 165
rect 54720 -505 54730 165
rect 54690 -520 54730 -505
rect 55370 165 55410 180
rect 55370 -505 55380 165
rect 55400 -505 55410 165
rect 56180 95 56190 315
rect 56210 95 56220 315
rect 56180 80 56220 95
rect 57525 315 57565 330
rect 57525 95 57535 315
rect 57555 95 57565 315
rect 57525 80 57565 95
rect 58390 165 58430 180
rect 56390 -340 56430 -325
rect 56390 -460 56400 -340
rect 56420 -460 56430 -340
rect 56390 -475 56430 -460
rect 56800 -340 56840 -325
rect 56800 -460 56810 -340
rect 56830 -460 56840 -340
rect 56800 -475 56840 -460
rect 55370 -520 55410 -505
rect 58390 -505 58400 165
rect 58420 -505 58430 165
rect 58390 -520 58430 -505
rect 59070 165 59110 180
rect 59070 -505 59080 165
rect 59100 -505 59110 165
rect 59070 -520 59110 -505
<< nsubdiff >>
rect 56045 4865 56085 4880
rect 56045 4545 56055 4865
rect 56075 4545 56085 4865
rect 56045 4530 56085 4545
rect 56305 4865 56345 4880
rect 56305 4545 56315 4865
rect 56335 4545 56345 4865
rect 56985 4865 57025 4880
rect 56305 4530 56345 4545
rect 56515 4695 56555 4710
rect 56515 4545 56525 4695
rect 56545 4545 56555 4695
rect 56515 4530 56555 4545
rect 56775 4695 56815 4710
rect 56775 4545 56785 4695
rect 56805 4545 56815 4695
rect 56775 4530 56815 4545
rect 56985 4545 56995 4865
rect 57015 4545 57025 4865
rect 56985 4530 57025 4545
rect 57245 4865 57285 4880
rect 57245 4545 57255 4865
rect 57275 4545 57285 4865
rect 57245 4530 57285 4545
rect 57455 4865 57495 4880
rect 57455 4545 57465 4865
rect 57485 4545 57495 4865
rect 57455 4530 57495 4545
rect 57715 4865 57755 4880
rect 57715 4545 57725 4865
rect 57745 4545 57755 4865
rect 57715 4530 57755 4545
rect 54630 4000 54670 4015
rect 54630 3680 54640 4000
rect 54660 3680 54670 4000
rect 54630 3665 54670 3680
rect 55430 4000 55470 4015
rect 55430 3680 55440 4000
rect 55460 3680 55470 4000
rect 55430 3665 55470 3680
rect 55965 4000 56005 4015
rect 55965 3680 55975 4000
rect 55995 3680 56005 4000
rect 55965 3665 56005 3680
rect 56765 4000 56805 4015
rect 56765 3680 56775 4000
rect 56795 3680 56805 4000
rect 56765 3665 56805 3680
rect 56995 4000 57035 4015
rect 56995 3680 57005 4000
rect 57025 3680 57035 4000
rect 56995 3665 57035 3680
rect 57795 4000 57835 4015
rect 57795 3680 57805 4000
rect 57825 3680 57835 4000
rect 57795 3665 57835 3680
rect 58330 4000 58370 4015
rect 58330 3680 58340 4000
rect 58360 3680 58370 4000
rect 58330 3665 58370 3680
rect 59130 4000 59170 4015
rect 59130 3680 59140 4000
rect 59160 3680 59170 4000
rect 59130 3665 59170 3680
rect 54660 3140 54700 3155
rect 54660 2570 54670 3140
rect 54690 2570 54700 3140
rect 54660 2555 54700 2570
rect 55400 3140 55440 3155
rect 55400 2570 55410 3140
rect 55430 2570 55440 3140
rect 56470 3145 56510 3160
rect 56470 3125 56480 3145
rect 56500 3125 56510 3145
rect 56470 3095 56510 3125
rect 56470 3075 56480 3095
rect 56500 3075 56510 3095
rect 56470 3045 56510 3075
rect 56470 3025 56480 3045
rect 56500 3025 56510 3045
rect 56470 2995 56510 3025
rect 56470 2975 56480 2995
rect 56500 2975 56510 2995
rect 56470 2945 56510 2975
rect 56470 2925 56480 2945
rect 56500 2925 56510 2945
rect 56470 2910 56510 2925
rect 56880 3145 56920 3160
rect 56880 3125 56890 3145
rect 56910 3125 56920 3145
rect 56880 3095 56920 3125
rect 56880 3075 56890 3095
rect 56910 3075 56920 3095
rect 56880 3045 56920 3075
rect 56880 3025 56890 3045
rect 56910 3025 56920 3045
rect 56880 2995 56920 3025
rect 56880 2975 56890 2995
rect 56910 2975 56920 2995
rect 56880 2945 56920 2975
rect 56880 2925 56890 2945
rect 56910 2925 56920 2945
rect 56880 2910 56920 2925
rect 57290 3145 57330 3160
rect 57290 3125 57300 3145
rect 57320 3125 57330 3145
rect 57290 3095 57330 3125
rect 57290 3075 57300 3095
rect 57320 3075 57330 3095
rect 57290 3045 57330 3075
rect 57290 3025 57300 3045
rect 57320 3025 57330 3045
rect 57290 2995 57330 3025
rect 57290 2975 57300 2995
rect 57320 2975 57330 2995
rect 57290 2945 57330 2975
rect 57290 2925 57300 2945
rect 57320 2925 57330 2945
rect 57290 2910 57330 2925
rect 58360 3140 58400 3155
rect 55400 2555 55440 2570
rect 58360 2570 58370 3140
rect 58390 2570 58400 3140
rect 58360 2555 58400 2570
rect 59100 3140 59140 3155
rect 59100 2570 59110 3140
rect 59130 2570 59140 3140
rect 59100 2555 59140 2570
rect 54660 1865 54700 1880
rect 54660 1695 54670 1865
rect 54690 1695 54700 1865
rect 54660 1680 54700 1695
rect 55400 1865 55440 1880
rect 55400 1695 55410 1865
rect 55430 1695 55440 1865
rect 58360 1865 58400 1880
rect 55400 1680 55440 1695
rect 58360 1695 58370 1865
rect 58390 1695 58400 1865
rect 58360 1680 58400 1695
rect 59100 1865 59140 1880
rect 59100 1695 59110 1865
rect 59130 1695 59140 1865
rect 59100 1680 59140 1695
<< psubdiffcont >>
rect 56740 2330 56760 2550
rect 57040 2330 57060 2550
rect 56000 1760 56020 1880
rect 56740 1760 56760 1880
rect 57040 1760 57060 1880
rect 57780 1760 57800 1880
rect 54670 1155 54690 1425
rect 55410 1155 55430 1425
rect 56000 1085 56020 1205
rect 56740 1085 56760 1205
rect 57040 1085 57060 1205
rect 57780 1085 57800 1205
rect 58370 1155 58390 1425
rect 59110 1155 59130 1425
rect 54700 -505 54720 165
rect 55380 -505 55400 165
rect 56190 95 56210 315
rect 57535 95 57555 315
rect 56400 -460 56420 -340
rect 56810 -460 56830 -340
rect 58400 -505 58420 165
rect 59080 -505 59100 165
<< nsubdiffcont >>
rect 56055 4545 56075 4865
rect 56315 4545 56335 4865
rect 56525 4545 56545 4695
rect 56785 4545 56805 4695
rect 56995 4545 57015 4865
rect 57255 4545 57275 4865
rect 57465 4545 57485 4865
rect 57725 4545 57745 4865
rect 54640 3680 54660 4000
rect 55440 3680 55460 4000
rect 55975 3680 55995 4000
rect 56775 3680 56795 4000
rect 57005 3680 57025 4000
rect 57805 3680 57825 4000
rect 58340 3680 58360 4000
rect 59140 3680 59160 4000
rect 54670 2570 54690 3140
rect 55410 2570 55430 3140
rect 56480 3125 56500 3145
rect 56480 3075 56500 3095
rect 56480 3025 56500 3045
rect 56480 2975 56500 2995
rect 56480 2925 56500 2945
rect 56890 3125 56910 3145
rect 56890 3075 56910 3095
rect 56890 3025 56910 3045
rect 56890 2975 56910 2995
rect 56890 2925 56910 2945
rect 57300 3125 57320 3145
rect 57300 3075 57320 3095
rect 57300 3025 57320 3045
rect 57300 2975 57320 2995
rect 57300 2925 57320 2945
rect 58370 2570 58390 3140
rect 59110 2570 59130 3140
rect 54670 1695 54690 1865
rect 55410 1695 55430 1865
rect 58370 1695 58390 1865
rect 59110 1695 59130 1865
<< poly >>
rect 56085 4925 56125 4935
rect 56085 4905 56095 4925
rect 56115 4910 56125 4925
rect 56265 4925 56305 4935
rect 56265 4910 56275 4925
rect 56115 4905 56145 4910
rect 56085 4895 56145 4905
rect 56245 4905 56275 4910
rect 56295 4905 56305 4925
rect 56245 4895 56305 4905
rect 57025 4925 57065 4935
rect 57025 4905 57035 4925
rect 57055 4910 57065 4925
rect 57205 4925 57245 4935
rect 57205 4910 57215 4925
rect 57055 4905 57085 4910
rect 57025 4895 57085 4905
rect 57185 4905 57215 4910
rect 57235 4905 57245 4925
rect 57185 4895 57245 4905
rect 57495 4925 57535 4935
rect 57495 4905 57505 4925
rect 57525 4910 57535 4925
rect 57675 4925 57715 4935
rect 57675 4910 57685 4925
rect 57525 4905 57555 4910
rect 57495 4895 57555 4905
rect 57655 4905 57685 4910
rect 57705 4905 57715 4925
rect 57655 4895 57715 4905
rect 56125 4880 56145 4895
rect 56185 4880 56205 4895
rect 56245 4880 56265 4895
rect 57065 4880 57085 4895
rect 57125 4880 57145 4895
rect 57185 4880 57205 4895
rect 57535 4880 57555 4895
rect 57595 4880 57615 4895
rect 57655 4880 57675 4895
rect 56555 4755 56595 4765
rect 56555 4735 56565 4755
rect 56585 4740 56595 4755
rect 56735 4755 56775 4765
rect 56735 4740 56745 4755
rect 56585 4735 56615 4740
rect 56555 4725 56615 4735
rect 56715 4735 56745 4740
rect 56765 4735 56775 4755
rect 56715 4725 56775 4735
rect 56595 4710 56615 4725
rect 56655 4710 56675 4725
rect 56715 4710 56735 4725
rect 56125 4515 56145 4530
rect 56185 4485 56205 4530
rect 56245 4515 56265 4530
rect 56595 4515 56615 4530
rect 56655 4485 56675 4530
rect 56715 4515 56735 4530
rect 57065 4515 57085 4530
rect 56150 4475 56205 4485
rect 56150 4455 56160 4475
rect 56180 4455 56205 4475
rect 56150 4445 56205 4455
rect 56630 4475 56675 4485
rect 56630 4455 56635 4475
rect 56655 4470 56675 4475
rect 57125 4485 57145 4530
rect 57185 4515 57205 4530
rect 57535 4515 57555 4530
rect 57125 4475 57170 4485
rect 57595 4475 57615 4530
rect 57655 4515 57675 4530
rect 57125 4470 57145 4475
rect 56655 4455 56660 4470
rect 56630 4445 56660 4455
rect 57140 4455 57145 4470
rect 57165 4455 57170 4475
rect 57140 4445 57170 4455
rect 57576 4465 57615 4475
rect 57576 4445 57581 4465
rect 57601 4460 57615 4465
rect 57601 4445 57606 4460
rect 57576 4435 57606 4445
rect 54710 4015 54730 4030
rect 54770 4015 54790 4030
rect 54830 4015 54850 4030
rect 54890 4015 54910 4030
rect 54950 4015 54970 4030
rect 55010 4015 55030 4030
rect 55070 4015 55090 4030
rect 55130 4015 55150 4030
rect 55190 4015 55210 4030
rect 55250 4015 55270 4030
rect 55310 4015 55330 4030
rect 55370 4015 55390 4030
rect 56045 4015 56065 4030
rect 56105 4015 56125 4030
rect 56165 4015 56185 4030
rect 56225 4015 56245 4030
rect 56285 4015 56305 4030
rect 56345 4015 56365 4030
rect 56405 4015 56425 4030
rect 56465 4015 56485 4030
rect 56525 4015 56545 4030
rect 56585 4015 56605 4030
rect 56645 4015 56665 4030
rect 56705 4015 56725 4030
rect 57075 4015 57095 4030
rect 57135 4015 57155 4030
rect 57195 4015 57215 4030
rect 57255 4015 57275 4030
rect 57315 4015 57335 4030
rect 57375 4015 57395 4030
rect 57435 4015 57455 4030
rect 57495 4015 57515 4030
rect 57555 4015 57575 4030
rect 57615 4015 57635 4030
rect 57675 4015 57695 4030
rect 57735 4015 57755 4030
rect 58410 4015 58430 4030
rect 58470 4015 58490 4030
rect 58530 4015 58550 4030
rect 58590 4015 58610 4030
rect 58650 4015 58670 4030
rect 58710 4015 58730 4030
rect 58770 4015 58790 4030
rect 58830 4015 58850 4030
rect 58890 4015 58910 4030
rect 58950 4015 58970 4030
rect 59010 4015 59030 4030
rect 59070 4015 59090 4030
rect 54710 3650 54730 3665
rect 54675 3640 54730 3650
rect 54770 3655 54790 3665
rect 54830 3655 54850 3665
rect 54890 3655 54910 3665
rect 54950 3655 54970 3665
rect 55010 3655 55030 3665
rect 55070 3655 55090 3665
rect 55130 3655 55150 3665
rect 55190 3655 55210 3665
rect 55250 3655 55270 3665
rect 55310 3655 55330 3665
rect 54770 3640 55330 3655
rect 55370 3650 55390 3665
rect 56045 3650 56065 3665
rect 55370 3640 55425 3650
rect 54675 3620 54680 3640
rect 54700 3635 54730 3640
rect 54700 3620 54705 3635
rect 54675 3610 54705 3620
rect 55035 3620 55040 3640
rect 55060 3620 55065 3640
rect 55370 3635 55400 3640
rect 55035 3610 55065 3620
rect 55395 3620 55400 3635
rect 55420 3620 55425 3640
rect 55395 3610 55425 3620
rect 56010 3640 56065 3650
rect 56105 3655 56125 3665
rect 56165 3655 56185 3665
rect 56225 3655 56245 3665
rect 56285 3655 56305 3665
rect 56345 3655 56365 3665
rect 56405 3655 56425 3665
rect 56465 3655 56485 3665
rect 56525 3655 56545 3665
rect 56585 3655 56605 3665
rect 56645 3655 56665 3665
rect 56105 3640 56665 3655
rect 56705 3650 56725 3665
rect 57075 3650 57095 3665
rect 56705 3640 56760 3650
rect 56010 3620 56015 3640
rect 56035 3635 56065 3640
rect 56035 3620 56040 3635
rect 56010 3610 56040 3620
rect 56370 3620 56375 3640
rect 56395 3620 56400 3640
rect 56705 3635 56735 3640
rect 56370 3610 56400 3620
rect 56730 3620 56735 3635
rect 56755 3620 56760 3640
rect 56730 3610 56760 3620
rect 57040 3640 57095 3650
rect 57135 3655 57155 3665
rect 57195 3655 57215 3665
rect 57255 3655 57275 3665
rect 57315 3655 57335 3665
rect 57375 3655 57395 3665
rect 57435 3655 57455 3665
rect 57495 3655 57515 3665
rect 57555 3655 57575 3665
rect 57615 3655 57635 3665
rect 57675 3655 57695 3665
rect 57135 3640 57695 3655
rect 57735 3650 57755 3665
rect 58410 3650 58430 3665
rect 57735 3640 57790 3650
rect 57040 3620 57045 3640
rect 57065 3635 57095 3640
rect 57065 3620 57070 3635
rect 57040 3610 57070 3620
rect 57400 3620 57405 3640
rect 57425 3620 57430 3640
rect 57735 3635 57765 3640
rect 57400 3610 57430 3620
rect 57760 3620 57765 3635
rect 57785 3620 57790 3640
rect 57760 3610 57790 3620
rect 58375 3640 58430 3650
rect 58470 3655 58490 3665
rect 58530 3655 58550 3665
rect 58590 3655 58610 3665
rect 58650 3655 58670 3665
rect 58710 3655 58730 3665
rect 58770 3655 58790 3665
rect 58830 3655 58850 3665
rect 58890 3655 58910 3665
rect 58950 3655 58970 3665
rect 59010 3655 59030 3665
rect 58470 3640 59030 3655
rect 59070 3650 59090 3665
rect 59070 3640 59125 3650
rect 58375 3620 58380 3640
rect 58400 3635 58430 3640
rect 58400 3620 58405 3635
rect 58375 3610 58405 3620
rect 58735 3620 58740 3640
rect 58760 3620 58765 3640
rect 59070 3635 59100 3640
rect 58735 3610 58765 3620
rect 59095 3620 59100 3635
rect 59120 3620 59125 3640
rect 59095 3610 59125 3620
rect 55040 3540 55060 3610
rect 56375 3585 56395 3610
rect 57405 3585 57425 3610
rect 56365 3575 56405 3585
rect 56365 3555 56375 3575
rect 56395 3555 56405 3575
rect 56365 3545 56405 3555
rect 57395 3575 57435 3585
rect 57395 3555 57405 3575
rect 57425 3555 57435 3575
rect 57395 3545 57435 3555
rect 58740 3540 58760 3610
rect 55030 3530 55070 3540
rect 55030 3510 55040 3530
rect 55060 3510 55070 3530
rect 55030 3500 55070 3510
rect 58730 3530 58770 3540
rect 58730 3510 58740 3530
rect 58760 3510 58770 3530
rect 58730 3500 58770 3510
rect 56510 3260 56550 3270
rect 56510 3240 56520 3260
rect 56540 3245 56550 3260
rect 56840 3260 56880 3270
rect 56840 3245 56850 3260
rect 56540 3240 56565 3245
rect 56510 3230 56565 3240
rect 54705 3200 54735 3210
rect 54705 3180 54710 3200
rect 54730 3185 54735 3200
rect 55365 3200 55395 3210
rect 55365 3185 55370 3200
rect 54730 3180 54755 3185
rect 54705 3170 54755 3180
rect 55345 3180 55370 3185
rect 55390 3180 55395 3200
rect 55345 3170 55395 3180
rect 54740 3155 54755 3170
rect 54795 3155 54810 3170
rect 54850 3155 54865 3170
rect 54905 3155 54920 3170
rect 54960 3155 54975 3170
rect 55015 3155 55030 3170
rect 55070 3155 55085 3170
rect 55125 3155 55140 3170
rect 55180 3155 55195 3170
rect 55235 3155 55250 3170
rect 55290 3155 55305 3170
rect 55345 3155 55360 3170
rect 56550 3160 56565 3230
rect 56825 3240 56850 3245
rect 56870 3240 56880 3260
rect 56825 3230 56880 3240
rect 56920 3260 56960 3270
rect 56920 3240 56930 3260
rect 56950 3245 56960 3260
rect 57250 3260 57290 3270
rect 57250 3245 57260 3260
rect 56950 3240 56975 3245
rect 56920 3230 56975 3240
rect 56605 3160 56620 3175
rect 56660 3160 56675 3175
rect 56715 3160 56730 3175
rect 56770 3160 56785 3175
rect 56825 3160 56840 3230
rect 56960 3160 56975 3230
rect 57235 3240 57260 3245
rect 57280 3240 57290 3260
rect 57235 3230 57290 3240
rect 57015 3160 57030 3175
rect 57070 3160 57085 3175
rect 57125 3160 57140 3175
rect 57180 3160 57195 3175
rect 57235 3160 57250 3230
rect 58405 3200 58435 3210
rect 58405 3180 58410 3200
rect 58430 3185 58435 3200
rect 59065 3200 59095 3210
rect 59065 3185 59070 3200
rect 58430 3180 58455 3185
rect 58405 3170 58455 3180
rect 59045 3180 59070 3185
rect 59090 3180 59095 3200
rect 59045 3170 59095 3180
rect 58440 3155 58455 3170
rect 58495 3155 58510 3170
rect 58550 3155 58565 3170
rect 58605 3155 58620 3170
rect 58660 3155 58675 3170
rect 58715 3155 58730 3170
rect 58770 3155 58785 3170
rect 58825 3155 58840 3170
rect 58880 3155 58895 3170
rect 58935 3155 58950 3170
rect 58990 3155 59005 3170
rect 59045 3155 59060 3170
rect 56550 2895 56565 2910
rect 56605 2895 56620 2910
rect 56660 2900 56675 2910
rect 56715 2900 56730 2910
rect 56605 2885 56637 2895
rect 56660 2885 56730 2900
rect 56770 2895 56785 2910
rect 56825 2895 56840 2910
rect 56960 2895 56975 2910
rect 57015 2895 57030 2910
rect 57070 2900 57085 2910
rect 57125 2900 57140 2910
rect 56753 2885 56785 2895
rect 57015 2885 57047 2895
rect 57070 2885 57140 2900
rect 57180 2895 57195 2910
rect 57235 2895 57250 2910
rect 57163 2885 57195 2895
rect 56607 2865 56612 2885
rect 56632 2865 56637 2885
rect 56607 2855 56637 2865
rect 56675 2865 56685 2885
rect 56705 2865 56715 2885
rect 56675 2855 56715 2865
rect 56753 2865 56758 2885
rect 56778 2865 56783 2885
rect 56753 2855 56783 2865
rect 57017 2865 57022 2885
rect 57042 2865 57047 2885
rect 57017 2855 57047 2865
rect 57085 2865 57095 2885
rect 57115 2865 57125 2885
rect 57085 2855 57125 2865
rect 57163 2865 57168 2885
rect 57188 2865 57193 2885
rect 57163 2855 57193 2865
rect 56850 2610 56890 2620
rect 56850 2590 56860 2610
rect 56880 2590 56890 2610
rect 56850 2580 56935 2590
rect 56810 2565 56825 2580
rect 56865 2575 56935 2580
rect 56865 2565 56880 2575
rect 56920 2565 56935 2575
rect 56975 2565 56990 2580
rect 54740 2540 54755 2555
rect 54795 2545 54810 2555
rect 54850 2545 54865 2555
rect 54905 2545 54920 2555
rect 54960 2545 54975 2555
rect 55015 2545 55030 2555
rect 55070 2545 55085 2555
rect 55125 2545 55140 2555
rect 55180 2545 55195 2555
rect 55235 2545 55250 2555
rect 55290 2545 55305 2555
rect 54795 2530 55305 2545
rect 55345 2540 55360 2555
rect 55035 2510 55040 2530
rect 55060 2510 55065 2530
rect 55035 2475 55065 2510
rect 55030 2465 55070 2475
rect 55030 2445 55040 2465
rect 55060 2445 55070 2465
rect 55030 2425 55070 2445
rect 55030 2405 55040 2425
rect 55060 2405 55070 2425
rect 55030 2385 55070 2405
rect 55030 2365 55040 2385
rect 55060 2365 55070 2385
rect 55030 2355 55070 2365
rect 58440 2540 58455 2555
rect 58495 2545 58510 2555
rect 58550 2545 58565 2555
rect 58605 2545 58620 2555
rect 58660 2545 58675 2555
rect 58715 2545 58730 2555
rect 58770 2545 58785 2555
rect 58825 2545 58840 2555
rect 58880 2545 58895 2555
rect 58935 2545 58950 2555
rect 58990 2545 59005 2555
rect 58495 2530 59005 2545
rect 59045 2540 59060 2555
rect 58735 2510 58740 2530
rect 58760 2510 58765 2530
rect 58735 2475 58765 2510
rect 58730 2465 58770 2475
rect 58730 2445 58740 2465
rect 58760 2445 58770 2465
rect 58730 2425 58770 2445
rect 58730 2405 58740 2425
rect 58760 2405 58770 2425
rect 58730 2385 58770 2405
rect 58730 2365 58740 2385
rect 58760 2365 58770 2385
rect 58730 2355 58770 2365
rect 56810 2300 56825 2315
rect 56865 2300 56880 2315
rect 56920 2300 56935 2315
rect 56975 2300 56990 2315
rect 56770 2290 56825 2300
rect 56770 2270 56780 2290
rect 56800 2285 56825 2290
rect 56975 2290 57030 2300
rect 56975 2285 57000 2290
rect 56800 2270 56810 2285
rect 56770 2260 56810 2270
rect 56990 2270 57000 2285
rect 57020 2270 57030 2290
rect 56990 2260 57030 2270
rect 55995 1980 56025 1990
rect 55995 1960 56000 1980
rect 56020 1965 56025 1980
rect 56690 1980 56720 1990
rect 56690 1965 56695 1980
rect 56020 1960 56140 1965
rect 55995 1950 56140 1960
rect 54705 1925 54735 1935
rect 54705 1905 54710 1925
rect 54730 1910 54735 1925
rect 55365 1925 55395 1935
rect 55365 1910 55370 1925
rect 54730 1905 54755 1910
rect 54705 1895 54755 1905
rect 55345 1905 55370 1910
rect 55390 1905 55395 1925
rect 56125 1920 56140 1950
rect 56620 1960 56695 1965
rect 56715 1960 56720 1980
rect 56620 1950 56720 1960
rect 57080 1980 57110 1990
rect 57080 1960 57085 1980
rect 57105 1965 57110 1980
rect 57105 1960 57180 1965
rect 57080 1950 57180 1960
rect 56620 1920 56635 1950
rect 55345 1895 55395 1905
rect 56070 1895 56085 1910
rect 56125 1905 56635 1920
rect 57165 1920 57180 1950
rect 58405 1925 58435 1935
rect 56125 1895 56140 1905
rect 56180 1895 56195 1905
rect 56235 1895 56250 1905
rect 56290 1895 56305 1905
rect 56345 1895 56360 1905
rect 56400 1895 56415 1905
rect 56455 1895 56470 1905
rect 56510 1895 56525 1905
rect 56565 1895 56580 1905
rect 56620 1895 56635 1905
rect 56675 1895 56690 1910
rect 57110 1895 57125 1910
rect 57165 1905 57675 1920
rect 57165 1895 57180 1905
rect 57220 1895 57235 1905
rect 57275 1895 57290 1905
rect 57330 1895 57345 1905
rect 57385 1895 57400 1905
rect 57440 1895 57455 1905
rect 57495 1895 57510 1905
rect 57550 1895 57565 1905
rect 57605 1895 57620 1905
rect 57660 1895 57675 1905
rect 57715 1895 57730 1910
rect 58405 1905 58410 1925
rect 58430 1910 58435 1925
rect 59065 1925 59095 1935
rect 59065 1910 59070 1925
rect 58430 1905 58455 1910
rect 58405 1895 58455 1905
rect 59045 1905 59070 1910
rect 59090 1905 59095 1925
rect 59045 1895 59095 1905
rect 54740 1880 54755 1895
rect 54795 1880 54810 1895
rect 54850 1880 54865 1895
rect 54905 1880 54920 1895
rect 54960 1880 54975 1895
rect 55015 1880 55030 1895
rect 55070 1880 55085 1895
rect 55125 1880 55140 1895
rect 55180 1880 55195 1895
rect 55235 1880 55250 1895
rect 55290 1880 55305 1895
rect 55345 1880 55360 1895
rect 58440 1880 58455 1895
rect 58495 1880 58510 1895
rect 58550 1880 58565 1895
rect 58605 1880 58620 1895
rect 58660 1880 58675 1895
rect 58715 1880 58730 1895
rect 58770 1880 58785 1895
rect 58825 1880 58840 1895
rect 58880 1880 58895 1895
rect 58935 1880 58950 1895
rect 58990 1880 59005 1895
rect 59045 1880 59060 1895
rect 56070 1730 56085 1745
rect 56125 1730 56140 1745
rect 56180 1730 56195 1745
rect 56235 1730 56250 1745
rect 56290 1730 56305 1745
rect 56345 1730 56360 1745
rect 56400 1730 56415 1745
rect 56455 1730 56470 1745
rect 56510 1730 56525 1745
rect 56565 1730 56580 1745
rect 56620 1730 56635 1745
rect 56675 1730 56690 1745
rect 57110 1730 57125 1745
rect 57165 1730 57180 1745
rect 57220 1730 57235 1745
rect 57275 1730 57290 1745
rect 57330 1730 57345 1745
rect 57385 1730 57400 1745
rect 57440 1730 57455 1745
rect 57495 1730 57510 1745
rect 57550 1730 57565 1745
rect 57605 1730 57620 1745
rect 57660 1730 57675 1745
rect 57715 1730 57730 1745
rect 56035 1720 56085 1730
rect 56035 1700 56040 1720
rect 56060 1715 56085 1720
rect 56675 1720 56725 1730
rect 56675 1715 56700 1720
rect 56060 1700 56065 1715
rect 56035 1690 56065 1700
rect 56695 1700 56700 1715
rect 56720 1700 56725 1720
rect 56695 1690 56725 1700
rect 57075 1720 57125 1730
rect 57075 1700 57080 1720
rect 57100 1715 57125 1720
rect 57715 1720 57765 1730
rect 57715 1715 57740 1720
rect 57100 1700 57105 1715
rect 57075 1690 57105 1700
rect 57735 1700 57740 1715
rect 57760 1700 57765 1720
rect 57735 1690 57765 1700
rect 54740 1665 54755 1680
rect 54795 1670 54810 1680
rect 54850 1670 54865 1680
rect 54905 1670 54920 1680
rect 54960 1670 54975 1680
rect 55015 1670 55030 1680
rect 55070 1670 55085 1680
rect 55125 1670 55140 1680
rect 55180 1670 55195 1680
rect 55235 1670 55250 1680
rect 55290 1670 55305 1680
rect 54795 1655 55305 1670
rect 55345 1665 55360 1680
rect 58440 1665 58455 1680
rect 58495 1670 58510 1680
rect 58550 1670 58565 1680
rect 58605 1670 58620 1680
rect 58660 1670 58675 1680
rect 58715 1670 58730 1680
rect 58770 1670 58785 1680
rect 58825 1670 58840 1680
rect 58880 1670 58895 1680
rect 58935 1670 58950 1680
rect 58990 1670 59005 1680
rect 58495 1655 59005 1670
rect 59045 1665 59060 1680
rect 55200 1635 55205 1655
rect 55225 1635 55230 1655
rect 55200 1625 55230 1635
rect 58570 1635 58575 1655
rect 58595 1635 58600 1655
rect 58570 1625 58600 1635
rect 55205 1600 55225 1625
rect 58575 1600 58595 1625
rect 55195 1590 55235 1600
rect 55195 1570 55205 1590
rect 55225 1570 55235 1590
rect 55195 1550 55235 1570
rect 55195 1530 55205 1550
rect 55225 1530 55235 1550
rect 55195 1520 55235 1530
rect 58565 1590 58605 1600
rect 58565 1570 58575 1590
rect 58595 1570 58605 1590
rect 58565 1550 58605 1570
rect 58565 1530 58575 1550
rect 58595 1530 58605 1550
rect 58565 1520 58605 1530
rect 55205 1495 55225 1520
rect 58575 1495 58595 1520
rect 55200 1485 55230 1495
rect 55200 1465 55205 1485
rect 55225 1465 55230 1485
rect 58570 1485 58600 1495
rect 58570 1465 58575 1485
rect 58595 1465 58600 1485
rect 54740 1440 54755 1455
rect 54795 1450 55305 1465
rect 54795 1440 54810 1450
rect 54850 1440 54865 1450
rect 54905 1440 54920 1450
rect 54960 1440 54975 1450
rect 55015 1440 55030 1450
rect 55070 1440 55085 1450
rect 55125 1440 55140 1450
rect 55180 1440 55195 1450
rect 55235 1440 55250 1450
rect 55290 1440 55305 1450
rect 55345 1440 55360 1455
rect 58440 1440 58455 1455
rect 58495 1450 59005 1465
rect 58495 1440 58510 1450
rect 58550 1440 58565 1450
rect 58605 1440 58620 1450
rect 58660 1440 58675 1450
rect 58715 1440 58730 1450
rect 58770 1440 58785 1450
rect 58825 1440 58840 1450
rect 58880 1440 58895 1450
rect 58935 1440 58950 1450
rect 58990 1440 59005 1450
rect 59045 1440 59060 1455
rect 56690 1300 56720 1310
rect 56040 1290 56070 1300
rect 56040 1270 56045 1290
rect 56065 1275 56070 1290
rect 56690 1285 56695 1300
rect 56620 1280 56695 1285
rect 56715 1280 56720 1300
rect 56065 1270 56140 1275
rect 56040 1260 56140 1270
rect 56125 1245 56140 1260
rect 56620 1270 56720 1280
rect 56840 1300 56870 1310
rect 56840 1280 56845 1300
rect 56865 1285 56870 1300
rect 56930 1300 56960 1310
rect 56930 1285 56935 1300
rect 56865 1280 56880 1285
rect 56840 1270 56880 1280
rect 56620 1245 56635 1270
rect 56070 1220 56085 1235
rect 56125 1230 56635 1245
rect 56125 1220 56140 1230
rect 56180 1220 56195 1230
rect 56235 1220 56250 1230
rect 56290 1220 56305 1230
rect 56345 1220 56360 1230
rect 56400 1220 56415 1230
rect 56455 1220 56470 1230
rect 56510 1220 56525 1230
rect 56565 1220 56580 1230
rect 56620 1220 56635 1230
rect 56675 1220 56690 1235
rect 56810 1220 56825 1235
rect 56865 1220 56880 1270
rect 56920 1280 56935 1285
rect 56955 1280 56960 1300
rect 56920 1270 56960 1280
rect 57080 1300 57110 1310
rect 57080 1280 57085 1300
rect 57105 1285 57110 1300
rect 57730 1290 57760 1300
rect 57105 1280 57180 1285
rect 57080 1270 57180 1280
rect 57730 1275 57735 1290
rect 56920 1220 56935 1270
rect 57165 1245 57180 1270
rect 57660 1270 57735 1275
rect 57755 1270 57760 1290
rect 57660 1260 57760 1270
rect 57660 1245 57675 1260
rect 56975 1220 56990 1235
rect 57110 1220 57125 1235
rect 57165 1230 57675 1245
rect 57165 1220 57180 1230
rect 57220 1220 57235 1230
rect 57275 1220 57290 1230
rect 57330 1220 57345 1230
rect 57385 1220 57400 1230
rect 57440 1220 57455 1230
rect 57495 1220 57510 1230
rect 57550 1220 57565 1230
rect 57605 1220 57620 1230
rect 57660 1220 57675 1230
rect 57715 1220 57730 1235
rect 54740 1125 54755 1140
rect 54795 1125 54810 1140
rect 54850 1125 54865 1140
rect 54905 1125 54920 1140
rect 54960 1125 54975 1140
rect 55015 1125 55030 1140
rect 55070 1125 55085 1140
rect 55125 1125 55140 1140
rect 55180 1125 55195 1140
rect 55235 1125 55250 1140
rect 55290 1125 55305 1140
rect 55345 1125 55360 1140
rect 54705 1115 54755 1125
rect 54705 1095 54710 1115
rect 54730 1110 54755 1115
rect 55345 1115 55395 1125
rect 55345 1110 55370 1115
rect 54730 1095 54735 1110
rect 54705 1080 54735 1095
rect 55365 1095 55370 1110
rect 55390 1095 55395 1115
rect 55365 1080 55395 1095
rect 58440 1125 58455 1140
rect 58495 1125 58510 1140
rect 58550 1125 58565 1140
rect 58605 1125 58620 1140
rect 58660 1125 58675 1140
rect 58715 1125 58730 1140
rect 58770 1125 58785 1140
rect 58825 1125 58840 1140
rect 58880 1125 58895 1140
rect 58935 1125 58950 1140
rect 58990 1125 59005 1140
rect 59045 1125 59060 1140
rect 58405 1115 58455 1125
rect 58405 1095 58410 1115
rect 58430 1110 58455 1115
rect 59045 1115 59095 1125
rect 59045 1110 59070 1115
rect 58430 1095 58435 1110
rect 58405 1080 58435 1095
rect 59065 1095 59070 1110
rect 59090 1095 59095 1115
rect 59065 1085 59095 1095
rect 56070 1055 56085 1070
rect 56125 1055 56140 1070
rect 56180 1055 56195 1070
rect 56235 1055 56250 1070
rect 56290 1055 56305 1070
rect 56345 1055 56360 1070
rect 56400 1055 56415 1070
rect 56455 1055 56470 1070
rect 56510 1055 56525 1070
rect 56565 1055 56580 1070
rect 56620 1055 56635 1070
rect 56675 1055 56690 1070
rect 56810 1055 56825 1070
rect 56865 1055 56880 1070
rect 56920 1055 56935 1070
rect 56975 1055 56990 1070
rect 57110 1055 57125 1070
rect 57165 1055 57180 1070
rect 57220 1055 57235 1070
rect 57275 1055 57290 1070
rect 57330 1055 57345 1070
rect 57385 1055 57400 1070
rect 57440 1055 57455 1070
rect 57495 1055 57510 1070
rect 57550 1055 57565 1070
rect 57605 1055 57620 1070
rect 57660 1055 57675 1070
rect 57715 1055 57730 1070
rect 56035 1045 56085 1055
rect 56035 1025 56040 1045
rect 56060 1040 56085 1045
rect 56675 1045 56825 1055
rect 56675 1040 56740 1045
rect 56060 1025 56065 1040
rect 56035 1015 56065 1025
rect 56735 1025 56740 1040
rect 56760 1040 56825 1045
rect 56975 1045 57125 1055
rect 56975 1040 57040 1045
rect 56760 1025 56765 1040
rect 56735 1015 56765 1025
rect 57035 1025 57040 1040
rect 57060 1040 57125 1045
rect 57715 1045 57765 1055
rect 57715 1040 57740 1045
rect 57060 1025 57065 1040
rect 57035 1015 57065 1025
rect 57735 1025 57740 1040
rect 57760 1025 57765 1045
rect 57735 1015 57765 1025
rect 55080 430 55120 440
rect 55080 410 55090 430
rect 55110 410 55120 430
rect 55080 400 55120 410
rect 58680 430 58720 440
rect 58680 410 58690 430
rect 58710 410 58720 430
rect 58680 400 58720 410
rect 55090 205 55110 400
rect 56825 375 56865 385
rect 56825 355 56835 375
rect 56855 355 56865 375
rect 56935 375 56975 385
rect 56935 355 56945 375
rect 56965 355 56975 375
rect 56260 330 56275 345
rect 56315 340 57375 355
rect 56315 330 56330 340
rect 56370 330 56385 340
rect 56425 330 56440 340
rect 56480 330 56495 340
rect 56535 330 56550 340
rect 56590 330 56605 340
rect 56645 330 56660 340
rect 56700 330 56715 340
rect 56755 330 56770 340
rect 56810 330 56825 340
rect 56865 330 56880 340
rect 56920 330 56935 340
rect 56975 330 56990 340
rect 57030 330 57045 340
rect 57085 330 57100 340
rect 57140 330 57155 340
rect 57195 330 57210 340
rect 57250 330 57265 340
rect 57305 330 57320 340
rect 57360 330 57375 340
rect 57415 330 57430 345
rect 57470 330 57485 345
rect 54770 180 54830 195
rect 54870 190 55230 205
rect 54870 180 54930 190
rect 54970 180 55030 190
rect 55070 180 55130 190
rect 55170 180 55230 190
rect 55270 180 55330 195
rect 58690 205 58710 400
rect 58470 180 58530 195
rect 58570 190 58930 205
rect 58570 180 58630 190
rect 58670 180 58730 190
rect 58770 180 58830 190
rect 58870 180 58930 190
rect 58970 180 59030 195
rect 56260 65 56275 80
rect 56315 65 56330 80
rect 56370 65 56385 80
rect 56425 65 56440 80
rect 56480 65 56495 80
rect 56535 65 56550 80
rect 56590 65 56605 80
rect 56645 65 56660 80
rect 56700 65 56715 80
rect 56755 65 56770 80
rect 56810 65 56825 80
rect 56865 65 56880 80
rect 56920 65 56935 80
rect 56975 65 56990 80
rect 57030 65 57045 80
rect 57085 65 57100 80
rect 57140 65 57155 80
rect 57195 65 57210 80
rect 57250 65 57265 80
rect 57305 65 57320 80
rect 57360 65 57375 80
rect 56220 55 56275 65
rect 56220 35 56230 55
rect 56250 50 56275 55
rect 56250 35 56260 50
rect 56220 25 56260 35
rect 57415 -35 57430 80
rect 57470 65 57485 80
rect 57470 55 57525 65
rect 57470 50 57495 55
rect 57485 35 57495 50
rect 57515 35 57525 55
rect 57485 25 57525 35
rect 57415 -45 57455 -35
rect 57415 -65 57425 -45
rect 57445 -65 57455 -45
rect 57415 -75 57455 -65
rect 56595 -280 56635 -270
rect 56595 -300 56605 -280
rect 56625 -300 56635 -280
rect 57040 -280 57080 -270
rect 57040 -300 57050 -280
rect 57070 -300 57080 -280
rect 56470 -325 56485 -310
rect 56525 -315 56705 -300
rect 57040 -310 57080 -300
rect 56525 -325 56540 -315
rect 56580 -325 56595 -315
rect 56635 -325 56650 -315
rect 56690 -325 56705 -315
rect 56745 -325 56760 -310
rect 56910 -325 57210 -310
rect 56470 -490 56485 -475
rect 56525 -490 56540 -475
rect 56580 -490 56595 -475
rect 56635 -490 56650 -475
rect 56690 -490 56705 -475
rect 56745 -490 56760 -475
rect 56910 -490 57210 -475
rect 56435 -500 56485 -490
rect 56435 -520 56440 -500
rect 56460 -505 56485 -500
rect 56745 -500 56795 -490
rect 56745 -505 56770 -500
rect 56460 -520 56465 -505
rect 54770 -535 54830 -520
rect 54870 -535 54930 -520
rect 54970 -535 55030 -520
rect 55070 -535 55130 -520
rect 55170 -535 55230 -520
rect 55270 -535 55330 -520
rect 56435 -530 56465 -520
rect 56765 -520 56770 -505
rect 56790 -520 56795 -500
rect 56765 -530 56795 -520
rect 58470 -535 58530 -520
rect 58570 -535 58630 -520
rect 58670 -535 58730 -520
rect 58770 -535 58830 -520
rect 58870 -535 58930 -520
rect 58970 -535 59030 -520
rect 54735 -545 54830 -535
rect 54735 -565 54740 -545
rect 54760 -550 54830 -545
rect 55270 -545 55365 -535
rect 55270 -550 55340 -545
rect 54760 -565 54765 -550
rect 54735 -575 54765 -565
rect 55335 -565 55340 -550
rect 55360 -565 55365 -545
rect 55335 -575 55365 -565
rect 58435 -545 58530 -535
rect 58435 -565 58440 -545
rect 58460 -550 58530 -545
rect 58970 -545 59065 -535
rect 58970 -550 59040 -545
rect 58460 -565 58465 -550
rect 58435 -575 58465 -565
rect 59035 -565 59040 -550
rect 59060 -565 59065 -545
rect 59035 -575 59065 -565
<< polycont >>
rect 56095 4905 56115 4925
rect 56275 4905 56295 4925
rect 57035 4905 57055 4925
rect 57215 4905 57235 4925
rect 57505 4905 57525 4925
rect 57685 4905 57705 4925
rect 56565 4735 56585 4755
rect 56745 4735 56765 4755
rect 56160 4455 56180 4475
rect 56635 4455 56655 4475
rect 57145 4455 57165 4475
rect 57581 4445 57601 4465
rect 54680 3620 54700 3640
rect 55040 3620 55060 3640
rect 55400 3620 55420 3640
rect 56015 3620 56035 3640
rect 56375 3620 56395 3640
rect 56735 3620 56755 3640
rect 57045 3620 57065 3640
rect 57405 3620 57425 3640
rect 57765 3620 57785 3640
rect 58380 3620 58400 3640
rect 58740 3620 58760 3640
rect 59100 3620 59120 3640
rect 56375 3555 56395 3575
rect 57405 3555 57425 3575
rect 55040 3510 55060 3530
rect 58740 3510 58760 3530
rect 56520 3240 56540 3260
rect 54710 3180 54730 3200
rect 55370 3180 55390 3200
rect 56850 3240 56870 3260
rect 56930 3240 56950 3260
rect 57260 3240 57280 3260
rect 58410 3180 58430 3200
rect 59070 3180 59090 3200
rect 56612 2865 56632 2885
rect 56685 2865 56705 2885
rect 56758 2865 56778 2885
rect 57022 2865 57042 2885
rect 57095 2865 57115 2885
rect 57168 2865 57188 2885
rect 56860 2590 56880 2610
rect 55040 2510 55060 2530
rect 55040 2445 55060 2465
rect 55040 2405 55060 2425
rect 55040 2365 55060 2385
rect 58740 2510 58760 2530
rect 58740 2445 58760 2465
rect 58740 2405 58760 2425
rect 58740 2365 58760 2385
rect 56780 2270 56800 2290
rect 57000 2270 57020 2290
rect 56000 1960 56020 1980
rect 54710 1905 54730 1925
rect 55370 1905 55390 1925
rect 56695 1960 56715 1980
rect 57085 1960 57105 1980
rect 58410 1905 58430 1925
rect 59070 1905 59090 1925
rect 56040 1700 56060 1720
rect 56700 1700 56720 1720
rect 57080 1700 57100 1720
rect 57740 1700 57760 1720
rect 55205 1635 55225 1655
rect 58575 1635 58595 1655
rect 55205 1570 55225 1590
rect 55205 1530 55225 1550
rect 58575 1570 58595 1590
rect 58575 1530 58595 1550
rect 55205 1465 55225 1485
rect 58575 1465 58595 1485
rect 56045 1270 56065 1290
rect 56695 1280 56715 1300
rect 56845 1280 56865 1300
rect 56935 1280 56955 1300
rect 57085 1280 57105 1300
rect 57735 1270 57755 1290
rect 54710 1095 54730 1115
rect 55370 1095 55390 1115
rect 58410 1095 58430 1115
rect 59070 1095 59090 1115
rect 56040 1025 56060 1045
rect 56740 1025 56760 1045
rect 57040 1025 57060 1045
rect 57740 1025 57760 1045
rect 55090 410 55110 430
rect 58690 410 58710 430
rect 56835 355 56855 375
rect 56945 355 56965 375
rect 56230 35 56250 55
rect 57495 35 57515 55
rect 57425 -65 57445 -45
rect 56605 -300 56625 -280
rect 57050 -300 57070 -280
rect 56440 -520 56460 -500
rect 56770 -520 56790 -500
rect 54740 -565 54760 -545
rect 55340 -565 55360 -545
rect 58440 -565 58460 -545
rect 59040 -565 59060 -545
<< xpolycontact >>
rect 54204 3040 54345 3260
rect 54204 2695 54345 2915
rect 59455 2955 59596 3175
rect 59455 2610 59596 2830
rect 54335 1544 54370 1764
rect 54335 1165 54370 1385
rect 54395 1544 54430 1764
rect 54395 1165 54430 1385
rect 54455 1544 54490 1764
rect 54455 1165 54490 1385
rect 54515 1544 54550 1764
rect 59250 1544 59285 1764
rect 54515 1165 54550 1385
rect 59250 1165 59285 1385
rect 59310 1544 59345 1764
rect 59310 1165 59345 1385
rect 59370 1544 59405 1764
rect 59370 1165 59405 1385
rect 59430 1544 59465 1764
rect 59430 1165 59465 1385
rect 54405 -85 54440 135
rect 54405 -552 54440 -332
rect 54465 -85 54500 135
rect 54465 -552 54500 -332
rect 59300 -85 59335 135
rect 59300 -552 59335 -332
rect 59360 -85 59395 135
rect 59360 -552 59395 -332
<< ppolyres >>
rect 54204 2915 54345 3040
rect 59455 2830 59596 2955
<< xpolyres >>
rect 54335 1385 54370 1544
rect 54395 1385 54430 1544
rect 54455 1385 54490 1544
rect 54515 1385 54550 1544
rect 59250 1385 59285 1544
rect 59310 1385 59345 1544
rect 59370 1385 59405 1544
rect 59430 1385 59465 1544
rect 54405 -332 54440 -85
rect 54465 -332 54500 -85
rect 59300 -332 59335 -85
rect 59360 -332 59395 -85
<< locali >>
rect 56085 4925 56125 4935
rect 56085 4905 56095 4925
rect 56115 4905 56125 4925
rect 56085 4895 56125 4905
rect 56265 4925 56305 4935
rect 56265 4905 56275 4925
rect 56295 4905 56305 4925
rect 56265 4895 56305 4905
rect 57025 4925 57065 4935
rect 57025 4905 57035 4925
rect 57055 4905 57065 4925
rect 57025 4895 57065 4905
rect 57205 4925 57245 4935
rect 57205 4905 57215 4925
rect 57235 4905 57245 4925
rect 57205 4895 57245 4905
rect 57495 4925 57535 4935
rect 57495 4905 57505 4925
rect 57525 4905 57535 4925
rect 57495 4895 57535 4905
rect 57675 4925 57715 4935
rect 57675 4905 57685 4925
rect 57705 4905 57715 4925
rect 57675 4895 57715 4905
rect 56050 4865 56120 4875
rect 56050 4545 56055 4865
rect 56075 4545 56095 4865
rect 56115 4545 56120 4865
rect 56050 4535 56120 4545
rect 56150 4865 56180 4875
rect 56150 4545 56155 4865
rect 56175 4545 56180 4865
rect 56150 4535 56180 4545
rect 56210 4865 56240 4875
rect 56210 4545 56215 4865
rect 56235 4545 56240 4865
rect 56210 4535 56240 4545
rect 56270 4865 56340 4875
rect 56270 4545 56275 4865
rect 56295 4545 56315 4865
rect 56335 4545 56340 4865
rect 56990 4865 57060 4875
rect 56555 4755 56595 4765
rect 56555 4735 56565 4755
rect 56585 4735 56595 4755
rect 56555 4725 56595 4735
rect 56735 4755 56775 4765
rect 56735 4735 56745 4755
rect 56765 4735 56775 4755
rect 56735 4725 56775 4735
rect 56270 4535 56340 4545
rect 56520 4695 56590 4705
rect 56520 4545 56525 4695
rect 56545 4545 56565 4695
rect 56585 4545 56590 4695
rect 56520 4535 56590 4545
rect 56620 4695 56650 4705
rect 56620 4545 56625 4695
rect 56645 4545 56650 4695
rect 56620 4535 56650 4545
rect 56680 4695 56710 4705
rect 56680 4545 56685 4695
rect 56705 4545 56710 4695
rect 56680 4535 56710 4545
rect 56740 4695 56810 4705
rect 56740 4545 56745 4695
rect 56765 4545 56785 4695
rect 56805 4545 56810 4695
rect 56740 4535 56810 4545
rect 56990 4545 56995 4865
rect 57015 4545 57035 4865
rect 57055 4545 57060 4865
rect 56990 4535 57060 4545
rect 57090 4865 57120 4875
rect 57090 4545 57095 4865
rect 57115 4545 57120 4865
rect 57090 4535 57120 4545
rect 57150 4865 57180 4875
rect 57150 4545 57155 4865
rect 57175 4545 57180 4865
rect 57150 4535 57180 4545
rect 57210 4865 57280 4875
rect 57210 4545 57215 4865
rect 57235 4545 57255 4865
rect 57275 4545 57280 4865
rect 57210 4535 57280 4545
rect 57460 4865 57530 4875
rect 57460 4545 57465 4865
rect 57485 4545 57505 4865
rect 57525 4545 57530 4865
rect 57460 4535 57530 4545
rect 57560 4865 57590 4875
rect 57560 4545 57565 4865
rect 57585 4545 57590 4865
rect 57560 4535 57590 4545
rect 57620 4865 57650 4875
rect 57620 4545 57625 4865
rect 57645 4545 57650 4865
rect 57620 4535 57650 4545
rect 57680 4865 57750 4875
rect 57680 4545 57685 4865
rect 57705 4545 57725 4865
rect 57745 4545 57750 4865
rect 57680 4535 57750 4545
rect 56150 4475 56190 4485
rect 56150 4455 56160 4475
rect 56180 4455 56190 4475
rect 56150 4445 56190 4455
rect 56630 4475 56660 4485
rect 56630 4455 56635 4475
rect 56655 4455 56660 4475
rect 56630 4445 56660 4455
rect 57140 4475 57170 4485
rect 57140 4455 57145 4475
rect 57165 4455 57170 4475
rect 57140 4445 57170 4455
rect 57576 4465 57606 4475
rect 57576 4445 57581 4465
rect 57601 4445 57606 4465
rect 57576 4435 57606 4445
rect 54635 4000 54705 4010
rect 54635 3680 54640 4000
rect 54660 3680 54680 4000
rect 54700 3680 54705 4000
rect 54635 3670 54705 3680
rect 54735 4000 54765 4010
rect 54735 3680 54740 4000
rect 54760 3680 54765 4000
rect 54735 3670 54765 3680
rect 54795 4000 54825 4010
rect 54795 3680 54800 4000
rect 54820 3680 54825 4000
rect 54795 3670 54825 3680
rect 54855 4000 54885 4010
rect 54855 3680 54860 4000
rect 54880 3680 54885 4000
rect 54855 3670 54885 3680
rect 54915 4000 54945 4010
rect 54915 3680 54920 4000
rect 54940 3680 54945 4000
rect 54915 3670 54945 3680
rect 54975 4000 55005 4010
rect 54975 3680 54980 4000
rect 55000 3680 55005 4000
rect 54975 3670 55005 3680
rect 55035 4000 55065 4010
rect 55035 3680 55040 4000
rect 55060 3680 55065 4000
rect 55035 3670 55065 3680
rect 55095 4000 55125 4010
rect 55095 3680 55100 4000
rect 55120 3680 55125 4000
rect 55095 3670 55125 3680
rect 55155 4000 55185 4010
rect 55155 3680 55160 4000
rect 55180 3680 55185 4000
rect 55155 3670 55185 3680
rect 55215 4000 55245 4010
rect 55215 3680 55220 4000
rect 55240 3680 55245 4000
rect 55215 3670 55245 3680
rect 55275 4000 55305 4010
rect 55275 3680 55280 4000
rect 55300 3680 55305 4000
rect 55275 3670 55305 3680
rect 55335 4000 55365 4010
rect 55335 3680 55340 4000
rect 55360 3680 55365 4000
rect 55335 3670 55365 3680
rect 55395 4000 55465 4010
rect 55395 3680 55400 4000
rect 55420 3680 55440 4000
rect 55460 3680 55465 4000
rect 55395 3670 55465 3680
rect 55970 4000 56040 4010
rect 55970 3680 55975 4000
rect 55995 3680 56015 4000
rect 56035 3680 56040 4000
rect 55970 3670 56040 3680
rect 56070 4000 56100 4010
rect 56070 3680 56075 4000
rect 56095 3680 56100 4000
rect 56070 3670 56100 3680
rect 56130 4000 56160 4010
rect 56130 3680 56135 4000
rect 56155 3680 56160 4000
rect 56130 3670 56160 3680
rect 56190 4000 56220 4010
rect 56190 3680 56195 4000
rect 56215 3680 56220 4000
rect 56190 3670 56220 3680
rect 56250 4000 56280 4010
rect 56250 3680 56255 4000
rect 56275 3680 56280 4000
rect 56250 3670 56280 3680
rect 56310 4000 56340 4010
rect 56310 3680 56315 4000
rect 56335 3680 56340 4000
rect 56310 3670 56340 3680
rect 56370 4000 56400 4010
rect 56370 3680 56375 4000
rect 56395 3680 56400 4000
rect 56370 3670 56400 3680
rect 56430 4000 56460 4010
rect 56430 3680 56435 4000
rect 56455 3680 56460 4000
rect 56430 3670 56460 3680
rect 56490 4000 56520 4010
rect 56490 3680 56495 4000
rect 56515 3680 56520 4000
rect 56490 3670 56520 3680
rect 56550 4000 56580 4010
rect 56550 3680 56555 4000
rect 56575 3680 56580 4000
rect 56550 3670 56580 3680
rect 56610 4000 56640 4010
rect 56610 3680 56615 4000
rect 56635 3680 56640 4000
rect 56610 3670 56640 3680
rect 56670 4000 56700 4010
rect 56670 3680 56675 4000
rect 56695 3680 56700 4000
rect 56670 3670 56700 3680
rect 56730 4000 56800 4010
rect 56730 3680 56735 4000
rect 56755 3680 56775 4000
rect 56795 3680 56800 4000
rect 56730 3670 56800 3680
rect 57000 4000 57070 4010
rect 57000 3680 57005 4000
rect 57025 3680 57045 4000
rect 57065 3680 57070 4000
rect 57000 3670 57070 3680
rect 57100 4000 57130 4010
rect 57100 3680 57105 4000
rect 57125 3680 57130 4000
rect 57100 3670 57130 3680
rect 57160 4000 57190 4010
rect 57160 3680 57165 4000
rect 57185 3680 57190 4000
rect 57160 3670 57190 3680
rect 57220 4000 57250 4010
rect 57220 3680 57225 4000
rect 57245 3680 57250 4000
rect 57220 3670 57250 3680
rect 57280 4000 57310 4010
rect 57280 3680 57285 4000
rect 57305 3680 57310 4000
rect 57280 3670 57310 3680
rect 57340 4000 57370 4010
rect 57340 3680 57345 4000
rect 57365 3680 57370 4000
rect 57340 3670 57370 3680
rect 57400 4000 57430 4010
rect 57400 3680 57405 4000
rect 57425 3680 57430 4000
rect 57400 3670 57430 3680
rect 57460 4000 57490 4010
rect 57460 3680 57465 4000
rect 57485 3680 57490 4000
rect 57460 3670 57490 3680
rect 57520 4000 57550 4010
rect 57520 3680 57525 4000
rect 57545 3680 57550 4000
rect 57520 3670 57550 3680
rect 57580 4000 57610 4010
rect 57580 3680 57585 4000
rect 57605 3680 57610 4000
rect 57580 3670 57610 3680
rect 57640 4000 57670 4010
rect 57640 3680 57645 4000
rect 57665 3680 57670 4000
rect 57640 3670 57670 3680
rect 57700 4000 57730 4010
rect 57700 3680 57705 4000
rect 57725 3680 57730 4000
rect 57700 3670 57730 3680
rect 57760 4000 57830 4010
rect 57760 3680 57765 4000
rect 57785 3680 57805 4000
rect 57825 3680 57830 4000
rect 57760 3670 57830 3680
rect 58335 4000 58405 4010
rect 58335 3680 58340 4000
rect 58360 3680 58380 4000
rect 58400 3680 58405 4000
rect 58335 3670 58405 3680
rect 58435 4000 58465 4010
rect 58435 3680 58440 4000
rect 58460 3680 58465 4000
rect 58435 3670 58465 3680
rect 58495 4000 58525 4010
rect 58495 3680 58500 4000
rect 58520 3680 58525 4000
rect 58495 3670 58525 3680
rect 58555 4000 58585 4010
rect 58555 3680 58560 4000
rect 58580 3680 58585 4000
rect 58555 3670 58585 3680
rect 58615 4000 58645 4010
rect 58615 3680 58620 4000
rect 58640 3680 58645 4000
rect 58615 3670 58645 3680
rect 58675 4000 58705 4010
rect 58675 3680 58680 4000
rect 58700 3680 58705 4000
rect 58675 3670 58705 3680
rect 58735 4000 58765 4010
rect 58735 3680 58740 4000
rect 58760 3680 58765 4000
rect 58735 3670 58765 3680
rect 58795 4000 58825 4010
rect 58795 3680 58800 4000
rect 58820 3680 58825 4000
rect 58795 3670 58825 3680
rect 58855 4000 58885 4010
rect 58855 3680 58860 4000
rect 58880 3680 58885 4000
rect 58855 3670 58885 3680
rect 58915 4000 58945 4010
rect 58915 3680 58920 4000
rect 58940 3680 58945 4000
rect 58915 3670 58945 3680
rect 58975 4000 59005 4010
rect 58975 3680 58980 4000
rect 59000 3680 59005 4000
rect 58975 3670 59005 3680
rect 59035 4000 59065 4010
rect 59035 3680 59040 4000
rect 59060 3680 59065 4000
rect 59035 3670 59065 3680
rect 59095 4000 59165 4010
rect 59095 3680 59100 4000
rect 59120 3680 59140 4000
rect 59160 3680 59165 4000
rect 59095 3670 59165 3680
rect 54675 3640 54705 3650
rect 54675 3620 54680 3640
rect 54700 3620 54705 3640
rect 54675 3610 54705 3620
rect 55035 3640 55065 3650
rect 55035 3620 55040 3640
rect 55060 3620 55065 3640
rect 55035 3610 55065 3620
rect 55395 3640 55425 3650
rect 55395 3620 55400 3640
rect 55420 3620 55425 3640
rect 55395 3610 55425 3620
rect 56010 3640 56040 3650
rect 56010 3620 56015 3640
rect 56035 3620 56040 3640
rect 56010 3610 56040 3620
rect 56370 3640 56400 3650
rect 56370 3620 56375 3640
rect 56395 3620 56400 3640
rect 56370 3610 56400 3620
rect 56730 3640 56760 3650
rect 56730 3620 56735 3640
rect 56755 3620 56760 3640
rect 56730 3610 56760 3620
rect 57040 3640 57070 3650
rect 57040 3620 57045 3640
rect 57065 3620 57070 3640
rect 57040 3610 57070 3620
rect 57400 3640 57430 3650
rect 57400 3620 57405 3640
rect 57425 3620 57430 3640
rect 57400 3610 57430 3620
rect 57760 3640 57790 3650
rect 57760 3620 57765 3640
rect 57785 3620 57790 3640
rect 57760 3610 57790 3620
rect 58375 3640 58405 3650
rect 58375 3620 58380 3640
rect 58400 3620 58405 3640
rect 58375 3610 58405 3620
rect 58735 3640 58765 3650
rect 58735 3620 58740 3640
rect 58760 3620 58765 3640
rect 58735 3610 58765 3620
rect 59095 3640 59125 3650
rect 59095 3620 59100 3640
rect 59120 3620 59125 3640
rect 59095 3610 59125 3620
rect 56365 3575 56405 3585
rect 56365 3555 56375 3575
rect 56395 3555 56405 3575
rect 56365 3545 56405 3555
rect 57395 3575 57435 3585
rect 57395 3555 57405 3575
rect 57425 3555 57435 3575
rect 57395 3545 57435 3555
rect 55030 3530 55070 3540
rect 55030 3510 55040 3530
rect 55060 3510 55070 3530
rect 55030 3500 55070 3510
rect 58730 3530 58770 3540
rect 58730 3510 58740 3530
rect 58760 3510 58770 3530
rect 58730 3500 58770 3510
rect 54204 3290 54345 3300
rect 54204 3270 54210 3290
rect 54230 3270 54265 3290
rect 54285 3270 54320 3290
rect 54340 3270 54345 3290
rect 54204 3260 54345 3270
rect 56510 3260 56550 3270
rect 56510 3240 56520 3260
rect 56540 3240 56550 3260
rect 56510 3230 56550 3240
rect 56680 3260 56710 3270
rect 56680 3240 56685 3260
rect 56705 3240 56710 3260
rect 56680 3230 56710 3240
rect 56840 3260 56880 3270
rect 56840 3240 56850 3260
rect 56870 3240 56880 3260
rect 56840 3230 56880 3240
rect 56920 3260 56960 3270
rect 56920 3240 56930 3260
rect 56950 3240 56960 3260
rect 56920 3230 56960 3240
rect 57090 3260 57120 3270
rect 57090 3240 57095 3260
rect 57115 3240 57120 3260
rect 57090 3230 57120 3240
rect 57250 3260 57290 3270
rect 57250 3240 57260 3260
rect 57280 3240 57290 3260
rect 57250 3230 57290 3240
rect 54705 3200 54735 3210
rect 54705 3180 54710 3200
rect 54730 3180 54735 3200
rect 54705 3170 54735 3180
rect 55365 3200 55395 3210
rect 55365 3180 55370 3200
rect 55390 3180 55395 3200
rect 55365 3170 55395 3180
rect 56520 3155 56540 3230
rect 56620 3205 56660 3215
rect 56620 3185 56630 3205
rect 56650 3185 56660 3205
rect 56620 3175 56660 3185
rect 56630 3155 56650 3175
rect 56685 3155 56705 3230
rect 56730 3205 56770 3215
rect 56730 3185 56740 3205
rect 56760 3185 56770 3205
rect 56730 3175 56770 3185
rect 56740 3155 56760 3175
rect 56850 3155 56870 3230
rect 56930 3155 56950 3230
rect 57030 3205 57070 3215
rect 57030 3185 57040 3205
rect 57060 3185 57070 3205
rect 57030 3175 57070 3185
rect 57040 3155 57060 3175
rect 57095 3155 57115 3230
rect 57140 3205 57180 3215
rect 57140 3185 57150 3205
rect 57170 3185 57180 3205
rect 57140 3175 57180 3185
rect 57150 3155 57170 3175
rect 57260 3155 57280 3230
rect 58405 3200 58435 3210
rect 58405 3180 58410 3200
rect 58430 3180 58435 3200
rect 58405 3170 58435 3180
rect 59065 3200 59095 3210
rect 59065 3180 59070 3200
rect 59090 3180 59095 3200
rect 59065 3170 59095 3180
rect 59455 3205 59596 3215
rect 59455 3185 59460 3205
rect 59480 3185 59515 3205
rect 59535 3185 59570 3205
rect 59590 3185 59596 3205
rect 59455 3175 59596 3185
rect 54665 3140 54735 3150
rect 54204 2685 54345 2695
rect 54204 2665 54210 2685
rect 54230 2665 54265 2685
rect 54285 2665 54320 2685
rect 54340 2665 54345 2685
rect 54204 2655 54345 2665
rect 54665 2570 54670 3140
rect 54690 2570 54710 3140
rect 54730 2570 54735 3140
rect 54665 2560 54735 2570
rect 54760 3140 54790 3150
rect 54760 2570 54765 3140
rect 54785 2570 54790 3140
rect 54760 2560 54790 2570
rect 54815 3140 54845 3150
rect 54815 2570 54820 3140
rect 54840 2570 54845 3140
rect 54815 2560 54845 2570
rect 54870 3140 54900 3150
rect 54870 2570 54875 3140
rect 54895 2570 54900 3140
rect 54870 2560 54900 2570
rect 54925 3140 54955 3150
rect 54925 2570 54930 3140
rect 54950 2570 54955 3140
rect 54925 2560 54955 2570
rect 54980 3140 55010 3150
rect 54980 2570 54985 3140
rect 55005 2570 55010 3140
rect 54980 2560 55010 2570
rect 55035 3140 55065 3150
rect 55035 2570 55040 3140
rect 55060 2570 55065 3140
rect 55035 2560 55065 2570
rect 55090 3140 55120 3150
rect 55090 2570 55095 3140
rect 55115 2570 55120 3140
rect 55090 2560 55120 2570
rect 55145 3140 55175 3150
rect 55145 2570 55150 3140
rect 55170 2570 55175 3140
rect 55145 2560 55175 2570
rect 55200 3140 55230 3150
rect 55200 2570 55205 3140
rect 55225 2570 55230 3140
rect 55200 2560 55230 2570
rect 55255 3140 55285 3150
rect 55255 2570 55260 3140
rect 55280 2570 55285 3140
rect 55255 2560 55285 2570
rect 55310 3140 55340 3150
rect 55310 2570 55315 3140
rect 55335 2570 55340 3140
rect 55310 2560 55340 2570
rect 55365 3140 55435 3150
rect 55365 2570 55370 3140
rect 55390 2570 55410 3140
rect 55430 2570 55435 3140
rect 56475 3145 56545 3155
rect 56475 3125 56480 3145
rect 56500 3125 56520 3145
rect 56540 3125 56545 3145
rect 56475 3095 56545 3125
rect 56475 3075 56480 3095
rect 56500 3075 56520 3095
rect 56540 3075 56545 3095
rect 56475 3045 56545 3075
rect 56475 3025 56480 3045
rect 56500 3025 56520 3045
rect 56540 3025 56545 3045
rect 56475 2995 56545 3025
rect 56475 2975 56480 2995
rect 56500 2975 56520 2995
rect 56540 2975 56545 2995
rect 56475 2945 56545 2975
rect 56475 2925 56480 2945
rect 56500 2925 56520 2945
rect 56540 2925 56545 2945
rect 56475 2915 56545 2925
rect 56570 3145 56600 3155
rect 56570 3125 56575 3145
rect 56595 3125 56600 3145
rect 56570 3095 56600 3125
rect 56570 3075 56575 3095
rect 56595 3075 56600 3095
rect 56570 3045 56600 3075
rect 56570 3025 56575 3045
rect 56595 3025 56600 3045
rect 56570 2995 56600 3025
rect 56570 2975 56575 2995
rect 56595 2975 56600 2995
rect 56570 2945 56600 2975
rect 56570 2925 56575 2945
rect 56595 2925 56600 2945
rect 56570 2915 56600 2925
rect 56625 3145 56655 3155
rect 56625 3125 56630 3145
rect 56650 3125 56655 3145
rect 56625 3095 56655 3125
rect 56625 3075 56630 3095
rect 56650 3075 56655 3095
rect 56625 3045 56655 3075
rect 56625 3025 56630 3045
rect 56650 3025 56655 3045
rect 56625 2995 56655 3025
rect 56625 2975 56630 2995
rect 56650 2975 56655 2995
rect 56625 2945 56655 2975
rect 56625 2925 56630 2945
rect 56650 2925 56655 2945
rect 56625 2915 56655 2925
rect 56680 3145 56710 3155
rect 56680 3125 56685 3145
rect 56705 3125 56710 3145
rect 56680 3095 56710 3125
rect 56680 3075 56685 3095
rect 56705 3075 56710 3095
rect 56680 3045 56710 3075
rect 56680 3025 56685 3045
rect 56705 3025 56710 3045
rect 56680 2995 56710 3025
rect 56680 2975 56685 2995
rect 56705 2975 56710 2995
rect 56680 2945 56710 2975
rect 56680 2925 56685 2945
rect 56705 2925 56710 2945
rect 56680 2915 56710 2925
rect 56735 3145 56765 3155
rect 56735 3125 56740 3145
rect 56760 3125 56765 3145
rect 56735 3095 56765 3125
rect 56735 3075 56740 3095
rect 56760 3075 56765 3095
rect 56735 3045 56765 3075
rect 56735 3025 56740 3045
rect 56760 3025 56765 3045
rect 56735 2995 56765 3025
rect 56735 2975 56740 2995
rect 56760 2975 56765 2995
rect 56735 2945 56765 2975
rect 56735 2925 56740 2945
rect 56760 2925 56765 2945
rect 56735 2915 56765 2925
rect 56790 3145 56820 3155
rect 56790 3125 56795 3145
rect 56815 3125 56820 3145
rect 56790 3095 56820 3125
rect 56790 3075 56795 3095
rect 56815 3075 56820 3095
rect 56790 3045 56820 3075
rect 56790 3025 56795 3045
rect 56815 3025 56820 3045
rect 56790 2995 56820 3025
rect 56790 2975 56795 2995
rect 56815 2975 56820 2995
rect 56790 2945 56820 2975
rect 56790 2925 56795 2945
rect 56815 2925 56820 2945
rect 56790 2915 56820 2925
rect 56845 3145 56955 3155
rect 56845 3125 56850 3145
rect 56870 3125 56890 3145
rect 56910 3125 56930 3145
rect 56950 3125 56955 3145
rect 56845 3095 56955 3125
rect 56845 3075 56850 3095
rect 56870 3075 56890 3095
rect 56910 3075 56930 3095
rect 56950 3075 56955 3095
rect 56845 3045 56955 3075
rect 56845 3025 56850 3045
rect 56870 3025 56890 3045
rect 56910 3025 56930 3045
rect 56950 3025 56955 3045
rect 56845 2995 56955 3025
rect 56845 2975 56850 2995
rect 56870 2975 56890 2995
rect 56910 2975 56930 2995
rect 56950 2975 56955 2995
rect 56845 2945 56955 2975
rect 56845 2925 56850 2945
rect 56870 2925 56890 2945
rect 56910 2925 56930 2945
rect 56950 2925 56955 2945
rect 56845 2915 56955 2925
rect 56980 3145 57010 3155
rect 56980 3125 56985 3145
rect 57005 3125 57010 3145
rect 56980 3095 57010 3125
rect 56980 3075 56985 3095
rect 57005 3075 57010 3095
rect 56980 3045 57010 3075
rect 56980 3025 56985 3045
rect 57005 3025 57010 3045
rect 56980 2995 57010 3025
rect 56980 2975 56985 2995
rect 57005 2975 57010 2995
rect 56980 2945 57010 2975
rect 56980 2925 56985 2945
rect 57005 2925 57010 2945
rect 56980 2915 57010 2925
rect 57035 3145 57065 3155
rect 57035 3125 57040 3145
rect 57060 3125 57065 3145
rect 57035 3095 57065 3125
rect 57035 3075 57040 3095
rect 57060 3075 57065 3095
rect 57035 3045 57065 3075
rect 57035 3025 57040 3045
rect 57060 3025 57065 3045
rect 57035 2995 57065 3025
rect 57035 2975 57040 2995
rect 57060 2975 57065 2995
rect 57035 2945 57065 2975
rect 57035 2925 57040 2945
rect 57060 2925 57065 2945
rect 57035 2915 57065 2925
rect 57090 3145 57120 3155
rect 57090 3125 57095 3145
rect 57115 3125 57120 3145
rect 57090 3095 57120 3125
rect 57090 3075 57095 3095
rect 57115 3075 57120 3095
rect 57090 3045 57120 3075
rect 57090 3025 57095 3045
rect 57115 3025 57120 3045
rect 57090 2995 57120 3025
rect 57090 2975 57095 2995
rect 57115 2975 57120 2995
rect 57090 2945 57120 2975
rect 57090 2925 57095 2945
rect 57115 2925 57120 2945
rect 57090 2915 57120 2925
rect 57145 3145 57175 3155
rect 57145 3125 57150 3145
rect 57170 3125 57175 3145
rect 57145 3095 57175 3125
rect 57145 3075 57150 3095
rect 57170 3075 57175 3095
rect 57145 3045 57175 3075
rect 57145 3025 57150 3045
rect 57170 3025 57175 3045
rect 57145 2995 57175 3025
rect 57145 2975 57150 2995
rect 57170 2975 57175 2995
rect 57145 2945 57175 2975
rect 57145 2925 57150 2945
rect 57170 2925 57175 2945
rect 57145 2915 57175 2925
rect 57200 3145 57230 3155
rect 57200 3125 57205 3145
rect 57225 3125 57230 3145
rect 57200 3095 57230 3125
rect 57200 3075 57205 3095
rect 57225 3075 57230 3095
rect 57200 3045 57230 3075
rect 57200 3025 57205 3045
rect 57225 3025 57230 3045
rect 57200 2995 57230 3025
rect 57200 2975 57205 2995
rect 57225 2975 57230 2995
rect 57200 2945 57230 2975
rect 57200 2925 57205 2945
rect 57225 2925 57230 2945
rect 57200 2915 57230 2925
rect 57255 3145 57325 3155
rect 57255 3125 57260 3145
rect 57280 3125 57300 3145
rect 57320 3125 57325 3145
rect 57255 3095 57325 3125
rect 57255 3075 57260 3095
rect 57280 3075 57300 3095
rect 57320 3075 57325 3095
rect 57255 3045 57325 3075
rect 57255 3025 57260 3045
rect 57280 3025 57300 3045
rect 57320 3025 57325 3045
rect 57255 2995 57325 3025
rect 57255 2975 57260 2995
rect 57280 2975 57300 2995
rect 57320 2975 57325 2995
rect 57255 2945 57325 2975
rect 57255 2925 57260 2945
rect 57280 2925 57300 2945
rect 57320 2925 57325 2945
rect 57255 2915 57325 2925
rect 58365 3140 58435 3150
rect 56570 2905 56590 2915
rect 56560 2895 56590 2905
rect 56800 2905 56820 2915
rect 56980 2905 57000 2915
rect 56800 2895 56830 2905
rect 56560 2875 56565 2895
rect 56585 2875 56590 2895
rect 56560 2865 56590 2875
rect 56607 2885 56637 2895
rect 56607 2865 56612 2885
rect 56632 2865 56637 2885
rect 56607 2855 56637 2865
rect 56675 2885 56715 2895
rect 56675 2865 56685 2885
rect 56705 2865 56715 2885
rect 56675 2855 56715 2865
rect 56753 2885 56783 2895
rect 56753 2865 56758 2885
rect 56778 2865 56783 2885
rect 56800 2875 56805 2895
rect 56825 2875 56830 2895
rect 56800 2865 56830 2875
rect 56970 2895 57000 2905
rect 57210 2905 57230 2915
rect 57210 2895 57240 2905
rect 56970 2875 56975 2895
rect 56995 2875 57000 2895
rect 56970 2865 57000 2875
rect 57017 2885 57047 2895
rect 57017 2865 57022 2885
rect 57042 2865 57047 2885
rect 56753 2855 56783 2865
rect 57017 2855 57047 2865
rect 57085 2885 57125 2895
rect 57085 2865 57095 2885
rect 57115 2865 57125 2885
rect 57085 2855 57125 2865
rect 57163 2885 57193 2895
rect 57163 2865 57168 2885
rect 57188 2865 57193 2885
rect 57210 2875 57215 2895
rect 57235 2875 57240 2895
rect 57210 2865 57240 2875
rect 57163 2855 57193 2865
rect 56600 2825 56640 2835
rect 56600 2805 56610 2825
rect 56630 2805 56640 2825
rect 56600 2795 56640 2805
rect 57160 2825 57200 2835
rect 57160 2805 57170 2825
rect 57190 2805 57200 2825
rect 57160 2795 57200 2805
rect 56850 2610 56890 2620
rect 56850 2590 56860 2610
rect 56880 2590 56890 2610
rect 56850 2580 56890 2590
rect 56935 2610 56975 2620
rect 56935 2590 56945 2610
rect 56965 2590 56975 2610
rect 56935 2580 56975 2590
rect 55365 2560 55435 2570
rect 58365 2570 58370 3140
rect 58390 2570 58410 3140
rect 58430 2570 58435 3140
rect 58365 2560 58435 2570
rect 58460 3140 58490 3150
rect 58460 2570 58465 3140
rect 58485 2570 58490 3140
rect 58460 2560 58490 2570
rect 58515 3140 58545 3150
rect 58515 2570 58520 3140
rect 58540 2570 58545 3140
rect 58515 2560 58545 2570
rect 58570 3140 58600 3150
rect 58570 2570 58575 3140
rect 58595 2570 58600 3140
rect 58570 2560 58600 2570
rect 58625 3140 58655 3150
rect 58625 2570 58630 3140
rect 58650 2570 58655 3140
rect 58625 2560 58655 2570
rect 58680 3140 58710 3150
rect 58680 2570 58685 3140
rect 58705 2570 58710 3140
rect 58680 2560 58710 2570
rect 58735 3140 58765 3150
rect 58735 2570 58740 3140
rect 58760 2570 58765 3140
rect 58735 2560 58765 2570
rect 58790 3140 58820 3150
rect 58790 2570 58795 3140
rect 58815 2570 58820 3140
rect 58790 2560 58820 2570
rect 58845 3140 58875 3150
rect 58845 2570 58850 3140
rect 58870 2570 58875 3140
rect 58845 2560 58875 2570
rect 58900 3140 58930 3150
rect 58900 2570 58905 3140
rect 58925 2570 58930 3140
rect 58900 2560 58930 2570
rect 58955 3140 58985 3150
rect 58955 2570 58960 3140
rect 58980 2570 58985 3140
rect 58955 2560 58985 2570
rect 59010 3140 59040 3150
rect 59010 2570 59015 3140
rect 59035 2570 59040 3140
rect 59010 2560 59040 2570
rect 59065 3140 59135 3150
rect 59065 2570 59070 3140
rect 59090 2570 59110 3140
rect 59130 2570 59135 3140
rect 59455 2600 59596 2610
rect 59455 2580 59460 2600
rect 59480 2580 59515 2600
rect 59535 2580 59570 2600
rect 59590 2580 59596 2600
rect 59455 2570 59596 2580
rect 59065 2560 59135 2570
rect 56735 2550 56805 2560
rect 55035 2530 55065 2540
rect 55035 2510 55040 2530
rect 55060 2510 55065 2530
rect 55035 2500 55065 2510
rect 55030 2465 55070 2475
rect 55030 2445 55040 2465
rect 55060 2445 55070 2465
rect 55030 2425 55070 2445
rect 55030 2405 55040 2425
rect 55060 2405 55070 2425
rect 55030 2385 55070 2405
rect 55030 2365 55040 2385
rect 55060 2365 55070 2385
rect 55030 2355 55070 2365
rect 56735 2330 56740 2550
rect 56760 2330 56780 2550
rect 56800 2330 56805 2550
rect 56735 2320 56805 2330
rect 56830 2550 56860 2560
rect 56830 2330 56835 2550
rect 56855 2330 56860 2550
rect 56830 2320 56860 2330
rect 56885 2550 56915 2560
rect 56885 2330 56890 2550
rect 56910 2330 56915 2550
rect 56885 2320 56915 2330
rect 56940 2550 56970 2560
rect 56940 2330 56945 2550
rect 56965 2330 56970 2550
rect 56940 2320 56970 2330
rect 56995 2550 57065 2560
rect 56995 2330 57000 2550
rect 57020 2330 57040 2550
rect 57060 2330 57065 2550
rect 58735 2530 58765 2540
rect 58735 2510 58740 2530
rect 58760 2510 58765 2530
rect 58735 2500 58765 2510
rect 58730 2465 58770 2475
rect 58730 2445 58740 2465
rect 58760 2445 58770 2465
rect 58730 2425 58770 2445
rect 58730 2405 58740 2425
rect 58760 2405 58770 2425
rect 58730 2385 58770 2405
rect 58730 2365 58740 2385
rect 58760 2365 58770 2385
rect 58730 2355 58770 2365
rect 56995 2320 57065 2330
rect 56770 2290 56810 2300
rect 56770 2270 56780 2290
rect 56800 2270 56810 2290
rect 56770 2260 56810 2270
rect 56990 2290 57030 2300
rect 56990 2270 57000 2290
rect 57020 2270 57030 2290
rect 56990 2260 57030 2270
rect 55995 1980 56025 1990
rect 55995 1960 56000 1980
rect 56020 1960 56025 1980
rect 55995 1950 56025 1960
rect 56690 1980 56720 1990
rect 56690 1960 56695 1980
rect 56715 1960 56720 1980
rect 56690 1950 56720 1960
rect 57080 1980 57110 1990
rect 57080 1960 57085 1980
rect 57105 1960 57110 1980
rect 57080 1950 57110 1960
rect 54705 1925 54735 1935
rect 54705 1905 54710 1925
rect 54730 1905 54735 1925
rect 54705 1895 54735 1905
rect 55365 1925 55395 1935
rect 55365 1905 55370 1925
rect 55390 1905 55395 1925
rect 55365 1895 55395 1905
rect 58405 1925 58435 1935
rect 58405 1905 58410 1925
rect 58430 1905 58435 1925
rect 58405 1895 58435 1905
rect 59065 1925 59095 1935
rect 59065 1905 59070 1925
rect 59090 1905 59095 1925
rect 59065 1895 59095 1905
rect 55995 1880 56065 1890
rect 54665 1865 54735 1875
rect 54335 1781 54550 1801
rect 54335 1764 54370 1781
rect 54515 1764 54550 1781
rect 54430 1714 54455 1764
rect 54665 1695 54670 1865
rect 54690 1695 54710 1865
rect 54730 1695 54735 1865
rect 54665 1685 54735 1695
rect 54760 1865 54790 1875
rect 54760 1695 54765 1865
rect 54785 1695 54790 1865
rect 54760 1685 54790 1695
rect 54815 1865 54845 1875
rect 54815 1695 54820 1865
rect 54840 1695 54845 1865
rect 54815 1685 54845 1695
rect 54870 1865 54900 1875
rect 54870 1695 54875 1865
rect 54895 1695 54900 1865
rect 54870 1685 54900 1695
rect 54925 1865 54955 1875
rect 54925 1695 54930 1865
rect 54950 1695 54955 1865
rect 54925 1685 54955 1695
rect 54980 1865 55010 1875
rect 54980 1695 54985 1865
rect 55005 1695 55010 1865
rect 54980 1685 55010 1695
rect 55035 1865 55065 1875
rect 55035 1695 55040 1865
rect 55060 1695 55065 1865
rect 55035 1685 55065 1695
rect 55090 1865 55120 1875
rect 55090 1695 55095 1865
rect 55115 1695 55120 1865
rect 55090 1685 55120 1695
rect 55145 1865 55175 1875
rect 55145 1695 55150 1865
rect 55170 1695 55175 1865
rect 55145 1685 55175 1695
rect 55200 1865 55230 1875
rect 55200 1695 55205 1865
rect 55225 1695 55230 1865
rect 55200 1685 55230 1695
rect 55255 1865 55285 1875
rect 55255 1695 55260 1865
rect 55280 1695 55285 1865
rect 55255 1685 55285 1695
rect 55310 1865 55340 1875
rect 55310 1695 55315 1865
rect 55335 1695 55340 1865
rect 55310 1685 55340 1695
rect 55365 1865 55435 1875
rect 55365 1695 55370 1865
rect 55390 1695 55410 1865
rect 55430 1695 55435 1865
rect 55995 1760 56000 1880
rect 56020 1760 56040 1880
rect 56060 1760 56065 1880
rect 55995 1750 56065 1760
rect 56090 1880 56120 1890
rect 56090 1760 56095 1880
rect 56115 1760 56120 1880
rect 56090 1750 56120 1760
rect 56145 1880 56175 1890
rect 56145 1760 56150 1880
rect 56170 1760 56175 1880
rect 56145 1750 56175 1760
rect 56200 1880 56230 1890
rect 56200 1760 56205 1880
rect 56225 1760 56230 1880
rect 56200 1750 56230 1760
rect 56255 1880 56285 1890
rect 56255 1760 56260 1880
rect 56280 1760 56285 1880
rect 56255 1750 56285 1760
rect 56310 1880 56340 1890
rect 56310 1760 56315 1880
rect 56335 1760 56340 1880
rect 56310 1750 56340 1760
rect 56365 1880 56395 1890
rect 56365 1760 56370 1880
rect 56390 1760 56395 1880
rect 56365 1750 56395 1760
rect 56420 1880 56450 1890
rect 56420 1760 56425 1880
rect 56445 1760 56450 1880
rect 56420 1750 56450 1760
rect 56475 1880 56505 1890
rect 56475 1760 56480 1880
rect 56500 1760 56505 1880
rect 56475 1750 56505 1760
rect 56530 1880 56560 1890
rect 56530 1760 56535 1880
rect 56555 1760 56560 1880
rect 56530 1750 56560 1760
rect 56585 1880 56615 1890
rect 56585 1760 56590 1880
rect 56610 1760 56615 1880
rect 56585 1750 56615 1760
rect 56640 1880 56670 1890
rect 56640 1760 56645 1880
rect 56665 1760 56670 1880
rect 56640 1750 56670 1760
rect 56695 1880 56765 1890
rect 56695 1760 56700 1880
rect 56720 1760 56740 1880
rect 56760 1760 56765 1880
rect 56695 1750 56765 1760
rect 57035 1880 57105 1890
rect 57035 1760 57040 1880
rect 57060 1760 57080 1880
rect 57100 1760 57105 1880
rect 57035 1750 57105 1760
rect 57130 1880 57160 1890
rect 57130 1760 57135 1880
rect 57155 1760 57160 1880
rect 57130 1750 57160 1760
rect 57185 1880 57215 1890
rect 57185 1760 57190 1880
rect 57210 1760 57215 1880
rect 57185 1750 57215 1760
rect 57240 1880 57270 1890
rect 57240 1760 57245 1880
rect 57265 1760 57270 1880
rect 57240 1750 57270 1760
rect 57295 1880 57325 1890
rect 57295 1760 57300 1880
rect 57320 1760 57325 1880
rect 57295 1750 57325 1760
rect 57350 1880 57380 1890
rect 57350 1760 57355 1880
rect 57375 1760 57380 1880
rect 57350 1750 57380 1760
rect 57405 1880 57435 1890
rect 57405 1760 57410 1880
rect 57430 1760 57435 1880
rect 57405 1750 57435 1760
rect 57460 1880 57490 1890
rect 57460 1760 57465 1880
rect 57485 1760 57490 1880
rect 57460 1750 57490 1760
rect 57515 1880 57545 1890
rect 57515 1760 57520 1880
rect 57540 1760 57545 1880
rect 57515 1750 57545 1760
rect 57570 1880 57600 1890
rect 57570 1760 57575 1880
rect 57595 1760 57600 1880
rect 57570 1750 57600 1760
rect 57625 1880 57655 1890
rect 57625 1760 57630 1880
rect 57650 1760 57655 1880
rect 57625 1750 57655 1760
rect 57680 1880 57710 1890
rect 57680 1760 57685 1880
rect 57705 1760 57710 1880
rect 57680 1750 57710 1760
rect 57735 1880 57805 1890
rect 57735 1760 57740 1880
rect 57760 1760 57780 1880
rect 57800 1760 57805 1880
rect 57735 1750 57805 1760
rect 58365 1865 58435 1875
rect 55365 1685 55435 1695
rect 56035 1720 56065 1750
rect 56035 1700 56040 1720
rect 56060 1700 56065 1720
rect 56035 1690 56065 1700
rect 56695 1720 56725 1730
rect 56695 1700 56700 1720
rect 56720 1700 56725 1720
rect 56695 1690 56725 1700
rect 57075 1720 57105 1730
rect 57075 1700 57080 1720
rect 57100 1700 57105 1720
rect 57075 1690 57105 1700
rect 57735 1720 57765 1750
rect 57735 1700 57740 1720
rect 57760 1700 57765 1720
rect 57735 1690 57765 1700
rect 58365 1695 58370 1865
rect 58390 1695 58410 1865
rect 58430 1695 58435 1865
rect 58365 1685 58435 1695
rect 58460 1865 58490 1875
rect 58460 1695 58465 1865
rect 58485 1695 58490 1865
rect 58460 1685 58490 1695
rect 58515 1865 58545 1875
rect 58515 1695 58520 1865
rect 58540 1695 58545 1865
rect 58515 1685 58545 1695
rect 58570 1865 58600 1875
rect 58570 1695 58575 1865
rect 58595 1695 58600 1865
rect 58570 1685 58600 1695
rect 58625 1865 58655 1875
rect 58625 1695 58630 1865
rect 58650 1695 58655 1865
rect 58625 1685 58655 1695
rect 58680 1865 58710 1875
rect 58680 1695 58685 1865
rect 58705 1695 58710 1865
rect 58680 1685 58710 1695
rect 58735 1865 58765 1875
rect 58735 1695 58740 1865
rect 58760 1695 58765 1865
rect 58735 1685 58765 1695
rect 58790 1865 58820 1875
rect 58790 1695 58795 1865
rect 58815 1695 58820 1865
rect 58790 1685 58820 1695
rect 58845 1865 58875 1875
rect 58845 1695 58850 1865
rect 58870 1695 58875 1865
rect 58845 1685 58875 1695
rect 58900 1865 58930 1875
rect 58900 1695 58905 1865
rect 58925 1695 58930 1865
rect 58900 1685 58930 1695
rect 58955 1865 58985 1875
rect 58955 1695 58960 1865
rect 58980 1695 58985 1865
rect 58955 1685 58985 1695
rect 59010 1865 59040 1875
rect 59010 1695 59015 1865
rect 59035 1695 59040 1865
rect 59010 1685 59040 1695
rect 59065 1865 59135 1875
rect 59065 1695 59070 1865
rect 59090 1695 59110 1865
rect 59130 1695 59135 1865
rect 59065 1685 59135 1695
rect 59250 1781 59465 1801
rect 59250 1764 59285 1781
rect 59430 1764 59465 1781
rect 54810 1655 54850 1665
rect 54810 1635 54820 1655
rect 54840 1635 54850 1655
rect 54810 1625 54850 1635
rect 54920 1655 54960 1665
rect 54920 1635 54930 1655
rect 54950 1635 54960 1655
rect 54920 1625 54960 1635
rect 55030 1655 55070 1665
rect 55030 1635 55040 1655
rect 55060 1635 55070 1655
rect 55030 1625 55070 1635
rect 55140 1655 55180 1665
rect 55140 1635 55150 1655
rect 55170 1635 55180 1655
rect 55140 1625 55180 1635
rect 55200 1655 55230 1665
rect 55200 1635 55205 1655
rect 55225 1635 55230 1655
rect 55200 1625 55230 1635
rect 55250 1655 55290 1665
rect 55250 1635 55260 1655
rect 55280 1635 55290 1655
rect 55250 1625 55290 1635
rect 58510 1655 58550 1665
rect 58510 1635 58520 1655
rect 58540 1635 58550 1655
rect 58510 1625 58550 1635
rect 58570 1655 58600 1665
rect 58570 1635 58575 1655
rect 58595 1635 58600 1655
rect 58570 1625 58600 1635
rect 58620 1655 58660 1665
rect 58620 1635 58630 1655
rect 58650 1635 58660 1655
rect 58620 1625 58660 1635
rect 58730 1655 58770 1665
rect 58730 1635 58740 1655
rect 58760 1635 58770 1655
rect 58730 1625 58770 1635
rect 58840 1655 58880 1665
rect 58840 1635 58850 1655
rect 58870 1635 58880 1655
rect 58840 1625 58880 1635
rect 58950 1655 58990 1665
rect 58950 1635 58960 1655
rect 58980 1635 58990 1655
rect 58950 1625 58990 1635
rect 55195 1590 55235 1600
rect 55195 1570 55205 1590
rect 55225 1570 55235 1590
rect 55195 1550 55235 1570
rect 55195 1530 55205 1550
rect 55225 1530 55235 1550
rect 55195 1520 55235 1530
rect 58565 1590 58605 1600
rect 58565 1570 58575 1590
rect 58595 1570 58605 1590
rect 58565 1550 58605 1570
rect 58565 1530 58575 1550
rect 58595 1530 58605 1550
rect 59345 1714 59370 1764
rect 58565 1520 58605 1530
rect 55200 1485 55230 1495
rect 55200 1465 55205 1485
rect 55225 1465 55230 1485
rect 55200 1455 55230 1465
rect 58570 1485 58600 1495
rect 58570 1465 58575 1485
rect 58595 1465 58600 1485
rect 58570 1455 58600 1465
rect 54665 1425 54735 1435
rect 54335 1155 54370 1165
rect 54335 1130 54340 1155
rect 54365 1130 54370 1155
rect 54335 1120 54370 1130
rect 54395 1155 54430 1165
rect 54395 1130 54400 1155
rect 54425 1130 54430 1155
rect 54395 1120 54430 1130
rect 54455 1155 54490 1165
rect 54455 1130 54460 1155
rect 54485 1130 54490 1155
rect 54455 1120 54490 1130
rect 54515 1155 54550 1165
rect 54515 1130 54520 1155
rect 54545 1130 54550 1155
rect 54665 1155 54670 1425
rect 54690 1155 54710 1425
rect 54730 1155 54735 1425
rect 54665 1145 54735 1155
rect 54760 1425 54790 1435
rect 54760 1155 54765 1425
rect 54785 1155 54790 1425
rect 54760 1145 54790 1155
rect 54815 1425 54845 1435
rect 54815 1155 54820 1425
rect 54840 1155 54845 1425
rect 54815 1145 54845 1155
rect 54870 1425 54900 1435
rect 54870 1155 54875 1425
rect 54895 1155 54900 1425
rect 54870 1145 54900 1155
rect 54925 1425 54955 1435
rect 54925 1155 54930 1425
rect 54950 1155 54955 1425
rect 54925 1145 54955 1155
rect 54980 1425 55010 1435
rect 54980 1155 54985 1425
rect 55005 1155 55010 1425
rect 54980 1145 55010 1155
rect 55035 1425 55065 1435
rect 55035 1155 55040 1425
rect 55060 1155 55065 1425
rect 55035 1145 55065 1155
rect 55090 1425 55120 1435
rect 55090 1155 55095 1425
rect 55115 1155 55120 1425
rect 55090 1145 55120 1155
rect 55145 1425 55175 1435
rect 55145 1155 55150 1425
rect 55170 1155 55175 1425
rect 55145 1145 55175 1155
rect 55200 1425 55230 1435
rect 55200 1155 55205 1425
rect 55225 1155 55230 1425
rect 55200 1145 55230 1155
rect 55255 1425 55285 1435
rect 55255 1155 55260 1425
rect 55280 1155 55285 1425
rect 55255 1145 55285 1155
rect 55310 1425 55340 1435
rect 55310 1155 55315 1425
rect 55335 1155 55340 1425
rect 55310 1145 55340 1155
rect 55365 1425 55435 1435
rect 55365 1155 55370 1425
rect 55390 1155 55410 1425
rect 55430 1155 55435 1425
rect 58365 1425 58435 1435
rect 56690 1300 56720 1310
rect 56040 1290 56070 1300
rect 56040 1270 56045 1290
rect 56065 1270 56070 1290
rect 56690 1280 56695 1300
rect 56715 1280 56720 1300
rect 56690 1270 56720 1280
rect 56840 1300 56870 1310
rect 56840 1280 56845 1300
rect 56865 1280 56870 1300
rect 56840 1270 56870 1280
rect 56930 1300 56960 1310
rect 56930 1280 56935 1300
rect 56955 1280 56960 1300
rect 56930 1270 56960 1280
rect 57080 1300 57110 1310
rect 57080 1280 57085 1300
rect 57105 1280 57110 1300
rect 57080 1270 57110 1280
rect 57730 1290 57760 1300
rect 57730 1270 57735 1290
rect 57755 1270 57760 1290
rect 56040 1260 56070 1270
rect 57730 1260 57760 1270
rect 55365 1145 55435 1155
rect 55995 1205 56065 1215
rect 54515 1120 54550 1130
rect 54705 1115 54735 1125
rect 54705 1095 54710 1115
rect 54730 1095 54735 1115
rect 54705 1080 54735 1095
rect 55365 1115 55395 1125
rect 55365 1095 55370 1115
rect 55390 1095 55395 1115
rect 55365 1080 55395 1095
rect 55995 1085 56000 1205
rect 56020 1085 56040 1205
rect 56060 1085 56065 1205
rect 55995 1075 56065 1085
rect 56090 1205 56120 1215
rect 56090 1085 56095 1205
rect 56115 1085 56120 1205
rect 56090 1075 56120 1085
rect 56145 1205 56175 1215
rect 56145 1085 56150 1205
rect 56170 1085 56175 1205
rect 56145 1075 56175 1085
rect 56200 1205 56230 1215
rect 56200 1085 56205 1205
rect 56225 1085 56230 1205
rect 56200 1075 56230 1085
rect 56255 1205 56285 1215
rect 56255 1085 56260 1205
rect 56280 1085 56285 1205
rect 56255 1075 56285 1085
rect 56310 1205 56340 1215
rect 56310 1085 56315 1205
rect 56335 1085 56340 1205
rect 56310 1075 56340 1085
rect 56365 1205 56395 1215
rect 56365 1085 56370 1205
rect 56390 1085 56395 1205
rect 56365 1075 56395 1085
rect 56420 1205 56450 1215
rect 56420 1085 56425 1205
rect 56445 1085 56450 1205
rect 56420 1075 56450 1085
rect 56475 1205 56505 1215
rect 56475 1085 56480 1205
rect 56500 1085 56505 1205
rect 56475 1075 56505 1085
rect 56530 1205 56560 1215
rect 56530 1085 56535 1205
rect 56555 1085 56560 1205
rect 56530 1075 56560 1085
rect 56585 1205 56615 1215
rect 56585 1085 56590 1205
rect 56610 1085 56615 1205
rect 56585 1075 56615 1085
rect 56640 1205 56670 1215
rect 56640 1085 56645 1205
rect 56665 1085 56670 1205
rect 56640 1075 56670 1085
rect 56695 1205 56805 1215
rect 56695 1085 56700 1205
rect 56720 1085 56740 1205
rect 56760 1085 56780 1205
rect 56800 1085 56805 1205
rect 56695 1075 56805 1085
rect 56830 1205 56860 1215
rect 56830 1085 56835 1205
rect 56855 1085 56860 1205
rect 56830 1075 56860 1085
rect 56885 1205 56915 1215
rect 56885 1085 56890 1205
rect 56910 1085 56915 1205
rect 56885 1075 56915 1085
rect 56940 1205 56970 1215
rect 56940 1085 56945 1205
rect 56965 1085 56970 1205
rect 56940 1075 56970 1085
rect 56995 1205 57105 1215
rect 56995 1085 57000 1205
rect 57020 1085 57040 1205
rect 57060 1085 57080 1205
rect 57100 1085 57105 1205
rect 56995 1075 57105 1085
rect 57130 1205 57160 1215
rect 57130 1085 57135 1205
rect 57155 1085 57160 1205
rect 57130 1075 57160 1085
rect 57185 1205 57215 1215
rect 57185 1085 57190 1205
rect 57210 1085 57215 1205
rect 57185 1075 57215 1085
rect 57240 1205 57270 1215
rect 57240 1085 57245 1205
rect 57265 1085 57270 1205
rect 57240 1075 57270 1085
rect 57295 1205 57325 1215
rect 57295 1085 57300 1205
rect 57320 1085 57325 1205
rect 57295 1075 57325 1085
rect 57350 1205 57380 1215
rect 57350 1085 57355 1205
rect 57375 1085 57380 1205
rect 57350 1075 57380 1085
rect 57405 1205 57435 1215
rect 57405 1085 57410 1205
rect 57430 1085 57435 1205
rect 57405 1075 57435 1085
rect 57460 1205 57490 1215
rect 57460 1085 57465 1205
rect 57485 1085 57490 1205
rect 57460 1075 57490 1085
rect 57515 1205 57545 1215
rect 57515 1085 57520 1205
rect 57540 1085 57545 1205
rect 57515 1075 57545 1085
rect 57570 1205 57600 1215
rect 57570 1085 57575 1205
rect 57595 1085 57600 1205
rect 57570 1075 57600 1085
rect 57625 1205 57655 1215
rect 57625 1085 57630 1205
rect 57650 1085 57655 1205
rect 57625 1075 57655 1085
rect 57680 1205 57710 1215
rect 57680 1085 57685 1205
rect 57705 1085 57710 1205
rect 57680 1075 57710 1085
rect 57735 1205 57805 1215
rect 57735 1085 57740 1205
rect 57760 1085 57780 1205
rect 57800 1085 57805 1205
rect 58365 1155 58370 1425
rect 58390 1155 58410 1425
rect 58430 1155 58435 1425
rect 58365 1145 58435 1155
rect 58460 1425 58490 1435
rect 58460 1155 58465 1425
rect 58485 1155 58490 1425
rect 58460 1145 58490 1155
rect 58515 1425 58545 1435
rect 58515 1155 58520 1425
rect 58540 1155 58545 1425
rect 58515 1145 58545 1155
rect 58570 1425 58600 1435
rect 58570 1155 58575 1425
rect 58595 1155 58600 1425
rect 58570 1145 58600 1155
rect 58625 1425 58655 1435
rect 58625 1155 58630 1425
rect 58650 1155 58655 1425
rect 58625 1145 58655 1155
rect 58680 1425 58710 1435
rect 58680 1155 58685 1425
rect 58705 1155 58710 1425
rect 58680 1145 58710 1155
rect 58735 1425 58765 1435
rect 58735 1155 58740 1425
rect 58760 1155 58765 1425
rect 58735 1145 58765 1155
rect 58790 1425 58820 1435
rect 58790 1155 58795 1425
rect 58815 1155 58820 1425
rect 58790 1145 58820 1155
rect 58845 1425 58875 1435
rect 58845 1155 58850 1425
rect 58870 1155 58875 1425
rect 58845 1145 58875 1155
rect 58900 1425 58930 1435
rect 58900 1155 58905 1425
rect 58925 1155 58930 1425
rect 58900 1145 58930 1155
rect 58955 1425 58985 1435
rect 58955 1155 58960 1425
rect 58980 1155 58985 1425
rect 58955 1145 58985 1155
rect 59010 1425 59040 1435
rect 59010 1155 59015 1425
rect 59035 1155 59040 1425
rect 59010 1145 59040 1155
rect 59065 1425 59135 1435
rect 59065 1155 59070 1425
rect 59090 1155 59110 1425
rect 59130 1155 59135 1425
rect 59065 1145 59135 1155
rect 59250 1155 59285 1165
rect 59250 1130 59255 1155
rect 59280 1130 59285 1155
rect 57735 1075 57805 1085
rect 58405 1115 58435 1125
rect 58405 1095 58410 1115
rect 58430 1095 58435 1115
rect 58405 1080 58435 1095
rect 59065 1115 59095 1125
rect 59250 1120 59285 1130
rect 59310 1155 59345 1165
rect 59310 1130 59315 1155
rect 59340 1130 59345 1155
rect 59310 1120 59345 1130
rect 59370 1155 59405 1165
rect 59370 1130 59375 1155
rect 59400 1130 59405 1155
rect 59370 1120 59405 1130
rect 59430 1155 59465 1165
rect 59430 1130 59435 1155
rect 59460 1130 59465 1155
rect 59430 1120 59465 1130
rect 59065 1095 59070 1115
rect 59090 1095 59095 1115
rect 59065 1085 59095 1095
rect 56040 1055 56065 1075
rect 56035 1045 56065 1055
rect 56035 1025 56040 1045
rect 56060 1025 56065 1045
rect 56035 1015 56065 1025
rect 56735 1045 56765 1055
rect 56735 1025 56740 1045
rect 56760 1025 56765 1045
rect 56735 1015 56765 1025
rect 57035 1045 57065 1055
rect 57035 1025 57040 1045
rect 57060 1025 57065 1045
rect 57035 1015 57065 1025
rect 57735 1045 57765 1075
rect 57735 1025 57740 1045
rect 57760 1025 57765 1045
rect 57735 1015 57765 1025
rect 55080 430 55120 440
rect 55080 410 55090 430
rect 55110 410 55120 430
rect 55080 400 55120 410
rect 58680 430 58720 440
rect 58680 410 58690 430
rect 58710 410 58720 430
rect 58680 400 58720 410
rect 56825 375 56865 385
rect 56825 355 56835 375
rect 56855 355 56865 375
rect 56825 345 56865 355
rect 56935 375 56975 385
rect 56935 355 56945 375
rect 56965 355 56975 375
rect 56935 345 56975 355
rect 56185 315 56255 325
rect 54405 170 54440 180
rect 54405 145 54410 170
rect 54435 145 54440 170
rect 54405 135 54440 145
rect 54465 170 54500 180
rect 54465 145 54470 170
rect 54495 145 54500 170
rect 54465 135 54500 145
rect 54695 165 54765 175
rect 54440 -552 54465 -502
rect 54695 -505 54700 165
rect 54720 -505 54740 165
rect 54760 -505 54765 165
rect 54695 -515 54765 -505
rect 54835 165 54865 175
rect 54835 -505 54840 165
rect 54860 -505 54865 165
rect 54835 -515 54865 -505
rect 54935 165 54965 175
rect 54935 -505 54940 165
rect 54960 -505 54965 165
rect 54935 -515 54965 -505
rect 55035 165 55065 175
rect 55035 -505 55040 165
rect 55060 -505 55065 165
rect 55035 -515 55065 -505
rect 55135 165 55165 175
rect 55135 -505 55140 165
rect 55160 -505 55165 165
rect 55135 -515 55165 -505
rect 55235 165 55265 175
rect 55235 -505 55240 165
rect 55260 -505 55265 165
rect 55235 -515 55265 -505
rect 55335 165 55405 175
rect 55335 -505 55340 165
rect 55360 -505 55380 165
rect 55400 -505 55405 165
rect 56185 95 56190 315
rect 56210 95 56230 315
rect 56250 95 56255 315
rect 56185 85 56255 95
rect 56280 315 56310 325
rect 56280 95 56285 315
rect 56305 95 56310 315
rect 56280 85 56310 95
rect 56335 315 56365 325
rect 56335 95 56340 315
rect 56360 95 56365 315
rect 56335 85 56365 95
rect 56390 315 56420 325
rect 56390 95 56395 315
rect 56415 95 56420 315
rect 56390 85 56420 95
rect 56445 315 56475 325
rect 56445 95 56450 315
rect 56470 95 56475 315
rect 56445 85 56475 95
rect 56500 315 56530 325
rect 56500 95 56505 315
rect 56525 95 56530 315
rect 56500 85 56530 95
rect 56555 315 56585 325
rect 56555 95 56560 315
rect 56580 95 56585 315
rect 56555 85 56585 95
rect 56610 315 56640 325
rect 56610 95 56615 315
rect 56635 95 56640 315
rect 56610 85 56640 95
rect 56665 315 56695 325
rect 56665 95 56670 315
rect 56690 95 56695 315
rect 56665 85 56695 95
rect 56720 315 56750 325
rect 56720 95 56725 315
rect 56745 95 56750 315
rect 56720 85 56750 95
rect 56775 315 56805 325
rect 56775 95 56780 315
rect 56800 95 56805 315
rect 56775 85 56805 95
rect 56830 315 56860 325
rect 56830 95 56835 315
rect 56855 95 56860 315
rect 56830 85 56860 95
rect 56885 315 56915 325
rect 56885 95 56890 315
rect 56910 95 56915 315
rect 56885 85 56915 95
rect 56940 315 56970 325
rect 56940 95 56945 315
rect 56965 95 56970 315
rect 56940 85 56970 95
rect 56995 315 57025 325
rect 56995 95 57000 315
rect 57020 95 57025 315
rect 56995 85 57025 95
rect 57050 315 57080 325
rect 57050 95 57055 315
rect 57075 95 57080 315
rect 57050 85 57080 95
rect 57105 315 57135 325
rect 57105 95 57110 315
rect 57130 95 57135 315
rect 57105 85 57135 95
rect 57160 315 57190 325
rect 57160 95 57165 315
rect 57185 95 57190 315
rect 57160 85 57190 95
rect 57215 315 57245 325
rect 57215 95 57220 315
rect 57240 95 57245 315
rect 57215 85 57245 95
rect 57270 315 57300 325
rect 57270 95 57275 315
rect 57295 95 57300 315
rect 57270 85 57300 95
rect 57325 315 57355 325
rect 57325 95 57330 315
rect 57350 95 57355 315
rect 57325 85 57355 95
rect 57380 315 57410 325
rect 57380 95 57385 315
rect 57405 95 57410 315
rect 57380 85 57410 95
rect 57435 315 57465 325
rect 57435 95 57440 315
rect 57460 95 57465 315
rect 57435 85 57465 95
rect 57490 315 57560 325
rect 57490 95 57495 315
rect 57515 95 57535 315
rect 57555 95 57560 315
rect 57490 85 57560 95
rect 58395 165 58465 175
rect 56220 55 56260 65
rect 56220 35 56230 55
rect 56250 35 56260 55
rect 56220 25 56260 35
rect 57485 55 57525 65
rect 57485 35 57495 55
rect 57515 35 57525 55
rect 57485 25 57525 35
rect 57415 -45 57455 -35
rect 57415 -65 57425 -45
rect 57445 -65 57455 -45
rect 57415 -75 57455 -65
rect 56595 -280 56635 -270
rect 56595 -300 56605 -280
rect 56625 -300 56635 -280
rect 56595 -310 56635 -300
rect 57040 -280 57080 -270
rect 57040 -300 57050 -280
rect 57070 -300 57080 -280
rect 57040 -310 57080 -300
rect 56395 -340 56465 -330
rect 56395 -460 56400 -340
rect 56420 -460 56440 -340
rect 56460 -460 56465 -340
rect 56395 -470 56465 -460
rect 56490 -340 56520 -330
rect 56490 -460 56495 -340
rect 56515 -460 56520 -340
rect 56490 -470 56520 -460
rect 56545 -340 56575 -330
rect 56545 -460 56550 -340
rect 56570 -460 56575 -340
rect 56545 -470 56575 -460
rect 56600 -340 56630 -330
rect 56600 -460 56605 -340
rect 56625 -460 56630 -340
rect 56600 -470 56630 -460
rect 56655 -340 56685 -330
rect 56655 -460 56660 -340
rect 56680 -460 56685 -340
rect 56655 -470 56685 -460
rect 56710 -340 56740 -330
rect 56710 -460 56715 -340
rect 56735 -460 56740 -340
rect 56710 -470 56740 -460
rect 56765 -340 56835 -330
rect 56765 -460 56770 -340
rect 56790 -460 56810 -340
rect 56830 -460 56835 -340
rect 56765 -470 56835 -460
rect 56875 -340 56905 -330
rect 56875 -460 56880 -340
rect 56900 -460 56905 -340
rect 56875 -470 56905 -460
rect 57215 -340 57245 -330
rect 57215 -460 57220 -340
rect 57240 -460 57245 -340
rect 57215 -470 57245 -460
rect 55335 -515 55405 -505
rect 56435 -500 56465 -490
rect 56435 -520 56440 -500
rect 56460 -520 56465 -500
rect 56435 -530 56465 -520
rect 56765 -500 56795 -490
rect 56765 -520 56770 -500
rect 56790 -520 56795 -500
rect 58395 -505 58400 165
rect 58420 -505 58440 165
rect 58460 -505 58465 165
rect 58395 -515 58465 -505
rect 58535 165 58565 175
rect 58535 -505 58540 165
rect 58560 -505 58565 165
rect 58535 -515 58565 -505
rect 58635 165 58665 175
rect 58635 -505 58640 165
rect 58660 -505 58665 165
rect 58635 -515 58665 -505
rect 58735 165 58765 175
rect 58735 -505 58740 165
rect 58760 -505 58765 165
rect 58735 -515 58765 -505
rect 58835 165 58865 175
rect 58835 -505 58840 165
rect 58860 -505 58865 165
rect 58835 -515 58865 -505
rect 58935 165 58965 175
rect 58935 -505 58940 165
rect 58960 -505 58965 165
rect 58935 -515 58965 -505
rect 59035 165 59105 175
rect 59035 -505 59040 165
rect 59060 -505 59080 165
rect 59100 -505 59105 165
rect 59300 170 59335 180
rect 59300 145 59305 170
rect 59330 145 59335 170
rect 59300 135 59335 145
rect 59360 170 59395 180
rect 59360 145 59365 170
rect 59390 145 59395 170
rect 59360 135 59395 145
rect 59035 -515 59105 -505
rect 56765 -530 56795 -520
rect 54735 -545 54765 -535
rect 54735 -565 54740 -545
rect 54760 -565 54765 -545
rect 54735 -575 54765 -565
rect 55335 -545 55365 -535
rect 55335 -565 55340 -545
rect 55360 -565 55365 -545
rect 55335 -575 55365 -565
rect 58435 -545 58465 -535
rect 58435 -565 58440 -545
rect 58460 -565 58465 -545
rect 58435 -575 58465 -565
rect 59035 -545 59065 -535
rect 59035 -565 59040 -545
rect 59060 -565 59065 -545
rect 59335 -552 59360 -502
rect 59035 -575 59065 -565
<< viali >>
rect 56095 4905 56115 4925
rect 56275 4905 56295 4925
rect 57035 4905 57055 4925
rect 57215 4905 57235 4925
rect 57505 4905 57525 4925
rect 57685 4905 57705 4925
rect 56095 4545 56115 4865
rect 56155 4545 56175 4865
rect 56215 4545 56235 4865
rect 56275 4545 56295 4865
rect 56565 4735 56585 4755
rect 56745 4735 56765 4755
rect 56565 4545 56585 4695
rect 56625 4545 56645 4695
rect 56685 4545 56705 4695
rect 56745 4545 56765 4695
rect 57035 4545 57055 4865
rect 57095 4545 57115 4865
rect 57155 4545 57175 4865
rect 57215 4545 57235 4865
rect 57505 4545 57525 4865
rect 57565 4545 57585 4865
rect 57625 4545 57645 4865
rect 57685 4545 57705 4865
rect 56160 4455 56180 4475
rect 56635 4455 56655 4475
rect 57145 4455 57165 4475
rect 57581 4445 57601 4465
rect 54680 3680 54700 4000
rect 54740 3680 54760 4000
rect 54800 3680 54820 4000
rect 54860 3680 54880 4000
rect 54920 3680 54940 4000
rect 54980 3680 55000 4000
rect 55040 3680 55060 4000
rect 55100 3680 55120 4000
rect 55160 3680 55180 4000
rect 55220 3680 55240 4000
rect 55280 3680 55300 4000
rect 55340 3680 55360 4000
rect 55400 3680 55420 4000
rect 56015 3680 56035 4000
rect 56075 3680 56095 4000
rect 56135 3680 56155 4000
rect 56195 3680 56215 4000
rect 56255 3680 56275 4000
rect 56315 3680 56335 4000
rect 56375 3680 56395 4000
rect 56435 3680 56455 4000
rect 56495 3680 56515 4000
rect 56555 3680 56575 4000
rect 56615 3680 56635 4000
rect 56675 3680 56695 4000
rect 56735 3680 56755 4000
rect 57045 3680 57065 4000
rect 57105 3680 57125 4000
rect 57165 3680 57185 4000
rect 57225 3680 57245 4000
rect 57285 3680 57305 4000
rect 57345 3680 57365 4000
rect 57405 3680 57425 4000
rect 57465 3680 57485 4000
rect 57525 3680 57545 4000
rect 57585 3680 57605 4000
rect 57645 3680 57665 4000
rect 57705 3680 57725 4000
rect 57765 3680 57785 4000
rect 58380 3680 58400 4000
rect 58440 3680 58460 4000
rect 58500 3680 58520 4000
rect 58560 3680 58580 4000
rect 58620 3680 58640 4000
rect 58680 3680 58700 4000
rect 58740 3680 58760 4000
rect 58800 3680 58820 4000
rect 58860 3680 58880 4000
rect 58920 3680 58940 4000
rect 58980 3680 59000 4000
rect 59040 3680 59060 4000
rect 59100 3680 59120 4000
rect 54680 3620 54700 3640
rect 55400 3620 55420 3640
rect 56015 3620 56035 3640
rect 56735 3620 56755 3640
rect 57045 3620 57065 3640
rect 57765 3620 57785 3640
rect 58380 3620 58400 3640
rect 59100 3620 59120 3640
rect 56375 3555 56395 3575
rect 57405 3555 57425 3575
rect 55040 3510 55060 3530
rect 58740 3510 58760 3530
rect 54210 3270 54230 3290
rect 54265 3270 54285 3290
rect 54320 3270 54340 3290
rect 56520 3240 56540 3260
rect 56685 3240 56705 3260
rect 56850 3240 56870 3260
rect 56930 3240 56950 3260
rect 57095 3240 57115 3260
rect 57260 3240 57280 3260
rect 54710 3180 54730 3200
rect 55370 3180 55390 3200
rect 56630 3185 56650 3205
rect 56740 3185 56760 3205
rect 57040 3185 57060 3205
rect 57150 3185 57170 3205
rect 58410 3180 58430 3200
rect 59070 3180 59090 3200
rect 59460 3185 59480 3205
rect 59515 3185 59535 3205
rect 59570 3185 59590 3205
rect 54210 2665 54230 2685
rect 54265 2665 54285 2685
rect 54320 2665 54340 2685
rect 54710 2570 54730 3140
rect 54765 2570 54785 3140
rect 54820 2570 54840 3140
rect 54875 2570 54895 3140
rect 54930 2570 54950 3140
rect 54985 2570 55005 3140
rect 55040 2570 55060 3140
rect 55095 2570 55115 3140
rect 55150 2570 55170 3140
rect 55205 2570 55225 3140
rect 55260 2570 55280 3140
rect 55315 2570 55335 3140
rect 55370 2570 55390 3140
rect 56565 2875 56585 2895
rect 56612 2865 56632 2885
rect 56685 2865 56705 2885
rect 56758 2865 56778 2885
rect 56805 2875 56825 2895
rect 56975 2875 56995 2895
rect 57022 2865 57042 2885
rect 57095 2865 57115 2885
rect 57168 2865 57188 2885
rect 57215 2875 57235 2895
rect 56610 2805 56630 2825
rect 57170 2805 57190 2825
rect 56860 2590 56880 2610
rect 56945 2590 56965 2610
rect 58410 2570 58430 3140
rect 58465 2570 58485 3140
rect 58520 2570 58540 3140
rect 58575 2570 58595 3140
rect 58630 2570 58650 3140
rect 58685 2570 58705 3140
rect 58740 2570 58760 3140
rect 58795 2570 58815 3140
rect 58850 2570 58870 3140
rect 58905 2570 58925 3140
rect 58960 2570 58980 3140
rect 59015 2570 59035 3140
rect 59070 2570 59090 3140
rect 59460 2580 59480 2600
rect 59515 2580 59535 2600
rect 59570 2580 59590 2600
rect 55040 2445 55060 2465
rect 55040 2405 55060 2425
rect 55040 2365 55060 2385
rect 56780 2330 56800 2550
rect 56835 2330 56855 2550
rect 56890 2330 56910 2550
rect 56945 2330 56965 2550
rect 57000 2330 57020 2550
rect 58740 2445 58760 2465
rect 58740 2405 58760 2425
rect 58740 2365 58760 2385
rect 56780 2270 56800 2290
rect 57000 2270 57020 2290
rect 56000 1960 56020 1980
rect 56695 1960 56715 1980
rect 57085 1960 57105 1980
rect 54710 1905 54730 1925
rect 55370 1905 55390 1925
rect 58410 1905 58430 1925
rect 59070 1905 59090 1925
rect 54710 1695 54730 1865
rect 54765 1695 54785 1865
rect 54820 1695 54840 1865
rect 54875 1695 54895 1865
rect 54930 1695 54950 1865
rect 54985 1695 55005 1865
rect 55040 1695 55060 1865
rect 55095 1695 55115 1865
rect 55150 1695 55170 1865
rect 55205 1695 55225 1865
rect 55260 1695 55280 1865
rect 55315 1695 55335 1865
rect 55370 1695 55390 1865
rect 56040 1760 56060 1880
rect 56095 1760 56115 1880
rect 56150 1760 56170 1880
rect 56205 1760 56225 1880
rect 56260 1760 56280 1880
rect 56315 1760 56335 1880
rect 56370 1760 56390 1880
rect 56425 1760 56445 1880
rect 56480 1760 56500 1880
rect 56535 1760 56555 1880
rect 56590 1760 56610 1880
rect 56645 1760 56665 1880
rect 56700 1760 56720 1880
rect 57080 1760 57100 1880
rect 57135 1760 57155 1880
rect 57190 1760 57210 1880
rect 57245 1760 57265 1880
rect 57300 1760 57320 1880
rect 57355 1760 57375 1880
rect 57410 1760 57430 1880
rect 57465 1760 57485 1880
rect 57520 1760 57540 1880
rect 57575 1760 57595 1880
rect 57630 1760 57650 1880
rect 57685 1760 57705 1880
rect 57740 1760 57760 1880
rect 56040 1700 56060 1720
rect 56700 1700 56720 1720
rect 57080 1700 57100 1720
rect 57740 1700 57760 1720
rect 58410 1695 58430 1865
rect 58465 1695 58485 1865
rect 58520 1695 58540 1865
rect 58575 1695 58595 1865
rect 58630 1695 58650 1865
rect 58685 1695 58705 1865
rect 58740 1695 58760 1865
rect 58795 1695 58815 1865
rect 58850 1695 58870 1865
rect 58905 1695 58925 1865
rect 58960 1695 58980 1865
rect 59015 1695 59035 1865
rect 59070 1695 59090 1865
rect 54820 1635 54840 1655
rect 54930 1635 54950 1655
rect 55040 1635 55060 1655
rect 55150 1635 55170 1655
rect 55260 1635 55280 1655
rect 58520 1635 58540 1655
rect 58630 1635 58650 1655
rect 58740 1635 58760 1655
rect 58850 1635 58870 1655
rect 58960 1635 58980 1655
rect 55205 1570 55225 1590
rect 55205 1530 55225 1550
rect 58575 1570 58595 1590
rect 58575 1530 58595 1550
rect 54340 1130 54365 1155
rect 54400 1130 54425 1155
rect 54460 1130 54485 1155
rect 54520 1130 54545 1155
rect 54710 1155 54730 1425
rect 54765 1155 54785 1425
rect 54820 1155 54840 1425
rect 54875 1155 54895 1425
rect 54930 1155 54950 1425
rect 54985 1155 55005 1425
rect 55040 1155 55060 1425
rect 55095 1155 55115 1425
rect 55150 1155 55170 1425
rect 55205 1155 55225 1425
rect 55260 1155 55280 1425
rect 55315 1155 55335 1425
rect 55370 1155 55390 1425
rect 56045 1270 56065 1290
rect 56695 1280 56715 1300
rect 56845 1280 56865 1300
rect 56935 1280 56955 1300
rect 57085 1280 57105 1300
rect 57735 1270 57755 1290
rect 54710 1095 54730 1115
rect 55370 1095 55390 1115
rect 56040 1085 56060 1205
rect 56095 1085 56115 1205
rect 56150 1085 56170 1205
rect 56205 1085 56225 1205
rect 56260 1085 56280 1205
rect 56315 1085 56335 1205
rect 56370 1085 56390 1205
rect 56425 1085 56445 1205
rect 56480 1085 56500 1205
rect 56535 1085 56555 1205
rect 56590 1085 56610 1205
rect 56645 1085 56665 1205
rect 56700 1085 56720 1205
rect 56780 1085 56800 1205
rect 56835 1085 56855 1205
rect 56890 1085 56910 1205
rect 56945 1085 56965 1205
rect 57000 1085 57020 1205
rect 57080 1085 57100 1205
rect 57135 1085 57155 1205
rect 57190 1085 57210 1205
rect 57245 1085 57265 1205
rect 57300 1085 57320 1205
rect 57355 1085 57375 1205
rect 57410 1085 57430 1205
rect 57465 1085 57485 1205
rect 57520 1085 57540 1205
rect 57575 1085 57595 1205
rect 57630 1085 57650 1205
rect 57685 1085 57705 1205
rect 57740 1085 57760 1205
rect 58410 1155 58430 1425
rect 58465 1155 58485 1425
rect 58520 1155 58540 1425
rect 58575 1155 58595 1425
rect 58630 1155 58650 1425
rect 58685 1155 58705 1425
rect 58740 1155 58760 1425
rect 58795 1155 58815 1425
rect 58850 1155 58870 1425
rect 58905 1155 58925 1425
rect 58960 1155 58980 1425
rect 59015 1155 59035 1425
rect 59070 1155 59090 1425
rect 59255 1130 59280 1155
rect 58410 1095 58430 1115
rect 59315 1130 59340 1155
rect 59375 1130 59400 1155
rect 59435 1130 59460 1155
rect 59070 1095 59090 1115
rect 56040 1025 56060 1045
rect 56740 1025 56760 1045
rect 57040 1025 57060 1045
rect 57740 1025 57760 1045
rect 55090 410 55110 430
rect 58690 410 58710 430
rect 56835 355 56855 375
rect 56945 355 56965 375
rect 54410 145 54435 170
rect 54470 145 54495 170
rect 54740 -505 54760 165
rect 54840 -505 54860 165
rect 54940 -505 54960 165
rect 55040 -505 55060 165
rect 55140 -505 55160 165
rect 55240 -505 55260 165
rect 55340 -505 55360 165
rect 56230 95 56250 315
rect 56285 95 56305 315
rect 56340 95 56360 315
rect 56395 95 56415 315
rect 56450 95 56470 315
rect 56505 95 56525 315
rect 56560 95 56580 315
rect 56615 95 56635 315
rect 56670 95 56690 315
rect 56725 95 56745 315
rect 56780 95 56800 315
rect 56835 95 56855 315
rect 56890 95 56910 315
rect 56945 95 56965 315
rect 57000 95 57020 315
rect 57055 95 57075 315
rect 57110 95 57130 315
rect 57165 95 57185 315
rect 57220 95 57240 315
rect 57275 95 57295 315
rect 57330 95 57350 315
rect 57385 95 57405 315
rect 57440 95 57460 315
rect 57495 95 57515 315
rect 56230 35 56250 55
rect 57495 35 57515 55
rect 57425 -65 57445 -45
rect 56605 -300 56625 -280
rect 57050 -300 57070 -280
rect 56440 -460 56460 -340
rect 56495 -460 56515 -340
rect 56550 -460 56570 -340
rect 56605 -460 56625 -340
rect 56660 -460 56680 -340
rect 56715 -460 56735 -340
rect 56770 -460 56790 -340
rect 56880 -460 56900 -340
rect 57220 -460 57240 -340
rect 56440 -520 56460 -500
rect 56770 -520 56790 -500
rect 58440 -505 58460 165
rect 58540 -505 58560 165
rect 58640 -505 58660 165
rect 58740 -505 58760 165
rect 58840 -505 58860 165
rect 58940 -505 58960 165
rect 59040 -505 59060 165
rect 59305 145 59330 170
rect 59365 145 59390 170
rect 54740 -565 54760 -545
rect 55340 -565 55360 -545
rect 58440 -565 58460 -545
rect 59040 -565 59060 -545
<< metal1 >>
rect 52290 4320 52410 6110
rect 52290 4290 52295 4320
rect 52325 4290 52335 4320
rect 52365 4290 52375 4320
rect 52405 4290 52410 4320
rect 52290 4280 52410 4290
rect 52290 4250 52295 4280
rect 52325 4250 52335 4280
rect 52365 4250 52375 4280
rect 52405 4250 52410 4280
rect 52290 4240 52410 4250
rect 52290 4210 52295 4240
rect 52325 4210 52335 4240
rect 52365 4210 52375 4240
rect 52405 4210 52410 4240
rect 52290 4205 52410 4210
rect 52640 4320 52760 6110
rect 52640 4290 52645 4320
rect 52675 4290 52685 4320
rect 52715 4290 52725 4320
rect 52755 4290 52760 4320
rect 52640 4280 52760 4290
rect 52640 4250 52645 4280
rect 52675 4250 52685 4280
rect 52715 4250 52725 4280
rect 52755 4250 52760 4280
rect 52640 4240 52760 4250
rect 52640 4210 52645 4240
rect 52675 4210 52685 4240
rect 52715 4210 52725 4240
rect 52755 4210 52760 4240
rect 52640 4205 52760 4210
rect 52990 4320 53110 6110
rect 52990 4290 52995 4320
rect 53025 4290 53035 4320
rect 53065 4290 53075 4320
rect 53105 4290 53110 4320
rect 52990 4280 53110 4290
rect 52990 4250 52995 4280
rect 53025 4250 53035 4280
rect 53065 4250 53075 4280
rect 53105 4250 53110 4280
rect 52990 4240 53110 4250
rect 52990 4210 52995 4240
rect 53025 4210 53035 4240
rect 53065 4210 53075 4240
rect 53105 4210 53110 4240
rect 52990 4205 53110 4210
rect 53690 4320 53810 6110
rect 53690 4290 53695 4320
rect 53725 4290 53735 4320
rect 53765 4290 53775 4320
rect 53805 4290 53810 4320
rect 53690 4280 53810 4290
rect 53690 4250 53695 4280
rect 53725 4250 53735 4280
rect 53765 4250 53775 4280
rect 53805 4250 53810 4280
rect 53690 4240 53810 4250
rect 53690 4210 53695 4240
rect 53725 4210 53735 4240
rect 53765 4210 53775 4240
rect 53805 4210 53810 4240
rect 53690 4205 53810 4210
rect 54040 4320 54160 6110
rect 56205 5065 56245 5070
rect 56205 5035 56210 5065
rect 56240 5035 56245 5065
rect 56085 4930 56125 4935
rect 56085 4900 56090 4930
rect 56120 4900 56125 4930
rect 56085 4895 56125 4900
rect 56205 4930 56245 5035
rect 56675 5065 56715 5070
rect 56675 5035 56680 5065
rect 56710 5035 56715 5065
rect 56675 5030 56715 5035
rect 57085 5065 57125 5070
rect 57085 5035 57090 5065
rect 57120 5035 57125 5065
rect 57085 5030 57125 5035
rect 57555 5065 57595 5070
rect 57555 5035 57560 5065
rect 57590 5035 57595 5065
rect 56205 4900 56210 4930
rect 56240 4900 56245 4930
rect 56205 4895 56245 4900
rect 56265 4930 56305 4935
rect 56265 4900 56270 4930
rect 56300 4900 56305 4930
rect 56265 4895 56305 4900
rect 56090 4865 56120 4895
rect 56090 4545 56095 4865
rect 56115 4545 56120 4865
rect 56090 4535 56120 4545
rect 56150 4865 56180 4875
rect 56150 4545 56155 4865
rect 56175 4545 56180 4865
rect 56150 4485 56180 4545
rect 56210 4865 56240 4895
rect 56210 4545 56215 4865
rect 56235 4545 56240 4865
rect 56210 4530 56240 4545
rect 56270 4865 56300 4895
rect 56270 4545 56275 4865
rect 56295 4545 56300 4865
rect 56555 4840 56595 4845
rect 56555 4810 56560 4840
rect 56590 4810 56595 4840
rect 56555 4800 56595 4810
rect 56555 4770 56560 4800
rect 56590 4770 56595 4800
rect 56555 4760 56595 4770
rect 56555 4730 56560 4760
rect 56590 4730 56595 4760
rect 56555 4725 56595 4730
rect 56615 4840 56655 4845
rect 56615 4810 56620 4840
rect 56650 4810 56655 4840
rect 56615 4800 56655 4810
rect 56615 4770 56620 4800
rect 56650 4770 56655 4800
rect 56615 4760 56655 4770
rect 56615 4730 56620 4760
rect 56650 4730 56655 4760
rect 56615 4725 56655 4730
rect 56270 4535 56300 4545
rect 56560 4695 56590 4725
rect 56560 4545 56565 4695
rect 56585 4545 56590 4695
rect 56560 4535 56590 4545
rect 56620 4695 56650 4725
rect 56620 4545 56625 4695
rect 56645 4545 56650 4695
rect 56620 4535 56650 4545
rect 56680 4695 56710 5030
rect 56880 5010 56920 5015
rect 56880 4980 56885 5010
rect 56915 4980 56920 5010
rect 56880 4970 56920 4980
rect 56880 4940 56885 4970
rect 56915 4940 56920 4970
rect 56880 4930 56920 4940
rect 56880 4900 56885 4930
rect 56915 4900 56920 4930
rect 56735 4840 56775 4845
rect 56735 4810 56740 4840
rect 56770 4810 56775 4840
rect 56735 4800 56775 4810
rect 56735 4770 56740 4800
rect 56770 4770 56775 4800
rect 56735 4760 56775 4770
rect 56735 4730 56740 4760
rect 56770 4730 56775 4760
rect 56735 4725 56775 4730
rect 56880 4840 56920 4900
rect 57025 5010 57065 5015
rect 57025 4980 57030 5010
rect 57060 4980 57065 5010
rect 57025 4970 57065 4980
rect 57025 4940 57030 4970
rect 57060 4940 57065 4970
rect 57025 4930 57065 4940
rect 57025 4900 57030 4930
rect 57060 4900 57065 4930
rect 57025 4895 57065 4900
rect 56880 4810 56885 4840
rect 56915 4810 56920 4840
rect 56880 4800 56920 4810
rect 56880 4770 56885 4800
rect 56915 4770 56920 4800
rect 56880 4760 56920 4770
rect 56880 4730 56885 4760
rect 56915 4730 56920 4760
rect 56680 4545 56685 4695
rect 56705 4545 56710 4695
rect 56680 4530 56710 4545
rect 56740 4695 56770 4725
rect 56740 4545 56745 4695
rect 56765 4545 56770 4695
rect 56740 4535 56770 4545
rect 56205 4525 56245 4530
rect 56205 4495 56210 4525
rect 56240 4495 56245 4525
rect 56205 4490 56245 4495
rect 56675 4525 56715 4530
rect 56675 4495 56680 4525
rect 56710 4495 56715 4525
rect 56675 4490 56715 4495
rect 56150 4480 56190 4485
rect 56150 4450 56155 4480
rect 56185 4450 56190 4480
rect 56150 4445 56190 4450
rect 56630 4480 56660 4485
rect 56630 4445 56660 4450
rect 56825 4480 56865 4485
rect 56825 4450 56830 4480
rect 56860 4450 56865 4480
rect 56825 4445 56865 4450
rect 54040 4290 54045 4320
rect 54075 4290 54085 4320
rect 54115 4290 54125 4320
rect 54155 4290 54160 4320
rect 54040 4280 54160 4290
rect 54040 4250 54045 4280
rect 54075 4250 54085 4280
rect 54115 4250 54125 4280
rect 54155 4250 54160 4280
rect 54040 4240 54160 4250
rect 54040 4210 54045 4240
rect 54075 4210 54085 4240
rect 54115 4210 54125 4240
rect 54155 4210 54160 4240
rect 54040 4205 54160 4210
rect 54670 4320 54710 4325
rect 54670 4290 54675 4320
rect 54705 4290 54710 4320
rect 54670 4280 54710 4290
rect 54670 4250 54675 4280
rect 54705 4250 54710 4280
rect 54670 4240 54710 4250
rect 54670 4210 54675 4240
rect 54705 4210 54710 4240
rect 54670 4050 54710 4210
rect 55030 4320 55070 4325
rect 55030 4290 55035 4320
rect 55065 4290 55070 4320
rect 55030 4280 55070 4290
rect 55030 4250 55035 4280
rect 55065 4250 55070 4280
rect 55030 4240 55070 4250
rect 55030 4210 55035 4240
rect 55065 4210 55070 4240
rect 54730 4185 55010 4190
rect 54730 4155 54735 4185
rect 54765 4155 54775 4185
rect 54805 4155 54815 4185
rect 54845 4155 54855 4185
rect 54885 4155 54895 4185
rect 54925 4155 54935 4185
rect 54965 4155 54975 4185
rect 55005 4155 55010 4185
rect 54730 4145 55010 4155
rect 54730 4115 54735 4145
rect 54765 4115 54775 4145
rect 54805 4115 54815 4145
rect 54845 4115 54855 4145
rect 54885 4115 54895 4145
rect 54925 4115 54935 4145
rect 54965 4115 54975 4145
rect 55005 4115 55010 4145
rect 54730 4105 55010 4115
rect 54730 4075 54735 4105
rect 54765 4075 54775 4105
rect 54805 4075 54815 4105
rect 54845 4075 54855 4105
rect 54885 4075 54895 4105
rect 54925 4075 54935 4105
rect 54965 4075 54975 4105
rect 55005 4075 55010 4105
rect 54730 4070 55010 4075
rect 54670 4020 54675 4050
rect 54705 4020 54710 4050
rect 54670 4015 54710 4020
rect 54675 4000 54705 4015
rect 54675 3680 54680 4000
rect 54700 3680 54705 4000
rect 54675 3640 54705 3680
rect 54735 4000 54765 4070
rect 54790 4050 54830 4055
rect 54790 4020 54795 4050
rect 54825 4020 54830 4050
rect 54790 4015 54830 4020
rect 54735 3680 54740 4000
rect 54760 3680 54765 4000
rect 54735 3665 54765 3680
rect 54795 4000 54825 4015
rect 54795 3680 54800 4000
rect 54820 3680 54825 4000
rect 54795 3670 54825 3680
rect 54855 4000 54885 4070
rect 54910 4050 54950 4055
rect 54910 4020 54915 4050
rect 54945 4020 54950 4050
rect 54910 4015 54950 4020
rect 54855 3680 54860 4000
rect 54880 3680 54885 4000
rect 54855 3665 54885 3680
rect 54915 4000 54945 4015
rect 54915 3680 54920 4000
rect 54940 3680 54945 4000
rect 54915 3670 54945 3680
rect 54975 4000 55005 4070
rect 55030 4050 55070 4210
rect 55390 4320 55430 4325
rect 55390 4290 55395 4320
rect 55425 4290 55430 4320
rect 55390 4280 55430 4290
rect 55390 4250 55395 4280
rect 55425 4250 55430 4280
rect 55390 4240 55430 4250
rect 55390 4210 55395 4240
rect 55425 4210 55430 4240
rect 55090 4185 55370 4190
rect 55090 4155 55095 4185
rect 55125 4155 55135 4185
rect 55165 4155 55175 4185
rect 55205 4155 55215 4185
rect 55245 4155 55255 4185
rect 55285 4155 55295 4185
rect 55325 4155 55335 4185
rect 55365 4155 55370 4185
rect 55090 4145 55370 4155
rect 55090 4115 55095 4145
rect 55125 4115 55135 4145
rect 55165 4115 55175 4145
rect 55205 4115 55215 4145
rect 55245 4115 55255 4145
rect 55285 4115 55295 4145
rect 55325 4115 55335 4145
rect 55365 4115 55370 4145
rect 55090 4105 55370 4115
rect 55090 4075 55095 4105
rect 55125 4075 55135 4105
rect 55165 4075 55175 4105
rect 55205 4075 55215 4105
rect 55245 4075 55255 4105
rect 55285 4075 55295 4105
rect 55325 4075 55335 4105
rect 55365 4075 55370 4105
rect 55090 4070 55370 4075
rect 55030 4020 55035 4050
rect 55065 4020 55070 4050
rect 55030 4015 55070 4020
rect 54975 3680 54980 4000
rect 55000 3680 55005 4000
rect 54975 3665 55005 3680
rect 55035 4000 55065 4015
rect 55035 3680 55040 4000
rect 55060 3680 55065 4000
rect 55035 3670 55065 3680
rect 55095 4000 55125 4070
rect 55150 4050 55190 4055
rect 55150 4020 55155 4050
rect 55185 4020 55190 4050
rect 55150 4015 55190 4020
rect 55095 3680 55100 4000
rect 55120 3680 55125 4000
rect 55095 3665 55125 3680
rect 55155 4000 55185 4015
rect 55155 3680 55160 4000
rect 55180 3680 55185 4000
rect 55155 3670 55185 3680
rect 55215 4000 55245 4070
rect 55270 4050 55310 4055
rect 55270 4020 55275 4050
rect 55305 4020 55310 4050
rect 55270 4015 55310 4020
rect 55215 3680 55220 4000
rect 55240 3680 55245 4000
rect 55215 3665 55245 3680
rect 55275 4000 55305 4015
rect 55275 3680 55280 4000
rect 55300 3680 55305 4000
rect 55275 3670 55305 3680
rect 55335 4000 55365 4070
rect 55390 4050 55430 4210
rect 55390 4020 55395 4050
rect 55425 4020 55430 4050
rect 55390 4015 55430 4020
rect 55620 4320 55740 4325
rect 55620 4290 55625 4320
rect 55655 4290 55665 4320
rect 55695 4290 55705 4320
rect 55735 4290 55740 4320
rect 55620 4280 55740 4290
rect 55620 4250 55625 4280
rect 55655 4250 55665 4280
rect 55695 4250 55705 4280
rect 55735 4250 55740 4280
rect 55620 4240 55740 4250
rect 55620 4210 55625 4240
rect 55655 4210 55665 4240
rect 55695 4210 55705 4240
rect 55735 4210 55740 4240
rect 55335 3680 55340 4000
rect 55360 3680 55365 4000
rect 55335 3665 55365 3680
rect 55395 4000 55425 4015
rect 55395 3680 55400 4000
rect 55420 3680 55425 4000
rect 54675 3620 54680 3640
rect 54700 3620 54705 3640
rect 54730 3660 54770 3665
rect 54730 3630 54735 3660
rect 54765 3630 54770 3660
rect 54730 3625 54770 3630
rect 54850 3660 54890 3665
rect 54850 3630 54855 3660
rect 54885 3630 54890 3660
rect 54850 3625 54890 3630
rect 54970 3660 55010 3665
rect 54970 3630 54975 3660
rect 55005 3630 55010 3660
rect 54970 3625 55010 3630
rect 55090 3660 55130 3665
rect 55090 3630 55095 3660
rect 55125 3630 55130 3660
rect 55090 3625 55130 3630
rect 55210 3660 55250 3665
rect 55210 3630 55215 3660
rect 55245 3630 55250 3660
rect 55210 3625 55250 3630
rect 55330 3660 55370 3665
rect 55330 3630 55335 3660
rect 55365 3630 55370 3660
rect 55330 3625 55370 3630
rect 55395 3640 55425 3680
rect 54675 3610 54705 3620
rect 55395 3620 55400 3640
rect 55420 3620 55425 3640
rect 55395 3610 55425 3620
rect 55030 3535 55070 3540
rect 55030 3505 55035 3535
rect 55065 3505 55070 3535
rect 55030 3500 55070 3505
rect 55480 3490 55600 3495
rect 55480 3460 55485 3490
rect 55515 3460 55525 3490
rect 55555 3460 55565 3490
rect 55595 3460 55600 3490
rect 55480 3450 55600 3460
rect 55480 3420 55485 3450
rect 55515 3420 55525 3450
rect 55555 3420 55565 3450
rect 55595 3420 55600 3450
rect 55480 3410 55600 3420
rect 55480 3380 55485 3410
rect 55515 3380 55525 3410
rect 55555 3380 55565 3410
rect 55595 3380 55600 3410
rect 54255 3375 54295 3380
rect 54255 3345 54260 3375
rect 54290 3345 54295 3375
rect 54255 3340 54295 3345
rect 54700 3355 54740 3360
rect 54265 3300 54285 3340
rect 54700 3325 54705 3355
rect 54735 3325 54740 3355
rect 54700 3315 54740 3325
rect 54204 3290 54345 3300
rect 54204 3270 54210 3290
rect 54230 3270 54265 3290
rect 54285 3270 54320 3290
rect 54340 3270 54345 3290
rect 54204 3260 54345 3270
rect 54700 3285 54705 3315
rect 54735 3285 54740 3315
rect 54700 3275 54740 3285
rect 54700 3245 54705 3275
rect 54735 3245 54740 3275
rect 54700 3240 54740 3245
rect 54810 3355 54850 3360
rect 54810 3325 54815 3355
rect 54845 3325 54850 3355
rect 54810 3315 54850 3325
rect 54810 3285 54815 3315
rect 54845 3285 54850 3315
rect 54810 3275 54850 3285
rect 54810 3245 54815 3275
rect 54845 3245 54850 3275
rect 54810 3240 54850 3245
rect 54920 3355 54960 3360
rect 54920 3325 54925 3355
rect 54955 3325 54960 3355
rect 54920 3315 54960 3325
rect 54920 3285 54925 3315
rect 54955 3285 54960 3315
rect 54920 3275 54960 3285
rect 54920 3245 54925 3275
rect 54955 3245 54960 3275
rect 54920 3240 54960 3245
rect 55030 3355 55070 3360
rect 55030 3325 55035 3355
rect 55065 3325 55070 3355
rect 55030 3315 55070 3325
rect 55030 3285 55035 3315
rect 55065 3285 55070 3315
rect 55030 3275 55070 3285
rect 55030 3245 55035 3275
rect 55065 3245 55070 3275
rect 55030 3240 55070 3245
rect 55140 3355 55180 3360
rect 55140 3325 55145 3355
rect 55175 3325 55180 3355
rect 55140 3315 55180 3325
rect 55140 3285 55145 3315
rect 55175 3285 55180 3315
rect 55140 3275 55180 3285
rect 55140 3245 55145 3275
rect 55175 3245 55180 3275
rect 55140 3240 55180 3245
rect 55250 3355 55290 3360
rect 55250 3325 55255 3355
rect 55285 3325 55290 3355
rect 55250 3315 55290 3325
rect 55250 3285 55255 3315
rect 55285 3285 55290 3315
rect 55250 3275 55290 3285
rect 55250 3245 55255 3275
rect 55285 3245 55290 3275
rect 55250 3240 55290 3245
rect 55360 3355 55400 3360
rect 55360 3325 55365 3355
rect 55395 3325 55400 3355
rect 55360 3315 55400 3325
rect 55360 3285 55365 3315
rect 55395 3285 55400 3315
rect 55360 3275 55400 3285
rect 55360 3245 55365 3275
rect 55395 3245 55400 3275
rect 55360 3240 55400 3245
rect 54705 3200 54735 3240
rect 54705 3180 54710 3200
rect 54730 3180 54735 3200
rect 54705 3140 54735 3180
rect 54755 3190 54795 3195
rect 54755 3160 54760 3190
rect 54790 3160 54795 3190
rect 54755 3155 54795 3160
rect 54204 2685 54345 2695
rect 54204 2665 54210 2685
rect 54230 2665 54265 2685
rect 54285 2665 54320 2685
rect 54340 2665 54345 2685
rect 54204 2655 54345 2665
rect 54215 2470 54335 2655
rect 54705 2570 54710 3140
rect 54730 2570 54735 3140
rect 54705 2560 54735 2570
rect 54760 3140 54790 3155
rect 54760 2570 54765 3140
rect 54785 2570 54790 3140
rect 54760 2555 54790 2570
rect 54815 3140 54845 3240
rect 54865 3190 54905 3195
rect 54865 3160 54870 3190
rect 54900 3160 54905 3190
rect 54865 3155 54905 3160
rect 54815 2570 54820 3140
rect 54840 2570 54845 3140
rect 54815 2560 54845 2570
rect 54870 3140 54900 3155
rect 54870 2570 54875 3140
rect 54895 2570 54900 3140
rect 54870 2555 54900 2570
rect 54925 3140 54955 3240
rect 54975 3190 55015 3195
rect 54975 3160 54980 3190
rect 55010 3160 55015 3190
rect 54975 3155 55015 3160
rect 54925 2570 54930 3140
rect 54950 2570 54955 3140
rect 54925 2560 54955 2570
rect 54980 3140 55010 3155
rect 54980 2570 54985 3140
rect 55005 2570 55010 3140
rect 54980 2555 55010 2570
rect 55035 3140 55065 3240
rect 55085 3190 55125 3195
rect 55085 3160 55090 3190
rect 55120 3160 55125 3190
rect 55085 3155 55125 3160
rect 55035 2570 55040 3140
rect 55060 2570 55065 3140
rect 55035 2560 55065 2570
rect 55090 3140 55120 3155
rect 55090 2570 55095 3140
rect 55115 2570 55120 3140
rect 55090 2555 55120 2570
rect 55145 3140 55175 3240
rect 55195 3190 55235 3195
rect 55195 3160 55200 3190
rect 55230 3160 55235 3190
rect 55195 3155 55235 3160
rect 55145 2570 55150 3140
rect 55170 2570 55175 3140
rect 55145 2560 55175 2570
rect 55200 3140 55230 3155
rect 55200 2570 55205 3140
rect 55225 2570 55230 3140
rect 55200 2555 55230 2570
rect 55255 3140 55285 3240
rect 55365 3200 55395 3240
rect 55305 3190 55345 3195
rect 55305 3160 55310 3190
rect 55340 3160 55345 3190
rect 55305 3155 55345 3160
rect 55365 3180 55370 3200
rect 55390 3180 55395 3200
rect 55255 2570 55260 3140
rect 55280 2570 55285 3140
rect 55255 2560 55285 2570
rect 55310 3140 55340 3155
rect 55310 2570 55315 3140
rect 55335 2570 55340 3140
rect 55310 2555 55340 2570
rect 55365 3140 55395 3180
rect 55365 2570 55370 3140
rect 55390 2570 55395 3140
rect 55365 2560 55395 2570
rect 54215 2440 54220 2470
rect 54250 2440 54260 2470
rect 54290 2440 54300 2470
rect 54330 2440 54335 2470
rect 54215 2430 54335 2440
rect 54215 2400 54220 2430
rect 54250 2400 54260 2430
rect 54290 2400 54300 2430
rect 54330 2400 54335 2430
rect 54215 2390 54335 2400
rect 54215 2360 54220 2390
rect 54250 2360 54260 2390
rect 54290 2360 54300 2390
rect 54330 2360 54335 2390
rect 54215 2355 54335 2360
rect 54755 2550 54795 2555
rect 54755 2520 54760 2550
rect 54790 2520 54795 2550
rect 54755 2325 54795 2520
rect 54865 2550 54905 2555
rect 54865 2520 54870 2550
rect 54900 2520 54905 2550
rect 54865 2325 54905 2520
rect 54975 2550 55015 2555
rect 54975 2520 54980 2550
rect 55010 2520 55015 2550
rect 54975 2325 55015 2520
rect 55085 2550 55125 2555
rect 55085 2520 55090 2550
rect 55120 2520 55125 2550
rect 55030 2470 55070 2475
rect 55030 2440 55035 2470
rect 55065 2440 55070 2470
rect 55030 2430 55070 2440
rect 55030 2400 55035 2430
rect 55065 2400 55070 2430
rect 55030 2390 55070 2400
rect 55030 2360 55035 2390
rect 55065 2360 55070 2390
rect 55030 2355 55070 2360
rect 55085 2325 55125 2520
rect 55195 2550 55235 2555
rect 55195 2520 55200 2550
rect 55230 2520 55235 2550
rect 55195 2325 55235 2520
rect 55305 2550 55345 2555
rect 55305 2520 55310 2550
rect 55340 2520 55345 2550
rect 55305 2325 55345 2520
rect 54070 2320 54320 2325
rect 54070 2290 54075 2320
rect 54105 2290 54115 2320
rect 54145 2290 54160 2320
rect 54190 2290 54200 2320
rect 54230 2290 54245 2320
rect 54275 2290 54285 2320
rect 54315 2290 54320 2320
rect 54070 2280 54320 2290
rect 54070 2250 54075 2280
rect 54105 2250 54115 2280
rect 54145 2250 54160 2280
rect 54190 2250 54200 2280
rect 54230 2250 54245 2280
rect 54275 2250 54285 2280
rect 54315 2250 54320 2280
rect 54070 2240 54320 2250
rect 54070 2210 54075 2240
rect 54105 2210 54115 2240
rect 54145 2210 54160 2240
rect 54190 2210 54200 2240
rect 54230 2210 54245 2240
rect 54275 2210 54285 2240
rect 54315 2210 54320 2240
rect 53920 2050 54040 2055
rect 53920 2020 53925 2050
rect 53955 2020 53965 2050
rect 53995 2020 54005 2050
rect 54035 2020 54040 2050
rect 53920 2010 54040 2020
rect 53920 1980 53925 2010
rect 53955 1980 53965 2010
rect 53995 1980 54005 2010
rect 54035 1980 54040 2010
rect 53920 1970 54040 1980
rect 53920 1940 53925 1970
rect 53955 1940 53965 1970
rect 53995 1940 54005 1970
rect 54035 1940 54040 1970
rect 53920 940 54040 1940
rect 53920 910 53925 940
rect 53955 910 53965 940
rect 53995 910 54005 940
rect 54035 910 54040 940
rect 53920 900 54040 910
rect 53920 870 53925 900
rect 53955 870 53965 900
rect 53995 870 54005 900
rect 54035 870 54040 900
rect 53920 860 54040 870
rect 53920 830 53925 860
rect 53955 830 53965 860
rect 53995 830 54005 860
rect 54035 830 54040 860
rect 53920 -575 54040 830
rect 54070 1710 54320 2210
rect 54755 2320 55345 2325
rect 54755 2290 54760 2320
rect 54790 2290 54815 2320
rect 54845 2290 54870 2320
rect 54900 2290 54925 2320
rect 54955 2290 54980 2320
rect 55010 2290 55035 2320
rect 55065 2290 55090 2320
rect 55120 2290 55145 2320
rect 55175 2290 55200 2320
rect 55230 2290 55255 2320
rect 55285 2290 55310 2320
rect 55340 2290 55345 2320
rect 54755 2280 55345 2290
rect 54755 2250 54760 2280
rect 54790 2250 54815 2280
rect 54845 2250 54870 2280
rect 54900 2250 54925 2280
rect 54955 2250 54980 2280
rect 55010 2250 55035 2280
rect 55065 2250 55090 2280
rect 55120 2250 55145 2280
rect 55175 2250 55200 2280
rect 55230 2250 55255 2280
rect 55285 2250 55310 2280
rect 55340 2250 55345 2280
rect 54755 2240 55345 2250
rect 54755 2210 54760 2240
rect 54790 2210 54815 2240
rect 54845 2210 54870 2240
rect 54900 2210 54925 2240
rect 54955 2210 54980 2240
rect 55010 2210 55035 2240
rect 55065 2210 55090 2240
rect 55120 2210 55145 2240
rect 55175 2210 55200 2240
rect 55230 2210 55255 2240
rect 55285 2210 55310 2240
rect 55340 2210 55345 2240
rect 54755 2205 55345 2210
rect 55480 2470 55600 3380
rect 55480 2440 55485 2470
rect 55515 2440 55525 2470
rect 55555 2440 55565 2470
rect 55595 2440 55600 2470
rect 55480 2430 55600 2440
rect 55480 2400 55485 2430
rect 55515 2400 55525 2430
rect 55555 2400 55565 2430
rect 55595 2400 55600 2430
rect 55480 2390 55600 2400
rect 55480 2360 55485 2390
rect 55515 2360 55525 2390
rect 55555 2360 55565 2390
rect 55595 2360 55600 2390
rect 54700 2185 54740 2190
rect 54700 2155 54705 2185
rect 54735 2155 54740 2185
rect 54700 2145 54740 2155
rect 54700 2115 54705 2145
rect 54735 2115 54740 2145
rect 54700 2105 54740 2115
rect 54700 2075 54705 2105
rect 54735 2075 54740 2105
rect 54700 2070 54740 2075
rect 55360 2185 55400 2190
rect 55360 2155 55365 2185
rect 55395 2155 55400 2185
rect 55360 2145 55400 2155
rect 55360 2115 55365 2145
rect 55395 2115 55400 2145
rect 55360 2105 55400 2115
rect 55360 2075 55365 2105
rect 55395 2075 55400 2105
rect 55360 2070 55400 2075
rect 54070 1680 54080 1710
rect 54110 1680 54130 1710
rect 54160 1680 54180 1710
rect 54210 1680 54230 1710
rect 54260 1680 54280 1710
rect 54310 1680 54320 1710
rect 54705 1925 54735 2070
rect 54755 2050 54795 2055
rect 54755 2020 54760 2050
rect 54790 2020 54795 2050
rect 54755 2010 54795 2020
rect 54755 1980 54760 2010
rect 54790 1980 54795 2010
rect 54755 1970 54795 1980
rect 54755 1940 54760 1970
rect 54790 1940 54795 1970
rect 54755 1935 54795 1940
rect 54865 2050 54905 2055
rect 54865 2020 54870 2050
rect 54900 2020 54905 2050
rect 54865 2010 54905 2020
rect 54865 1980 54870 2010
rect 54900 1980 54905 2010
rect 54865 1970 54905 1980
rect 54865 1940 54870 1970
rect 54900 1940 54905 1970
rect 54865 1935 54905 1940
rect 54975 2050 55015 2055
rect 54975 2020 54980 2050
rect 55010 2020 55015 2050
rect 54975 2010 55015 2020
rect 54975 1980 54980 2010
rect 55010 1980 55015 2010
rect 54975 1970 55015 1980
rect 54975 1940 54980 1970
rect 55010 1940 55015 1970
rect 54975 1935 55015 1940
rect 55085 2050 55125 2055
rect 55085 2020 55090 2050
rect 55120 2020 55125 2050
rect 55085 2010 55125 2020
rect 55085 1980 55090 2010
rect 55120 1980 55125 2010
rect 55085 1970 55125 1980
rect 55085 1940 55090 1970
rect 55120 1940 55125 1970
rect 55085 1935 55125 1940
rect 55195 2050 55235 2055
rect 55195 2020 55200 2050
rect 55230 2020 55235 2050
rect 55195 2010 55235 2020
rect 55195 1980 55200 2010
rect 55230 1980 55235 2010
rect 55195 1970 55235 1980
rect 55195 1940 55200 1970
rect 55230 1940 55235 1970
rect 55195 1935 55235 1940
rect 55305 2050 55345 2055
rect 55305 2020 55310 2050
rect 55340 2020 55345 2050
rect 55305 2010 55345 2020
rect 55305 1980 55310 2010
rect 55340 1980 55345 2010
rect 55305 1970 55345 1980
rect 55305 1940 55310 1970
rect 55340 1940 55345 1970
rect 55305 1935 55345 1940
rect 54705 1905 54710 1925
rect 54730 1905 54735 1925
rect 54705 1865 54735 1905
rect 54705 1695 54710 1865
rect 54730 1695 54735 1865
rect 54705 1685 54735 1695
rect 54760 1865 54790 1935
rect 54810 1915 54850 1920
rect 54810 1885 54815 1915
rect 54845 1885 54850 1915
rect 54810 1880 54850 1885
rect 54760 1695 54765 1865
rect 54785 1695 54790 1865
rect 54760 1685 54790 1695
rect 54815 1865 54845 1880
rect 54815 1695 54820 1865
rect 54840 1695 54845 1865
rect 54070 1660 54320 1680
rect 54815 1665 54845 1695
rect 54870 1865 54900 1935
rect 54920 1915 54960 1920
rect 54920 1885 54925 1915
rect 54955 1885 54960 1915
rect 54920 1880 54960 1885
rect 54870 1695 54875 1865
rect 54895 1695 54900 1865
rect 54870 1685 54900 1695
rect 54925 1865 54955 1880
rect 54925 1695 54930 1865
rect 54950 1695 54955 1865
rect 54925 1665 54955 1695
rect 54980 1865 55010 1935
rect 55030 1915 55070 1920
rect 55030 1885 55035 1915
rect 55065 1885 55070 1915
rect 55030 1880 55070 1885
rect 54980 1695 54985 1865
rect 55005 1695 55010 1865
rect 54980 1685 55010 1695
rect 55035 1865 55065 1880
rect 55035 1695 55040 1865
rect 55060 1695 55065 1865
rect 55035 1665 55065 1695
rect 55090 1865 55120 1935
rect 55140 1915 55180 1920
rect 55140 1885 55145 1915
rect 55175 1885 55180 1915
rect 55140 1880 55180 1885
rect 55090 1695 55095 1865
rect 55115 1695 55120 1865
rect 55090 1685 55120 1695
rect 55145 1865 55175 1880
rect 55145 1695 55150 1865
rect 55170 1695 55175 1865
rect 55145 1665 55175 1695
rect 55200 1865 55230 1935
rect 55250 1915 55290 1920
rect 55250 1885 55255 1915
rect 55285 1885 55290 1915
rect 55250 1880 55290 1885
rect 55200 1695 55205 1865
rect 55225 1695 55230 1865
rect 55200 1685 55230 1695
rect 55255 1865 55285 1880
rect 55255 1695 55260 1865
rect 55280 1695 55285 1865
rect 55255 1665 55285 1695
rect 55310 1865 55340 1935
rect 55310 1695 55315 1865
rect 55335 1695 55340 1865
rect 55310 1685 55340 1695
rect 55365 1925 55395 2070
rect 55365 1905 55370 1925
rect 55390 1905 55395 1925
rect 55365 1865 55395 1905
rect 55365 1695 55370 1865
rect 55390 1695 55395 1865
rect 55365 1685 55395 1695
rect 54070 1630 54080 1660
rect 54110 1630 54130 1660
rect 54160 1630 54180 1660
rect 54210 1630 54230 1660
rect 54260 1630 54280 1660
rect 54310 1630 54320 1660
rect 54070 1610 54320 1630
rect 54565 1660 54605 1665
rect 54565 1630 54570 1660
rect 54600 1630 54605 1660
rect 54565 1625 54605 1630
rect 54810 1660 54850 1665
rect 54810 1630 54815 1660
rect 54845 1630 54850 1660
rect 54810 1625 54850 1630
rect 54920 1660 54960 1665
rect 54920 1630 54925 1660
rect 54955 1630 54960 1660
rect 54920 1625 54960 1630
rect 55030 1660 55070 1665
rect 55030 1630 55035 1660
rect 55065 1630 55070 1660
rect 55030 1625 55070 1630
rect 55140 1660 55180 1665
rect 55140 1630 55145 1660
rect 55175 1630 55180 1660
rect 55140 1625 55180 1630
rect 55250 1660 55290 1665
rect 55250 1630 55255 1660
rect 55285 1630 55290 1660
rect 55250 1625 55290 1630
rect 54070 1580 54080 1610
rect 54110 1580 54130 1610
rect 54160 1580 54180 1610
rect 54210 1580 54230 1610
rect 54260 1580 54280 1610
rect 54310 1580 54320 1610
rect 54070 310 54320 1580
rect 54335 1160 54370 1166
rect 54335 1120 54370 1125
rect 54395 1160 54430 1165
rect 54395 1120 54430 1125
rect 54455 1160 54490 1165
rect 54455 1120 54490 1125
rect 54515 1160 54550 1165
rect 54515 1120 54550 1125
rect 54345 810 54365 1120
rect 54465 1090 54485 1120
rect 54575 1090 54595 1625
rect 55195 1595 55235 1600
rect 55195 1565 55200 1595
rect 55230 1565 55235 1595
rect 55195 1555 55235 1565
rect 55195 1525 55200 1555
rect 55230 1525 55235 1555
rect 55195 1520 55235 1525
rect 55480 1595 55600 2360
rect 55480 1565 55485 1595
rect 55515 1565 55525 1595
rect 55555 1565 55565 1595
rect 55595 1565 55600 1595
rect 55480 1555 55600 1565
rect 55480 1525 55485 1555
rect 55515 1525 55525 1555
rect 55555 1525 55565 1555
rect 55595 1525 55600 1555
rect 55480 1520 55600 1525
rect 55620 3355 55740 4210
rect 56005 4185 56765 4190
rect 56005 4155 56010 4185
rect 56040 4155 56050 4185
rect 56080 4155 56090 4185
rect 56120 4155 56130 4185
rect 56160 4155 56170 4185
rect 56200 4155 56210 4185
rect 56240 4155 56250 4185
rect 56280 4155 56290 4185
rect 56320 4155 56330 4185
rect 56360 4155 56370 4185
rect 56400 4155 56410 4185
rect 56440 4155 56450 4185
rect 56480 4155 56490 4185
rect 56520 4155 56530 4185
rect 56560 4155 56570 4185
rect 56600 4155 56610 4185
rect 56640 4155 56650 4185
rect 56680 4155 56690 4185
rect 56720 4155 56730 4185
rect 56760 4155 56765 4185
rect 56005 4145 56765 4155
rect 56005 4115 56010 4145
rect 56040 4115 56050 4145
rect 56080 4115 56090 4145
rect 56120 4115 56130 4145
rect 56160 4115 56170 4145
rect 56200 4115 56210 4145
rect 56240 4115 56250 4145
rect 56280 4115 56290 4145
rect 56320 4115 56330 4145
rect 56360 4115 56370 4145
rect 56400 4115 56410 4145
rect 56440 4115 56450 4145
rect 56480 4115 56490 4145
rect 56520 4115 56530 4145
rect 56560 4115 56570 4145
rect 56600 4115 56610 4145
rect 56640 4115 56650 4145
rect 56680 4115 56690 4145
rect 56720 4115 56730 4145
rect 56760 4115 56765 4145
rect 56005 4105 56765 4115
rect 56005 4075 56010 4105
rect 56040 4075 56050 4105
rect 56080 4075 56090 4105
rect 56120 4075 56130 4105
rect 56160 4075 56170 4105
rect 56200 4075 56210 4105
rect 56240 4075 56250 4105
rect 56280 4075 56290 4105
rect 56320 4075 56330 4105
rect 56360 4075 56370 4105
rect 56400 4075 56410 4105
rect 56440 4075 56450 4105
rect 56480 4075 56490 4105
rect 56520 4075 56530 4105
rect 56560 4075 56570 4105
rect 56600 4075 56610 4105
rect 56640 4075 56650 4105
rect 56680 4075 56690 4105
rect 56720 4075 56730 4105
rect 56760 4075 56765 4105
rect 56005 4070 56765 4075
rect 56010 4000 56040 4070
rect 56065 4050 56105 4055
rect 56065 4020 56070 4050
rect 56100 4020 56105 4050
rect 56065 4015 56105 4020
rect 56010 3680 56015 4000
rect 56035 3680 56040 4000
rect 56010 3640 56040 3680
rect 56070 4000 56100 4015
rect 56070 3680 56075 4000
rect 56095 3680 56100 4000
rect 56070 3665 56100 3680
rect 56130 4000 56160 4070
rect 56185 4050 56225 4055
rect 56185 4020 56190 4050
rect 56220 4020 56225 4050
rect 56185 4015 56225 4020
rect 56130 3680 56135 4000
rect 56155 3680 56160 4000
rect 56130 3670 56160 3680
rect 56190 4000 56220 4015
rect 56190 3680 56195 4000
rect 56215 3680 56220 4000
rect 56190 3665 56220 3680
rect 56250 4000 56280 4070
rect 56305 4050 56345 4055
rect 56305 4020 56310 4050
rect 56340 4020 56345 4050
rect 56305 4015 56345 4020
rect 56250 3680 56255 4000
rect 56275 3680 56280 4000
rect 56250 3670 56280 3680
rect 56310 4000 56340 4015
rect 56310 3680 56315 4000
rect 56335 3680 56340 4000
rect 56310 3665 56340 3680
rect 56370 4000 56400 4070
rect 56425 4050 56465 4055
rect 56425 4020 56430 4050
rect 56460 4020 56465 4050
rect 56425 4015 56465 4020
rect 56370 3680 56375 4000
rect 56395 3680 56400 4000
rect 56370 3670 56400 3680
rect 56430 4000 56460 4015
rect 56430 3680 56435 4000
rect 56455 3680 56460 4000
rect 56430 3665 56460 3680
rect 56490 4000 56520 4070
rect 56545 4050 56585 4055
rect 56545 4020 56550 4050
rect 56580 4020 56585 4050
rect 56545 4015 56585 4020
rect 56490 3680 56495 4000
rect 56515 3680 56520 4000
rect 56490 3670 56520 3680
rect 56550 4000 56580 4015
rect 56550 3680 56555 4000
rect 56575 3680 56580 4000
rect 56550 3665 56580 3680
rect 56610 4000 56640 4070
rect 56665 4050 56705 4055
rect 56665 4020 56670 4050
rect 56700 4020 56705 4050
rect 56665 4015 56705 4020
rect 56610 3680 56615 4000
rect 56635 3680 56640 4000
rect 56610 3670 56640 3680
rect 56670 4000 56700 4015
rect 56670 3680 56675 4000
rect 56695 3680 56700 4000
rect 56670 3665 56700 3680
rect 56730 4000 56760 4070
rect 56730 3680 56735 4000
rect 56755 3680 56760 4000
rect 56010 3620 56015 3640
rect 56035 3620 56040 3640
rect 56010 3610 56040 3620
rect 56065 3660 56105 3665
rect 56065 3630 56070 3660
rect 56100 3630 56105 3660
rect 56065 3495 56105 3630
rect 56185 3660 56225 3665
rect 56185 3630 56190 3660
rect 56220 3630 56225 3660
rect 56185 3495 56225 3630
rect 56305 3660 56345 3665
rect 56305 3630 56310 3660
rect 56340 3630 56345 3660
rect 56305 3495 56345 3630
rect 56425 3660 56465 3665
rect 56425 3630 56430 3660
rect 56460 3630 56465 3660
rect 56365 3580 56405 3585
rect 56365 3550 56370 3580
rect 56400 3550 56405 3580
rect 56365 3545 56405 3550
rect 56425 3495 56465 3630
rect 56545 3660 56585 3665
rect 56545 3630 56550 3660
rect 56580 3630 56585 3660
rect 56545 3495 56585 3630
rect 56665 3660 56705 3665
rect 56665 3630 56670 3660
rect 56700 3630 56705 3660
rect 56665 3495 56705 3630
rect 56730 3640 56760 3680
rect 56730 3620 56735 3640
rect 56755 3620 56760 3640
rect 56730 3610 56760 3620
rect 56845 3585 56865 4445
rect 56880 4320 56920 4730
rect 57030 4865 57060 4895
rect 57030 4545 57035 4865
rect 57055 4545 57060 4865
rect 57030 4535 57060 4545
rect 57090 4865 57120 5030
rect 57145 5010 57185 5015
rect 57145 4980 57150 5010
rect 57180 4980 57185 5010
rect 57145 4970 57185 4980
rect 57145 4940 57150 4970
rect 57180 4940 57185 4970
rect 57145 4930 57185 4940
rect 57145 4900 57150 4930
rect 57180 4900 57185 4930
rect 57145 4895 57185 4900
rect 57205 5010 57245 5015
rect 57205 4980 57210 5010
rect 57240 4980 57245 5010
rect 57205 4970 57245 4980
rect 57205 4940 57210 4970
rect 57240 4940 57245 4970
rect 57205 4930 57245 4940
rect 57205 4900 57210 4930
rect 57240 4900 57245 4930
rect 57205 4895 57245 4900
rect 57495 4930 57535 4935
rect 57495 4900 57500 4930
rect 57530 4900 57535 4930
rect 57495 4895 57535 4900
rect 57555 4930 57595 5035
rect 57555 4900 57560 4930
rect 57590 4900 57595 4930
rect 57555 4895 57595 4900
rect 57675 4930 57715 4935
rect 57675 4900 57680 4930
rect 57710 4900 57715 4930
rect 57675 4895 57715 4900
rect 57090 4545 57095 4865
rect 57115 4545 57120 4865
rect 57090 4530 57120 4545
rect 57150 4865 57180 4895
rect 57150 4545 57155 4865
rect 57175 4545 57180 4865
rect 57150 4535 57180 4545
rect 57210 4865 57240 4895
rect 57210 4545 57215 4865
rect 57235 4545 57240 4865
rect 57210 4535 57240 4545
rect 57500 4865 57530 4895
rect 57500 4545 57505 4865
rect 57525 4545 57530 4865
rect 57500 4535 57530 4545
rect 57560 4865 57590 4895
rect 57560 4545 57565 4865
rect 57585 4545 57590 4865
rect 57560 4530 57590 4545
rect 57620 4865 57650 4875
rect 57620 4545 57625 4865
rect 57645 4545 57650 4865
rect 57085 4525 57125 4530
rect 57085 4495 57090 4525
rect 57120 4495 57125 4525
rect 57085 4490 57125 4495
rect 57555 4525 57595 4530
rect 57555 4495 57560 4525
rect 57590 4495 57595 4525
rect 57555 4490 57595 4495
rect 57140 4475 57170 4485
rect 57140 4455 57145 4475
rect 57165 4455 57170 4475
rect 56880 4290 56885 4320
rect 56915 4290 56920 4320
rect 56880 4280 56920 4290
rect 56880 4250 56885 4280
rect 56915 4250 56920 4280
rect 56880 4240 56920 4250
rect 56880 4210 56885 4240
rect 56915 4210 56920 4240
rect 56880 4205 56920 4210
rect 56935 4425 56975 4430
rect 56935 4395 56940 4425
rect 56970 4395 56975 4425
rect 57140 4420 57170 4455
rect 57576 4470 57606 4475
rect 57576 4435 57606 4440
rect 57620 4420 57650 4545
rect 57680 4865 57710 4895
rect 57680 4545 57685 4865
rect 57705 4545 57710 4865
rect 57680 4535 57710 4545
rect 56935 4390 56975 4395
rect 57135 4415 57175 4420
rect 56835 3580 56875 3585
rect 56835 3550 56840 3580
rect 56870 3550 56875 3580
rect 56835 3545 56875 3550
rect 56935 3540 56955 4390
rect 57135 4385 57140 4415
rect 57170 4385 57175 4415
rect 57135 4380 57175 4385
rect 57615 4415 57655 4420
rect 57615 4385 57620 4415
rect 57650 4385 57655 4415
rect 57615 4380 57655 4385
rect 58055 4320 58175 4325
rect 58055 4290 58060 4320
rect 58090 4290 58100 4320
rect 58130 4290 58140 4320
rect 58170 4290 58175 4320
rect 58055 4280 58175 4290
rect 58055 4250 58060 4280
rect 58090 4250 58100 4280
rect 58130 4250 58140 4280
rect 58170 4250 58175 4280
rect 58055 4240 58175 4250
rect 58055 4210 58060 4240
rect 58090 4210 58100 4240
rect 58130 4210 58140 4240
rect 58170 4210 58175 4240
rect 57035 4185 57795 4190
rect 57035 4155 57040 4185
rect 57070 4155 57080 4185
rect 57110 4155 57120 4185
rect 57150 4155 57160 4185
rect 57190 4155 57200 4185
rect 57230 4155 57240 4185
rect 57270 4155 57280 4185
rect 57310 4155 57320 4185
rect 57350 4155 57360 4185
rect 57390 4155 57400 4185
rect 57430 4155 57440 4185
rect 57470 4155 57480 4185
rect 57510 4155 57520 4185
rect 57550 4155 57560 4185
rect 57590 4155 57600 4185
rect 57630 4155 57640 4185
rect 57670 4155 57680 4185
rect 57710 4155 57720 4185
rect 57750 4155 57760 4185
rect 57790 4155 57795 4185
rect 57035 4145 57795 4155
rect 57035 4115 57040 4145
rect 57070 4115 57080 4145
rect 57110 4115 57120 4145
rect 57150 4115 57160 4145
rect 57190 4115 57200 4145
rect 57230 4115 57240 4145
rect 57270 4115 57280 4145
rect 57310 4115 57320 4145
rect 57350 4115 57360 4145
rect 57390 4115 57400 4145
rect 57430 4115 57440 4145
rect 57470 4115 57480 4145
rect 57510 4115 57520 4145
rect 57550 4115 57560 4145
rect 57590 4115 57600 4145
rect 57630 4115 57640 4145
rect 57670 4115 57680 4145
rect 57710 4115 57720 4145
rect 57750 4115 57760 4145
rect 57790 4115 57795 4145
rect 57035 4105 57795 4115
rect 57035 4075 57040 4105
rect 57070 4075 57080 4105
rect 57110 4075 57120 4105
rect 57150 4075 57160 4105
rect 57190 4075 57200 4105
rect 57230 4075 57240 4105
rect 57270 4075 57280 4105
rect 57310 4075 57320 4105
rect 57350 4075 57360 4105
rect 57390 4075 57400 4105
rect 57430 4075 57440 4105
rect 57470 4075 57480 4105
rect 57510 4075 57520 4105
rect 57550 4075 57560 4105
rect 57590 4075 57600 4105
rect 57630 4075 57640 4105
rect 57670 4075 57680 4105
rect 57710 4075 57720 4105
rect 57750 4075 57760 4105
rect 57790 4075 57795 4105
rect 57035 4070 57795 4075
rect 57040 4000 57070 4070
rect 57095 4050 57135 4055
rect 57095 4020 57100 4050
rect 57130 4020 57135 4050
rect 57095 4015 57135 4020
rect 57040 3680 57045 4000
rect 57065 3680 57070 4000
rect 57040 3640 57070 3680
rect 57100 4000 57130 4015
rect 57100 3680 57105 4000
rect 57125 3680 57130 4000
rect 57100 3665 57130 3680
rect 57160 4000 57190 4070
rect 57215 4050 57255 4055
rect 57215 4020 57220 4050
rect 57250 4020 57255 4050
rect 57215 4015 57255 4020
rect 57160 3680 57165 4000
rect 57185 3680 57190 4000
rect 57160 3670 57190 3680
rect 57220 4000 57250 4015
rect 57220 3680 57225 4000
rect 57245 3680 57250 4000
rect 57220 3665 57250 3680
rect 57280 4000 57310 4070
rect 57335 4050 57375 4055
rect 57335 4020 57340 4050
rect 57370 4020 57375 4050
rect 57335 4015 57375 4020
rect 57280 3680 57285 4000
rect 57305 3680 57310 4000
rect 57280 3670 57310 3680
rect 57340 4000 57370 4015
rect 57340 3680 57345 4000
rect 57365 3680 57370 4000
rect 57340 3665 57370 3680
rect 57400 4000 57430 4070
rect 57455 4050 57495 4055
rect 57455 4020 57460 4050
rect 57490 4020 57495 4050
rect 57455 4015 57495 4020
rect 57400 3680 57405 4000
rect 57425 3680 57430 4000
rect 57400 3670 57430 3680
rect 57460 4000 57490 4015
rect 57460 3680 57465 4000
rect 57485 3680 57490 4000
rect 57460 3665 57490 3680
rect 57520 4000 57550 4070
rect 57575 4050 57615 4055
rect 57575 4020 57580 4050
rect 57610 4020 57615 4050
rect 57575 4015 57615 4020
rect 57520 3680 57525 4000
rect 57545 3680 57550 4000
rect 57520 3670 57550 3680
rect 57580 4000 57610 4015
rect 57580 3680 57585 4000
rect 57605 3680 57610 4000
rect 57580 3665 57610 3680
rect 57640 4000 57670 4070
rect 57695 4050 57735 4055
rect 57695 4020 57700 4050
rect 57730 4020 57735 4050
rect 57695 4015 57735 4020
rect 57640 3680 57645 4000
rect 57665 3680 57670 4000
rect 57640 3670 57670 3680
rect 57700 4000 57730 4015
rect 57700 3680 57705 4000
rect 57725 3680 57730 4000
rect 57700 3665 57730 3680
rect 57760 4000 57790 4070
rect 57760 3680 57765 4000
rect 57785 3680 57790 4000
rect 57040 3620 57045 3640
rect 57065 3620 57070 3640
rect 57040 3610 57070 3620
rect 57095 3660 57135 3665
rect 57095 3630 57100 3660
rect 57130 3630 57135 3660
rect 56925 3535 56965 3540
rect 56925 3505 56930 3535
rect 56960 3505 56965 3535
rect 56925 3500 56965 3505
rect 56065 3490 56705 3495
rect 56065 3460 56070 3490
rect 56100 3460 56110 3490
rect 56140 3460 56150 3490
rect 56180 3460 56190 3490
rect 56220 3460 56230 3490
rect 56260 3460 56270 3490
rect 56300 3460 56310 3490
rect 56340 3460 56350 3490
rect 56380 3460 56390 3490
rect 56420 3460 56430 3490
rect 56460 3460 56470 3490
rect 56500 3460 56510 3490
rect 56540 3460 56550 3490
rect 56580 3460 56590 3490
rect 56620 3460 56630 3490
rect 56660 3460 56670 3490
rect 56700 3460 56705 3490
rect 56065 3450 56705 3460
rect 56065 3420 56070 3450
rect 56100 3420 56110 3450
rect 56140 3420 56150 3450
rect 56180 3420 56190 3450
rect 56220 3420 56230 3450
rect 56260 3420 56270 3450
rect 56300 3420 56310 3450
rect 56340 3420 56350 3450
rect 56380 3420 56390 3450
rect 56420 3420 56430 3450
rect 56460 3420 56470 3450
rect 56500 3420 56510 3450
rect 56540 3420 56550 3450
rect 56580 3420 56590 3450
rect 56620 3420 56630 3450
rect 56660 3420 56670 3450
rect 56700 3420 56705 3450
rect 56065 3410 56705 3420
rect 56065 3380 56070 3410
rect 56100 3380 56110 3410
rect 56140 3380 56150 3410
rect 56180 3380 56190 3410
rect 56220 3380 56230 3410
rect 56260 3380 56270 3410
rect 56300 3380 56310 3410
rect 56340 3380 56350 3410
rect 56380 3380 56390 3410
rect 56420 3380 56430 3410
rect 56460 3380 56470 3410
rect 56500 3380 56510 3410
rect 56540 3380 56550 3410
rect 56580 3380 56590 3410
rect 56620 3380 56630 3410
rect 56660 3380 56670 3410
rect 56700 3380 56705 3410
rect 56065 3375 56705 3380
rect 57095 3495 57135 3630
rect 57215 3660 57255 3665
rect 57215 3630 57220 3660
rect 57250 3630 57255 3660
rect 57215 3495 57255 3630
rect 57335 3660 57375 3665
rect 57335 3630 57340 3660
rect 57370 3630 57375 3660
rect 57335 3495 57375 3630
rect 57455 3660 57495 3665
rect 57455 3630 57460 3660
rect 57490 3630 57495 3660
rect 57395 3580 57435 3585
rect 57395 3550 57400 3580
rect 57430 3550 57435 3580
rect 57395 3545 57435 3550
rect 57455 3495 57495 3630
rect 57575 3660 57615 3665
rect 57575 3630 57580 3660
rect 57610 3630 57615 3660
rect 57575 3495 57615 3630
rect 57695 3660 57735 3665
rect 57695 3630 57700 3660
rect 57730 3630 57735 3660
rect 57695 3495 57735 3630
rect 57760 3640 57790 3680
rect 57760 3620 57765 3640
rect 57785 3620 57790 3640
rect 57760 3610 57790 3620
rect 57095 3490 57735 3495
rect 57095 3460 57100 3490
rect 57130 3460 57140 3490
rect 57170 3460 57180 3490
rect 57210 3460 57220 3490
rect 57250 3460 57260 3490
rect 57290 3460 57300 3490
rect 57330 3460 57340 3490
rect 57370 3460 57380 3490
rect 57410 3460 57420 3490
rect 57450 3460 57460 3490
rect 57490 3460 57500 3490
rect 57530 3460 57540 3490
rect 57570 3460 57580 3490
rect 57610 3460 57620 3490
rect 57650 3460 57660 3490
rect 57690 3460 57700 3490
rect 57730 3460 57735 3490
rect 57095 3450 57735 3460
rect 57095 3420 57100 3450
rect 57130 3420 57140 3450
rect 57170 3420 57180 3450
rect 57210 3420 57220 3450
rect 57250 3420 57260 3450
rect 57290 3420 57300 3450
rect 57330 3420 57340 3450
rect 57370 3420 57380 3450
rect 57410 3420 57420 3450
rect 57450 3420 57460 3450
rect 57490 3420 57500 3450
rect 57530 3420 57540 3450
rect 57570 3420 57580 3450
rect 57610 3420 57620 3450
rect 57650 3420 57660 3450
rect 57690 3420 57700 3450
rect 57730 3420 57735 3450
rect 57095 3410 57735 3420
rect 57095 3380 57100 3410
rect 57130 3380 57140 3410
rect 57170 3380 57180 3410
rect 57210 3380 57220 3410
rect 57250 3380 57260 3410
rect 57290 3380 57300 3410
rect 57330 3380 57340 3410
rect 57370 3380 57380 3410
rect 57410 3380 57420 3410
rect 57450 3380 57460 3410
rect 57490 3380 57500 3410
rect 57530 3380 57540 3410
rect 57570 3380 57580 3410
rect 57610 3380 57620 3410
rect 57650 3380 57660 3410
rect 57690 3380 57700 3410
rect 57730 3380 57735 3410
rect 57095 3375 57735 3380
rect 55620 3325 55625 3355
rect 55655 3325 55665 3355
rect 55695 3325 55705 3355
rect 55735 3325 55740 3355
rect 58055 3355 58175 4210
rect 58370 4320 58410 4325
rect 58370 4290 58375 4320
rect 58405 4290 58410 4320
rect 58370 4280 58410 4290
rect 58370 4250 58375 4280
rect 58405 4250 58410 4280
rect 58370 4240 58410 4250
rect 58370 4210 58375 4240
rect 58405 4210 58410 4240
rect 58370 4050 58410 4210
rect 58730 4320 58770 4325
rect 58730 4290 58735 4320
rect 58765 4290 58770 4320
rect 58730 4280 58770 4290
rect 58730 4250 58735 4280
rect 58765 4250 58770 4280
rect 58730 4240 58770 4250
rect 58730 4210 58735 4240
rect 58765 4210 58770 4240
rect 58430 4185 58710 4190
rect 58430 4155 58435 4185
rect 58465 4155 58475 4185
rect 58505 4155 58515 4185
rect 58545 4155 58555 4185
rect 58585 4155 58595 4185
rect 58625 4155 58635 4185
rect 58665 4155 58675 4185
rect 58705 4155 58710 4185
rect 58430 4145 58710 4155
rect 58430 4115 58435 4145
rect 58465 4115 58475 4145
rect 58505 4115 58515 4145
rect 58545 4115 58555 4145
rect 58585 4115 58595 4145
rect 58625 4115 58635 4145
rect 58665 4115 58675 4145
rect 58705 4115 58710 4145
rect 58430 4105 58710 4115
rect 58430 4075 58435 4105
rect 58465 4075 58475 4105
rect 58505 4075 58515 4105
rect 58545 4075 58555 4105
rect 58585 4075 58595 4105
rect 58625 4075 58635 4105
rect 58665 4075 58675 4105
rect 58705 4075 58710 4105
rect 58430 4070 58710 4075
rect 58370 4020 58375 4050
rect 58405 4020 58410 4050
rect 58370 4015 58410 4020
rect 58375 4000 58405 4015
rect 58375 3680 58380 4000
rect 58400 3680 58405 4000
rect 58375 3640 58405 3680
rect 58435 4000 58465 4070
rect 58490 4050 58530 4055
rect 58490 4020 58495 4050
rect 58525 4020 58530 4050
rect 58490 4015 58530 4020
rect 58435 3680 58440 4000
rect 58460 3680 58465 4000
rect 58435 3665 58465 3680
rect 58495 4000 58525 4015
rect 58495 3680 58500 4000
rect 58520 3680 58525 4000
rect 58495 3670 58525 3680
rect 58555 4000 58585 4070
rect 58610 4050 58650 4055
rect 58610 4020 58615 4050
rect 58645 4020 58650 4050
rect 58610 4015 58650 4020
rect 58555 3680 58560 4000
rect 58580 3680 58585 4000
rect 58555 3665 58585 3680
rect 58615 4000 58645 4015
rect 58615 3680 58620 4000
rect 58640 3680 58645 4000
rect 58615 3670 58645 3680
rect 58675 4000 58705 4070
rect 58730 4050 58770 4210
rect 59090 4320 59130 4325
rect 59090 4290 59095 4320
rect 59125 4290 59130 4320
rect 59090 4280 59130 4290
rect 59090 4250 59095 4280
rect 59125 4250 59130 4280
rect 59090 4240 59130 4250
rect 59090 4210 59095 4240
rect 59125 4210 59130 4240
rect 58790 4185 59070 4190
rect 58790 4155 58795 4185
rect 58825 4155 58835 4185
rect 58865 4155 58875 4185
rect 58905 4155 58915 4185
rect 58945 4155 58955 4185
rect 58985 4155 58995 4185
rect 59025 4155 59035 4185
rect 59065 4155 59070 4185
rect 58790 4145 59070 4155
rect 58790 4115 58795 4145
rect 58825 4115 58835 4145
rect 58865 4115 58875 4145
rect 58905 4115 58915 4145
rect 58945 4115 58955 4145
rect 58985 4115 58995 4145
rect 59025 4115 59035 4145
rect 59065 4115 59070 4145
rect 58790 4105 59070 4115
rect 58790 4075 58795 4105
rect 58825 4075 58835 4105
rect 58865 4075 58875 4105
rect 58905 4075 58915 4105
rect 58945 4075 58955 4105
rect 58985 4075 58995 4105
rect 59025 4075 59035 4105
rect 59065 4075 59070 4105
rect 58790 4070 59070 4075
rect 58730 4020 58735 4050
rect 58765 4020 58770 4050
rect 58730 4015 58770 4020
rect 58675 3680 58680 4000
rect 58700 3680 58705 4000
rect 58675 3665 58705 3680
rect 58735 4000 58765 4015
rect 58735 3680 58740 4000
rect 58760 3680 58765 4000
rect 58735 3670 58765 3680
rect 58795 4000 58825 4070
rect 58850 4050 58890 4055
rect 58850 4020 58855 4050
rect 58885 4020 58890 4050
rect 58850 4015 58890 4020
rect 58795 3680 58800 4000
rect 58820 3680 58825 4000
rect 58795 3665 58825 3680
rect 58855 4000 58885 4015
rect 58855 3680 58860 4000
rect 58880 3680 58885 4000
rect 58855 3670 58885 3680
rect 58915 4000 58945 4070
rect 58970 4050 59010 4055
rect 58970 4020 58975 4050
rect 59005 4020 59010 4050
rect 58970 4015 59010 4020
rect 58915 3680 58920 4000
rect 58940 3680 58945 4000
rect 58915 3665 58945 3680
rect 58975 4000 59005 4015
rect 58975 3680 58980 4000
rect 59000 3680 59005 4000
rect 58975 3670 59005 3680
rect 59035 4000 59065 4070
rect 59090 4050 59130 4210
rect 59640 4320 59760 6110
rect 59640 4290 59645 4320
rect 59675 4290 59685 4320
rect 59715 4290 59725 4320
rect 59755 4290 59760 4320
rect 59640 4280 59760 4290
rect 59640 4250 59645 4280
rect 59675 4250 59685 4280
rect 59715 4250 59725 4280
rect 59755 4250 59760 4280
rect 59640 4240 59760 4250
rect 59640 4210 59645 4240
rect 59675 4210 59685 4240
rect 59715 4210 59725 4240
rect 59755 4210 59760 4240
rect 59640 4195 59760 4210
rect 59990 4320 60110 6110
rect 59990 4290 59995 4320
rect 60025 4290 60035 4320
rect 60065 4290 60075 4320
rect 60105 4290 60110 4320
rect 59990 4280 60110 4290
rect 59990 4250 59995 4280
rect 60025 4250 60035 4280
rect 60065 4250 60075 4280
rect 60105 4250 60110 4280
rect 59990 4240 60110 4250
rect 59990 4210 59995 4240
rect 60025 4210 60035 4240
rect 60065 4210 60075 4240
rect 60105 4210 60110 4240
rect 59990 4205 60110 4210
rect 60690 4320 60810 6110
rect 60690 4290 60695 4320
rect 60725 4290 60735 4320
rect 60765 4290 60775 4320
rect 60805 4290 60810 4320
rect 60690 4280 60810 4290
rect 60690 4250 60695 4280
rect 60725 4250 60735 4280
rect 60765 4250 60775 4280
rect 60805 4250 60810 4280
rect 60690 4240 60810 4250
rect 60690 4210 60695 4240
rect 60725 4210 60735 4240
rect 60765 4210 60775 4240
rect 60805 4210 60810 4240
rect 60690 4205 60810 4210
rect 61040 4320 61160 6110
rect 61040 4290 61045 4320
rect 61075 4290 61085 4320
rect 61115 4290 61125 4320
rect 61155 4290 61160 4320
rect 61040 4280 61160 4290
rect 61040 4250 61045 4280
rect 61075 4250 61085 4280
rect 61115 4250 61125 4280
rect 61155 4250 61160 4280
rect 61040 4240 61160 4250
rect 61040 4210 61045 4240
rect 61075 4210 61085 4240
rect 61115 4210 61125 4240
rect 61155 4210 61160 4240
rect 61040 4205 61160 4210
rect 61390 4320 61510 6110
rect 61390 4290 61395 4320
rect 61425 4290 61435 4320
rect 61465 4290 61475 4320
rect 61505 4290 61510 4320
rect 61390 4280 61510 4290
rect 61390 4250 61395 4280
rect 61425 4250 61435 4280
rect 61465 4250 61475 4280
rect 61505 4250 61510 4280
rect 61390 4240 61510 4250
rect 61390 4210 61395 4240
rect 61425 4210 61435 4240
rect 61465 4210 61475 4240
rect 61505 4210 61510 4240
rect 61390 4205 61510 4210
rect 59090 4020 59095 4050
rect 59125 4020 59130 4050
rect 59090 4015 59130 4020
rect 59035 3680 59040 4000
rect 59060 3680 59065 4000
rect 59035 3665 59065 3680
rect 59095 4000 59125 4015
rect 59095 3680 59100 4000
rect 59120 3680 59125 4000
rect 58375 3620 58380 3640
rect 58400 3620 58405 3640
rect 58430 3660 58470 3665
rect 58430 3630 58435 3660
rect 58465 3630 58470 3660
rect 58430 3625 58470 3630
rect 58550 3660 58590 3665
rect 58550 3630 58555 3660
rect 58585 3630 58590 3660
rect 58550 3625 58590 3630
rect 58670 3660 58710 3665
rect 58670 3630 58675 3660
rect 58705 3630 58710 3660
rect 58670 3625 58710 3630
rect 58790 3660 58830 3665
rect 58790 3630 58795 3660
rect 58825 3630 58830 3660
rect 58790 3625 58830 3630
rect 58910 3660 58950 3665
rect 58910 3630 58915 3660
rect 58945 3630 58950 3660
rect 58910 3625 58950 3630
rect 59030 3660 59070 3665
rect 59030 3630 59035 3660
rect 59065 3630 59070 3660
rect 59030 3625 59070 3630
rect 59095 3640 59125 3680
rect 58375 3610 58405 3620
rect 59095 3620 59100 3640
rect 59120 3620 59125 3640
rect 59095 3610 59125 3620
rect 58730 3535 58770 3540
rect 58730 3505 58735 3535
rect 58765 3505 58770 3535
rect 58730 3500 58770 3505
rect 55620 3315 55740 3325
rect 55620 3285 55625 3315
rect 55655 3285 55665 3315
rect 55695 3285 55705 3315
rect 55735 3285 55740 3315
rect 55620 3275 55740 3285
rect 55620 3245 55625 3275
rect 55655 3245 55665 3275
rect 55695 3245 55705 3275
rect 55735 3245 55740 3275
rect 55620 2185 55740 3245
rect 56510 3345 56550 3350
rect 56510 3315 56515 3345
rect 56545 3315 56550 3345
rect 56510 3305 56550 3315
rect 56510 3275 56515 3305
rect 56545 3275 56550 3305
rect 56510 3265 56550 3275
rect 56510 3235 56515 3265
rect 56545 3235 56550 3265
rect 56510 3230 56550 3235
rect 56680 3345 56710 3350
rect 56680 3305 56710 3315
rect 56680 3265 56710 3275
rect 56680 3230 56710 3235
rect 56840 3345 56880 3350
rect 56840 3315 56845 3345
rect 56875 3315 56880 3345
rect 56840 3305 56880 3315
rect 56840 3275 56845 3305
rect 56875 3275 56880 3305
rect 56840 3265 56880 3275
rect 56840 3235 56845 3265
rect 56875 3235 56880 3265
rect 56840 3230 56880 3235
rect 56920 3345 56960 3350
rect 56920 3315 56925 3345
rect 56955 3315 56960 3345
rect 56920 3305 56960 3315
rect 56920 3275 56925 3305
rect 56955 3275 56960 3305
rect 56920 3265 56960 3275
rect 56920 3235 56925 3265
rect 56955 3235 56960 3265
rect 56920 3230 56960 3235
rect 57090 3345 57120 3350
rect 57090 3305 57120 3315
rect 57090 3265 57120 3275
rect 57090 3230 57120 3235
rect 57250 3345 57290 3350
rect 57250 3315 57255 3345
rect 57285 3315 57290 3345
rect 57250 3305 57290 3315
rect 57250 3275 57255 3305
rect 57285 3275 57290 3305
rect 57250 3265 57290 3275
rect 57250 3235 57255 3265
rect 57285 3235 57290 3265
rect 57250 3230 57290 3235
rect 58055 3325 58060 3355
rect 58090 3325 58100 3355
rect 58130 3325 58140 3355
rect 58170 3325 58175 3355
rect 58055 3315 58175 3325
rect 58055 3285 58060 3315
rect 58090 3285 58100 3315
rect 58130 3285 58140 3315
rect 58170 3285 58175 3315
rect 58055 3275 58175 3285
rect 58055 3245 58060 3275
rect 58090 3245 58100 3275
rect 58130 3245 58140 3275
rect 58170 3245 58175 3275
rect 56620 3210 56660 3215
rect 56620 3180 56625 3210
rect 56655 3180 56660 3210
rect 56620 3175 56660 3180
rect 56730 3210 56770 3215
rect 56730 3180 56735 3210
rect 56765 3180 56770 3210
rect 56730 3175 56770 3180
rect 57030 3210 57070 3215
rect 57030 3180 57035 3210
rect 57065 3180 57070 3210
rect 57030 3175 57070 3180
rect 57140 3210 57180 3215
rect 57140 3180 57145 3210
rect 57175 3180 57180 3210
rect 57140 3175 57180 3180
rect 56560 2900 56590 2905
rect 56800 2900 56830 2905
rect 56560 2865 56590 2870
rect 56607 2885 56637 2895
rect 56607 2865 56612 2885
rect 56632 2865 56637 2885
rect 56607 2855 56637 2865
rect 56675 2890 56715 2895
rect 56675 2860 56680 2890
rect 56710 2860 56715 2890
rect 56675 2855 56715 2860
rect 56753 2885 56783 2895
rect 56753 2865 56758 2885
rect 56778 2865 56783 2885
rect 56800 2865 56830 2870
rect 56970 2895 57000 2905
rect 57210 2895 57240 2905
rect 56970 2875 56975 2895
rect 56995 2875 57000 2895
rect 56970 2865 57000 2875
rect 57017 2885 57047 2895
rect 57017 2865 57022 2885
rect 57042 2865 57047 2885
rect 56753 2855 56783 2865
rect 56610 2835 56630 2855
rect 56600 2830 56640 2835
rect 56600 2800 56605 2830
rect 56635 2800 56640 2830
rect 56600 2795 56640 2800
rect 56760 2785 56780 2855
rect 55940 2780 55980 2785
rect 55940 2750 55945 2780
rect 55975 2750 55980 2780
rect 55940 2745 55980 2750
rect 56745 2780 56785 2785
rect 56745 2750 56750 2780
rect 56780 2750 56785 2780
rect 56745 2745 56785 2750
rect 55620 2155 55625 2185
rect 55655 2155 55665 2185
rect 55695 2155 55705 2185
rect 55735 2155 55740 2185
rect 55620 2145 55740 2155
rect 55620 2115 55625 2145
rect 55655 2115 55665 2145
rect 55695 2115 55705 2145
rect 55735 2115 55740 2145
rect 55620 2105 55740 2115
rect 55620 2075 55625 2105
rect 55655 2075 55665 2105
rect 55695 2075 55705 2105
rect 55735 2075 55740 2105
rect 54610 1475 54650 1480
rect 54610 1445 54615 1475
rect 54645 1445 54650 1475
rect 54610 1440 54650 1445
rect 54810 1475 54850 1480
rect 54810 1445 54815 1475
rect 54845 1445 54850 1475
rect 54810 1440 54850 1445
rect 54920 1475 54960 1480
rect 54920 1445 54925 1475
rect 54955 1445 54960 1475
rect 54920 1440 54960 1445
rect 55030 1475 55070 1480
rect 55030 1445 55035 1475
rect 55065 1445 55070 1475
rect 55030 1440 55070 1445
rect 55140 1475 55180 1480
rect 55140 1445 55145 1475
rect 55175 1445 55180 1475
rect 55140 1440 55180 1445
rect 55250 1475 55290 1480
rect 55250 1445 55255 1475
rect 55285 1445 55290 1475
rect 55250 1440 55290 1445
rect 54620 1160 54640 1440
rect 54705 1425 54735 1435
rect 54610 1155 54650 1160
rect 54610 1125 54615 1155
rect 54645 1125 54650 1155
rect 54610 1120 54650 1125
rect 54705 1155 54710 1425
rect 54730 1155 54735 1425
rect 54705 1115 54735 1155
rect 54705 1095 54710 1115
rect 54730 1095 54735 1115
rect 54455 1085 54495 1090
rect 54455 1055 54460 1085
rect 54490 1055 54495 1085
rect 54455 1050 54495 1055
rect 54565 1085 54605 1090
rect 54565 1055 54570 1085
rect 54600 1055 54605 1085
rect 54565 1050 54605 1055
rect 54705 945 54735 1095
rect 54760 1425 54790 1435
rect 54760 1155 54765 1425
rect 54785 1155 54790 1425
rect 54760 1080 54790 1155
rect 54815 1425 54845 1440
rect 54815 1155 54820 1425
rect 54840 1155 54845 1425
rect 54815 1140 54845 1155
rect 54870 1425 54900 1435
rect 54870 1155 54875 1425
rect 54895 1155 54900 1425
rect 54810 1135 54850 1140
rect 54810 1105 54815 1135
rect 54845 1105 54850 1135
rect 54810 1100 54850 1105
rect 54870 1080 54900 1155
rect 54925 1425 54955 1440
rect 54925 1155 54930 1425
rect 54950 1155 54955 1425
rect 54925 1140 54955 1155
rect 54980 1425 55010 1435
rect 54980 1155 54985 1425
rect 55005 1155 55010 1425
rect 54920 1135 54960 1140
rect 54920 1105 54925 1135
rect 54955 1105 54960 1135
rect 54920 1100 54960 1105
rect 54980 1080 55010 1155
rect 55035 1425 55065 1440
rect 55035 1155 55040 1425
rect 55060 1155 55065 1425
rect 55035 1140 55065 1155
rect 55090 1425 55120 1435
rect 55090 1155 55095 1425
rect 55115 1155 55120 1425
rect 55030 1135 55070 1140
rect 55030 1105 55035 1135
rect 55065 1105 55070 1135
rect 55030 1100 55070 1105
rect 55090 1080 55120 1155
rect 55145 1425 55175 1440
rect 55145 1155 55150 1425
rect 55170 1155 55175 1425
rect 55145 1140 55175 1155
rect 55200 1425 55230 1435
rect 55200 1155 55205 1425
rect 55225 1155 55230 1425
rect 55140 1135 55180 1140
rect 55140 1105 55145 1135
rect 55175 1105 55180 1135
rect 55140 1100 55180 1105
rect 55200 1080 55230 1155
rect 55255 1425 55285 1440
rect 55255 1155 55260 1425
rect 55280 1155 55285 1425
rect 55255 1140 55285 1155
rect 55310 1425 55340 1435
rect 55310 1155 55315 1425
rect 55335 1155 55340 1425
rect 55250 1135 55290 1140
rect 55250 1105 55255 1135
rect 55285 1105 55290 1135
rect 55250 1100 55290 1105
rect 55310 1080 55340 1155
rect 55365 1425 55395 1435
rect 55365 1155 55370 1425
rect 55390 1155 55395 1425
rect 55365 1115 55395 1155
rect 55365 1095 55370 1115
rect 55390 1095 55395 1115
rect 54755 1075 54795 1080
rect 54755 1045 54760 1075
rect 54790 1045 54795 1075
rect 54755 1035 54795 1045
rect 54755 1005 54760 1035
rect 54790 1005 54795 1035
rect 54755 995 54795 1005
rect 54755 965 54760 995
rect 54790 965 54795 995
rect 54755 960 54795 965
rect 54865 1075 54905 1080
rect 54865 1045 54870 1075
rect 54900 1045 54905 1075
rect 54865 1035 54905 1045
rect 54865 1005 54870 1035
rect 54900 1005 54905 1035
rect 54865 995 54905 1005
rect 54865 965 54870 995
rect 54900 965 54905 995
rect 54865 960 54905 965
rect 54975 1075 55015 1080
rect 54975 1045 54980 1075
rect 55010 1045 55015 1075
rect 54975 1035 55015 1045
rect 54975 1005 54980 1035
rect 55010 1005 55015 1035
rect 54975 995 55015 1005
rect 54975 965 54980 995
rect 55010 965 55015 995
rect 54975 960 55015 965
rect 55085 1075 55125 1080
rect 55085 1045 55090 1075
rect 55120 1045 55125 1075
rect 55085 1035 55125 1045
rect 55085 1005 55090 1035
rect 55120 1005 55125 1035
rect 55085 995 55125 1005
rect 55085 965 55090 995
rect 55120 965 55125 995
rect 55085 960 55125 965
rect 55195 1075 55235 1080
rect 55195 1045 55200 1075
rect 55230 1045 55235 1075
rect 55195 1035 55235 1045
rect 55195 1005 55200 1035
rect 55230 1005 55235 1035
rect 55195 995 55235 1005
rect 55195 965 55200 995
rect 55230 965 55235 995
rect 55195 960 55235 965
rect 55305 1075 55345 1080
rect 55305 1045 55310 1075
rect 55340 1045 55345 1075
rect 55305 1035 55345 1045
rect 55305 1005 55310 1035
rect 55340 1005 55345 1035
rect 55305 995 55345 1005
rect 55305 965 55310 995
rect 55340 965 55345 995
rect 55305 960 55345 965
rect 55365 945 55395 1095
rect 55620 1075 55740 2075
rect 55895 1985 55935 1990
rect 55895 1955 55900 1985
rect 55930 1955 55935 1985
rect 55895 1950 55935 1955
rect 55620 1045 55625 1075
rect 55655 1045 55665 1075
rect 55695 1045 55705 1075
rect 55735 1045 55740 1075
rect 55620 1035 55740 1045
rect 55620 1005 55625 1035
rect 55655 1005 55665 1035
rect 55695 1005 55705 1035
rect 55735 1005 55740 1035
rect 55620 995 55740 1005
rect 55620 965 55625 995
rect 55655 965 55665 995
rect 55695 965 55705 995
rect 55735 965 55740 995
rect 55620 960 55740 965
rect 55755 1485 55875 1490
rect 55755 1455 55760 1485
rect 55790 1455 55800 1485
rect 55830 1455 55840 1485
rect 55870 1455 55875 1485
rect 55755 1445 55875 1455
rect 55755 1415 55760 1445
rect 55790 1415 55800 1445
rect 55830 1415 55840 1445
rect 55870 1415 55875 1445
rect 55755 1405 55875 1415
rect 55755 1375 55760 1405
rect 55790 1375 55800 1405
rect 55830 1375 55840 1405
rect 55870 1375 55875 1405
rect 54700 940 54740 945
rect 54700 910 54705 940
rect 54735 910 54740 940
rect 54700 900 54740 910
rect 54700 870 54705 900
rect 54735 870 54740 900
rect 54700 860 54740 870
rect 54700 830 54705 860
rect 54735 830 54740 860
rect 54700 825 54740 830
rect 55360 940 55400 945
rect 55360 910 55365 940
rect 55395 910 55400 940
rect 55360 900 55400 910
rect 55360 870 55365 900
rect 55395 870 55400 900
rect 55360 860 55400 870
rect 55360 830 55365 860
rect 55395 830 55400 860
rect 55360 825 55400 830
rect 54335 805 54375 810
rect 54335 775 54340 805
rect 54370 775 54375 805
rect 54335 770 54375 775
rect 54400 435 54440 440
rect 54400 405 54405 435
rect 54435 405 54440 435
rect 54400 400 54440 405
rect 55080 435 55120 440
rect 55080 405 55085 435
rect 55115 405 55120 435
rect 55080 400 55120 405
rect 54070 280 54075 310
rect 54105 280 54115 310
rect 54145 280 54160 310
rect 54190 280 54200 310
rect 54230 280 54245 310
rect 54275 280 54285 310
rect 54315 280 54320 310
rect 54070 270 54320 280
rect 54070 240 54075 270
rect 54105 240 54115 270
rect 54145 240 54160 270
rect 54190 240 54200 270
rect 54230 240 54245 270
rect 54275 240 54285 270
rect 54315 240 54320 270
rect 54070 230 54320 240
rect 54070 200 54075 230
rect 54105 200 54115 230
rect 54145 200 54160 230
rect 54190 200 54200 230
rect 54230 200 54245 230
rect 54275 200 54285 230
rect 54315 200 54320 230
rect 54070 195 54320 200
rect 54410 180 54430 400
rect 54465 310 54505 315
rect 54465 280 54470 310
rect 54500 280 54505 310
rect 54465 270 54505 280
rect 54465 240 54470 270
rect 54500 240 54505 270
rect 54465 230 54505 240
rect 54465 200 54470 230
rect 54500 200 54505 230
rect 54465 195 54505 200
rect 54830 310 55270 315
rect 54830 280 54835 310
rect 54865 280 54875 310
rect 54905 280 54915 310
rect 54945 280 54955 310
rect 54985 280 54995 310
rect 55025 280 55035 310
rect 55065 280 55075 310
rect 55105 280 55115 310
rect 55145 280 55155 310
rect 55185 280 55195 310
rect 55225 280 55235 310
rect 55265 280 55270 310
rect 54830 270 55270 280
rect 54830 240 54835 270
rect 54865 240 54875 270
rect 54905 240 54915 270
rect 54945 240 54955 270
rect 54985 240 54995 270
rect 55025 240 55035 270
rect 55065 240 55075 270
rect 55105 240 55115 270
rect 55145 240 55155 270
rect 55185 240 55195 270
rect 55225 240 55235 270
rect 55265 240 55270 270
rect 54830 230 55270 240
rect 54830 200 54835 230
rect 54865 200 54875 230
rect 54905 200 54915 230
rect 54945 200 54955 230
rect 54985 200 54995 230
rect 55025 200 55035 230
rect 55065 200 55075 230
rect 55105 200 55115 230
rect 55145 200 55155 230
rect 55185 200 55195 230
rect 55225 200 55235 230
rect 55265 200 55270 230
rect 54830 195 55270 200
rect 54405 175 54440 180
rect 54405 135 54440 140
rect 54465 175 54500 195
rect 54465 135 54500 140
rect 54735 165 54765 175
rect 54735 -505 54740 165
rect 54760 -505 54765 165
rect 54735 -545 54765 -505
rect 54835 165 54865 195
rect 54835 -505 54840 165
rect 54860 -505 54865 165
rect 54835 -520 54865 -505
rect 54935 165 54965 175
rect 54935 -505 54940 165
rect 54960 -505 54965 165
rect 54735 -565 54740 -545
rect 54760 -565 54765 -545
rect 54830 -525 54870 -520
rect 54830 -555 54835 -525
rect 54865 -555 54870 -525
rect 54830 -560 54870 -555
rect 54735 -575 54765 -565
rect 54935 -575 54965 -505
rect 55035 165 55065 195
rect 55035 -505 55040 165
rect 55060 -505 55065 165
rect 55035 -520 55065 -505
rect 55135 165 55165 175
rect 55135 -505 55140 165
rect 55160 -505 55165 165
rect 55030 -525 55070 -520
rect 55030 -555 55035 -525
rect 55065 -555 55070 -525
rect 55030 -560 55070 -555
rect 55135 -575 55165 -505
rect 55235 165 55265 195
rect 55235 -505 55240 165
rect 55260 -505 55265 165
rect 55235 -520 55265 -505
rect 55335 165 55365 175
rect 55335 -505 55340 165
rect 55360 -505 55365 165
rect 55755 -95 55875 1375
rect 55755 -125 55760 -95
rect 55790 -125 55800 -95
rect 55830 -125 55840 -95
rect 55870 -125 55875 -95
rect 55755 -135 55875 -125
rect 55755 -165 55760 -135
rect 55790 -165 55800 -135
rect 55830 -165 55840 -135
rect 55870 -165 55875 -135
rect 55755 -175 55875 -165
rect 55755 -205 55760 -175
rect 55790 -205 55800 -175
rect 55830 -205 55840 -175
rect 55870 -205 55875 -175
rect 55755 -210 55875 -205
rect 55905 -270 55925 1950
rect 55950 810 55970 2745
rect 56970 2730 56990 2865
rect 57017 2855 57047 2865
rect 57085 2890 57125 2895
rect 57085 2860 57090 2890
rect 57120 2860 57125 2890
rect 57085 2855 57125 2860
rect 57163 2885 57193 2895
rect 57163 2865 57168 2885
rect 57188 2865 57193 2885
rect 57210 2875 57215 2895
rect 57235 2875 57240 2895
rect 57210 2865 57240 2875
rect 57163 2855 57193 2865
rect 57020 2785 57040 2855
rect 57170 2835 57190 2855
rect 57160 2830 57200 2835
rect 57160 2800 57165 2830
rect 57195 2800 57200 2830
rect 57160 2795 57200 2800
rect 57015 2780 57055 2785
rect 57015 2750 57020 2780
rect 57050 2750 57055 2780
rect 57015 2745 57055 2750
rect 56850 2725 56890 2730
rect 56850 2695 56855 2725
rect 56885 2695 56890 2725
rect 56850 2690 56890 2695
rect 56960 2725 57000 2730
rect 56960 2695 56965 2725
rect 56995 2695 57000 2725
rect 56960 2690 57000 2695
rect 56860 2620 56880 2690
rect 57220 2675 57240 2865
rect 57820 2780 57860 2785
rect 57820 2750 57825 2780
rect 57855 2750 57860 2780
rect 57820 2745 57860 2750
rect 56935 2670 56975 2675
rect 56935 2640 56940 2670
rect 56970 2640 56975 2670
rect 56935 2635 56975 2640
rect 57210 2670 57250 2675
rect 57210 2640 57215 2670
rect 57245 2640 57250 2670
rect 57210 2635 57250 2640
rect 56945 2620 56965 2635
rect 56830 2615 56890 2620
rect 56830 2585 56855 2615
rect 56885 2585 56890 2615
rect 56830 2580 56890 2585
rect 56935 2610 56975 2620
rect 56935 2590 56945 2610
rect 56965 2590 56975 2610
rect 56935 2580 56975 2590
rect 56775 2550 56805 2560
rect 56085 2470 56675 2475
rect 56085 2440 56090 2470
rect 56120 2440 56145 2470
rect 56175 2440 56200 2470
rect 56230 2440 56255 2470
rect 56285 2440 56310 2470
rect 56340 2440 56365 2470
rect 56395 2440 56420 2470
rect 56450 2440 56475 2470
rect 56505 2440 56530 2470
rect 56560 2440 56585 2470
rect 56615 2440 56640 2470
rect 56670 2440 56675 2470
rect 56085 2430 56675 2440
rect 56085 2400 56090 2430
rect 56120 2400 56145 2430
rect 56175 2400 56200 2430
rect 56230 2400 56255 2430
rect 56285 2400 56310 2430
rect 56340 2400 56365 2430
rect 56395 2400 56420 2430
rect 56450 2400 56475 2430
rect 56505 2400 56530 2430
rect 56560 2400 56585 2430
rect 56615 2400 56640 2430
rect 56670 2400 56675 2430
rect 56085 2390 56675 2400
rect 56085 2360 56090 2390
rect 56120 2360 56145 2390
rect 56175 2360 56200 2390
rect 56230 2360 56255 2390
rect 56285 2360 56310 2390
rect 56340 2360 56365 2390
rect 56395 2360 56420 2390
rect 56450 2360 56475 2390
rect 56505 2360 56530 2390
rect 56560 2360 56585 2390
rect 56615 2360 56640 2390
rect 56670 2360 56675 2390
rect 56085 2355 56675 2360
rect 55995 1985 56025 1990
rect 55995 1950 56025 1955
rect 56085 1930 56125 2355
rect 56140 1975 56180 1980
rect 56140 1945 56145 1975
rect 56175 1945 56180 1975
rect 56140 1940 56180 1945
rect 56085 1900 56090 1930
rect 56120 1900 56125 1930
rect 56085 1895 56125 1900
rect 56030 1880 56065 1890
rect 56030 1760 56040 1880
rect 56060 1760 56065 1880
rect 56030 1750 56065 1760
rect 56035 1745 56065 1750
rect 56090 1880 56120 1895
rect 56090 1760 56095 1880
rect 56115 1760 56120 1880
rect 56035 1720 56065 1730
rect 56035 1700 56040 1720
rect 56060 1700 56065 1720
rect 56090 1700 56120 1760
rect 56145 1880 56175 1940
rect 56195 1930 56235 2355
rect 56250 1975 56290 1980
rect 56250 1945 56255 1975
rect 56285 1945 56290 1975
rect 56250 1940 56290 1945
rect 56195 1900 56200 1930
rect 56230 1900 56235 1930
rect 56195 1895 56235 1900
rect 56145 1760 56150 1880
rect 56170 1760 56175 1880
rect 56145 1745 56175 1760
rect 56200 1880 56230 1895
rect 56200 1760 56205 1880
rect 56225 1760 56230 1880
rect 56140 1740 56180 1745
rect 56140 1710 56145 1740
rect 56175 1710 56180 1740
rect 56140 1705 56180 1710
rect 56035 1645 56065 1700
rect 56085 1695 56125 1700
rect 56085 1665 56090 1695
rect 56120 1665 56125 1695
rect 56085 1660 56125 1665
rect 56030 1640 56070 1645
rect 56030 1610 56035 1640
rect 56065 1610 56070 1640
rect 56030 1600 56070 1610
rect 56030 1570 56035 1600
rect 56065 1570 56070 1600
rect 56030 1560 56070 1570
rect 56030 1530 56035 1560
rect 56065 1530 56070 1560
rect 56030 1525 56070 1530
rect 56145 1315 56175 1705
rect 56200 1700 56230 1760
rect 56255 1880 56285 1940
rect 56305 1930 56345 2355
rect 56360 1975 56400 1980
rect 56360 1945 56365 1975
rect 56395 1945 56400 1975
rect 56360 1940 56400 1945
rect 56305 1900 56310 1930
rect 56340 1900 56345 1930
rect 56305 1895 56345 1900
rect 56255 1760 56260 1880
rect 56280 1760 56285 1880
rect 56255 1745 56285 1760
rect 56310 1880 56340 1895
rect 56310 1760 56315 1880
rect 56335 1760 56340 1880
rect 56250 1740 56290 1745
rect 56250 1710 56255 1740
rect 56285 1710 56290 1740
rect 56250 1705 56290 1710
rect 56195 1695 56235 1700
rect 56195 1665 56200 1695
rect 56230 1665 56235 1695
rect 56195 1660 56235 1665
rect 56085 1305 56125 1310
rect 56040 1295 56070 1300
rect 56085 1275 56090 1305
rect 56120 1275 56125 1305
rect 56255 1315 56285 1705
rect 56310 1700 56340 1760
rect 56365 1880 56395 1940
rect 56415 1930 56455 2355
rect 56470 1975 56510 1980
rect 56470 1945 56475 1975
rect 56505 1945 56510 1975
rect 56470 1940 56510 1945
rect 56415 1900 56420 1930
rect 56450 1900 56455 1930
rect 56415 1895 56455 1900
rect 56365 1760 56370 1880
rect 56390 1760 56395 1880
rect 56365 1745 56395 1760
rect 56420 1880 56450 1895
rect 56420 1760 56425 1880
rect 56445 1760 56450 1880
rect 56360 1740 56400 1745
rect 56360 1710 56365 1740
rect 56395 1710 56400 1740
rect 56360 1705 56400 1710
rect 56305 1695 56345 1700
rect 56305 1665 56310 1695
rect 56340 1665 56345 1695
rect 56305 1660 56345 1665
rect 56145 1280 56175 1285
rect 56195 1305 56235 1310
rect 56085 1270 56125 1275
rect 56195 1275 56200 1305
rect 56230 1275 56235 1305
rect 56365 1315 56395 1705
rect 56420 1700 56450 1760
rect 56475 1880 56505 1940
rect 56525 1930 56565 2355
rect 56580 1975 56620 1980
rect 56580 1945 56585 1975
rect 56615 1945 56620 1975
rect 56580 1940 56620 1945
rect 56525 1900 56530 1930
rect 56560 1900 56565 1930
rect 56525 1895 56565 1900
rect 56475 1760 56480 1880
rect 56500 1760 56505 1880
rect 56475 1745 56505 1760
rect 56530 1880 56560 1895
rect 56530 1760 56535 1880
rect 56555 1760 56560 1880
rect 56470 1740 56510 1745
rect 56470 1710 56475 1740
rect 56505 1710 56510 1740
rect 56470 1705 56510 1710
rect 56415 1695 56455 1700
rect 56415 1665 56420 1695
rect 56450 1665 56455 1695
rect 56415 1660 56455 1665
rect 56255 1280 56285 1285
rect 56305 1305 56345 1310
rect 56195 1270 56235 1275
rect 56305 1275 56310 1305
rect 56340 1275 56345 1305
rect 56475 1315 56505 1705
rect 56530 1700 56560 1760
rect 56585 1880 56615 1940
rect 56635 1930 56675 2355
rect 56775 2330 56780 2550
rect 56800 2330 56805 2550
rect 56775 2300 56805 2330
rect 56830 2550 56860 2580
rect 56830 2330 56835 2550
rect 56855 2330 56860 2550
rect 56830 2320 56860 2330
rect 56885 2550 56915 2560
rect 56885 2330 56890 2550
rect 56910 2330 56915 2550
rect 56885 2300 56915 2330
rect 56940 2550 56970 2580
rect 56940 2330 56945 2550
rect 56965 2330 56970 2550
rect 56940 2320 56970 2330
rect 56995 2550 57025 2560
rect 56995 2330 57000 2550
rect 57020 2330 57025 2550
rect 56995 2300 57025 2330
rect 57125 2470 57715 2475
rect 57125 2440 57130 2470
rect 57160 2440 57185 2470
rect 57215 2440 57240 2470
rect 57270 2440 57295 2470
rect 57325 2440 57350 2470
rect 57380 2440 57405 2470
rect 57435 2440 57460 2470
rect 57490 2440 57515 2470
rect 57545 2440 57570 2470
rect 57600 2440 57625 2470
rect 57655 2440 57680 2470
rect 57710 2440 57715 2470
rect 57125 2430 57715 2440
rect 57125 2400 57130 2430
rect 57160 2400 57185 2430
rect 57215 2400 57240 2430
rect 57270 2400 57295 2430
rect 57325 2400 57350 2430
rect 57380 2400 57405 2430
rect 57435 2400 57460 2430
rect 57490 2400 57515 2430
rect 57545 2400 57570 2430
rect 57600 2400 57625 2430
rect 57655 2400 57680 2430
rect 57710 2400 57715 2430
rect 57125 2390 57715 2400
rect 57125 2360 57130 2390
rect 57160 2360 57185 2390
rect 57215 2360 57240 2390
rect 57270 2360 57295 2390
rect 57325 2360 57350 2390
rect 57380 2360 57405 2390
rect 57435 2360 57460 2390
rect 57490 2360 57515 2390
rect 57545 2360 57570 2390
rect 57600 2360 57625 2390
rect 57655 2360 57680 2390
rect 57710 2360 57715 2390
rect 57125 2355 57715 2360
rect 56770 2295 56810 2300
rect 56770 2265 56775 2295
rect 56805 2265 56810 2295
rect 56770 2255 56810 2265
rect 56770 2225 56775 2255
rect 56805 2225 56810 2255
rect 56770 2215 56810 2225
rect 56770 2185 56775 2215
rect 56805 2185 56810 2215
rect 56770 2180 56810 2185
rect 56880 2295 56920 2300
rect 56880 2265 56885 2295
rect 56915 2265 56920 2295
rect 56880 2255 56920 2265
rect 56880 2225 56885 2255
rect 56915 2225 56920 2255
rect 56880 2215 56920 2225
rect 56880 2185 56885 2215
rect 56915 2185 56920 2215
rect 56880 2180 56920 2185
rect 56990 2295 57030 2300
rect 56990 2265 56995 2295
rect 57025 2265 57030 2295
rect 56990 2255 57030 2265
rect 56990 2225 56995 2255
rect 57025 2225 57030 2255
rect 56990 2215 57030 2225
rect 56990 2185 56995 2215
rect 57025 2185 57030 2215
rect 56990 2180 57030 2185
rect 56690 1985 56720 1990
rect 56690 1950 56720 1955
rect 57080 1985 57110 1990
rect 57080 1950 57110 1955
rect 56635 1900 56640 1930
rect 56670 1900 56675 1930
rect 56635 1895 56675 1900
rect 57125 1930 57165 2355
rect 57180 1975 57220 1980
rect 57180 1945 57185 1975
rect 57215 1945 57220 1975
rect 57180 1940 57220 1945
rect 57125 1900 57130 1930
rect 57160 1900 57165 1930
rect 57125 1895 57165 1900
rect 56585 1760 56590 1880
rect 56610 1760 56615 1880
rect 56585 1745 56615 1760
rect 56640 1880 56670 1895
rect 56640 1760 56645 1880
rect 56665 1760 56670 1880
rect 56580 1740 56620 1745
rect 56580 1710 56585 1740
rect 56615 1710 56620 1740
rect 56580 1705 56620 1710
rect 56525 1695 56565 1700
rect 56525 1665 56530 1695
rect 56560 1665 56565 1695
rect 56525 1660 56565 1665
rect 56365 1280 56395 1285
rect 56415 1305 56455 1310
rect 56305 1270 56345 1275
rect 56415 1275 56420 1305
rect 56450 1275 56455 1305
rect 56585 1315 56615 1705
rect 56640 1700 56670 1760
rect 56695 1880 56765 1890
rect 56695 1760 56700 1880
rect 56720 1760 56765 1880
rect 56695 1750 56765 1760
rect 57035 1880 57105 1890
rect 57035 1760 57080 1880
rect 57100 1760 57105 1880
rect 57035 1750 57105 1760
rect 56695 1720 56725 1750
rect 56695 1700 56700 1720
rect 56720 1700 56725 1720
rect 56635 1695 56675 1700
rect 56635 1665 56640 1695
rect 56670 1665 56675 1695
rect 56635 1660 56675 1665
rect 56695 1645 56725 1700
rect 57075 1720 57105 1750
rect 57075 1700 57080 1720
rect 57100 1700 57105 1720
rect 57130 1880 57160 1895
rect 57130 1760 57135 1880
rect 57155 1760 57160 1880
rect 57130 1700 57160 1760
rect 57185 1880 57215 1940
rect 57235 1930 57275 2355
rect 57290 1975 57330 1980
rect 57290 1945 57295 1975
rect 57325 1945 57330 1975
rect 57290 1940 57330 1945
rect 57235 1900 57240 1930
rect 57270 1900 57275 1930
rect 57235 1895 57275 1900
rect 57185 1760 57190 1880
rect 57210 1760 57215 1880
rect 57185 1745 57215 1760
rect 57240 1880 57270 1895
rect 57240 1760 57245 1880
rect 57265 1760 57270 1880
rect 57180 1740 57220 1745
rect 57180 1710 57185 1740
rect 57215 1710 57220 1740
rect 57180 1705 57220 1710
rect 57075 1645 57105 1700
rect 57125 1695 57165 1700
rect 57125 1665 57130 1695
rect 57160 1665 57165 1695
rect 57125 1660 57165 1665
rect 56690 1640 56730 1645
rect 56690 1610 56695 1640
rect 56725 1610 56730 1640
rect 56690 1600 56730 1610
rect 56690 1570 56695 1600
rect 56725 1570 56730 1600
rect 56690 1560 56730 1570
rect 56690 1530 56695 1560
rect 56725 1530 56730 1560
rect 56690 1525 56730 1530
rect 57070 1640 57110 1645
rect 57070 1610 57075 1640
rect 57105 1610 57110 1640
rect 57070 1600 57110 1610
rect 57070 1570 57075 1600
rect 57105 1570 57110 1600
rect 57070 1560 57110 1570
rect 57070 1530 57075 1560
rect 57105 1530 57110 1560
rect 57070 1525 57110 1530
rect 56880 1485 56920 1490
rect 56880 1455 56885 1485
rect 56915 1455 56920 1485
rect 56880 1445 56920 1455
rect 56880 1415 56885 1445
rect 56915 1415 56920 1445
rect 56880 1405 56920 1415
rect 56880 1375 56885 1405
rect 56915 1375 56920 1405
rect 56880 1370 56920 1375
rect 56475 1280 56505 1285
rect 56525 1305 56565 1310
rect 56415 1270 56455 1275
rect 56525 1275 56530 1305
rect 56560 1275 56565 1305
rect 56585 1280 56615 1285
rect 56635 1305 56675 1310
rect 56525 1270 56565 1275
rect 56635 1275 56640 1305
rect 56670 1275 56675 1305
rect 56635 1270 56675 1275
rect 56690 1305 56720 1310
rect 56690 1270 56720 1275
rect 56840 1305 56870 1310
rect 56840 1270 56870 1275
rect 56040 1260 56070 1265
rect 56035 1205 56065 1215
rect 56035 1085 56040 1205
rect 56060 1085 56065 1205
rect 56035 1075 56065 1085
rect 56090 1205 56120 1270
rect 56140 1260 56180 1265
rect 56140 1230 56145 1260
rect 56175 1230 56180 1260
rect 56140 1225 56180 1230
rect 56090 1085 56095 1205
rect 56115 1085 56120 1205
rect 56090 1070 56120 1085
rect 56145 1205 56175 1225
rect 56145 1085 56150 1205
rect 56170 1085 56175 1205
rect 56085 1065 56125 1070
rect 56035 1045 56065 1055
rect 56035 1025 56040 1045
rect 56060 1025 56065 1045
rect 56085 1035 56090 1065
rect 56120 1035 56125 1065
rect 56085 1030 56125 1035
rect 56035 1015 56065 1025
rect 56040 945 56060 1015
rect 56145 1000 56175 1085
rect 56200 1205 56230 1270
rect 56250 1260 56290 1265
rect 56250 1230 56255 1260
rect 56285 1230 56290 1260
rect 56250 1225 56290 1230
rect 56200 1085 56205 1205
rect 56225 1085 56230 1205
rect 56200 1070 56230 1085
rect 56255 1205 56285 1225
rect 56255 1085 56260 1205
rect 56280 1085 56285 1205
rect 56195 1065 56235 1070
rect 56195 1035 56200 1065
rect 56230 1035 56235 1065
rect 56195 1030 56235 1035
rect 56255 1000 56285 1085
rect 56310 1205 56340 1270
rect 56360 1260 56400 1265
rect 56360 1230 56365 1260
rect 56395 1230 56400 1260
rect 56360 1225 56400 1230
rect 56310 1085 56315 1205
rect 56335 1085 56340 1205
rect 56310 1070 56340 1085
rect 56365 1205 56395 1225
rect 56365 1085 56370 1205
rect 56390 1085 56395 1205
rect 56305 1065 56345 1070
rect 56305 1035 56310 1065
rect 56340 1035 56345 1065
rect 56305 1030 56345 1035
rect 56365 1000 56395 1085
rect 56420 1205 56450 1270
rect 56470 1260 56510 1265
rect 56470 1230 56475 1260
rect 56505 1230 56510 1260
rect 56470 1225 56510 1230
rect 56420 1085 56425 1205
rect 56445 1085 56450 1205
rect 56420 1070 56450 1085
rect 56475 1205 56505 1225
rect 56475 1085 56480 1205
rect 56500 1085 56505 1205
rect 56415 1065 56455 1070
rect 56415 1035 56420 1065
rect 56450 1035 56455 1065
rect 56415 1030 56455 1035
rect 56475 1000 56505 1085
rect 56530 1205 56560 1270
rect 56580 1260 56620 1265
rect 56580 1230 56585 1260
rect 56615 1230 56620 1260
rect 56580 1225 56620 1230
rect 56530 1085 56535 1205
rect 56555 1085 56560 1205
rect 56530 1070 56560 1085
rect 56585 1205 56615 1225
rect 56585 1085 56590 1205
rect 56610 1085 56615 1205
rect 56525 1065 56565 1070
rect 56525 1035 56530 1065
rect 56560 1035 56565 1065
rect 56525 1030 56565 1035
rect 56585 1000 56615 1085
rect 56640 1205 56670 1270
rect 56640 1085 56645 1205
rect 56665 1085 56670 1205
rect 56640 1070 56670 1085
rect 56695 1205 56805 1215
rect 56695 1085 56700 1205
rect 56720 1085 56780 1205
rect 56800 1085 56805 1205
rect 56695 1075 56805 1085
rect 56830 1205 56860 1215
rect 56830 1085 56835 1205
rect 56855 1085 56860 1205
rect 56635 1065 56675 1070
rect 56635 1035 56640 1065
rect 56670 1035 56675 1065
rect 56740 1055 56760 1075
rect 56830 1070 56860 1085
rect 56885 1205 56915 1370
rect 57185 1315 57215 1705
rect 57240 1700 57270 1760
rect 57295 1880 57325 1940
rect 57345 1930 57385 2355
rect 57400 1975 57440 1980
rect 57400 1945 57405 1975
rect 57435 1945 57440 1975
rect 57400 1940 57440 1945
rect 57345 1900 57350 1930
rect 57380 1900 57385 1930
rect 57345 1895 57385 1900
rect 57295 1760 57300 1880
rect 57320 1760 57325 1880
rect 57295 1745 57325 1760
rect 57350 1880 57380 1895
rect 57350 1760 57355 1880
rect 57375 1760 57380 1880
rect 57290 1740 57330 1745
rect 57290 1710 57295 1740
rect 57325 1710 57330 1740
rect 57290 1705 57330 1710
rect 57235 1695 57275 1700
rect 57235 1665 57240 1695
rect 57270 1665 57275 1695
rect 57235 1660 57275 1665
rect 56930 1305 56960 1310
rect 56930 1270 56960 1275
rect 57080 1305 57110 1310
rect 57080 1270 57110 1275
rect 57125 1305 57165 1310
rect 57125 1275 57130 1305
rect 57160 1275 57165 1305
rect 57295 1315 57325 1705
rect 57350 1700 57380 1760
rect 57405 1880 57435 1940
rect 57455 1930 57495 2355
rect 57510 1975 57550 1980
rect 57510 1945 57515 1975
rect 57545 1945 57550 1975
rect 57510 1940 57550 1945
rect 57455 1900 57460 1930
rect 57490 1900 57495 1930
rect 57455 1895 57495 1900
rect 57405 1760 57410 1880
rect 57430 1760 57435 1880
rect 57405 1745 57435 1760
rect 57460 1880 57490 1895
rect 57460 1760 57465 1880
rect 57485 1760 57490 1880
rect 57400 1740 57440 1745
rect 57400 1710 57405 1740
rect 57435 1710 57440 1740
rect 57400 1705 57440 1710
rect 57345 1695 57385 1700
rect 57345 1665 57350 1695
rect 57380 1665 57385 1695
rect 57345 1660 57385 1665
rect 57185 1280 57215 1285
rect 57235 1305 57275 1310
rect 57125 1270 57165 1275
rect 57235 1275 57240 1305
rect 57270 1275 57275 1305
rect 57405 1315 57435 1705
rect 57460 1700 57490 1760
rect 57515 1880 57545 1940
rect 57565 1930 57605 2355
rect 57620 1975 57660 1980
rect 57620 1945 57625 1975
rect 57655 1945 57660 1975
rect 57620 1940 57660 1945
rect 57565 1900 57570 1930
rect 57600 1900 57605 1930
rect 57565 1895 57605 1900
rect 57515 1760 57520 1880
rect 57540 1760 57545 1880
rect 57515 1745 57545 1760
rect 57570 1880 57600 1895
rect 57570 1760 57575 1880
rect 57595 1760 57600 1880
rect 57510 1740 57550 1745
rect 57510 1710 57515 1740
rect 57545 1710 57550 1740
rect 57510 1705 57550 1710
rect 57455 1695 57495 1700
rect 57455 1665 57460 1695
rect 57490 1665 57495 1695
rect 57455 1660 57495 1665
rect 57295 1280 57325 1285
rect 57345 1305 57385 1310
rect 57235 1270 57275 1275
rect 57345 1275 57350 1305
rect 57380 1275 57385 1305
rect 57515 1315 57545 1705
rect 57570 1700 57600 1760
rect 57625 1880 57655 1940
rect 57675 1930 57715 2355
rect 57675 1900 57680 1930
rect 57710 1900 57715 1930
rect 57675 1895 57715 1900
rect 57625 1760 57630 1880
rect 57650 1760 57655 1880
rect 57625 1745 57655 1760
rect 57680 1880 57710 1895
rect 57680 1760 57685 1880
rect 57705 1760 57710 1880
rect 57620 1740 57660 1745
rect 57620 1710 57625 1740
rect 57655 1710 57660 1740
rect 57620 1705 57660 1710
rect 57565 1695 57605 1700
rect 57565 1665 57570 1695
rect 57600 1665 57605 1695
rect 57565 1660 57605 1665
rect 57405 1280 57435 1285
rect 57455 1305 57495 1310
rect 57345 1270 57385 1275
rect 57455 1275 57460 1305
rect 57490 1275 57495 1305
rect 57625 1315 57655 1705
rect 57680 1700 57710 1760
rect 57735 1880 57765 1890
rect 57735 1760 57740 1880
rect 57760 1760 57765 1880
rect 57735 1750 57765 1760
rect 57735 1720 57765 1730
rect 57735 1700 57740 1720
rect 57760 1700 57765 1720
rect 57675 1695 57715 1700
rect 57675 1665 57680 1695
rect 57710 1665 57715 1695
rect 57675 1660 57715 1665
rect 57735 1645 57765 1700
rect 57730 1640 57770 1645
rect 57730 1610 57735 1640
rect 57765 1610 57770 1640
rect 57730 1600 57770 1610
rect 57730 1570 57735 1600
rect 57765 1570 57770 1600
rect 57730 1560 57770 1570
rect 57730 1530 57735 1560
rect 57765 1530 57770 1560
rect 57730 1525 57770 1530
rect 57515 1280 57545 1285
rect 57565 1305 57605 1310
rect 57455 1270 57495 1275
rect 57565 1275 57570 1305
rect 57600 1275 57605 1305
rect 57625 1280 57655 1285
rect 57675 1305 57715 1310
rect 57565 1270 57605 1275
rect 57675 1275 57680 1305
rect 57710 1275 57715 1305
rect 57675 1270 57715 1275
rect 57730 1295 57760 1300
rect 56885 1085 56890 1205
rect 56910 1085 56915 1205
rect 56885 1075 56915 1085
rect 56940 1205 56970 1215
rect 56940 1085 56945 1205
rect 56965 1085 56970 1205
rect 56940 1070 56970 1085
rect 56995 1205 57105 1215
rect 56995 1085 57000 1205
rect 57020 1085 57080 1205
rect 57100 1085 57105 1205
rect 56995 1075 57105 1085
rect 57130 1205 57160 1270
rect 57180 1260 57220 1265
rect 57180 1230 57185 1260
rect 57215 1230 57220 1260
rect 57180 1225 57220 1230
rect 57130 1085 57135 1205
rect 57155 1085 57160 1205
rect 56825 1065 56865 1070
rect 56635 1030 56675 1035
rect 56735 1045 56765 1055
rect 56735 1025 56740 1045
rect 56760 1025 56765 1045
rect 56735 1015 56765 1025
rect 56825 1035 56830 1065
rect 56860 1035 56865 1065
rect 56140 995 56180 1000
rect 56140 965 56145 995
rect 56175 965 56180 995
rect 56140 960 56180 965
rect 56250 995 56290 1000
rect 56250 965 56255 995
rect 56285 965 56290 995
rect 56250 960 56290 965
rect 56360 995 56400 1000
rect 56360 965 56365 995
rect 56395 965 56400 995
rect 56360 960 56400 965
rect 56440 995 56700 1000
rect 56440 965 56475 995
rect 56505 965 56585 995
rect 56615 965 56700 995
rect 56030 940 56070 945
rect 56030 910 56035 940
rect 56065 910 56070 940
rect 56030 900 56070 910
rect 56030 870 56035 900
rect 56065 870 56070 900
rect 56030 860 56070 870
rect 56030 830 56035 860
rect 56065 830 56070 860
rect 56030 825 56070 830
rect 55940 805 55980 810
rect 55940 775 55945 805
rect 55975 775 55980 805
rect 55940 770 55980 775
rect 56440 390 56700 965
rect 56740 945 56760 1015
rect 56730 940 56770 945
rect 56730 910 56735 940
rect 56765 910 56770 940
rect 56730 900 56770 910
rect 56730 870 56735 900
rect 56765 870 56770 900
rect 56730 860 56770 870
rect 56730 830 56735 860
rect 56765 830 56770 860
rect 56730 825 56770 830
rect 56440 360 56445 390
rect 56475 360 56555 390
rect 56585 360 56665 390
rect 56695 360 56700 390
rect 56440 355 56700 360
rect 56770 390 56810 395
rect 56770 360 56775 390
rect 56805 360 56810 390
rect 56770 355 56810 360
rect 56825 375 56865 1035
rect 56935 1065 56975 1070
rect 56935 1035 56940 1065
rect 56970 1035 56975 1065
rect 57040 1055 57060 1075
rect 57130 1070 57160 1085
rect 57185 1205 57215 1225
rect 57185 1085 57190 1205
rect 57210 1085 57215 1205
rect 57125 1065 57165 1070
rect 56825 355 56835 375
rect 56855 355 56865 375
rect 56880 390 56920 395
rect 56880 360 56885 390
rect 56915 360 56920 390
rect 56880 355 56920 360
rect 56935 375 56975 1035
rect 57035 1045 57065 1055
rect 57035 1025 57040 1045
rect 57060 1025 57065 1045
rect 57125 1035 57130 1065
rect 57160 1035 57165 1065
rect 57125 1030 57165 1035
rect 57035 1015 57065 1025
rect 57040 945 57060 1015
rect 57185 1000 57215 1085
rect 57240 1205 57270 1270
rect 57290 1260 57330 1265
rect 57290 1230 57295 1260
rect 57325 1230 57330 1260
rect 57290 1225 57330 1230
rect 57240 1085 57245 1205
rect 57265 1085 57270 1205
rect 57240 1070 57270 1085
rect 57295 1205 57325 1225
rect 57295 1085 57300 1205
rect 57320 1085 57325 1205
rect 57235 1065 57275 1070
rect 57235 1035 57240 1065
rect 57270 1035 57275 1065
rect 57235 1030 57275 1035
rect 57295 1000 57325 1085
rect 57350 1205 57380 1270
rect 57400 1260 57440 1265
rect 57400 1230 57405 1260
rect 57435 1230 57440 1260
rect 57400 1225 57440 1230
rect 57350 1085 57355 1205
rect 57375 1085 57380 1205
rect 57350 1070 57380 1085
rect 57405 1205 57435 1225
rect 57405 1085 57410 1205
rect 57430 1085 57435 1205
rect 57345 1065 57385 1070
rect 57345 1035 57350 1065
rect 57380 1035 57385 1065
rect 57345 1030 57385 1035
rect 57405 1000 57435 1085
rect 57460 1205 57490 1270
rect 57510 1260 57550 1265
rect 57510 1230 57515 1260
rect 57545 1230 57550 1260
rect 57510 1225 57550 1230
rect 57460 1085 57465 1205
rect 57485 1085 57490 1205
rect 57460 1070 57490 1085
rect 57515 1205 57545 1225
rect 57515 1085 57520 1205
rect 57540 1085 57545 1205
rect 57455 1065 57495 1070
rect 57455 1035 57460 1065
rect 57490 1035 57495 1065
rect 57455 1030 57495 1035
rect 57515 1000 57545 1085
rect 57570 1205 57600 1270
rect 57620 1260 57660 1265
rect 57620 1230 57625 1260
rect 57655 1230 57660 1260
rect 57620 1225 57660 1230
rect 57570 1085 57575 1205
rect 57595 1085 57600 1205
rect 57570 1070 57600 1085
rect 57625 1205 57655 1225
rect 57625 1085 57630 1205
rect 57650 1085 57655 1205
rect 57565 1065 57605 1070
rect 57565 1035 57570 1065
rect 57600 1035 57605 1065
rect 57565 1030 57605 1035
rect 57625 1000 57655 1085
rect 57680 1205 57710 1270
rect 57730 1260 57760 1265
rect 57680 1085 57685 1205
rect 57705 1085 57710 1205
rect 57680 1070 57710 1085
rect 57735 1205 57765 1215
rect 57735 1085 57740 1205
rect 57760 1085 57765 1205
rect 57735 1075 57765 1085
rect 57675 1065 57715 1070
rect 57675 1035 57680 1065
rect 57710 1035 57715 1065
rect 57675 1030 57715 1035
rect 57735 1045 57765 1055
rect 57735 1025 57740 1045
rect 57760 1025 57765 1045
rect 57735 1015 57765 1025
rect 57100 995 57360 1000
rect 57100 965 57185 995
rect 57215 965 57295 995
rect 57325 965 57360 995
rect 57030 940 57070 945
rect 57030 910 57035 940
rect 57065 910 57070 940
rect 57030 900 57070 910
rect 57030 870 57035 900
rect 57065 870 57070 900
rect 57030 860 57070 870
rect 57030 830 57035 860
rect 57065 830 57070 860
rect 57030 825 57070 830
rect 56935 355 56945 375
rect 56965 355 56975 375
rect 56990 390 57030 395
rect 56990 360 56995 390
rect 57025 360 57030 390
rect 56990 355 57030 360
rect 57100 390 57360 965
rect 57400 995 57440 1000
rect 57400 965 57405 995
rect 57435 965 57440 995
rect 57400 960 57440 965
rect 57510 995 57550 1000
rect 57510 965 57515 995
rect 57545 965 57550 995
rect 57510 960 57550 965
rect 57620 995 57660 1000
rect 57620 965 57625 995
rect 57655 965 57660 995
rect 57620 960 57660 965
rect 57740 945 57760 1015
rect 57730 940 57770 945
rect 57730 910 57735 940
rect 57765 910 57770 940
rect 57730 900 57770 910
rect 57730 870 57735 900
rect 57765 870 57770 900
rect 57730 860 57770 870
rect 57730 830 57735 860
rect 57765 830 57770 860
rect 57730 825 57770 830
rect 57830 810 57850 2745
rect 57865 2670 57905 2675
rect 57865 2640 57870 2670
rect 57900 2640 57905 2670
rect 57865 2635 57905 2640
rect 57820 805 57860 810
rect 57820 775 57825 805
rect 57855 775 57860 805
rect 57820 770 57860 775
rect 57100 360 57105 390
rect 57135 360 57215 390
rect 57245 360 57325 390
rect 57355 360 57360 390
rect 57100 355 57360 360
rect 57430 390 57470 395
rect 57430 360 57435 390
rect 57465 360 57470 390
rect 57430 355 57470 360
rect 56185 315 56255 325
rect 56185 95 56230 315
rect 56250 95 56255 315
rect 56185 85 56255 95
rect 56225 65 56255 85
rect 56280 315 56310 325
rect 56280 95 56285 315
rect 56305 95 56310 315
rect 56280 65 56310 95
rect 56335 315 56365 325
rect 56335 95 56340 315
rect 56360 95 56365 315
rect 56220 60 56260 65
rect 56220 30 56225 60
rect 56255 30 56260 60
rect 55895 -275 55935 -270
rect 55895 -305 55900 -275
rect 55930 -305 55935 -275
rect 55895 -310 55935 -305
rect 55230 -525 55270 -520
rect 55230 -555 55235 -525
rect 55265 -555 55270 -525
rect 55230 -560 55270 -555
rect 55335 -545 55365 -505
rect 55335 -565 55340 -545
rect 55360 -565 55365 -545
rect 55335 -575 55365 -565
rect 56220 -575 56260 30
rect 56275 60 56315 65
rect 56275 30 56280 60
rect 56310 30 56315 60
rect 56275 25 56315 30
rect 56335 -90 56365 95
rect 56390 315 56420 325
rect 56390 95 56395 315
rect 56415 95 56420 315
rect 56390 65 56420 95
rect 56445 315 56475 355
rect 56445 95 56450 315
rect 56470 95 56475 315
rect 56385 60 56425 65
rect 56385 30 56390 60
rect 56420 30 56425 60
rect 56385 25 56425 30
rect 56445 20 56475 95
rect 56500 315 56530 325
rect 56500 95 56505 315
rect 56525 95 56530 315
rect 56500 65 56530 95
rect 56555 315 56585 355
rect 56555 95 56560 315
rect 56580 95 56585 315
rect 56495 60 56535 65
rect 56495 30 56500 60
rect 56530 30 56535 60
rect 56495 25 56535 30
rect 56555 20 56585 95
rect 56610 315 56640 325
rect 56610 95 56615 315
rect 56635 95 56640 315
rect 56610 65 56640 95
rect 56665 315 56695 355
rect 56665 95 56670 315
rect 56690 95 56695 315
rect 56605 60 56645 65
rect 56605 30 56610 60
rect 56640 30 56645 60
rect 56605 25 56645 30
rect 56665 20 56695 95
rect 56720 315 56750 325
rect 56720 95 56725 315
rect 56745 95 56750 315
rect 56720 65 56750 95
rect 56775 315 56805 355
rect 56825 345 56865 355
rect 56775 95 56780 315
rect 56800 95 56805 315
rect 56715 60 56755 65
rect 56715 30 56720 60
rect 56750 30 56755 60
rect 56715 25 56755 30
rect 56775 20 56805 95
rect 56830 315 56860 325
rect 56830 95 56835 315
rect 56855 95 56860 315
rect 56830 65 56860 95
rect 56885 315 56915 355
rect 56935 345 56975 355
rect 56885 95 56890 315
rect 56910 95 56915 315
rect 56825 60 56865 65
rect 56825 30 56830 60
rect 56860 30 56865 60
rect 56825 25 56865 30
rect 56885 20 56915 95
rect 56940 315 56970 325
rect 56940 95 56945 315
rect 56965 95 56970 315
rect 56940 65 56970 95
rect 56995 315 57025 355
rect 56995 95 57000 315
rect 57020 95 57025 315
rect 56935 60 56975 65
rect 56935 30 56940 60
rect 56970 30 56975 60
rect 56935 25 56975 30
rect 56995 20 57025 95
rect 57050 315 57080 325
rect 57050 95 57055 315
rect 57075 95 57080 315
rect 57050 65 57080 95
rect 57105 315 57135 355
rect 57105 95 57110 315
rect 57130 95 57135 315
rect 57045 60 57085 65
rect 57045 30 57050 60
rect 57080 30 57085 60
rect 57045 25 57085 30
rect 57105 20 57135 95
rect 57160 315 57190 325
rect 57160 95 57165 315
rect 57185 95 57190 315
rect 57160 65 57190 95
rect 57215 315 57245 355
rect 57215 95 57220 315
rect 57240 95 57245 315
rect 57155 60 57195 65
rect 57155 30 57160 60
rect 57190 30 57195 60
rect 57155 25 57195 30
rect 57215 20 57245 95
rect 57270 315 57300 325
rect 57270 95 57275 315
rect 57295 95 57300 315
rect 57270 65 57300 95
rect 57325 315 57355 355
rect 57325 95 57330 315
rect 57350 95 57355 315
rect 57265 60 57305 65
rect 57265 30 57270 60
rect 57300 30 57305 60
rect 57265 25 57305 30
rect 57325 20 57355 95
rect 57380 315 57410 325
rect 57380 95 57385 315
rect 57405 95 57410 315
rect 57380 65 57410 95
rect 57435 315 57465 355
rect 57435 95 57440 315
rect 57460 95 57465 315
rect 57375 60 57415 65
rect 57375 30 57380 60
rect 57410 30 57415 60
rect 57375 25 57415 30
rect 57435 20 57465 95
rect 57490 315 57520 325
rect 57490 95 57495 315
rect 57515 95 57520 315
rect 57490 65 57520 95
rect 57485 60 57525 65
rect 57485 30 57490 60
rect 57520 30 57525 60
rect 56440 15 56480 20
rect 56440 -15 56445 15
rect 56475 -15 56480 15
rect 56440 -20 56480 -15
rect 56550 15 56590 20
rect 56550 -15 56555 15
rect 56585 -15 56590 15
rect 56550 -20 56590 -15
rect 56660 15 56700 20
rect 56660 -15 56665 15
rect 56695 -15 56700 15
rect 56660 -20 56700 -15
rect 56770 15 56810 20
rect 56770 -15 56775 15
rect 56805 -15 56810 15
rect 56770 -20 56810 -15
rect 56880 15 56920 20
rect 56880 -15 56885 15
rect 56915 -15 56920 15
rect 56880 -20 56920 -15
rect 56990 15 57030 20
rect 56990 -15 56995 15
rect 57025 -15 57030 15
rect 56990 -20 57030 -15
rect 57100 15 57140 20
rect 57100 -15 57105 15
rect 57135 -15 57140 15
rect 57100 -20 57140 -15
rect 57210 15 57250 20
rect 57210 -15 57215 15
rect 57245 -15 57250 15
rect 57210 -20 57250 -15
rect 57320 15 57360 20
rect 57320 -15 57325 15
rect 57355 -15 57360 15
rect 57320 -20 57360 -15
rect 57430 15 57470 20
rect 57430 -15 57435 15
rect 57465 -15 57470 15
rect 57430 -20 57470 -15
rect 56330 -95 56370 -90
rect 56330 -125 56335 -95
rect 56365 -125 56370 -95
rect 56330 -135 56370 -125
rect 56330 -165 56335 -135
rect 56365 -165 56370 -135
rect 56330 -175 56370 -165
rect 56330 -205 56335 -175
rect 56365 -205 56370 -175
rect 56330 -210 56370 -205
rect 56540 -230 56580 -225
rect 56540 -260 56545 -230
rect 56575 -260 56580 -230
rect 56540 -265 56580 -260
rect 56650 -230 56690 -225
rect 56650 -260 56655 -230
rect 56685 -260 56690 -230
rect 56650 -265 56690 -260
rect 56870 -230 56910 -225
rect 56870 -260 56875 -230
rect 56905 -260 56910 -230
rect 56870 -265 56910 -260
rect 56485 -275 56525 -270
rect 56485 -305 56490 -275
rect 56520 -305 56525 -275
rect 56485 -310 56525 -305
rect 56395 -340 56465 -330
rect 56395 -460 56440 -340
rect 56460 -460 56465 -340
rect 56395 -470 56465 -460
rect 56435 -500 56465 -470
rect 56435 -520 56440 -500
rect 56460 -520 56465 -500
rect 56490 -340 56520 -310
rect 56490 -460 56495 -340
rect 56515 -460 56520 -340
rect 56490 -520 56520 -460
rect 56545 -340 56575 -265
rect 56595 -275 56635 -270
rect 56595 -305 56600 -275
rect 56630 -305 56635 -275
rect 56595 -310 56635 -305
rect 56545 -460 56550 -340
rect 56570 -460 56575 -340
rect 56545 -475 56575 -460
rect 56600 -340 56630 -310
rect 56600 -460 56605 -340
rect 56625 -460 56630 -340
rect 56540 -480 56580 -475
rect 56540 -510 56545 -480
rect 56575 -510 56580 -480
rect 56540 -515 56580 -510
rect 56600 -520 56630 -460
rect 56655 -340 56685 -265
rect 56705 -275 56745 -270
rect 56705 -305 56710 -275
rect 56740 -305 56745 -275
rect 56705 -310 56745 -305
rect 56655 -460 56660 -340
rect 56680 -460 56685 -340
rect 56655 -475 56685 -460
rect 56710 -340 56740 -310
rect 56710 -460 56715 -340
rect 56735 -460 56740 -340
rect 56650 -480 56690 -475
rect 56650 -510 56655 -480
rect 56685 -510 56690 -480
rect 56650 -515 56690 -510
rect 56710 -520 56740 -460
rect 56765 -340 56835 -330
rect 56765 -460 56770 -340
rect 56790 -460 56835 -340
rect 56765 -470 56835 -460
rect 56875 -340 56905 -265
rect 57040 -275 57080 -270
rect 57040 -305 57045 -275
rect 57075 -305 57080 -275
rect 57040 -310 57080 -305
rect 56875 -460 56880 -340
rect 56900 -460 56905 -340
rect 56765 -500 56795 -470
rect 56875 -475 56905 -460
rect 57215 -340 57245 -20
rect 57415 -40 57455 -35
rect 57415 -70 57420 -40
rect 57450 -70 57455 -40
rect 57415 -75 57455 -70
rect 57215 -460 57220 -340
rect 57240 -460 57245 -340
rect 57215 -470 57245 -460
rect 56765 -520 56770 -500
rect 56790 -520 56795 -500
rect 56870 -480 56910 -475
rect 56870 -510 56875 -480
rect 56905 -510 56910 -480
rect 56870 -515 56910 -510
rect 56435 -575 56465 -520
rect 56485 -525 56525 -520
rect 56485 -555 56490 -525
rect 56520 -555 56525 -525
rect 56485 -560 56525 -555
rect 56595 -525 56635 -520
rect 56595 -555 56600 -525
rect 56630 -555 56635 -525
rect 56595 -560 56635 -555
rect 56705 -525 56745 -520
rect 56705 -555 56710 -525
rect 56740 -555 56745 -525
rect 56705 -560 56745 -555
rect 56765 -575 56795 -520
rect 52290 -580 52410 -575
rect 52290 -610 52295 -580
rect 52325 -610 52335 -580
rect 52365 -610 52375 -580
rect 52405 -610 52410 -580
rect 52290 -620 52410 -610
rect 52290 -650 52295 -620
rect 52325 -650 52335 -620
rect 52365 -650 52375 -620
rect 52405 -650 52410 -620
rect 52290 -660 52410 -650
rect 52290 -690 52295 -660
rect 52325 -690 52335 -660
rect 52365 -690 52375 -660
rect 52405 -690 52410 -660
rect 52290 -1500 52410 -690
rect 52640 -580 52760 -575
rect 52640 -610 52645 -580
rect 52675 -610 52685 -580
rect 52715 -610 52725 -580
rect 52755 -610 52760 -580
rect 52640 -620 52760 -610
rect 52640 -650 52645 -620
rect 52675 -650 52685 -620
rect 52715 -650 52725 -620
rect 52755 -650 52760 -620
rect 52640 -660 52760 -650
rect 52640 -690 52645 -660
rect 52675 -690 52685 -660
rect 52715 -690 52725 -660
rect 52755 -690 52760 -660
rect 52640 -1500 52760 -690
rect 52990 -580 53110 -575
rect 52990 -610 52995 -580
rect 53025 -610 53035 -580
rect 53065 -610 53075 -580
rect 53105 -610 53110 -580
rect 52990 -620 53110 -610
rect 52990 -650 52995 -620
rect 53025 -650 53035 -620
rect 53065 -650 53075 -620
rect 53105 -650 53110 -620
rect 52990 -660 53110 -650
rect 52990 -690 52995 -660
rect 53025 -690 53035 -660
rect 53065 -690 53075 -660
rect 53105 -690 53110 -660
rect 52990 -1500 53110 -690
rect 53340 -580 53460 -575
rect 53340 -610 53345 -580
rect 53375 -610 53385 -580
rect 53415 -610 53425 -580
rect 53455 -610 53460 -580
rect 53340 -620 53460 -610
rect 53340 -650 53345 -620
rect 53375 -650 53385 -620
rect 53415 -650 53425 -620
rect 53455 -650 53460 -620
rect 53340 -660 53460 -650
rect 53340 -690 53345 -660
rect 53375 -690 53385 -660
rect 53415 -690 53425 -660
rect 53455 -690 53460 -660
rect 53340 -1500 53460 -690
rect 53690 -580 54160 -575
rect 53690 -610 53695 -580
rect 53725 -610 53735 -580
rect 53765 -610 53775 -580
rect 53805 -610 53925 -580
rect 53955 -610 53965 -580
rect 53995 -610 54005 -580
rect 54035 -610 54045 -580
rect 54075 -610 54085 -580
rect 54115 -610 54125 -580
rect 54155 -610 54160 -580
rect 53690 -620 54160 -610
rect 53690 -650 53695 -620
rect 53725 -650 53735 -620
rect 53765 -650 53775 -620
rect 53805 -650 53925 -620
rect 53955 -650 53965 -620
rect 53995 -650 54005 -620
rect 54035 -650 54045 -620
rect 54075 -650 54085 -620
rect 54115 -650 54125 -620
rect 54155 -650 54160 -620
rect 53690 -660 54160 -650
rect 53690 -690 53695 -660
rect 53725 -690 53735 -660
rect 53765 -690 53775 -660
rect 53805 -690 53925 -660
rect 53955 -690 53965 -660
rect 53995 -690 54005 -660
rect 54035 -690 54045 -660
rect 54075 -690 54085 -660
rect 54115 -690 54125 -660
rect 54155 -690 54160 -660
rect 53690 -695 54160 -690
rect 53690 -1500 53810 -695
rect 54040 -1500 54160 -695
rect 54390 -580 54510 -575
rect 54390 -610 54395 -580
rect 54425 -610 54435 -580
rect 54465 -610 54475 -580
rect 54505 -610 54510 -580
rect 54390 -620 54510 -610
rect 54390 -650 54395 -620
rect 54425 -650 54435 -620
rect 54465 -650 54475 -620
rect 54505 -650 54510 -620
rect 54390 -660 54510 -650
rect 54390 -690 54395 -660
rect 54425 -690 54435 -660
rect 54465 -690 54475 -660
rect 54505 -690 54510 -660
rect 54390 -1500 54510 -690
rect 54735 -580 54860 -575
rect 54735 -610 54745 -580
rect 54775 -610 54785 -580
rect 54815 -610 54825 -580
rect 54855 -610 54860 -580
rect 54735 -620 54860 -610
rect 54735 -650 54745 -620
rect 54775 -650 54785 -620
rect 54815 -650 54825 -620
rect 54855 -650 54860 -620
rect 54735 -660 54860 -650
rect 54735 -690 54745 -660
rect 54775 -690 54785 -660
rect 54815 -690 54825 -660
rect 54855 -690 54860 -660
rect 54735 -695 54860 -690
rect 54930 -580 54970 -575
rect 54930 -610 54935 -580
rect 54965 -610 54970 -580
rect 54930 -620 54970 -610
rect 54930 -650 54935 -620
rect 54965 -650 54970 -620
rect 54930 -660 54970 -650
rect 54930 -690 54935 -660
rect 54965 -690 54970 -660
rect 54930 -695 54970 -690
rect 55090 -580 55210 -575
rect 55090 -610 55095 -580
rect 55125 -610 55135 -580
rect 55165 -610 55175 -580
rect 55205 -610 55210 -580
rect 55090 -620 55210 -610
rect 55090 -650 55095 -620
rect 55125 -650 55135 -620
rect 55165 -650 55175 -620
rect 55205 -650 55210 -620
rect 55090 -660 55210 -650
rect 55090 -690 55095 -660
rect 55125 -690 55135 -660
rect 55165 -690 55175 -660
rect 55205 -690 55210 -660
rect 54740 -1500 54860 -695
rect 55090 -1500 55210 -690
rect 55320 -580 55560 -575
rect 55320 -610 55325 -580
rect 55355 -610 55365 -580
rect 55395 -610 55405 -580
rect 55435 -610 55445 -580
rect 55475 -610 55485 -580
rect 55515 -610 55525 -580
rect 55555 -610 55560 -580
rect 55320 -620 55560 -610
rect 55320 -650 55325 -620
rect 55355 -650 55365 -620
rect 55395 -650 55405 -620
rect 55435 -650 55445 -620
rect 55475 -650 55485 -620
rect 55515 -650 55525 -620
rect 55555 -650 55560 -620
rect 55320 -660 55560 -650
rect 55320 -690 55325 -660
rect 55355 -690 55365 -660
rect 55395 -690 55405 -660
rect 55435 -690 55445 -660
rect 55475 -690 55485 -660
rect 55515 -690 55525 -660
rect 55555 -690 55560 -660
rect 55320 -695 55560 -690
rect 55440 -1500 55560 -695
rect 55790 -580 55910 -575
rect 55790 -610 55795 -580
rect 55825 -610 55835 -580
rect 55865 -610 55875 -580
rect 55905 -610 55910 -580
rect 55790 -620 55910 -610
rect 55790 -650 55795 -620
rect 55825 -650 55835 -620
rect 55865 -650 55875 -620
rect 55905 -650 55910 -620
rect 55790 -660 55910 -650
rect 55790 -690 55795 -660
rect 55825 -690 55835 -660
rect 55865 -690 55875 -660
rect 55905 -690 55910 -660
rect 55790 -1500 55910 -690
rect 56140 -580 56260 -575
rect 56140 -610 56145 -580
rect 56175 -610 56185 -580
rect 56215 -610 56225 -580
rect 56255 -610 56260 -580
rect 56140 -620 56260 -610
rect 56140 -650 56145 -620
rect 56175 -650 56185 -620
rect 56215 -650 56225 -620
rect 56255 -650 56260 -620
rect 56140 -660 56260 -650
rect 56140 -690 56145 -660
rect 56175 -690 56185 -660
rect 56215 -690 56225 -660
rect 56255 -690 56260 -660
rect 56140 -1500 56260 -690
rect 56430 -580 56470 -575
rect 56430 -610 56435 -580
rect 56465 -610 56470 -580
rect 56430 -620 56470 -610
rect 56430 -650 56435 -620
rect 56465 -650 56470 -620
rect 56430 -660 56470 -650
rect 56430 -690 56435 -660
rect 56465 -690 56470 -660
rect 56430 -695 56470 -690
rect 56490 -580 56610 -575
rect 56490 -610 56495 -580
rect 56525 -610 56535 -580
rect 56565 -610 56575 -580
rect 56605 -610 56610 -580
rect 56490 -620 56610 -610
rect 56490 -650 56495 -620
rect 56525 -650 56535 -620
rect 56565 -650 56575 -620
rect 56605 -650 56610 -620
rect 56490 -660 56610 -650
rect 56490 -690 56495 -660
rect 56525 -690 56535 -660
rect 56565 -690 56575 -660
rect 56605 -690 56610 -660
rect 56490 -1500 56610 -690
rect 56760 -580 56800 -575
rect 56760 -610 56765 -580
rect 56795 -610 56800 -580
rect 56760 -620 56800 -610
rect 56760 -650 56765 -620
rect 56795 -650 56800 -620
rect 56760 -660 56800 -650
rect 56760 -690 56765 -660
rect 56795 -690 56800 -660
rect 56760 -695 56800 -690
rect 56840 -580 56960 -575
rect 56840 -610 56845 -580
rect 56875 -610 56885 -580
rect 56915 -610 56925 -580
rect 56955 -610 56960 -580
rect 56840 -620 56960 -610
rect 56840 -650 56845 -620
rect 56875 -650 56885 -620
rect 56915 -650 56925 -620
rect 56955 -650 56960 -620
rect 56840 -660 56960 -650
rect 56840 -690 56845 -660
rect 56875 -690 56885 -660
rect 56915 -690 56925 -660
rect 56955 -690 56960 -660
rect 56840 -1500 56960 -690
rect 57190 -580 57310 -575
rect 57190 -610 57195 -580
rect 57225 -610 57235 -580
rect 57265 -610 57275 -580
rect 57305 -610 57310 -580
rect 57190 -620 57310 -610
rect 57190 -650 57195 -620
rect 57225 -650 57235 -620
rect 57265 -650 57275 -620
rect 57305 -650 57310 -620
rect 57190 -660 57310 -650
rect 57190 -690 57195 -660
rect 57225 -690 57235 -660
rect 57265 -690 57275 -660
rect 57305 -690 57310 -660
rect 57190 -1500 57310 -690
rect 57485 -580 57525 30
rect 57875 -35 57895 2635
rect 57920 2295 58040 2300
rect 57920 2265 57925 2295
rect 57955 2265 57965 2295
rect 57995 2265 58005 2295
rect 58035 2265 58040 2295
rect 57920 2255 58040 2265
rect 57920 2225 57925 2255
rect 57955 2225 57965 2255
rect 57995 2225 58005 2255
rect 58035 2225 58040 2255
rect 57920 2215 58040 2225
rect 57920 2185 57925 2215
rect 57955 2185 57965 2215
rect 57995 2185 58005 2215
rect 58035 2185 58040 2215
rect 57920 2050 58040 2185
rect 57920 2020 57925 2050
rect 57955 2020 57965 2050
rect 57995 2020 58005 2050
rect 58035 2020 58040 2050
rect 57920 2010 58040 2020
rect 57920 1980 57925 2010
rect 57955 1980 57965 2010
rect 57995 1980 58005 2010
rect 58035 1980 58040 2010
rect 57920 1970 58040 1980
rect 57920 1940 57925 1970
rect 57955 1940 57965 1970
rect 57995 1940 58005 1970
rect 58035 1940 58040 1970
rect 57920 1640 58040 1940
rect 57920 1610 57925 1640
rect 57955 1610 57965 1640
rect 57995 1610 58005 1640
rect 58035 1610 58040 1640
rect 57920 1600 58040 1610
rect 57920 1570 57925 1600
rect 57955 1570 57965 1600
rect 57995 1570 58005 1600
rect 58035 1570 58040 1600
rect 57920 1560 58040 1570
rect 57920 1530 57925 1560
rect 57955 1530 57965 1560
rect 57995 1530 58005 1560
rect 58035 1530 58040 1560
rect 57920 1525 58040 1530
rect 58055 2185 58175 3245
rect 58055 2155 58060 2185
rect 58090 2155 58100 2185
rect 58130 2155 58140 2185
rect 58170 2155 58175 2185
rect 58055 2145 58175 2155
rect 58055 2115 58060 2145
rect 58090 2115 58100 2145
rect 58130 2115 58140 2145
rect 58170 2115 58175 2145
rect 58055 2105 58175 2115
rect 58055 2075 58060 2105
rect 58090 2075 58100 2105
rect 58130 2075 58140 2105
rect 58170 2075 58175 2105
rect 57920 1485 58040 1490
rect 57920 1455 57925 1485
rect 57955 1455 57965 1485
rect 57995 1455 58005 1485
rect 58035 1455 58040 1485
rect 57920 1445 58040 1455
rect 57920 1415 57925 1445
rect 57955 1415 57965 1445
rect 57995 1415 58005 1445
rect 58035 1415 58040 1445
rect 57920 1405 58040 1415
rect 57920 1375 57925 1405
rect 57955 1375 57965 1405
rect 57995 1375 58005 1405
rect 58035 1375 58040 1405
rect 57865 -40 57905 -35
rect 57865 -70 57870 -40
rect 57900 -70 57905 -40
rect 57865 -75 57905 -70
rect 57920 -95 58040 1375
rect 58055 1080 58175 2075
rect 58190 3490 58310 3495
rect 58190 3460 58195 3490
rect 58225 3460 58235 3490
rect 58265 3460 58275 3490
rect 58305 3460 58310 3490
rect 58190 3450 58310 3460
rect 58190 3420 58195 3450
rect 58225 3420 58235 3450
rect 58265 3420 58275 3450
rect 58305 3420 58310 3450
rect 58190 3410 58310 3420
rect 58190 3380 58195 3410
rect 58225 3380 58235 3410
rect 58265 3380 58275 3410
rect 58305 3380 58310 3410
rect 58190 2470 58310 3380
rect 59505 3375 59545 3380
rect 58400 3355 58440 3360
rect 58400 3325 58405 3355
rect 58435 3325 58440 3355
rect 58400 3315 58440 3325
rect 58400 3285 58405 3315
rect 58435 3285 58440 3315
rect 58400 3275 58440 3285
rect 58400 3245 58405 3275
rect 58435 3245 58440 3275
rect 58400 3240 58440 3245
rect 58510 3355 58550 3360
rect 58510 3325 58515 3355
rect 58545 3325 58550 3355
rect 58510 3315 58550 3325
rect 58510 3285 58515 3315
rect 58545 3285 58550 3315
rect 58510 3275 58550 3285
rect 58510 3245 58515 3275
rect 58545 3245 58550 3275
rect 58510 3240 58550 3245
rect 58620 3355 58660 3360
rect 58620 3325 58625 3355
rect 58655 3325 58660 3355
rect 58620 3315 58660 3325
rect 58620 3285 58625 3315
rect 58655 3285 58660 3315
rect 58620 3275 58660 3285
rect 58620 3245 58625 3275
rect 58655 3245 58660 3275
rect 58620 3240 58660 3245
rect 58730 3355 58770 3360
rect 58730 3325 58735 3355
rect 58765 3325 58770 3355
rect 58730 3315 58770 3325
rect 58730 3285 58735 3315
rect 58765 3285 58770 3315
rect 58730 3275 58770 3285
rect 58730 3245 58735 3275
rect 58765 3245 58770 3275
rect 58730 3240 58770 3245
rect 58840 3355 58880 3360
rect 58840 3325 58845 3355
rect 58875 3325 58880 3355
rect 58840 3315 58880 3325
rect 58840 3285 58845 3315
rect 58875 3285 58880 3315
rect 58840 3275 58880 3285
rect 58840 3245 58845 3275
rect 58875 3245 58880 3275
rect 58840 3240 58880 3245
rect 58950 3355 58990 3360
rect 58950 3325 58955 3355
rect 58985 3325 58990 3355
rect 58950 3315 58990 3325
rect 58950 3285 58955 3315
rect 58985 3285 58990 3315
rect 58950 3275 58990 3285
rect 58950 3245 58955 3275
rect 58985 3245 58990 3275
rect 58950 3240 58990 3245
rect 59060 3355 59100 3360
rect 59060 3325 59065 3355
rect 59095 3325 59100 3355
rect 59505 3345 59510 3375
rect 59540 3345 59545 3375
rect 59505 3340 59545 3345
rect 59060 3315 59100 3325
rect 59060 3285 59065 3315
rect 59095 3285 59100 3315
rect 59060 3275 59100 3285
rect 59060 3245 59065 3275
rect 59095 3245 59100 3275
rect 59060 3240 59100 3245
rect 58405 3200 58435 3240
rect 58405 3180 58410 3200
rect 58430 3180 58435 3200
rect 58405 3140 58435 3180
rect 58455 3190 58495 3195
rect 58455 3160 58460 3190
rect 58490 3160 58495 3190
rect 58455 3155 58495 3160
rect 58405 2570 58410 3140
rect 58430 2570 58435 3140
rect 58405 2560 58435 2570
rect 58460 3140 58490 3155
rect 58460 2570 58465 3140
rect 58485 2570 58490 3140
rect 58460 2555 58490 2570
rect 58515 3140 58545 3240
rect 58565 3190 58605 3195
rect 58565 3160 58570 3190
rect 58600 3160 58605 3190
rect 58565 3155 58605 3160
rect 58515 2570 58520 3140
rect 58540 2570 58545 3140
rect 58515 2560 58545 2570
rect 58570 3140 58600 3155
rect 58570 2570 58575 3140
rect 58595 2570 58600 3140
rect 58570 2555 58600 2570
rect 58625 3140 58655 3240
rect 58675 3190 58715 3195
rect 58675 3160 58680 3190
rect 58710 3160 58715 3190
rect 58675 3155 58715 3160
rect 58625 2570 58630 3140
rect 58650 2570 58655 3140
rect 58625 2560 58655 2570
rect 58680 3140 58710 3155
rect 58680 2570 58685 3140
rect 58705 2570 58710 3140
rect 58680 2555 58710 2570
rect 58735 3140 58765 3240
rect 58785 3190 58825 3195
rect 58785 3160 58790 3190
rect 58820 3160 58825 3190
rect 58785 3155 58825 3160
rect 58735 2570 58740 3140
rect 58760 2570 58765 3140
rect 58735 2560 58765 2570
rect 58790 3140 58820 3155
rect 58790 2570 58795 3140
rect 58815 2570 58820 3140
rect 58790 2555 58820 2570
rect 58845 3140 58875 3240
rect 58895 3190 58935 3195
rect 58895 3160 58900 3190
rect 58930 3160 58935 3190
rect 58895 3155 58935 3160
rect 58845 2570 58850 3140
rect 58870 2570 58875 3140
rect 58845 2560 58875 2570
rect 58900 3140 58930 3155
rect 58900 2570 58905 3140
rect 58925 2570 58930 3140
rect 58900 2555 58930 2570
rect 58955 3140 58985 3240
rect 59065 3200 59095 3240
rect 59515 3215 59535 3340
rect 59005 3190 59045 3195
rect 59005 3160 59010 3190
rect 59040 3160 59045 3190
rect 59005 3155 59045 3160
rect 59065 3180 59070 3200
rect 59090 3180 59095 3200
rect 58955 2570 58960 3140
rect 58980 2570 58985 3140
rect 58955 2560 58985 2570
rect 59010 3140 59040 3155
rect 59010 2570 59015 3140
rect 59035 2570 59040 3140
rect 59010 2555 59040 2570
rect 59065 3140 59095 3180
rect 59455 3205 59596 3215
rect 59455 3185 59460 3205
rect 59480 3185 59515 3205
rect 59535 3185 59570 3205
rect 59590 3185 59596 3205
rect 59455 3175 59596 3185
rect 59065 2570 59070 3140
rect 59090 2570 59095 3140
rect 59455 2600 59596 2610
rect 59455 2580 59460 2600
rect 59480 2580 59515 2600
rect 59535 2580 59570 2600
rect 59590 2580 59596 2600
rect 59455 2570 59596 2580
rect 59065 2560 59095 2570
rect 58190 2440 58195 2470
rect 58225 2440 58235 2470
rect 58265 2440 58275 2470
rect 58305 2440 58310 2470
rect 58190 2430 58310 2440
rect 58190 2400 58195 2430
rect 58225 2400 58235 2430
rect 58265 2400 58275 2430
rect 58305 2400 58310 2430
rect 58190 2390 58310 2400
rect 58190 2360 58195 2390
rect 58225 2360 58235 2390
rect 58265 2360 58275 2390
rect 58305 2360 58310 2390
rect 58190 1595 58310 2360
rect 58455 2550 58495 2555
rect 58455 2520 58460 2550
rect 58490 2520 58495 2550
rect 58455 2325 58495 2520
rect 58565 2550 58605 2555
rect 58565 2520 58570 2550
rect 58600 2520 58605 2550
rect 58565 2325 58605 2520
rect 58675 2550 58715 2555
rect 58675 2520 58680 2550
rect 58710 2520 58715 2550
rect 58675 2325 58715 2520
rect 58785 2550 58825 2555
rect 58785 2520 58790 2550
rect 58820 2520 58825 2550
rect 58730 2470 58770 2475
rect 58730 2440 58735 2470
rect 58765 2440 58770 2470
rect 58730 2430 58770 2440
rect 58730 2400 58735 2430
rect 58765 2400 58770 2430
rect 58730 2390 58770 2400
rect 58730 2360 58735 2390
rect 58765 2360 58770 2390
rect 58730 2355 58770 2360
rect 58785 2325 58825 2520
rect 58895 2550 58935 2555
rect 58895 2520 58900 2550
rect 58930 2520 58935 2550
rect 58895 2325 58935 2520
rect 59005 2550 59045 2555
rect 59005 2520 59010 2550
rect 59040 2520 59045 2550
rect 59005 2325 59045 2520
rect 59465 2470 59585 2570
rect 59465 2440 59470 2470
rect 59500 2440 59510 2470
rect 59540 2440 59550 2470
rect 59580 2440 59585 2470
rect 59465 2430 59585 2440
rect 59465 2400 59470 2430
rect 59500 2400 59510 2430
rect 59540 2400 59550 2430
rect 59580 2400 59585 2430
rect 59465 2390 59585 2400
rect 59465 2360 59470 2390
rect 59500 2360 59510 2390
rect 59540 2360 59550 2390
rect 59580 2360 59585 2390
rect 59465 2355 59585 2360
rect 58455 2320 59045 2325
rect 58455 2290 58460 2320
rect 58490 2290 58515 2320
rect 58545 2290 58570 2320
rect 58600 2290 58625 2320
rect 58655 2290 58680 2320
rect 58710 2290 58735 2320
rect 58765 2290 58790 2320
rect 58820 2290 58845 2320
rect 58875 2290 58900 2320
rect 58930 2290 58955 2320
rect 58985 2290 59010 2320
rect 59040 2290 59045 2320
rect 58455 2280 59045 2290
rect 58455 2250 58460 2280
rect 58490 2250 58515 2280
rect 58545 2250 58570 2280
rect 58600 2250 58625 2280
rect 58655 2250 58680 2280
rect 58710 2250 58735 2280
rect 58765 2250 58790 2280
rect 58820 2250 58845 2280
rect 58875 2250 58900 2280
rect 58930 2250 58955 2280
rect 58985 2250 59010 2280
rect 59040 2250 59045 2280
rect 58455 2240 59045 2250
rect 58455 2210 58460 2240
rect 58490 2210 58515 2240
rect 58545 2210 58570 2240
rect 58600 2210 58625 2240
rect 58655 2210 58680 2240
rect 58710 2210 58735 2240
rect 58765 2210 58790 2240
rect 58820 2210 58845 2240
rect 58875 2210 58900 2240
rect 58930 2210 58955 2240
rect 58985 2210 59010 2240
rect 59040 2210 59045 2240
rect 58455 2205 59045 2210
rect 59480 2320 59730 2325
rect 59480 2290 59485 2320
rect 59515 2290 59525 2320
rect 59555 2290 59570 2320
rect 59600 2290 59610 2320
rect 59640 2290 59655 2320
rect 59685 2290 59695 2320
rect 59725 2290 59730 2320
rect 59480 2280 59730 2290
rect 59480 2250 59485 2280
rect 59515 2250 59525 2280
rect 59555 2250 59570 2280
rect 59600 2250 59610 2280
rect 59640 2250 59655 2280
rect 59685 2250 59695 2280
rect 59725 2250 59730 2280
rect 59480 2240 59730 2250
rect 59480 2210 59485 2240
rect 59515 2210 59525 2240
rect 59555 2210 59570 2240
rect 59600 2210 59610 2240
rect 59640 2210 59655 2240
rect 59685 2210 59695 2240
rect 59725 2210 59730 2240
rect 58400 2185 58440 2190
rect 58400 2155 58405 2185
rect 58435 2155 58440 2185
rect 58400 2145 58440 2155
rect 58400 2115 58405 2145
rect 58435 2115 58440 2145
rect 58400 2105 58440 2115
rect 58400 2075 58405 2105
rect 58435 2075 58440 2105
rect 58400 2070 58440 2075
rect 59060 2185 59100 2190
rect 59060 2155 59065 2185
rect 59095 2155 59100 2185
rect 59060 2145 59100 2155
rect 59060 2115 59065 2145
rect 59095 2115 59100 2145
rect 59060 2105 59100 2115
rect 59060 2075 59065 2105
rect 59095 2075 59100 2105
rect 59060 2070 59100 2075
rect 58405 1925 58435 2070
rect 58455 2050 58495 2055
rect 58455 2020 58460 2050
rect 58490 2020 58495 2050
rect 58455 2010 58495 2020
rect 58455 1980 58460 2010
rect 58490 1980 58495 2010
rect 58455 1970 58495 1980
rect 58455 1940 58460 1970
rect 58490 1940 58495 1970
rect 58455 1935 58495 1940
rect 58565 2050 58605 2055
rect 58565 2020 58570 2050
rect 58600 2020 58605 2050
rect 58565 2010 58605 2020
rect 58565 1980 58570 2010
rect 58600 1980 58605 2010
rect 58565 1970 58605 1980
rect 58565 1940 58570 1970
rect 58600 1940 58605 1970
rect 58565 1935 58605 1940
rect 58675 2050 58715 2055
rect 58675 2020 58680 2050
rect 58710 2020 58715 2050
rect 58675 2010 58715 2020
rect 58675 1980 58680 2010
rect 58710 1980 58715 2010
rect 58675 1970 58715 1980
rect 58675 1940 58680 1970
rect 58710 1940 58715 1970
rect 58675 1935 58715 1940
rect 58785 2050 58825 2055
rect 58785 2020 58790 2050
rect 58820 2020 58825 2050
rect 58785 2010 58825 2020
rect 58785 1980 58790 2010
rect 58820 1980 58825 2010
rect 58785 1970 58825 1980
rect 58785 1940 58790 1970
rect 58820 1940 58825 1970
rect 58785 1935 58825 1940
rect 58895 2050 58935 2055
rect 58895 2020 58900 2050
rect 58930 2020 58935 2050
rect 58895 2010 58935 2020
rect 58895 1980 58900 2010
rect 58930 1980 58935 2010
rect 58895 1970 58935 1980
rect 58895 1940 58900 1970
rect 58930 1940 58935 1970
rect 58895 1935 58935 1940
rect 59005 2050 59045 2055
rect 59005 2020 59010 2050
rect 59040 2020 59045 2050
rect 59005 2010 59045 2020
rect 59005 1980 59010 2010
rect 59040 1980 59045 2010
rect 59005 1970 59045 1980
rect 59005 1940 59010 1970
rect 59040 1940 59045 1970
rect 59005 1935 59045 1940
rect 58405 1905 58410 1925
rect 58430 1905 58435 1925
rect 58405 1865 58435 1905
rect 58405 1695 58410 1865
rect 58430 1695 58435 1865
rect 58405 1685 58435 1695
rect 58460 1865 58490 1935
rect 58510 1915 58550 1920
rect 58510 1885 58515 1915
rect 58545 1885 58550 1915
rect 58510 1880 58550 1885
rect 58460 1695 58465 1865
rect 58485 1695 58490 1865
rect 58460 1685 58490 1695
rect 58515 1865 58545 1880
rect 58515 1695 58520 1865
rect 58540 1695 58545 1865
rect 58515 1665 58545 1695
rect 58570 1865 58600 1935
rect 58620 1915 58660 1920
rect 58620 1885 58625 1915
rect 58655 1885 58660 1915
rect 58620 1880 58660 1885
rect 58570 1695 58575 1865
rect 58595 1695 58600 1865
rect 58570 1685 58600 1695
rect 58625 1865 58655 1880
rect 58625 1695 58630 1865
rect 58650 1695 58655 1865
rect 58625 1665 58655 1695
rect 58680 1865 58710 1935
rect 58730 1915 58770 1920
rect 58730 1885 58735 1915
rect 58765 1885 58770 1915
rect 58730 1880 58770 1885
rect 58680 1695 58685 1865
rect 58705 1695 58710 1865
rect 58680 1685 58710 1695
rect 58735 1865 58765 1880
rect 58735 1695 58740 1865
rect 58760 1695 58765 1865
rect 58735 1665 58765 1695
rect 58790 1865 58820 1935
rect 58840 1915 58880 1920
rect 58840 1885 58845 1915
rect 58875 1885 58880 1915
rect 58840 1880 58880 1885
rect 58790 1695 58795 1865
rect 58815 1695 58820 1865
rect 58790 1685 58820 1695
rect 58845 1865 58875 1880
rect 58845 1695 58850 1865
rect 58870 1695 58875 1865
rect 58845 1665 58875 1695
rect 58900 1865 58930 1935
rect 58950 1915 58990 1920
rect 58950 1885 58955 1915
rect 58985 1885 58990 1915
rect 58950 1880 58990 1885
rect 58900 1695 58905 1865
rect 58925 1695 58930 1865
rect 58900 1685 58930 1695
rect 58955 1865 58985 1880
rect 58955 1695 58960 1865
rect 58980 1695 58985 1865
rect 58955 1665 58985 1695
rect 59010 1865 59040 1935
rect 59010 1695 59015 1865
rect 59035 1695 59040 1865
rect 59010 1685 59040 1695
rect 59065 1925 59095 2070
rect 59065 1905 59070 1925
rect 59090 1905 59095 1925
rect 59065 1865 59095 1905
rect 59065 1695 59070 1865
rect 59090 1695 59095 1865
rect 59065 1685 59095 1695
rect 59480 1710 59730 2210
rect 59480 1680 59490 1710
rect 59520 1680 59540 1710
rect 59570 1680 59590 1710
rect 59620 1680 59640 1710
rect 59670 1680 59690 1710
rect 59720 1680 59730 1710
rect 58510 1660 58550 1665
rect 58510 1630 58515 1660
rect 58545 1630 58550 1660
rect 58510 1625 58550 1630
rect 58620 1660 58660 1665
rect 58620 1630 58625 1660
rect 58655 1630 58660 1660
rect 58620 1625 58660 1630
rect 58730 1660 58770 1665
rect 58730 1630 58735 1660
rect 58765 1630 58770 1660
rect 58730 1625 58770 1630
rect 58840 1660 58880 1665
rect 58840 1630 58845 1660
rect 58875 1630 58880 1660
rect 58840 1625 58880 1630
rect 58950 1660 58990 1665
rect 58950 1630 58955 1660
rect 58985 1630 58990 1660
rect 58950 1625 58990 1630
rect 59195 1660 59235 1665
rect 59195 1630 59200 1660
rect 59230 1630 59235 1660
rect 59195 1625 59235 1630
rect 59480 1660 59730 1680
rect 59480 1630 59490 1660
rect 59520 1630 59540 1660
rect 59570 1630 59590 1660
rect 59620 1630 59640 1660
rect 59670 1630 59690 1660
rect 59720 1630 59730 1660
rect 58190 1565 58195 1595
rect 58225 1565 58235 1595
rect 58265 1565 58275 1595
rect 58305 1565 58310 1595
rect 58190 1555 58310 1565
rect 58190 1525 58195 1555
rect 58225 1525 58235 1555
rect 58265 1525 58275 1555
rect 58305 1525 58310 1555
rect 58190 1520 58310 1525
rect 58565 1595 58605 1600
rect 58565 1565 58570 1595
rect 58600 1565 58605 1595
rect 58565 1555 58605 1565
rect 58565 1525 58570 1555
rect 58600 1525 58605 1555
rect 58565 1520 58605 1525
rect 58510 1475 58550 1480
rect 58510 1445 58515 1475
rect 58545 1445 58550 1475
rect 58510 1440 58550 1445
rect 58620 1475 58660 1480
rect 58620 1445 58625 1475
rect 58655 1445 58660 1475
rect 58620 1440 58660 1445
rect 58730 1475 58770 1480
rect 58730 1445 58735 1475
rect 58765 1445 58770 1475
rect 58730 1440 58770 1445
rect 58840 1475 58880 1480
rect 58840 1445 58845 1475
rect 58875 1445 58880 1475
rect 58840 1440 58880 1445
rect 58950 1475 58990 1480
rect 58950 1445 58955 1475
rect 58985 1445 58990 1475
rect 58950 1440 58990 1445
rect 59150 1475 59190 1480
rect 59150 1445 59155 1475
rect 59185 1445 59190 1475
rect 59150 1440 59190 1445
rect 58055 1050 58060 1080
rect 58090 1050 58100 1080
rect 58130 1050 58140 1080
rect 58170 1050 58175 1080
rect 58055 1040 58175 1050
rect 58055 1010 58060 1040
rect 58090 1010 58100 1040
rect 58130 1010 58140 1040
rect 58170 1010 58175 1040
rect 58055 1000 58175 1010
rect 58055 970 58060 1000
rect 58090 970 58100 1000
rect 58130 970 58140 1000
rect 58170 970 58175 1000
rect 58055 965 58175 970
rect 58405 1425 58435 1435
rect 58405 1155 58410 1425
rect 58430 1155 58435 1425
rect 58405 1115 58435 1155
rect 58405 1095 58410 1115
rect 58430 1095 58435 1115
rect 58405 945 58435 1095
rect 58460 1425 58490 1435
rect 58460 1155 58465 1425
rect 58485 1155 58490 1425
rect 58460 1085 58490 1155
rect 58515 1425 58545 1440
rect 58515 1155 58520 1425
rect 58540 1155 58545 1425
rect 58515 1140 58545 1155
rect 58570 1425 58600 1435
rect 58570 1155 58575 1425
rect 58595 1155 58600 1425
rect 58510 1135 58550 1140
rect 58510 1105 58515 1135
rect 58545 1105 58550 1135
rect 58510 1100 58550 1105
rect 58570 1085 58600 1155
rect 58625 1425 58655 1440
rect 58625 1155 58630 1425
rect 58650 1155 58655 1425
rect 58625 1140 58655 1155
rect 58680 1425 58710 1435
rect 58680 1155 58685 1425
rect 58705 1155 58710 1425
rect 58620 1135 58660 1140
rect 58620 1105 58625 1135
rect 58655 1105 58660 1135
rect 58620 1100 58660 1105
rect 58680 1085 58710 1155
rect 58735 1425 58765 1440
rect 58735 1155 58740 1425
rect 58760 1155 58765 1425
rect 58735 1140 58765 1155
rect 58790 1425 58820 1435
rect 58790 1155 58795 1425
rect 58815 1155 58820 1425
rect 58730 1135 58770 1140
rect 58730 1105 58735 1135
rect 58765 1105 58770 1135
rect 58730 1100 58770 1105
rect 58790 1085 58820 1155
rect 58845 1425 58875 1440
rect 58845 1155 58850 1425
rect 58870 1155 58875 1425
rect 58845 1140 58875 1155
rect 58900 1425 58930 1435
rect 58900 1155 58905 1425
rect 58925 1155 58930 1425
rect 58840 1135 58880 1140
rect 58840 1105 58845 1135
rect 58875 1105 58880 1135
rect 58840 1100 58880 1105
rect 58900 1085 58930 1155
rect 58955 1425 58985 1440
rect 58955 1155 58960 1425
rect 58980 1155 58985 1425
rect 58955 1140 58985 1155
rect 59010 1425 59040 1435
rect 59010 1155 59015 1425
rect 59035 1155 59040 1425
rect 58950 1135 58990 1140
rect 58950 1105 58955 1135
rect 58985 1105 58990 1135
rect 58950 1100 58990 1105
rect 59010 1085 59040 1155
rect 59065 1425 59095 1435
rect 59065 1155 59070 1425
rect 59090 1155 59095 1425
rect 59160 1160 59180 1440
rect 59065 1115 59095 1155
rect 59150 1155 59190 1160
rect 59150 1125 59155 1155
rect 59185 1125 59190 1155
rect 59150 1120 59190 1125
rect 59065 1095 59070 1115
rect 59090 1095 59095 1115
rect 58455 1080 58495 1085
rect 58455 1050 58460 1080
rect 58490 1050 58495 1080
rect 58455 1040 58495 1050
rect 58455 1010 58460 1040
rect 58490 1010 58495 1040
rect 58455 1000 58495 1010
rect 58455 970 58460 1000
rect 58490 970 58495 1000
rect 58455 965 58495 970
rect 58565 1080 58605 1085
rect 58565 1050 58570 1080
rect 58600 1050 58605 1080
rect 58565 1040 58605 1050
rect 58565 1010 58570 1040
rect 58600 1010 58605 1040
rect 58565 1000 58605 1010
rect 58565 970 58570 1000
rect 58600 970 58605 1000
rect 58565 965 58605 970
rect 58675 1080 58715 1085
rect 58675 1050 58680 1080
rect 58710 1050 58715 1080
rect 58675 1040 58715 1050
rect 58675 1010 58680 1040
rect 58710 1010 58715 1040
rect 58675 1000 58715 1010
rect 58675 970 58680 1000
rect 58710 970 58715 1000
rect 58675 965 58715 970
rect 58785 1080 58825 1085
rect 58785 1050 58790 1080
rect 58820 1050 58825 1080
rect 58785 1040 58825 1050
rect 58785 1010 58790 1040
rect 58820 1010 58825 1040
rect 58785 1000 58825 1010
rect 58785 970 58790 1000
rect 58820 970 58825 1000
rect 58785 965 58825 970
rect 58895 1080 58935 1085
rect 58895 1050 58900 1080
rect 58930 1050 58935 1080
rect 58895 1040 58935 1050
rect 58895 1010 58900 1040
rect 58930 1010 58935 1040
rect 58895 1000 58935 1010
rect 58895 970 58900 1000
rect 58930 970 58935 1000
rect 58895 965 58935 970
rect 59005 1080 59045 1085
rect 59005 1050 59010 1080
rect 59040 1050 59045 1080
rect 59005 1040 59045 1050
rect 59005 1010 59010 1040
rect 59040 1010 59045 1040
rect 59005 1000 59045 1010
rect 59005 970 59010 1000
rect 59040 970 59045 1000
rect 59005 965 59045 970
rect 59065 945 59095 1095
rect 59205 1090 59225 1625
rect 59480 1610 59730 1630
rect 59480 1580 59490 1610
rect 59520 1580 59540 1610
rect 59570 1580 59590 1610
rect 59620 1580 59640 1610
rect 59670 1580 59690 1610
rect 59720 1580 59730 1610
rect 59250 1160 59285 1165
rect 59250 1120 59285 1125
rect 59310 1160 59345 1165
rect 59310 1120 59345 1125
rect 59370 1160 59405 1165
rect 59370 1120 59405 1125
rect 59430 1160 59465 1166
rect 59430 1120 59465 1125
rect 59315 1090 59335 1120
rect 59195 1085 59235 1090
rect 59195 1055 59200 1085
rect 59230 1055 59235 1085
rect 59195 1050 59235 1055
rect 59305 1085 59345 1090
rect 59305 1055 59310 1085
rect 59340 1055 59345 1085
rect 59305 1050 59345 1055
rect 58400 940 58440 945
rect 58400 910 58405 940
rect 58435 910 58440 940
rect 58400 900 58440 910
rect 58400 870 58405 900
rect 58435 870 58440 900
rect 58400 860 58440 870
rect 58400 830 58405 860
rect 58435 830 58440 860
rect 58400 825 58440 830
rect 59060 940 59100 945
rect 59060 910 59065 940
rect 59095 910 59100 940
rect 59060 900 59100 910
rect 59060 870 59065 900
rect 59095 870 59100 900
rect 59060 860 59100 870
rect 59060 830 59065 860
rect 59095 830 59100 860
rect 59060 825 59100 830
rect 59435 810 59455 1120
rect 59425 805 59465 810
rect 59425 775 59430 805
rect 59460 775 59465 805
rect 59425 770 59465 775
rect 58680 435 58720 440
rect 58680 405 58685 435
rect 58715 405 58720 435
rect 58680 400 58720 405
rect 59360 435 59400 440
rect 59360 405 59365 435
rect 59395 405 59400 435
rect 59360 400 59400 405
rect 58530 310 58970 315
rect 58530 280 58535 310
rect 58565 280 58575 310
rect 58605 280 58615 310
rect 58645 280 58655 310
rect 58685 280 58695 310
rect 58725 280 58735 310
rect 58765 280 58775 310
rect 58805 280 58815 310
rect 58845 280 58855 310
rect 58885 280 58895 310
rect 58925 280 58935 310
rect 58965 280 58970 310
rect 58530 270 58970 280
rect 58530 240 58535 270
rect 58565 240 58575 270
rect 58605 240 58615 270
rect 58645 240 58655 270
rect 58685 240 58695 270
rect 58725 240 58735 270
rect 58765 240 58775 270
rect 58805 240 58815 270
rect 58845 240 58855 270
rect 58885 240 58895 270
rect 58925 240 58935 270
rect 58965 240 58970 270
rect 58530 230 58970 240
rect 58530 200 58535 230
rect 58565 200 58575 230
rect 58605 200 58615 230
rect 58645 200 58655 230
rect 58685 200 58695 230
rect 58725 200 58735 230
rect 58765 200 58775 230
rect 58805 200 58815 230
rect 58845 200 58855 230
rect 58885 200 58895 230
rect 58925 200 58935 230
rect 58965 200 58970 230
rect 58530 195 58970 200
rect 59295 310 59335 315
rect 59295 280 59300 310
rect 59330 280 59335 310
rect 59295 270 59335 280
rect 59295 240 59300 270
rect 59330 240 59335 270
rect 59295 230 59335 240
rect 59295 200 59300 230
rect 59330 200 59335 230
rect 59295 195 59335 200
rect 57920 -125 57925 -95
rect 57955 -125 57965 -95
rect 57995 -125 58005 -95
rect 58035 -125 58040 -95
rect 57920 -135 58040 -125
rect 57920 -165 57925 -135
rect 57955 -165 57965 -135
rect 57995 -165 58005 -135
rect 58035 -165 58040 -135
rect 57920 -175 58040 -165
rect 57920 -205 57925 -175
rect 57955 -205 57965 -175
rect 57995 -205 58005 -175
rect 58035 -205 58040 -175
rect 57920 -210 58040 -205
rect 58435 165 58465 175
rect 58435 -505 58440 165
rect 58460 -505 58465 165
rect 58435 -545 58465 -505
rect 58535 165 58565 195
rect 58535 -505 58540 165
rect 58560 -505 58565 165
rect 58535 -520 58565 -505
rect 58635 165 58665 175
rect 58635 -505 58640 165
rect 58660 -505 58665 165
rect 58435 -565 58440 -545
rect 58460 -565 58465 -545
rect 58530 -525 58570 -520
rect 58530 -555 58535 -525
rect 58565 -555 58570 -525
rect 58530 -560 58570 -555
rect 58435 -575 58465 -565
rect 58635 -575 58665 -505
rect 58735 165 58765 195
rect 58735 -505 58740 165
rect 58760 -505 58765 165
rect 58735 -520 58765 -505
rect 58835 165 58865 175
rect 58835 -505 58840 165
rect 58860 -505 58865 165
rect 58730 -525 58770 -520
rect 58730 -555 58735 -525
rect 58765 -555 58770 -525
rect 58730 -560 58770 -555
rect 58835 -575 58865 -505
rect 58935 165 58965 195
rect 59300 175 59335 195
rect 59370 180 59390 400
rect 59480 310 59730 1580
rect 59480 280 59485 310
rect 59515 280 59525 310
rect 59555 280 59570 310
rect 59600 280 59610 310
rect 59640 280 59655 310
rect 59685 280 59695 310
rect 59725 280 59730 310
rect 59480 270 59730 280
rect 59480 240 59485 270
rect 59515 240 59525 270
rect 59555 240 59570 270
rect 59600 240 59610 270
rect 59640 240 59655 270
rect 59685 240 59695 270
rect 59725 240 59730 270
rect 59480 230 59730 240
rect 59480 200 59485 230
rect 59515 200 59525 230
rect 59555 200 59570 230
rect 59600 200 59610 230
rect 59640 200 59655 230
rect 59685 200 59695 230
rect 59725 200 59730 230
rect 59480 195 59730 200
rect 59760 2050 59880 2055
rect 59760 2020 59765 2050
rect 59795 2020 59805 2050
rect 59835 2020 59845 2050
rect 59875 2020 59880 2050
rect 59760 2010 59880 2020
rect 59760 1980 59765 2010
rect 59795 1980 59805 2010
rect 59835 1980 59845 2010
rect 59875 1980 59880 2010
rect 59760 1970 59880 1980
rect 59760 1940 59765 1970
rect 59795 1940 59805 1970
rect 59835 1940 59845 1970
rect 59875 1940 59880 1970
rect 59760 940 59880 1940
rect 59760 910 59765 940
rect 59795 910 59805 940
rect 59835 910 59845 940
rect 59875 910 59880 940
rect 59760 900 59880 910
rect 59760 870 59765 900
rect 59795 870 59805 900
rect 59835 870 59845 900
rect 59875 870 59880 900
rect 59760 860 59880 870
rect 59760 830 59765 860
rect 59795 830 59805 860
rect 59835 830 59845 860
rect 59875 830 59880 860
rect 58935 -505 58940 165
rect 58960 -505 58965 165
rect 58935 -520 58965 -505
rect 59035 165 59065 175
rect 59035 -505 59040 165
rect 59060 -505 59065 165
rect 59300 135 59335 140
rect 59360 175 59395 180
rect 59360 135 59395 140
rect 58930 -525 58970 -520
rect 58930 -555 58935 -525
rect 58965 -555 58970 -525
rect 58930 -560 58970 -555
rect 59035 -545 59065 -505
rect 59035 -565 59040 -545
rect 59060 -565 59065 -545
rect 59035 -575 59065 -565
rect 59760 -575 59880 830
rect 57485 -610 57490 -580
rect 57520 -610 57525 -580
rect 57485 -620 57525 -610
rect 57485 -650 57490 -620
rect 57520 -650 57525 -620
rect 57485 -660 57525 -650
rect 57485 -690 57490 -660
rect 57520 -690 57525 -660
rect 57485 -695 57525 -690
rect 57540 -580 57660 -575
rect 57540 -610 57545 -580
rect 57575 -610 57585 -580
rect 57615 -610 57625 -580
rect 57655 -610 57660 -580
rect 57540 -620 57660 -610
rect 57540 -650 57545 -620
rect 57575 -650 57585 -620
rect 57615 -650 57625 -620
rect 57655 -650 57660 -620
rect 57540 -660 57660 -650
rect 57540 -690 57545 -660
rect 57575 -690 57585 -660
rect 57615 -690 57625 -660
rect 57655 -690 57660 -660
rect 57540 -1500 57660 -690
rect 57890 -580 58010 -575
rect 57890 -610 57895 -580
rect 57925 -610 57935 -580
rect 57965 -610 57975 -580
rect 58005 -610 58010 -580
rect 57890 -620 58010 -610
rect 57890 -650 57895 -620
rect 57925 -650 57935 -620
rect 57965 -650 57975 -620
rect 58005 -650 58010 -620
rect 57890 -660 58010 -650
rect 57890 -690 57895 -660
rect 57925 -690 57935 -660
rect 57965 -690 57975 -660
rect 58005 -690 58010 -660
rect 57890 -1500 58010 -690
rect 58240 -580 58480 -575
rect 58240 -610 58245 -580
rect 58275 -610 58285 -580
rect 58315 -610 58325 -580
rect 58355 -610 58365 -580
rect 58395 -610 58405 -580
rect 58435 -610 58445 -580
rect 58475 -610 58480 -580
rect 58240 -620 58480 -610
rect 58240 -650 58245 -620
rect 58275 -650 58285 -620
rect 58315 -650 58325 -620
rect 58355 -650 58365 -620
rect 58395 -650 58405 -620
rect 58435 -650 58445 -620
rect 58475 -650 58480 -620
rect 58240 -660 58480 -650
rect 58240 -690 58245 -660
rect 58275 -690 58285 -660
rect 58315 -690 58325 -660
rect 58355 -690 58365 -660
rect 58395 -690 58405 -660
rect 58435 -690 58445 -660
rect 58475 -690 58480 -660
rect 58240 -695 58480 -690
rect 58590 -580 58710 -575
rect 58590 -610 58595 -580
rect 58625 -610 58635 -580
rect 58665 -610 58675 -580
rect 58705 -610 58710 -580
rect 58590 -620 58710 -610
rect 58590 -650 58595 -620
rect 58625 -650 58635 -620
rect 58665 -650 58675 -620
rect 58705 -650 58710 -620
rect 58590 -660 58710 -650
rect 58590 -690 58595 -660
rect 58625 -690 58635 -660
rect 58665 -690 58675 -660
rect 58705 -690 58710 -660
rect 58240 -1500 58360 -695
rect 58590 -1500 58710 -690
rect 58830 -580 58870 -575
rect 58830 -610 58835 -580
rect 58865 -610 58870 -580
rect 58830 -620 58870 -610
rect 58830 -650 58835 -620
rect 58865 -650 58870 -620
rect 58830 -660 58870 -650
rect 58830 -690 58835 -660
rect 58865 -690 58870 -660
rect 58830 -695 58870 -690
rect 58940 -580 59065 -575
rect 58940 -610 58945 -580
rect 58975 -610 58985 -580
rect 59015 -610 59025 -580
rect 59055 -610 59065 -580
rect 58940 -620 59065 -610
rect 58940 -650 58945 -620
rect 58975 -650 58985 -620
rect 59015 -650 59025 -620
rect 59055 -650 59065 -620
rect 58940 -660 59065 -650
rect 58940 -690 58945 -660
rect 58975 -690 58985 -660
rect 59015 -690 59025 -660
rect 59055 -690 59065 -660
rect 58940 -695 59065 -690
rect 59290 -580 59410 -575
rect 59290 -610 59295 -580
rect 59325 -610 59335 -580
rect 59365 -610 59375 -580
rect 59405 -610 59410 -580
rect 59290 -620 59410 -610
rect 59290 -650 59295 -620
rect 59325 -650 59335 -620
rect 59365 -650 59375 -620
rect 59405 -650 59410 -620
rect 59290 -660 59410 -650
rect 59290 -690 59295 -660
rect 59325 -690 59335 -660
rect 59365 -690 59375 -660
rect 59405 -690 59410 -660
rect 58940 -1500 59060 -695
rect 59290 -1500 59410 -690
rect 59640 -580 59880 -575
rect 59640 -610 59645 -580
rect 59675 -610 59685 -580
rect 59715 -610 59725 -580
rect 59755 -610 59765 -580
rect 59795 -610 59805 -580
rect 59835 -610 59845 -580
rect 59875 -610 59880 -580
rect 59640 -620 59880 -610
rect 59640 -650 59645 -620
rect 59675 -650 59685 -620
rect 59715 -650 59725 -620
rect 59755 -650 59765 -620
rect 59795 -650 59805 -620
rect 59835 -650 59845 -620
rect 59875 -650 59880 -620
rect 59640 -660 59880 -650
rect 59640 -690 59645 -660
rect 59675 -690 59685 -660
rect 59715 -690 59725 -660
rect 59755 -690 59765 -660
rect 59795 -690 59805 -660
rect 59835 -690 59845 -660
rect 59875 -690 59880 -660
rect 59640 -695 59880 -690
rect 59990 -580 60110 -575
rect 59990 -610 59995 -580
rect 60025 -610 60035 -580
rect 60065 -610 60075 -580
rect 60105 -610 60110 -580
rect 59990 -620 60110 -610
rect 59990 -650 59995 -620
rect 60025 -650 60035 -620
rect 60065 -650 60075 -620
rect 60105 -650 60110 -620
rect 59990 -660 60110 -650
rect 59990 -690 59995 -660
rect 60025 -690 60035 -660
rect 60065 -690 60075 -660
rect 60105 -690 60110 -660
rect 59640 -1500 59760 -695
rect 59990 -1500 60110 -690
rect 60340 -580 60460 -575
rect 60340 -610 60345 -580
rect 60375 -610 60385 -580
rect 60415 -610 60425 -580
rect 60455 -610 60460 -580
rect 60340 -620 60460 -610
rect 60340 -650 60345 -620
rect 60375 -650 60385 -620
rect 60415 -650 60425 -620
rect 60455 -650 60460 -620
rect 60340 -660 60460 -650
rect 60340 -690 60345 -660
rect 60375 -690 60385 -660
rect 60415 -690 60425 -660
rect 60455 -690 60460 -660
rect 60340 -1500 60460 -690
rect 60690 -580 60810 -575
rect 60690 -610 60695 -580
rect 60725 -610 60735 -580
rect 60765 -610 60775 -580
rect 60805 -610 60810 -580
rect 60690 -620 60810 -610
rect 60690 -650 60695 -620
rect 60725 -650 60735 -620
rect 60765 -650 60775 -620
rect 60805 -650 60810 -620
rect 60690 -660 60810 -650
rect 60690 -690 60695 -660
rect 60725 -690 60735 -660
rect 60765 -690 60775 -660
rect 60805 -690 60810 -660
rect 60690 -1500 60810 -690
rect 61040 -580 61160 -575
rect 61040 -610 61045 -580
rect 61075 -610 61085 -580
rect 61115 -610 61125 -580
rect 61155 -610 61160 -580
rect 61040 -620 61160 -610
rect 61040 -650 61045 -620
rect 61075 -650 61085 -620
rect 61115 -650 61125 -620
rect 61155 -650 61160 -620
rect 61040 -660 61160 -650
rect 61040 -690 61045 -660
rect 61075 -690 61085 -660
rect 61115 -690 61125 -660
rect 61155 -690 61160 -660
rect 61040 -1500 61160 -690
rect 61390 -580 61510 -575
rect 61390 -610 61395 -580
rect 61425 -610 61435 -580
rect 61465 -610 61475 -580
rect 61505 -610 61510 -580
rect 61390 -620 61510 -610
rect 61390 -650 61395 -620
rect 61425 -650 61435 -620
rect 61465 -650 61475 -620
rect 61505 -650 61510 -620
rect 61390 -660 61510 -650
rect 61390 -690 61395 -660
rect 61425 -690 61435 -660
rect 61465 -690 61475 -660
rect 61505 -690 61510 -660
rect 61390 -1500 61510 -690
<< via1 >>
rect 52295 4290 52325 4320
rect 52335 4290 52365 4320
rect 52375 4290 52405 4320
rect 52295 4250 52325 4280
rect 52335 4250 52365 4280
rect 52375 4250 52405 4280
rect 52295 4210 52325 4240
rect 52335 4210 52365 4240
rect 52375 4210 52405 4240
rect 52645 4290 52675 4320
rect 52685 4290 52715 4320
rect 52725 4290 52755 4320
rect 52645 4250 52675 4280
rect 52685 4250 52715 4280
rect 52725 4250 52755 4280
rect 52645 4210 52675 4240
rect 52685 4210 52715 4240
rect 52725 4210 52755 4240
rect 52995 4290 53025 4320
rect 53035 4290 53065 4320
rect 53075 4290 53105 4320
rect 52995 4250 53025 4280
rect 53035 4250 53065 4280
rect 53075 4250 53105 4280
rect 52995 4210 53025 4240
rect 53035 4210 53065 4240
rect 53075 4210 53105 4240
rect 53695 4290 53725 4320
rect 53735 4290 53765 4320
rect 53775 4290 53805 4320
rect 53695 4250 53725 4280
rect 53735 4250 53765 4280
rect 53775 4250 53805 4280
rect 53695 4210 53725 4240
rect 53735 4210 53765 4240
rect 53775 4210 53805 4240
rect 56210 5035 56240 5065
rect 56090 4925 56120 4930
rect 56090 4905 56095 4925
rect 56095 4905 56115 4925
rect 56115 4905 56120 4925
rect 56090 4900 56120 4905
rect 56680 5035 56710 5065
rect 57090 5035 57120 5065
rect 57560 5035 57590 5065
rect 56210 4900 56240 4930
rect 56270 4925 56300 4930
rect 56270 4905 56275 4925
rect 56275 4905 56295 4925
rect 56295 4905 56300 4925
rect 56270 4900 56300 4905
rect 56560 4810 56590 4840
rect 56560 4770 56590 4800
rect 56560 4755 56590 4760
rect 56560 4735 56565 4755
rect 56565 4735 56585 4755
rect 56585 4735 56590 4755
rect 56560 4730 56590 4735
rect 56620 4810 56650 4840
rect 56620 4770 56650 4800
rect 56620 4730 56650 4760
rect 56885 4980 56915 5010
rect 56885 4940 56915 4970
rect 56885 4900 56915 4930
rect 56740 4810 56770 4840
rect 56740 4770 56770 4800
rect 56740 4755 56770 4760
rect 56740 4735 56745 4755
rect 56745 4735 56765 4755
rect 56765 4735 56770 4755
rect 56740 4730 56770 4735
rect 57030 4980 57060 5010
rect 57030 4940 57060 4970
rect 57030 4925 57060 4930
rect 57030 4905 57035 4925
rect 57035 4905 57055 4925
rect 57055 4905 57060 4925
rect 57030 4900 57060 4905
rect 56885 4810 56915 4840
rect 56885 4770 56915 4800
rect 56885 4730 56915 4760
rect 56210 4495 56240 4525
rect 56680 4495 56710 4525
rect 56155 4475 56185 4480
rect 56155 4455 56160 4475
rect 56160 4455 56180 4475
rect 56180 4455 56185 4475
rect 56155 4450 56185 4455
rect 56630 4475 56660 4480
rect 56630 4455 56635 4475
rect 56635 4455 56655 4475
rect 56655 4455 56660 4475
rect 56630 4450 56660 4455
rect 56830 4450 56860 4480
rect 54045 4290 54075 4320
rect 54085 4290 54115 4320
rect 54125 4290 54155 4320
rect 54045 4250 54075 4280
rect 54085 4250 54115 4280
rect 54125 4250 54155 4280
rect 54045 4210 54075 4240
rect 54085 4210 54115 4240
rect 54125 4210 54155 4240
rect 54675 4290 54705 4320
rect 54675 4250 54705 4280
rect 54675 4210 54705 4240
rect 55035 4290 55065 4320
rect 55035 4250 55065 4280
rect 55035 4210 55065 4240
rect 54735 4155 54765 4185
rect 54775 4155 54805 4185
rect 54815 4155 54845 4185
rect 54855 4155 54885 4185
rect 54895 4155 54925 4185
rect 54935 4155 54965 4185
rect 54975 4155 55005 4185
rect 54735 4115 54765 4145
rect 54775 4115 54805 4145
rect 54815 4115 54845 4145
rect 54855 4115 54885 4145
rect 54895 4115 54925 4145
rect 54935 4115 54965 4145
rect 54975 4115 55005 4145
rect 54735 4075 54765 4105
rect 54775 4075 54805 4105
rect 54815 4075 54845 4105
rect 54855 4075 54885 4105
rect 54895 4075 54925 4105
rect 54935 4075 54965 4105
rect 54975 4075 55005 4105
rect 54675 4020 54705 4050
rect 54795 4020 54825 4050
rect 54915 4020 54945 4050
rect 55395 4290 55425 4320
rect 55395 4250 55425 4280
rect 55395 4210 55425 4240
rect 55095 4155 55125 4185
rect 55135 4155 55165 4185
rect 55175 4155 55205 4185
rect 55215 4155 55245 4185
rect 55255 4155 55285 4185
rect 55295 4155 55325 4185
rect 55335 4155 55365 4185
rect 55095 4115 55125 4145
rect 55135 4115 55165 4145
rect 55175 4115 55205 4145
rect 55215 4115 55245 4145
rect 55255 4115 55285 4145
rect 55295 4115 55325 4145
rect 55335 4115 55365 4145
rect 55095 4075 55125 4105
rect 55135 4075 55165 4105
rect 55175 4075 55205 4105
rect 55215 4075 55245 4105
rect 55255 4075 55285 4105
rect 55295 4075 55325 4105
rect 55335 4075 55365 4105
rect 55035 4020 55065 4050
rect 55155 4020 55185 4050
rect 55275 4020 55305 4050
rect 55395 4020 55425 4050
rect 55625 4290 55655 4320
rect 55665 4290 55695 4320
rect 55705 4290 55735 4320
rect 55625 4250 55655 4280
rect 55665 4250 55695 4280
rect 55705 4250 55735 4280
rect 55625 4210 55655 4240
rect 55665 4210 55695 4240
rect 55705 4210 55735 4240
rect 54735 3630 54765 3660
rect 54855 3630 54885 3660
rect 54975 3630 55005 3660
rect 55095 3630 55125 3660
rect 55215 3630 55245 3660
rect 55335 3630 55365 3660
rect 55035 3530 55065 3535
rect 55035 3510 55040 3530
rect 55040 3510 55060 3530
rect 55060 3510 55065 3530
rect 55035 3505 55065 3510
rect 55485 3460 55515 3490
rect 55525 3460 55555 3490
rect 55565 3460 55595 3490
rect 55485 3420 55515 3450
rect 55525 3420 55555 3450
rect 55565 3420 55595 3450
rect 55485 3380 55515 3410
rect 55525 3380 55555 3410
rect 55565 3380 55595 3410
rect 54260 3345 54290 3375
rect 54705 3325 54735 3355
rect 54705 3285 54735 3315
rect 54705 3245 54735 3275
rect 54815 3325 54845 3355
rect 54815 3285 54845 3315
rect 54815 3245 54845 3275
rect 54925 3325 54955 3355
rect 54925 3285 54955 3315
rect 54925 3245 54955 3275
rect 55035 3325 55065 3355
rect 55035 3285 55065 3315
rect 55035 3245 55065 3275
rect 55145 3325 55175 3355
rect 55145 3285 55175 3315
rect 55145 3245 55175 3275
rect 55255 3325 55285 3355
rect 55255 3285 55285 3315
rect 55255 3245 55285 3275
rect 55365 3325 55395 3355
rect 55365 3285 55395 3315
rect 55365 3245 55395 3275
rect 54760 3160 54790 3190
rect 54870 3160 54900 3190
rect 54980 3160 55010 3190
rect 55090 3160 55120 3190
rect 55200 3160 55230 3190
rect 55310 3160 55340 3190
rect 54220 2440 54250 2470
rect 54260 2440 54290 2470
rect 54300 2440 54330 2470
rect 54220 2400 54250 2430
rect 54260 2400 54290 2430
rect 54300 2400 54330 2430
rect 54220 2360 54250 2390
rect 54260 2360 54290 2390
rect 54300 2360 54330 2390
rect 54760 2520 54790 2550
rect 54870 2520 54900 2550
rect 54980 2520 55010 2550
rect 55090 2520 55120 2550
rect 55035 2465 55065 2470
rect 55035 2445 55040 2465
rect 55040 2445 55060 2465
rect 55060 2445 55065 2465
rect 55035 2440 55065 2445
rect 55035 2425 55065 2430
rect 55035 2405 55040 2425
rect 55040 2405 55060 2425
rect 55060 2405 55065 2425
rect 55035 2400 55065 2405
rect 55035 2385 55065 2390
rect 55035 2365 55040 2385
rect 55040 2365 55060 2385
rect 55060 2365 55065 2385
rect 55035 2360 55065 2365
rect 55200 2520 55230 2550
rect 55310 2520 55340 2550
rect 54075 2290 54105 2320
rect 54115 2290 54145 2320
rect 54160 2290 54190 2320
rect 54200 2290 54230 2320
rect 54245 2290 54275 2320
rect 54285 2290 54315 2320
rect 54075 2250 54105 2280
rect 54115 2250 54145 2280
rect 54160 2250 54190 2280
rect 54200 2250 54230 2280
rect 54245 2250 54275 2280
rect 54285 2250 54315 2280
rect 54075 2210 54105 2240
rect 54115 2210 54145 2240
rect 54160 2210 54190 2240
rect 54200 2210 54230 2240
rect 54245 2210 54275 2240
rect 54285 2210 54315 2240
rect 53925 2020 53955 2050
rect 53965 2020 53995 2050
rect 54005 2020 54035 2050
rect 53925 1980 53955 2010
rect 53965 1980 53995 2010
rect 54005 1980 54035 2010
rect 53925 1940 53955 1970
rect 53965 1940 53995 1970
rect 54005 1940 54035 1970
rect 53925 910 53955 940
rect 53965 910 53995 940
rect 54005 910 54035 940
rect 53925 870 53955 900
rect 53965 870 53995 900
rect 54005 870 54035 900
rect 53925 830 53955 860
rect 53965 830 53995 860
rect 54005 830 54035 860
rect 54760 2290 54790 2320
rect 54815 2290 54845 2320
rect 54870 2290 54900 2320
rect 54925 2290 54955 2320
rect 54980 2290 55010 2320
rect 55035 2290 55065 2320
rect 55090 2290 55120 2320
rect 55145 2290 55175 2320
rect 55200 2290 55230 2320
rect 55255 2290 55285 2320
rect 55310 2290 55340 2320
rect 54760 2250 54790 2280
rect 54815 2250 54845 2280
rect 54870 2250 54900 2280
rect 54925 2250 54955 2280
rect 54980 2250 55010 2280
rect 55035 2250 55065 2280
rect 55090 2250 55120 2280
rect 55145 2250 55175 2280
rect 55200 2250 55230 2280
rect 55255 2250 55285 2280
rect 55310 2250 55340 2280
rect 54760 2210 54790 2240
rect 54815 2210 54845 2240
rect 54870 2210 54900 2240
rect 54925 2210 54955 2240
rect 54980 2210 55010 2240
rect 55035 2210 55065 2240
rect 55090 2210 55120 2240
rect 55145 2210 55175 2240
rect 55200 2210 55230 2240
rect 55255 2210 55285 2240
rect 55310 2210 55340 2240
rect 55485 2440 55515 2470
rect 55525 2440 55555 2470
rect 55565 2440 55595 2470
rect 55485 2400 55515 2430
rect 55525 2400 55555 2430
rect 55565 2400 55595 2430
rect 55485 2360 55515 2390
rect 55525 2360 55555 2390
rect 55565 2360 55595 2390
rect 54705 2155 54735 2185
rect 54705 2115 54735 2145
rect 54705 2075 54735 2105
rect 55365 2155 55395 2185
rect 55365 2115 55395 2145
rect 55365 2075 55395 2105
rect 54080 1680 54110 1710
rect 54130 1680 54160 1710
rect 54180 1680 54210 1710
rect 54230 1680 54260 1710
rect 54280 1680 54310 1710
rect 54760 2020 54790 2050
rect 54760 1980 54790 2010
rect 54760 1940 54790 1970
rect 54870 2020 54900 2050
rect 54870 1980 54900 2010
rect 54870 1940 54900 1970
rect 54980 2020 55010 2050
rect 54980 1980 55010 2010
rect 54980 1940 55010 1970
rect 55090 2020 55120 2050
rect 55090 1980 55120 2010
rect 55090 1940 55120 1970
rect 55200 2020 55230 2050
rect 55200 1980 55230 2010
rect 55200 1940 55230 1970
rect 55310 2020 55340 2050
rect 55310 1980 55340 2010
rect 55310 1940 55340 1970
rect 54815 1885 54845 1915
rect 54925 1885 54955 1915
rect 55035 1885 55065 1915
rect 55145 1885 55175 1915
rect 55255 1885 55285 1915
rect 54080 1630 54110 1660
rect 54130 1630 54160 1660
rect 54180 1630 54210 1660
rect 54230 1630 54260 1660
rect 54280 1630 54310 1660
rect 54570 1630 54600 1660
rect 54815 1655 54845 1660
rect 54815 1635 54820 1655
rect 54820 1635 54840 1655
rect 54840 1635 54845 1655
rect 54815 1630 54845 1635
rect 54925 1655 54955 1660
rect 54925 1635 54930 1655
rect 54930 1635 54950 1655
rect 54950 1635 54955 1655
rect 54925 1630 54955 1635
rect 55035 1655 55065 1660
rect 55035 1635 55040 1655
rect 55040 1635 55060 1655
rect 55060 1635 55065 1655
rect 55035 1630 55065 1635
rect 55145 1655 55175 1660
rect 55145 1635 55150 1655
rect 55150 1635 55170 1655
rect 55170 1635 55175 1655
rect 55145 1630 55175 1635
rect 55255 1655 55285 1660
rect 55255 1635 55260 1655
rect 55260 1635 55280 1655
rect 55280 1635 55285 1655
rect 55255 1630 55285 1635
rect 54080 1580 54110 1610
rect 54130 1580 54160 1610
rect 54180 1580 54210 1610
rect 54230 1580 54260 1610
rect 54280 1580 54310 1610
rect 54335 1155 54370 1160
rect 54335 1130 54340 1155
rect 54340 1130 54365 1155
rect 54365 1130 54370 1155
rect 54335 1125 54370 1130
rect 54395 1155 54430 1160
rect 54395 1130 54400 1155
rect 54400 1130 54425 1155
rect 54425 1130 54430 1155
rect 54395 1125 54430 1130
rect 54455 1155 54490 1160
rect 54455 1130 54460 1155
rect 54460 1130 54485 1155
rect 54485 1130 54490 1155
rect 54455 1125 54490 1130
rect 54515 1155 54550 1160
rect 54515 1130 54520 1155
rect 54520 1130 54545 1155
rect 54545 1130 54550 1155
rect 54515 1125 54550 1130
rect 55200 1590 55230 1595
rect 55200 1570 55205 1590
rect 55205 1570 55225 1590
rect 55225 1570 55230 1590
rect 55200 1565 55230 1570
rect 55200 1550 55230 1555
rect 55200 1530 55205 1550
rect 55205 1530 55225 1550
rect 55225 1530 55230 1550
rect 55200 1525 55230 1530
rect 55485 1565 55515 1595
rect 55525 1565 55555 1595
rect 55565 1565 55595 1595
rect 55485 1525 55515 1555
rect 55525 1525 55555 1555
rect 55565 1525 55595 1555
rect 56010 4155 56040 4185
rect 56050 4155 56080 4185
rect 56090 4155 56120 4185
rect 56130 4155 56160 4185
rect 56170 4155 56200 4185
rect 56210 4155 56240 4185
rect 56250 4155 56280 4185
rect 56290 4155 56320 4185
rect 56330 4155 56360 4185
rect 56370 4155 56400 4185
rect 56410 4155 56440 4185
rect 56450 4155 56480 4185
rect 56490 4155 56520 4185
rect 56530 4155 56560 4185
rect 56570 4155 56600 4185
rect 56610 4155 56640 4185
rect 56650 4155 56680 4185
rect 56690 4155 56720 4185
rect 56730 4155 56760 4185
rect 56010 4115 56040 4145
rect 56050 4115 56080 4145
rect 56090 4115 56120 4145
rect 56130 4115 56160 4145
rect 56170 4115 56200 4145
rect 56210 4115 56240 4145
rect 56250 4115 56280 4145
rect 56290 4115 56320 4145
rect 56330 4115 56360 4145
rect 56370 4115 56400 4145
rect 56410 4115 56440 4145
rect 56450 4115 56480 4145
rect 56490 4115 56520 4145
rect 56530 4115 56560 4145
rect 56570 4115 56600 4145
rect 56610 4115 56640 4145
rect 56650 4115 56680 4145
rect 56690 4115 56720 4145
rect 56730 4115 56760 4145
rect 56010 4075 56040 4105
rect 56050 4075 56080 4105
rect 56090 4075 56120 4105
rect 56130 4075 56160 4105
rect 56170 4075 56200 4105
rect 56210 4075 56240 4105
rect 56250 4075 56280 4105
rect 56290 4075 56320 4105
rect 56330 4075 56360 4105
rect 56370 4075 56400 4105
rect 56410 4075 56440 4105
rect 56450 4075 56480 4105
rect 56490 4075 56520 4105
rect 56530 4075 56560 4105
rect 56570 4075 56600 4105
rect 56610 4075 56640 4105
rect 56650 4075 56680 4105
rect 56690 4075 56720 4105
rect 56730 4075 56760 4105
rect 56070 4020 56100 4050
rect 56190 4020 56220 4050
rect 56310 4020 56340 4050
rect 56430 4020 56460 4050
rect 56550 4020 56580 4050
rect 56670 4020 56700 4050
rect 56070 3630 56100 3660
rect 56190 3630 56220 3660
rect 56310 3630 56340 3660
rect 56430 3630 56460 3660
rect 56370 3575 56400 3580
rect 56370 3555 56375 3575
rect 56375 3555 56395 3575
rect 56395 3555 56400 3575
rect 56370 3550 56400 3555
rect 56550 3630 56580 3660
rect 56670 3630 56700 3660
rect 57150 4980 57180 5010
rect 57150 4940 57180 4970
rect 57150 4900 57180 4930
rect 57210 4980 57240 5010
rect 57210 4940 57240 4970
rect 57210 4925 57240 4930
rect 57210 4905 57215 4925
rect 57215 4905 57235 4925
rect 57235 4905 57240 4925
rect 57210 4900 57240 4905
rect 57500 4925 57530 4930
rect 57500 4905 57505 4925
rect 57505 4905 57525 4925
rect 57525 4905 57530 4925
rect 57500 4900 57530 4905
rect 57560 4900 57590 4930
rect 57680 4925 57710 4930
rect 57680 4905 57685 4925
rect 57685 4905 57705 4925
rect 57705 4905 57710 4925
rect 57680 4900 57710 4905
rect 57090 4495 57120 4525
rect 57560 4495 57590 4525
rect 56885 4290 56915 4320
rect 56885 4250 56915 4280
rect 56885 4210 56915 4240
rect 56940 4395 56970 4425
rect 57576 4465 57606 4470
rect 57576 4445 57581 4465
rect 57581 4445 57601 4465
rect 57601 4445 57606 4465
rect 57576 4440 57606 4445
rect 56840 3550 56870 3580
rect 57140 4385 57170 4415
rect 57620 4385 57650 4415
rect 58060 4290 58090 4320
rect 58100 4290 58130 4320
rect 58140 4290 58170 4320
rect 58060 4250 58090 4280
rect 58100 4250 58130 4280
rect 58140 4250 58170 4280
rect 58060 4210 58090 4240
rect 58100 4210 58130 4240
rect 58140 4210 58170 4240
rect 57040 4155 57070 4185
rect 57080 4155 57110 4185
rect 57120 4155 57150 4185
rect 57160 4155 57190 4185
rect 57200 4155 57230 4185
rect 57240 4155 57270 4185
rect 57280 4155 57310 4185
rect 57320 4155 57350 4185
rect 57360 4155 57390 4185
rect 57400 4155 57430 4185
rect 57440 4155 57470 4185
rect 57480 4155 57510 4185
rect 57520 4155 57550 4185
rect 57560 4155 57590 4185
rect 57600 4155 57630 4185
rect 57640 4155 57670 4185
rect 57680 4155 57710 4185
rect 57720 4155 57750 4185
rect 57760 4155 57790 4185
rect 57040 4115 57070 4145
rect 57080 4115 57110 4145
rect 57120 4115 57150 4145
rect 57160 4115 57190 4145
rect 57200 4115 57230 4145
rect 57240 4115 57270 4145
rect 57280 4115 57310 4145
rect 57320 4115 57350 4145
rect 57360 4115 57390 4145
rect 57400 4115 57430 4145
rect 57440 4115 57470 4145
rect 57480 4115 57510 4145
rect 57520 4115 57550 4145
rect 57560 4115 57590 4145
rect 57600 4115 57630 4145
rect 57640 4115 57670 4145
rect 57680 4115 57710 4145
rect 57720 4115 57750 4145
rect 57760 4115 57790 4145
rect 57040 4075 57070 4105
rect 57080 4075 57110 4105
rect 57120 4075 57150 4105
rect 57160 4075 57190 4105
rect 57200 4075 57230 4105
rect 57240 4075 57270 4105
rect 57280 4075 57310 4105
rect 57320 4075 57350 4105
rect 57360 4075 57390 4105
rect 57400 4075 57430 4105
rect 57440 4075 57470 4105
rect 57480 4075 57510 4105
rect 57520 4075 57550 4105
rect 57560 4075 57590 4105
rect 57600 4075 57630 4105
rect 57640 4075 57670 4105
rect 57680 4075 57710 4105
rect 57720 4075 57750 4105
rect 57760 4075 57790 4105
rect 57100 4020 57130 4050
rect 57220 4020 57250 4050
rect 57340 4020 57370 4050
rect 57460 4020 57490 4050
rect 57580 4020 57610 4050
rect 57700 4020 57730 4050
rect 57100 3630 57130 3660
rect 56930 3505 56960 3535
rect 56070 3460 56100 3490
rect 56110 3460 56140 3490
rect 56150 3460 56180 3490
rect 56190 3460 56220 3490
rect 56230 3460 56260 3490
rect 56270 3460 56300 3490
rect 56310 3460 56340 3490
rect 56350 3460 56380 3490
rect 56390 3460 56420 3490
rect 56430 3460 56460 3490
rect 56470 3460 56500 3490
rect 56510 3460 56540 3490
rect 56550 3460 56580 3490
rect 56590 3460 56620 3490
rect 56630 3460 56660 3490
rect 56670 3460 56700 3490
rect 56070 3420 56100 3450
rect 56110 3420 56140 3450
rect 56150 3420 56180 3450
rect 56190 3420 56220 3450
rect 56230 3420 56260 3450
rect 56270 3420 56300 3450
rect 56310 3420 56340 3450
rect 56350 3420 56380 3450
rect 56390 3420 56420 3450
rect 56430 3420 56460 3450
rect 56470 3420 56500 3450
rect 56510 3420 56540 3450
rect 56550 3420 56580 3450
rect 56590 3420 56620 3450
rect 56630 3420 56660 3450
rect 56670 3420 56700 3450
rect 56070 3380 56100 3410
rect 56110 3380 56140 3410
rect 56150 3380 56180 3410
rect 56190 3380 56220 3410
rect 56230 3380 56260 3410
rect 56270 3380 56300 3410
rect 56310 3380 56340 3410
rect 56350 3380 56380 3410
rect 56390 3380 56420 3410
rect 56430 3380 56460 3410
rect 56470 3380 56500 3410
rect 56510 3380 56540 3410
rect 56550 3380 56580 3410
rect 56590 3380 56620 3410
rect 56630 3380 56660 3410
rect 56670 3380 56700 3410
rect 57220 3630 57250 3660
rect 57340 3630 57370 3660
rect 57460 3630 57490 3660
rect 57400 3575 57430 3580
rect 57400 3555 57405 3575
rect 57405 3555 57425 3575
rect 57425 3555 57430 3575
rect 57400 3550 57430 3555
rect 57580 3630 57610 3660
rect 57700 3630 57730 3660
rect 57100 3460 57130 3490
rect 57140 3460 57170 3490
rect 57180 3460 57210 3490
rect 57220 3460 57250 3490
rect 57260 3460 57290 3490
rect 57300 3460 57330 3490
rect 57340 3460 57370 3490
rect 57380 3460 57410 3490
rect 57420 3460 57450 3490
rect 57460 3460 57490 3490
rect 57500 3460 57530 3490
rect 57540 3460 57570 3490
rect 57580 3460 57610 3490
rect 57620 3460 57650 3490
rect 57660 3460 57690 3490
rect 57700 3460 57730 3490
rect 57100 3420 57130 3450
rect 57140 3420 57170 3450
rect 57180 3420 57210 3450
rect 57220 3420 57250 3450
rect 57260 3420 57290 3450
rect 57300 3420 57330 3450
rect 57340 3420 57370 3450
rect 57380 3420 57410 3450
rect 57420 3420 57450 3450
rect 57460 3420 57490 3450
rect 57500 3420 57530 3450
rect 57540 3420 57570 3450
rect 57580 3420 57610 3450
rect 57620 3420 57650 3450
rect 57660 3420 57690 3450
rect 57700 3420 57730 3450
rect 57100 3380 57130 3410
rect 57140 3380 57170 3410
rect 57180 3380 57210 3410
rect 57220 3380 57250 3410
rect 57260 3380 57290 3410
rect 57300 3380 57330 3410
rect 57340 3380 57370 3410
rect 57380 3380 57410 3410
rect 57420 3380 57450 3410
rect 57460 3380 57490 3410
rect 57500 3380 57530 3410
rect 57540 3380 57570 3410
rect 57580 3380 57610 3410
rect 57620 3380 57650 3410
rect 57660 3380 57690 3410
rect 57700 3380 57730 3410
rect 55625 3325 55655 3355
rect 55665 3325 55695 3355
rect 55705 3325 55735 3355
rect 58375 4290 58405 4320
rect 58375 4250 58405 4280
rect 58375 4210 58405 4240
rect 58735 4290 58765 4320
rect 58735 4250 58765 4280
rect 58735 4210 58765 4240
rect 58435 4155 58465 4185
rect 58475 4155 58505 4185
rect 58515 4155 58545 4185
rect 58555 4155 58585 4185
rect 58595 4155 58625 4185
rect 58635 4155 58665 4185
rect 58675 4155 58705 4185
rect 58435 4115 58465 4145
rect 58475 4115 58505 4145
rect 58515 4115 58545 4145
rect 58555 4115 58585 4145
rect 58595 4115 58625 4145
rect 58635 4115 58665 4145
rect 58675 4115 58705 4145
rect 58435 4075 58465 4105
rect 58475 4075 58505 4105
rect 58515 4075 58545 4105
rect 58555 4075 58585 4105
rect 58595 4075 58625 4105
rect 58635 4075 58665 4105
rect 58675 4075 58705 4105
rect 58375 4020 58405 4050
rect 58495 4020 58525 4050
rect 58615 4020 58645 4050
rect 59095 4290 59125 4320
rect 59095 4250 59125 4280
rect 59095 4210 59125 4240
rect 58795 4155 58825 4185
rect 58835 4155 58865 4185
rect 58875 4155 58905 4185
rect 58915 4155 58945 4185
rect 58955 4155 58985 4185
rect 58995 4155 59025 4185
rect 59035 4155 59065 4185
rect 58795 4115 58825 4145
rect 58835 4115 58865 4145
rect 58875 4115 58905 4145
rect 58915 4115 58945 4145
rect 58955 4115 58985 4145
rect 58995 4115 59025 4145
rect 59035 4115 59065 4145
rect 58795 4075 58825 4105
rect 58835 4075 58865 4105
rect 58875 4075 58905 4105
rect 58915 4075 58945 4105
rect 58955 4075 58985 4105
rect 58995 4075 59025 4105
rect 59035 4075 59065 4105
rect 58735 4020 58765 4050
rect 58855 4020 58885 4050
rect 58975 4020 59005 4050
rect 59645 4290 59675 4320
rect 59685 4290 59715 4320
rect 59725 4290 59755 4320
rect 59645 4250 59675 4280
rect 59685 4250 59715 4280
rect 59725 4250 59755 4280
rect 59645 4210 59675 4240
rect 59685 4210 59715 4240
rect 59725 4210 59755 4240
rect 59995 4290 60025 4320
rect 60035 4290 60065 4320
rect 60075 4290 60105 4320
rect 59995 4250 60025 4280
rect 60035 4250 60065 4280
rect 60075 4250 60105 4280
rect 59995 4210 60025 4240
rect 60035 4210 60065 4240
rect 60075 4210 60105 4240
rect 60695 4290 60725 4320
rect 60735 4290 60765 4320
rect 60775 4290 60805 4320
rect 60695 4250 60725 4280
rect 60735 4250 60765 4280
rect 60775 4250 60805 4280
rect 60695 4210 60725 4240
rect 60735 4210 60765 4240
rect 60775 4210 60805 4240
rect 61045 4290 61075 4320
rect 61085 4290 61115 4320
rect 61125 4290 61155 4320
rect 61045 4250 61075 4280
rect 61085 4250 61115 4280
rect 61125 4250 61155 4280
rect 61045 4210 61075 4240
rect 61085 4210 61115 4240
rect 61125 4210 61155 4240
rect 61395 4290 61425 4320
rect 61435 4290 61465 4320
rect 61475 4290 61505 4320
rect 61395 4250 61425 4280
rect 61435 4250 61465 4280
rect 61475 4250 61505 4280
rect 61395 4210 61425 4240
rect 61435 4210 61465 4240
rect 61475 4210 61505 4240
rect 59095 4020 59125 4050
rect 58435 3630 58465 3660
rect 58555 3630 58585 3660
rect 58675 3630 58705 3660
rect 58795 3630 58825 3660
rect 58915 3630 58945 3660
rect 59035 3630 59065 3660
rect 58735 3530 58765 3535
rect 58735 3510 58740 3530
rect 58740 3510 58760 3530
rect 58760 3510 58765 3530
rect 58735 3505 58765 3510
rect 55625 3285 55655 3315
rect 55665 3285 55695 3315
rect 55705 3285 55735 3315
rect 55625 3245 55655 3275
rect 55665 3245 55695 3275
rect 55705 3245 55735 3275
rect 56515 3315 56545 3345
rect 56515 3275 56545 3305
rect 56515 3260 56545 3265
rect 56515 3240 56520 3260
rect 56520 3240 56540 3260
rect 56540 3240 56545 3260
rect 56515 3235 56545 3240
rect 56680 3315 56710 3345
rect 56680 3275 56710 3305
rect 56680 3260 56710 3265
rect 56680 3240 56685 3260
rect 56685 3240 56705 3260
rect 56705 3240 56710 3260
rect 56680 3235 56710 3240
rect 56845 3315 56875 3345
rect 56845 3275 56875 3305
rect 56845 3260 56875 3265
rect 56845 3240 56850 3260
rect 56850 3240 56870 3260
rect 56870 3240 56875 3260
rect 56845 3235 56875 3240
rect 56925 3315 56955 3345
rect 56925 3275 56955 3305
rect 56925 3260 56955 3265
rect 56925 3240 56930 3260
rect 56930 3240 56950 3260
rect 56950 3240 56955 3260
rect 56925 3235 56955 3240
rect 57090 3315 57120 3345
rect 57090 3275 57120 3305
rect 57090 3260 57120 3265
rect 57090 3240 57095 3260
rect 57095 3240 57115 3260
rect 57115 3240 57120 3260
rect 57090 3235 57120 3240
rect 57255 3315 57285 3345
rect 57255 3275 57285 3305
rect 57255 3260 57285 3265
rect 57255 3240 57260 3260
rect 57260 3240 57280 3260
rect 57280 3240 57285 3260
rect 57255 3235 57285 3240
rect 58060 3325 58090 3355
rect 58100 3325 58130 3355
rect 58140 3325 58170 3355
rect 58060 3285 58090 3315
rect 58100 3285 58130 3315
rect 58140 3285 58170 3315
rect 58060 3245 58090 3275
rect 58100 3245 58130 3275
rect 58140 3245 58170 3275
rect 56625 3205 56655 3210
rect 56625 3185 56630 3205
rect 56630 3185 56650 3205
rect 56650 3185 56655 3205
rect 56625 3180 56655 3185
rect 56735 3205 56765 3210
rect 56735 3185 56740 3205
rect 56740 3185 56760 3205
rect 56760 3185 56765 3205
rect 56735 3180 56765 3185
rect 57035 3205 57065 3210
rect 57035 3185 57040 3205
rect 57040 3185 57060 3205
rect 57060 3185 57065 3205
rect 57035 3180 57065 3185
rect 57145 3205 57175 3210
rect 57145 3185 57150 3205
rect 57150 3185 57170 3205
rect 57170 3185 57175 3205
rect 57145 3180 57175 3185
rect 56560 2895 56590 2900
rect 56800 2895 56830 2900
rect 56560 2875 56565 2895
rect 56565 2875 56585 2895
rect 56585 2875 56590 2895
rect 56560 2870 56590 2875
rect 56680 2885 56710 2890
rect 56680 2865 56685 2885
rect 56685 2865 56705 2885
rect 56705 2865 56710 2885
rect 56680 2860 56710 2865
rect 56800 2875 56805 2895
rect 56805 2875 56825 2895
rect 56825 2875 56830 2895
rect 56800 2870 56830 2875
rect 56605 2825 56635 2830
rect 56605 2805 56610 2825
rect 56610 2805 56630 2825
rect 56630 2805 56635 2825
rect 56605 2800 56635 2805
rect 55945 2750 55975 2780
rect 56750 2750 56780 2780
rect 55625 2155 55655 2185
rect 55665 2155 55695 2185
rect 55705 2155 55735 2185
rect 55625 2115 55655 2145
rect 55665 2115 55695 2145
rect 55705 2115 55735 2145
rect 55625 2075 55655 2105
rect 55665 2075 55695 2105
rect 55705 2075 55735 2105
rect 54615 1445 54645 1475
rect 54815 1445 54845 1475
rect 54925 1445 54955 1475
rect 55035 1445 55065 1475
rect 55145 1445 55175 1475
rect 55255 1445 55285 1475
rect 54615 1125 54645 1155
rect 54460 1055 54490 1085
rect 54570 1055 54600 1085
rect 54815 1105 54845 1135
rect 54925 1105 54955 1135
rect 55035 1105 55065 1135
rect 55145 1105 55175 1135
rect 55255 1105 55285 1135
rect 54760 1045 54790 1075
rect 54760 1005 54790 1035
rect 54760 965 54790 995
rect 54870 1045 54900 1075
rect 54870 1005 54900 1035
rect 54870 965 54900 995
rect 54980 1045 55010 1075
rect 54980 1005 55010 1035
rect 54980 965 55010 995
rect 55090 1045 55120 1075
rect 55090 1005 55120 1035
rect 55090 965 55120 995
rect 55200 1045 55230 1075
rect 55200 1005 55230 1035
rect 55200 965 55230 995
rect 55310 1045 55340 1075
rect 55310 1005 55340 1035
rect 55310 965 55340 995
rect 55900 1955 55930 1985
rect 55625 1045 55655 1075
rect 55665 1045 55695 1075
rect 55705 1045 55735 1075
rect 55625 1005 55655 1035
rect 55665 1005 55695 1035
rect 55705 1005 55735 1035
rect 55625 965 55655 995
rect 55665 965 55695 995
rect 55705 965 55735 995
rect 55760 1455 55790 1485
rect 55800 1455 55830 1485
rect 55840 1455 55870 1485
rect 55760 1415 55790 1445
rect 55800 1415 55830 1445
rect 55840 1415 55870 1445
rect 55760 1375 55790 1405
rect 55800 1375 55830 1405
rect 55840 1375 55870 1405
rect 54705 910 54735 940
rect 54705 870 54735 900
rect 54705 830 54735 860
rect 55365 910 55395 940
rect 55365 870 55395 900
rect 55365 830 55395 860
rect 54340 775 54370 805
rect 54405 405 54435 435
rect 55085 430 55115 435
rect 55085 410 55090 430
rect 55090 410 55110 430
rect 55110 410 55115 430
rect 55085 405 55115 410
rect 54075 280 54105 310
rect 54115 280 54145 310
rect 54160 280 54190 310
rect 54200 280 54230 310
rect 54245 280 54275 310
rect 54285 280 54315 310
rect 54075 240 54105 270
rect 54115 240 54145 270
rect 54160 240 54190 270
rect 54200 240 54230 270
rect 54245 240 54275 270
rect 54285 240 54315 270
rect 54075 200 54105 230
rect 54115 200 54145 230
rect 54160 200 54190 230
rect 54200 200 54230 230
rect 54245 200 54275 230
rect 54285 200 54315 230
rect 54470 280 54500 310
rect 54470 240 54500 270
rect 54470 200 54500 230
rect 54835 280 54865 310
rect 54875 280 54905 310
rect 54915 280 54945 310
rect 54955 280 54985 310
rect 54995 280 55025 310
rect 55035 280 55065 310
rect 55075 280 55105 310
rect 55115 280 55145 310
rect 55155 280 55185 310
rect 55195 280 55225 310
rect 55235 280 55265 310
rect 54835 240 54865 270
rect 54875 240 54905 270
rect 54915 240 54945 270
rect 54955 240 54985 270
rect 54995 240 55025 270
rect 55035 240 55065 270
rect 55075 240 55105 270
rect 55115 240 55145 270
rect 55155 240 55185 270
rect 55195 240 55225 270
rect 55235 240 55265 270
rect 54835 200 54865 230
rect 54875 200 54905 230
rect 54915 200 54945 230
rect 54955 200 54985 230
rect 54995 200 55025 230
rect 55035 200 55065 230
rect 55075 200 55105 230
rect 55115 200 55145 230
rect 55155 200 55185 230
rect 55195 200 55225 230
rect 55235 200 55265 230
rect 54405 170 54440 175
rect 54405 145 54410 170
rect 54410 145 54435 170
rect 54435 145 54440 170
rect 54405 140 54440 145
rect 54465 170 54500 175
rect 54465 145 54470 170
rect 54470 145 54495 170
rect 54495 145 54500 170
rect 54465 140 54500 145
rect 54835 -555 54865 -525
rect 55035 -555 55065 -525
rect 55760 -125 55790 -95
rect 55800 -125 55830 -95
rect 55840 -125 55870 -95
rect 55760 -165 55790 -135
rect 55800 -165 55830 -135
rect 55840 -165 55870 -135
rect 55760 -205 55790 -175
rect 55800 -205 55830 -175
rect 55840 -205 55870 -175
rect 57090 2885 57120 2890
rect 57090 2865 57095 2885
rect 57095 2865 57115 2885
rect 57115 2865 57120 2885
rect 57090 2860 57120 2865
rect 57165 2825 57195 2830
rect 57165 2805 57170 2825
rect 57170 2805 57190 2825
rect 57190 2805 57195 2825
rect 57165 2800 57195 2805
rect 57020 2750 57050 2780
rect 56855 2695 56885 2725
rect 56965 2695 56995 2725
rect 57825 2750 57855 2780
rect 56940 2640 56970 2670
rect 57215 2640 57245 2670
rect 56855 2610 56885 2615
rect 56855 2590 56860 2610
rect 56860 2590 56880 2610
rect 56880 2590 56885 2610
rect 56855 2585 56885 2590
rect 56090 2440 56120 2470
rect 56145 2440 56175 2470
rect 56200 2440 56230 2470
rect 56255 2440 56285 2470
rect 56310 2440 56340 2470
rect 56365 2440 56395 2470
rect 56420 2440 56450 2470
rect 56475 2440 56505 2470
rect 56530 2440 56560 2470
rect 56585 2440 56615 2470
rect 56640 2440 56670 2470
rect 56090 2400 56120 2430
rect 56145 2400 56175 2430
rect 56200 2400 56230 2430
rect 56255 2400 56285 2430
rect 56310 2400 56340 2430
rect 56365 2400 56395 2430
rect 56420 2400 56450 2430
rect 56475 2400 56505 2430
rect 56530 2400 56560 2430
rect 56585 2400 56615 2430
rect 56640 2400 56670 2430
rect 56090 2360 56120 2390
rect 56145 2360 56175 2390
rect 56200 2360 56230 2390
rect 56255 2360 56285 2390
rect 56310 2360 56340 2390
rect 56365 2360 56395 2390
rect 56420 2360 56450 2390
rect 56475 2360 56505 2390
rect 56530 2360 56560 2390
rect 56585 2360 56615 2390
rect 56640 2360 56670 2390
rect 55995 1980 56025 1985
rect 55995 1960 56000 1980
rect 56000 1960 56020 1980
rect 56020 1960 56025 1980
rect 55995 1955 56025 1960
rect 56145 1945 56175 1975
rect 56090 1900 56120 1930
rect 56255 1945 56285 1975
rect 56200 1900 56230 1930
rect 56145 1710 56175 1740
rect 56090 1665 56120 1695
rect 56035 1610 56065 1640
rect 56035 1570 56065 1600
rect 56035 1530 56065 1560
rect 56365 1945 56395 1975
rect 56310 1900 56340 1930
rect 56255 1710 56285 1740
rect 56200 1665 56230 1695
rect 56040 1290 56070 1295
rect 56040 1270 56045 1290
rect 56045 1270 56065 1290
rect 56065 1270 56070 1290
rect 56090 1275 56120 1305
rect 56145 1285 56175 1315
rect 56475 1945 56505 1975
rect 56420 1900 56450 1930
rect 56365 1710 56395 1740
rect 56310 1665 56340 1695
rect 56200 1275 56230 1305
rect 56255 1285 56285 1315
rect 56585 1945 56615 1975
rect 56530 1900 56560 1930
rect 56475 1710 56505 1740
rect 56420 1665 56450 1695
rect 56310 1275 56340 1305
rect 56365 1285 56395 1315
rect 57130 2440 57160 2470
rect 57185 2440 57215 2470
rect 57240 2440 57270 2470
rect 57295 2440 57325 2470
rect 57350 2440 57380 2470
rect 57405 2440 57435 2470
rect 57460 2440 57490 2470
rect 57515 2440 57545 2470
rect 57570 2440 57600 2470
rect 57625 2440 57655 2470
rect 57680 2440 57710 2470
rect 57130 2400 57160 2430
rect 57185 2400 57215 2430
rect 57240 2400 57270 2430
rect 57295 2400 57325 2430
rect 57350 2400 57380 2430
rect 57405 2400 57435 2430
rect 57460 2400 57490 2430
rect 57515 2400 57545 2430
rect 57570 2400 57600 2430
rect 57625 2400 57655 2430
rect 57680 2400 57710 2430
rect 57130 2360 57160 2390
rect 57185 2360 57215 2390
rect 57240 2360 57270 2390
rect 57295 2360 57325 2390
rect 57350 2360 57380 2390
rect 57405 2360 57435 2390
rect 57460 2360 57490 2390
rect 57515 2360 57545 2390
rect 57570 2360 57600 2390
rect 57625 2360 57655 2390
rect 57680 2360 57710 2390
rect 56775 2290 56805 2295
rect 56775 2270 56780 2290
rect 56780 2270 56800 2290
rect 56800 2270 56805 2290
rect 56775 2265 56805 2270
rect 56775 2225 56805 2255
rect 56775 2185 56805 2215
rect 56885 2265 56915 2295
rect 56885 2225 56915 2255
rect 56885 2185 56915 2215
rect 56995 2290 57025 2295
rect 56995 2270 57000 2290
rect 57000 2270 57020 2290
rect 57020 2270 57025 2290
rect 56995 2265 57025 2270
rect 56995 2225 57025 2255
rect 56995 2185 57025 2215
rect 56690 1980 56720 1985
rect 56690 1960 56695 1980
rect 56695 1960 56715 1980
rect 56715 1960 56720 1980
rect 56690 1955 56720 1960
rect 57080 1980 57110 1985
rect 57080 1960 57085 1980
rect 57085 1960 57105 1980
rect 57105 1960 57110 1980
rect 57080 1955 57110 1960
rect 56640 1900 56670 1930
rect 57185 1945 57215 1975
rect 57130 1900 57160 1930
rect 56585 1710 56615 1740
rect 56530 1665 56560 1695
rect 56420 1275 56450 1305
rect 56475 1285 56505 1315
rect 56640 1665 56670 1695
rect 57295 1945 57325 1975
rect 57240 1900 57270 1930
rect 57185 1710 57215 1740
rect 57130 1665 57160 1695
rect 56695 1610 56725 1640
rect 56695 1570 56725 1600
rect 56695 1530 56725 1560
rect 57075 1610 57105 1640
rect 57075 1570 57105 1600
rect 57075 1530 57105 1560
rect 56885 1455 56915 1485
rect 56885 1415 56915 1445
rect 56885 1375 56915 1405
rect 56530 1275 56560 1305
rect 56585 1285 56615 1315
rect 56640 1275 56670 1305
rect 56690 1300 56720 1305
rect 56690 1280 56695 1300
rect 56695 1280 56715 1300
rect 56715 1280 56720 1300
rect 56690 1275 56720 1280
rect 56840 1300 56870 1305
rect 56840 1280 56845 1300
rect 56845 1280 56865 1300
rect 56865 1280 56870 1300
rect 56840 1275 56870 1280
rect 56040 1265 56070 1270
rect 56145 1230 56175 1260
rect 56090 1035 56120 1065
rect 56255 1230 56285 1260
rect 56200 1035 56230 1065
rect 56365 1230 56395 1260
rect 56310 1035 56340 1065
rect 56475 1230 56505 1260
rect 56420 1035 56450 1065
rect 56585 1230 56615 1260
rect 56530 1035 56560 1065
rect 56640 1035 56670 1065
rect 57405 1945 57435 1975
rect 57350 1900 57380 1930
rect 57295 1710 57325 1740
rect 57240 1665 57270 1695
rect 56930 1300 56960 1305
rect 56930 1280 56935 1300
rect 56935 1280 56955 1300
rect 56955 1280 56960 1300
rect 56930 1275 56960 1280
rect 57080 1300 57110 1305
rect 57080 1280 57085 1300
rect 57085 1280 57105 1300
rect 57105 1280 57110 1300
rect 57080 1275 57110 1280
rect 57130 1275 57160 1305
rect 57185 1285 57215 1315
rect 57515 1945 57545 1975
rect 57460 1900 57490 1930
rect 57405 1710 57435 1740
rect 57350 1665 57380 1695
rect 57240 1275 57270 1305
rect 57295 1285 57325 1315
rect 57625 1945 57655 1975
rect 57570 1900 57600 1930
rect 57515 1710 57545 1740
rect 57460 1665 57490 1695
rect 57350 1275 57380 1305
rect 57405 1285 57435 1315
rect 57680 1900 57710 1930
rect 57625 1710 57655 1740
rect 57570 1665 57600 1695
rect 57460 1275 57490 1305
rect 57515 1285 57545 1315
rect 57680 1665 57710 1695
rect 57735 1610 57765 1640
rect 57735 1570 57765 1600
rect 57735 1530 57765 1560
rect 57570 1275 57600 1305
rect 57625 1285 57655 1315
rect 57680 1275 57710 1305
rect 57730 1290 57760 1295
rect 57730 1270 57735 1290
rect 57735 1270 57755 1290
rect 57755 1270 57760 1290
rect 57185 1230 57215 1260
rect 56830 1035 56860 1065
rect 56145 965 56175 995
rect 56255 965 56285 995
rect 56365 965 56395 995
rect 56475 965 56505 995
rect 56585 965 56615 995
rect 56035 910 56065 940
rect 56035 870 56065 900
rect 56035 830 56065 860
rect 55945 775 55975 805
rect 56735 910 56765 940
rect 56735 870 56765 900
rect 56735 830 56765 860
rect 56445 360 56475 390
rect 56555 360 56585 390
rect 56665 360 56695 390
rect 56775 360 56805 390
rect 56940 1035 56970 1065
rect 56885 360 56915 390
rect 57130 1035 57160 1065
rect 57295 1230 57325 1260
rect 57240 1035 57270 1065
rect 57405 1230 57435 1260
rect 57350 1035 57380 1065
rect 57515 1230 57545 1260
rect 57460 1035 57490 1065
rect 57625 1230 57655 1260
rect 57570 1035 57600 1065
rect 57730 1265 57760 1270
rect 57680 1035 57710 1065
rect 57185 965 57215 995
rect 57295 965 57325 995
rect 57035 910 57065 940
rect 57035 870 57065 900
rect 57035 830 57065 860
rect 56995 360 57025 390
rect 57405 965 57435 995
rect 57515 965 57545 995
rect 57625 965 57655 995
rect 57735 910 57765 940
rect 57735 870 57765 900
rect 57735 830 57765 860
rect 57870 2640 57900 2670
rect 57825 775 57855 805
rect 57105 360 57135 390
rect 57215 360 57245 390
rect 57325 360 57355 390
rect 57435 360 57465 390
rect 56225 55 56255 60
rect 56225 35 56230 55
rect 56230 35 56250 55
rect 56250 35 56255 55
rect 56225 30 56255 35
rect 55900 -305 55930 -275
rect 55235 -555 55265 -525
rect 56280 30 56310 60
rect 56390 30 56420 60
rect 56500 30 56530 60
rect 56610 30 56640 60
rect 56720 30 56750 60
rect 56830 30 56860 60
rect 56940 30 56970 60
rect 57050 30 57080 60
rect 57160 30 57190 60
rect 57270 30 57300 60
rect 57380 30 57410 60
rect 57490 55 57520 60
rect 57490 35 57495 55
rect 57495 35 57515 55
rect 57515 35 57520 55
rect 57490 30 57520 35
rect 56445 -15 56475 15
rect 56555 -15 56585 15
rect 56665 -15 56695 15
rect 56775 -15 56805 15
rect 56885 -15 56915 15
rect 56995 -15 57025 15
rect 57105 -15 57135 15
rect 57215 -15 57245 15
rect 57325 -15 57355 15
rect 57435 -15 57465 15
rect 56335 -125 56365 -95
rect 56335 -165 56365 -135
rect 56335 -205 56365 -175
rect 56545 -260 56575 -230
rect 56655 -260 56685 -230
rect 56875 -260 56905 -230
rect 56490 -305 56520 -275
rect 56600 -280 56630 -275
rect 56600 -300 56605 -280
rect 56605 -300 56625 -280
rect 56625 -300 56630 -280
rect 56600 -305 56630 -300
rect 56545 -510 56575 -480
rect 56710 -305 56740 -275
rect 56655 -510 56685 -480
rect 57045 -280 57075 -275
rect 57045 -300 57050 -280
rect 57050 -300 57070 -280
rect 57070 -300 57075 -280
rect 57045 -305 57075 -300
rect 57420 -45 57450 -40
rect 57420 -65 57425 -45
rect 57425 -65 57445 -45
rect 57445 -65 57450 -45
rect 57420 -70 57450 -65
rect 56875 -510 56905 -480
rect 56490 -555 56520 -525
rect 56600 -555 56630 -525
rect 56710 -555 56740 -525
rect 52295 -610 52325 -580
rect 52335 -610 52365 -580
rect 52375 -610 52405 -580
rect 52295 -650 52325 -620
rect 52335 -650 52365 -620
rect 52375 -650 52405 -620
rect 52295 -690 52325 -660
rect 52335 -690 52365 -660
rect 52375 -690 52405 -660
rect 52645 -610 52675 -580
rect 52685 -610 52715 -580
rect 52725 -610 52755 -580
rect 52645 -650 52675 -620
rect 52685 -650 52715 -620
rect 52725 -650 52755 -620
rect 52645 -690 52675 -660
rect 52685 -690 52715 -660
rect 52725 -690 52755 -660
rect 52995 -610 53025 -580
rect 53035 -610 53065 -580
rect 53075 -610 53105 -580
rect 52995 -650 53025 -620
rect 53035 -650 53065 -620
rect 53075 -650 53105 -620
rect 52995 -690 53025 -660
rect 53035 -690 53065 -660
rect 53075 -690 53105 -660
rect 53345 -610 53375 -580
rect 53385 -610 53415 -580
rect 53425 -610 53455 -580
rect 53345 -650 53375 -620
rect 53385 -650 53415 -620
rect 53425 -650 53455 -620
rect 53345 -690 53375 -660
rect 53385 -690 53415 -660
rect 53425 -690 53455 -660
rect 53695 -610 53725 -580
rect 53735 -610 53765 -580
rect 53775 -610 53805 -580
rect 53925 -610 53955 -580
rect 53965 -610 53995 -580
rect 54005 -610 54035 -580
rect 54045 -610 54075 -580
rect 54085 -610 54115 -580
rect 54125 -610 54155 -580
rect 53695 -650 53725 -620
rect 53735 -650 53765 -620
rect 53775 -650 53805 -620
rect 53925 -650 53955 -620
rect 53965 -650 53995 -620
rect 54005 -650 54035 -620
rect 54045 -650 54075 -620
rect 54085 -650 54115 -620
rect 54125 -650 54155 -620
rect 53695 -690 53725 -660
rect 53735 -690 53765 -660
rect 53775 -690 53805 -660
rect 53925 -690 53955 -660
rect 53965 -690 53995 -660
rect 54005 -690 54035 -660
rect 54045 -690 54075 -660
rect 54085 -690 54115 -660
rect 54125 -690 54155 -660
rect 54395 -610 54425 -580
rect 54435 -610 54465 -580
rect 54475 -610 54505 -580
rect 54395 -650 54425 -620
rect 54435 -650 54465 -620
rect 54475 -650 54505 -620
rect 54395 -690 54425 -660
rect 54435 -690 54465 -660
rect 54475 -690 54505 -660
rect 54745 -610 54775 -580
rect 54785 -610 54815 -580
rect 54825 -610 54855 -580
rect 54745 -650 54775 -620
rect 54785 -650 54815 -620
rect 54825 -650 54855 -620
rect 54745 -690 54775 -660
rect 54785 -690 54815 -660
rect 54825 -690 54855 -660
rect 54935 -610 54965 -580
rect 54935 -650 54965 -620
rect 54935 -690 54965 -660
rect 55095 -610 55125 -580
rect 55135 -610 55165 -580
rect 55175 -610 55205 -580
rect 55095 -650 55125 -620
rect 55135 -650 55165 -620
rect 55175 -650 55205 -620
rect 55095 -690 55125 -660
rect 55135 -690 55165 -660
rect 55175 -690 55205 -660
rect 55325 -610 55355 -580
rect 55365 -610 55395 -580
rect 55405 -610 55435 -580
rect 55445 -610 55475 -580
rect 55485 -610 55515 -580
rect 55525 -610 55555 -580
rect 55325 -650 55355 -620
rect 55365 -650 55395 -620
rect 55405 -650 55435 -620
rect 55445 -650 55475 -620
rect 55485 -650 55515 -620
rect 55525 -650 55555 -620
rect 55325 -690 55355 -660
rect 55365 -690 55395 -660
rect 55405 -690 55435 -660
rect 55445 -690 55475 -660
rect 55485 -690 55515 -660
rect 55525 -690 55555 -660
rect 55795 -610 55825 -580
rect 55835 -610 55865 -580
rect 55875 -610 55905 -580
rect 55795 -650 55825 -620
rect 55835 -650 55865 -620
rect 55875 -650 55905 -620
rect 55795 -690 55825 -660
rect 55835 -690 55865 -660
rect 55875 -690 55905 -660
rect 56145 -610 56175 -580
rect 56185 -610 56215 -580
rect 56225 -610 56255 -580
rect 56145 -650 56175 -620
rect 56185 -650 56215 -620
rect 56225 -650 56255 -620
rect 56145 -690 56175 -660
rect 56185 -690 56215 -660
rect 56225 -690 56255 -660
rect 56435 -610 56465 -580
rect 56435 -650 56465 -620
rect 56435 -690 56465 -660
rect 56495 -610 56525 -580
rect 56535 -610 56565 -580
rect 56575 -610 56605 -580
rect 56495 -650 56525 -620
rect 56535 -650 56565 -620
rect 56575 -650 56605 -620
rect 56495 -690 56525 -660
rect 56535 -690 56565 -660
rect 56575 -690 56605 -660
rect 56765 -610 56795 -580
rect 56765 -650 56795 -620
rect 56765 -690 56795 -660
rect 56845 -610 56875 -580
rect 56885 -610 56915 -580
rect 56925 -610 56955 -580
rect 56845 -650 56875 -620
rect 56885 -650 56915 -620
rect 56925 -650 56955 -620
rect 56845 -690 56875 -660
rect 56885 -690 56915 -660
rect 56925 -690 56955 -660
rect 57195 -610 57225 -580
rect 57235 -610 57265 -580
rect 57275 -610 57305 -580
rect 57195 -650 57225 -620
rect 57235 -650 57265 -620
rect 57275 -650 57305 -620
rect 57195 -690 57225 -660
rect 57235 -690 57265 -660
rect 57275 -690 57305 -660
rect 57925 2265 57955 2295
rect 57965 2265 57995 2295
rect 58005 2265 58035 2295
rect 57925 2225 57955 2255
rect 57965 2225 57995 2255
rect 58005 2225 58035 2255
rect 57925 2185 57955 2215
rect 57965 2185 57995 2215
rect 58005 2185 58035 2215
rect 57925 2020 57955 2050
rect 57965 2020 57995 2050
rect 58005 2020 58035 2050
rect 57925 1980 57955 2010
rect 57965 1980 57995 2010
rect 58005 1980 58035 2010
rect 57925 1940 57955 1970
rect 57965 1940 57995 1970
rect 58005 1940 58035 1970
rect 57925 1610 57955 1640
rect 57965 1610 57995 1640
rect 58005 1610 58035 1640
rect 57925 1570 57955 1600
rect 57965 1570 57995 1600
rect 58005 1570 58035 1600
rect 57925 1530 57955 1560
rect 57965 1530 57995 1560
rect 58005 1530 58035 1560
rect 58060 2155 58090 2185
rect 58100 2155 58130 2185
rect 58140 2155 58170 2185
rect 58060 2115 58090 2145
rect 58100 2115 58130 2145
rect 58140 2115 58170 2145
rect 58060 2075 58090 2105
rect 58100 2075 58130 2105
rect 58140 2075 58170 2105
rect 57925 1455 57955 1485
rect 57965 1455 57995 1485
rect 58005 1455 58035 1485
rect 57925 1415 57955 1445
rect 57965 1415 57995 1445
rect 58005 1415 58035 1445
rect 57925 1375 57955 1405
rect 57965 1375 57995 1405
rect 58005 1375 58035 1405
rect 57870 -70 57900 -40
rect 58195 3460 58225 3490
rect 58235 3460 58265 3490
rect 58275 3460 58305 3490
rect 58195 3420 58225 3450
rect 58235 3420 58265 3450
rect 58275 3420 58305 3450
rect 58195 3380 58225 3410
rect 58235 3380 58265 3410
rect 58275 3380 58305 3410
rect 58405 3325 58435 3355
rect 58405 3285 58435 3315
rect 58405 3245 58435 3275
rect 58515 3325 58545 3355
rect 58515 3285 58545 3315
rect 58515 3245 58545 3275
rect 58625 3325 58655 3355
rect 58625 3285 58655 3315
rect 58625 3245 58655 3275
rect 58735 3325 58765 3355
rect 58735 3285 58765 3315
rect 58735 3245 58765 3275
rect 58845 3325 58875 3355
rect 58845 3285 58875 3315
rect 58845 3245 58875 3275
rect 58955 3325 58985 3355
rect 58955 3285 58985 3315
rect 58955 3245 58985 3275
rect 59065 3325 59095 3355
rect 59510 3345 59540 3375
rect 59065 3285 59095 3315
rect 59065 3245 59095 3275
rect 58460 3160 58490 3190
rect 58570 3160 58600 3190
rect 58680 3160 58710 3190
rect 58790 3160 58820 3190
rect 58900 3160 58930 3190
rect 59010 3160 59040 3190
rect 58195 2440 58225 2470
rect 58235 2440 58265 2470
rect 58275 2440 58305 2470
rect 58195 2400 58225 2430
rect 58235 2400 58265 2430
rect 58275 2400 58305 2430
rect 58195 2360 58225 2390
rect 58235 2360 58265 2390
rect 58275 2360 58305 2390
rect 58460 2520 58490 2550
rect 58570 2520 58600 2550
rect 58680 2520 58710 2550
rect 58790 2520 58820 2550
rect 58735 2465 58765 2470
rect 58735 2445 58740 2465
rect 58740 2445 58760 2465
rect 58760 2445 58765 2465
rect 58735 2440 58765 2445
rect 58735 2425 58765 2430
rect 58735 2405 58740 2425
rect 58740 2405 58760 2425
rect 58760 2405 58765 2425
rect 58735 2400 58765 2405
rect 58735 2385 58765 2390
rect 58735 2365 58740 2385
rect 58740 2365 58760 2385
rect 58760 2365 58765 2385
rect 58735 2360 58765 2365
rect 58900 2520 58930 2550
rect 59010 2520 59040 2550
rect 59470 2440 59500 2470
rect 59510 2440 59540 2470
rect 59550 2440 59580 2470
rect 59470 2400 59500 2430
rect 59510 2400 59540 2430
rect 59550 2400 59580 2430
rect 59470 2360 59500 2390
rect 59510 2360 59540 2390
rect 59550 2360 59580 2390
rect 58460 2290 58490 2320
rect 58515 2290 58545 2320
rect 58570 2290 58600 2320
rect 58625 2290 58655 2320
rect 58680 2290 58710 2320
rect 58735 2290 58765 2320
rect 58790 2290 58820 2320
rect 58845 2290 58875 2320
rect 58900 2290 58930 2320
rect 58955 2290 58985 2320
rect 59010 2290 59040 2320
rect 58460 2250 58490 2280
rect 58515 2250 58545 2280
rect 58570 2250 58600 2280
rect 58625 2250 58655 2280
rect 58680 2250 58710 2280
rect 58735 2250 58765 2280
rect 58790 2250 58820 2280
rect 58845 2250 58875 2280
rect 58900 2250 58930 2280
rect 58955 2250 58985 2280
rect 59010 2250 59040 2280
rect 58460 2210 58490 2240
rect 58515 2210 58545 2240
rect 58570 2210 58600 2240
rect 58625 2210 58655 2240
rect 58680 2210 58710 2240
rect 58735 2210 58765 2240
rect 58790 2210 58820 2240
rect 58845 2210 58875 2240
rect 58900 2210 58930 2240
rect 58955 2210 58985 2240
rect 59010 2210 59040 2240
rect 59485 2290 59515 2320
rect 59525 2290 59555 2320
rect 59570 2290 59600 2320
rect 59610 2290 59640 2320
rect 59655 2290 59685 2320
rect 59695 2290 59725 2320
rect 59485 2250 59515 2280
rect 59525 2250 59555 2280
rect 59570 2250 59600 2280
rect 59610 2250 59640 2280
rect 59655 2250 59685 2280
rect 59695 2250 59725 2280
rect 59485 2210 59515 2240
rect 59525 2210 59555 2240
rect 59570 2210 59600 2240
rect 59610 2210 59640 2240
rect 59655 2210 59685 2240
rect 59695 2210 59725 2240
rect 58405 2155 58435 2185
rect 58405 2115 58435 2145
rect 58405 2075 58435 2105
rect 59065 2155 59095 2185
rect 59065 2115 59095 2145
rect 59065 2075 59095 2105
rect 58460 2020 58490 2050
rect 58460 1980 58490 2010
rect 58460 1940 58490 1970
rect 58570 2020 58600 2050
rect 58570 1980 58600 2010
rect 58570 1940 58600 1970
rect 58680 2020 58710 2050
rect 58680 1980 58710 2010
rect 58680 1940 58710 1970
rect 58790 2020 58820 2050
rect 58790 1980 58820 2010
rect 58790 1940 58820 1970
rect 58900 2020 58930 2050
rect 58900 1980 58930 2010
rect 58900 1940 58930 1970
rect 59010 2020 59040 2050
rect 59010 1980 59040 2010
rect 59010 1940 59040 1970
rect 58515 1885 58545 1915
rect 58625 1885 58655 1915
rect 58735 1885 58765 1915
rect 58845 1885 58875 1915
rect 58955 1885 58985 1915
rect 59490 1680 59520 1710
rect 59540 1680 59570 1710
rect 59590 1680 59620 1710
rect 59640 1680 59670 1710
rect 59690 1680 59720 1710
rect 58515 1655 58545 1660
rect 58515 1635 58520 1655
rect 58520 1635 58540 1655
rect 58540 1635 58545 1655
rect 58515 1630 58545 1635
rect 58625 1655 58655 1660
rect 58625 1635 58630 1655
rect 58630 1635 58650 1655
rect 58650 1635 58655 1655
rect 58625 1630 58655 1635
rect 58735 1655 58765 1660
rect 58735 1635 58740 1655
rect 58740 1635 58760 1655
rect 58760 1635 58765 1655
rect 58735 1630 58765 1635
rect 58845 1655 58875 1660
rect 58845 1635 58850 1655
rect 58850 1635 58870 1655
rect 58870 1635 58875 1655
rect 58845 1630 58875 1635
rect 58955 1655 58985 1660
rect 58955 1635 58960 1655
rect 58960 1635 58980 1655
rect 58980 1635 58985 1655
rect 58955 1630 58985 1635
rect 59200 1630 59230 1660
rect 59490 1630 59520 1660
rect 59540 1630 59570 1660
rect 59590 1630 59620 1660
rect 59640 1630 59670 1660
rect 59690 1630 59720 1660
rect 58195 1565 58225 1595
rect 58235 1565 58265 1595
rect 58275 1565 58305 1595
rect 58195 1525 58225 1555
rect 58235 1525 58265 1555
rect 58275 1525 58305 1555
rect 58570 1590 58600 1595
rect 58570 1570 58575 1590
rect 58575 1570 58595 1590
rect 58595 1570 58600 1590
rect 58570 1565 58600 1570
rect 58570 1550 58600 1555
rect 58570 1530 58575 1550
rect 58575 1530 58595 1550
rect 58595 1530 58600 1550
rect 58570 1525 58600 1530
rect 58515 1445 58545 1475
rect 58625 1445 58655 1475
rect 58735 1445 58765 1475
rect 58845 1445 58875 1475
rect 58955 1445 58985 1475
rect 59155 1445 59185 1475
rect 58060 1050 58090 1080
rect 58100 1050 58130 1080
rect 58140 1050 58170 1080
rect 58060 1010 58090 1040
rect 58100 1010 58130 1040
rect 58140 1010 58170 1040
rect 58060 970 58090 1000
rect 58100 970 58130 1000
rect 58140 970 58170 1000
rect 58515 1105 58545 1135
rect 58625 1105 58655 1135
rect 58735 1105 58765 1135
rect 58845 1105 58875 1135
rect 58955 1105 58985 1135
rect 59155 1125 59185 1155
rect 58460 1050 58490 1080
rect 58460 1010 58490 1040
rect 58460 970 58490 1000
rect 58570 1050 58600 1080
rect 58570 1010 58600 1040
rect 58570 970 58600 1000
rect 58680 1050 58710 1080
rect 58680 1010 58710 1040
rect 58680 970 58710 1000
rect 58790 1050 58820 1080
rect 58790 1010 58820 1040
rect 58790 970 58820 1000
rect 58900 1050 58930 1080
rect 58900 1010 58930 1040
rect 58900 970 58930 1000
rect 59010 1050 59040 1080
rect 59010 1010 59040 1040
rect 59010 970 59040 1000
rect 59490 1580 59520 1610
rect 59540 1580 59570 1610
rect 59590 1580 59620 1610
rect 59640 1580 59670 1610
rect 59690 1580 59720 1610
rect 59250 1155 59285 1160
rect 59250 1130 59255 1155
rect 59255 1130 59280 1155
rect 59280 1130 59285 1155
rect 59250 1125 59285 1130
rect 59310 1155 59345 1160
rect 59310 1130 59315 1155
rect 59315 1130 59340 1155
rect 59340 1130 59345 1155
rect 59310 1125 59345 1130
rect 59370 1155 59405 1160
rect 59370 1130 59375 1155
rect 59375 1130 59400 1155
rect 59400 1130 59405 1155
rect 59370 1125 59405 1130
rect 59430 1155 59465 1160
rect 59430 1130 59435 1155
rect 59435 1130 59460 1155
rect 59460 1130 59465 1155
rect 59430 1125 59465 1130
rect 59200 1055 59230 1085
rect 59310 1055 59340 1085
rect 58405 910 58435 940
rect 58405 870 58435 900
rect 58405 830 58435 860
rect 59065 910 59095 940
rect 59065 870 59095 900
rect 59065 830 59095 860
rect 59430 775 59460 805
rect 58685 430 58715 435
rect 58685 410 58690 430
rect 58690 410 58710 430
rect 58710 410 58715 430
rect 58685 405 58715 410
rect 59365 405 59395 435
rect 58535 280 58565 310
rect 58575 280 58605 310
rect 58615 280 58645 310
rect 58655 280 58685 310
rect 58695 280 58725 310
rect 58735 280 58765 310
rect 58775 280 58805 310
rect 58815 280 58845 310
rect 58855 280 58885 310
rect 58895 280 58925 310
rect 58935 280 58965 310
rect 58535 240 58565 270
rect 58575 240 58605 270
rect 58615 240 58645 270
rect 58655 240 58685 270
rect 58695 240 58725 270
rect 58735 240 58765 270
rect 58775 240 58805 270
rect 58815 240 58845 270
rect 58855 240 58885 270
rect 58895 240 58925 270
rect 58935 240 58965 270
rect 58535 200 58565 230
rect 58575 200 58605 230
rect 58615 200 58645 230
rect 58655 200 58685 230
rect 58695 200 58725 230
rect 58735 200 58765 230
rect 58775 200 58805 230
rect 58815 200 58845 230
rect 58855 200 58885 230
rect 58895 200 58925 230
rect 58935 200 58965 230
rect 59300 280 59330 310
rect 59300 240 59330 270
rect 59300 200 59330 230
rect 57925 -125 57955 -95
rect 57965 -125 57995 -95
rect 58005 -125 58035 -95
rect 57925 -165 57955 -135
rect 57965 -165 57995 -135
rect 58005 -165 58035 -135
rect 57925 -205 57955 -175
rect 57965 -205 57995 -175
rect 58005 -205 58035 -175
rect 58535 -555 58565 -525
rect 58735 -555 58765 -525
rect 59485 280 59515 310
rect 59525 280 59555 310
rect 59570 280 59600 310
rect 59610 280 59640 310
rect 59655 280 59685 310
rect 59695 280 59725 310
rect 59485 240 59515 270
rect 59525 240 59555 270
rect 59570 240 59600 270
rect 59610 240 59640 270
rect 59655 240 59685 270
rect 59695 240 59725 270
rect 59485 200 59515 230
rect 59525 200 59555 230
rect 59570 200 59600 230
rect 59610 200 59640 230
rect 59655 200 59685 230
rect 59695 200 59725 230
rect 59765 2020 59795 2050
rect 59805 2020 59835 2050
rect 59845 2020 59875 2050
rect 59765 1980 59795 2010
rect 59805 1980 59835 2010
rect 59845 1980 59875 2010
rect 59765 1940 59795 1970
rect 59805 1940 59835 1970
rect 59845 1940 59875 1970
rect 59765 910 59795 940
rect 59805 910 59835 940
rect 59845 910 59875 940
rect 59765 870 59795 900
rect 59805 870 59835 900
rect 59845 870 59875 900
rect 59765 830 59795 860
rect 59805 830 59835 860
rect 59845 830 59875 860
rect 59300 170 59335 175
rect 59300 145 59305 170
rect 59305 145 59330 170
rect 59330 145 59335 170
rect 59300 140 59335 145
rect 59360 170 59395 175
rect 59360 145 59365 170
rect 59365 145 59390 170
rect 59390 145 59395 170
rect 59360 140 59395 145
rect 58935 -555 58965 -525
rect 57490 -610 57520 -580
rect 57490 -650 57520 -620
rect 57490 -690 57520 -660
rect 57545 -610 57575 -580
rect 57585 -610 57615 -580
rect 57625 -610 57655 -580
rect 57545 -650 57575 -620
rect 57585 -650 57615 -620
rect 57625 -650 57655 -620
rect 57545 -690 57575 -660
rect 57585 -690 57615 -660
rect 57625 -690 57655 -660
rect 57895 -610 57925 -580
rect 57935 -610 57965 -580
rect 57975 -610 58005 -580
rect 57895 -650 57925 -620
rect 57935 -650 57965 -620
rect 57975 -650 58005 -620
rect 57895 -690 57925 -660
rect 57935 -690 57965 -660
rect 57975 -690 58005 -660
rect 58245 -610 58275 -580
rect 58285 -610 58315 -580
rect 58325 -610 58355 -580
rect 58365 -610 58395 -580
rect 58405 -610 58435 -580
rect 58445 -610 58475 -580
rect 58245 -650 58275 -620
rect 58285 -650 58315 -620
rect 58325 -650 58355 -620
rect 58365 -650 58395 -620
rect 58405 -650 58435 -620
rect 58445 -650 58475 -620
rect 58245 -690 58275 -660
rect 58285 -690 58315 -660
rect 58325 -690 58355 -660
rect 58365 -690 58395 -660
rect 58405 -690 58435 -660
rect 58445 -690 58475 -660
rect 58595 -610 58625 -580
rect 58635 -610 58665 -580
rect 58675 -610 58705 -580
rect 58595 -650 58625 -620
rect 58635 -650 58665 -620
rect 58675 -650 58705 -620
rect 58595 -690 58625 -660
rect 58635 -690 58665 -660
rect 58675 -690 58705 -660
rect 58835 -610 58865 -580
rect 58835 -650 58865 -620
rect 58835 -690 58865 -660
rect 58945 -610 58975 -580
rect 58985 -610 59015 -580
rect 59025 -610 59055 -580
rect 58945 -650 58975 -620
rect 58985 -650 59015 -620
rect 59025 -650 59055 -620
rect 58945 -690 58975 -660
rect 58985 -690 59015 -660
rect 59025 -690 59055 -660
rect 59295 -610 59325 -580
rect 59335 -610 59365 -580
rect 59375 -610 59405 -580
rect 59295 -650 59325 -620
rect 59335 -650 59365 -620
rect 59375 -650 59405 -620
rect 59295 -690 59325 -660
rect 59335 -690 59365 -660
rect 59375 -690 59405 -660
rect 59645 -610 59675 -580
rect 59685 -610 59715 -580
rect 59725 -610 59755 -580
rect 59765 -610 59795 -580
rect 59805 -610 59835 -580
rect 59845 -610 59875 -580
rect 59645 -650 59675 -620
rect 59685 -650 59715 -620
rect 59725 -650 59755 -620
rect 59765 -650 59795 -620
rect 59805 -650 59835 -620
rect 59845 -650 59875 -620
rect 59645 -690 59675 -660
rect 59685 -690 59715 -660
rect 59725 -690 59755 -660
rect 59765 -690 59795 -660
rect 59805 -690 59835 -660
rect 59845 -690 59875 -660
rect 59995 -610 60025 -580
rect 60035 -610 60065 -580
rect 60075 -610 60105 -580
rect 59995 -650 60025 -620
rect 60035 -650 60065 -620
rect 60075 -650 60105 -620
rect 59995 -690 60025 -660
rect 60035 -690 60065 -660
rect 60075 -690 60105 -660
rect 60345 -610 60375 -580
rect 60385 -610 60415 -580
rect 60425 -610 60455 -580
rect 60345 -650 60375 -620
rect 60385 -650 60415 -620
rect 60425 -650 60455 -620
rect 60345 -690 60375 -660
rect 60385 -690 60415 -660
rect 60425 -690 60455 -660
rect 60695 -610 60725 -580
rect 60735 -610 60765 -580
rect 60775 -610 60805 -580
rect 60695 -650 60725 -620
rect 60735 -650 60765 -620
rect 60775 -650 60805 -620
rect 60695 -690 60725 -660
rect 60735 -690 60765 -660
rect 60775 -690 60805 -660
rect 61045 -610 61075 -580
rect 61085 -610 61115 -580
rect 61125 -610 61155 -580
rect 61045 -650 61075 -620
rect 61085 -650 61115 -620
rect 61125 -650 61155 -620
rect 61045 -690 61075 -660
rect 61085 -690 61115 -660
rect 61125 -690 61155 -660
rect 61395 -610 61425 -580
rect 61435 -610 61465 -580
rect 61475 -610 61505 -580
rect 61395 -650 61425 -620
rect 61435 -650 61465 -620
rect 61475 -650 61505 -620
rect 61395 -690 61425 -660
rect 61435 -690 61465 -660
rect 61475 -690 61505 -660
<< metal2 >>
rect 56205 5065 56245 5070
rect 56205 5035 56210 5065
rect 56240 5060 56245 5065
rect 56675 5065 56715 5070
rect 56675 5060 56680 5065
rect 56240 5040 56680 5060
rect 56240 5035 56245 5040
rect 56205 5030 56245 5035
rect 56675 5035 56680 5040
rect 56710 5035 56715 5065
rect 56675 5030 56715 5035
rect 57085 5065 57125 5070
rect 57085 5035 57090 5065
rect 57120 5060 57125 5065
rect 57555 5065 57595 5070
rect 57555 5060 57560 5065
rect 57120 5040 57560 5060
rect 57120 5035 57125 5040
rect 57085 5030 57125 5035
rect 57555 5035 57560 5040
rect 57590 5035 57595 5065
rect 57555 5030 57595 5035
rect 56880 5010 57245 5015
rect 56880 4980 56885 5010
rect 56915 4980 57030 5010
rect 57060 4980 57150 5010
rect 57180 4980 57210 5010
rect 57240 4980 57245 5010
rect 56880 4970 57245 4980
rect 56880 4940 56885 4970
rect 56915 4940 57030 4970
rect 57060 4940 57150 4970
rect 57180 4940 57210 4970
rect 57240 4940 57245 4970
rect 56085 4930 56125 4935
rect 56085 4900 56090 4930
rect 56120 4925 56125 4930
rect 56205 4930 56245 4935
rect 56205 4925 56210 4930
rect 56120 4905 56210 4925
rect 56120 4900 56125 4905
rect 56085 4895 56125 4900
rect 56205 4900 56210 4905
rect 56240 4925 56245 4930
rect 56265 4930 56305 4935
rect 56265 4925 56270 4930
rect 56240 4905 56270 4925
rect 56240 4900 56245 4905
rect 56205 4895 56245 4900
rect 56265 4900 56270 4905
rect 56300 4900 56305 4930
rect 56265 4895 56305 4900
rect 56880 4930 57245 4940
rect 56880 4900 56885 4930
rect 56915 4900 57030 4930
rect 57060 4900 57150 4930
rect 57180 4900 57210 4930
rect 57240 4900 57245 4930
rect 56880 4895 57245 4900
rect 57495 4930 57535 4935
rect 57495 4900 57500 4930
rect 57530 4925 57535 4930
rect 57555 4930 57595 4935
rect 57555 4925 57560 4930
rect 57530 4905 57560 4925
rect 57530 4900 57535 4905
rect 57495 4895 57535 4900
rect 57555 4900 57560 4905
rect 57590 4925 57595 4930
rect 57675 4930 57715 4935
rect 57675 4925 57680 4930
rect 57590 4905 57680 4925
rect 57590 4900 57595 4905
rect 57555 4895 57595 4900
rect 57675 4900 57680 4905
rect 57710 4900 57715 4930
rect 57675 4895 57715 4900
rect 56555 4840 56920 4845
rect 56555 4810 56560 4840
rect 56590 4810 56620 4840
rect 56650 4810 56740 4840
rect 56770 4810 56885 4840
rect 56915 4810 56920 4840
rect 56555 4800 56920 4810
rect 56555 4770 56560 4800
rect 56590 4770 56620 4800
rect 56650 4770 56740 4800
rect 56770 4770 56885 4800
rect 56915 4770 56920 4800
rect 56555 4760 56920 4770
rect 56555 4730 56560 4760
rect 56590 4730 56620 4760
rect 56650 4730 56740 4760
rect 56770 4730 56885 4760
rect 56915 4730 56920 4760
rect 56555 4725 56920 4730
rect 56205 4525 56245 4530
rect 56205 4495 56210 4525
rect 56240 4520 56245 4525
rect 56675 4525 56715 4530
rect 56675 4520 56680 4525
rect 56240 4500 56680 4520
rect 56240 4495 56245 4500
rect 56205 4490 56245 4495
rect 56675 4495 56680 4500
rect 56710 4495 56715 4525
rect 56675 4490 56715 4495
rect 57085 4525 57125 4530
rect 57085 4495 57090 4525
rect 57120 4520 57125 4525
rect 57555 4525 57595 4530
rect 57555 4520 57560 4525
rect 57120 4500 57560 4520
rect 57120 4495 57125 4500
rect 57085 4490 57125 4495
rect 57555 4495 57560 4500
rect 57590 4495 57595 4525
rect 57555 4490 57595 4495
rect 56150 4480 56190 4485
rect 56150 4450 56155 4480
rect 56185 4475 56190 4480
rect 56630 4480 56660 4485
rect 56185 4455 56630 4475
rect 56185 4450 56190 4455
rect 56150 4445 56190 4450
rect 56825 4480 56865 4485
rect 56825 4475 56830 4480
rect 56660 4455 56830 4475
rect 56630 4445 56660 4450
rect 56825 4450 56830 4455
rect 56860 4475 56865 4480
rect 56860 4470 57606 4475
rect 56860 4455 57576 4470
rect 56860 4450 56865 4455
rect 56825 4445 56865 4450
rect 57576 4435 57606 4440
rect 56935 4425 56975 4430
rect 56935 4395 56940 4425
rect 56970 4410 56975 4425
rect 57135 4415 57175 4420
rect 57135 4410 57140 4415
rect 56970 4395 57140 4410
rect 56935 4390 57140 4395
rect 57135 4385 57140 4390
rect 57170 4410 57175 4415
rect 57615 4415 57655 4420
rect 57615 4410 57620 4415
rect 57170 4390 57620 4410
rect 57170 4385 57175 4390
rect 57135 4380 57175 4385
rect 57615 4385 57620 4390
rect 57650 4385 57655 4415
rect 57615 4380 57655 4385
rect 52290 4320 61510 4325
rect 52290 4290 52295 4320
rect 52325 4290 52335 4320
rect 52365 4290 52375 4320
rect 52405 4290 52645 4320
rect 52675 4290 52685 4320
rect 52715 4290 52725 4320
rect 52755 4290 52995 4320
rect 53025 4290 53035 4320
rect 53065 4290 53075 4320
rect 53105 4290 53695 4320
rect 53725 4290 53735 4320
rect 53765 4290 53775 4320
rect 53805 4290 54045 4320
rect 54075 4290 54085 4320
rect 54115 4290 54125 4320
rect 54155 4290 54675 4320
rect 54705 4290 55035 4320
rect 55065 4290 55395 4320
rect 55425 4290 55625 4320
rect 55655 4290 55665 4320
rect 55695 4290 55705 4320
rect 55735 4290 56885 4320
rect 56915 4290 58060 4320
rect 58090 4290 58100 4320
rect 58130 4290 58140 4320
rect 58170 4290 58375 4320
rect 58405 4290 58735 4320
rect 58765 4290 59095 4320
rect 59125 4290 59645 4320
rect 59675 4290 59685 4320
rect 59715 4290 59725 4320
rect 59755 4290 59995 4320
rect 60025 4290 60035 4320
rect 60065 4290 60075 4320
rect 60105 4290 60695 4320
rect 60725 4290 60735 4320
rect 60765 4290 60775 4320
rect 60805 4290 61045 4320
rect 61075 4290 61085 4320
rect 61115 4290 61125 4320
rect 61155 4290 61395 4320
rect 61425 4290 61435 4320
rect 61465 4290 61475 4320
rect 61505 4290 61510 4320
rect 52290 4280 61510 4290
rect 52290 4250 52295 4280
rect 52325 4250 52335 4280
rect 52365 4250 52375 4280
rect 52405 4250 52645 4280
rect 52675 4250 52685 4280
rect 52715 4250 52725 4280
rect 52755 4250 52995 4280
rect 53025 4250 53035 4280
rect 53065 4250 53075 4280
rect 53105 4250 53695 4280
rect 53725 4250 53735 4280
rect 53765 4250 53775 4280
rect 53805 4250 54045 4280
rect 54075 4250 54085 4280
rect 54115 4250 54125 4280
rect 54155 4250 54675 4280
rect 54705 4250 55035 4280
rect 55065 4250 55395 4280
rect 55425 4250 55625 4280
rect 55655 4250 55665 4280
rect 55695 4250 55705 4280
rect 55735 4250 56885 4280
rect 56915 4250 58060 4280
rect 58090 4250 58100 4280
rect 58130 4250 58140 4280
rect 58170 4250 58375 4280
rect 58405 4250 58735 4280
rect 58765 4250 59095 4280
rect 59125 4250 59645 4280
rect 59675 4250 59685 4280
rect 59715 4250 59725 4280
rect 59755 4250 59995 4280
rect 60025 4250 60035 4280
rect 60065 4250 60075 4280
rect 60105 4250 60695 4280
rect 60725 4250 60735 4280
rect 60765 4250 60775 4280
rect 60805 4250 61045 4280
rect 61075 4250 61085 4280
rect 61115 4250 61125 4280
rect 61155 4250 61395 4280
rect 61425 4250 61435 4280
rect 61465 4250 61475 4280
rect 61505 4250 61510 4280
rect 52290 4240 61510 4250
rect 52290 4210 52295 4240
rect 52325 4210 52335 4240
rect 52365 4210 52375 4240
rect 52405 4210 52645 4240
rect 52675 4210 52685 4240
rect 52715 4210 52725 4240
rect 52755 4210 52995 4240
rect 53025 4210 53035 4240
rect 53065 4210 53075 4240
rect 53105 4210 53695 4240
rect 53725 4210 53735 4240
rect 53765 4210 53775 4240
rect 53805 4210 54045 4240
rect 54075 4210 54085 4240
rect 54115 4210 54125 4240
rect 54155 4210 54675 4240
rect 54705 4210 55035 4240
rect 55065 4210 55395 4240
rect 55425 4210 55625 4240
rect 55655 4210 55665 4240
rect 55695 4210 55705 4240
rect 55735 4210 56885 4240
rect 56915 4210 58060 4240
rect 58090 4210 58100 4240
rect 58130 4210 58140 4240
rect 58170 4210 58375 4240
rect 58405 4210 58735 4240
rect 58765 4210 59095 4240
rect 59125 4210 59645 4240
rect 59675 4210 59685 4240
rect 59715 4210 59725 4240
rect 59755 4210 59995 4240
rect 60025 4210 60035 4240
rect 60065 4210 60075 4240
rect 60105 4210 60695 4240
rect 60725 4210 60735 4240
rect 60765 4210 60775 4240
rect 60805 4210 61045 4240
rect 61075 4210 61085 4240
rect 61115 4210 61125 4240
rect 61155 4210 61395 4240
rect 61425 4210 61435 4240
rect 61465 4210 61475 4240
rect 61505 4210 61510 4240
rect 52290 4205 61510 4210
rect 54730 4185 56765 4190
rect 54730 4155 54735 4185
rect 54765 4155 54775 4185
rect 54805 4155 54815 4185
rect 54845 4155 54855 4185
rect 54885 4155 54895 4185
rect 54925 4155 54935 4185
rect 54965 4155 54975 4185
rect 55005 4155 55095 4185
rect 55125 4155 55135 4185
rect 55165 4155 55175 4185
rect 55205 4155 55215 4185
rect 55245 4155 55255 4185
rect 55285 4155 55295 4185
rect 55325 4155 55335 4185
rect 55365 4155 56010 4185
rect 56040 4155 56050 4185
rect 56080 4155 56090 4185
rect 56120 4155 56130 4185
rect 56160 4155 56170 4185
rect 56200 4155 56210 4185
rect 56240 4155 56250 4185
rect 56280 4155 56290 4185
rect 56320 4155 56330 4185
rect 56360 4155 56370 4185
rect 56400 4155 56410 4185
rect 56440 4155 56450 4185
rect 56480 4155 56490 4185
rect 56520 4155 56530 4185
rect 56560 4155 56570 4185
rect 56600 4155 56610 4185
rect 56640 4155 56650 4185
rect 56680 4155 56690 4185
rect 56720 4155 56730 4185
rect 56760 4155 56765 4185
rect 54730 4145 56765 4155
rect 54730 4115 54735 4145
rect 54765 4115 54775 4145
rect 54805 4115 54815 4145
rect 54845 4115 54855 4145
rect 54885 4115 54895 4145
rect 54925 4115 54935 4145
rect 54965 4115 54975 4145
rect 55005 4115 55095 4145
rect 55125 4115 55135 4145
rect 55165 4115 55175 4145
rect 55205 4115 55215 4145
rect 55245 4115 55255 4145
rect 55285 4115 55295 4145
rect 55325 4115 55335 4145
rect 55365 4115 56010 4145
rect 56040 4115 56050 4145
rect 56080 4115 56090 4145
rect 56120 4115 56130 4145
rect 56160 4115 56170 4145
rect 56200 4115 56210 4145
rect 56240 4115 56250 4145
rect 56280 4115 56290 4145
rect 56320 4115 56330 4145
rect 56360 4115 56370 4145
rect 56400 4115 56410 4145
rect 56440 4115 56450 4145
rect 56480 4115 56490 4145
rect 56520 4115 56530 4145
rect 56560 4115 56570 4145
rect 56600 4115 56610 4145
rect 56640 4115 56650 4145
rect 56680 4115 56690 4145
rect 56720 4115 56730 4145
rect 56760 4115 56765 4145
rect 54730 4105 56765 4115
rect 54730 4075 54735 4105
rect 54765 4075 54775 4105
rect 54805 4075 54815 4105
rect 54845 4075 54855 4105
rect 54885 4075 54895 4105
rect 54925 4075 54935 4105
rect 54965 4075 54975 4105
rect 55005 4075 55095 4105
rect 55125 4075 55135 4105
rect 55165 4075 55175 4105
rect 55205 4075 55215 4105
rect 55245 4075 55255 4105
rect 55285 4075 55295 4105
rect 55325 4075 55335 4105
rect 55365 4075 56010 4105
rect 56040 4075 56050 4105
rect 56080 4075 56090 4105
rect 56120 4075 56130 4105
rect 56160 4075 56170 4105
rect 56200 4075 56210 4105
rect 56240 4075 56250 4105
rect 56280 4075 56290 4105
rect 56320 4075 56330 4105
rect 56360 4075 56370 4105
rect 56400 4075 56410 4105
rect 56440 4075 56450 4105
rect 56480 4075 56490 4105
rect 56520 4075 56530 4105
rect 56560 4075 56570 4105
rect 56600 4075 56610 4105
rect 56640 4075 56650 4105
rect 56680 4075 56690 4105
rect 56720 4075 56730 4105
rect 56760 4075 56765 4105
rect 54730 4070 56765 4075
rect 57035 4185 59070 4190
rect 57035 4155 57040 4185
rect 57070 4155 57080 4185
rect 57110 4155 57120 4185
rect 57150 4155 57160 4185
rect 57190 4155 57200 4185
rect 57230 4155 57240 4185
rect 57270 4155 57280 4185
rect 57310 4155 57320 4185
rect 57350 4155 57360 4185
rect 57390 4155 57400 4185
rect 57430 4155 57440 4185
rect 57470 4155 57480 4185
rect 57510 4155 57520 4185
rect 57550 4155 57560 4185
rect 57590 4155 57600 4185
rect 57630 4155 57640 4185
rect 57670 4155 57680 4185
rect 57710 4155 57720 4185
rect 57750 4155 57760 4185
rect 57790 4155 58435 4185
rect 58465 4155 58475 4185
rect 58505 4155 58515 4185
rect 58545 4155 58555 4185
rect 58585 4155 58595 4185
rect 58625 4155 58635 4185
rect 58665 4155 58675 4185
rect 58705 4155 58795 4185
rect 58825 4155 58835 4185
rect 58865 4155 58875 4185
rect 58905 4155 58915 4185
rect 58945 4155 58955 4185
rect 58985 4155 58995 4185
rect 59025 4155 59035 4185
rect 59065 4155 59070 4185
rect 57035 4145 59070 4155
rect 57035 4115 57040 4145
rect 57070 4115 57080 4145
rect 57110 4115 57120 4145
rect 57150 4115 57160 4145
rect 57190 4115 57200 4145
rect 57230 4115 57240 4145
rect 57270 4115 57280 4145
rect 57310 4115 57320 4145
rect 57350 4115 57360 4145
rect 57390 4115 57400 4145
rect 57430 4115 57440 4145
rect 57470 4115 57480 4145
rect 57510 4115 57520 4145
rect 57550 4115 57560 4145
rect 57590 4115 57600 4145
rect 57630 4115 57640 4145
rect 57670 4115 57680 4145
rect 57710 4115 57720 4145
rect 57750 4115 57760 4145
rect 57790 4115 58435 4145
rect 58465 4115 58475 4145
rect 58505 4115 58515 4145
rect 58545 4115 58555 4145
rect 58585 4115 58595 4145
rect 58625 4115 58635 4145
rect 58665 4115 58675 4145
rect 58705 4115 58795 4145
rect 58825 4115 58835 4145
rect 58865 4115 58875 4145
rect 58905 4115 58915 4145
rect 58945 4115 58955 4145
rect 58985 4115 58995 4145
rect 59025 4115 59035 4145
rect 59065 4115 59070 4145
rect 57035 4105 59070 4115
rect 57035 4075 57040 4105
rect 57070 4075 57080 4105
rect 57110 4075 57120 4105
rect 57150 4075 57160 4105
rect 57190 4075 57200 4105
rect 57230 4075 57240 4105
rect 57270 4075 57280 4105
rect 57310 4075 57320 4105
rect 57350 4075 57360 4105
rect 57390 4075 57400 4105
rect 57430 4075 57440 4105
rect 57470 4075 57480 4105
rect 57510 4075 57520 4105
rect 57550 4075 57560 4105
rect 57590 4075 57600 4105
rect 57630 4075 57640 4105
rect 57670 4075 57680 4105
rect 57710 4075 57720 4105
rect 57750 4075 57760 4105
rect 57790 4075 58435 4105
rect 58465 4075 58475 4105
rect 58505 4075 58515 4105
rect 58545 4075 58555 4105
rect 58585 4075 58595 4105
rect 58625 4075 58635 4105
rect 58665 4075 58675 4105
rect 58705 4075 58795 4105
rect 58825 4075 58835 4105
rect 58865 4075 58875 4105
rect 58905 4075 58915 4105
rect 58945 4075 58955 4105
rect 58985 4075 58995 4105
rect 59025 4075 59035 4105
rect 59065 4075 59070 4105
rect 57035 4070 59070 4075
rect 54670 4050 54710 4055
rect 54670 4020 54675 4050
rect 54705 4045 54710 4050
rect 54790 4050 54830 4055
rect 54790 4045 54795 4050
rect 54705 4025 54795 4045
rect 54705 4020 54710 4025
rect 54670 4015 54710 4020
rect 54790 4020 54795 4025
rect 54825 4045 54830 4050
rect 54910 4050 54950 4055
rect 54910 4045 54915 4050
rect 54825 4025 54915 4045
rect 54825 4020 54830 4025
rect 54790 4015 54830 4020
rect 54910 4020 54915 4025
rect 54945 4045 54950 4050
rect 55030 4050 55070 4055
rect 55030 4045 55035 4050
rect 54945 4025 55035 4045
rect 54945 4020 54950 4025
rect 54910 4015 54950 4020
rect 55030 4020 55035 4025
rect 55065 4045 55070 4050
rect 55150 4050 55190 4055
rect 55150 4045 55155 4050
rect 55065 4025 55155 4045
rect 55065 4020 55070 4025
rect 55030 4015 55070 4020
rect 55150 4020 55155 4025
rect 55185 4045 55190 4050
rect 55270 4050 55310 4055
rect 55270 4045 55275 4050
rect 55185 4025 55275 4045
rect 55185 4020 55190 4025
rect 55150 4015 55190 4020
rect 55270 4020 55275 4025
rect 55305 4045 55310 4050
rect 55390 4050 55430 4055
rect 55390 4045 55395 4050
rect 55305 4025 55395 4045
rect 55305 4020 55310 4025
rect 55270 4015 55310 4020
rect 55390 4020 55395 4025
rect 55425 4020 55430 4050
rect 55390 4015 55430 4020
rect 56065 4050 56105 4055
rect 56065 4020 56070 4050
rect 56100 4045 56105 4050
rect 56185 4050 56225 4055
rect 56185 4045 56190 4050
rect 56100 4025 56190 4045
rect 56100 4020 56105 4025
rect 56065 4015 56105 4020
rect 56185 4020 56190 4025
rect 56220 4045 56225 4050
rect 56305 4050 56345 4055
rect 56305 4045 56310 4050
rect 56220 4025 56310 4045
rect 56220 4020 56225 4025
rect 56185 4015 56225 4020
rect 56305 4020 56310 4025
rect 56340 4045 56345 4050
rect 56425 4050 56465 4055
rect 56425 4045 56430 4050
rect 56340 4025 56430 4045
rect 56340 4020 56345 4025
rect 56305 4015 56345 4020
rect 56425 4020 56430 4025
rect 56460 4045 56465 4050
rect 56545 4050 56585 4055
rect 56545 4045 56550 4050
rect 56460 4025 56550 4045
rect 56460 4020 56465 4025
rect 56425 4015 56465 4020
rect 56545 4020 56550 4025
rect 56580 4045 56585 4050
rect 56665 4050 56705 4055
rect 56665 4045 56670 4050
rect 56580 4025 56670 4045
rect 56580 4020 56585 4025
rect 56545 4015 56585 4020
rect 56665 4020 56670 4025
rect 56700 4020 56705 4050
rect 56665 4015 56705 4020
rect 57095 4050 57135 4055
rect 57095 4020 57100 4050
rect 57130 4045 57135 4050
rect 57215 4050 57255 4055
rect 57215 4045 57220 4050
rect 57130 4025 57220 4045
rect 57130 4020 57135 4025
rect 57095 4015 57135 4020
rect 57215 4020 57220 4025
rect 57250 4045 57255 4050
rect 57335 4050 57375 4055
rect 57335 4045 57340 4050
rect 57250 4025 57340 4045
rect 57250 4020 57255 4025
rect 57215 4015 57255 4020
rect 57335 4020 57340 4025
rect 57370 4045 57375 4050
rect 57455 4050 57495 4055
rect 57455 4045 57460 4050
rect 57370 4025 57460 4045
rect 57370 4020 57375 4025
rect 57335 4015 57375 4020
rect 57455 4020 57460 4025
rect 57490 4045 57495 4050
rect 57575 4050 57615 4055
rect 57575 4045 57580 4050
rect 57490 4025 57580 4045
rect 57490 4020 57495 4025
rect 57455 4015 57495 4020
rect 57575 4020 57580 4025
rect 57610 4045 57615 4050
rect 57695 4050 57735 4055
rect 57695 4045 57700 4050
rect 57610 4025 57700 4045
rect 57610 4020 57615 4025
rect 57575 4015 57615 4020
rect 57695 4020 57700 4025
rect 57730 4020 57735 4050
rect 57695 4015 57735 4020
rect 58370 4050 58410 4055
rect 58370 4020 58375 4050
rect 58405 4045 58410 4050
rect 58490 4050 58530 4055
rect 58490 4045 58495 4050
rect 58405 4025 58495 4045
rect 58405 4020 58410 4025
rect 58370 4015 58410 4020
rect 58490 4020 58495 4025
rect 58525 4045 58530 4050
rect 58610 4050 58650 4055
rect 58610 4045 58615 4050
rect 58525 4025 58615 4045
rect 58525 4020 58530 4025
rect 58490 4015 58530 4020
rect 58610 4020 58615 4025
rect 58645 4045 58650 4050
rect 58730 4050 58770 4055
rect 58730 4045 58735 4050
rect 58645 4025 58735 4045
rect 58645 4020 58650 4025
rect 58610 4015 58650 4020
rect 58730 4020 58735 4025
rect 58765 4045 58770 4050
rect 58850 4050 58890 4055
rect 58850 4045 58855 4050
rect 58765 4025 58855 4045
rect 58765 4020 58770 4025
rect 58730 4015 58770 4020
rect 58850 4020 58855 4025
rect 58885 4045 58890 4050
rect 58970 4050 59010 4055
rect 58970 4045 58975 4050
rect 58885 4025 58975 4045
rect 58885 4020 58890 4025
rect 58850 4015 58890 4020
rect 58970 4020 58975 4025
rect 59005 4045 59010 4050
rect 59090 4050 59130 4055
rect 59090 4045 59095 4050
rect 59005 4025 59095 4045
rect 59005 4020 59010 4025
rect 58970 4015 59010 4020
rect 59090 4020 59095 4025
rect 59125 4020 59130 4050
rect 59090 4015 59130 4020
rect 54730 3660 54770 3665
rect 54730 3630 54735 3660
rect 54765 3655 54770 3660
rect 54850 3660 54890 3665
rect 54850 3655 54855 3660
rect 54765 3635 54855 3655
rect 54765 3630 54770 3635
rect 54730 3625 54770 3630
rect 54850 3630 54855 3635
rect 54885 3655 54890 3660
rect 54970 3660 55010 3665
rect 54970 3655 54975 3660
rect 54885 3635 54975 3655
rect 54885 3630 54890 3635
rect 54850 3625 54890 3630
rect 54970 3630 54975 3635
rect 55005 3655 55010 3660
rect 55090 3660 55130 3665
rect 55090 3655 55095 3660
rect 55005 3635 55095 3655
rect 55005 3630 55010 3635
rect 54970 3625 55010 3630
rect 55090 3630 55095 3635
rect 55125 3655 55130 3660
rect 55210 3660 55250 3665
rect 55210 3655 55215 3660
rect 55125 3635 55215 3655
rect 55125 3630 55130 3635
rect 55090 3625 55130 3630
rect 55210 3630 55215 3635
rect 55245 3655 55250 3660
rect 55330 3660 55370 3665
rect 55330 3655 55335 3660
rect 55245 3635 55335 3655
rect 55245 3630 55250 3635
rect 55210 3625 55250 3630
rect 55330 3630 55335 3635
rect 55365 3630 55370 3660
rect 55330 3625 55370 3630
rect 56065 3660 56105 3665
rect 56065 3630 56070 3660
rect 56100 3655 56105 3660
rect 56185 3660 56225 3665
rect 56185 3655 56190 3660
rect 56100 3635 56190 3655
rect 56100 3630 56105 3635
rect 56065 3625 56105 3630
rect 56185 3630 56190 3635
rect 56220 3655 56225 3660
rect 56305 3660 56345 3665
rect 56305 3655 56310 3660
rect 56220 3635 56310 3655
rect 56220 3630 56225 3635
rect 56185 3625 56225 3630
rect 56305 3630 56310 3635
rect 56340 3655 56345 3660
rect 56425 3660 56465 3665
rect 56425 3655 56430 3660
rect 56340 3635 56430 3655
rect 56340 3630 56345 3635
rect 56305 3625 56345 3630
rect 56425 3630 56430 3635
rect 56460 3655 56465 3660
rect 56545 3660 56585 3665
rect 56545 3655 56550 3660
rect 56460 3635 56550 3655
rect 56460 3630 56465 3635
rect 56425 3625 56465 3630
rect 56545 3630 56550 3635
rect 56580 3655 56585 3660
rect 56665 3660 56705 3665
rect 56665 3655 56670 3660
rect 56580 3635 56670 3655
rect 56580 3630 56585 3635
rect 56545 3625 56585 3630
rect 56665 3630 56670 3635
rect 56700 3630 56705 3660
rect 56665 3625 56705 3630
rect 57095 3660 57135 3665
rect 57095 3630 57100 3660
rect 57130 3655 57135 3660
rect 57215 3660 57255 3665
rect 57215 3655 57220 3660
rect 57130 3635 57220 3655
rect 57130 3630 57135 3635
rect 57095 3625 57135 3630
rect 57215 3630 57220 3635
rect 57250 3655 57255 3660
rect 57335 3660 57375 3665
rect 57335 3655 57340 3660
rect 57250 3635 57340 3655
rect 57250 3630 57255 3635
rect 57215 3625 57255 3630
rect 57335 3630 57340 3635
rect 57370 3655 57375 3660
rect 57455 3660 57495 3665
rect 57455 3655 57460 3660
rect 57370 3635 57460 3655
rect 57370 3630 57375 3635
rect 57335 3625 57375 3630
rect 57455 3630 57460 3635
rect 57490 3655 57495 3660
rect 57575 3660 57615 3665
rect 57575 3655 57580 3660
rect 57490 3635 57580 3655
rect 57490 3630 57495 3635
rect 57455 3625 57495 3630
rect 57575 3630 57580 3635
rect 57610 3655 57615 3660
rect 57695 3660 57735 3665
rect 57695 3655 57700 3660
rect 57610 3635 57700 3655
rect 57610 3630 57615 3635
rect 57575 3625 57615 3630
rect 57695 3630 57700 3635
rect 57730 3630 57735 3660
rect 57695 3625 57735 3630
rect 58430 3660 58470 3665
rect 58430 3630 58435 3660
rect 58465 3655 58470 3660
rect 58550 3660 58590 3665
rect 58550 3655 58555 3660
rect 58465 3635 58555 3655
rect 58465 3630 58470 3635
rect 58430 3625 58470 3630
rect 58550 3630 58555 3635
rect 58585 3655 58590 3660
rect 58670 3660 58710 3665
rect 58670 3655 58675 3660
rect 58585 3635 58675 3655
rect 58585 3630 58590 3635
rect 58550 3625 58590 3630
rect 58670 3630 58675 3635
rect 58705 3655 58710 3660
rect 58790 3660 58830 3665
rect 58790 3655 58795 3660
rect 58705 3635 58795 3655
rect 58705 3630 58710 3635
rect 58670 3625 58710 3630
rect 58790 3630 58795 3635
rect 58825 3655 58830 3660
rect 58910 3660 58950 3665
rect 58910 3655 58915 3660
rect 58825 3635 58915 3655
rect 58825 3630 58830 3635
rect 58790 3625 58830 3630
rect 58910 3630 58915 3635
rect 58945 3655 58950 3660
rect 59030 3660 59070 3665
rect 59030 3655 59035 3660
rect 58945 3635 59035 3655
rect 58945 3630 58950 3635
rect 58910 3625 58950 3630
rect 59030 3630 59035 3635
rect 59065 3630 59070 3660
rect 59030 3625 59070 3630
rect 56365 3580 56405 3585
rect 56365 3550 56370 3580
rect 56400 3575 56405 3580
rect 56835 3580 56875 3585
rect 56835 3575 56840 3580
rect 56400 3555 56840 3575
rect 56400 3550 56405 3555
rect 56365 3545 56405 3550
rect 56835 3550 56840 3555
rect 56870 3575 56875 3580
rect 57395 3580 57435 3585
rect 57395 3575 57400 3580
rect 56870 3555 57400 3575
rect 56870 3550 56875 3555
rect 56835 3545 56875 3550
rect 57395 3550 57400 3555
rect 57430 3550 57435 3580
rect 57395 3545 57435 3550
rect 55030 3535 55070 3540
rect 55030 3505 55035 3535
rect 55065 3530 55070 3535
rect 56925 3535 56965 3540
rect 56925 3530 56930 3535
rect 55065 3510 56930 3530
rect 55065 3505 55070 3510
rect 55030 3500 55070 3505
rect 56925 3505 56930 3510
rect 56960 3530 56965 3535
rect 58730 3535 58770 3540
rect 58730 3530 58735 3535
rect 56960 3510 58735 3530
rect 56960 3505 56965 3510
rect 56925 3500 56965 3505
rect 58730 3505 58735 3510
rect 58765 3505 58770 3535
rect 58730 3500 58770 3505
rect 55480 3490 56705 3495
rect 55480 3460 55485 3490
rect 55515 3460 55525 3490
rect 55555 3460 55565 3490
rect 55595 3460 56070 3490
rect 56100 3460 56110 3490
rect 56140 3460 56150 3490
rect 56180 3460 56190 3490
rect 56220 3460 56230 3490
rect 56260 3460 56270 3490
rect 56300 3460 56310 3490
rect 56340 3460 56350 3490
rect 56380 3460 56390 3490
rect 56420 3460 56430 3490
rect 56460 3460 56470 3490
rect 56500 3460 56510 3490
rect 56540 3460 56550 3490
rect 56580 3460 56590 3490
rect 56620 3460 56630 3490
rect 56660 3460 56670 3490
rect 56700 3460 56705 3490
rect 55480 3450 56705 3460
rect 55480 3420 55485 3450
rect 55515 3420 55525 3450
rect 55555 3420 55565 3450
rect 55595 3420 56070 3450
rect 56100 3420 56110 3450
rect 56140 3420 56150 3450
rect 56180 3420 56190 3450
rect 56220 3420 56230 3450
rect 56260 3420 56270 3450
rect 56300 3420 56310 3450
rect 56340 3420 56350 3450
rect 56380 3420 56390 3450
rect 56420 3420 56430 3450
rect 56460 3420 56470 3450
rect 56500 3420 56510 3450
rect 56540 3420 56550 3450
rect 56580 3420 56590 3450
rect 56620 3420 56630 3450
rect 56660 3420 56670 3450
rect 56700 3420 56705 3450
rect 55480 3410 56705 3420
rect 55480 3380 55485 3410
rect 55515 3380 55525 3410
rect 55555 3380 55565 3410
rect 55595 3380 56070 3410
rect 56100 3380 56110 3410
rect 56140 3380 56150 3410
rect 56180 3380 56190 3410
rect 56220 3380 56230 3410
rect 56260 3380 56270 3410
rect 56300 3380 56310 3410
rect 56340 3380 56350 3410
rect 56380 3380 56390 3410
rect 56420 3380 56430 3410
rect 56460 3380 56470 3410
rect 56500 3380 56510 3410
rect 56540 3380 56550 3410
rect 56580 3380 56590 3410
rect 56620 3380 56630 3410
rect 56660 3380 56670 3410
rect 56700 3380 56705 3410
rect 54255 3375 54295 3380
rect 55480 3375 56705 3380
rect 57095 3490 58310 3495
rect 57095 3460 57100 3490
rect 57130 3460 57140 3490
rect 57170 3460 57180 3490
rect 57210 3460 57220 3490
rect 57250 3460 57260 3490
rect 57290 3460 57300 3490
rect 57330 3460 57340 3490
rect 57370 3460 57380 3490
rect 57410 3460 57420 3490
rect 57450 3460 57460 3490
rect 57490 3460 57500 3490
rect 57530 3460 57540 3490
rect 57570 3460 57580 3490
rect 57610 3460 57620 3490
rect 57650 3460 57660 3490
rect 57690 3460 57700 3490
rect 57730 3460 58195 3490
rect 58225 3460 58235 3490
rect 58265 3460 58275 3490
rect 58305 3460 58310 3490
rect 57095 3450 58310 3460
rect 57095 3420 57100 3450
rect 57130 3420 57140 3450
rect 57170 3420 57180 3450
rect 57210 3420 57220 3450
rect 57250 3420 57260 3450
rect 57290 3420 57300 3450
rect 57330 3420 57340 3450
rect 57370 3420 57380 3450
rect 57410 3420 57420 3450
rect 57450 3420 57460 3450
rect 57490 3420 57500 3450
rect 57530 3420 57540 3450
rect 57570 3420 57580 3450
rect 57610 3420 57620 3450
rect 57650 3420 57660 3450
rect 57690 3420 57700 3450
rect 57730 3420 58195 3450
rect 58225 3420 58235 3450
rect 58265 3420 58275 3450
rect 58305 3420 58310 3450
rect 57095 3410 58310 3420
rect 57095 3380 57100 3410
rect 57130 3380 57140 3410
rect 57170 3380 57180 3410
rect 57210 3380 57220 3410
rect 57250 3380 57260 3410
rect 57290 3380 57300 3410
rect 57330 3380 57340 3410
rect 57370 3380 57380 3410
rect 57410 3380 57420 3410
rect 57450 3380 57460 3410
rect 57490 3380 57500 3410
rect 57530 3380 57540 3410
rect 57570 3380 57580 3410
rect 57610 3380 57620 3410
rect 57650 3380 57660 3410
rect 57690 3380 57700 3410
rect 57730 3380 58195 3410
rect 58225 3380 58235 3410
rect 58265 3380 58275 3410
rect 58305 3380 58310 3410
rect 57095 3375 58310 3380
rect 59505 3375 59545 3380
rect 54255 3345 54260 3375
rect 54290 3345 54295 3375
rect 54255 3340 54295 3345
rect 54700 3355 55740 3360
rect 54700 3325 54705 3355
rect 54735 3325 54815 3355
rect 54845 3325 54925 3355
rect 54955 3325 55035 3355
rect 55065 3325 55145 3355
rect 55175 3325 55255 3355
rect 55285 3325 55365 3355
rect 55395 3325 55625 3355
rect 55655 3325 55665 3355
rect 55695 3325 55705 3355
rect 55735 3325 55740 3355
rect 57290 3355 59100 3360
rect 57290 3350 58060 3355
rect 54700 3315 55740 3325
rect 54700 3285 54705 3315
rect 54735 3285 54815 3315
rect 54845 3285 54925 3315
rect 54955 3285 55035 3315
rect 55065 3285 55145 3315
rect 55175 3285 55255 3315
rect 55285 3285 55365 3315
rect 55395 3285 55625 3315
rect 55655 3285 55665 3315
rect 55695 3285 55705 3315
rect 55735 3285 55740 3315
rect 54700 3275 55740 3285
rect 54700 3245 54705 3275
rect 54735 3245 54815 3275
rect 54845 3245 54925 3275
rect 54955 3245 55035 3275
rect 55065 3245 55145 3275
rect 55175 3245 55255 3275
rect 55285 3245 55365 3275
rect 55395 3245 55625 3275
rect 55655 3245 55665 3275
rect 55695 3245 55705 3275
rect 55735 3245 55740 3275
rect 54700 3240 55740 3245
rect 56510 3345 58060 3350
rect 56510 3315 56515 3345
rect 56545 3315 56680 3345
rect 56710 3315 56845 3345
rect 56875 3315 56925 3345
rect 56955 3315 57090 3345
rect 57120 3315 57255 3345
rect 57285 3325 58060 3345
rect 58090 3325 58100 3355
rect 58130 3325 58140 3355
rect 58170 3325 58405 3355
rect 58435 3325 58515 3355
rect 58545 3325 58625 3355
rect 58655 3325 58735 3355
rect 58765 3325 58845 3355
rect 58875 3325 58955 3355
rect 58985 3325 59065 3355
rect 59095 3325 59100 3355
rect 59505 3345 59510 3375
rect 59540 3345 59545 3375
rect 59505 3340 59545 3345
rect 57285 3315 59100 3325
rect 56510 3305 58060 3315
rect 56510 3275 56515 3305
rect 56545 3275 56680 3305
rect 56710 3275 56845 3305
rect 56875 3275 56925 3305
rect 56955 3275 57090 3305
rect 57120 3275 57255 3305
rect 57285 3285 58060 3305
rect 58090 3285 58100 3315
rect 58130 3285 58140 3315
rect 58170 3285 58405 3315
rect 58435 3285 58515 3315
rect 58545 3285 58625 3315
rect 58655 3285 58735 3315
rect 58765 3285 58845 3315
rect 58875 3285 58955 3315
rect 58985 3285 59065 3315
rect 59095 3285 59100 3315
rect 57285 3275 59100 3285
rect 56510 3265 58060 3275
rect 56510 3235 56515 3265
rect 56545 3235 56680 3265
rect 56710 3235 56845 3265
rect 56875 3235 56925 3265
rect 56955 3235 57090 3265
rect 57120 3235 57255 3265
rect 57285 3245 58060 3265
rect 58090 3245 58100 3275
rect 58130 3245 58140 3275
rect 58170 3245 58405 3275
rect 58435 3245 58515 3275
rect 58545 3245 58625 3275
rect 58655 3245 58735 3275
rect 58765 3245 58845 3275
rect 58875 3245 58955 3275
rect 58985 3245 59065 3275
rect 59095 3245 59100 3275
rect 57285 3240 59100 3245
rect 57285 3235 57290 3240
rect 56510 3230 57290 3235
rect 56620 3210 56660 3215
rect 54755 3190 54795 3195
rect 54755 3160 54760 3190
rect 54790 3185 54795 3190
rect 54865 3190 54905 3195
rect 54865 3185 54870 3190
rect 54790 3165 54870 3185
rect 54790 3160 54795 3165
rect 54755 3155 54795 3160
rect 54865 3160 54870 3165
rect 54900 3185 54905 3190
rect 54975 3190 55015 3195
rect 54975 3185 54980 3190
rect 54900 3165 54980 3185
rect 54900 3160 54905 3165
rect 54865 3155 54905 3160
rect 54975 3160 54980 3165
rect 55010 3185 55015 3190
rect 55085 3190 55125 3195
rect 55085 3185 55090 3190
rect 55010 3165 55090 3185
rect 55010 3160 55015 3165
rect 54975 3155 55015 3160
rect 55085 3160 55090 3165
rect 55120 3185 55125 3190
rect 55195 3190 55235 3195
rect 55195 3185 55200 3190
rect 55120 3165 55200 3185
rect 55120 3160 55125 3165
rect 55085 3155 55125 3160
rect 55195 3160 55200 3165
rect 55230 3185 55235 3190
rect 55305 3190 55345 3195
rect 55305 3185 55310 3190
rect 55230 3165 55310 3185
rect 55230 3160 55235 3165
rect 55195 3155 55235 3160
rect 55305 3160 55310 3165
rect 55340 3160 55345 3190
rect 56620 3180 56625 3210
rect 56655 3205 56660 3210
rect 56730 3210 56770 3215
rect 56730 3205 56735 3210
rect 56655 3185 56735 3205
rect 56655 3180 56660 3185
rect 56620 3175 56660 3180
rect 56730 3180 56735 3185
rect 56765 3180 56770 3210
rect 56730 3175 56770 3180
rect 57030 3210 57070 3215
rect 57030 3180 57035 3210
rect 57065 3205 57070 3210
rect 57140 3210 57180 3215
rect 57140 3205 57145 3210
rect 57065 3185 57145 3205
rect 57065 3180 57070 3185
rect 57030 3175 57070 3180
rect 57140 3180 57145 3185
rect 57175 3180 57180 3210
rect 57140 3175 57180 3180
rect 58455 3190 58495 3195
rect 55305 3155 55345 3160
rect 58455 3160 58460 3190
rect 58490 3185 58495 3190
rect 58565 3190 58605 3195
rect 58565 3185 58570 3190
rect 58490 3165 58570 3185
rect 58490 3160 58495 3165
rect 58455 3155 58495 3160
rect 58565 3160 58570 3165
rect 58600 3185 58605 3190
rect 58675 3190 58715 3195
rect 58675 3185 58680 3190
rect 58600 3165 58680 3185
rect 58600 3160 58605 3165
rect 58565 3155 58605 3160
rect 58675 3160 58680 3165
rect 58710 3185 58715 3190
rect 58785 3190 58825 3195
rect 58785 3185 58790 3190
rect 58710 3165 58790 3185
rect 58710 3160 58715 3165
rect 58675 3155 58715 3160
rect 58785 3160 58790 3165
rect 58820 3185 58825 3190
rect 58895 3190 58935 3195
rect 58895 3185 58900 3190
rect 58820 3165 58900 3185
rect 58820 3160 58825 3165
rect 58785 3155 58825 3160
rect 58895 3160 58900 3165
rect 58930 3185 58935 3190
rect 59005 3190 59045 3195
rect 59005 3185 59010 3190
rect 58930 3165 59010 3185
rect 58930 3160 58935 3165
rect 58895 3155 58935 3160
rect 59005 3160 59010 3165
rect 59040 3160 59045 3190
rect 59005 3155 59045 3160
rect 56560 2900 56590 2905
rect 56800 2900 56830 2905
rect 56675 2890 56715 2895
rect 56675 2885 56680 2890
rect 56590 2870 56680 2885
rect 56560 2865 56680 2870
rect 56675 2860 56680 2865
rect 56710 2885 56715 2890
rect 56710 2870 56800 2885
rect 57085 2890 57125 2895
rect 57085 2885 57090 2890
rect 56830 2870 57090 2885
rect 56710 2865 57090 2870
rect 56710 2860 56715 2865
rect 56675 2855 56715 2860
rect 57085 2860 57090 2865
rect 57120 2885 57125 2890
rect 57120 2865 57130 2885
rect 57120 2860 57125 2865
rect 57085 2855 57125 2860
rect 56600 2830 56640 2835
rect 56600 2825 56605 2830
rect 56365 2805 56605 2825
rect 56600 2800 56605 2805
rect 56635 2825 56640 2830
rect 57160 2830 57200 2835
rect 57160 2825 57165 2830
rect 56635 2805 57165 2825
rect 56635 2800 56640 2805
rect 56600 2795 56640 2800
rect 57160 2800 57165 2805
rect 57195 2800 57200 2830
rect 57160 2795 57200 2800
rect 55940 2780 55980 2785
rect 55940 2750 55945 2780
rect 55975 2775 55980 2780
rect 56745 2780 56785 2785
rect 56745 2775 56750 2780
rect 55975 2755 56750 2775
rect 55975 2750 55980 2755
rect 55940 2745 55980 2750
rect 56745 2750 56750 2755
rect 56780 2775 56785 2780
rect 57015 2780 57055 2785
rect 57015 2775 57020 2780
rect 56780 2755 57020 2775
rect 56780 2750 56785 2755
rect 56745 2745 56785 2750
rect 57015 2750 57020 2755
rect 57050 2775 57055 2780
rect 57820 2780 57860 2785
rect 57820 2775 57825 2780
rect 57050 2755 57825 2775
rect 57050 2750 57055 2755
rect 57015 2745 57055 2750
rect 57820 2750 57825 2755
rect 57855 2750 57860 2780
rect 57820 2745 57860 2750
rect 56850 2725 56890 2730
rect 56850 2695 56855 2725
rect 56885 2720 56890 2725
rect 56960 2725 57000 2730
rect 56960 2720 56965 2725
rect 56885 2700 56965 2720
rect 56885 2695 56890 2700
rect 56850 2690 56890 2695
rect 56960 2695 56965 2700
rect 56995 2695 57000 2725
rect 56960 2690 57000 2695
rect 56935 2670 56975 2675
rect 56935 2640 56940 2670
rect 56970 2665 56975 2670
rect 57210 2670 57250 2675
rect 57210 2665 57215 2670
rect 56970 2645 57215 2665
rect 56970 2640 56975 2645
rect 56935 2635 56975 2640
rect 57210 2640 57215 2645
rect 57245 2665 57250 2670
rect 57865 2670 57905 2675
rect 57865 2665 57870 2670
rect 57245 2645 57870 2665
rect 57245 2640 57250 2645
rect 57210 2635 57250 2640
rect 57865 2640 57870 2645
rect 57900 2640 57905 2670
rect 57865 2635 57905 2640
rect 56850 2615 56890 2620
rect 56850 2585 56855 2615
rect 56885 2585 56890 2615
rect 56850 2580 56890 2585
rect 54755 2550 54795 2555
rect 54755 2520 54760 2550
rect 54790 2545 54795 2550
rect 54865 2550 54905 2555
rect 54865 2545 54870 2550
rect 54790 2525 54870 2545
rect 54790 2520 54795 2525
rect 54755 2515 54795 2520
rect 54865 2520 54870 2525
rect 54900 2545 54905 2550
rect 54975 2550 55015 2555
rect 54975 2545 54980 2550
rect 54900 2525 54980 2545
rect 54900 2520 54905 2525
rect 54865 2515 54905 2520
rect 54975 2520 54980 2525
rect 55010 2545 55015 2550
rect 55085 2550 55125 2555
rect 55085 2545 55090 2550
rect 55010 2525 55090 2545
rect 55010 2520 55015 2525
rect 54975 2515 55015 2520
rect 55085 2520 55090 2525
rect 55120 2545 55125 2550
rect 55195 2550 55235 2555
rect 55195 2545 55200 2550
rect 55120 2525 55200 2545
rect 55120 2520 55125 2525
rect 55085 2515 55125 2520
rect 55195 2520 55200 2525
rect 55230 2545 55235 2550
rect 55305 2550 55345 2555
rect 55305 2545 55310 2550
rect 55230 2525 55310 2545
rect 55230 2520 55235 2525
rect 55195 2515 55235 2520
rect 55305 2520 55310 2525
rect 55340 2520 55345 2550
rect 55305 2515 55345 2520
rect 58455 2550 58495 2555
rect 58455 2520 58460 2550
rect 58490 2545 58495 2550
rect 58565 2550 58605 2555
rect 58565 2545 58570 2550
rect 58490 2525 58570 2545
rect 58490 2520 58495 2525
rect 58455 2515 58495 2520
rect 58565 2520 58570 2525
rect 58600 2545 58605 2550
rect 58675 2550 58715 2555
rect 58675 2545 58680 2550
rect 58600 2525 58680 2545
rect 58600 2520 58605 2525
rect 58565 2515 58605 2520
rect 58675 2520 58680 2525
rect 58710 2545 58715 2550
rect 58785 2550 58825 2555
rect 58785 2545 58790 2550
rect 58710 2525 58790 2545
rect 58710 2520 58715 2525
rect 58675 2515 58715 2520
rect 58785 2520 58790 2525
rect 58820 2545 58825 2550
rect 58895 2550 58935 2555
rect 58895 2545 58900 2550
rect 58820 2525 58900 2545
rect 58820 2520 58825 2525
rect 58785 2515 58825 2520
rect 58895 2520 58900 2525
rect 58930 2545 58935 2550
rect 59005 2550 59045 2555
rect 59005 2545 59010 2550
rect 58930 2525 59010 2545
rect 58930 2520 58935 2525
rect 58895 2515 58935 2520
rect 59005 2520 59010 2525
rect 59040 2520 59045 2550
rect 59005 2515 59045 2520
rect 54215 2470 56675 2475
rect 54215 2440 54220 2470
rect 54250 2440 54260 2470
rect 54290 2440 54300 2470
rect 54330 2440 55035 2470
rect 55065 2440 55485 2470
rect 55515 2440 55525 2470
rect 55555 2440 55565 2470
rect 55595 2440 56090 2470
rect 56120 2440 56145 2470
rect 56175 2440 56200 2470
rect 56230 2440 56255 2470
rect 56285 2440 56310 2470
rect 56340 2440 56365 2470
rect 56395 2440 56420 2470
rect 56450 2440 56475 2470
rect 56505 2440 56530 2470
rect 56560 2440 56585 2470
rect 56615 2440 56640 2470
rect 56670 2440 56675 2470
rect 54215 2430 56675 2440
rect 54215 2400 54220 2430
rect 54250 2400 54260 2430
rect 54290 2400 54300 2430
rect 54330 2400 55035 2430
rect 55065 2400 55485 2430
rect 55515 2400 55525 2430
rect 55555 2400 55565 2430
rect 55595 2400 56090 2430
rect 56120 2400 56145 2430
rect 56175 2400 56200 2430
rect 56230 2400 56255 2430
rect 56285 2400 56310 2430
rect 56340 2400 56365 2430
rect 56395 2400 56420 2430
rect 56450 2400 56475 2430
rect 56505 2400 56530 2430
rect 56560 2400 56585 2430
rect 56615 2400 56640 2430
rect 56670 2400 56675 2430
rect 54215 2390 56675 2400
rect 54215 2360 54220 2390
rect 54250 2360 54260 2390
rect 54290 2360 54300 2390
rect 54330 2360 55035 2390
rect 55065 2360 55485 2390
rect 55515 2360 55525 2390
rect 55555 2360 55565 2390
rect 55595 2360 56090 2390
rect 56120 2360 56145 2390
rect 56175 2360 56200 2390
rect 56230 2360 56255 2390
rect 56285 2360 56310 2390
rect 56340 2360 56365 2390
rect 56395 2360 56420 2390
rect 56450 2360 56475 2390
rect 56505 2360 56530 2390
rect 56560 2360 56585 2390
rect 56615 2360 56640 2390
rect 56670 2360 56675 2390
rect 54215 2355 56675 2360
rect 57125 2470 59585 2475
rect 57125 2440 57130 2470
rect 57160 2440 57185 2470
rect 57215 2440 57240 2470
rect 57270 2440 57295 2470
rect 57325 2440 57350 2470
rect 57380 2440 57405 2470
rect 57435 2440 57460 2470
rect 57490 2440 57515 2470
rect 57545 2440 57570 2470
rect 57600 2440 57625 2470
rect 57655 2440 57680 2470
rect 57710 2440 58195 2470
rect 58225 2440 58235 2470
rect 58265 2440 58275 2470
rect 58305 2440 58735 2470
rect 58765 2440 59470 2470
rect 59500 2440 59510 2470
rect 59540 2440 59550 2470
rect 59580 2440 59585 2470
rect 57125 2430 59585 2440
rect 57125 2400 57130 2430
rect 57160 2400 57185 2430
rect 57215 2400 57240 2430
rect 57270 2400 57295 2430
rect 57325 2400 57350 2430
rect 57380 2400 57405 2430
rect 57435 2400 57460 2430
rect 57490 2400 57515 2430
rect 57545 2400 57570 2430
rect 57600 2400 57625 2430
rect 57655 2400 57680 2430
rect 57710 2400 58195 2430
rect 58225 2400 58235 2430
rect 58265 2400 58275 2430
rect 58305 2400 58735 2430
rect 58765 2400 59470 2430
rect 59500 2400 59510 2430
rect 59540 2400 59550 2430
rect 59580 2400 59585 2430
rect 57125 2390 59585 2400
rect 57125 2360 57130 2390
rect 57160 2360 57185 2390
rect 57215 2360 57240 2390
rect 57270 2360 57295 2390
rect 57325 2360 57350 2390
rect 57380 2360 57405 2390
rect 57435 2360 57460 2390
rect 57490 2360 57515 2390
rect 57545 2360 57570 2390
rect 57600 2360 57625 2390
rect 57655 2360 57680 2390
rect 57710 2360 58195 2390
rect 58225 2360 58235 2390
rect 58265 2360 58275 2390
rect 58305 2360 58735 2390
rect 58765 2360 59470 2390
rect 59500 2360 59510 2390
rect 59540 2360 59550 2390
rect 59580 2360 59585 2390
rect 57125 2355 59585 2360
rect 54070 2320 55345 2325
rect 54070 2290 54075 2320
rect 54105 2290 54115 2320
rect 54145 2290 54160 2320
rect 54190 2290 54200 2320
rect 54230 2290 54245 2320
rect 54275 2290 54285 2320
rect 54315 2290 54760 2320
rect 54790 2290 54815 2320
rect 54845 2290 54870 2320
rect 54900 2290 54925 2320
rect 54955 2290 54980 2320
rect 55010 2290 55035 2320
rect 55065 2290 55090 2320
rect 55120 2290 55145 2320
rect 55175 2290 55200 2320
rect 55230 2290 55255 2320
rect 55285 2290 55310 2320
rect 55340 2290 55345 2320
rect 58455 2320 59730 2325
rect 54070 2280 55345 2290
rect 54070 2250 54075 2280
rect 54105 2250 54115 2280
rect 54145 2250 54160 2280
rect 54190 2250 54200 2280
rect 54230 2250 54245 2280
rect 54275 2250 54285 2280
rect 54315 2250 54760 2280
rect 54790 2250 54815 2280
rect 54845 2250 54870 2280
rect 54900 2250 54925 2280
rect 54955 2250 54980 2280
rect 55010 2250 55035 2280
rect 55065 2250 55090 2280
rect 55120 2250 55145 2280
rect 55175 2250 55200 2280
rect 55230 2250 55255 2280
rect 55285 2250 55310 2280
rect 55340 2250 55345 2280
rect 54070 2240 55345 2250
rect 54070 2210 54075 2240
rect 54105 2210 54115 2240
rect 54145 2210 54160 2240
rect 54190 2210 54200 2240
rect 54230 2210 54245 2240
rect 54275 2210 54285 2240
rect 54315 2210 54760 2240
rect 54790 2210 54815 2240
rect 54845 2210 54870 2240
rect 54900 2210 54925 2240
rect 54955 2210 54980 2240
rect 55010 2210 55035 2240
rect 55065 2210 55090 2240
rect 55120 2210 55145 2240
rect 55175 2210 55200 2240
rect 55230 2210 55255 2240
rect 55285 2210 55310 2240
rect 55340 2210 55345 2240
rect 54070 2205 55345 2210
rect 56770 2295 58040 2300
rect 56770 2265 56775 2295
rect 56805 2265 56885 2295
rect 56915 2265 56995 2295
rect 57025 2265 57925 2295
rect 57955 2265 57965 2295
rect 57995 2265 58005 2295
rect 58035 2265 58040 2295
rect 56770 2255 58040 2265
rect 56770 2225 56775 2255
rect 56805 2225 56885 2255
rect 56915 2225 56995 2255
rect 57025 2225 57925 2255
rect 57955 2225 57965 2255
rect 57995 2225 58005 2255
rect 58035 2225 58040 2255
rect 56770 2215 58040 2225
rect 54700 2185 55740 2190
rect 54700 2155 54705 2185
rect 54735 2155 55365 2185
rect 55395 2155 55625 2185
rect 55655 2155 55665 2185
rect 55695 2155 55705 2185
rect 55735 2155 55740 2185
rect 56770 2185 56775 2215
rect 56805 2185 56885 2215
rect 56915 2185 56995 2215
rect 57025 2185 57925 2215
rect 57955 2185 57965 2215
rect 57995 2185 58005 2215
rect 58035 2185 58040 2215
rect 58455 2290 58460 2320
rect 58490 2290 58515 2320
rect 58545 2290 58570 2320
rect 58600 2290 58625 2320
rect 58655 2290 58680 2320
rect 58710 2290 58735 2320
rect 58765 2290 58790 2320
rect 58820 2290 58845 2320
rect 58875 2290 58900 2320
rect 58930 2290 58955 2320
rect 58985 2290 59010 2320
rect 59040 2290 59485 2320
rect 59515 2290 59525 2320
rect 59555 2290 59570 2320
rect 59600 2290 59610 2320
rect 59640 2290 59655 2320
rect 59685 2290 59695 2320
rect 59725 2290 59730 2320
rect 58455 2280 59730 2290
rect 58455 2250 58460 2280
rect 58490 2250 58515 2280
rect 58545 2250 58570 2280
rect 58600 2250 58625 2280
rect 58655 2250 58680 2280
rect 58710 2250 58735 2280
rect 58765 2250 58790 2280
rect 58820 2250 58845 2280
rect 58875 2250 58900 2280
rect 58930 2250 58955 2280
rect 58985 2250 59010 2280
rect 59040 2250 59485 2280
rect 59515 2250 59525 2280
rect 59555 2250 59570 2280
rect 59600 2250 59610 2280
rect 59640 2250 59655 2280
rect 59685 2250 59695 2280
rect 59725 2250 59730 2280
rect 58455 2240 59730 2250
rect 58455 2210 58460 2240
rect 58490 2210 58515 2240
rect 58545 2210 58570 2240
rect 58600 2210 58625 2240
rect 58655 2210 58680 2240
rect 58710 2210 58735 2240
rect 58765 2210 58790 2240
rect 58820 2210 58845 2240
rect 58875 2210 58900 2240
rect 58930 2210 58955 2240
rect 58985 2210 59010 2240
rect 59040 2210 59485 2240
rect 59515 2210 59525 2240
rect 59555 2210 59570 2240
rect 59600 2210 59610 2240
rect 59640 2210 59655 2240
rect 59685 2210 59695 2240
rect 59725 2210 59730 2240
rect 58455 2205 59730 2210
rect 56770 2180 58040 2185
rect 58055 2185 59100 2190
rect 54700 2145 55740 2155
rect 54700 2115 54705 2145
rect 54735 2115 55365 2145
rect 55395 2115 55625 2145
rect 55655 2115 55665 2145
rect 55695 2115 55705 2145
rect 55735 2115 55740 2145
rect 54700 2105 55740 2115
rect 54700 2075 54705 2105
rect 54735 2075 55365 2105
rect 55395 2075 55625 2105
rect 55655 2075 55665 2105
rect 55695 2075 55705 2105
rect 55735 2075 55740 2105
rect 54700 2070 55740 2075
rect 58055 2155 58060 2185
rect 58090 2155 58100 2185
rect 58130 2155 58140 2185
rect 58170 2155 58405 2185
rect 58435 2155 59065 2185
rect 59095 2155 59100 2185
rect 58055 2145 59100 2155
rect 58055 2115 58060 2145
rect 58090 2115 58100 2145
rect 58130 2115 58140 2145
rect 58170 2115 58405 2145
rect 58435 2115 59065 2145
rect 59095 2115 59100 2145
rect 58055 2105 59100 2115
rect 58055 2075 58060 2105
rect 58090 2075 58100 2105
rect 58130 2075 58140 2105
rect 58170 2075 58405 2105
rect 58435 2075 59065 2105
rect 59095 2075 59100 2105
rect 58055 2070 59100 2075
rect 53920 2050 55345 2055
rect 53920 2020 53925 2050
rect 53955 2020 53965 2050
rect 53995 2020 54005 2050
rect 54035 2020 54760 2050
rect 54790 2020 54870 2050
rect 54900 2020 54980 2050
rect 55010 2020 55090 2050
rect 55120 2020 55200 2050
rect 55230 2020 55310 2050
rect 55340 2020 55345 2050
rect 53920 2010 55345 2020
rect 53920 1980 53925 2010
rect 53955 1980 53965 2010
rect 53995 1980 54005 2010
rect 54035 1980 54760 2010
rect 54790 1980 54870 2010
rect 54900 1980 54980 2010
rect 55010 1980 55090 2010
rect 55120 1980 55200 2010
rect 55230 1980 55310 2010
rect 55340 1980 55345 2010
rect 57920 2050 59880 2055
rect 57920 2020 57925 2050
rect 57955 2020 57965 2050
rect 57995 2020 58005 2050
rect 58035 2020 58460 2050
rect 58490 2020 58570 2050
rect 58600 2020 58680 2050
rect 58710 2020 58790 2050
rect 58820 2020 58900 2050
rect 58930 2020 59010 2050
rect 59040 2020 59765 2050
rect 59795 2020 59805 2050
rect 59835 2020 59845 2050
rect 59875 2020 59880 2050
rect 57920 2010 59880 2020
rect 53920 1970 55345 1980
rect 53920 1940 53925 1970
rect 53955 1940 53965 1970
rect 53995 1940 54005 1970
rect 54035 1940 54760 1970
rect 54790 1940 54870 1970
rect 54900 1940 54980 1970
rect 55010 1940 55090 1970
rect 55120 1940 55200 1970
rect 55230 1940 55310 1970
rect 55340 1940 55345 1970
rect 55895 1985 55935 1990
rect 55895 1955 55900 1985
rect 55930 1980 55935 1985
rect 55995 1985 56025 1990
rect 55930 1960 55995 1980
rect 55930 1955 55935 1960
rect 55895 1950 55935 1955
rect 56690 1985 56720 1990
rect 55995 1950 56025 1955
rect 56140 1975 56180 1980
rect 56140 1945 56145 1975
rect 56175 1970 56180 1975
rect 56250 1975 56290 1980
rect 56250 1970 56255 1975
rect 56175 1950 56255 1970
rect 56175 1945 56180 1950
rect 56140 1940 56180 1945
rect 56250 1945 56255 1950
rect 56285 1970 56290 1975
rect 56360 1975 56400 1980
rect 56360 1970 56365 1975
rect 56285 1950 56365 1970
rect 56285 1945 56290 1950
rect 56250 1940 56290 1945
rect 56360 1945 56365 1950
rect 56395 1970 56400 1975
rect 56470 1975 56510 1980
rect 56470 1970 56475 1975
rect 56395 1950 56475 1970
rect 56395 1945 56400 1950
rect 56360 1940 56400 1945
rect 56470 1945 56475 1950
rect 56505 1970 56510 1975
rect 56580 1975 56620 1980
rect 56580 1970 56585 1975
rect 56505 1950 56585 1970
rect 56505 1945 56510 1950
rect 56470 1940 56510 1945
rect 56580 1945 56585 1950
rect 56615 1945 56620 1975
rect 57080 1985 57110 1990
rect 56720 1960 57080 1980
rect 56690 1950 56720 1955
rect 57920 1980 57925 2010
rect 57955 1980 57965 2010
rect 57995 1980 58005 2010
rect 58035 1980 58460 2010
rect 58490 1980 58570 2010
rect 58600 1980 58680 2010
rect 58710 1980 58790 2010
rect 58820 1980 58900 2010
rect 58930 1980 59010 2010
rect 59040 1980 59765 2010
rect 59795 1980 59805 2010
rect 59835 1980 59845 2010
rect 59875 1980 59880 2010
rect 57080 1950 57110 1955
rect 57180 1975 57220 1980
rect 56580 1940 56620 1945
rect 57180 1945 57185 1975
rect 57215 1970 57220 1975
rect 57290 1975 57330 1980
rect 57290 1970 57295 1975
rect 57215 1950 57295 1970
rect 57215 1945 57220 1950
rect 57180 1940 57220 1945
rect 57290 1945 57295 1950
rect 57325 1970 57330 1975
rect 57400 1975 57440 1980
rect 57400 1970 57405 1975
rect 57325 1950 57405 1970
rect 57325 1945 57330 1950
rect 57290 1940 57330 1945
rect 57400 1945 57405 1950
rect 57435 1970 57440 1975
rect 57510 1975 57550 1980
rect 57510 1970 57515 1975
rect 57435 1950 57515 1970
rect 57435 1945 57440 1950
rect 57400 1940 57440 1945
rect 57510 1945 57515 1950
rect 57545 1970 57550 1975
rect 57620 1975 57660 1980
rect 57620 1970 57625 1975
rect 57545 1950 57625 1970
rect 57545 1945 57550 1950
rect 57510 1940 57550 1945
rect 57620 1945 57625 1950
rect 57655 1945 57660 1975
rect 57620 1940 57660 1945
rect 57920 1970 59880 1980
rect 57920 1940 57925 1970
rect 57955 1940 57965 1970
rect 57995 1940 58005 1970
rect 58035 1940 58460 1970
rect 58490 1940 58570 1970
rect 58600 1940 58680 1970
rect 58710 1940 58790 1970
rect 58820 1940 58900 1970
rect 58930 1940 59010 1970
rect 59040 1940 59765 1970
rect 59795 1940 59805 1970
rect 59835 1940 59845 1970
rect 59875 1940 59880 1970
rect 53920 1935 55345 1940
rect 57920 1935 59880 1940
rect 54705 1930 54735 1935
rect 56085 1930 56125 1935
rect 54810 1915 54850 1920
rect 54810 1885 54815 1915
rect 54845 1910 54850 1915
rect 54920 1915 54960 1920
rect 54920 1910 54925 1915
rect 54845 1890 54925 1910
rect 54845 1885 54850 1890
rect 54810 1880 54850 1885
rect 54920 1885 54925 1890
rect 54955 1910 54960 1915
rect 55030 1915 55070 1920
rect 55030 1910 55035 1915
rect 54955 1890 55035 1910
rect 54955 1885 54960 1890
rect 54920 1880 54960 1885
rect 55030 1885 55035 1890
rect 55065 1910 55070 1915
rect 55140 1915 55180 1920
rect 55140 1910 55145 1915
rect 55065 1890 55145 1910
rect 55065 1885 55070 1890
rect 55030 1880 55070 1885
rect 55140 1885 55145 1890
rect 55175 1910 55180 1915
rect 55250 1915 55290 1920
rect 55250 1910 55255 1915
rect 55175 1890 55255 1910
rect 55175 1885 55180 1890
rect 55140 1880 55180 1885
rect 55250 1885 55255 1890
rect 55285 1885 55290 1915
rect 56085 1900 56090 1930
rect 56120 1925 56125 1930
rect 56195 1930 56235 1935
rect 56195 1925 56200 1930
rect 56120 1905 56200 1925
rect 56120 1900 56125 1905
rect 56085 1895 56125 1900
rect 56195 1900 56200 1905
rect 56230 1925 56235 1930
rect 56305 1930 56345 1935
rect 56305 1925 56310 1930
rect 56230 1905 56310 1925
rect 56230 1900 56235 1905
rect 56195 1895 56235 1900
rect 56305 1900 56310 1905
rect 56340 1925 56345 1930
rect 56415 1930 56455 1935
rect 56415 1925 56420 1930
rect 56340 1905 56420 1925
rect 56340 1900 56345 1905
rect 56305 1895 56345 1900
rect 56415 1900 56420 1905
rect 56450 1925 56455 1930
rect 56525 1930 56565 1935
rect 56525 1925 56530 1930
rect 56450 1905 56530 1925
rect 56450 1900 56455 1905
rect 56415 1895 56455 1900
rect 56525 1900 56530 1905
rect 56560 1925 56565 1930
rect 56635 1930 56675 1935
rect 56635 1925 56640 1930
rect 56560 1905 56640 1925
rect 56560 1900 56565 1905
rect 56525 1895 56565 1900
rect 56635 1900 56640 1905
rect 56670 1900 56675 1930
rect 56635 1895 56675 1900
rect 57125 1930 57165 1935
rect 57125 1900 57130 1930
rect 57160 1925 57165 1930
rect 57235 1930 57275 1935
rect 57235 1925 57240 1930
rect 57160 1905 57240 1925
rect 57160 1900 57165 1905
rect 57125 1895 57165 1900
rect 57235 1900 57240 1905
rect 57270 1925 57275 1930
rect 57345 1930 57385 1935
rect 57345 1925 57350 1930
rect 57270 1905 57350 1925
rect 57270 1900 57275 1905
rect 57235 1895 57275 1900
rect 57345 1900 57350 1905
rect 57380 1925 57385 1930
rect 57455 1930 57495 1935
rect 57455 1925 57460 1930
rect 57380 1905 57460 1925
rect 57380 1900 57385 1905
rect 57345 1895 57385 1900
rect 57455 1900 57460 1905
rect 57490 1925 57495 1930
rect 57565 1930 57605 1935
rect 57565 1925 57570 1930
rect 57490 1905 57570 1925
rect 57490 1900 57495 1905
rect 57455 1895 57495 1900
rect 57565 1900 57570 1905
rect 57600 1925 57605 1930
rect 57675 1930 57715 1935
rect 58405 1930 58435 1935
rect 59065 1930 59095 1935
rect 57675 1925 57680 1930
rect 57600 1905 57680 1925
rect 57600 1900 57605 1905
rect 57565 1895 57605 1900
rect 57675 1900 57680 1905
rect 57710 1900 57715 1930
rect 57675 1895 57715 1900
rect 58510 1915 58550 1920
rect 55250 1880 55290 1885
rect 58510 1885 58515 1915
rect 58545 1910 58550 1915
rect 58620 1915 58660 1920
rect 58620 1910 58625 1915
rect 58545 1890 58625 1910
rect 58545 1885 58550 1890
rect 58510 1880 58550 1885
rect 58620 1885 58625 1890
rect 58655 1910 58660 1915
rect 58730 1915 58770 1920
rect 58730 1910 58735 1915
rect 58655 1890 58735 1910
rect 58655 1885 58660 1890
rect 58620 1880 58660 1885
rect 58730 1885 58735 1890
rect 58765 1910 58770 1915
rect 58840 1915 58880 1920
rect 58840 1910 58845 1915
rect 58765 1890 58845 1910
rect 58765 1885 58770 1890
rect 58730 1880 58770 1885
rect 58840 1885 58845 1890
rect 58875 1910 58880 1915
rect 58950 1915 58990 1920
rect 58950 1910 58955 1915
rect 58875 1890 58955 1910
rect 58875 1885 58880 1890
rect 58840 1880 58880 1885
rect 58950 1885 58955 1890
rect 58985 1885 58990 1915
rect 58950 1880 58990 1885
rect 56140 1740 56180 1745
rect 54070 1710 54320 1720
rect 54070 1680 54080 1710
rect 54110 1680 54130 1710
rect 54160 1680 54180 1710
rect 54210 1680 54230 1710
rect 54260 1680 54280 1710
rect 54310 1680 54320 1710
rect 56140 1710 56145 1740
rect 56175 1735 56180 1740
rect 56250 1740 56290 1745
rect 56250 1735 56255 1740
rect 56175 1715 56255 1735
rect 56175 1710 56180 1715
rect 56140 1705 56180 1710
rect 56250 1710 56255 1715
rect 56285 1735 56290 1740
rect 56360 1740 56400 1745
rect 56360 1735 56365 1740
rect 56285 1715 56365 1735
rect 56285 1710 56290 1715
rect 56250 1705 56290 1710
rect 56360 1710 56365 1715
rect 56395 1735 56400 1740
rect 56470 1740 56510 1745
rect 56470 1735 56475 1740
rect 56395 1715 56475 1735
rect 56395 1710 56400 1715
rect 56360 1705 56400 1710
rect 56470 1710 56475 1715
rect 56505 1735 56510 1740
rect 56580 1740 56620 1745
rect 56580 1735 56585 1740
rect 56505 1715 56585 1735
rect 56505 1710 56510 1715
rect 56470 1705 56510 1710
rect 56580 1710 56585 1715
rect 56615 1710 56620 1740
rect 56580 1705 56620 1710
rect 57180 1740 57220 1745
rect 57180 1710 57185 1740
rect 57215 1735 57220 1740
rect 57290 1740 57330 1745
rect 57290 1735 57295 1740
rect 57215 1715 57295 1735
rect 57215 1710 57220 1715
rect 57180 1705 57220 1710
rect 57290 1710 57295 1715
rect 57325 1735 57330 1740
rect 57400 1740 57440 1745
rect 57400 1735 57405 1740
rect 57325 1715 57405 1735
rect 57325 1710 57330 1715
rect 57290 1705 57330 1710
rect 57400 1710 57405 1715
rect 57435 1735 57440 1740
rect 57510 1740 57550 1745
rect 57510 1735 57515 1740
rect 57435 1715 57515 1735
rect 57435 1710 57440 1715
rect 57400 1705 57440 1710
rect 57510 1710 57515 1715
rect 57545 1735 57550 1740
rect 57620 1740 57660 1745
rect 57620 1735 57625 1740
rect 57545 1715 57625 1735
rect 57545 1710 57550 1715
rect 57510 1705 57550 1710
rect 57620 1710 57625 1715
rect 57655 1710 57660 1740
rect 57620 1705 57660 1710
rect 59480 1710 59730 1720
rect 54070 1660 54320 1680
rect 56085 1695 56125 1700
rect 56085 1665 56090 1695
rect 56120 1690 56125 1695
rect 56195 1695 56235 1700
rect 56195 1690 56200 1695
rect 56120 1670 56200 1690
rect 56120 1665 56125 1670
rect 54070 1630 54080 1660
rect 54110 1630 54130 1660
rect 54160 1630 54180 1660
rect 54210 1630 54230 1660
rect 54260 1630 54280 1660
rect 54310 1630 54320 1660
rect 54070 1610 54320 1630
rect 54565 1660 54605 1665
rect 54565 1630 54570 1660
rect 54600 1655 54605 1660
rect 54810 1660 54850 1665
rect 54810 1655 54815 1660
rect 54600 1635 54815 1655
rect 54600 1630 54605 1635
rect 54565 1625 54605 1630
rect 54810 1630 54815 1635
rect 54845 1655 54850 1660
rect 54920 1660 54960 1665
rect 54920 1655 54925 1660
rect 54845 1635 54925 1655
rect 54845 1630 54850 1635
rect 54810 1625 54850 1630
rect 54920 1630 54925 1635
rect 54955 1655 54960 1660
rect 55030 1660 55070 1665
rect 55030 1655 55035 1660
rect 54955 1635 55035 1655
rect 54955 1630 54960 1635
rect 54920 1625 54960 1630
rect 55030 1630 55035 1635
rect 55065 1655 55070 1660
rect 55140 1660 55180 1665
rect 55140 1655 55145 1660
rect 55065 1635 55145 1655
rect 55065 1630 55070 1635
rect 55030 1625 55070 1630
rect 55140 1630 55145 1635
rect 55175 1655 55180 1660
rect 55250 1660 55290 1665
rect 56085 1660 56125 1665
rect 56195 1665 56200 1670
rect 56230 1690 56235 1695
rect 56305 1695 56345 1700
rect 56305 1690 56310 1695
rect 56230 1670 56310 1690
rect 56230 1665 56235 1670
rect 56195 1660 56235 1665
rect 56305 1665 56310 1670
rect 56340 1690 56345 1695
rect 56415 1695 56455 1700
rect 56415 1690 56420 1695
rect 56340 1670 56420 1690
rect 56340 1665 56345 1670
rect 56305 1660 56345 1665
rect 56415 1665 56420 1670
rect 56450 1690 56455 1695
rect 56525 1695 56565 1700
rect 56525 1690 56530 1695
rect 56450 1670 56530 1690
rect 56450 1665 56455 1670
rect 56415 1660 56455 1665
rect 56525 1665 56530 1670
rect 56560 1690 56565 1695
rect 56635 1695 56675 1700
rect 56635 1690 56640 1695
rect 56560 1670 56640 1690
rect 56560 1665 56565 1670
rect 56525 1660 56565 1665
rect 56635 1665 56640 1670
rect 56670 1665 56675 1695
rect 56635 1660 56675 1665
rect 57125 1695 57165 1700
rect 57125 1665 57130 1695
rect 57160 1690 57165 1695
rect 57235 1695 57275 1700
rect 57235 1690 57240 1695
rect 57160 1670 57240 1690
rect 57160 1665 57165 1670
rect 57125 1660 57165 1665
rect 57235 1665 57240 1670
rect 57270 1690 57275 1695
rect 57345 1695 57385 1700
rect 57345 1690 57350 1695
rect 57270 1670 57350 1690
rect 57270 1665 57275 1670
rect 57235 1660 57275 1665
rect 57345 1665 57350 1670
rect 57380 1690 57385 1695
rect 57455 1695 57495 1700
rect 57455 1690 57460 1695
rect 57380 1670 57460 1690
rect 57380 1665 57385 1670
rect 57345 1660 57385 1665
rect 57455 1665 57460 1670
rect 57490 1690 57495 1695
rect 57565 1695 57605 1700
rect 57565 1690 57570 1695
rect 57490 1670 57570 1690
rect 57490 1665 57495 1670
rect 57455 1660 57495 1665
rect 57565 1665 57570 1670
rect 57600 1690 57605 1695
rect 57675 1695 57715 1700
rect 57675 1690 57680 1695
rect 57600 1670 57680 1690
rect 57600 1665 57605 1670
rect 57565 1660 57605 1665
rect 57675 1665 57680 1670
rect 57710 1665 57715 1695
rect 59480 1680 59490 1710
rect 59520 1680 59540 1710
rect 59570 1680 59590 1710
rect 59620 1680 59640 1710
rect 59670 1680 59690 1710
rect 59720 1680 59730 1710
rect 57675 1660 57715 1665
rect 58510 1660 58550 1665
rect 55250 1655 55255 1660
rect 55175 1635 55255 1655
rect 55175 1630 55180 1635
rect 55140 1625 55180 1630
rect 55250 1630 55255 1635
rect 55285 1630 55290 1660
rect 55250 1625 55290 1630
rect 56030 1640 58040 1645
rect 54070 1580 54080 1610
rect 54110 1580 54130 1610
rect 54160 1580 54180 1610
rect 54210 1580 54230 1610
rect 54260 1580 54280 1610
rect 54310 1580 54320 1610
rect 56030 1610 56035 1640
rect 56065 1610 56695 1640
rect 56725 1610 57075 1640
rect 57105 1610 57735 1640
rect 57765 1610 57925 1640
rect 57955 1610 57965 1640
rect 57995 1610 58005 1640
rect 58035 1610 58040 1640
rect 58510 1630 58515 1660
rect 58545 1655 58550 1660
rect 58620 1660 58660 1665
rect 58620 1655 58625 1660
rect 58545 1635 58625 1655
rect 58545 1630 58550 1635
rect 58510 1625 58550 1630
rect 58620 1630 58625 1635
rect 58655 1655 58660 1660
rect 58730 1660 58770 1665
rect 58730 1655 58735 1660
rect 58655 1635 58735 1655
rect 58655 1630 58660 1635
rect 58620 1625 58660 1630
rect 58730 1630 58735 1635
rect 58765 1655 58770 1660
rect 58840 1660 58880 1665
rect 58840 1655 58845 1660
rect 58765 1635 58845 1655
rect 58765 1630 58770 1635
rect 58730 1625 58770 1630
rect 58840 1630 58845 1635
rect 58875 1655 58880 1660
rect 58950 1660 58990 1665
rect 58950 1655 58955 1660
rect 58875 1635 58955 1655
rect 58875 1630 58880 1635
rect 58840 1625 58880 1630
rect 58950 1630 58955 1635
rect 58985 1655 58990 1660
rect 59195 1660 59235 1665
rect 59195 1655 59200 1660
rect 58985 1635 59200 1655
rect 58985 1630 58990 1635
rect 58950 1625 58990 1630
rect 59195 1630 59200 1635
rect 59230 1630 59235 1660
rect 59195 1625 59235 1630
rect 59480 1660 59730 1680
rect 59480 1630 59490 1660
rect 59520 1630 59540 1660
rect 59570 1630 59590 1660
rect 59620 1630 59640 1660
rect 59670 1630 59690 1660
rect 59720 1630 59730 1660
rect 56030 1600 58040 1610
rect 59480 1610 59730 1630
rect 54070 1570 54320 1580
rect 55195 1595 55600 1600
rect 55195 1565 55200 1595
rect 55230 1565 55485 1595
rect 55515 1565 55525 1595
rect 55555 1565 55565 1595
rect 55595 1565 55600 1595
rect 55195 1555 55600 1565
rect 55195 1525 55200 1555
rect 55230 1525 55485 1555
rect 55515 1525 55525 1555
rect 55555 1525 55565 1555
rect 55595 1525 55600 1555
rect 56030 1570 56035 1600
rect 56065 1570 56695 1600
rect 56725 1570 57075 1600
rect 57105 1570 57735 1600
rect 57765 1570 57925 1600
rect 57955 1570 57965 1600
rect 57995 1570 58005 1600
rect 58035 1570 58040 1600
rect 56030 1560 58040 1570
rect 56030 1530 56035 1560
rect 56065 1530 56695 1560
rect 56725 1530 57075 1560
rect 57105 1530 57735 1560
rect 57765 1530 57925 1560
rect 57955 1530 57965 1560
rect 57995 1530 58005 1560
rect 58035 1530 58040 1560
rect 56030 1525 58040 1530
rect 58190 1595 58605 1600
rect 58190 1565 58195 1595
rect 58225 1565 58235 1595
rect 58265 1565 58275 1595
rect 58305 1565 58570 1595
rect 58600 1565 58605 1595
rect 59480 1580 59490 1610
rect 59520 1580 59540 1610
rect 59570 1580 59590 1610
rect 59620 1580 59640 1610
rect 59670 1580 59690 1610
rect 59720 1580 59730 1610
rect 59480 1570 59730 1580
rect 58190 1555 58605 1565
rect 58190 1525 58195 1555
rect 58225 1525 58235 1555
rect 58265 1525 58275 1555
rect 58305 1525 58570 1555
rect 58600 1525 58605 1555
rect 55195 1520 55600 1525
rect 58190 1520 58605 1525
rect 55755 1485 58040 1490
rect 54610 1475 54650 1480
rect 54610 1445 54615 1475
rect 54645 1470 54650 1475
rect 54810 1475 54850 1480
rect 54810 1470 54815 1475
rect 54645 1450 54815 1470
rect 54645 1445 54650 1450
rect 54610 1440 54650 1445
rect 54810 1445 54815 1450
rect 54845 1470 54850 1475
rect 54920 1475 54960 1480
rect 54920 1470 54925 1475
rect 54845 1450 54925 1470
rect 54845 1445 54850 1450
rect 54810 1440 54850 1445
rect 54920 1445 54925 1450
rect 54955 1470 54960 1475
rect 55030 1475 55070 1480
rect 55030 1470 55035 1475
rect 54955 1450 55035 1470
rect 54955 1445 54960 1450
rect 54920 1440 54960 1445
rect 55030 1445 55035 1450
rect 55065 1470 55070 1475
rect 55140 1475 55180 1480
rect 55140 1470 55145 1475
rect 55065 1450 55145 1470
rect 55065 1445 55070 1450
rect 55030 1440 55070 1445
rect 55140 1445 55145 1450
rect 55175 1470 55180 1475
rect 55250 1475 55290 1480
rect 55250 1470 55255 1475
rect 55175 1450 55255 1470
rect 55175 1445 55180 1450
rect 55140 1440 55180 1445
rect 55250 1445 55255 1450
rect 55285 1445 55290 1475
rect 55250 1440 55290 1445
rect 55755 1455 55760 1485
rect 55790 1455 55800 1485
rect 55830 1455 55840 1485
rect 55870 1455 56885 1485
rect 56915 1455 57925 1485
rect 57955 1455 57965 1485
rect 57995 1455 58005 1485
rect 58035 1455 58040 1485
rect 55755 1445 58040 1455
rect 55755 1415 55760 1445
rect 55790 1415 55800 1445
rect 55830 1415 55840 1445
rect 55870 1415 56885 1445
rect 56915 1415 57925 1445
rect 57955 1415 57965 1445
rect 57995 1415 58005 1445
rect 58035 1415 58040 1445
rect 58510 1475 58550 1480
rect 58510 1445 58515 1475
rect 58545 1470 58550 1475
rect 58620 1475 58660 1480
rect 58620 1470 58625 1475
rect 58545 1450 58625 1470
rect 58545 1445 58550 1450
rect 58510 1440 58550 1445
rect 58620 1445 58625 1450
rect 58655 1470 58660 1475
rect 58730 1475 58770 1480
rect 58730 1470 58735 1475
rect 58655 1450 58735 1470
rect 58655 1445 58660 1450
rect 58620 1440 58660 1445
rect 58730 1445 58735 1450
rect 58765 1470 58770 1475
rect 58840 1475 58880 1480
rect 58840 1470 58845 1475
rect 58765 1450 58845 1470
rect 58765 1445 58770 1450
rect 58730 1440 58770 1445
rect 58840 1445 58845 1450
rect 58875 1470 58880 1475
rect 58950 1475 58990 1480
rect 58950 1470 58955 1475
rect 58875 1450 58955 1470
rect 58875 1445 58880 1450
rect 58840 1440 58880 1445
rect 58950 1445 58955 1450
rect 58985 1470 58990 1475
rect 59150 1475 59190 1480
rect 59150 1470 59155 1475
rect 58985 1450 59155 1470
rect 58985 1445 58990 1450
rect 58950 1440 58990 1445
rect 59150 1445 59155 1450
rect 59185 1445 59190 1475
rect 59150 1440 59190 1445
rect 55755 1405 58040 1415
rect 55755 1375 55760 1405
rect 55790 1375 55800 1405
rect 55830 1375 55840 1405
rect 55870 1375 56885 1405
rect 56915 1375 57925 1405
rect 57955 1375 57965 1405
rect 57995 1375 58005 1405
rect 58035 1375 58040 1405
rect 55755 1370 58040 1375
rect 56145 1315 56175 1320
rect 56085 1305 56125 1310
rect 56040 1295 56070 1300
rect 56030 1270 56040 1290
rect 56085 1275 56090 1305
rect 56120 1300 56125 1305
rect 56120 1285 56145 1300
rect 56255 1315 56285 1320
rect 56195 1305 56235 1310
rect 56195 1300 56200 1305
rect 56175 1285 56200 1300
rect 56120 1280 56200 1285
rect 56120 1275 56125 1280
rect 56085 1270 56125 1275
rect 56195 1275 56200 1280
rect 56230 1300 56235 1305
rect 56230 1285 56255 1300
rect 56365 1315 56395 1320
rect 56305 1305 56345 1310
rect 56305 1300 56310 1305
rect 56285 1285 56310 1300
rect 56230 1280 56310 1285
rect 56230 1275 56235 1280
rect 56195 1270 56235 1275
rect 56305 1275 56310 1280
rect 56340 1300 56345 1305
rect 56340 1285 56365 1300
rect 56475 1315 56505 1320
rect 56415 1305 56455 1310
rect 56415 1300 56420 1305
rect 56395 1285 56420 1300
rect 56340 1280 56420 1285
rect 56340 1275 56345 1280
rect 56305 1270 56345 1275
rect 56415 1275 56420 1280
rect 56450 1300 56455 1305
rect 56450 1285 56475 1300
rect 56585 1315 56615 1320
rect 56525 1305 56565 1310
rect 56525 1300 56530 1305
rect 56505 1285 56530 1300
rect 56450 1280 56530 1285
rect 56450 1275 56455 1280
rect 56415 1270 56455 1275
rect 56525 1275 56530 1280
rect 56560 1300 56565 1305
rect 56560 1285 56585 1300
rect 57185 1315 57215 1320
rect 56635 1305 56675 1310
rect 56635 1300 56640 1305
rect 56615 1285 56640 1300
rect 56560 1280 56640 1285
rect 56560 1275 56565 1280
rect 56525 1270 56565 1275
rect 56635 1275 56640 1280
rect 56670 1275 56675 1305
rect 56635 1270 56675 1275
rect 56690 1305 56720 1310
rect 56840 1305 56870 1310
rect 56720 1280 56840 1300
rect 56690 1270 56720 1275
rect 56840 1270 56870 1275
rect 56930 1305 56960 1310
rect 57080 1305 57110 1310
rect 56960 1280 57080 1300
rect 56930 1270 56960 1275
rect 57080 1270 57110 1275
rect 57125 1305 57165 1310
rect 57125 1275 57130 1305
rect 57160 1300 57165 1305
rect 57160 1285 57185 1300
rect 57295 1315 57325 1320
rect 57235 1305 57275 1310
rect 57235 1300 57240 1305
rect 57215 1285 57240 1300
rect 57160 1280 57240 1285
rect 57160 1275 57165 1280
rect 57125 1270 57165 1275
rect 57235 1275 57240 1280
rect 57270 1300 57275 1305
rect 57270 1285 57295 1300
rect 57405 1315 57435 1320
rect 57345 1305 57385 1310
rect 57345 1300 57350 1305
rect 57325 1285 57350 1300
rect 57270 1280 57350 1285
rect 57270 1275 57275 1280
rect 57235 1270 57275 1275
rect 57345 1275 57350 1280
rect 57380 1300 57385 1305
rect 57380 1285 57405 1300
rect 57515 1315 57545 1320
rect 57455 1305 57495 1310
rect 57455 1300 57460 1305
rect 57435 1285 57460 1300
rect 57380 1280 57460 1285
rect 57380 1275 57385 1280
rect 57345 1270 57385 1275
rect 57455 1275 57460 1280
rect 57490 1300 57495 1305
rect 57490 1285 57515 1300
rect 57625 1315 57655 1320
rect 57565 1305 57605 1310
rect 57565 1300 57570 1305
rect 57545 1285 57570 1300
rect 57490 1280 57570 1285
rect 57490 1275 57495 1280
rect 57455 1270 57495 1275
rect 57565 1275 57570 1280
rect 57600 1300 57605 1305
rect 57600 1285 57625 1300
rect 57675 1305 57715 1310
rect 57675 1300 57680 1305
rect 57655 1285 57680 1300
rect 57600 1280 57680 1285
rect 57600 1275 57605 1280
rect 57565 1270 57605 1275
rect 57675 1275 57680 1280
rect 57710 1275 57715 1305
rect 57675 1270 57715 1275
rect 57730 1295 57760 1300
rect 57760 1270 57770 1290
rect 56040 1260 56070 1265
rect 56140 1260 56180 1265
rect 56140 1230 56145 1260
rect 56175 1255 56180 1260
rect 56250 1260 56290 1265
rect 56250 1255 56255 1260
rect 56175 1235 56255 1255
rect 56175 1230 56180 1235
rect 56140 1225 56180 1230
rect 56250 1230 56255 1235
rect 56285 1255 56290 1260
rect 56360 1260 56400 1265
rect 56360 1255 56365 1260
rect 56285 1235 56365 1255
rect 56285 1230 56290 1235
rect 56250 1225 56290 1230
rect 56360 1230 56365 1235
rect 56395 1255 56400 1260
rect 56470 1260 56510 1265
rect 56470 1255 56475 1260
rect 56395 1235 56475 1255
rect 56395 1230 56400 1235
rect 56360 1225 56400 1230
rect 56470 1230 56475 1235
rect 56505 1255 56510 1260
rect 56580 1260 56620 1265
rect 56580 1255 56585 1260
rect 56505 1235 56585 1255
rect 56505 1230 56510 1235
rect 56470 1225 56510 1230
rect 56580 1230 56585 1235
rect 56615 1255 56620 1260
rect 57180 1260 57220 1265
rect 57180 1255 57185 1260
rect 56615 1235 57185 1255
rect 56615 1230 56620 1235
rect 56580 1225 56620 1230
rect 57180 1230 57185 1235
rect 57215 1255 57220 1260
rect 57290 1260 57330 1265
rect 57290 1255 57295 1260
rect 57215 1235 57295 1255
rect 57215 1230 57220 1235
rect 57180 1225 57220 1230
rect 57290 1230 57295 1235
rect 57325 1255 57330 1260
rect 57400 1260 57440 1265
rect 57400 1255 57405 1260
rect 57325 1235 57405 1255
rect 57325 1230 57330 1235
rect 57290 1225 57330 1230
rect 57400 1230 57405 1235
rect 57435 1255 57440 1260
rect 57510 1260 57550 1265
rect 57510 1255 57515 1260
rect 57435 1235 57515 1255
rect 57435 1230 57440 1235
rect 57400 1225 57440 1230
rect 57510 1230 57515 1235
rect 57545 1255 57550 1260
rect 57620 1260 57660 1265
rect 57730 1260 57760 1265
rect 57620 1255 57625 1260
rect 57545 1235 57625 1255
rect 57545 1230 57550 1235
rect 57510 1225 57550 1230
rect 57620 1230 57625 1235
rect 57655 1230 57660 1260
rect 57620 1225 57660 1230
rect 54335 1165 54370 1166
rect 59430 1165 59465 1166
rect 54335 1160 54430 1165
rect 54370 1125 54395 1160
rect 54335 1120 54430 1125
rect 54455 1160 54490 1165
rect 54455 1120 54490 1125
rect 54515 1160 54550 1165
rect 59250 1160 59285 1165
rect 54610 1155 54650 1160
rect 54610 1150 54615 1155
rect 54550 1130 54615 1150
rect 54515 1120 54550 1125
rect 54610 1125 54615 1130
rect 54645 1125 54650 1155
rect 59150 1155 59190 1160
rect 54610 1120 54650 1125
rect 54810 1135 54850 1140
rect 54810 1105 54815 1135
rect 54845 1130 54850 1135
rect 54920 1135 54960 1140
rect 54920 1130 54925 1135
rect 54845 1110 54925 1130
rect 54845 1105 54850 1110
rect 54810 1100 54850 1105
rect 54920 1105 54925 1110
rect 54955 1130 54960 1135
rect 55030 1135 55070 1140
rect 55030 1130 55035 1135
rect 54955 1110 55035 1130
rect 54955 1105 54960 1110
rect 54920 1100 54960 1105
rect 55030 1105 55035 1110
rect 55065 1130 55070 1135
rect 55140 1135 55180 1140
rect 55140 1130 55145 1135
rect 55065 1110 55145 1130
rect 55065 1105 55070 1110
rect 55030 1100 55070 1105
rect 55140 1105 55145 1110
rect 55175 1130 55180 1135
rect 55250 1135 55290 1140
rect 55250 1130 55255 1135
rect 55175 1110 55255 1130
rect 55175 1105 55180 1110
rect 55140 1100 55180 1105
rect 55250 1105 55255 1110
rect 55285 1105 55290 1135
rect 55250 1100 55290 1105
rect 58510 1135 58550 1140
rect 58510 1105 58515 1135
rect 58545 1130 58550 1135
rect 58620 1135 58660 1140
rect 58620 1130 58625 1135
rect 58545 1110 58625 1130
rect 58545 1105 58550 1110
rect 58510 1100 58550 1105
rect 58620 1105 58625 1110
rect 58655 1130 58660 1135
rect 58730 1135 58770 1140
rect 58730 1130 58735 1135
rect 58655 1110 58735 1130
rect 58655 1105 58660 1110
rect 58620 1100 58660 1105
rect 58730 1105 58735 1110
rect 58765 1130 58770 1135
rect 58840 1135 58880 1140
rect 58840 1130 58845 1135
rect 58765 1110 58845 1130
rect 58765 1105 58770 1110
rect 58730 1100 58770 1105
rect 58840 1105 58845 1110
rect 58875 1130 58880 1135
rect 58950 1135 58990 1140
rect 58950 1130 58955 1135
rect 58875 1110 58955 1130
rect 58875 1105 58880 1110
rect 58840 1100 58880 1105
rect 58950 1105 58955 1110
rect 58985 1105 58990 1135
rect 59150 1125 59155 1155
rect 59185 1150 59190 1155
rect 59185 1130 59250 1150
rect 59185 1125 59190 1130
rect 59150 1120 59190 1125
rect 59250 1120 59285 1125
rect 59310 1160 59345 1165
rect 59310 1120 59345 1125
rect 59370 1160 59465 1165
rect 59405 1125 59430 1160
rect 59370 1120 59465 1125
rect 58950 1100 58990 1105
rect 54455 1085 54495 1090
rect 54455 1055 54460 1085
rect 54490 1075 54495 1085
rect 54565 1085 54605 1090
rect 59195 1085 59235 1090
rect 54565 1075 54570 1085
rect 54490 1060 54570 1075
rect 54490 1055 54495 1060
rect 54455 1050 54495 1055
rect 54565 1055 54570 1060
rect 54600 1055 54605 1085
rect 58055 1080 59045 1085
rect 54565 1050 54605 1055
rect 54755 1075 55740 1080
rect 54755 1045 54760 1075
rect 54790 1045 54870 1075
rect 54900 1045 54980 1075
rect 55010 1045 55090 1075
rect 55120 1045 55200 1075
rect 55230 1045 55310 1075
rect 55340 1045 55625 1075
rect 55655 1045 55665 1075
rect 55695 1045 55705 1075
rect 55735 1045 55740 1075
rect 54755 1035 55740 1045
rect 54755 1005 54760 1035
rect 54790 1005 54870 1035
rect 54900 1005 54980 1035
rect 55010 1005 55090 1035
rect 55120 1005 55200 1035
rect 55230 1005 55310 1035
rect 55340 1005 55625 1035
rect 55655 1005 55665 1035
rect 55695 1005 55705 1035
rect 55735 1005 55740 1035
rect 56085 1065 56125 1070
rect 56085 1035 56090 1065
rect 56120 1060 56125 1065
rect 56195 1065 56235 1070
rect 56195 1060 56200 1065
rect 56120 1040 56200 1060
rect 56120 1035 56125 1040
rect 56085 1030 56125 1035
rect 56195 1035 56200 1040
rect 56230 1060 56235 1065
rect 56305 1065 56345 1070
rect 56305 1060 56310 1065
rect 56230 1040 56310 1060
rect 56230 1035 56235 1040
rect 56195 1030 56235 1035
rect 56305 1035 56310 1040
rect 56340 1060 56345 1065
rect 56415 1065 56455 1070
rect 56415 1060 56420 1065
rect 56340 1040 56420 1060
rect 56340 1035 56345 1040
rect 56305 1030 56345 1035
rect 56415 1035 56420 1040
rect 56450 1060 56455 1065
rect 56525 1065 56565 1070
rect 56525 1060 56530 1065
rect 56450 1040 56530 1060
rect 56450 1035 56455 1040
rect 56415 1030 56455 1035
rect 56525 1035 56530 1040
rect 56560 1060 56565 1065
rect 56635 1065 56675 1070
rect 56635 1060 56640 1065
rect 56560 1040 56640 1060
rect 56560 1035 56565 1040
rect 56525 1030 56565 1035
rect 56635 1035 56640 1040
rect 56670 1035 56675 1065
rect 56635 1030 56675 1035
rect 56825 1065 56865 1070
rect 56825 1035 56830 1065
rect 56860 1060 56865 1065
rect 56935 1065 56975 1070
rect 56935 1060 56940 1065
rect 56860 1040 56940 1060
rect 56860 1035 56865 1040
rect 56825 1030 56865 1035
rect 56935 1035 56940 1040
rect 56970 1035 56975 1065
rect 56935 1030 56975 1035
rect 57125 1065 57165 1070
rect 57125 1035 57130 1065
rect 57160 1060 57165 1065
rect 57235 1065 57275 1070
rect 57235 1060 57240 1065
rect 57160 1040 57240 1060
rect 57160 1035 57165 1040
rect 57125 1030 57165 1035
rect 57235 1035 57240 1040
rect 57270 1060 57275 1065
rect 57345 1065 57385 1070
rect 57345 1060 57350 1065
rect 57270 1040 57350 1060
rect 57270 1035 57275 1040
rect 57235 1030 57275 1035
rect 57345 1035 57350 1040
rect 57380 1060 57385 1065
rect 57455 1065 57495 1070
rect 57455 1060 57460 1065
rect 57380 1040 57460 1060
rect 57380 1035 57385 1040
rect 57345 1030 57385 1035
rect 57455 1035 57460 1040
rect 57490 1060 57495 1065
rect 57565 1065 57605 1070
rect 57565 1060 57570 1065
rect 57490 1040 57570 1060
rect 57490 1035 57495 1040
rect 57455 1030 57495 1035
rect 57565 1035 57570 1040
rect 57600 1060 57605 1065
rect 57675 1065 57715 1070
rect 57675 1060 57680 1065
rect 57600 1040 57680 1060
rect 57600 1035 57605 1040
rect 57565 1030 57605 1035
rect 57675 1035 57680 1040
rect 57710 1035 57715 1065
rect 57675 1030 57715 1035
rect 58055 1050 58060 1080
rect 58090 1050 58100 1080
rect 58130 1050 58140 1080
rect 58170 1050 58460 1080
rect 58490 1050 58570 1080
rect 58600 1050 58680 1080
rect 58710 1050 58790 1080
rect 58820 1050 58900 1080
rect 58930 1050 59010 1080
rect 59040 1050 59045 1080
rect 59195 1055 59200 1085
rect 59230 1080 59235 1085
rect 59305 1085 59345 1090
rect 59305 1080 59310 1085
rect 59230 1060 59310 1080
rect 59230 1055 59235 1060
rect 59195 1050 59235 1055
rect 59305 1055 59310 1060
rect 59340 1055 59345 1085
rect 59305 1050 59345 1055
rect 58055 1040 59045 1050
rect 54755 995 55740 1005
rect 58055 1010 58060 1040
rect 58090 1010 58100 1040
rect 58130 1010 58140 1040
rect 58170 1010 58460 1040
rect 58490 1010 58570 1040
rect 58600 1010 58680 1040
rect 58710 1010 58790 1040
rect 58820 1010 58900 1040
rect 58930 1010 59010 1040
rect 59040 1010 59045 1040
rect 58055 1000 59045 1010
rect 54755 965 54760 995
rect 54790 965 54870 995
rect 54900 965 54980 995
rect 55010 965 55090 995
rect 55120 965 55200 995
rect 55230 965 55310 995
rect 55340 965 55625 995
rect 55655 965 55665 995
rect 55695 965 55705 995
rect 55735 965 55740 995
rect 54755 960 55740 965
rect 56140 995 57660 1000
rect 56140 965 56145 995
rect 56175 965 56255 995
rect 56285 965 56365 995
rect 56395 965 56475 995
rect 56505 965 56585 995
rect 56615 965 57185 995
rect 57215 965 57295 995
rect 57325 965 57405 995
rect 57435 965 57515 995
rect 57545 965 57625 995
rect 57655 965 57660 995
rect 58055 970 58060 1000
rect 58090 970 58100 1000
rect 58130 970 58140 1000
rect 58170 970 58460 1000
rect 58490 970 58570 1000
rect 58600 970 58680 1000
rect 58710 970 58790 1000
rect 58820 970 58900 1000
rect 58930 970 59010 1000
rect 59040 970 59045 1000
rect 58055 965 59045 970
rect 56140 960 57660 965
rect 53920 940 59880 945
rect 53920 910 53925 940
rect 53955 910 53965 940
rect 53995 910 54005 940
rect 54035 910 54705 940
rect 54735 910 55365 940
rect 55395 910 56035 940
rect 56065 910 56735 940
rect 56765 910 57035 940
rect 57065 910 57735 940
rect 57765 910 58405 940
rect 58435 910 59065 940
rect 59095 910 59765 940
rect 59795 910 59805 940
rect 59835 910 59845 940
rect 59875 910 59880 940
rect 53920 900 59880 910
rect 53920 870 53925 900
rect 53955 870 53965 900
rect 53995 870 54005 900
rect 54035 870 54705 900
rect 54735 870 55365 900
rect 55395 870 56035 900
rect 56065 870 56735 900
rect 56765 870 57035 900
rect 57065 870 57735 900
rect 57765 870 58405 900
rect 58435 870 59065 900
rect 59095 870 59765 900
rect 59795 870 59805 900
rect 59835 870 59845 900
rect 59875 870 59880 900
rect 53920 860 59880 870
rect 53920 830 53925 860
rect 53955 830 53965 860
rect 53995 830 54005 860
rect 54035 830 54705 860
rect 54735 830 55365 860
rect 55395 830 56035 860
rect 56065 830 56735 860
rect 56765 830 57035 860
rect 57065 830 57735 860
rect 57765 830 58405 860
rect 58435 830 59065 860
rect 59095 830 59765 860
rect 59795 830 59805 860
rect 59835 830 59845 860
rect 59875 830 59880 860
rect 53920 825 59880 830
rect 54335 805 54375 810
rect 54335 775 54340 805
rect 54370 800 54375 805
rect 55940 805 55980 810
rect 55940 800 55945 805
rect 54370 780 55945 800
rect 54370 775 54375 780
rect 54335 770 54375 775
rect 55940 775 55945 780
rect 55975 775 55980 805
rect 55940 770 55980 775
rect 57820 805 57860 810
rect 57820 775 57825 805
rect 57855 800 57860 805
rect 59425 805 59465 810
rect 59425 800 59430 805
rect 57855 780 59430 800
rect 57855 775 57860 780
rect 57820 770 57860 775
rect 59425 775 59430 780
rect 59460 775 59465 805
rect 59425 770 59465 775
rect 54400 435 54440 440
rect 54400 405 54405 435
rect 54435 430 54440 435
rect 55080 435 55120 440
rect 55080 430 55085 435
rect 54435 410 55085 430
rect 54435 405 54440 410
rect 54400 400 54440 405
rect 55080 405 55085 410
rect 55115 430 55120 435
rect 58680 435 58720 440
rect 58680 430 58685 435
rect 55115 410 58685 430
rect 55115 405 55120 410
rect 55080 400 55120 405
rect 58680 405 58685 410
rect 58715 430 58720 435
rect 59360 435 59400 440
rect 59360 430 59365 435
rect 58715 410 59365 430
rect 58715 405 58720 410
rect 58680 400 58720 405
rect 59360 405 59365 410
rect 59395 405 59400 435
rect 59360 400 59400 405
rect 56440 390 57470 395
rect 56440 360 56445 390
rect 56475 360 56555 390
rect 56585 360 56665 390
rect 56695 360 56775 390
rect 56805 360 56885 390
rect 56915 360 56995 390
rect 57025 360 57105 390
rect 57135 360 57215 390
rect 57245 360 57325 390
rect 57355 360 57435 390
rect 57465 360 57470 390
rect 56440 355 57470 360
rect 54070 310 55270 315
rect 54070 280 54075 310
rect 54105 280 54115 310
rect 54145 280 54160 310
rect 54190 280 54200 310
rect 54230 280 54245 310
rect 54275 280 54285 310
rect 54315 280 54470 310
rect 54500 280 54835 310
rect 54865 280 54875 310
rect 54905 280 54915 310
rect 54945 280 54955 310
rect 54985 280 54995 310
rect 55025 280 55035 310
rect 55065 280 55075 310
rect 55105 280 55115 310
rect 55145 280 55155 310
rect 55185 280 55195 310
rect 55225 280 55235 310
rect 55265 280 55270 310
rect 54070 270 55270 280
rect 54070 240 54075 270
rect 54105 240 54115 270
rect 54145 240 54160 270
rect 54190 240 54200 270
rect 54230 240 54245 270
rect 54275 240 54285 270
rect 54315 240 54470 270
rect 54500 240 54835 270
rect 54865 240 54875 270
rect 54905 240 54915 270
rect 54945 240 54955 270
rect 54985 240 54995 270
rect 55025 240 55035 270
rect 55065 240 55075 270
rect 55105 240 55115 270
rect 55145 240 55155 270
rect 55185 240 55195 270
rect 55225 240 55235 270
rect 55265 240 55270 270
rect 54070 230 55270 240
rect 54070 200 54075 230
rect 54105 200 54115 230
rect 54145 200 54160 230
rect 54190 200 54200 230
rect 54230 200 54245 230
rect 54275 200 54285 230
rect 54315 200 54470 230
rect 54500 200 54835 230
rect 54865 200 54875 230
rect 54905 200 54915 230
rect 54945 200 54955 230
rect 54985 200 54995 230
rect 55025 200 55035 230
rect 55065 200 55075 230
rect 55105 200 55115 230
rect 55145 200 55155 230
rect 55185 200 55195 230
rect 55225 200 55235 230
rect 55265 200 55270 230
rect 54070 195 55270 200
rect 58530 310 59730 315
rect 58530 280 58535 310
rect 58565 280 58575 310
rect 58605 280 58615 310
rect 58645 280 58655 310
rect 58685 280 58695 310
rect 58725 280 58735 310
rect 58765 280 58775 310
rect 58805 280 58815 310
rect 58845 280 58855 310
rect 58885 280 58895 310
rect 58925 280 58935 310
rect 58965 280 59300 310
rect 59330 280 59485 310
rect 59515 280 59525 310
rect 59555 280 59570 310
rect 59600 280 59610 310
rect 59640 280 59655 310
rect 59685 280 59695 310
rect 59725 280 59730 310
rect 58530 270 59730 280
rect 58530 240 58535 270
rect 58565 240 58575 270
rect 58605 240 58615 270
rect 58645 240 58655 270
rect 58685 240 58695 270
rect 58725 240 58735 270
rect 58765 240 58775 270
rect 58805 240 58815 270
rect 58845 240 58855 270
rect 58885 240 58895 270
rect 58925 240 58935 270
rect 58965 240 59300 270
rect 59330 240 59485 270
rect 59515 240 59525 270
rect 59555 240 59570 270
rect 59600 240 59610 270
rect 59640 240 59655 270
rect 59685 240 59695 270
rect 59725 240 59730 270
rect 58530 230 59730 240
rect 58530 200 58535 230
rect 58565 200 58575 230
rect 58605 200 58615 230
rect 58645 200 58655 230
rect 58685 200 58695 230
rect 58725 200 58735 230
rect 58765 200 58775 230
rect 58805 200 58815 230
rect 58845 200 58855 230
rect 58885 200 58895 230
rect 58925 200 58935 230
rect 58965 200 59300 230
rect 59330 200 59485 230
rect 59515 200 59525 230
rect 59555 200 59570 230
rect 59600 200 59610 230
rect 59640 200 59655 230
rect 59685 200 59695 230
rect 59725 200 59730 230
rect 58530 195 59730 200
rect 54405 175 54440 180
rect 54405 135 54440 140
rect 54465 175 54500 180
rect 54465 135 54500 140
rect 59300 175 59335 180
rect 59300 135 59335 140
rect 59360 175 59395 180
rect 59360 135 59395 140
rect 56220 60 56260 65
rect 56220 30 56225 60
rect 56255 55 56260 60
rect 56275 60 56315 65
rect 56275 55 56280 60
rect 56255 35 56280 55
rect 56255 30 56260 35
rect 56220 25 56260 30
rect 56275 30 56280 35
rect 56310 55 56315 60
rect 56385 60 56425 65
rect 56385 55 56390 60
rect 56310 35 56390 55
rect 56310 30 56315 35
rect 56275 25 56315 30
rect 56385 30 56390 35
rect 56420 55 56425 60
rect 56495 60 56535 65
rect 56495 55 56500 60
rect 56420 35 56500 55
rect 56420 30 56425 35
rect 56385 25 56425 30
rect 56495 30 56500 35
rect 56530 55 56535 60
rect 56605 60 56645 65
rect 56605 55 56610 60
rect 56530 35 56610 55
rect 56530 30 56535 35
rect 56495 25 56535 30
rect 56605 30 56610 35
rect 56640 55 56645 60
rect 56715 60 56755 65
rect 56715 55 56720 60
rect 56640 35 56720 55
rect 56640 30 56645 35
rect 56605 25 56645 30
rect 56715 30 56720 35
rect 56750 55 56755 60
rect 56825 60 56865 65
rect 56825 55 56830 60
rect 56750 35 56830 55
rect 56750 30 56755 35
rect 56715 25 56755 30
rect 56825 30 56830 35
rect 56860 55 56865 60
rect 56935 60 56975 65
rect 56935 55 56940 60
rect 56860 35 56940 55
rect 56860 30 56865 35
rect 56825 25 56865 30
rect 56935 30 56940 35
rect 56970 55 56975 60
rect 57045 60 57085 65
rect 57045 55 57050 60
rect 56970 35 57050 55
rect 56970 30 56975 35
rect 56935 25 56975 30
rect 57045 30 57050 35
rect 57080 55 57085 60
rect 57155 60 57195 65
rect 57155 55 57160 60
rect 57080 35 57160 55
rect 57080 30 57085 35
rect 57045 25 57085 30
rect 57155 30 57160 35
rect 57190 55 57195 60
rect 57265 60 57305 65
rect 57265 55 57270 60
rect 57190 35 57270 55
rect 57190 30 57195 35
rect 57155 25 57195 30
rect 57265 30 57270 35
rect 57300 55 57305 60
rect 57375 60 57415 65
rect 57375 55 57380 60
rect 57300 35 57380 55
rect 57300 30 57305 35
rect 57265 25 57305 30
rect 57375 30 57380 35
rect 57410 55 57415 60
rect 57485 60 57525 65
rect 57485 55 57490 60
rect 57410 35 57490 55
rect 57410 30 57415 35
rect 57375 25 57415 30
rect 57485 30 57490 35
rect 57520 30 57525 60
rect 57485 25 57525 30
rect 56440 15 56480 20
rect 56440 -15 56445 15
rect 56475 10 56480 15
rect 56550 15 56590 20
rect 56550 10 56555 15
rect 56475 -10 56555 10
rect 56475 -15 56480 -10
rect 56440 -20 56480 -15
rect 56550 -15 56555 -10
rect 56585 10 56590 15
rect 56660 15 56700 20
rect 56660 10 56665 15
rect 56585 -10 56665 10
rect 56585 -15 56590 -10
rect 56550 -20 56590 -15
rect 56660 -15 56665 -10
rect 56695 10 56700 15
rect 56770 15 56810 20
rect 56770 10 56775 15
rect 56695 -10 56775 10
rect 56695 -15 56700 -10
rect 56660 -20 56700 -15
rect 56770 -15 56775 -10
rect 56805 10 56810 15
rect 56880 15 56920 20
rect 56880 10 56885 15
rect 56805 -10 56885 10
rect 56805 -15 56810 -10
rect 56770 -20 56810 -15
rect 56880 -15 56885 -10
rect 56915 10 56920 15
rect 56990 15 57030 20
rect 56990 10 56995 15
rect 56915 -10 56995 10
rect 56915 -15 56920 -10
rect 56880 -20 56920 -15
rect 56990 -15 56995 -10
rect 57025 10 57030 15
rect 57100 15 57140 20
rect 57100 10 57105 15
rect 57025 -10 57105 10
rect 57025 -15 57030 -10
rect 56990 -20 57030 -15
rect 57100 -15 57105 -10
rect 57135 10 57140 15
rect 57210 15 57250 20
rect 57210 10 57215 15
rect 57135 -10 57215 10
rect 57135 -15 57140 -10
rect 57100 -20 57140 -15
rect 57210 -15 57215 -10
rect 57245 10 57250 15
rect 57320 15 57360 20
rect 57320 10 57325 15
rect 57245 -10 57325 10
rect 57245 -15 57250 -10
rect 57210 -20 57250 -15
rect 57320 -15 57325 -10
rect 57355 10 57360 15
rect 57430 15 57470 20
rect 57430 10 57435 15
rect 57355 -10 57435 10
rect 57355 -15 57360 -10
rect 57320 -20 57360 -15
rect 57430 -15 57435 -10
rect 57465 -15 57470 15
rect 57430 -20 57470 -15
rect 57415 -40 57455 -35
rect 57415 -70 57420 -40
rect 57450 -45 57455 -40
rect 57865 -40 57905 -35
rect 57865 -45 57870 -40
rect 57450 -65 57870 -45
rect 57450 -70 57455 -65
rect 57415 -75 57455 -70
rect 57865 -70 57870 -65
rect 57900 -70 57905 -40
rect 57865 -75 57905 -70
rect 55755 -95 58040 -90
rect 55755 -125 55760 -95
rect 55790 -125 55800 -95
rect 55830 -125 55840 -95
rect 55870 -125 56335 -95
rect 56365 -125 57925 -95
rect 57955 -125 57965 -95
rect 57995 -125 58005 -95
rect 58035 -125 58040 -95
rect 55755 -135 58040 -125
rect 55755 -165 55760 -135
rect 55790 -165 55800 -135
rect 55830 -165 55840 -135
rect 55870 -165 56335 -135
rect 56365 -165 57925 -135
rect 57955 -165 57965 -135
rect 57995 -165 58005 -135
rect 58035 -165 58040 -135
rect 55755 -175 58040 -165
rect 55755 -205 55760 -175
rect 55790 -205 55800 -175
rect 55830 -205 55840 -175
rect 55870 -205 56335 -175
rect 56365 -205 57925 -175
rect 57955 -205 57965 -175
rect 57995 -205 58005 -175
rect 58035 -205 58040 -175
rect 55755 -210 58040 -205
rect 56540 -230 56580 -225
rect 56540 -260 56545 -230
rect 56575 -235 56580 -230
rect 56650 -230 56690 -225
rect 56650 -235 56655 -230
rect 56575 -255 56655 -235
rect 56575 -260 56580 -255
rect 56540 -265 56580 -260
rect 56650 -260 56655 -255
rect 56685 -235 56690 -230
rect 56870 -230 56910 -225
rect 56870 -235 56875 -230
rect 56685 -255 56875 -235
rect 56685 -260 56690 -255
rect 56650 -265 56690 -260
rect 56870 -260 56875 -255
rect 56905 -260 56910 -230
rect 56870 -265 56910 -260
rect 55895 -275 55935 -270
rect 55895 -305 55900 -275
rect 55930 -280 55935 -275
rect 56485 -275 56525 -270
rect 56485 -280 56490 -275
rect 55930 -300 56490 -280
rect 55930 -305 55935 -300
rect 55895 -310 55935 -305
rect 56485 -305 56490 -300
rect 56520 -280 56525 -275
rect 56595 -275 56635 -270
rect 56595 -280 56600 -275
rect 56520 -300 56600 -280
rect 56520 -305 56525 -300
rect 56485 -310 56525 -305
rect 56595 -305 56600 -300
rect 56630 -280 56635 -275
rect 56705 -275 56745 -270
rect 56705 -280 56710 -275
rect 56630 -300 56710 -280
rect 56630 -305 56635 -300
rect 56595 -310 56635 -305
rect 56705 -305 56710 -300
rect 56740 -280 56745 -275
rect 57040 -275 57080 -270
rect 57040 -280 57045 -275
rect 56740 -300 57045 -280
rect 56740 -305 56745 -300
rect 56705 -310 56745 -305
rect 57040 -305 57045 -300
rect 57075 -305 57080 -275
rect 57040 -310 57080 -305
rect 56540 -480 56580 -475
rect 56540 -510 56545 -480
rect 56575 -485 56580 -480
rect 56650 -480 56690 -475
rect 56650 -485 56655 -480
rect 56575 -505 56655 -485
rect 56575 -510 56580 -505
rect 56540 -515 56580 -510
rect 56650 -510 56655 -505
rect 56685 -485 56690 -480
rect 56870 -480 56910 -475
rect 56870 -485 56875 -480
rect 56685 -505 56875 -485
rect 56685 -510 56690 -505
rect 56650 -515 56690 -510
rect 56870 -510 56875 -505
rect 56905 -510 56910 -480
rect 56870 -515 56910 -510
rect 54830 -525 55270 -520
rect 54830 -555 54835 -525
rect 54865 -555 55035 -525
rect 55065 -555 55235 -525
rect 55265 -555 55270 -525
rect 54830 -560 55270 -555
rect 56485 -525 56525 -520
rect 56485 -555 56490 -525
rect 56520 -530 56525 -525
rect 56595 -525 56635 -520
rect 56595 -530 56600 -525
rect 56520 -550 56600 -530
rect 56520 -555 56525 -550
rect 56485 -560 56525 -555
rect 56595 -555 56600 -550
rect 56630 -530 56635 -525
rect 56705 -525 56745 -520
rect 56705 -530 56710 -525
rect 56630 -550 56710 -530
rect 56630 -555 56635 -550
rect 56595 -560 56635 -555
rect 56705 -555 56710 -550
rect 56740 -555 56745 -525
rect 56705 -560 56745 -555
rect 58530 -525 58970 -520
rect 58530 -555 58535 -525
rect 58565 -555 58735 -525
rect 58765 -555 58935 -525
rect 58965 -555 58970 -525
rect 58530 -560 58970 -555
rect 52290 -580 61510 -575
rect 52290 -610 52295 -580
rect 52325 -610 52335 -580
rect 52365 -610 52375 -580
rect 52405 -610 52645 -580
rect 52675 -610 52685 -580
rect 52715 -610 52725 -580
rect 52755 -610 52995 -580
rect 53025 -610 53035 -580
rect 53065 -610 53075 -580
rect 53105 -610 53345 -580
rect 53375 -610 53385 -580
rect 53415 -610 53425 -580
rect 53455 -610 53695 -580
rect 53725 -610 53735 -580
rect 53765 -610 53775 -580
rect 53805 -610 53925 -580
rect 53955 -610 53965 -580
rect 53995 -610 54005 -580
rect 54035 -610 54045 -580
rect 54075 -610 54085 -580
rect 54115 -610 54125 -580
rect 54155 -610 54395 -580
rect 54425 -610 54435 -580
rect 54465 -610 54475 -580
rect 54505 -610 54745 -580
rect 54775 -610 54785 -580
rect 54815 -610 54825 -580
rect 54855 -610 54935 -580
rect 54965 -610 55095 -580
rect 55125 -610 55135 -580
rect 55165 -610 55175 -580
rect 55205 -610 55325 -580
rect 55355 -610 55365 -580
rect 55395 -610 55405 -580
rect 55435 -610 55445 -580
rect 55475 -610 55485 -580
rect 55515 -610 55525 -580
rect 55555 -610 55795 -580
rect 55825 -610 55835 -580
rect 55865 -610 55875 -580
rect 55905 -610 56145 -580
rect 56175 -610 56185 -580
rect 56215 -610 56225 -580
rect 56255 -610 56435 -580
rect 56465 -610 56495 -580
rect 56525 -610 56535 -580
rect 56565 -610 56575 -580
rect 56605 -610 56765 -580
rect 56795 -610 56845 -580
rect 56875 -610 56885 -580
rect 56915 -610 56925 -580
rect 56955 -610 57195 -580
rect 57225 -610 57235 -580
rect 57265 -610 57275 -580
rect 57305 -610 57490 -580
rect 57520 -610 57545 -580
rect 57575 -610 57585 -580
rect 57615 -610 57625 -580
rect 57655 -610 57895 -580
rect 57925 -610 57935 -580
rect 57965 -610 57975 -580
rect 58005 -610 58245 -580
rect 58275 -610 58285 -580
rect 58315 -610 58325 -580
rect 58355 -610 58365 -580
rect 58395 -610 58405 -580
rect 58435 -610 58445 -580
rect 58475 -610 58595 -580
rect 58625 -610 58635 -580
rect 58665 -610 58675 -580
rect 58705 -610 58835 -580
rect 58865 -610 58945 -580
rect 58975 -610 58985 -580
rect 59015 -610 59025 -580
rect 59055 -610 59295 -580
rect 59325 -610 59335 -580
rect 59365 -610 59375 -580
rect 59405 -610 59645 -580
rect 59675 -610 59685 -580
rect 59715 -610 59725 -580
rect 59755 -610 59765 -580
rect 59795 -610 59805 -580
rect 59835 -610 59845 -580
rect 59875 -610 59995 -580
rect 60025 -610 60035 -580
rect 60065 -610 60075 -580
rect 60105 -610 60345 -580
rect 60375 -610 60385 -580
rect 60415 -610 60425 -580
rect 60455 -610 60695 -580
rect 60725 -610 60735 -580
rect 60765 -610 60775 -580
rect 60805 -610 61045 -580
rect 61075 -610 61085 -580
rect 61115 -610 61125 -580
rect 61155 -610 61395 -580
rect 61425 -610 61435 -580
rect 61465 -610 61475 -580
rect 61505 -610 61510 -580
rect 52290 -620 61510 -610
rect 52290 -650 52295 -620
rect 52325 -650 52335 -620
rect 52365 -650 52375 -620
rect 52405 -650 52645 -620
rect 52675 -650 52685 -620
rect 52715 -650 52725 -620
rect 52755 -650 52995 -620
rect 53025 -650 53035 -620
rect 53065 -650 53075 -620
rect 53105 -650 53345 -620
rect 53375 -650 53385 -620
rect 53415 -650 53425 -620
rect 53455 -650 53695 -620
rect 53725 -650 53735 -620
rect 53765 -650 53775 -620
rect 53805 -650 53925 -620
rect 53955 -650 53965 -620
rect 53995 -650 54005 -620
rect 54035 -650 54045 -620
rect 54075 -650 54085 -620
rect 54115 -650 54125 -620
rect 54155 -650 54395 -620
rect 54425 -650 54435 -620
rect 54465 -650 54475 -620
rect 54505 -650 54745 -620
rect 54775 -650 54785 -620
rect 54815 -650 54825 -620
rect 54855 -650 54935 -620
rect 54965 -650 55095 -620
rect 55125 -650 55135 -620
rect 55165 -650 55175 -620
rect 55205 -650 55325 -620
rect 55355 -650 55365 -620
rect 55395 -650 55405 -620
rect 55435 -650 55445 -620
rect 55475 -650 55485 -620
rect 55515 -650 55525 -620
rect 55555 -650 55795 -620
rect 55825 -650 55835 -620
rect 55865 -650 55875 -620
rect 55905 -650 56145 -620
rect 56175 -650 56185 -620
rect 56215 -650 56225 -620
rect 56255 -650 56435 -620
rect 56465 -650 56495 -620
rect 56525 -650 56535 -620
rect 56565 -650 56575 -620
rect 56605 -650 56765 -620
rect 56795 -650 56845 -620
rect 56875 -650 56885 -620
rect 56915 -650 56925 -620
rect 56955 -650 57195 -620
rect 57225 -650 57235 -620
rect 57265 -650 57275 -620
rect 57305 -650 57490 -620
rect 57520 -650 57545 -620
rect 57575 -650 57585 -620
rect 57615 -650 57625 -620
rect 57655 -650 57895 -620
rect 57925 -650 57935 -620
rect 57965 -650 57975 -620
rect 58005 -650 58245 -620
rect 58275 -650 58285 -620
rect 58315 -650 58325 -620
rect 58355 -650 58365 -620
rect 58395 -650 58405 -620
rect 58435 -650 58445 -620
rect 58475 -650 58595 -620
rect 58625 -650 58635 -620
rect 58665 -650 58675 -620
rect 58705 -650 58835 -620
rect 58865 -650 58945 -620
rect 58975 -650 58985 -620
rect 59015 -650 59025 -620
rect 59055 -650 59295 -620
rect 59325 -650 59335 -620
rect 59365 -650 59375 -620
rect 59405 -650 59645 -620
rect 59675 -650 59685 -620
rect 59715 -650 59725 -620
rect 59755 -650 59765 -620
rect 59795 -650 59805 -620
rect 59835 -650 59845 -620
rect 59875 -650 59995 -620
rect 60025 -650 60035 -620
rect 60065 -650 60075 -620
rect 60105 -650 60345 -620
rect 60375 -650 60385 -620
rect 60415 -650 60425 -620
rect 60455 -650 60695 -620
rect 60725 -650 60735 -620
rect 60765 -650 60775 -620
rect 60805 -650 61045 -620
rect 61075 -650 61085 -620
rect 61115 -650 61125 -620
rect 61155 -650 61395 -620
rect 61425 -650 61435 -620
rect 61465 -650 61475 -620
rect 61505 -650 61510 -620
rect 52290 -660 61510 -650
rect 52290 -690 52295 -660
rect 52325 -690 52335 -660
rect 52365 -690 52375 -660
rect 52405 -690 52645 -660
rect 52675 -690 52685 -660
rect 52715 -690 52725 -660
rect 52755 -690 52995 -660
rect 53025 -690 53035 -660
rect 53065 -690 53075 -660
rect 53105 -690 53345 -660
rect 53375 -690 53385 -660
rect 53415 -690 53425 -660
rect 53455 -690 53695 -660
rect 53725 -690 53735 -660
rect 53765 -690 53775 -660
rect 53805 -690 53925 -660
rect 53955 -690 53965 -660
rect 53995 -690 54005 -660
rect 54035 -690 54045 -660
rect 54075 -690 54085 -660
rect 54115 -690 54125 -660
rect 54155 -690 54395 -660
rect 54425 -690 54435 -660
rect 54465 -690 54475 -660
rect 54505 -690 54745 -660
rect 54775 -690 54785 -660
rect 54815 -690 54825 -660
rect 54855 -690 54935 -660
rect 54965 -690 55095 -660
rect 55125 -690 55135 -660
rect 55165 -690 55175 -660
rect 55205 -690 55325 -660
rect 55355 -690 55365 -660
rect 55395 -690 55405 -660
rect 55435 -690 55445 -660
rect 55475 -690 55485 -660
rect 55515 -690 55525 -660
rect 55555 -690 55795 -660
rect 55825 -690 55835 -660
rect 55865 -690 55875 -660
rect 55905 -690 56145 -660
rect 56175 -690 56185 -660
rect 56215 -690 56225 -660
rect 56255 -690 56435 -660
rect 56465 -690 56495 -660
rect 56525 -690 56535 -660
rect 56565 -690 56575 -660
rect 56605 -690 56765 -660
rect 56795 -690 56845 -660
rect 56875 -690 56885 -660
rect 56915 -690 56925 -660
rect 56955 -690 57195 -660
rect 57225 -690 57235 -660
rect 57265 -690 57275 -660
rect 57305 -690 57490 -660
rect 57520 -690 57545 -660
rect 57575 -690 57585 -660
rect 57615 -690 57625 -660
rect 57655 -690 57895 -660
rect 57925 -690 57935 -660
rect 57965 -690 57975 -660
rect 58005 -690 58245 -660
rect 58275 -690 58285 -660
rect 58315 -690 58325 -660
rect 58355 -690 58365 -660
rect 58395 -690 58405 -660
rect 58435 -690 58445 -660
rect 58475 -690 58595 -660
rect 58625 -690 58635 -660
rect 58665 -690 58675 -660
rect 58705 -690 58835 -660
rect 58865 -690 58945 -660
rect 58975 -690 58985 -660
rect 59015 -690 59025 -660
rect 59055 -690 59295 -660
rect 59325 -690 59335 -660
rect 59365 -690 59375 -660
rect 59405 -690 59645 -660
rect 59675 -690 59685 -660
rect 59715 -690 59725 -660
rect 59755 -690 59765 -660
rect 59795 -690 59805 -660
rect 59835 -690 59845 -660
rect 59875 -690 59995 -660
rect 60025 -690 60035 -660
rect 60065 -690 60075 -660
rect 60105 -690 60345 -660
rect 60375 -690 60385 -660
rect 60415 -690 60425 -660
rect 60455 -690 60695 -660
rect 60725 -690 60735 -660
rect 60765 -690 60775 -660
rect 60805 -690 61045 -660
rect 61075 -690 61085 -660
rect 61115 -690 61125 -660
rect 61155 -690 61395 -660
rect 61425 -690 61435 -660
rect 61465 -690 61475 -660
rect 61505 -690 61510 -660
rect 52290 -695 61510 -690
<< via2 >>
rect 54260 3345 54290 3375
rect 59510 3345 59540 3375
rect 54080 1680 54110 1710
rect 54130 1680 54160 1710
rect 54180 1680 54210 1710
rect 54230 1680 54260 1710
rect 54280 1680 54310 1710
rect 54080 1630 54110 1660
rect 54130 1630 54160 1660
rect 54180 1630 54210 1660
rect 54230 1630 54260 1660
rect 54280 1630 54310 1660
rect 59490 1680 59520 1710
rect 59540 1680 59570 1710
rect 59590 1680 59620 1710
rect 59640 1680 59670 1710
rect 59690 1680 59720 1710
rect 54080 1580 54110 1610
rect 54130 1580 54160 1610
rect 54180 1580 54210 1610
rect 54230 1580 54260 1610
rect 54280 1580 54310 1610
rect 59490 1630 59520 1660
rect 59540 1630 59570 1660
rect 59590 1630 59620 1660
rect 59640 1630 59670 1660
rect 59690 1630 59720 1660
rect 59490 1580 59520 1610
rect 59540 1580 59570 1610
rect 59590 1580 59620 1610
rect 59640 1580 59670 1610
rect 59690 1580 59720 1610
<< metal3 >>
rect 52060 5520 52290 5605
rect 52410 5520 52640 5605
rect 52760 5520 52990 5605
rect 53110 5520 53340 5605
rect 53460 5520 53690 5605
rect 53810 5520 54040 5605
rect 54160 5520 54390 5605
rect 54510 5520 54740 5605
rect 54860 5520 55090 5605
rect 55210 5520 55440 5605
rect 55560 5520 55790 5605
rect 55910 5520 56140 5605
rect 56260 5520 56490 5605
rect 56610 5520 56840 5605
rect 52060 5470 56840 5520
rect 52060 5375 52290 5470
rect 52410 5375 52640 5470
rect 52760 5375 52990 5470
rect 53110 5375 53340 5470
rect 53460 5375 53690 5470
rect 53810 5375 54040 5470
rect 54160 5375 54390 5470
rect 54510 5375 54740 5470
rect 54860 5375 55090 5470
rect 55210 5375 55440 5470
rect 55560 5375 55790 5470
rect 55910 5375 56140 5470
rect 56260 5375 56490 5470
rect 56610 5375 56840 5470
rect 56960 5520 57190 5605
rect 57310 5520 57540 5605
rect 57660 5520 57890 5605
rect 58010 5520 58240 5605
rect 58360 5520 58590 5605
rect 58710 5520 58940 5605
rect 59060 5520 59290 5605
rect 59410 5520 59640 5605
rect 59760 5520 59990 5605
rect 60110 5520 60340 5605
rect 60460 5520 60690 5605
rect 60810 5520 61040 5605
rect 61160 5520 61390 5605
rect 61510 5520 61740 5605
rect 56960 5470 61740 5520
rect 56960 5375 57190 5470
rect 57310 5375 57540 5470
rect 57660 5375 57890 5470
rect 58010 5375 58240 5470
rect 58360 5375 58590 5470
rect 58710 5375 58940 5470
rect 59060 5375 59290 5470
rect 59410 5375 59640 5470
rect 59760 5375 59990 5470
rect 60110 5375 60340 5470
rect 60460 5375 60690 5470
rect 60810 5375 61040 5470
rect 61160 5375 61390 5470
rect 61510 5375 61740 5470
rect 52850 5255 52900 5375
rect 53900 5255 53950 5375
rect 54250 5255 54300 5375
rect 54600 5255 54650 5375
rect 54950 5255 55000 5375
rect 55300 5255 55350 5375
rect 55650 5255 55700 5375
rect 58100 5255 58150 5375
rect 58450 5255 58500 5375
rect 58800 5255 58850 5375
rect 59150 5255 59200 5375
rect 59500 5255 59550 5375
rect 59850 5255 59900 5375
rect 60900 5255 60950 5375
rect 52060 5170 52290 5255
rect 52410 5170 52640 5255
rect 52760 5170 52990 5255
rect 53110 5170 53340 5255
rect 53460 5170 53690 5255
rect 52060 5120 53690 5170
rect 52060 5025 52290 5120
rect 52410 5025 52640 5120
rect 52760 5025 52990 5120
rect 53110 5025 53340 5120
rect 53460 5025 53690 5120
rect 53810 5025 54040 5255
rect 54160 5025 54390 5255
rect 54510 5025 54740 5255
rect 54860 5025 55090 5255
rect 55210 5025 55440 5255
rect 55560 5025 55790 5255
rect 58010 5025 58240 5255
rect 58360 5025 58590 5255
rect 58710 5025 58940 5255
rect 59060 5025 59290 5255
rect 59410 5025 59640 5255
rect 59760 5025 59990 5255
rect 60110 5170 60340 5255
rect 60460 5170 60690 5255
rect 60810 5170 61040 5255
rect 61160 5170 61390 5255
rect 61510 5170 61740 5255
rect 60110 5120 61740 5170
rect 60110 5025 60340 5120
rect 60460 5025 60690 5120
rect 60810 5025 61040 5120
rect 61160 5025 61390 5120
rect 61510 5025 61740 5120
rect 52850 4905 52900 5025
rect 53900 4905 53950 5025
rect 54250 4905 54300 5025
rect 54600 4905 54650 5025
rect 54950 4905 55000 5025
rect 55300 4905 55350 5025
rect 58450 4905 58500 5025
rect 58800 4905 58850 5025
rect 59150 4905 59200 5025
rect 59500 4905 59550 5025
rect 59850 4905 59900 5025
rect 60900 4905 60950 5025
rect 52060 4820 52290 4905
rect 52410 4820 52640 4905
rect 52760 4820 52990 4905
rect 53110 4820 53340 4905
rect 53460 4820 53690 4905
rect 52060 4770 53690 4820
rect 52060 4675 52290 4770
rect 52410 4675 52640 4770
rect 52760 4675 52990 4770
rect 53110 4675 53340 4770
rect 53460 4675 53690 4770
rect 53810 4675 54040 4905
rect 54160 4675 54390 4905
rect 54510 4675 54740 4905
rect 54860 4675 55090 4905
rect 55210 4675 55440 4905
rect 58360 4675 58590 4905
rect 58710 4675 58940 4905
rect 59060 4675 59290 4905
rect 59410 4675 59640 4905
rect 59760 4675 59990 4905
rect 60110 4820 60340 4905
rect 60460 4820 60690 4905
rect 60810 4820 61040 4905
rect 61160 4820 61390 4905
rect 61510 4820 61740 4905
rect 60110 4770 61740 4820
rect 60110 4675 60340 4770
rect 60460 4675 60690 4770
rect 60810 4675 61040 4770
rect 61160 4675 61390 4770
rect 61510 4675 61740 4770
rect 52850 4555 52900 4675
rect 52060 4470 52290 4555
rect 52410 4470 52640 4555
rect 52760 4470 52990 4555
rect 53110 4470 53340 4555
rect 53460 4470 53690 4555
rect 52060 4420 53690 4470
rect 52060 4325 52290 4420
rect 52410 4325 52640 4420
rect 52760 4325 52990 4420
rect 53110 4325 53340 4420
rect 53460 4325 53690 4420
rect 52850 4205 52900 4325
rect 52060 4120 52290 4205
rect 52410 4120 52640 4205
rect 52760 4120 52990 4205
rect 53110 4120 53340 4205
rect 53460 4120 53690 4205
rect 52060 4070 53690 4120
rect 52060 3975 52290 4070
rect 52410 3975 52640 4070
rect 52760 3975 52990 4070
rect 53110 3975 53340 4070
rect 53460 3975 53690 4070
rect 52850 3855 52900 3975
rect 52060 3770 52290 3855
rect 52410 3770 52640 3855
rect 52760 3770 52990 3855
rect 53110 3770 53340 3855
rect 53460 3770 53690 3855
rect 52060 3720 53690 3770
rect 52060 3625 52290 3720
rect 52410 3625 52640 3720
rect 52760 3625 52990 3720
rect 53110 3625 53340 3720
rect 53460 3625 53690 3720
rect 52850 3505 52900 3625
rect 52060 3420 52290 3505
rect 52410 3420 52640 3505
rect 52760 3420 52990 3505
rect 53110 3420 53340 3505
rect 53460 3420 53690 3505
rect 52060 3370 53690 3420
rect 52060 3275 52290 3370
rect 52410 3275 52640 3370
rect 52760 3275 52990 3370
rect 53110 3275 53340 3370
rect 53460 3275 53690 3370
rect 54255 3375 54295 4675
rect 54255 3345 54260 3375
rect 54290 3345 54295 3375
rect 54255 3340 54295 3345
rect 59505 3375 59545 4675
rect 60900 4555 60950 4675
rect 60110 4470 60340 4555
rect 60460 4470 60690 4555
rect 60810 4470 61040 4555
rect 61160 4470 61390 4555
rect 61510 4470 61740 4555
rect 60110 4420 61740 4470
rect 60110 4325 60340 4420
rect 60460 4325 60690 4420
rect 60810 4325 61040 4420
rect 61160 4325 61390 4420
rect 61510 4325 61740 4420
rect 60900 4205 60950 4325
rect 60110 4120 60340 4205
rect 60460 4120 60690 4205
rect 60810 4120 61040 4205
rect 61160 4120 61390 4205
rect 61510 4120 61740 4205
rect 60110 4070 61740 4120
rect 60110 3975 60340 4070
rect 60460 3975 60690 4070
rect 60810 3975 61040 4070
rect 61160 3975 61390 4070
rect 61510 3975 61740 4070
rect 60900 3855 60950 3975
rect 60110 3770 60340 3855
rect 60460 3770 60690 3855
rect 60810 3770 61040 3855
rect 61160 3770 61390 3855
rect 61510 3770 61740 3855
rect 60110 3720 61740 3770
rect 60110 3625 60340 3720
rect 60460 3625 60690 3720
rect 60810 3625 61040 3720
rect 61160 3625 61390 3720
rect 61510 3625 61740 3720
rect 60900 3505 60950 3625
rect 59505 3345 59510 3375
rect 59540 3345 59545 3375
rect 59505 3340 59545 3345
rect 60110 3420 60340 3505
rect 60460 3420 60690 3505
rect 60810 3420 61040 3505
rect 61160 3420 61390 3505
rect 61510 3420 61740 3505
rect 60110 3370 61740 3420
rect 60110 3275 60340 3370
rect 60460 3275 60690 3370
rect 60810 3275 61040 3370
rect 61160 3275 61390 3370
rect 61510 3275 61740 3370
rect 52850 3155 52900 3275
rect 60900 3155 60950 3275
rect 52060 3070 52290 3155
rect 52410 3070 52640 3155
rect 52760 3070 52990 3155
rect 53110 3070 53340 3155
rect 53460 3070 53690 3155
rect 52060 3020 53690 3070
rect 52060 2925 52290 3020
rect 52410 2925 52640 3020
rect 52760 2925 52990 3020
rect 53110 2925 53340 3020
rect 53460 2925 53690 3020
rect 60110 3070 60340 3155
rect 60460 3070 60690 3155
rect 60810 3070 61040 3155
rect 61160 3070 61390 3155
rect 61510 3070 61740 3155
rect 60110 3020 61740 3070
rect 60110 2925 60340 3020
rect 60460 2925 60690 3020
rect 60810 2925 61040 3020
rect 61160 2925 61390 3020
rect 61510 2925 61740 3020
rect 52850 2805 52900 2925
rect 60900 2805 60950 2925
rect 52060 2720 52290 2805
rect 52410 2720 52640 2805
rect 52760 2720 52990 2805
rect 53110 2720 53340 2805
rect 53460 2720 53690 2805
rect 52060 2670 53690 2720
rect 52060 2575 52290 2670
rect 52410 2575 52640 2670
rect 52760 2575 52990 2670
rect 53110 2575 53340 2670
rect 53460 2575 53690 2670
rect 60110 2720 60340 2805
rect 60460 2720 60690 2805
rect 60810 2720 61040 2805
rect 61160 2720 61390 2805
rect 61510 2720 61740 2805
rect 60110 2670 61740 2720
rect 60110 2575 60340 2670
rect 60460 2575 60690 2670
rect 60810 2575 61040 2670
rect 61160 2575 61390 2670
rect 61510 2575 61740 2670
rect 52850 2455 52900 2575
rect 60900 2455 60950 2575
rect 52060 2370 52290 2455
rect 52410 2370 52640 2455
rect 52760 2370 52990 2455
rect 53110 2370 53340 2455
rect 53460 2370 53690 2455
rect 52060 2320 53690 2370
rect 52060 2225 52290 2320
rect 52410 2225 52640 2320
rect 52760 2225 52990 2320
rect 53110 2225 53340 2320
rect 53460 2225 53690 2320
rect 60110 2370 60340 2455
rect 60460 2370 60690 2455
rect 60810 2370 61040 2455
rect 61160 2370 61390 2455
rect 61510 2370 61740 2455
rect 60110 2320 61740 2370
rect 60110 2225 60340 2320
rect 60460 2225 60690 2320
rect 60810 2225 61040 2320
rect 61160 2225 61390 2320
rect 61510 2225 61740 2320
rect 52850 2105 52900 2225
rect 60900 2105 60950 2225
rect 52060 2020 52290 2105
rect 52410 2020 52640 2105
rect 52760 2020 52990 2105
rect 53110 2020 53340 2105
rect 53460 2020 53690 2105
rect 52060 1970 53690 2020
rect 52060 1875 52290 1970
rect 52410 1875 52640 1970
rect 52760 1875 52990 1970
rect 53110 1875 53340 1970
rect 53460 1875 53690 1970
rect 60110 2020 60340 2105
rect 60460 2020 60690 2105
rect 60810 2020 61040 2105
rect 61160 2020 61390 2105
rect 61510 2020 61740 2105
rect 60110 1970 61740 2020
rect 60110 1875 60340 1970
rect 60460 1875 60690 1970
rect 60810 1875 61040 1970
rect 61160 1875 61390 1970
rect 61510 1875 61740 1970
rect 52850 1755 52900 1875
rect 60900 1755 60950 1875
rect 52060 1670 52290 1755
rect 52410 1670 52640 1755
rect 52760 1670 52990 1755
rect 53110 1670 53340 1755
rect 53460 1670 53690 1755
rect 52060 1620 53690 1670
rect 52060 1525 52290 1620
rect 52410 1525 52640 1620
rect 52760 1525 52990 1620
rect 53110 1525 53340 1620
rect 53460 1525 53690 1620
rect 54070 1715 54320 1720
rect 54070 1675 54075 1715
rect 54115 1675 54125 1715
rect 54165 1675 54175 1715
rect 54215 1675 54225 1715
rect 54265 1675 54275 1715
rect 54315 1675 54320 1715
rect 54070 1665 54320 1675
rect 54070 1625 54075 1665
rect 54115 1625 54125 1665
rect 54165 1625 54175 1665
rect 54215 1625 54225 1665
rect 54265 1625 54275 1665
rect 54315 1625 54320 1665
rect 54070 1615 54320 1625
rect 54070 1575 54075 1615
rect 54115 1575 54125 1615
rect 54165 1575 54175 1615
rect 54215 1575 54225 1615
rect 54265 1575 54275 1615
rect 54315 1575 54320 1615
rect 54070 1570 54320 1575
rect 59480 1715 59730 1720
rect 59480 1675 59485 1715
rect 59525 1675 59535 1715
rect 59575 1675 59585 1715
rect 59625 1675 59635 1715
rect 59675 1675 59685 1715
rect 59725 1675 59730 1715
rect 59480 1665 59730 1675
rect 59480 1625 59485 1665
rect 59525 1625 59535 1665
rect 59575 1625 59585 1665
rect 59625 1625 59635 1665
rect 59675 1625 59685 1665
rect 59725 1625 59730 1665
rect 59480 1615 59730 1625
rect 59480 1575 59485 1615
rect 59525 1575 59535 1615
rect 59575 1575 59585 1615
rect 59625 1575 59635 1615
rect 59675 1575 59685 1615
rect 59725 1575 59730 1615
rect 59480 1570 59730 1575
rect 60110 1670 60340 1755
rect 60460 1670 60690 1755
rect 60810 1670 61040 1755
rect 61160 1670 61390 1755
rect 61510 1670 61740 1755
rect 60110 1620 61740 1670
rect 60110 1525 60340 1620
rect 60460 1525 60690 1620
rect 60810 1525 61040 1620
rect 61160 1525 61390 1620
rect 61510 1525 61740 1620
rect 52850 1405 52900 1525
rect 60900 1405 60950 1525
rect 52060 1320 52290 1405
rect 52410 1320 52640 1405
rect 52760 1320 52990 1405
rect 53110 1320 53340 1405
rect 53460 1320 53690 1405
rect 52060 1270 53690 1320
rect 52060 1175 52290 1270
rect 52410 1175 52640 1270
rect 52760 1175 52990 1270
rect 53110 1175 53340 1270
rect 53460 1175 53690 1270
rect 60110 1320 60340 1405
rect 60460 1320 60690 1405
rect 60810 1320 61040 1405
rect 61160 1320 61390 1405
rect 61510 1320 61740 1405
rect 60110 1270 61740 1320
rect 60110 1175 60340 1270
rect 60460 1175 60690 1270
rect 60810 1175 61040 1270
rect 61160 1175 61390 1270
rect 61510 1175 61740 1270
rect 52850 1055 52900 1175
rect 60900 1055 60950 1175
rect 52060 970 52290 1055
rect 52410 970 52640 1055
rect 52760 970 52990 1055
rect 53110 970 53340 1055
rect 53460 970 53690 1055
rect 52060 920 53690 970
rect 52060 825 52290 920
rect 52410 825 52640 920
rect 52760 825 52990 920
rect 53110 825 53340 920
rect 53460 825 53690 920
rect 60110 970 60340 1055
rect 60460 970 60690 1055
rect 60810 970 61040 1055
rect 61160 970 61390 1055
rect 61510 970 61740 1055
rect 60110 920 61740 970
rect 60110 825 60340 920
rect 60460 825 60690 920
rect 60810 825 61040 920
rect 61160 825 61390 920
rect 61510 825 61740 920
rect 52850 705 52900 825
rect 60900 705 60950 825
rect 52060 620 52290 705
rect 52410 620 52640 705
rect 52760 620 52990 705
rect 53110 620 53340 705
rect 53460 620 53690 705
rect 52060 570 53690 620
rect 52060 475 52290 570
rect 52410 475 52640 570
rect 52760 475 52990 570
rect 53110 475 53340 570
rect 53460 475 53690 570
rect 60110 620 60340 705
rect 60460 620 60690 705
rect 60810 620 61040 705
rect 61160 620 61390 705
rect 61510 620 61740 705
rect 60110 570 61740 620
rect 60110 475 60340 570
rect 60460 475 60690 570
rect 60810 475 61040 570
rect 61160 475 61390 570
rect 61510 475 61740 570
rect 52850 355 52900 475
rect 60900 355 60950 475
rect 52060 270 52290 355
rect 52410 270 52640 355
rect 52760 270 52990 355
rect 53110 270 53340 355
rect 53460 270 53690 355
rect 52060 220 53690 270
rect 52060 125 52290 220
rect 52410 125 52640 220
rect 52760 125 52990 220
rect 53110 125 53340 220
rect 53460 125 53690 220
rect 60110 270 60340 355
rect 60460 270 60690 355
rect 60810 270 61040 355
rect 61160 270 61390 355
rect 61510 270 61740 355
rect 60110 220 61740 270
rect 60110 125 60340 220
rect 60460 125 60690 220
rect 60810 125 61040 220
rect 61160 125 61390 220
rect 61510 125 61740 220
rect 52850 5 52900 125
rect 60900 5 60950 125
rect 52060 -80 52290 5
rect 52410 -80 52640 5
rect 52760 -80 52990 5
rect 53110 -80 53340 5
rect 53460 -80 53690 5
rect 52060 -130 53690 -80
rect 52060 -225 52290 -130
rect 52410 -225 52640 -130
rect 52760 -225 52990 -130
rect 53110 -225 53340 -130
rect 53460 -225 53690 -130
rect 60110 -80 60340 5
rect 60460 -80 60690 5
rect 60810 -80 61040 5
rect 61160 -80 61390 5
rect 61510 -80 61740 5
rect 60110 -130 61740 -80
rect 60110 -225 60340 -130
rect 60460 -225 60690 -130
rect 60810 -225 61040 -130
rect 61160 -225 61390 -130
rect 61510 -225 61740 -130
rect 52850 -345 52900 -225
rect 60900 -345 60950 -225
rect 52060 -430 52290 -345
rect 52410 -430 52640 -345
rect 52760 -430 52990 -345
rect 53110 -430 53340 -345
rect 53460 -430 53690 -345
rect 52060 -480 53690 -430
rect 52060 -575 52290 -480
rect 52410 -575 52640 -480
rect 52760 -575 52990 -480
rect 53110 -575 53340 -480
rect 53460 -575 53690 -480
rect 60110 -430 60340 -345
rect 60460 -430 60690 -345
rect 60810 -430 61040 -345
rect 61160 -430 61390 -345
rect 61510 -430 61740 -345
rect 60110 -480 61740 -430
rect 60110 -575 60340 -480
rect 60460 -575 60690 -480
rect 60810 -575 61040 -480
rect 61160 -575 61390 -480
rect 61510 -575 61740 -480
rect 52850 -695 52900 -575
rect 60900 -695 60950 -575
rect 52060 -780 52290 -695
rect 52410 -780 52640 -695
rect 52760 -780 52990 -695
rect 53110 -780 53340 -695
rect 53460 -780 53690 -695
rect 53810 -780 54040 -695
rect 54160 -780 54390 -695
rect 54510 -780 54740 -695
rect 54860 -780 55090 -695
rect 55210 -780 55440 -695
rect 55560 -780 55790 -695
rect 55910 -780 56140 -695
rect 56260 -780 56490 -695
rect 56610 -780 56840 -695
rect 52060 -830 56840 -780
rect 52060 -925 52290 -830
rect 52410 -925 52640 -830
rect 52760 -925 52990 -830
rect 53110 -925 53340 -830
rect 53460 -925 53690 -830
rect 53810 -925 54040 -830
rect 54160 -925 54390 -830
rect 54510 -925 54740 -830
rect 54860 -925 55090 -830
rect 55210 -925 55440 -830
rect 55560 -925 55790 -830
rect 55910 -925 56140 -830
rect 56260 -925 56490 -830
rect 56610 -925 56840 -830
rect 56960 -780 57190 -695
rect 57310 -780 57540 -695
rect 57660 -780 57890 -695
rect 58010 -780 58240 -695
rect 58360 -780 58590 -695
rect 58710 -780 58940 -695
rect 59060 -780 59290 -695
rect 59410 -780 59640 -695
rect 59760 -780 59990 -695
rect 60110 -780 60340 -695
rect 60460 -780 60690 -695
rect 60810 -780 61040 -695
rect 61160 -780 61390 -695
rect 61510 -780 61740 -695
rect 56960 -830 61740 -780
rect 56960 -925 57190 -830
rect 57310 -925 57540 -830
rect 57660 -925 57890 -830
rect 58010 -925 58240 -830
rect 58360 -925 58590 -830
rect 58710 -925 58940 -830
rect 59060 -925 59290 -830
rect 59410 -925 59640 -830
rect 59760 -925 59990 -830
rect 60110 -925 60340 -830
rect 60460 -925 60690 -830
rect 60810 -925 61040 -830
rect 61160 -925 61390 -830
rect 61510 -925 61740 -830
rect 52850 -1045 52900 -925
rect 53200 -1045 53250 -925
rect 53550 -1045 53600 -925
rect 53900 -1045 53950 -925
rect 54250 -1045 54300 -925
rect 54600 -1045 54650 -925
rect 54950 -1045 55000 -925
rect 55300 -1045 55350 -925
rect 55650 -1045 55700 -925
rect 56000 -1045 56050 -925
rect 56350 -1045 56400 -925
rect 56700 -1045 56750 -925
rect 57050 -1045 57100 -925
rect 57400 -1045 57450 -925
rect 57750 -1045 57800 -925
rect 58100 -1045 58150 -925
rect 58450 -1045 58500 -925
rect 58800 -1045 58850 -925
rect 59150 -1045 59200 -925
rect 59500 -1045 59550 -925
rect 59850 -1045 59900 -925
rect 60200 -1045 60250 -925
rect 60550 -1045 60600 -925
rect 60900 -1045 60950 -925
rect 52060 -1130 52290 -1045
rect 52410 -1130 52640 -1045
rect 52760 -1130 52990 -1045
rect 52060 -1180 52990 -1130
rect 52060 -1275 52290 -1180
rect 52410 -1275 52640 -1180
rect 52760 -1275 52990 -1180
rect 53110 -1275 53340 -1045
rect 53460 -1275 53690 -1045
rect 53810 -1275 54040 -1045
rect 54160 -1275 54390 -1045
rect 54510 -1275 54740 -1045
rect 54860 -1275 55090 -1045
rect 55210 -1275 55440 -1045
rect 55560 -1275 55790 -1045
rect 55910 -1275 56140 -1045
rect 56260 -1275 56490 -1045
rect 56610 -1275 56840 -1045
rect 56960 -1275 57190 -1045
rect 57310 -1275 57540 -1045
rect 57660 -1275 57890 -1045
rect 58010 -1275 58240 -1045
rect 58360 -1275 58590 -1045
rect 58710 -1275 58940 -1045
rect 59060 -1275 59290 -1045
rect 59410 -1275 59640 -1045
rect 59760 -1275 59990 -1045
rect 60110 -1275 60340 -1045
rect 60460 -1275 60690 -1045
rect 60810 -1130 61040 -1045
rect 61160 -1130 61390 -1045
rect 61510 -1130 61740 -1045
rect 60810 -1180 61740 -1130
rect 60810 -1275 61040 -1180
rect 61160 -1275 61390 -1180
rect 61510 -1275 61740 -1180
<< via3 >>
rect 54075 1710 54115 1715
rect 54075 1680 54080 1710
rect 54080 1680 54110 1710
rect 54110 1680 54115 1710
rect 54075 1675 54115 1680
rect 54125 1710 54165 1715
rect 54125 1680 54130 1710
rect 54130 1680 54160 1710
rect 54160 1680 54165 1710
rect 54125 1675 54165 1680
rect 54175 1710 54215 1715
rect 54175 1680 54180 1710
rect 54180 1680 54210 1710
rect 54210 1680 54215 1710
rect 54175 1675 54215 1680
rect 54225 1710 54265 1715
rect 54225 1680 54230 1710
rect 54230 1680 54260 1710
rect 54260 1680 54265 1710
rect 54225 1675 54265 1680
rect 54275 1710 54315 1715
rect 54275 1680 54280 1710
rect 54280 1680 54310 1710
rect 54310 1680 54315 1710
rect 54275 1675 54315 1680
rect 54075 1660 54115 1665
rect 54075 1630 54080 1660
rect 54080 1630 54110 1660
rect 54110 1630 54115 1660
rect 54075 1625 54115 1630
rect 54125 1660 54165 1665
rect 54125 1630 54130 1660
rect 54130 1630 54160 1660
rect 54160 1630 54165 1660
rect 54125 1625 54165 1630
rect 54175 1660 54215 1665
rect 54175 1630 54180 1660
rect 54180 1630 54210 1660
rect 54210 1630 54215 1660
rect 54175 1625 54215 1630
rect 54225 1660 54265 1665
rect 54225 1630 54230 1660
rect 54230 1630 54260 1660
rect 54260 1630 54265 1660
rect 54225 1625 54265 1630
rect 54275 1660 54315 1665
rect 54275 1630 54280 1660
rect 54280 1630 54310 1660
rect 54310 1630 54315 1660
rect 54275 1625 54315 1630
rect 54075 1610 54115 1615
rect 54075 1580 54080 1610
rect 54080 1580 54110 1610
rect 54110 1580 54115 1610
rect 54075 1575 54115 1580
rect 54125 1610 54165 1615
rect 54125 1580 54130 1610
rect 54130 1580 54160 1610
rect 54160 1580 54165 1610
rect 54125 1575 54165 1580
rect 54175 1610 54215 1615
rect 54175 1580 54180 1610
rect 54180 1580 54210 1610
rect 54210 1580 54215 1610
rect 54175 1575 54215 1580
rect 54225 1610 54265 1615
rect 54225 1580 54230 1610
rect 54230 1580 54260 1610
rect 54260 1580 54265 1610
rect 54225 1575 54265 1580
rect 54275 1610 54315 1615
rect 54275 1580 54280 1610
rect 54280 1580 54310 1610
rect 54310 1580 54315 1610
rect 54275 1575 54315 1580
rect 59485 1710 59525 1715
rect 59485 1680 59490 1710
rect 59490 1680 59520 1710
rect 59520 1680 59525 1710
rect 59485 1675 59525 1680
rect 59535 1710 59575 1715
rect 59535 1680 59540 1710
rect 59540 1680 59570 1710
rect 59570 1680 59575 1710
rect 59535 1675 59575 1680
rect 59585 1710 59625 1715
rect 59585 1680 59590 1710
rect 59590 1680 59620 1710
rect 59620 1680 59625 1710
rect 59585 1675 59625 1680
rect 59635 1710 59675 1715
rect 59635 1680 59640 1710
rect 59640 1680 59670 1710
rect 59670 1680 59675 1710
rect 59635 1675 59675 1680
rect 59685 1710 59725 1715
rect 59685 1680 59690 1710
rect 59690 1680 59720 1710
rect 59720 1680 59725 1710
rect 59685 1675 59725 1680
rect 59485 1660 59525 1665
rect 59485 1630 59490 1660
rect 59490 1630 59520 1660
rect 59520 1630 59525 1660
rect 59485 1625 59525 1630
rect 59535 1660 59575 1665
rect 59535 1630 59540 1660
rect 59540 1630 59570 1660
rect 59570 1630 59575 1660
rect 59535 1625 59575 1630
rect 59585 1660 59625 1665
rect 59585 1630 59590 1660
rect 59590 1630 59620 1660
rect 59620 1630 59625 1660
rect 59585 1625 59625 1630
rect 59635 1660 59675 1665
rect 59635 1630 59640 1660
rect 59640 1630 59670 1660
rect 59670 1630 59675 1660
rect 59635 1625 59675 1630
rect 59685 1660 59725 1665
rect 59685 1630 59690 1660
rect 59690 1630 59720 1660
rect 59720 1630 59725 1660
rect 59685 1625 59725 1630
rect 59485 1610 59525 1615
rect 59485 1580 59490 1610
rect 59490 1580 59520 1610
rect 59520 1580 59525 1610
rect 59485 1575 59525 1580
rect 59535 1610 59575 1615
rect 59535 1580 59540 1610
rect 59540 1580 59570 1610
rect 59570 1580 59575 1610
rect 59535 1575 59575 1580
rect 59585 1610 59625 1615
rect 59585 1580 59590 1610
rect 59590 1580 59620 1610
rect 59620 1580 59625 1610
rect 59585 1575 59625 1580
rect 59635 1610 59675 1615
rect 59635 1580 59640 1610
rect 59640 1580 59670 1610
rect 59670 1580 59675 1610
rect 59635 1575 59675 1580
rect 59685 1610 59725 1615
rect 59685 1580 59690 1610
rect 59690 1580 59720 1610
rect 59720 1580 59725 1610
rect 59685 1575 59725 1580
<< mimcap >>
rect 52075 5515 52275 5590
rect 52075 5475 52155 5515
rect 52195 5475 52275 5515
rect 52075 5390 52275 5475
rect 52425 5515 52625 5590
rect 52425 5475 52505 5515
rect 52545 5475 52625 5515
rect 52425 5390 52625 5475
rect 52775 5515 52975 5590
rect 52775 5475 52855 5515
rect 52895 5475 52975 5515
rect 52775 5390 52975 5475
rect 53125 5515 53325 5590
rect 53125 5475 53205 5515
rect 53245 5475 53325 5515
rect 53125 5390 53325 5475
rect 53475 5515 53675 5590
rect 53475 5475 53555 5515
rect 53595 5475 53675 5515
rect 53475 5390 53675 5475
rect 53825 5515 54025 5590
rect 53825 5475 53905 5515
rect 53945 5475 54025 5515
rect 53825 5390 54025 5475
rect 54175 5515 54375 5590
rect 54175 5475 54255 5515
rect 54295 5475 54375 5515
rect 54175 5390 54375 5475
rect 54525 5515 54725 5590
rect 54525 5475 54605 5515
rect 54645 5475 54725 5515
rect 54525 5390 54725 5475
rect 54875 5515 55075 5590
rect 54875 5475 54955 5515
rect 54995 5475 55075 5515
rect 54875 5390 55075 5475
rect 55225 5515 55425 5590
rect 55225 5475 55305 5515
rect 55345 5475 55425 5515
rect 55225 5390 55425 5475
rect 55575 5515 55775 5590
rect 55575 5475 55655 5515
rect 55695 5475 55775 5515
rect 55575 5390 55775 5475
rect 55925 5515 56125 5590
rect 55925 5475 56005 5515
rect 56045 5475 56125 5515
rect 55925 5390 56125 5475
rect 56275 5515 56475 5590
rect 56275 5475 56355 5515
rect 56395 5475 56475 5515
rect 56275 5390 56475 5475
rect 56625 5515 56825 5590
rect 56625 5475 56705 5515
rect 56745 5475 56825 5515
rect 56625 5390 56825 5475
rect 56975 5515 57175 5590
rect 56975 5475 57055 5515
rect 57095 5475 57175 5515
rect 56975 5390 57175 5475
rect 57325 5515 57525 5590
rect 57325 5475 57405 5515
rect 57445 5475 57525 5515
rect 57325 5390 57525 5475
rect 57675 5515 57875 5590
rect 57675 5475 57755 5515
rect 57795 5475 57875 5515
rect 57675 5390 57875 5475
rect 58025 5515 58225 5590
rect 58025 5475 58105 5515
rect 58145 5475 58225 5515
rect 58025 5390 58225 5475
rect 58375 5515 58575 5590
rect 58375 5475 58455 5515
rect 58495 5475 58575 5515
rect 58375 5390 58575 5475
rect 58725 5515 58925 5590
rect 58725 5475 58805 5515
rect 58845 5475 58925 5515
rect 58725 5390 58925 5475
rect 59075 5515 59275 5590
rect 59075 5475 59155 5515
rect 59195 5475 59275 5515
rect 59075 5390 59275 5475
rect 59425 5515 59625 5590
rect 59425 5475 59505 5515
rect 59545 5475 59625 5515
rect 59425 5390 59625 5475
rect 59775 5515 59975 5590
rect 59775 5475 59855 5515
rect 59895 5475 59975 5515
rect 59775 5390 59975 5475
rect 60125 5515 60325 5590
rect 60125 5475 60205 5515
rect 60245 5475 60325 5515
rect 60125 5390 60325 5475
rect 60475 5515 60675 5590
rect 60475 5475 60555 5515
rect 60595 5475 60675 5515
rect 60475 5390 60675 5475
rect 60825 5515 61025 5590
rect 60825 5475 60905 5515
rect 60945 5475 61025 5515
rect 60825 5390 61025 5475
rect 61175 5515 61375 5590
rect 61175 5475 61255 5515
rect 61295 5475 61375 5515
rect 61175 5390 61375 5475
rect 61525 5515 61725 5590
rect 61525 5475 61605 5515
rect 61645 5475 61725 5515
rect 61525 5390 61725 5475
rect 52075 5165 52275 5240
rect 52075 5125 52155 5165
rect 52195 5125 52275 5165
rect 52075 5040 52275 5125
rect 52425 5165 52625 5240
rect 52425 5125 52505 5165
rect 52545 5125 52625 5165
rect 52425 5040 52625 5125
rect 52775 5165 52975 5240
rect 52775 5125 52855 5165
rect 52895 5125 52975 5165
rect 52775 5040 52975 5125
rect 53125 5165 53325 5240
rect 53125 5125 53205 5165
rect 53245 5125 53325 5165
rect 53125 5040 53325 5125
rect 53475 5165 53675 5240
rect 53475 5125 53555 5165
rect 53595 5125 53675 5165
rect 53475 5040 53675 5125
rect 53825 5165 54025 5240
rect 53825 5125 53905 5165
rect 53945 5125 54025 5165
rect 53825 5040 54025 5125
rect 54175 5165 54375 5240
rect 54175 5125 54255 5165
rect 54295 5125 54375 5165
rect 54175 5040 54375 5125
rect 54525 5165 54725 5240
rect 54525 5125 54605 5165
rect 54645 5125 54725 5165
rect 54525 5040 54725 5125
rect 54875 5165 55075 5240
rect 54875 5125 54955 5165
rect 54995 5125 55075 5165
rect 54875 5040 55075 5125
rect 55225 5155 55425 5240
rect 55225 5115 55305 5155
rect 55345 5115 55425 5155
rect 55225 5040 55425 5115
rect 55575 5155 55775 5240
rect 55575 5115 55655 5155
rect 55695 5115 55775 5155
rect 55575 5040 55775 5115
rect 58025 5155 58225 5240
rect 58025 5115 58105 5155
rect 58145 5115 58225 5155
rect 58025 5040 58225 5115
rect 58375 5155 58575 5240
rect 58375 5115 58455 5155
rect 58495 5115 58575 5155
rect 58375 5040 58575 5115
rect 58725 5165 58925 5240
rect 58725 5125 58805 5165
rect 58845 5125 58925 5165
rect 58725 5040 58925 5125
rect 59075 5165 59275 5240
rect 59075 5125 59155 5165
rect 59195 5125 59275 5165
rect 59075 5040 59275 5125
rect 59425 5165 59625 5240
rect 59425 5125 59505 5165
rect 59545 5125 59625 5165
rect 59425 5040 59625 5125
rect 59775 5165 59975 5240
rect 59775 5125 59855 5165
rect 59895 5125 59975 5165
rect 59775 5040 59975 5125
rect 60125 5165 60325 5240
rect 60125 5125 60205 5165
rect 60245 5125 60325 5165
rect 60125 5040 60325 5125
rect 60475 5165 60675 5240
rect 60475 5125 60555 5165
rect 60595 5125 60675 5165
rect 60475 5040 60675 5125
rect 60825 5165 61025 5240
rect 60825 5125 60905 5165
rect 60945 5125 61025 5165
rect 60825 5040 61025 5125
rect 61175 5165 61375 5240
rect 61175 5125 61255 5165
rect 61295 5125 61375 5165
rect 61175 5040 61375 5125
rect 61525 5165 61725 5240
rect 61525 5125 61605 5165
rect 61645 5125 61725 5165
rect 61525 5040 61725 5125
rect 52075 4815 52275 4890
rect 52075 4775 52155 4815
rect 52195 4775 52275 4815
rect 52075 4690 52275 4775
rect 52425 4815 52625 4890
rect 52425 4775 52505 4815
rect 52545 4775 52625 4815
rect 52425 4690 52625 4775
rect 52775 4815 52975 4890
rect 52775 4775 52855 4815
rect 52895 4775 52975 4815
rect 52775 4690 52975 4775
rect 53125 4815 53325 4890
rect 53125 4775 53205 4815
rect 53245 4775 53325 4815
rect 53125 4690 53325 4775
rect 53475 4815 53675 4890
rect 53475 4775 53555 4815
rect 53595 4775 53675 4815
rect 53475 4690 53675 4775
rect 53825 4815 54025 4890
rect 53825 4775 53905 4815
rect 53945 4775 54025 4815
rect 53825 4690 54025 4775
rect 54175 4815 54375 4890
rect 54175 4775 54255 4815
rect 54295 4775 54375 4815
rect 54175 4690 54375 4775
rect 54525 4815 54725 4890
rect 54525 4775 54605 4815
rect 54645 4775 54725 4815
rect 54525 4690 54725 4775
rect 54875 4815 55075 4890
rect 54875 4775 54955 4815
rect 54995 4775 55075 4815
rect 54875 4690 55075 4775
rect 55225 4805 55425 4890
rect 55225 4765 55305 4805
rect 55345 4765 55425 4805
rect 55225 4690 55425 4765
rect 58375 4805 58575 4890
rect 58375 4765 58455 4805
rect 58495 4765 58575 4805
rect 58375 4690 58575 4765
rect 58725 4815 58925 4890
rect 58725 4775 58805 4815
rect 58845 4775 58925 4815
rect 58725 4690 58925 4775
rect 59075 4815 59275 4890
rect 59075 4775 59155 4815
rect 59195 4775 59275 4815
rect 59075 4690 59275 4775
rect 59425 4815 59625 4890
rect 59425 4775 59505 4815
rect 59545 4775 59625 4815
rect 59425 4690 59625 4775
rect 59775 4815 59975 4890
rect 59775 4775 59855 4815
rect 59895 4775 59975 4815
rect 59775 4690 59975 4775
rect 60125 4815 60325 4890
rect 60125 4775 60205 4815
rect 60245 4775 60325 4815
rect 60125 4690 60325 4775
rect 60475 4815 60675 4890
rect 60475 4775 60555 4815
rect 60595 4775 60675 4815
rect 60475 4690 60675 4775
rect 60825 4815 61025 4890
rect 60825 4775 60905 4815
rect 60945 4775 61025 4815
rect 60825 4690 61025 4775
rect 61175 4815 61375 4890
rect 61175 4775 61255 4815
rect 61295 4775 61375 4815
rect 61175 4690 61375 4775
rect 61525 4815 61725 4890
rect 61525 4775 61605 4815
rect 61645 4775 61725 4815
rect 61525 4690 61725 4775
rect 52075 4465 52275 4540
rect 52075 4425 52155 4465
rect 52195 4425 52275 4465
rect 52075 4340 52275 4425
rect 52425 4465 52625 4540
rect 52425 4425 52505 4465
rect 52545 4425 52625 4465
rect 52425 4340 52625 4425
rect 52775 4465 52975 4540
rect 52775 4425 52855 4465
rect 52895 4425 52975 4465
rect 52775 4340 52975 4425
rect 53125 4465 53325 4540
rect 53125 4425 53205 4465
rect 53245 4425 53325 4465
rect 53125 4340 53325 4425
rect 53475 4465 53675 4540
rect 53475 4425 53555 4465
rect 53595 4425 53675 4465
rect 53475 4340 53675 4425
rect 60125 4465 60325 4540
rect 60125 4425 60205 4465
rect 60245 4425 60325 4465
rect 60125 4340 60325 4425
rect 60475 4465 60675 4540
rect 60475 4425 60555 4465
rect 60595 4425 60675 4465
rect 60475 4340 60675 4425
rect 60825 4465 61025 4540
rect 60825 4425 60905 4465
rect 60945 4425 61025 4465
rect 60825 4340 61025 4425
rect 61175 4465 61375 4540
rect 61175 4425 61255 4465
rect 61295 4425 61375 4465
rect 61175 4340 61375 4425
rect 61525 4465 61725 4540
rect 61525 4425 61605 4465
rect 61645 4425 61725 4465
rect 61525 4340 61725 4425
rect 52075 4115 52275 4190
rect 52075 4075 52155 4115
rect 52195 4075 52275 4115
rect 52075 3990 52275 4075
rect 52425 4115 52625 4190
rect 52425 4075 52505 4115
rect 52545 4075 52625 4115
rect 52425 3990 52625 4075
rect 52775 4115 52975 4190
rect 52775 4075 52855 4115
rect 52895 4075 52975 4115
rect 52775 3990 52975 4075
rect 53125 4115 53325 4190
rect 53125 4075 53205 4115
rect 53245 4075 53325 4115
rect 53125 3990 53325 4075
rect 53475 4115 53675 4190
rect 53475 4075 53555 4115
rect 53595 4075 53675 4115
rect 53475 3990 53675 4075
rect 60125 4115 60325 4190
rect 60125 4075 60205 4115
rect 60245 4075 60325 4115
rect 60125 3990 60325 4075
rect 60475 4115 60675 4190
rect 60475 4075 60555 4115
rect 60595 4075 60675 4115
rect 60475 3990 60675 4075
rect 60825 4115 61025 4190
rect 60825 4075 60905 4115
rect 60945 4075 61025 4115
rect 60825 3990 61025 4075
rect 61175 4115 61375 4190
rect 61175 4075 61255 4115
rect 61295 4075 61375 4115
rect 61175 3990 61375 4075
rect 61525 4115 61725 4190
rect 61525 4075 61605 4115
rect 61645 4075 61725 4115
rect 61525 3990 61725 4075
rect 52075 3765 52275 3840
rect 52075 3725 52155 3765
rect 52195 3725 52275 3765
rect 52075 3640 52275 3725
rect 52425 3765 52625 3840
rect 52425 3725 52505 3765
rect 52545 3725 52625 3765
rect 52425 3640 52625 3725
rect 52775 3765 52975 3840
rect 52775 3725 52855 3765
rect 52895 3725 52975 3765
rect 52775 3640 52975 3725
rect 53125 3765 53325 3840
rect 53125 3725 53205 3765
rect 53245 3725 53325 3765
rect 53125 3640 53325 3725
rect 53475 3765 53675 3840
rect 53475 3725 53555 3765
rect 53595 3725 53675 3765
rect 53475 3640 53675 3725
rect 60125 3765 60325 3840
rect 60125 3725 60205 3765
rect 60245 3725 60325 3765
rect 60125 3640 60325 3725
rect 60475 3765 60675 3840
rect 60475 3725 60555 3765
rect 60595 3725 60675 3765
rect 60475 3640 60675 3725
rect 60825 3765 61025 3840
rect 60825 3725 60905 3765
rect 60945 3725 61025 3765
rect 60825 3640 61025 3725
rect 61175 3765 61375 3840
rect 61175 3725 61255 3765
rect 61295 3725 61375 3765
rect 61175 3640 61375 3725
rect 61525 3765 61725 3840
rect 61525 3725 61605 3765
rect 61645 3725 61725 3765
rect 61525 3640 61725 3725
rect 52075 3415 52275 3490
rect 52075 3375 52155 3415
rect 52195 3375 52275 3415
rect 52075 3290 52275 3375
rect 52425 3415 52625 3490
rect 52425 3375 52505 3415
rect 52545 3375 52625 3415
rect 52425 3290 52625 3375
rect 52775 3415 52975 3490
rect 52775 3375 52855 3415
rect 52895 3375 52975 3415
rect 52775 3290 52975 3375
rect 53125 3415 53325 3490
rect 53125 3375 53205 3415
rect 53245 3375 53325 3415
rect 53125 3290 53325 3375
rect 53475 3415 53675 3490
rect 53475 3375 53555 3415
rect 53595 3375 53675 3415
rect 53475 3290 53675 3375
rect 60125 3415 60325 3490
rect 60125 3375 60205 3415
rect 60245 3375 60325 3415
rect 60125 3290 60325 3375
rect 60475 3415 60675 3490
rect 60475 3375 60555 3415
rect 60595 3375 60675 3415
rect 60475 3290 60675 3375
rect 60825 3415 61025 3490
rect 60825 3375 60905 3415
rect 60945 3375 61025 3415
rect 60825 3290 61025 3375
rect 61175 3415 61375 3490
rect 61175 3375 61255 3415
rect 61295 3375 61375 3415
rect 61175 3290 61375 3375
rect 61525 3415 61725 3490
rect 61525 3375 61605 3415
rect 61645 3375 61725 3415
rect 61525 3290 61725 3375
rect 52075 3065 52275 3140
rect 52075 3025 52155 3065
rect 52195 3025 52275 3065
rect 52075 2940 52275 3025
rect 52425 3065 52625 3140
rect 52425 3025 52505 3065
rect 52545 3025 52625 3065
rect 52425 2940 52625 3025
rect 52775 3065 52975 3140
rect 52775 3025 52855 3065
rect 52895 3025 52975 3065
rect 52775 2940 52975 3025
rect 53125 3065 53325 3140
rect 53125 3025 53205 3065
rect 53245 3025 53325 3065
rect 53125 2940 53325 3025
rect 53475 3065 53675 3140
rect 53475 3025 53555 3065
rect 53595 3025 53675 3065
rect 53475 2940 53675 3025
rect 60125 3065 60325 3140
rect 60125 3025 60205 3065
rect 60245 3025 60325 3065
rect 60125 2940 60325 3025
rect 60475 3065 60675 3140
rect 60475 3025 60555 3065
rect 60595 3025 60675 3065
rect 60475 2940 60675 3025
rect 60825 3065 61025 3140
rect 60825 3025 60905 3065
rect 60945 3025 61025 3065
rect 60825 2940 61025 3025
rect 61175 3065 61375 3140
rect 61175 3025 61255 3065
rect 61295 3025 61375 3065
rect 61175 2940 61375 3025
rect 61525 3065 61725 3140
rect 61525 3025 61605 3065
rect 61645 3025 61725 3065
rect 61525 2940 61725 3025
rect 52075 2715 52275 2790
rect 52075 2675 52155 2715
rect 52195 2675 52275 2715
rect 52075 2590 52275 2675
rect 52425 2715 52625 2790
rect 52425 2675 52505 2715
rect 52545 2675 52625 2715
rect 52425 2590 52625 2675
rect 52775 2715 52975 2790
rect 52775 2675 52855 2715
rect 52895 2675 52975 2715
rect 52775 2590 52975 2675
rect 53125 2715 53325 2790
rect 53125 2675 53205 2715
rect 53245 2675 53325 2715
rect 53125 2590 53325 2675
rect 53475 2715 53675 2790
rect 53475 2675 53555 2715
rect 53595 2675 53675 2715
rect 53475 2590 53675 2675
rect 60125 2715 60325 2790
rect 60125 2675 60205 2715
rect 60245 2675 60325 2715
rect 60125 2590 60325 2675
rect 60475 2715 60675 2790
rect 60475 2675 60555 2715
rect 60595 2675 60675 2715
rect 60475 2590 60675 2675
rect 60825 2715 61025 2790
rect 60825 2675 60905 2715
rect 60945 2675 61025 2715
rect 60825 2590 61025 2675
rect 61175 2715 61375 2790
rect 61175 2675 61255 2715
rect 61295 2675 61375 2715
rect 61175 2590 61375 2675
rect 61525 2715 61725 2790
rect 61525 2675 61605 2715
rect 61645 2675 61725 2715
rect 61525 2590 61725 2675
rect 52075 2365 52275 2440
rect 52075 2325 52155 2365
rect 52195 2325 52275 2365
rect 52075 2240 52275 2325
rect 52425 2365 52625 2440
rect 52425 2325 52505 2365
rect 52545 2325 52625 2365
rect 52425 2240 52625 2325
rect 52775 2365 52975 2440
rect 52775 2325 52855 2365
rect 52895 2325 52975 2365
rect 52775 2240 52975 2325
rect 53125 2365 53325 2440
rect 53125 2325 53205 2365
rect 53245 2325 53325 2365
rect 53125 2240 53325 2325
rect 53475 2365 53675 2440
rect 53475 2325 53555 2365
rect 53595 2325 53675 2365
rect 53475 2240 53675 2325
rect 60125 2365 60325 2440
rect 60125 2325 60205 2365
rect 60245 2325 60325 2365
rect 60125 2240 60325 2325
rect 60475 2365 60675 2440
rect 60475 2325 60555 2365
rect 60595 2325 60675 2365
rect 60475 2240 60675 2325
rect 60825 2365 61025 2440
rect 60825 2325 60905 2365
rect 60945 2325 61025 2365
rect 60825 2240 61025 2325
rect 61175 2365 61375 2440
rect 61175 2325 61255 2365
rect 61295 2325 61375 2365
rect 61175 2240 61375 2325
rect 61525 2365 61725 2440
rect 61525 2325 61605 2365
rect 61645 2325 61725 2365
rect 61525 2240 61725 2325
rect 52075 2015 52275 2090
rect 52075 1975 52155 2015
rect 52195 1975 52275 2015
rect 52075 1890 52275 1975
rect 52425 2015 52625 2090
rect 52425 1975 52505 2015
rect 52545 1975 52625 2015
rect 52425 1890 52625 1975
rect 52775 2015 52975 2090
rect 52775 1975 52855 2015
rect 52895 1975 52975 2015
rect 52775 1890 52975 1975
rect 53125 2015 53325 2090
rect 53125 1975 53205 2015
rect 53245 1975 53325 2015
rect 53125 1890 53325 1975
rect 53475 2015 53675 2090
rect 53475 1975 53555 2015
rect 53595 1975 53675 2015
rect 53475 1890 53675 1975
rect 60125 2015 60325 2090
rect 60125 1975 60205 2015
rect 60245 1975 60325 2015
rect 60125 1890 60325 1975
rect 60475 2015 60675 2090
rect 60475 1975 60555 2015
rect 60595 1975 60675 2015
rect 60475 1890 60675 1975
rect 60825 2015 61025 2090
rect 60825 1975 60905 2015
rect 60945 1975 61025 2015
rect 60825 1890 61025 1975
rect 61175 2015 61375 2090
rect 61175 1975 61255 2015
rect 61295 1975 61375 2015
rect 61175 1890 61375 1975
rect 61525 2015 61725 2090
rect 61525 1975 61605 2015
rect 61645 1975 61725 2015
rect 61525 1890 61725 1975
rect 52075 1665 52275 1740
rect 52075 1625 52155 1665
rect 52195 1625 52275 1665
rect 52075 1540 52275 1625
rect 52425 1665 52625 1740
rect 52425 1625 52505 1665
rect 52545 1625 52625 1665
rect 52425 1540 52625 1625
rect 52775 1665 52975 1740
rect 52775 1625 52855 1665
rect 52895 1625 52975 1665
rect 52775 1540 52975 1625
rect 53125 1665 53325 1740
rect 53125 1625 53205 1665
rect 53245 1625 53325 1665
rect 53125 1540 53325 1625
rect 53475 1665 53675 1740
rect 53475 1625 53555 1665
rect 53595 1625 53675 1665
rect 53475 1540 53675 1625
rect 60125 1665 60325 1740
rect 60125 1625 60205 1665
rect 60245 1625 60325 1665
rect 60125 1540 60325 1625
rect 60475 1665 60675 1740
rect 60475 1625 60555 1665
rect 60595 1625 60675 1665
rect 60475 1540 60675 1625
rect 60825 1665 61025 1740
rect 60825 1625 60905 1665
rect 60945 1625 61025 1665
rect 60825 1540 61025 1625
rect 61175 1665 61375 1740
rect 61175 1625 61255 1665
rect 61295 1625 61375 1665
rect 61175 1540 61375 1625
rect 61525 1665 61725 1740
rect 61525 1625 61605 1665
rect 61645 1625 61725 1665
rect 61525 1540 61725 1625
rect 52075 1315 52275 1390
rect 52075 1275 52155 1315
rect 52195 1275 52275 1315
rect 52075 1190 52275 1275
rect 52425 1315 52625 1390
rect 52425 1275 52505 1315
rect 52545 1275 52625 1315
rect 52425 1190 52625 1275
rect 52775 1315 52975 1390
rect 52775 1275 52855 1315
rect 52895 1275 52975 1315
rect 52775 1190 52975 1275
rect 53125 1315 53325 1390
rect 53125 1275 53205 1315
rect 53245 1275 53325 1315
rect 53125 1190 53325 1275
rect 53475 1315 53675 1390
rect 53475 1275 53555 1315
rect 53595 1275 53675 1315
rect 53475 1190 53675 1275
rect 60125 1315 60325 1390
rect 60125 1275 60205 1315
rect 60245 1275 60325 1315
rect 60125 1190 60325 1275
rect 60475 1315 60675 1390
rect 60475 1275 60555 1315
rect 60595 1275 60675 1315
rect 60475 1190 60675 1275
rect 60825 1315 61025 1390
rect 60825 1275 60905 1315
rect 60945 1275 61025 1315
rect 60825 1190 61025 1275
rect 61175 1315 61375 1390
rect 61175 1275 61255 1315
rect 61295 1275 61375 1315
rect 61175 1190 61375 1275
rect 61525 1315 61725 1390
rect 61525 1275 61605 1315
rect 61645 1275 61725 1315
rect 61525 1190 61725 1275
rect 52075 965 52275 1040
rect 52075 925 52155 965
rect 52195 925 52275 965
rect 52075 840 52275 925
rect 52425 965 52625 1040
rect 52425 925 52505 965
rect 52545 925 52625 965
rect 52425 840 52625 925
rect 52775 965 52975 1040
rect 52775 925 52855 965
rect 52895 925 52975 965
rect 52775 840 52975 925
rect 53125 965 53325 1040
rect 53125 925 53205 965
rect 53245 925 53325 965
rect 53125 840 53325 925
rect 53475 965 53675 1040
rect 53475 925 53555 965
rect 53595 925 53675 965
rect 53475 840 53675 925
rect 60125 965 60325 1040
rect 60125 925 60205 965
rect 60245 925 60325 965
rect 60125 840 60325 925
rect 60475 965 60675 1040
rect 60475 925 60555 965
rect 60595 925 60675 965
rect 60475 840 60675 925
rect 60825 965 61025 1040
rect 60825 925 60905 965
rect 60945 925 61025 965
rect 60825 840 61025 925
rect 61175 965 61375 1040
rect 61175 925 61255 965
rect 61295 925 61375 965
rect 61175 840 61375 925
rect 61525 965 61725 1040
rect 61525 925 61605 965
rect 61645 925 61725 965
rect 61525 840 61725 925
rect 52075 615 52275 690
rect 52075 575 52155 615
rect 52195 575 52275 615
rect 52075 490 52275 575
rect 52425 615 52625 690
rect 52425 575 52505 615
rect 52545 575 52625 615
rect 52425 490 52625 575
rect 52775 615 52975 690
rect 52775 575 52855 615
rect 52895 575 52975 615
rect 52775 490 52975 575
rect 53125 615 53325 690
rect 53125 575 53205 615
rect 53245 575 53325 615
rect 53125 490 53325 575
rect 53475 615 53675 690
rect 53475 575 53555 615
rect 53595 575 53675 615
rect 53475 490 53675 575
rect 60125 615 60325 690
rect 60125 575 60205 615
rect 60245 575 60325 615
rect 60125 490 60325 575
rect 60475 615 60675 690
rect 60475 575 60555 615
rect 60595 575 60675 615
rect 60475 490 60675 575
rect 60825 615 61025 690
rect 60825 575 60905 615
rect 60945 575 61025 615
rect 60825 490 61025 575
rect 61175 615 61375 690
rect 61175 575 61255 615
rect 61295 575 61375 615
rect 61175 490 61375 575
rect 61525 615 61725 690
rect 61525 575 61605 615
rect 61645 575 61725 615
rect 61525 490 61725 575
rect 52075 265 52275 340
rect 52075 225 52155 265
rect 52195 225 52275 265
rect 52075 140 52275 225
rect 52425 265 52625 340
rect 52425 225 52505 265
rect 52545 225 52625 265
rect 52425 140 52625 225
rect 52775 265 52975 340
rect 52775 225 52855 265
rect 52895 225 52975 265
rect 52775 140 52975 225
rect 53125 265 53325 340
rect 53125 225 53205 265
rect 53245 225 53325 265
rect 53125 140 53325 225
rect 53475 265 53675 340
rect 53475 225 53555 265
rect 53595 225 53675 265
rect 53475 140 53675 225
rect 60125 265 60325 340
rect 60125 225 60205 265
rect 60245 225 60325 265
rect 60125 140 60325 225
rect 60475 265 60675 340
rect 60475 225 60555 265
rect 60595 225 60675 265
rect 60475 140 60675 225
rect 60825 265 61025 340
rect 60825 225 60905 265
rect 60945 225 61025 265
rect 60825 140 61025 225
rect 61175 265 61375 340
rect 61175 225 61255 265
rect 61295 225 61375 265
rect 61175 140 61375 225
rect 61525 265 61725 340
rect 61525 225 61605 265
rect 61645 225 61725 265
rect 61525 140 61725 225
rect 52075 -85 52275 -10
rect 52075 -125 52155 -85
rect 52195 -125 52275 -85
rect 52075 -210 52275 -125
rect 52425 -85 52625 -10
rect 52425 -125 52505 -85
rect 52545 -125 52625 -85
rect 52425 -210 52625 -125
rect 52775 -85 52975 -10
rect 52775 -125 52855 -85
rect 52895 -125 52975 -85
rect 52775 -210 52975 -125
rect 53125 -85 53325 -10
rect 53125 -125 53205 -85
rect 53245 -125 53325 -85
rect 53125 -210 53325 -125
rect 53475 -85 53675 -10
rect 53475 -125 53555 -85
rect 53595 -125 53675 -85
rect 53475 -210 53675 -125
rect 60125 -85 60325 -10
rect 60125 -125 60205 -85
rect 60245 -125 60325 -85
rect 60125 -210 60325 -125
rect 60475 -85 60675 -10
rect 60475 -125 60555 -85
rect 60595 -125 60675 -85
rect 60475 -210 60675 -125
rect 60825 -85 61025 -10
rect 60825 -125 60905 -85
rect 60945 -125 61025 -85
rect 60825 -210 61025 -125
rect 61175 -85 61375 -10
rect 61175 -125 61255 -85
rect 61295 -125 61375 -85
rect 61175 -210 61375 -125
rect 61525 -85 61725 -10
rect 61525 -125 61605 -85
rect 61645 -125 61725 -85
rect 61525 -210 61725 -125
rect 52075 -435 52275 -360
rect 52075 -475 52155 -435
rect 52195 -475 52275 -435
rect 52075 -560 52275 -475
rect 52425 -435 52625 -360
rect 52425 -475 52505 -435
rect 52545 -475 52625 -435
rect 52425 -560 52625 -475
rect 52775 -435 52975 -360
rect 52775 -475 52855 -435
rect 52895 -475 52975 -435
rect 52775 -560 52975 -475
rect 53125 -435 53325 -360
rect 53125 -475 53205 -435
rect 53245 -475 53325 -435
rect 53125 -560 53325 -475
rect 53475 -435 53675 -360
rect 53475 -475 53555 -435
rect 53595 -475 53675 -435
rect 53475 -560 53675 -475
rect 60125 -435 60325 -360
rect 60125 -475 60205 -435
rect 60245 -475 60325 -435
rect 60125 -560 60325 -475
rect 60475 -435 60675 -360
rect 60475 -475 60555 -435
rect 60595 -475 60675 -435
rect 60475 -560 60675 -475
rect 60825 -435 61025 -360
rect 60825 -475 60905 -435
rect 60945 -475 61025 -435
rect 60825 -560 61025 -475
rect 61175 -435 61375 -360
rect 61175 -475 61255 -435
rect 61295 -475 61375 -435
rect 61175 -560 61375 -475
rect 61525 -435 61725 -360
rect 61525 -475 61605 -435
rect 61645 -475 61725 -435
rect 61525 -560 61725 -475
rect 52075 -785 52275 -710
rect 52075 -825 52155 -785
rect 52195 -825 52275 -785
rect 52075 -910 52275 -825
rect 52425 -785 52625 -710
rect 52425 -825 52505 -785
rect 52545 -825 52625 -785
rect 52425 -910 52625 -825
rect 52775 -785 52975 -710
rect 52775 -825 52855 -785
rect 52895 -825 52975 -785
rect 52775 -910 52975 -825
rect 53125 -785 53325 -710
rect 53125 -825 53205 -785
rect 53245 -825 53325 -785
rect 53125 -910 53325 -825
rect 53475 -785 53675 -710
rect 53475 -825 53555 -785
rect 53595 -825 53675 -785
rect 53475 -910 53675 -825
rect 53825 -785 54025 -710
rect 53825 -825 53905 -785
rect 53945 -825 54025 -785
rect 53825 -910 54025 -825
rect 54175 -785 54375 -710
rect 54175 -825 54255 -785
rect 54295 -825 54375 -785
rect 54175 -910 54375 -825
rect 54525 -785 54725 -710
rect 54525 -825 54605 -785
rect 54645 -825 54725 -785
rect 54525 -910 54725 -825
rect 54875 -785 55075 -710
rect 54875 -825 54955 -785
rect 54995 -825 55075 -785
rect 54875 -910 55075 -825
rect 55225 -785 55425 -710
rect 55225 -825 55305 -785
rect 55345 -825 55425 -785
rect 55225 -910 55425 -825
rect 55575 -785 55775 -710
rect 55575 -825 55655 -785
rect 55695 -825 55775 -785
rect 55575 -910 55775 -825
rect 55925 -785 56125 -710
rect 55925 -825 56005 -785
rect 56045 -825 56125 -785
rect 55925 -910 56125 -825
rect 56275 -785 56475 -710
rect 56275 -825 56355 -785
rect 56395 -825 56475 -785
rect 56275 -910 56475 -825
rect 56625 -785 56825 -710
rect 56625 -825 56705 -785
rect 56745 -825 56825 -785
rect 56625 -910 56825 -825
rect 56975 -785 57175 -710
rect 56975 -825 57055 -785
rect 57095 -825 57175 -785
rect 56975 -910 57175 -825
rect 57325 -785 57525 -710
rect 57325 -825 57405 -785
rect 57445 -825 57525 -785
rect 57325 -910 57525 -825
rect 57675 -785 57875 -710
rect 57675 -825 57755 -785
rect 57795 -825 57875 -785
rect 57675 -910 57875 -825
rect 58025 -785 58225 -710
rect 58025 -825 58105 -785
rect 58145 -825 58225 -785
rect 58025 -910 58225 -825
rect 58375 -785 58575 -710
rect 58375 -825 58455 -785
rect 58495 -825 58575 -785
rect 58375 -910 58575 -825
rect 58725 -785 58925 -710
rect 58725 -825 58805 -785
rect 58845 -825 58925 -785
rect 58725 -910 58925 -825
rect 59075 -785 59275 -710
rect 59075 -825 59155 -785
rect 59195 -825 59275 -785
rect 59075 -910 59275 -825
rect 59425 -785 59625 -710
rect 59425 -825 59505 -785
rect 59545 -825 59625 -785
rect 59425 -910 59625 -825
rect 59775 -785 59975 -710
rect 59775 -825 59855 -785
rect 59895 -825 59975 -785
rect 59775 -910 59975 -825
rect 60125 -785 60325 -710
rect 60125 -825 60205 -785
rect 60245 -825 60325 -785
rect 60125 -910 60325 -825
rect 60475 -785 60675 -710
rect 60475 -825 60555 -785
rect 60595 -825 60675 -785
rect 60475 -910 60675 -825
rect 60825 -785 61025 -710
rect 60825 -825 60905 -785
rect 60945 -825 61025 -785
rect 60825 -910 61025 -825
rect 61175 -785 61375 -710
rect 61175 -825 61255 -785
rect 61295 -825 61375 -785
rect 61175 -910 61375 -825
rect 61525 -785 61725 -710
rect 61525 -825 61605 -785
rect 61645 -825 61725 -785
rect 61525 -910 61725 -825
rect 52075 -1135 52275 -1060
rect 52075 -1175 52155 -1135
rect 52195 -1175 52275 -1135
rect 52075 -1260 52275 -1175
rect 52425 -1135 52625 -1060
rect 52425 -1175 52505 -1135
rect 52545 -1175 52625 -1135
rect 52425 -1260 52625 -1175
rect 52775 -1135 52975 -1060
rect 52775 -1175 52855 -1135
rect 52895 -1175 52975 -1135
rect 52775 -1260 52975 -1175
rect 53125 -1135 53325 -1060
rect 53125 -1175 53205 -1135
rect 53245 -1175 53325 -1135
rect 53125 -1260 53325 -1175
rect 53475 -1135 53675 -1060
rect 53475 -1175 53555 -1135
rect 53595 -1175 53675 -1135
rect 53475 -1260 53675 -1175
rect 53825 -1135 54025 -1060
rect 53825 -1175 53905 -1135
rect 53945 -1175 54025 -1135
rect 53825 -1260 54025 -1175
rect 54175 -1135 54375 -1060
rect 54175 -1175 54255 -1135
rect 54295 -1175 54375 -1135
rect 54175 -1260 54375 -1175
rect 54525 -1135 54725 -1060
rect 54525 -1175 54605 -1135
rect 54645 -1175 54725 -1135
rect 54525 -1260 54725 -1175
rect 54875 -1135 55075 -1060
rect 54875 -1175 54955 -1135
rect 54995 -1175 55075 -1135
rect 54875 -1260 55075 -1175
rect 55225 -1135 55425 -1060
rect 55225 -1175 55305 -1135
rect 55345 -1175 55425 -1135
rect 55225 -1260 55425 -1175
rect 55575 -1135 55775 -1060
rect 55575 -1175 55655 -1135
rect 55695 -1175 55775 -1135
rect 55575 -1260 55775 -1175
rect 55925 -1135 56125 -1060
rect 55925 -1175 56005 -1135
rect 56045 -1175 56125 -1135
rect 55925 -1260 56125 -1175
rect 56275 -1135 56475 -1060
rect 56275 -1175 56355 -1135
rect 56395 -1175 56475 -1135
rect 56275 -1260 56475 -1175
rect 56625 -1135 56825 -1060
rect 56625 -1175 56705 -1135
rect 56745 -1175 56825 -1135
rect 56625 -1260 56825 -1175
rect 56975 -1135 57175 -1060
rect 56975 -1175 57055 -1135
rect 57095 -1175 57175 -1135
rect 56975 -1260 57175 -1175
rect 57325 -1135 57525 -1060
rect 57325 -1175 57405 -1135
rect 57445 -1175 57525 -1135
rect 57325 -1260 57525 -1175
rect 57675 -1135 57875 -1060
rect 57675 -1175 57755 -1135
rect 57795 -1175 57875 -1135
rect 57675 -1260 57875 -1175
rect 58025 -1135 58225 -1060
rect 58025 -1175 58105 -1135
rect 58145 -1175 58225 -1135
rect 58025 -1260 58225 -1175
rect 58375 -1135 58575 -1060
rect 58375 -1175 58455 -1135
rect 58495 -1175 58575 -1135
rect 58375 -1260 58575 -1175
rect 58725 -1135 58925 -1060
rect 58725 -1175 58805 -1135
rect 58845 -1175 58925 -1135
rect 58725 -1260 58925 -1175
rect 59075 -1135 59275 -1060
rect 59075 -1175 59155 -1135
rect 59195 -1175 59275 -1135
rect 59075 -1260 59275 -1175
rect 59425 -1135 59625 -1060
rect 59425 -1175 59505 -1135
rect 59545 -1175 59625 -1135
rect 59425 -1260 59625 -1175
rect 59775 -1135 59975 -1060
rect 59775 -1175 59855 -1135
rect 59895 -1175 59975 -1135
rect 59775 -1260 59975 -1175
rect 60125 -1135 60325 -1060
rect 60125 -1175 60205 -1135
rect 60245 -1175 60325 -1135
rect 60125 -1260 60325 -1175
rect 60475 -1135 60675 -1060
rect 60475 -1175 60555 -1135
rect 60595 -1175 60675 -1135
rect 60475 -1260 60675 -1175
rect 60825 -1135 61025 -1060
rect 60825 -1175 60905 -1135
rect 60945 -1175 61025 -1135
rect 60825 -1260 61025 -1175
rect 61175 -1135 61375 -1060
rect 61175 -1175 61255 -1135
rect 61295 -1175 61375 -1135
rect 61175 -1260 61375 -1175
rect 61525 -1135 61725 -1060
rect 61525 -1175 61605 -1135
rect 61645 -1175 61725 -1135
rect 61525 -1260 61725 -1175
<< mimcapcontact >>
rect 52155 5475 52195 5515
rect 52505 5475 52545 5515
rect 52855 5475 52895 5515
rect 53205 5475 53245 5515
rect 53555 5475 53595 5515
rect 53905 5475 53945 5515
rect 54255 5475 54295 5515
rect 54605 5475 54645 5515
rect 54955 5475 54995 5515
rect 55305 5475 55345 5515
rect 55655 5475 55695 5515
rect 56005 5475 56045 5515
rect 56355 5475 56395 5515
rect 56705 5475 56745 5515
rect 57055 5475 57095 5515
rect 57405 5475 57445 5515
rect 57755 5475 57795 5515
rect 58105 5475 58145 5515
rect 58455 5475 58495 5515
rect 58805 5475 58845 5515
rect 59155 5475 59195 5515
rect 59505 5475 59545 5515
rect 59855 5475 59895 5515
rect 60205 5475 60245 5515
rect 60555 5475 60595 5515
rect 60905 5475 60945 5515
rect 61255 5475 61295 5515
rect 61605 5475 61645 5515
rect 52155 5125 52195 5165
rect 52505 5125 52545 5165
rect 52855 5125 52895 5165
rect 53205 5125 53245 5165
rect 53555 5125 53595 5165
rect 53905 5125 53945 5165
rect 54255 5125 54295 5165
rect 54605 5125 54645 5165
rect 54955 5125 54995 5165
rect 55305 5115 55345 5155
rect 55655 5115 55695 5155
rect 58105 5115 58145 5155
rect 58455 5115 58495 5155
rect 58805 5125 58845 5165
rect 59155 5125 59195 5165
rect 59505 5125 59545 5165
rect 59855 5125 59895 5165
rect 60205 5125 60245 5165
rect 60555 5125 60595 5165
rect 60905 5125 60945 5165
rect 61255 5125 61295 5165
rect 61605 5125 61645 5165
rect 52155 4775 52195 4815
rect 52505 4775 52545 4815
rect 52855 4775 52895 4815
rect 53205 4775 53245 4815
rect 53555 4775 53595 4815
rect 53905 4775 53945 4815
rect 54255 4775 54295 4815
rect 54605 4775 54645 4815
rect 54955 4775 54995 4815
rect 55305 4765 55345 4805
rect 58455 4765 58495 4805
rect 58805 4775 58845 4815
rect 59155 4775 59195 4815
rect 59505 4775 59545 4815
rect 59855 4775 59895 4815
rect 60205 4775 60245 4815
rect 60555 4775 60595 4815
rect 60905 4775 60945 4815
rect 61255 4775 61295 4815
rect 61605 4775 61645 4815
rect 52155 4425 52195 4465
rect 52505 4425 52545 4465
rect 52855 4425 52895 4465
rect 53205 4425 53245 4465
rect 53555 4425 53595 4465
rect 60205 4425 60245 4465
rect 60555 4425 60595 4465
rect 60905 4425 60945 4465
rect 61255 4425 61295 4465
rect 61605 4425 61645 4465
rect 52155 4075 52195 4115
rect 52505 4075 52545 4115
rect 52855 4075 52895 4115
rect 53205 4075 53245 4115
rect 53555 4075 53595 4115
rect 60205 4075 60245 4115
rect 60555 4075 60595 4115
rect 60905 4075 60945 4115
rect 61255 4075 61295 4115
rect 61605 4075 61645 4115
rect 52155 3725 52195 3765
rect 52505 3725 52545 3765
rect 52855 3725 52895 3765
rect 53205 3725 53245 3765
rect 53555 3725 53595 3765
rect 60205 3725 60245 3765
rect 60555 3725 60595 3765
rect 60905 3725 60945 3765
rect 61255 3725 61295 3765
rect 61605 3725 61645 3765
rect 52155 3375 52195 3415
rect 52505 3375 52545 3415
rect 52855 3375 52895 3415
rect 53205 3375 53245 3415
rect 53555 3375 53595 3415
rect 60205 3375 60245 3415
rect 60555 3375 60595 3415
rect 60905 3375 60945 3415
rect 61255 3375 61295 3415
rect 61605 3375 61645 3415
rect 52155 3025 52195 3065
rect 52505 3025 52545 3065
rect 52855 3025 52895 3065
rect 53205 3025 53245 3065
rect 53555 3025 53595 3065
rect 60205 3025 60245 3065
rect 60555 3025 60595 3065
rect 60905 3025 60945 3065
rect 61255 3025 61295 3065
rect 61605 3025 61645 3065
rect 52155 2675 52195 2715
rect 52505 2675 52545 2715
rect 52855 2675 52895 2715
rect 53205 2675 53245 2715
rect 53555 2675 53595 2715
rect 60205 2675 60245 2715
rect 60555 2675 60595 2715
rect 60905 2675 60945 2715
rect 61255 2675 61295 2715
rect 61605 2675 61645 2715
rect 52155 2325 52195 2365
rect 52505 2325 52545 2365
rect 52855 2325 52895 2365
rect 53205 2325 53245 2365
rect 53555 2325 53595 2365
rect 60205 2325 60245 2365
rect 60555 2325 60595 2365
rect 60905 2325 60945 2365
rect 61255 2325 61295 2365
rect 61605 2325 61645 2365
rect 52155 1975 52195 2015
rect 52505 1975 52545 2015
rect 52855 1975 52895 2015
rect 53205 1975 53245 2015
rect 53555 1975 53595 2015
rect 60205 1975 60245 2015
rect 60555 1975 60595 2015
rect 60905 1975 60945 2015
rect 61255 1975 61295 2015
rect 61605 1975 61645 2015
rect 52155 1625 52195 1665
rect 52505 1625 52545 1665
rect 52855 1625 52895 1665
rect 53205 1625 53245 1665
rect 53555 1625 53595 1665
rect 60205 1625 60245 1665
rect 60555 1625 60595 1665
rect 60905 1625 60945 1665
rect 61255 1625 61295 1665
rect 61605 1625 61645 1665
rect 52155 1275 52195 1315
rect 52505 1275 52545 1315
rect 52855 1275 52895 1315
rect 53205 1275 53245 1315
rect 53555 1275 53595 1315
rect 60205 1275 60245 1315
rect 60555 1275 60595 1315
rect 60905 1275 60945 1315
rect 61255 1275 61295 1315
rect 61605 1275 61645 1315
rect 52155 925 52195 965
rect 52505 925 52545 965
rect 52855 925 52895 965
rect 53205 925 53245 965
rect 53555 925 53595 965
rect 60205 925 60245 965
rect 60555 925 60595 965
rect 60905 925 60945 965
rect 61255 925 61295 965
rect 61605 925 61645 965
rect 52155 575 52195 615
rect 52505 575 52545 615
rect 52855 575 52895 615
rect 53205 575 53245 615
rect 53555 575 53595 615
rect 60205 575 60245 615
rect 60555 575 60595 615
rect 60905 575 60945 615
rect 61255 575 61295 615
rect 61605 575 61645 615
rect 52155 225 52195 265
rect 52505 225 52545 265
rect 52855 225 52895 265
rect 53205 225 53245 265
rect 53555 225 53595 265
rect 60205 225 60245 265
rect 60555 225 60595 265
rect 60905 225 60945 265
rect 61255 225 61295 265
rect 61605 225 61645 265
rect 52155 -125 52195 -85
rect 52505 -125 52545 -85
rect 52855 -125 52895 -85
rect 53205 -125 53245 -85
rect 53555 -125 53595 -85
rect 60205 -125 60245 -85
rect 60555 -125 60595 -85
rect 60905 -125 60945 -85
rect 61255 -125 61295 -85
rect 61605 -125 61645 -85
rect 52155 -475 52195 -435
rect 52505 -475 52545 -435
rect 52855 -475 52895 -435
rect 53205 -475 53245 -435
rect 53555 -475 53595 -435
rect 60205 -475 60245 -435
rect 60555 -475 60595 -435
rect 60905 -475 60945 -435
rect 61255 -475 61295 -435
rect 61605 -475 61645 -435
rect 52155 -825 52195 -785
rect 52505 -825 52545 -785
rect 52855 -825 52895 -785
rect 53205 -825 53245 -785
rect 53555 -825 53595 -785
rect 53905 -825 53945 -785
rect 54255 -825 54295 -785
rect 54605 -825 54645 -785
rect 54955 -825 54995 -785
rect 55305 -825 55345 -785
rect 55655 -825 55695 -785
rect 56005 -825 56045 -785
rect 56355 -825 56395 -785
rect 56705 -825 56745 -785
rect 57055 -825 57095 -785
rect 57405 -825 57445 -785
rect 57755 -825 57795 -785
rect 58105 -825 58145 -785
rect 58455 -825 58495 -785
rect 58805 -825 58845 -785
rect 59155 -825 59195 -785
rect 59505 -825 59545 -785
rect 59855 -825 59895 -785
rect 60205 -825 60245 -785
rect 60555 -825 60595 -785
rect 60905 -825 60945 -785
rect 61255 -825 61295 -785
rect 61605 -825 61645 -785
rect 52155 -1175 52195 -1135
rect 52505 -1175 52545 -1135
rect 52855 -1175 52895 -1135
rect 53205 -1175 53245 -1135
rect 53555 -1175 53595 -1135
rect 53905 -1175 53945 -1135
rect 54255 -1175 54295 -1135
rect 54605 -1175 54645 -1135
rect 54955 -1175 54995 -1135
rect 55305 -1175 55345 -1135
rect 55655 -1175 55695 -1135
rect 56005 -1175 56045 -1135
rect 56355 -1175 56395 -1135
rect 56705 -1175 56745 -1135
rect 57055 -1175 57095 -1135
rect 57405 -1175 57445 -1135
rect 57755 -1175 57795 -1135
rect 58105 -1175 58145 -1135
rect 58455 -1175 58495 -1135
rect 58805 -1175 58845 -1135
rect 59155 -1175 59195 -1135
rect 59505 -1175 59545 -1135
rect 59855 -1175 59895 -1135
rect 60205 -1175 60245 -1135
rect 60555 -1175 60595 -1135
rect 60905 -1175 60945 -1135
rect 61255 -1175 61295 -1135
rect 61605 -1175 61645 -1135
<< metal4 >>
rect 52150 5515 56750 5520
rect 52150 5475 52155 5515
rect 52195 5475 52505 5515
rect 52545 5475 52855 5515
rect 52895 5475 53205 5515
rect 53245 5475 53555 5515
rect 53595 5475 53905 5515
rect 53945 5475 54255 5515
rect 54295 5475 54605 5515
rect 54645 5475 54955 5515
rect 54995 5475 55305 5515
rect 55345 5475 55655 5515
rect 55695 5475 56005 5515
rect 56045 5475 56355 5515
rect 56395 5475 56705 5515
rect 56745 5475 56750 5515
rect 52150 5470 56750 5475
rect 57050 5515 61650 5520
rect 57050 5475 57055 5515
rect 57095 5475 57405 5515
rect 57445 5475 57755 5515
rect 57795 5475 58105 5515
rect 58145 5475 58455 5515
rect 58495 5475 58805 5515
rect 58845 5475 59155 5515
rect 59195 5475 59505 5515
rect 59545 5475 59855 5515
rect 59895 5475 60205 5515
rect 60245 5475 60555 5515
rect 60595 5475 60905 5515
rect 60945 5475 61255 5515
rect 61295 5475 61605 5515
rect 61645 5475 61650 5515
rect 57050 5470 61650 5475
rect 52850 5170 52900 5470
rect 52150 5165 53600 5170
rect 52150 5125 52155 5165
rect 52195 5125 52505 5165
rect 52545 5125 52855 5165
rect 52895 5125 53205 5165
rect 53245 5125 53555 5165
rect 53595 5125 53600 5165
rect 52150 5120 53600 5125
rect 53900 5165 53950 5470
rect 53900 5125 53905 5165
rect 53945 5125 53950 5165
rect 52850 4820 52900 5120
rect 52150 4815 53600 4820
rect 52150 4775 52155 4815
rect 52195 4775 52505 4815
rect 52545 4775 52855 4815
rect 52895 4775 53205 4815
rect 53245 4775 53555 4815
rect 53595 4775 53600 4815
rect 52150 4770 53600 4775
rect 53900 4815 53950 5125
rect 53900 4775 53905 4815
rect 53945 4775 53950 4815
rect 53900 4770 53950 4775
rect 54250 5165 54300 5470
rect 54250 5125 54255 5165
rect 54295 5125 54300 5165
rect 54250 4815 54300 5125
rect 54250 4775 54255 4815
rect 54295 4775 54300 4815
rect 54250 4770 54300 4775
rect 54600 5165 54650 5470
rect 54600 5125 54605 5165
rect 54645 5125 54650 5165
rect 54600 4815 54650 5125
rect 54600 4775 54605 4815
rect 54645 4775 54650 4815
rect 54600 4770 54650 4775
rect 54950 5165 55000 5470
rect 54950 5125 54955 5165
rect 54995 5125 55000 5165
rect 54950 4815 55000 5125
rect 54950 4775 54955 4815
rect 54995 4775 55000 4815
rect 54950 4770 55000 4775
rect 55300 5155 55350 5470
rect 55300 5115 55305 5155
rect 55345 5115 55350 5155
rect 55300 4805 55350 5115
rect 55650 5155 55700 5470
rect 55650 5115 55655 5155
rect 55695 5115 55700 5155
rect 55650 5110 55700 5115
rect 58100 5155 58150 5470
rect 58100 5115 58105 5155
rect 58145 5115 58150 5155
rect 58100 5110 58150 5115
rect 58450 5155 58500 5470
rect 58450 5115 58455 5155
rect 58495 5115 58500 5155
rect 52850 4470 52900 4770
rect 55300 4765 55305 4805
rect 55345 4765 55350 4805
rect 55300 4760 55350 4765
rect 58450 4805 58500 5115
rect 58450 4765 58455 4805
rect 58495 4765 58500 4805
rect 58800 5165 58850 5470
rect 58800 5125 58805 5165
rect 58845 5125 58850 5165
rect 58800 4815 58850 5125
rect 58800 4775 58805 4815
rect 58845 4775 58850 4815
rect 58800 4770 58850 4775
rect 59150 5165 59200 5470
rect 59150 5125 59155 5165
rect 59195 5125 59200 5165
rect 59150 4815 59200 5125
rect 59150 4775 59155 4815
rect 59195 4775 59200 4815
rect 59150 4770 59200 4775
rect 59500 5165 59550 5470
rect 59500 5125 59505 5165
rect 59545 5125 59550 5165
rect 59500 4815 59550 5125
rect 59500 4775 59505 4815
rect 59545 4775 59550 4815
rect 59500 4770 59550 4775
rect 59850 5165 59900 5470
rect 60900 5170 60950 5470
rect 59850 5125 59855 5165
rect 59895 5125 59900 5165
rect 59850 4815 59900 5125
rect 60200 5165 61650 5170
rect 60200 5125 60205 5165
rect 60245 5125 60555 5165
rect 60595 5125 60905 5165
rect 60945 5125 61255 5165
rect 61295 5125 61605 5165
rect 61645 5125 61650 5165
rect 60200 5120 61650 5125
rect 60900 4820 60950 5120
rect 59850 4775 59855 4815
rect 59895 4775 59900 4815
rect 59850 4770 59900 4775
rect 60200 4815 61650 4820
rect 60200 4775 60205 4815
rect 60245 4775 60555 4815
rect 60595 4775 60905 4815
rect 60945 4775 61255 4815
rect 61295 4775 61605 4815
rect 61645 4775 61650 4815
rect 60200 4770 61650 4775
rect 58450 4760 58500 4765
rect 60900 4470 60950 4770
rect 52150 4465 53600 4470
rect 52150 4425 52155 4465
rect 52195 4425 52505 4465
rect 52545 4425 52855 4465
rect 52895 4425 53205 4465
rect 53245 4425 53555 4465
rect 53595 4425 53600 4465
rect 52150 4420 53600 4425
rect 60200 4465 61650 4470
rect 60200 4425 60205 4465
rect 60245 4425 60555 4465
rect 60595 4425 60905 4465
rect 60945 4425 61255 4465
rect 61295 4425 61605 4465
rect 61645 4425 61650 4465
rect 60200 4420 61650 4425
rect 52850 4120 52900 4420
rect 60900 4120 60950 4420
rect 52150 4115 53600 4120
rect 52150 4075 52155 4115
rect 52195 4075 52505 4115
rect 52545 4075 52855 4115
rect 52895 4075 53205 4115
rect 53245 4075 53555 4115
rect 53595 4075 53600 4115
rect 52150 4070 53600 4075
rect 60200 4115 61650 4120
rect 60200 4075 60205 4115
rect 60245 4075 60555 4115
rect 60595 4075 60905 4115
rect 60945 4075 61255 4115
rect 61295 4075 61605 4115
rect 61645 4075 61650 4115
rect 60200 4070 61650 4075
rect 52850 3770 52900 4070
rect 60900 3770 60950 4070
rect 52150 3765 53600 3770
rect 52150 3725 52155 3765
rect 52195 3725 52505 3765
rect 52545 3725 52855 3765
rect 52895 3725 53205 3765
rect 53245 3725 53555 3765
rect 53595 3725 53600 3765
rect 52150 3720 53600 3725
rect 60200 3765 61650 3770
rect 60200 3725 60205 3765
rect 60245 3725 60555 3765
rect 60595 3725 60905 3765
rect 60945 3725 61255 3765
rect 61295 3725 61605 3765
rect 61645 3725 61650 3765
rect 60200 3720 61650 3725
rect 52850 3420 52900 3720
rect 60900 3420 60950 3720
rect 52150 3415 53600 3420
rect 52150 3375 52155 3415
rect 52195 3375 52505 3415
rect 52545 3375 52855 3415
rect 52895 3375 53205 3415
rect 53245 3375 53555 3415
rect 53595 3375 53600 3415
rect 52150 3370 53600 3375
rect 60200 3415 61650 3420
rect 60200 3375 60205 3415
rect 60245 3375 60555 3415
rect 60595 3375 60905 3415
rect 60945 3375 61255 3415
rect 61295 3375 61605 3415
rect 61645 3375 61650 3415
rect 60200 3370 61650 3375
rect 52850 3070 52900 3370
rect 60900 3070 60950 3370
rect 52150 3065 53600 3070
rect 52150 3025 52155 3065
rect 52195 3025 52505 3065
rect 52545 3025 52855 3065
rect 52895 3025 53205 3065
rect 53245 3025 53555 3065
rect 53595 3025 53600 3065
rect 52150 3020 53600 3025
rect 60200 3065 61650 3070
rect 60200 3025 60205 3065
rect 60245 3025 60555 3065
rect 60595 3025 60905 3065
rect 60945 3025 61255 3065
rect 61295 3025 61605 3065
rect 61645 3025 61650 3065
rect 60200 3020 61650 3025
rect 52850 2720 52900 3020
rect 60900 2720 60950 3020
rect 52150 2715 53600 2720
rect 52150 2675 52155 2715
rect 52195 2675 52505 2715
rect 52545 2675 52855 2715
rect 52895 2675 53205 2715
rect 53245 2675 53555 2715
rect 53595 2675 53600 2715
rect 52150 2670 53600 2675
rect 60200 2715 61650 2720
rect 60200 2675 60205 2715
rect 60245 2675 60555 2715
rect 60595 2675 60905 2715
rect 60945 2675 61255 2715
rect 61295 2675 61605 2715
rect 61645 2675 61650 2715
rect 60200 2670 61650 2675
rect 52850 2370 52900 2670
rect 60900 2370 60950 2670
rect 52150 2365 53600 2370
rect 52150 2325 52155 2365
rect 52195 2325 52505 2365
rect 52545 2325 52855 2365
rect 52895 2325 53205 2365
rect 53245 2325 53555 2365
rect 53595 2325 53600 2365
rect 52150 2320 53600 2325
rect 60200 2365 61650 2370
rect 60200 2325 60205 2365
rect 60245 2325 60555 2365
rect 60595 2325 60905 2365
rect 60945 2325 61255 2365
rect 61295 2325 61605 2365
rect 61645 2325 61650 2365
rect 60200 2320 61650 2325
rect 52850 2020 52900 2320
rect 60900 2020 60950 2320
rect 52150 2015 53600 2020
rect 52150 1975 52155 2015
rect 52195 1975 52505 2015
rect 52545 1975 52855 2015
rect 52895 1975 53205 2015
rect 53245 1975 53555 2015
rect 53595 1975 53600 2015
rect 52150 1970 53600 1975
rect 60200 2015 61650 2020
rect 60200 1975 60205 2015
rect 60245 1975 60555 2015
rect 60595 1975 60905 2015
rect 60945 1975 61255 2015
rect 61295 1975 61605 2015
rect 61645 1975 61650 2015
rect 60200 1970 61650 1975
rect 52850 1670 52900 1970
rect 53550 1715 54320 1720
rect 53550 1675 54075 1715
rect 54115 1675 54125 1715
rect 54165 1675 54175 1715
rect 54215 1675 54225 1715
rect 54265 1675 54275 1715
rect 54315 1675 54320 1715
rect 53550 1670 54320 1675
rect 52150 1665 54320 1670
rect 52150 1625 52155 1665
rect 52195 1625 52505 1665
rect 52545 1625 52855 1665
rect 52895 1625 53205 1665
rect 53245 1625 53555 1665
rect 53595 1625 54075 1665
rect 54115 1625 54125 1665
rect 54165 1625 54175 1665
rect 54215 1625 54225 1665
rect 54265 1625 54275 1665
rect 54315 1625 54320 1665
rect 52150 1620 54320 1625
rect 52850 1320 52900 1620
rect 53550 1615 54320 1620
rect 53550 1575 54075 1615
rect 54115 1575 54125 1615
rect 54165 1575 54175 1615
rect 54215 1575 54225 1615
rect 54265 1575 54275 1615
rect 54315 1575 54320 1615
rect 53550 1570 54320 1575
rect 59480 1715 60255 1720
rect 59480 1675 59485 1715
rect 59525 1675 59535 1715
rect 59575 1675 59585 1715
rect 59625 1675 59635 1715
rect 59675 1675 59685 1715
rect 59725 1675 60255 1715
rect 59480 1670 60255 1675
rect 60900 1670 60950 1970
rect 59480 1665 61650 1670
rect 59480 1625 59485 1665
rect 59525 1625 59535 1665
rect 59575 1625 59585 1665
rect 59625 1625 59635 1665
rect 59675 1625 59685 1665
rect 59725 1625 60205 1665
rect 60245 1625 60555 1665
rect 60595 1625 60905 1665
rect 60945 1625 61255 1665
rect 61295 1625 61605 1665
rect 61645 1625 61650 1665
rect 59480 1620 61650 1625
rect 59480 1615 60255 1620
rect 59480 1575 59485 1615
rect 59525 1575 59535 1615
rect 59575 1575 59585 1615
rect 59625 1575 59635 1615
rect 59675 1575 59685 1615
rect 59725 1575 60255 1615
rect 59480 1570 60255 1575
rect 60900 1320 60950 1620
rect 52150 1315 53600 1320
rect 52150 1275 52155 1315
rect 52195 1275 52505 1315
rect 52545 1275 52855 1315
rect 52895 1275 53205 1315
rect 53245 1275 53555 1315
rect 53595 1275 53600 1315
rect 52150 1270 53600 1275
rect 60200 1315 61650 1320
rect 60200 1275 60205 1315
rect 60245 1275 60555 1315
rect 60595 1275 60905 1315
rect 60945 1275 61255 1315
rect 61295 1275 61605 1315
rect 61645 1275 61650 1315
rect 60200 1270 61650 1275
rect 52850 970 52900 1270
rect 60900 970 60950 1270
rect 52150 965 53600 970
rect 52150 925 52155 965
rect 52195 925 52505 965
rect 52545 925 52855 965
rect 52895 925 53205 965
rect 53245 925 53555 965
rect 53595 925 53600 965
rect 52150 920 53600 925
rect 60200 965 61650 970
rect 60200 925 60205 965
rect 60245 925 60555 965
rect 60595 925 60905 965
rect 60945 925 61255 965
rect 61295 925 61605 965
rect 61645 925 61650 965
rect 60200 920 61650 925
rect 52850 620 52900 920
rect 60900 620 60950 920
rect 52150 615 53600 620
rect 52150 575 52155 615
rect 52195 575 52505 615
rect 52545 575 52855 615
rect 52895 575 53205 615
rect 53245 575 53555 615
rect 53595 575 53600 615
rect 52150 570 53600 575
rect 60200 615 61650 620
rect 60200 575 60205 615
rect 60245 575 60555 615
rect 60595 575 60905 615
rect 60945 575 61255 615
rect 61295 575 61605 615
rect 61645 575 61650 615
rect 60200 570 61650 575
rect 52850 270 52900 570
rect 60900 270 60950 570
rect 52150 265 53600 270
rect 52150 225 52155 265
rect 52195 225 52505 265
rect 52545 225 52855 265
rect 52895 225 53205 265
rect 53245 225 53555 265
rect 53595 225 53600 265
rect 52150 220 53600 225
rect 60200 265 61650 270
rect 60200 225 60205 265
rect 60245 225 60555 265
rect 60595 225 60905 265
rect 60945 225 61255 265
rect 61295 225 61605 265
rect 61645 225 61650 265
rect 60200 220 61650 225
rect 52850 -80 52900 220
rect 60900 -80 60950 220
rect 52150 -85 53600 -80
rect 52150 -125 52155 -85
rect 52195 -125 52505 -85
rect 52545 -125 52855 -85
rect 52895 -125 53205 -85
rect 53245 -125 53555 -85
rect 53595 -125 53600 -85
rect 52150 -130 53600 -125
rect 60200 -85 61650 -80
rect 60200 -125 60205 -85
rect 60245 -125 60555 -85
rect 60595 -125 60905 -85
rect 60945 -125 61255 -85
rect 61295 -125 61605 -85
rect 61645 -125 61650 -85
rect 60200 -130 61650 -125
rect 52850 -430 52900 -130
rect 60900 -430 60950 -130
rect 52150 -435 53600 -430
rect 52150 -475 52155 -435
rect 52195 -475 52505 -435
rect 52545 -475 52855 -435
rect 52895 -475 53205 -435
rect 53245 -475 53555 -435
rect 53595 -475 53600 -435
rect 52150 -480 53600 -475
rect 60200 -435 61650 -430
rect 60200 -475 60205 -435
rect 60245 -475 60555 -435
rect 60595 -475 60905 -435
rect 60945 -475 61255 -435
rect 61295 -475 61605 -435
rect 61645 -475 61650 -435
rect 60200 -480 61650 -475
rect 52850 -780 52900 -480
rect 60900 -780 60950 -480
rect 52150 -785 56750 -780
rect 52150 -825 52155 -785
rect 52195 -825 52505 -785
rect 52545 -825 52855 -785
rect 52895 -825 53205 -785
rect 53245 -825 53555 -785
rect 53595 -825 53905 -785
rect 53945 -825 54255 -785
rect 54295 -825 54605 -785
rect 54645 -825 54955 -785
rect 54995 -825 55305 -785
rect 55345 -825 55655 -785
rect 55695 -825 56005 -785
rect 56045 -825 56355 -785
rect 56395 -825 56705 -785
rect 56745 -825 56750 -785
rect 52150 -830 56750 -825
rect 52850 -1130 52900 -830
rect 52150 -1135 52900 -1130
rect 52150 -1175 52155 -1135
rect 52195 -1175 52505 -1135
rect 52545 -1175 52855 -1135
rect 52895 -1175 52900 -1135
rect 52150 -1180 52900 -1175
rect 53200 -1135 53250 -830
rect 53200 -1175 53205 -1135
rect 53245 -1175 53250 -1135
rect 53200 -1180 53250 -1175
rect 53550 -1135 53600 -830
rect 53550 -1175 53555 -1135
rect 53595 -1175 53600 -1135
rect 53550 -1180 53600 -1175
rect 53900 -1135 53950 -830
rect 53900 -1175 53905 -1135
rect 53945 -1175 53950 -1135
rect 53900 -1180 53950 -1175
rect 54250 -1135 54300 -830
rect 54250 -1175 54255 -1135
rect 54295 -1175 54300 -1135
rect 54250 -1180 54300 -1175
rect 54600 -1135 54650 -830
rect 54600 -1175 54605 -1135
rect 54645 -1175 54650 -1135
rect 54600 -1180 54650 -1175
rect 54950 -1135 55000 -830
rect 54950 -1175 54955 -1135
rect 54995 -1175 55000 -1135
rect 54950 -1180 55000 -1175
rect 55300 -1135 55350 -830
rect 55300 -1175 55305 -1135
rect 55345 -1175 55350 -1135
rect 55300 -1180 55350 -1175
rect 55650 -1135 55700 -830
rect 55650 -1175 55655 -1135
rect 55695 -1175 55700 -1135
rect 55650 -1180 55700 -1175
rect 56000 -1135 56050 -830
rect 56000 -1175 56005 -1135
rect 56045 -1175 56050 -1135
rect 56000 -1180 56050 -1175
rect 56350 -1135 56400 -830
rect 56350 -1175 56355 -1135
rect 56395 -1175 56400 -1135
rect 56350 -1180 56400 -1175
rect 56700 -1135 56750 -830
rect 56700 -1175 56705 -1135
rect 56745 -1175 56750 -1135
rect 56700 -1180 56750 -1175
rect 57050 -785 61650 -780
rect 57050 -825 57055 -785
rect 57095 -825 57405 -785
rect 57445 -825 57755 -785
rect 57795 -825 58105 -785
rect 58145 -825 58455 -785
rect 58495 -825 58805 -785
rect 58845 -825 59155 -785
rect 59195 -825 59505 -785
rect 59545 -825 59855 -785
rect 59895 -825 60205 -785
rect 60245 -825 60555 -785
rect 60595 -825 60905 -785
rect 60945 -825 61255 -785
rect 61295 -825 61605 -785
rect 61645 -825 61650 -785
rect 57050 -830 61650 -825
rect 57050 -1135 57100 -830
rect 57050 -1175 57055 -1135
rect 57095 -1175 57100 -1135
rect 57050 -1180 57100 -1175
rect 57400 -1135 57450 -830
rect 57400 -1175 57405 -1135
rect 57445 -1175 57450 -1135
rect 57400 -1180 57450 -1175
rect 57750 -1135 57800 -830
rect 57750 -1175 57755 -1135
rect 57795 -1175 57800 -1135
rect 57750 -1180 57800 -1175
rect 58100 -1135 58150 -830
rect 58100 -1175 58105 -1135
rect 58145 -1175 58150 -1135
rect 58100 -1180 58150 -1175
rect 58450 -1135 58500 -830
rect 58450 -1175 58455 -1135
rect 58495 -1175 58500 -1135
rect 58450 -1180 58500 -1175
rect 58800 -1135 58850 -830
rect 58800 -1175 58805 -1135
rect 58845 -1175 58850 -1135
rect 58800 -1180 58850 -1175
rect 59150 -1135 59200 -830
rect 59150 -1175 59155 -1135
rect 59195 -1175 59200 -1135
rect 59150 -1180 59200 -1175
rect 59500 -1135 59550 -830
rect 59500 -1175 59505 -1135
rect 59545 -1175 59550 -1135
rect 59500 -1180 59550 -1175
rect 59850 -1135 59900 -830
rect 59850 -1175 59855 -1135
rect 59895 -1175 59900 -1135
rect 59850 -1180 59900 -1175
rect 60200 -1135 60250 -830
rect 60200 -1175 60205 -1135
rect 60245 -1175 60250 -1135
rect 60200 -1180 60250 -1175
rect 60550 -1135 60600 -830
rect 60550 -1175 60555 -1135
rect 60595 -1175 60600 -1135
rect 60550 -1180 60600 -1175
rect 60900 -1130 60950 -830
rect 60900 -1135 61650 -1130
rect 60900 -1175 60905 -1135
rect 60945 -1175 61255 -1135
rect 61295 -1175 61605 -1135
rect 61645 -1175 61650 -1135
rect 60900 -1180 61650 -1175
<< labels >>
flabel metal2 57365 5060 57365 5060 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 56455 5060 56455 5060 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 56800 -235 56800 -235 1 FreeSans 240 0 0 80 Vb1_2
flabel metal2 56460 -90 56460 -90 1 FreeSans 240 0 0 80 V_p_mir
flabel metal2 57000 3510 57000 3510 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56855 3545 56855 3545 5 FreeSans 200 0 0 -80 Vb2
port 5 s
flabel metal2 57950 4070 57950 4070 5 FreeSans 240 0 0 -80 VD3
flabel metal2 55865 4070 55865 4070 5 FreeSans 240 0 0 -80 VD4
flabel metal1 56945 655 56945 655 7 FreeSans 240 0 -80 0 V_tail_gate
port 11 w
flabel metal2 57770 1280 57770 1280 3 FreeSans 240 0 80 0 VIN-
flabel metal2 56030 1280 56030 1280 7 FreeSans 240 0 -80 0 VIN+
flabel metal1 57430 1325 57430 1325 3 FreeSans 240 0 80 0 VD1
flabel metal1 56370 1325 56370 1325 7 FreeSans 240 0 -80 0 VD2
flabel metal2 56900 1960 56900 1960 5 FreeSans 240 0 0 -80 Vb1
flabel metal2 57455 2465 57455 2465 7 FreeSans 240 0 -80 0 X
flabel metal2 57525 2665 57525 2665 1 FreeSans 240 0 0 80 err_amp_out
flabel metal2 57000 2710 57000 2710 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal2 57125 2875 57125 2875 3 FreeSans 240 0 80 0 V_err_gate
port 13 e
flabel metal2 56365 2815 56365 2815 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal1 56620 3195 56620 3195 7 FreeSans 240 0 -80 0 V_err_mir_p
flabel metal2 57180 3195 57180 3195 3 FreeSans 240 0 80 0 V_err_p
flabel metal2 57580 2775 57580 2775 1 FreeSans 240 0 0 160 V_tot
flabel metal1 56345 2455 56345 2455 3 FreeSans 240 0 80 0 Y
flabel metal3 59545 3435 59545 3435 3 FreeSans 240 0 80 0 cap_res_X
flabel metal3 54255 3435 54255 3435 7 FreeSans 240 0 -80 0 cap_res_Y
flabel metal2 57720 410 57720 410 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal1 57220 440 57220 440 3 FreeSans 240 0 80 0 V_source
flabel metal1 59625 195 59625 195 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 59215 1665 59215 1665 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 59170 1480 59170 1480 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal2 54630 1480 54630 1480 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal2 54585 1665 54585 1665 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal2 54175 195 54175 195 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
<< end >>
