* PEX produced on Sat Feb  1 08:41:07 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from div4.ext - technology: sky130A

.subckt div4 VOUT VIN VDDA GNDA
X0 VDDA.t17 div2.t2 div2_3_1.A.t1 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X1 div2.t1 div2_3_1.C.t4 GNDA.t25 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X2 VDDA.t15 div2.t3 div2_3_2.CLK.t2 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X3 GNDA.t15 div2_3_1.CLK.t3 div2_3_1.C.t2 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X4 div2_3_1.C.t0 div2_3_1.CLK.t4 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X5 div2_3_2.C.t3 div2_3_2.A.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X6 GNDA.t8 div2_3_1.CLK.t5 div2_3_1.C.t1 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 VDDA.t1 VIN.t0 div2_3_1.CLK.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X8 div2_3_1.C.t3 div2_3_1.A.t2 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 GNDA.t17 div2_3_2.CLK.t3 div2_3_2.C.t2 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X10 VOUT.t1 div2_3_2.C.t4 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X11 VOUT.t0 div2_3_2.CLK.t4 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X12 GNDA.t19 div2_3_2.CLK.t5 div2_3_2.C.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X13 div2_3_1.A.t0 div2_3_1.CLK.t6 div2_3_1.B.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X14 div2_3_2.C.t0 div2_3_2.CLK.t6 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 div2_3_2.A.t0 div2_3_2.CLK.t7 div2_3_2.B.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X16 div2_3_1.B.t1 div2.t4 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X17 div2_3_2.B.t1 VOUT.t2 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X18 div2.t0 div2_3_1.CLK.t7 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X19 GNDA.t3 VIN.t1 div2_3_1.CLK.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X20 div2_3_2.CLK.t1 div2.t5 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X21 GNDA.t21 div2.t6 div2_3_2.CLK.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X22 div2_3_1.CLK.t2 VIN.t2 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 VDDA.t11 VOUT.t3 div2_3_2.A.t1 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
R0 div2.t2 div2.t4 819.4
R1 div2.n0 div2.t0 663.801
R2 div2.n0 div2.t2 489.168
R3 div2.t3 div2.t5 401.668
R4 div2.n1 div2.t1 270.12
R5 div2.n2 div2.t3 257.067
R6 div2_3_2.VIN div2.n2 216.9
R7 div2.n2 div2.t6 208.868
R8 div2.n3 div2_3_2.VIN 192.167
R9 div2.n1 div2.n0 67.2005
R10 div2.n3 div2.n1 25.6005
R11 div2_3_1.VOUT div2.n3 4.8005
R12 div2_3_1.A.n0 div2_3_1.A.t1 713.933
R13 div2_3_1.A.n0 div2_3_1.A.t2 314.233
R14 div2_3_1.A.t0 div2_3_1.A.n0 308.2
R15 VDDA.t4 VDDA.t14 2080.95
R16 VDDA.t12 VDDA.t10 1130.95
R17 VDDA.t16 VDDA.t6 1130.95
R18 VDDA.t2 VDDA.n7 927.381
R19 VDDA.n8 VDDA.t18 927.381
R20 VDDA.n6 VDDA.t9 667.62
R21 VDDA.n1 VDDA.t5 663.801
R22 VDDA.n7 VDDA.t8 610.715
R23 VDDA.n8 VDDA.t4 610.715
R24 VDDA.n14 VDDA.n13 594.301
R25 VDDA.n12 VDDA.n11 594.301
R26 VDDA.n3 VDDA.n2 594.301
R27 VDDA.n5 VDDA.n4 594.301
R28 VDDA.t10 VDDA.t2 497.62
R29 VDDA.t14 VDDA.t12 497.62
R30 VDDA.t18 VDDA.t16 497.62
R31 VDDA.t6 VDDA.t0 497.62
R32 VDDA.n7 VDDA.n6 373.781
R33 VDDA.n9 VDDA.n8 370
R34 VDDA.n13 VDDA.t7 78.8005
R35 VDDA.n13 VDDA.t1 78.8005
R36 VDDA.n11 VDDA.t19 78.8005
R37 VDDA.n11 VDDA.t17 78.8005
R38 VDDA.n2 VDDA.t13 78.8005
R39 VDDA.n2 VDDA.t15 78.8005
R40 VDDA.n4 VDDA.t3 78.8005
R41 VDDA.n4 VDDA.t11 78.8005
R42 VDDA.n9 VDDA.n1 12.8005
R43 VDDA.n1 VDDA.n0 9.3005
R44 VDDA.n10 VDDA.n9 9.3005
R45 VDDA.n6 VDDA.n5 3.10124
R46 VDDA VDDA.n0 0.4755
R47 VDDA.n5 VDDA.n3 0.4505
R48 VDDA.n14 VDDA.n12 0.4505
R49 VDDA.n12 VDDA.n10 0.3255
R50 VDDA.n3 VDDA 0.238
R51 VDDA VDDA.n14 0.238
R52 VDDA.n10 VDDA.n0 0.1005
R53 div2_3_1.C.n0 div2_3_1.C.t3 721.4
R54 div2_3_1.C.n1 div2_3_1.C.t4 349.433
R55 div2_3_1.C.n0 div2_3_1.C.t1 276.733
R56 div2_3_1.C.n2 div2_3_1.C.n1 206.333
R57 div2_3_1.C.n1 div2_3_1.C.n0 48.0005
R58 div2_3_1.C.n2 div2_3_1.C.t2 48.0005
R59 div2_3_1.C.t0 div2_3_1.C.n2 48.0005
R60 GNDA.t6 GNDA.t16 4683.87
R61 GNDA.t7 GNDA.t13 4683.87
R62 GNDA.t9 GNDA.n5 3947.35
R63 GNDA.n6 GNDA.t20 2767.74
R64 GNDA.n6 GNDA.t24 2767.74
R65 GNDA.t18 GNDA.t9 1561.29
R66 GNDA.t0 GNDA.t18 1561.29
R67 GNDA.t16 GNDA.t0 1561.29
R68 GNDA.t11 GNDA.t6 1561.29
R69 GNDA.t20 GNDA.t11 1561.29
R70 GNDA.t24 GNDA.t14 1561.29
R71 GNDA.t14 GNDA.t4 1561.29
R72 GNDA.t4 GNDA.t7 1561.29
R73 GNDA.t13 GNDA.t22 1561.29
R74 GNDA.t22 GNDA.t2 1561.29
R75 GNDA.n7 GNDA.n6 1179.3
R76 GNDA.n13 GNDA.n12 194.3
R77 GNDA.n11 GNDA.n10 194.3
R78 GNDA.n9 GNDA.n8 194.3
R79 GNDA.n1 GNDA.n0 194.3
R80 GNDA.n3 GNDA.n2 194.3
R81 GNDA.n5 GNDA.n4 194.3
R82 GNDA.n12 GNDA.t23 48.0005
R83 GNDA.n12 GNDA.t3 48.0005
R84 GNDA.n10 GNDA.t5 48.0005
R85 GNDA.n10 GNDA.t8 48.0005
R86 GNDA.n8 GNDA.t25 48.0005
R87 GNDA.n8 GNDA.t15 48.0005
R88 GNDA.n0 GNDA.t12 48.0005
R89 GNDA.n0 GNDA.t21 48.0005
R90 GNDA.n2 GNDA.t1 48.0005
R91 GNDA.n2 GNDA.t17 48.0005
R92 GNDA.n4 GNDA.t10 48.0005
R93 GNDA.n4 GNDA.t19 48.0005
R94 GNDA.n3 GNDA.n1 0.688
R95 GNDA.n13 GNDA.n11 0.688
R96 GNDA.n9 GNDA.n7 0.313
R97 GNDA.n5 GNDA.n3 0.2755
R98 GNDA.n11 GNDA.n9 0.2755
R99 GNDA.n1 GNDA 0.238
R100 GNDA GNDA.n13 0.238
R101 GNDA.n7 GNDA 0.0755
R102 div2_3_2.CLK.n4 div2_3_2.CLK.t1 723.534
R103 div2_3_2.CLK.t2 div2_3_2.CLK.n5 723.534
R104 div2_3_2.CLK.n0 div2_3_2.CLK.t4 369.534
R105 div2_3_2.CLK.n3 div2_3_2.CLK.n2 366.856
R106 div2_3_2.CLK.n5 div2_3_2.CLK.t0 254.333
R107 div2_3_2.CLK.n3 div2_3_2.CLK.t7 190.123
R108 div2_3_2.CLK.n4 div2_3_2.CLK.n3 187.201
R109 div2_3_2.CLK.n1 div2_3_2.CLK.n0 176.733
R110 div2_3_2.CLK.n2 div2_3_2.CLK.n1 176.733
R111 div2_3_2.CLK.n0 div2_3_2.CLK.t5 112.468
R112 div2_3_2.CLK.n2 div2_3_2.CLK.t3 112.468
R113 div2_3_2.CLK.n1 div2_3_2.CLK.t6 112.468
R114 div2_3_2.CLK.n5 div2_3_2.CLK.n4 70.4005
R115 div2_3_1.CLK.n5 div2_3_1.CLK.t0 723.534
R116 div2_3_1.CLK.n4 div2_3_1.CLK.t2 723.534
R117 div2_3_1.CLK.n0 div2_3_1.CLK.t7 369.534
R118 div2_3_1.CLK.n3 div2_3_1.CLK.n2 366.856
R119 div2_3_1.CLK.t1 div2_3_1.CLK.n5 254.333
R120 div2_3_1.CLK.n3 div2_3_1.CLK.t6 190.123
R121 div2_3_1.CLK.n4 div2_3_1.CLK.n3 187.201
R122 div2_3_1.CLK.n1 div2_3_1.CLK.n0 176.733
R123 div2_3_1.CLK.n2 div2_3_1.CLK.n1 176.733
R124 div2_3_1.CLK.n0 div2_3_1.CLK.t3 112.468
R125 div2_3_1.CLK.n2 div2_3_1.CLK.t5 112.468
R126 div2_3_1.CLK.n1 div2_3_1.CLK.t4 112.468
R127 div2_3_1.CLK.n5 div2_3_1.CLK.n4 70.4005
R128 div2_3_2.A.n0 div2_3_2.A.t1 713.933
R129 div2_3_2.A.n0 div2_3_2.A.t2 314.233
R130 div2_3_2.A.t0 div2_3_2.A.n0 308.2
R131 div2_3_2.C.n2 div2_3_2.C.t3 721.4
R132 div2_3_2.C.n1 div2_3_2.C.t4 349.433
R133 div2_3_2.C.t2 div2_3_2.C.n2 276.733
R134 div2_3_2.C.n1 div2_3_2.C.n0 206.333
R135 div2_3_2.C.n0 div2_3_2.C.t1 48.0005
R136 div2_3_2.C.n0 div2_3_2.C.t0 48.0005
R137 div2_3_2.C.n2 div2_3_2.C.n1 48.0005
R138 VIN.t0 VIN.t2 401.668
R139 VIN.n0 VIN.t0 257.067
R140 VIN VIN.n0 216.9
R141 VIN.n0 VIN.t1 208.868
R142 VOUT.t3 VOUT.t2 819.4
R143 VOUT.n0 VOUT.t0 663.801
R144 VOUT.n0 VOUT.t3 489.168
R145 VOUT.n1 VOUT.t1 270.12
R146 VOUT.n2 VOUT 192.167
R147 VOUT.n1 VOUT.n0 67.2005
R148 VOUT.n2 VOUT.n1 25.6005
R149 VOUT VOUT.n2 4.8005
R150 div2_3_1.B.t0 div2_3_1.B.t1 96.0005
R151 div2_3_2.B.t0 div2_3_2.B.t1 96.0005
C0 VIN VDDA 0.125773f
C1 VDDA VOUT 0.488631f
C2 VIN GNDA 0.304628f
C3 VOUT GNDA 0.785902f
C4 VDDA GNDA 2.66524f
.ends

