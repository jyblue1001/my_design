magic
tech sky130A
magscale 1 2
timestamp 1746385583
<< error_p >>
rect 3991 142 4024 146
rect 8071 142 8104 146
rect 2590 92 2634 124
rect 2766 92 2814 124
rect 2946 92 2990 124
rect 3126 92 3170 124
rect 3306 92 3350 124
rect 3486 92 3530 124
rect 3666 92 3710 124
rect 3846 92 3890 124
rect 3972 114 4024 142
rect 4026 114 4074 124
rect 3972 92 4074 114
rect 2620 58 2634 92
rect 2800 58 2814 92
rect 3980 58 4004 92
rect 4024 58 4094 92
rect 4096 58 4124 142
rect 4206 92 4254 124
rect 4386 92 4434 124
rect 4566 92 4614 124
rect 4746 92 4794 124
rect 4926 92 4974 124
rect 5106 92 5154 124
rect 5286 92 5334 124
rect 5356 92 5384 142
rect 5456 124 5484 142
rect 5406 92 5434 116
rect 5456 92 5514 124
rect 4160 58 4184 92
rect 5330 58 5334 92
rect 5386 58 5454 92
rect 5456 58 5484 92
rect 5510 58 5514 92
rect 5646 92 5694 124
rect 5826 92 5874 124
rect 6006 92 6054 124
rect 6186 92 6234 124
rect 6366 92 6414 124
rect 6546 92 6594 124
rect 6726 92 6774 124
rect 5646 90 5654 92
rect 5826 90 5834 92
rect 6006 90 6014 92
rect 6186 90 6194 92
rect 6366 90 6374 92
rect 6546 90 6554 92
rect 6700 58 6704 92
rect 6726 90 6734 92
rect 6770 58 6794 92
rect 6816 58 6824 127
rect 6906 92 6954 124
rect 7086 92 7134 124
rect 7266 92 7314 124
rect 7446 92 7494 124
rect 7626 92 7674 124
rect 7806 92 7854 124
rect 7986 92 8034 124
rect 8056 92 8104 142
rect 8176 124 8204 142
rect 8106 114 8150 124
rect 8166 114 8214 124
rect 8106 92 8214 114
rect 6880 58 6884 92
rect 6906 90 6914 92
rect 7086 90 7104 92
rect 7266 90 7284 92
rect 7446 90 7464 92
rect 7626 90 7644 92
rect 7806 90 7824 92
rect 7986 90 8004 92
rect 7100 58 7104 90
rect 7280 58 7284 90
rect 7460 58 7464 90
rect 7640 58 7644 90
rect 7820 58 7824 90
rect 8000 58 8004 90
rect 8030 58 8034 92
rect 8104 90 8204 92
rect 8104 68 8194 90
rect 8104 58 8164 68
rect 8166 66 8194 68
rect 8176 58 8194 66
rect 8210 58 8214 92
rect 8346 92 8394 124
rect 8526 92 8574 124
rect 8706 92 8754 124
rect 8886 92 8934 124
rect 9066 92 9114 124
rect 9246 92 9294 124
rect 9366 92 9420 124
rect 9426 92 9474 124
rect 8346 90 8374 92
rect 8360 58 8374 90
rect 8390 58 8394 92
rect 8396 58 8424 92
rect 8526 90 8554 92
rect 8540 58 8554 90
rect 8570 58 8574 92
rect 8576 58 8604 92
rect 8706 90 8734 92
rect 8720 58 8734 90
rect 8750 58 8754 92
rect 8756 58 8784 92
rect 8886 90 8914 92
rect 8900 58 8914 90
rect 8930 58 8934 92
rect 8936 58 8964 92
rect 9066 90 9094 92
rect 9080 58 9094 90
rect 9110 58 9114 92
rect 9116 58 9144 92
rect 9246 90 9274 92
rect 9260 58 9274 90
rect 9290 58 9294 92
rect 9296 58 9324 92
rect 9366 90 9370 92
rect 9426 90 9454 92
rect 9400 58 9404 90
rect 9470 58 9494 92
rect 4040 34 4070 58
rect 5406 34 5434 58
rect 6746 34 6770 58
rect 8110 34 8140 58
rect 9464 34 9470 58
<< error_s >>
rect 2586 92 2590 124
<< nwell >>
rect 4300 3690 9310 5480
<< pwell >>
rect 1350 1187 2690 1340
rect 1350 153 1503 1187
rect 2537 153 2690 1187
rect 40 50 80 90
rect 1350 0 2690 153
rect 2710 1187 4050 1340
rect 2710 153 2863 1187
rect 3897 153 4050 1187
rect 2710 0 4050 153
rect 4070 1320 5400 1340
rect 5440 1320 6770 1340
rect 4070 1187 5410 1320
rect 4070 153 4223 1187
rect 5257 153 5410 1187
rect 4070 0 5410 153
rect 5430 1187 6770 1320
rect 5430 153 5583 1187
rect 6617 153 6770 1187
rect 5430 0 6770 153
rect 6790 1187 8130 1340
rect 6790 153 6943 1187
rect 7977 153 8130 1187
rect 6790 0 8130 153
rect 8150 1187 9490 1340
rect 8150 153 8303 1187
rect 9337 153 9490 1187
rect 8150 0 9490 153
<< nbase >>
rect 1503 153 2537 1187
rect 2863 153 3897 1187
rect 4223 153 5257 1187
rect 5583 153 6617 1187
rect 6943 153 7977 1187
rect 8303 153 9337 1187
<< nmos >>
rect 5220 3120 5340 3320
rect 5420 3120 5540 3320
rect 5620 3120 5740 3320
rect 5820 3120 5940 3320
rect 6020 3120 6140 3320
rect 6220 3120 6340 3320
rect 6580 3120 6700 3320
rect 6780 3120 6900 3320
rect 6980 3120 7100 3320
rect 7180 3120 7300 3320
rect 7380 3120 7500 3320
rect 7580 3120 7700 3320
rect 4740 1970 5540 2770
rect 5620 1970 6420 2770
rect 6500 1970 7300 2770
rect 7380 1970 8180 2770
rect 5440 1510 7440 1710
<< pmos >>
rect 4500 4640 4620 5440
rect 4700 4640 4820 5440
rect 4900 4640 5020 5440
rect 5100 4640 5220 5440
rect 5300 4640 5420 5440
rect 5500 4640 5620 5440
rect 5700 4640 5820 5440
rect 5900 4640 6020 5440
rect 6100 4640 6220 5440
rect 6300 4640 6420 5440
rect 6500 4640 6620 5440
rect 6700 4640 6820 5440
rect 6900 4640 7020 5440
rect 7100 4640 7220 5440
rect 7300 4640 7420 5440
rect 7500 4640 7620 5440
rect 7700 4640 7820 5440
rect 7900 4640 8020 5440
rect 8100 4640 8220 5440
rect 8300 4640 8420 5440
rect 4540 3730 4660 4130
rect 4740 3730 4860 4130
rect 4940 3730 5060 4130
rect 5140 3730 5260 4130
rect 5340 3730 5460 4130
rect 5540 3730 5660 4130
rect 5900 3730 6020 4130
rect 6100 3730 6220 4130
rect 6300 3730 6420 4130
rect 6500 3730 6620 4130
rect 6700 3730 6820 4130
rect 6900 3730 7020 4130
rect 7260 3730 7380 4130
rect 7460 3730 7580 4130
rect 7660 3730 7780 4130
rect 7860 3730 7980 4130
rect 8060 3730 8180 4130
rect 8260 3730 8380 4130
rect 8830 3730 8860 4130
rect 9080 3730 9110 4130
<< ndiff >>
rect 5140 3290 5220 3320
rect 5140 3250 5160 3290
rect 5200 3250 5220 3290
rect 5140 3190 5220 3250
rect 5140 3150 5160 3190
rect 5200 3150 5220 3190
rect 5140 3120 5220 3150
rect 5340 3290 5420 3320
rect 5340 3250 5360 3290
rect 5400 3250 5420 3290
rect 5340 3190 5420 3250
rect 5340 3150 5360 3190
rect 5400 3150 5420 3190
rect 5340 3120 5420 3150
rect 5540 3290 5620 3320
rect 5540 3250 5560 3290
rect 5600 3250 5620 3290
rect 5540 3190 5620 3250
rect 5540 3150 5560 3190
rect 5600 3150 5620 3190
rect 5540 3120 5620 3150
rect 5740 3290 5820 3320
rect 5740 3250 5760 3290
rect 5800 3250 5820 3290
rect 5740 3190 5820 3250
rect 5740 3150 5760 3190
rect 5800 3150 5820 3190
rect 5740 3120 5820 3150
rect 5940 3290 6020 3320
rect 5940 3250 5960 3290
rect 6000 3250 6020 3290
rect 5940 3190 6020 3250
rect 5940 3150 5960 3190
rect 6000 3150 6020 3190
rect 5940 3120 6020 3150
rect 6140 3290 6220 3320
rect 6140 3250 6160 3290
rect 6200 3250 6220 3290
rect 6140 3190 6220 3250
rect 6140 3150 6160 3190
rect 6200 3150 6220 3190
rect 6140 3120 6220 3150
rect 6340 3290 6420 3320
rect 6500 3290 6580 3320
rect 6340 3250 6360 3290
rect 6400 3250 6420 3290
rect 6500 3250 6520 3290
rect 6560 3250 6580 3290
rect 6340 3190 6420 3250
rect 6500 3190 6580 3250
rect 6340 3150 6360 3190
rect 6400 3150 6420 3190
rect 6500 3150 6520 3190
rect 6560 3150 6580 3190
rect 6340 3120 6420 3150
rect 6500 3120 6580 3150
rect 6700 3290 6780 3320
rect 6700 3250 6720 3290
rect 6760 3250 6780 3290
rect 6700 3190 6780 3250
rect 6700 3150 6720 3190
rect 6760 3150 6780 3190
rect 6700 3120 6780 3150
rect 6900 3290 6980 3320
rect 6900 3250 6920 3290
rect 6960 3250 6980 3290
rect 6900 3190 6980 3250
rect 6900 3150 6920 3190
rect 6960 3150 6980 3190
rect 6900 3120 6980 3150
rect 7100 3290 7180 3320
rect 7100 3250 7120 3290
rect 7160 3250 7180 3290
rect 7100 3190 7180 3250
rect 7100 3150 7120 3190
rect 7160 3150 7180 3190
rect 7100 3120 7180 3150
rect 7300 3290 7380 3320
rect 7300 3250 7320 3290
rect 7360 3250 7380 3290
rect 7300 3190 7380 3250
rect 7300 3150 7320 3190
rect 7360 3150 7380 3190
rect 7300 3120 7380 3150
rect 7500 3290 7580 3320
rect 7500 3250 7520 3290
rect 7560 3250 7580 3290
rect 7500 3190 7580 3250
rect 7500 3150 7520 3190
rect 7560 3150 7580 3190
rect 7500 3120 7580 3150
rect 7700 3290 7780 3320
rect 7700 3250 7720 3290
rect 7760 3250 7780 3290
rect 7700 3190 7780 3250
rect 7700 3150 7720 3190
rect 7760 3150 7780 3190
rect 7700 3120 7780 3150
rect 4660 2740 4740 2770
rect 4660 2700 4680 2740
rect 4720 2700 4740 2740
rect 4660 2640 4740 2700
rect 4660 2600 4680 2640
rect 4720 2600 4740 2640
rect 4660 2540 4740 2600
rect 4660 2500 4680 2540
rect 4720 2500 4740 2540
rect 4660 2440 4740 2500
rect 4660 2400 4680 2440
rect 4720 2400 4740 2440
rect 4660 2340 4740 2400
rect 4660 2300 4680 2340
rect 4720 2300 4740 2340
rect 4660 2240 4740 2300
rect 4660 2200 4680 2240
rect 4720 2200 4740 2240
rect 4660 2140 4740 2200
rect 4660 2100 4680 2140
rect 4720 2100 4740 2140
rect 4660 2040 4740 2100
rect 4660 2000 4680 2040
rect 4720 2000 4740 2040
rect 4660 1970 4740 2000
rect 5540 2740 5620 2770
rect 5540 2700 5560 2740
rect 5600 2700 5620 2740
rect 5540 2640 5620 2700
rect 5540 2600 5560 2640
rect 5600 2600 5620 2640
rect 5540 2540 5620 2600
rect 5540 2500 5560 2540
rect 5600 2500 5620 2540
rect 5540 2440 5620 2500
rect 5540 2400 5560 2440
rect 5600 2400 5620 2440
rect 5540 2340 5620 2400
rect 5540 2300 5560 2340
rect 5600 2300 5620 2340
rect 5540 2240 5620 2300
rect 5540 2200 5560 2240
rect 5600 2200 5620 2240
rect 5540 2140 5620 2200
rect 5540 2100 5560 2140
rect 5600 2100 5620 2140
rect 5540 2040 5620 2100
rect 5540 2000 5560 2040
rect 5600 2000 5620 2040
rect 5540 1970 5620 2000
rect 6420 2740 6500 2770
rect 6420 2700 6440 2740
rect 6480 2700 6500 2740
rect 6420 2640 6500 2700
rect 6420 2600 6440 2640
rect 6480 2600 6500 2640
rect 6420 2540 6500 2600
rect 6420 2500 6440 2540
rect 6480 2500 6500 2540
rect 6420 2440 6500 2500
rect 6420 2400 6440 2440
rect 6480 2400 6500 2440
rect 6420 2340 6500 2400
rect 6420 2300 6440 2340
rect 6480 2300 6500 2340
rect 6420 2240 6500 2300
rect 6420 2200 6440 2240
rect 6480 2200 6500 2240
rect 6420 2140 6500 2200
rect 6420 2100 6440 2140
rect 6480 2100 6500 2140
rect 6420 2040 6500 2100
rect 6420 2000 6440 2040
rect 6480 2000 6500 2040
rect 6420 1970 6500 2000
rect 7300 2740 7380 2770
rect 7300 2700 7320 2740
rect 7360 2700 7380 2740
rect 7300 2640 7380 2700
rect 7300 2600 7320 2640
rect 7360 2600 7380 2640
rect 7300 2540 7380 2600
rect 7300 2500 7320 2540
rect 7360 2500 7380 2540
rect 7300 2440 7380 2500
rect 7300 2400 7320 2440
rect 7360 2400 7380 2440
rect 7300 2340 7380 2400
rect 7300 2300 7320 2340
rect 7360 2300 7380 2340
rect 7300 2240 7380 2300
rect 7300 2200 7320 2240
rect 7360 2200 7380 2240
rect 7300 2140 7380 2200
rect 7300 2100 7320 2140
rect 7360 2100 7380 2140
rect 7300 2040 7380 2100
rect 7300 2000 7320 2040
rect 7360 2000 7380 2040
rect 7300 1970 7380 2000
rect 8180 2740 8260 2770
rect 8180 2700 8200 2740
rect 8240 2700 8260 2740
rect 8180 2640 8260 2700
rect 8180 2600 8200 2640
rect 8240 2600 8260 2640
rect 8180 2540 8260 2600
rect 8180 2500 8200 2540
rect 8240 2500 8260 2540
rect 8180 2440 8260 2500
rect 8180 2400 8200 2440
rect 8240 2400 8260 2440
rect 8180 2340 8260 2400
rect 8180 2300 8200 2340
rect 8240 2300 8260 2340
rect 8180 2240 8260 2300
rect 8180 2200 8200 2240
rect 8240 2200 8260 2240
rect 8180 2140 8260 2200
rect 8180 2100 8200 2140
rect 8240 2100 8260 2140
rect 8180 2040 8260 2100
rect 8180 2000 8200 2040
rect 8240 2000 8260 2040
rect 8180 1970 8260 2000
rect 5360 1680 5440 1710
rect 5360 1640 5380 1680
rect 5420 1640 5440 1680
rect 5360 1580 5440 1640
rect 5360 1540 5380 1580
rect 5420 1540 5440 1580
rect 5360 1510 5440 1540
rect 7440 1680 7520 1710
rect 7440 1640 7460 1680
rect 7500 1640 7520 1680
rect 7440 1580 7520 1640
rect 7440 1540 7460 1580
rect 7500 1540 7520 1580
rect 7440 1510 7520 1540
<< pdiff >>
rect 4420 5410 4500 5440
rect 4420 5370 4440 5410
rect 4480 5370 4500 5410
rect 4420 5310 4500 5370
rect 4420 5270 4440 5310
rect 4480 5270 4500 5310
rect 4420 5210 4500 5270
rect 4420 5170 4440 5210
rect 4480 5170 4500 5210
rect 4420 5110 4500 5170
rect 4420 5070 4440 5110
rect 4480 5070 4500 5110
rect 4420 5010 4500 5070
rect 4420 4970 4440 5010
rect 4480 4970 4500 5010
rect 4420 4910 4500 4970
rect 4420 4870 4440 4910
rect 4480 4870 4500 4910
rect 4420 4810 4500 4870
rect 4420 4770 4440 4810
rect 4480 4770 4500 4810
rect 4420 4710 4500 4770
rect 4420 4670 4440 4710
rect 4480 4670 4500 4710
rect 4420 4640 4500 4670
rect 4620 5410 4700 5440
rect 4620 5370 4640 5410
rect 4680 5370 4700 5410
rect 4620 5310 4700 5370
rect 4620 5270 4640 5310
rect 4680 5270 4700 5310
rect 4620 5210 4700 5270
rect 4620 5170 4640 5210
rect 4680 5170 4700 5210
rect 4620 5110 4700 5170
rect 4620 5070 4640 5110
rect 4680 5070 4700 5110
rect 4620 5010 4700 5070
rect 4620 4970 4640 5010
rect 4680 4970 4700 5010
rect 4620 4910 4700 4970
rect 4620 4870 4640 4910
rect 4680 4870 4700 4910
rect 4620 4810 4700 4870
rect 4620 4770 4640 4810
rect 4680 4770 4700 4810
rect 4620 4710 4700 4770
rect 4620 4670 4640 4710
rect 4680 4670 4700 4710
rect 4620 4640 4700 4670
rect 4820 5410 4900 5440
rect 4820 5370 4840 5410
rect 4880 5370 4900 5410
rect 4820 5310 4900 5370
rect 4820 5270 4840 5310
rect 4880 5270 4900 5310
rect 4820 5210 4900 5270
rect 4820 5170 4840 5210
rect 4880 5170 4900 5210
rect 4820 5110 4900 5170
rect 4820 5070 4840 5110
rect 4880 5070 4900 5110
rect 4820 5010 4900 5070
rect 4820 4970 4840 5010
rect 4880 4970 4900 5010
rect 4820 4910 4900 4970
rect 4820 4870 4840 4910
rect 4880 4870 4900 4910
rect 4820 4810 4900 4870
rect 4820 4770 4840 4810
rect 4880 4770 4900 4810
rect 4820 4710 4900 4770
rect 4820 4670 4840 4710
rect 4880 4670 4900 4710
rect 4820 4640 4900 4670
rect 5020 5410 5100 5440
rect 5020 5370 5040 5410
rect 5080 5370 5100 5410
rect 5020 5310 5100 5370
rect 5020 5270 5040 5310
rect 5080 5270 5100 5310
rect 5020 5210 5100 5270
rect 5020 5170 5040 5210
rect 5080 5170 5100 5210
rect 5020 5110 5100 5170
rect 5020 5070 5040 5110
rect 5080 5070 5100 5110
rect 5020 5010 5100 5070
rect 5020 4970 5040 5010
rect 5080 4970 5100 5010
rect 5020 4910 5100 4970
rect 5020 4870 5040 4910
rect 5080 4870 5100 4910
rect 5020 4810 5100 4870
rect 5020 4770 5040 4810
rect 5080 4770 5100 4810
rect 5020 4710 5100 4770
rect 5020 4670 5040 4710
rect 5080 4670 5100 4710
rect 5020 4640 5100 4670
rect 5220 5410 5300 5440
rect 5220 5370 5240 5410
rect 5280 5370 5300 5410
rect 5220 5310 5300 5370
rect 5220 5270 5240 5310
rect 5280 5270 5300 5310
rect 5220 5210 5300 5270
rect 5220 5170 5240 5210
rect 5280 5170 5300 5210
rect 5220 5110 5300 5170
rect 5220 5070 5240 5110
rect 5280 5070 5300 5110
rect 5220 5010 5300 5070
rect 5220 4970 5240 5010
rect 5280 4970 5300 5010
rect 5220 4910 5300 4970
rect 5220 4870 5240 4910
rect 5280 4870 5300 4910
rect 5220 4810 5300 4870
rect 5220 4770 5240 4810
rect 5280 4770 5300 4810
rect 5220 4710 5300 4770
rect 5220 4670 5240 4710
rect 5280 4670 5300 4710
rect 5220 4640 5300 4670
rect 5420 5410 5500 5440
rect 5420 5370 5440 5410
rect 5480 5370 5500 5410
rect 5420 5310 5500 5370
rect 5420 5270 5440 5310
rect 5480 5270 5500 5310
rect 5420 5210 5500 5270
rect 5420 5170 5440 5210
rect 5480 5170 5500 5210
rect 5420 5110 5500 5170
rect 5420 5070 5440 5110
rect 5480 5070 5500 5110
rect 5420 5010 5500 5070
rect 5420 4970 5440 5010
rect 5480 4970 5500 5010
rect 5420 4910 5500 4970
rect 5420 4870 5440 4910
rect 5480 4870 5500 4910
rect 5420 4810 5500 4870
rect 5420 4770 5440 4810
rect 5480 4770 5500 4810
rect 5420 4710 5500 4770
rect 5420 4670 5440 4710
rect 5480 4670 5500 4710
rect 5420 4640 5500 4670
rect 5620 5410 5700 5440
rect 5620 5370 5640 5410
rect 5680 5370 5700 5410
rect 5620 5310 5700 5370
rect 5620 5270 5640 5310
rect 5680 5270 5700 5310
rect 5620 5210 5700 5270
rect 5620 5170 5640 5210
rect 5680 5170 5700 5210
rect 5620 5110 5700 5170
rect 5620 5070 5640 5110
rect 5680 5070 5700 5110
rect 5620 5010 5700 5070
rect 5620 4970 5640 5010
rect 5680 4970 5700 5010
rect 5620 4910 5700 4970
rect 5620 4870 5640 4910
rect 5680 4870 5700 4910
rect 5620 4810 5700 4870
rect 5620 4770 5640 4810
rect 5680 4770 5700 4810
rect 5620 4710 5700 4770
rect 5620 4670 5640 4710
rect 5680 4670 5700 4710
rect 5620 4640 5700 4670
rect 5820 5410 5900 5440
rect 5820 5370 5840 5410
rect 5880 5370 5900 5410
rect 5820 5310 5900 5370
rect 5820 5270 5840 5310
rect 5880 5270 5900 5310
rect 5820 5210 5900 5270
rect 5820 5170 5840 5210
rect 5880 5170 5900 5210
rect 5820 5110 5900 5170
rect 5820 5070 5840 5110
rect 5880 5070 5900 5110
rect 5820 5010 5900 5070
rect 5820 4970 5840 5010
rect 5880 4970 5900 5010
rect 5820 4910 5900 4970
rect 5820 4870 5840 4910
rect 5880 4870 5900 4910
rect 5820 4810 5900 4870
rect 5820 4770 5840 4810
rect 5880 4770 5900 4810
rect 5820 4710 5900 4770
rect 5820 4670 5840 4710
rect 5880 4670 5900 4710
rect 5820 4640 5900 4670
rect 6020 5410 6100 5440
rect 6020 5370 6040 5410
rect 6080 5370 6100 5410
rect 6020 5310 6100 5370
rect 6020 5270 6040 5310
rect 6080 5270 6100 5310
rect 6020 5210 6100 5270
rect 6020 5170 6040 5210
rect 6080 5170 6100 5210
rect 6020 5110 6100 5170
rect 6020 5070 6040 5110
rect 6080 5070 6100 5110
rect 6020 5010 6100 5070
rect 6020 4970 6040 5010
rect 6080 4970 6100 5010
rect 6020 4910 6100 4970
rect 6020 4870 6040 4910
rect 6080 4870 6100 4910
rect 6020 4810 6100 4870
rect 6020 4770 6040 4810
rect 6080 4770 6100 4810
rect 6020 4710 6100 4770
rect 6020 4670 6040 4710
rect 6080 4670 6100 4710
rect 6020 4640 6100 4670
rect 6220 5410 6300 5440
rect 6220 5370 6240 5410
rect 6280 5370 6300 5410
rect 6220 5310 6300 5370
rect 6220 5270 6240 5310
rect 6280 5270 6300 5310
rect 6220 5210 6300 5270
rect 6220 5170 6240 5210
rect 6280 5170 6300 5210
rect 6220 5110 6300 5170
rect 6220 5070 6240 5110
rect 6280 5070 6300 5110
rect 6220 5010 6300 5070
rect 6220 4970 6240 5010
rect 6280 4970 6300 5010
rect 6220 4910 6300 4970
rect 6220 4870 6240 4910
rect 6280 4870 6300 4910
rect 6220 4810 6300 4870
rect 6220 4770 6240 4810
rect 6280 4770 6300 4810
rect 6220 4710 6300 4770
rect 6220 4670 6240 4710
rect 6280 4670 6300 4710
rect 6220 4640 6300 4670
rect 6420 5410 6500 5440
rect 6420 5370 6440 5410
rect 6480 5370 6500 5410
rect 6420 5310 6500 5370
rect 6420 5270 6440 5310
rect 6480 5270 6500 5310
rect 6420 5210 6500 5270
rect 6420 5170 6440 5210
rect 6480 5170 6500 5210
rect 6420 5110 6500 5170
rect 6420 5070 6440 5110
rect 6480 5070 6500 5110
rect 6420 5010 6500 5070
rect 6420 4970 6440 5010
rect 6480 4970 6500 5010
rect 6420 4910 6500 4970
rect 6420 4870 6440 4910
rect 6480 4870 6500 4910
rect 6420 4810 6500 4870
rect 6420 4770 6440 4810
rect 6480 4770 6500 4810
rect 6420 4710 6500 4770
rect 6420 4670 6440 4710
rect 6480 4670 6500 4710
rect 6420 4640 6500 4670
rect 6620 5410 6700 5440
rect 6620 5370 6640 5410
rect 6680 5370 6700 5410
rect 6620 5310 6700 5370
rect 6620 5270 6640 5310
rect 6680 5270 6700 5310
rect 6620 5210 6700 5270
rect 6620 5170 6640 5210
rect 6680 5170 6700 5210
rect 6620 5110 6700 5170
rect 6620 5070 6640 5110
rect 6680 5070 6700 5110
rect 6620 5010 6700 5070
rect 6620 4970 6640 5010
rect 6680 4970 6700 5010
rect 6620 4910 6700 4970
rect 6620 4870 6640 4910
rect 6680 4870 6700 4910
rect 6620 4810 6700 4870
rect 6620 4770 6640 4810
rect 6680 4770 6700 4810
rect 6620 4710 6700 4770
rect 6620 4670 6640 4710
rect 6680 4670 6700 4710
rect 6620 4640 6700 4670
rect 6820 5410 6900 5440
rect 6820 5370 6840 5410
rect 6880 5370 6900 5410
rect 6820 5310 6900 5370
rect 6820 5270 6840 5310
rect 6880 5270 6900 5310
rect 6820 5210 6900 5270
rect 6820 5170 6840 5210
rect 6880 5170 6900 5210
rect 6820 5110 6900 5170
rect 6820 5070 6840 5110
rect 6880 5070 6900 5110
rect 6820 5010 6900 5070
rect 6820 4970 6840 5010
rect 6880 4970 6900 5010
rect 6820 4910 6900 4970
rect 6820 4870 6840 4910
rect 6880 4870 6900 4910
rect 6820 4810 6900 4870
rect 6820 4770 6840 4810
rect 6880 4770 6900 4810
rect 6820 4710 6900 4770
rect 6820 4670 6840 4710
rect 6880 4670 6900 4710
rect 6820 4640 6900 4670
rect 7020 5410 7100 5440
rect 7020 5370 7040 5410
rect 7080 5370 7100 5410
rect 7020 5310 7100 5370
rect 7020 5270 7040 5310
rect 7080 5270 7100 5310
rect 7020 5210 7100 5270
rect 7020 5170 7040 5210
rect 7080 5170 7100 5210
rect 7020 5110 7100 5170
rect 7020 5070 7040 5110
rect 7080 5070 7100 5110
rect 7020 5010 7100 5070
rect 7020 4970 7040 5010
rect 7080 4970 7100 5010
rect 7020 4910 7100 4970
rect 7020 4870 7040 4910
rect 7080 4870 7100 4910
rect 7020 4810 7100 4870
rect 7020 4770 7040 4810
rect 7080 4770 7100 4810
rect 7020 4710 7100 4770
rect 7020 4670 7040 4710
rect 7080 4670 7100 4710
rect 7020 4640 7100 4670
rect 7220 5410 7300 5440
rect 7220 5370 7240 5410
rect 7280 5370 7300 5410
rect 7220 5310 7300 5370
rect 7220 5270 7240 5310
rect 7280 5270 7300 5310
rect 7220 5210 7300 5270
rect 7220 5170 7240 5210
rect 7280 5170 7300 5210
rect 7220 5110 7300 5170
rect 7220 5070 7240 5110
rect 7280 5070 7300 5110
rect 7220 5010 7300 5070
rect 7220 4970 7240 5010
rect 7280 4970 7300 5010
rect 7220 4910 7300 4970
rect 7220 4870 7240 4910
rect 7280 4870 7300 4910
rect 7220 4810 7300 4870
rect 7220 4770 7240 4810
rect 7280 4770 7300 4810
rect 7220 4710 7300 4770
rect 7220 4670 7240 4710
rect 7280 4670 7300 4710
rect 7220 4640 7300 4670
rect 7420 5410 7500 5440
rect 7420 5370 7440 5410
rect 7480 5370 7500 5410
rect 7420 5310 7500 5370
rect 7420 5270 7440 5310
rect 7480 5270 7500 5310
rect 7420 5210 7500 5270
rect 7420 5170 7440 5210
rect 7480 5170 7500 5210
rect 7420 5110 7500 5170
rect 7420 5070 7440 5110
rect 7480 5070 7500 5110
rect 7420 5010 7500 5070
rect 7420 4970 7440 5010
rect 7480 4970 7500 5010
rect 7420 4910 7500 4970
rect 7420 4870 7440 4910
rect 7480 4870 7500 4910
rect 7420 4810 7500 4870
rect 7420 4770 7440 4810
rect 7480 4770 7500 4810
rect 7420 4710 7500 4770
rect 7420 4670 7440 4710
rect 7480 4670 7500 4710
rect 7420 4640 7500 4670
rect 7620 5410 7700 5440
rect 7620 5370 7640 5410
rect 7680 5370 7700 5410
rect 7620 5310 7700 5370
rect 7620 5270 7640 5310
rect 7680 5270 7700 5310
rect 7620 5210 7700 5270
rect 7620 5170 7640 5210
rect 7680 5170 7700 5210
rect 7620 5110 7700 5170
rect 7620 5070 7640 5110
rect 7680 5070 7700 5110
rect 7620 5010 7700 5070
rect 7620 4970 7640 5010
rect 7680 4970 7700 5010
rect 7620 4910 7700 4970
rect 7620 4870 7640 4910
rect 7680 4870 7700 4910
rect 7620 4810 7700 4870
rect 7620 4770 7640 4810
rect 7680 4770 7700 4810
rect 7620 4710 7700 4770
rect 7620 4670 7640 4710
rect 7680 4670 7700 4710
rect 7620 4640 7700 4670
rect 7820 5410 7900 5440
rect 7820 5370 7840 5410
rect 7880 5370 7900 5410
rect 7820 5310 7900 5370
rect 7820 5270 7840 5310
rect 7880 5270 7900 5310
rect 7820 5210 7900 5270
rect 7820 5170 7840 5210
rect 7880 5170 7900 5210
rect 7820 5110 7900 5170
rect 7820 5070 7840 5110
rect 7880 5070 7900 5110
rect 7820 5010 7900 5070
rect 7820 4970 7840 5010
rect 7880 4970 7900 5010
rect 7820 4910 7900 4970
rect 7820 4870 7840 4910
rect 7880 4870 7900 4910
rect 7820 4810 7900 4870
rect 7820 4770 7840 4810
rect 7880 4770 7900 4810
rect 7820 4710 7900 4770
rect 7820 4670 7840 4710
rect 7880 4670 7900 4710
rect 7820 4640 7900 4670
rect 8020 5410 8100 5440
rect 8020 5370 8040 5410
rect 8080 5370 8100 5410
rect 8020 5310 8100 5370
rect 8020 5270 8040 5310
rect 8080 5270 8100 5310
rect 8020 5210 8100 5270
rect 8020 5170 8040 5210
rect 8080 5170 8100 5210
rect 8020 5110 8100 5170
rect 8020 5070 8040 5110
rect 8080 5070 8100 5110
rect 8020 5010 8100 5070
rect 8020 4970 8040 5010
rect 8080 4970 8100 5010
rect 8020 4910 8100 4970
rect 8020 4870 8040 4910
rect 8080 4870 8100 4910
rect 8020 4810 8100 4870
rect 8020 4770 8040 4810
rect 8080 4770 8100 4810
rect 8020 4710 8100 4770
rect 8020 4670 8040 4710
rect 8080 4670 8100 4710
rect 8020 4640 8100 4670
rect 8220 5410 8300 5440
rect 8220 5370 8240 5410
rect 8280 5370 8300 5410
rect 8220 5310 8300 5370
rect 8220 5270 8240 5310
rect 8280 5270 8300 5310
rect 8220 5210 8300 5270
rect 8220 5170 8240 5210
rect 8280 5170 8300 5210
rect 8220 5110 8300 5170
rect 8220 5070 8240 5110
rect 8280 5070 8300 5110
rect 8220 5010 8300 5070
rect 8220 4970 8240 5010
rect 8280 4970 8300 5010
rect 8220 4910 8300 4970
rect 8220 4870 8240 4910
rect 8280 4870 8300 4910
rect 8220 4810 8300 4870
rect 8220 4770 8240 4810
rect 8280 4770 8300 4810
rect 8220 4710 8300 4770
rect 8220 4670 8240 4710
rect 8280 4670 8300 4710
rect 8220 4640 8300 4670
rect 8420 5410 8500 5440
rect 8420 5370 8440 5410
rect 8480 5370 8500 5410
rect 8420 5310 8500 5370
rect 8420 5270 8440 5310
rect 8480 5270 8500 5310
rect 8420 5210 8500 5270
rect 8420 5170 8440 5210
rect 8480 5170 8500 5210
rect 8420 5110 8500 5170
rect 8420 5070 8440 5110
rect 8480 5070 8500 5110
rect 8420 5010 8500 5070
rect 8420 4970 8440 5010
rect 8480 4970 8500 5010
rect 8420 4910 8500 4970
rect 8420 4870 8440 4910
rect 8480 4870 8500 4910
rect 8420 4810 8500 4870
rect 8420 4770 8440 4810
rect 8480 4770 8500 4810
rect 8420 4710 8500 4770
rect 8420 4670 8440 4710
rect 8480 4670 8500 4710
rect 8420 4640 8500 4670
rect 4460 4100 4540 4130
rect 4460 4060 4480 4100
rect 4520 4060 4540 4100
rect 4460 4000 4540 4060
rect 4460 3960 4480 4000
rect 4520 3960 4540 4000
rect 4460 3900 4540 3960
rect 4460 3860 4480 3900
rect 4520 3860 4540 3900
rect 4460 3800 4540 3860
rect 4460 3760 4480 3800
rect 4520 3760 4540 3800
rect 4460 3730 4540 3760
rect 4660 4100 4740 4130
rect 4660 4060 4680 4100
rect 4720 4060 4740 4100
rect 4660 4000 4740 4060
rect 4660 3960 4680 4000
rect 4720 3960 4740 4000
rect 4660 3900 4740 3960
rect 4660 3860 4680 3900
rect 4720 3860 4740 3900
rect 4660 3800 4740 3860
rect 4660 3760 4680 3800
rect 4720 3760 4740 3800
rect 4660 3730 4740 3760
rect 4860 4100 4940 4130
rect 4860 4060 4880 4100
rect 4920 4060 4940 4100
rect 4860 4000 4940 4060
rect 4860 3960 4880 4000
rect 4920 3960 4940 4000
rect 4860 3900 4940 3960
rect 4860 3860 4880 3900
rect 4920 3860 4940 3900
rect 4860 3800 4940 3860
rect 4860 3760 4880 3800
rect 4920 3760 4940 3800
rect 4860 3730 4940 3760
rect 5060 4100 5140 4130
rect 5060 4060 5080 4100
rect 5120 4060 5140 4100
rect 5060 4000 5140 4060
rect 5060 3960 5080 4000
rect 5120 3960 5140 4000
rect 5060 3900 5140 3960
rect 5060 3860 5080 3900
rect 5120 3860 5140 3900
rect 5060 3800 5140 3860
rect 5060 3760 5080 3800
rect 5120 3760 5140 3800
rect 5060 3730 5140 3760
rect 5260 4100 5340 4130
rect 5260 4060 5280 4100
rect 5320 4060 5340 4100
rect 5260 4000 5340 4060
rect 5260 3960 5280 4000
rect 5320 3960 5340 4000
rect 5260 3900 5340 3960
rect 5260 3860 5280 3900
rect 5320 3860 5340 3900
rect 5260 3800 5340 3860
rect 5260 3760 5280 3800
rect 5320 3760 5340 3800
rect 5260 3730 5340 3760
rect 5460 4100 5540 4130
rect 5460 4060 5480 4100
rect 5520 4060 5540 4100
rect 5460 4000 5540 4060
rect 5460 3960 5480 4000
rect 5520 3960 5540 4000
rect 5460 3900 5540 3960
rect 5460 3860 5480 3900
rect 5520 3860 5540 3900
rect 5460 3800 5540 3860
rect 5460 3760 5480 3800
rect 5520 3760 5540 3800
rect 5460 3730 5540 3760
rect 5660 4100 5740 4130
rect 5820 4100 5900 4130
rect 5660 4060 5680 4100
rect 5720 4060 5740 4100
rect 5820 4060 5840 4100
rect 5880 4060 5900 4100
rect 5660 4000 5740 4060
rect 5820 4000 5900 4060
rect 5660 3960 5680 4000
rect 5720 3960 5740 4000
rect 5820 3960 5840 4000
rect 5880 3960 5900 4000
rect 5660 3900 5740 3960
rect 5820 3900 5900 3960
rect 5660 3860 5680 3900
rect 5720 3860 5740 3900
rect 5820 3860 5840 3900
rect 5880 3860 5900 3900
rect 5660 3800 5740 3860
rect 5820 3800 5900 3860
rect 5660 3760 5680 3800
rect 5720 3760 5740 3800
rect 5820 3760 5840 3800
rect 5880 3760 5900 3800
rect 5660 3730 5740 3760
rect 5820 3730 5900 3760
rect 6020 4100 6100 4130
rect 6020 4060 6040 4100
rect 6080 4060 6100 4100
rect 6020 4000 6100 4060
rect 6020 3960 6040 4000
rect 6080 3960 6100 4000
rect 6020 3900 6100 3960
rect 6020 3860 6040 3900
rect 6080 3860 6100 3900
rect 6020 3800 6100 3860
rect 6020 3760 6040 3800
rect 6080 3760 6100 3800
rect 6020 3730 6100 3760
rect 6220 4100 6300 4130
rect 6220 4060 6240 4100
rect 6280 4060 6300 4100
rect 6220 4000 6300 4060
rect 6220 3960 6240 4000
rect 6280 3960 6300 4000
rect 6220 3900 6300 3960
rect 6220 3860 6240 3900
rect 6280 3860 6300 3900
rect 6220 3800 6300 3860
rect 6220 3760 6240 3800
rect 6280 3760 6300 3800
rect 6220 3730 6300 3760
rect 6420 4100 6500 4130
rect 6420 4060 6440 4100
rect 6480 4060 6500 4100
rect 6420 4000 6500 4060
rect 6420 3960 6440 4000
rect 6480 3960 6500 4000
rect 6420 3900 6500 3960
rect 6420 3860 6440 3900
rect 6480 3860 6500 3900
rect 6420 3800 6500 3860
rect 6420 3760 6440 3800
rect 6480 3760 6500 3800
rect 6420 3730 6500 3760
rect 6620 4100 6700 4130
rect 6620 4060 6640 4100
rect 6680 4060 6700 4100
rect 6620 4000 6700 4060
rect 6620 3960 6640 4000
rect 6680 3960 6700 4000
rect 6620 3900 6700 3960
rect 6620 3860 6640 3900
rect 6680 3860 6700 3900
rect 6620 3800 6700 3860
rect 6620 3760 6640 3800
rect 6680 3760 6700 3800
rect 6620 3730 6700 3760
rect 6820 4100 6900 4130
rect 6820 4060 6840 4100
rect 6880 4060 6900 4100
rect 6820 4000 6900 4060
rect 6820 3960 6840 4000
rect 6880 3960 6900 4000
rect 6820 3900 6900 3960
rect 6820 3860 6840 3900
rect 6880 3860 6900 3900
rect 6820 3800 6900 3860
rect 6820 3760 6840 3800
rect 6880 3760 6900 3800
rect 6820 3730 6900 3760
rect 7020 4100 7100 4130
rect 7180 4100 7260 4130
rect 7020 4060 7040 4100
rect 7080 4060 7100 4100
rect 7180 4060 7200 4100
rect 7240 4060 7260 4100
rect 7020 4000 7100 4060
rect 7180 4000 7260 4060
rect 7020 3960 7040 4000
rect 7080 3960 7100 4000
rect 7180 3960 7200 4000
rect 7240 3960 7260 4000
rect 7020 3900 7100 3960
rect 7180 3900 7260 3960
rect 7020 3860 7040 3900
rect 7080 3860 7100 3900
rect 7180 3860 7200 3900
rect 7240 3860 7260 3900
rect 7020 3800 7100 3860
rect 7180 3800 7260 3860
rect 7020 3760 7040 3800
rect 7080 3760 7100 3800
rect 7180 3760 7200 3800
rect 7240 3760 7260 3800
rect 7020 3730 7100 3760
rect 7180 3730 7260 3760
rect 7380 4100 7460 4130
rect 7380 4060 7400 4100
rect 7440 4060 7460 4100
rect 7380 4000 7460 4060
rect 7380 3960 7400 4000
rect 7440 3960 7460 4000
rect 7380 3900 7460 3960
rect 7380 3860 7400 3900
rect 7440 3860 7460 3900
rect 7380 3800 7460 3860
rect 7380 3760 7400 3800
rect 7440 3760 7460 3800
rect 7380 3730 7460 3760
rect 7580 4100 7660 4130
rect 7580 4060 7600 4100
rect 7640 4060 7660 4100
rect 7580 4000 7660 4060
rect 7580 3960 7600 4000
rect 7640 3960 7660 4000
rect 7580 3900 7660 3960
rect 7580 3860 7600 3900
rect 7640 3860 7660 3900
rect 7580 3800 7660 3860
rect 7580 3760 7600 3800
rect 7640 3760 7660 3800
rect 7580 3730 7660 3760
rect 7780 4100 7860 4130
rect 7780 4060 7800 4100
rect 7840 4060 7860 4100
rect 7780 4000 7860 4060
rect 7780 3960 7800 4000
rect 7840 3960 7860 4000
rect 7780 3900 7860 3960
rect 7780 3860 7800 3900
rect 7840 3860 7860 3900
rect 7780 3800 7860 3860
rect 7780 3760 7800 3800
rect 7840 3760 7860 3800
rect 7780 3730 7860 3760
rect 7980 4100 8060 4130
rect 7980 4060 8000 4100
rect 8040 4060 8060 4100
rect 7980 4000 8060 4060
rect 7980 3960 8000 4000
rect 8040 3960 8060 4000
rect 7980 3900 8060 3960
rect 7980 3860 8000 3900
rect 8040 3860 8060 3900
rect 7980 3800 8060 3860
rect 7980 3760 8000 3800
rect 8040 3760 8060 3800
rect 7980 3730 8060 3760
rect 8180 4100 8260 4130
rect 8180 4060 8200 4100
rect 8240 4060 8260 4100
rect 8180 4000 8260 4060
rect 8180 3960 8200 4000
rect 8240 3960 8260 4000
rect 8180 3900 8260 3960
rect 8180 3860 8200 3900
rect 8240 3860 8260 3900
rect 8180 3800 8260 3860
rect 8180 3760 8200 3800
rect 8240 3760 8260 3800
rect 8180 3730 8260 3760
rect 8380 4100 8460 4130
rect 8380 4060 8400 4100
rect 8440 4060 8460 4100
rect 8380 4000 8460 4060
rect 8380 3960 8400 4000
rect 8440 3960 8460 4000
rect 8380 3900 8460 3960
rect 8380 3860 8400 3900
rect 8440 3860 8460 3900
rect 8380 3800 8460 3860
rect 8380 3760 8400 3800
rect 8440 3760 8460 3800
rect 8380 3730 8460 3760
rect 8750 4100 8830 4130
rect 8750 4060 8770 4100
rect 8810 4060 8830 4100
rect 8750 4000 8830 4060
rect 8750 3960 8770 4000
rect 8810 3960 8830 4000
rect 8750 3900 8830 3960
rect 8750 3860 8770 3900
rect 8810 3860 8830 3900
rect 8750 3800 8830 3860
rect 8750 3760 8770 3800
rect 8810 3760 8830 3800
rect 8750 3730 8830 3760
rect 8860 4100 8940 4130
rect 8860 4060 8880 4100
rect 8920 4060 8940 4100
rect 8860 4000 8940 4060
rect 8860 3960 8880 4000
rect 8920 3960 8940 4000
rect 8860 3900 8940 3960
rect 8860 3860 8880 3900
rect 8920 3860 8940 3900
rect 8860 3800 8940 3860
rect 8860 3760 8880 3800
rect 8920 3760 8940 3800
rect 8860 3730 8940 3760
rect 9000 4100 9080 4130
rect 9000 4060 9020 4100
rect 9060 4060 9080 4100
rect 9000 4000 9080 4060
rect 9000 3960 9020 4000
rect 9060 3960 9080 4000
rect 9000 3900 9080 3960
rect 9000 3860 9020 3900
rect 9060 3860 9080 3900
rect 9000 3800 9080 3860
rect 9000 3760 9020 3800
rect 9060 3760 9080 3800
rect 9000 3730 9080 3760
rect 9110 4100 9190 4130
rect 9110 4060 9130 4100
rect 9170 4060 9190 4100
rect 9110 4000 9190 4060
rect 9110 3960 9130 4000
rect 9170 3960 9190 4000
rect 9110 3900 9190 3960
rect 9110 3860 9130 3900
rect 9170 3860 9190 3900
rect 9110 3800 9190 3860
rect 9110 3760 9130 3800
rect 9170 3760 9190 3800
rect 9110 3730 9190 3760
rect 1680 958 2360 1010
rect 1680 924 1734 958
rect 1768 924 1824 958
rect 1858 924 1914 958
rect 1948 924 2004 958
rect 2038 924 2094 958
rect 2128 924 2184 958
rect 2218 924 2274 958
rect 2308 924 2360 958
rect 1680 868 2360 924
rect 1680 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2360 868
rect 1680 778 2360 834
rect 1680 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2360 778
rect 1680 688 2360 744
rect 1680 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2360 688
rect 1680 598 2360 654
rect 1680 564 1734 598
rect 1768 564 1824 598
rect 1858 564 1914 598
rect 1948 564 2004 598
rect 2038 564 2094 598
rect 2128 564 2184 598
rect 2218 564 2274 598
rect 2308 564 2360 598
rect 1680 508 2360 564
rect 1680 474 1734 508
rect 1768 474 1824 508
rect 1858 474 1914 508
rect 1948 474 2004 508
rect 2038 474 2094 508
rect 2128 474 2184 508
rect 2218 474 2274 508
rect 2308 474 2360 508
rect 1680 418 2360 474
rect 1680 384 1734 418
rect 1768 384 1824 418
rect 1858 384 1914 418
rect 1948 384 2004 418
rect 2038 384 2094 418
rect 2128 384 2184 418
rect 2218 384 2274 418
rect 2308 384 2360 418
rect 1680 330 2360 384
rect 3040 958 3720 1010
rect 3040 924 3094 958
rect 3128 924 3184 958
rect 3218 924 3274 958
rect 3308 924 3364 958
rect 3398 924 3454 958
rect 3488 924 3544 958
rect 3578 924 3634 958
rect 3668 924 3720 958
rect 3040 868 3720 924
rect 3040 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3720 868
rect 3040 778 3720 834
rect 3040 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3720 778
rect 3040 688 3720 744
rect 3040 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3720 688
rect 3040 598 3720 654
rect 3040 564 3094 598
rect 3128 564 3184 598
rect 3218 564 3274 598
rect 3308 564 3364 598
rect 3398 564 3454 598
rect 3488 564 3544 598
rect 3578 564 3634 598
rect 3668 564 3720 598
rect 3040 508 3720 564
rect 3040 474 3094 508
rect 3128 474 3184 508
rect 3218 474 3274 508
rect 3308 474 3364 508
rect 3398 474 3454 508
rect 3488 474 3544 508
rect 3578 474 3634 508
rect 3668 474 3720 508
rect 3040 418 3720 474
rect 3040 384 3094 418
rect 3128 384 3184 418
rect 3218 384 3274 418
rect 3308 384 3364 418
rect 3398 384 3454 418
rect 3488 384 3544 418
rect 3578 384 3634 418
rect 3668 384 3720 418
rect 3040 330 3720 384
rect 4400 958 5080 1010
rect 4400 924 4454 958
rect 4488 924 4544 958
rect 4578 924 4634 958
rect 4668 924 4724 958
rect 4758 924 4814 958
rect 4848 924 4904 958
rect 4938 924 4994 958
rect 5028 924 5080 958
rect 4400 868 5080 924
rect 4400 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5080 868
rect 4400 778 5080 834
rect 4400 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5080 778
rect 4400 688 5080 744
rect 4400 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5080 688
rect 4400 598 5080 654
rect 4400 564 4454 598
rect 4488 564 4544 598
rect 4578 564 4634 598
rect 4668 564 4724 598
rect 4758 564 4814 598
rect 4848 564 4904 598
rect 4938 564 4994 598
rect 5028 564 5080 598
rect 4400 508 5080 564
rect 4400 474 4454 508
rect 4488 474 4544 508
rect 4578 474 4634 508
rect 4668 474 4724 508
rect 4758 474 4814 508
rect 4848 474 4904 508
rect 4938 474 4994 508
rect 5028 474 5080 508
rect 4400 418 5080 474
rect 4400 384 4454 418
rect 4488 384 4544 418
rect 4578 384 4634 418
rect 4668 384 4724 418
rect 4758 384 4814 418
rect 4848 384 4904 418
rect 4938 384 4994 418
rect 5028 384 5080 418
rect 4400 330 5080 384
rect 5760 958 6440 1010
rect 5760 924 5814 958
rect 5848 924 5904 958
rect 5938 924 5994 958
rect 6028 924 6084 958
rect 6118 924 6174 958
rect 6208 924 6264 958
rect 6298 924 6354 958
rect 6388 924 6440 958
rect 5760 868 6440 924
rect 5760 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6440 868
rect 5760 778 6440 834
rect 5760 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6440 778
rect 5760 688 6440 744
rect 5760 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6440 688
rect 5760 598 6440 654
rect 5760 564 5814 598
rect 5848 564 5904 598
rect 5938 564 5994 598
rect 6028 564 6084 598
rect 6118 564 6174 598
rect 6208 564 6264 598
rect 6298 564 6354 598
rect 6388 564 6440 598
rect 5760 508 6440 564
rect 5760 474 5814 508
rect 5848 474 5904 508
rect 5938 474 5994 508
rect 6028 474 6084 508
rect 6118 474 6174 508
rect 6208 474 6264 508
rect 6298 474 6354 508
rect 6388 474 6440 508
rect 5760 418 6440 474
rect 5760 384 5814 418
rect 5848 384 5904 418
rect 5938 384 5994 418
rect 6028 384 6084 418
rect 6118 384 6174 418
rect 6208 384 6264 418
rect 6298 384 6354 418
rect 6388 384 6440 418
rect 5760 330 6440 384
rect 7120 958 7800 1010
rect 7120 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7714 958
rect 7748 924 7800 958
rect 7120 868 7800 924
rect 7120 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7800 868
rect 7120 778 7800 834
rect 7120 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7800 778
rect 7120 688 7800 744
rect 7120 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7800 688
rect 7120 598 7800 654
rect 7120 564 7174 598
rect 7208 564 7264 598
rect 7298 564 7354 598
rect 7388 564 7444 598
rect 7478 564 7534 598
rect 7568 564 7624 598
rect 7658 564 7714 598
rect 7748 564 7800 598
rect 7120 508 7800 564
rect 7120 474 7174 508
rect 7208 474 7264 508
rect 7298 474 7354 508
rect 7388 474 7444 508
rect 7478 474 7534 508
rect 7568 474 7624 508
rect 7658 474 7714 508
rect 7748 474 7800 508
rect 7120 418 7800 474
rect 7120 384 7174 418
rect 7208 384 7264 418
rect 7298 384 7354 418
rect 7388 384 7444 418
rect 7478 384 7534 418
rect 7568 384 7624 418
rect 7658 384 7714 418
rect 7748 384 7800 418
rect 7120 330 7800 384
rect 8480 958 9160 1010
rect 8480 924 8534 958
rect 8568 924 8624 958
rect 8658 924 8714 958
rect 8748 924 8804 958
rect 8838 924 8894 958
rect 8928 924 8984 958
rect 9018 924 9074 958
rect 9108 924 9160 958
rect 8480 868 9160 924
rect 8480 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9160 868
rect 8480 778 9160 834
rect 8480 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9160 778
rect 8480 688 9160 744
rect 8480 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9160 688
rect 8480 598 9160 654
rect 8480 564 8534 598
rect 8568 564 8624 598
rect 8658 564 8714 598
rect 8748 564 8804 598
rect 8838 564 8894 598
rect 8928 564 8984 598
rect 9018 564 9074 598
rect 9108 564 9160 598
rect 8480 508 9160 564
rect 8480 474 8534 508
rect 8568 474 8624 508
rect 8658 474 8714 508
rect 8748 474 8804 508
rect 8838 474 8894 508
rect 8928 474 8984 508
rect 9018 474 9074 508
rect 9108 474 9160 508
rect 8480 418 9160 474
rect 8480 384 8534 418
rect 8568 384 8624 418
rect 8658 384 8714 418
rect 8748 384 8804 418
rect 8838 384 8894 418
rect 8928 384 8984 418
rect 9018 384 9074 418
rect 9108 384 9160 418
rect 8480 330 9160 384
<< ndiffc >>
rect 5160 3250 5200 3290
rect 5160 3150 5200 3190
rect 5360 3250 5400 3290
rect 5360 3150 5400 3190
rect 5560 3250 5600 3290
rect 5560 3150 5600 3190
rect 5760 3250 5800 3290
rect 5760 3150 5800 3190
rect 5960 3250 6000 3290
rect 5960 3150 6000 3190
rect 6160 3250 6200 3290
rect 6160 3150 6200 3190
rect 6360 3250 6400 3290
rect 6520 3250 6560 3290
rect 6360 3150 6400 3190
rect 6520 3150 6560 3190
rect 6720 3250 6760 3290
rect 6720 3150 6760 3190
rect 6920 3250 6960 3290
rect 6920 3150 6960 3190
rect 7120 3250 7160 3290
rect 7120 3150 7160 3190
rect 7320 3250 7360 3290
rect 7320 3150 7360 3190
rect 7520 3250 7560 3290
rect 7520 3150 7560 3190
rect 7720 3250 7760 3290
rect 7720 3150 7760 3190
rect 4680 2700 4720 2740
rect 4680 2600 4720 2640
rect 4680 2500 4720 2540
rect 4680 2400 4720 2440
rect 4680 2300 4720 2340
rect 4680 2200 4720 2240
rect 4680 2100 4720 2140
rect 4680 2000 4720 2040
rect 5560 2700 5600 2740
rect 5560 2600 5600 2640
rect 5560 2500 5600 2540
rect 5560 2400 5600 2440
rect 5560 2300 5600 2340
rect 5560 2200 5600 2240
rect 5560 2100 5600 2140
rect 5560 2000 5600 2040
rect 6440 2700 6480 2740
rect 6440 2600 6480 2640
rect 6440 2500 6480 2540
rect 6440 2400 6480 2440
rect 6440 2300 6480 2340
rect 6440 2200 6480 2240
rect 6440 2100 6480 2140
rect 6440 2000 6480 2040
rect 7320 2700 7360 2740
rect 7320 2600 7360 2640
rect 7320 2500 7360 2540
rect 7320 2400 7360 2440
rect 7320 2300 7360 2340
rect 7320 2200 7360 2240
rect 7320 2100 7360 2140
rect 7320 2000 7360 2040
rect 8200 2700 8240 2740
rect 8200 2600 8240 2640
rect 8200 2500 8240 2540
rect 8200 2400 8240 2440
rect 8200 2300 8240 2340
rect 8200 2200 8240 2240
rect 8200 2100 8240 2140
rect 8200 2000 8240 2040
rect 5380 1640 5420 1680
rect 5380 1540 5420 1580
rect 7460 1640 7500 1680
rect 7460 1540 7500 1580
<< pdiffc >>
rect 4440 5370 4480 5410
rect 4440 5270 4480 5310
rect 4440 5170 4480 5210
rect 4440 5070 4480 5110
rect 4440 4970 4480 5010
rect 4440 4870 4480 4910
rect 4440 4770 4480 4810
rect 4440 4670 4480 4710
rect 4640 5370 4680 5410
rect 4640 5270 4680 5310
rect 4640 5170 4680 5210
rect 4640 5070 4680 5110
rect 4640 4970 4680 5010
rect 4640 4870 4680 4910
rect 4640 4770 4680 4810
rect 4640 4670 4680 4710
rect 4840 5370 4880 5410
rect 4840 5270 4880 5310
rect 4840 5170 4880 5210
rect 4840 5070 4880 5110
rect 4840 4970 4880 5010
rect 4840 4870 4880 4910
rect 4840 4770 4880 4810
rect 4840 4670 4880 4710
rect 5040 5370 5080 5410
rect 5040 5270 5080 5310
rect 5040 5170 5080 5210
rect 5040 5070 5080 5110
rect 5040 4970 5080 5010
rect 5040 4870 5080 4910
rect 5040 4770 5080 4810
rect 5040 4670 5080 4710
rect 5240 5370 5280 5410
rect 5240 5270 5280 5310
rect 5240 5170 5280 5210
rect 5240 5070 5280 5110
rect 5240 4970 5280 5010
rect 5240 4870 5280 4910
rect 5240 4770 5280 4810
rect 5240 4670 5280 4710
rect 5440 5370 5480 5410
rect 5440 5270 5480 5310
rect 5440 5170 5480 5210
rect 5440 5070 5480 5110
rect 5440 4970 5480 5010
rect 5440 4870 5480 4910
rect 5440 4770 5480 4810
rect 5440 4670 5480 4710
rect 5640 5370 5680 5410
rect 5640 5270 5680 5310
rect 5640 5170 5680 5210
rect 5640 5070 5680 5110
rect 5640 4970 5680 5010
rect 5640 4870 5680 4910
rect 5640 4770 5680 4810
rect 5640 4670 5680 4710
rect 5840 5370 5880 5410
rect 5840 5270 5880 5310
rect 5840 5170 5880 5210
rect 5840 5070 5880 5110
rect 5840 4970 5880 5010
rect 5840 4870 5880 4910
rect 5840 4770 5880 4810
rect 5840 4670 5880 4710
rect 6040 5370 6080 5410
rect 6040 5270 6080 5310
rect 6040 5170 6080 5210
rect 6040 5070 6080 5110
rect 6040 4970 6080 5010
rect 6040 4870 6080 4910
rect 6040 4770 6080 4810
rect 6040 4670 6080 4710
rect 6240 5370 6280 5410
rect 6240 5270 6280 5310
rect 6240 5170 6280 5210
rect 6240 5070 6280 5110
rect 6240 4970 6280 5010
rect 6240 4870 6280 4910
rect 6240 4770 6280 4810
rect 6240 4670 6280 4710
rect 6440 5370 6480 5410
rect 6440 5270 6480 5310
rect 6440 5170 6480 5210
rect 6440 5070 6480 5110
rect 6440 4970 6480 5010
rect 6440 4870 6480 4910
rect 6440 4770 6480 4810
rect 6440 4670 6480 4710
rect 6640 5370 6680 5410
rect 6640 5270 6680 5310
rect 6640 5170 6680 5210
rect 6640 5070 6680 5110
rect 6640 4970 6680 5010
rect 6640 4870 6680 4910
rect 6640 4770 6680 4810
rect 6640 4670 6680 4710
rect 6840 5370 6880 5410
rect 6840 5270 6880 5310
rect 6840 5170 6880 5210
rect 6840 5070 6880 5110
rect 6840 4970 6880 5010
rect 6840 4870 6880 4910
rect 6840 4770 6880 4810
rect 6840 4670 6880 4710
rect 7040 5370 7080 5410
rect 7040 5270 7080 5310
rect 7040 5170 7080 5210
rect 7040 5070 7080 5110
rect 7040 4970 7080 5010
rect 7040 4870 7080 4910
rect 7040 4770 7080 4810
rect 7040 4670 7080 4710
rect 7240 5370 7280 5410
rect 7240 5270 7280 5310
rect 7240 5170 7280 5210
rect 7240 5070 7280 5110
rect 7240 4970 7280 5010
rect 7240 4870 7280 4910
rect 7240 4770 7280 4810
rect 7240 4670 7280 4710
rect 7440 5370 7480 5410
rect 7440 5270 7480 5310
rect 7440 5170 7480 5210
rect 7440 5070 7480 5110
rect 7440 4970 7480 5010
rect 7440 4870 7480 4910
rect 7440 4770 7480 4810
rect 7440 4670 7480 4710
rect 7640 5370 7680 5410
rect 7640 5270 7680 5310
rect 7640 5170 7680 5210
rect 7640 5070 7680 5110
rect 7640 4970 7680 5010
rect 7640 4870 7680 4910
rect 7640 4770 7680 4810
rect 7640 4670 7680 4710
rect 7840 5370 7880 5410
rect 7840 5270 7880 5310
rect 7840 5170 7880 5210
rect 7840 5070 7880 5110
rect 7840 4970 7880 5010
rect 7840 4870 7880 4910
rect 7840 4770 7880 4810
rect 7840 4670 7880 4710
rect 8040 5370 8080 5410
rect 8040 5270 8080 5310
rect 8040 5170 8080 5210
rect 8040 5070 8080 5110
rect 8040 4970 8080 5010
rect 8040 4870 8080 4910
rect 8040 4770 8080 4810
rect 8040 4670 8080 4710
rect 8240 5370 8280 5410
rect 8240 5270 8280 5310
rect 8240 5170 8280 5210
rect 8240 5070 8280 5110
rect 8240 4970 8280 5010
rect 8240 4870 8280 4910
rect 8240 4770 8280 4810
rect 8240 4670 8280 4710
rect 8440 5370 8480 5410
rect 8440 5270 8480 5310
rect 8440 5170 8480 5210
rect 8440 5070 8480 5110
rect 8440 4970 8480 5010
rect 8440 4870 8480 4910
rect 8440 4770 8480 4810
rect 8440 4670 8480 4710
rect 4480 4060 4520 4100
rect 4480 3960 4520 4000
rect 4480 3860 4520 3900
rect 4480 3760 4520 3800
rect 4680 4060 4720 4100
rect 4680 3960 4720 4000
rect 4680 3860 4720 3900
rect 4680 3760 4720 3800
rect 4880 4060 4920 4100
rect 4880 3960 4920 4000
rect 4880 3860 4920 3900
rect 4880 3760 4920 3800
rect 5080 4060 5120 4100
rect 5080 3960 5120 4000
rect 5080 3860 5120 3900
rect 5080 3760 5120 3800
rect 5280 4060 5320 4100
rect 5280 3960 5320 4000
rect 5280 3860 5320 3900
rect 5280 3760 5320 3800
rect 5480 4060 5520 4100
rect 5480 3960 5520 4000
rect 5480 3860 5520 3900
rect 5480 3760 5520 3800
rect 5680 4060 5720 4100
rect 5840 4060 5880 4100
rect 5680 3960 5720 4000
rect 5840 3960 5880 4000
rect 5680 3860 5720 3900
rect 5840 3860 5880 3900
rect 5680 3760 5720 3800
rect 5840 3760 5880 3800
rect 6040 4060 6080 4100
rect 6040 3960 6080 4000
rect 6040 3860 6080 3900
rect 6040 3760 6080 3800
rect 6240 4060 6280 4100
rect 6240 3960 6280 4000
rect 6240 3860 6280 3900
rect 6240 3760 6280 3800
rect 6440 4060 6480 4100
rect 6440 3960 6480 4000
rect 6440 3860 6480 3900
rect 6440 3760 6480 3800
rect 6640 4060 6680 4100
rect 6640 3960 6680 4000
rect 6640 3860 6680 3900
rect 6640 3760 6680 3800
rect 6840 4060 6880 4100
rect 6840 3960 6880 4000
rect 6840 3860 6880 3900
rect 6840 3760 6880 3800
rect 7040 4060 7080 4100
rect 7200 4060 7240 4100
rect 7040 3960 7080 4000
rect 7200 3960 7240 4000
rect 7040 3860 7080 3900
rect 7200 3860 7240 3900
rect 7040 3760 7080 3800
rect 7200 3760 7240 3800
rect 7400 4060 7440 4100
rect 7400 3960 7440 4000
rect 7400 3860 7440 3900
rect 7400 3760 7440 3800
rect 7600 4060 7640 4100
rect 7600 3960 7640 4000
rect 7600 3860 7640 3900
rect 7600 3760 7640 3800
rect 7800 4060 7840 4100
rect 7800 3960 7840 4000
rect 7800 3860 7840 3900
rect 7800 3760 7840 3800
rect 8000 4060 8040 4100
rect 8000 3960 8040 4000
rect 8000 3860 8040 3900
rect 8000 3760 8040 3800
rect 8200 4060 8240 4100
rect 8200 3960 8240 4000
rect 8200 3860 8240 3900
rect 8200 3760 8240 3800
rect 8400 4060 8440 4100
rect 8400 3960 8440 4000
rect 8400 3860 8440 3900
rect 8400 3760 8440 3800
rect 8770 4060 8810 4100
rect 8770 3960 8810 4000
rect 8770 3860 8810 3900
rect 8770 3760 8810 3800
rect 8880 4060 8920 4100
rect 8880 3960 8920 4000
rect 8880 3860 8920 3900
rect 8880 3760 8920 3800
rect 9020 4060 9060 4100
rect 9020 3960 9060 4000
rect 9020 3860 9060 3900
rect 9020 3760 9060 3800
rect 9130 4060 9170 4100
rect 9130 3960 9170 4000
rect 9130 3860 9170 3900
rect 9130 3760 9170 3800
rect 1734 924 1768 958
rect 1824 924 1858 958
rect 1914 924 1948 958
rect 2004 924 2038 958
rect 2094 924 2128 958
rect 2184 924 2218 958
rect 2274 924 2308 958
rect 1734 834 1768 868
rect 1824 834 1858 868
rect 1914 834 1948 868
rect 2004 834 2038 868
rect 2094 834 2128 868
rect 2184 834 2218 868
rect 2274 834 2308 868
rect 1734 744 1768 778
rect 1824 744 1858 778
rect 1914 744 1948 778
rect 2004 744 2038 778
rect 2094 744 2128 778
rect 2184 744 2218 778
rect 2274 744 2308 778
rect 1734 654 1768 688
rect 1824 654 1858 688
rect 1914 654 1948 688
rect 2004 654 2038 688
rect 2094 654 2128 688
rect 2184 654 2218 688
rect 2274 654 2308 688
rect 1734 564 1768 598
rect 1824 564 1858 598
rect 1914 564 1948 598
rect 2004 564 2038 598
rect 2094 564 2128 598
rect 2184 564 2218 598
rect 2274 564 2308 598
rect 1734 474 1768 508
rect 1824 474 1858 508
rect 1914 474 1948 508
rect 2004 474 2038 508
rect 2094 474 2128 508
rect 2184 474 2218 508
rect 2274 474 2308 508
rect 1734 384 1768 418
rect 1824 384 1858 418
rect 1914 384 1948 418
rect 2004 384 2038 418
rect 2094 384 2128 418
rect 2184 384 2218 418
rect 2274 384 2308 418
rect 3094 924 3128 958
rect 3184 924 3218 958
rect 3274 924 3308 958
rect 3364 924 3398 958
rect 3454 924 3488 958
rect 3544 924 3578 958
rect 3634 924 3668 958
rect 3094 834 3128 868
rect 3184 834 3218 868
rect 3274 834 3308 868
rect 3364 834 3398 868
rect 3454 834 3488 868
rect 3544 834 3578 868
rect 3634 834 3668 868
rect 3094 744 3128 778
rect 3184 744 3218 778
rect 3274 744 3308 778
rect 3364 744 3398 778
rect 3454 744 3488 778
rect 3544 744 3578 778
rect 3634 744 3668 778
rect 3094 654 3128 688
rect 3184 654 3218 688
rect 3274 654 3308 688
rect 3364 654 3398 688
rect 3454 654 3488 688
rect 3544 654 3578 688
rect 3634 654 3668 688
rect 3094 564 3128 598
rect 3184 564 3218 598
rect 3274 564 3308 598
rect 3364 564 3398 598
rect 3454 564 3488 598
rect 3544 564 3578 598
rect 3634 564 3668 598
rect 3094 474 3128 508
rect 3184 474 3218 508
rect 3274 474 3308 508
rect 3364 474 3398 508
rect 3454 474 3488 508
rect 3544 474 3578 508
rect 3634 474 3668 508
rect 3094 384 3128 418
rect 3184 384 3218 418
rect 3274 384 3308 418
rect 3364 384 3398 418
rect 3454 384 3488 418
rect 3544 384 3578 418
rect 3634 384 3668 418
rect 4454 924 4488 958
rect 4544 924 4578 958
rect 4634 924 4668 958
rect 4724 924 4758 958
rect 4814 924 4848 958
rect 4904 924 4938 958
rect 4994 924 5028 958
rect 4454 834 4488 868
rect 4544 834 4578 868
rect 4634 834 4668 868
rect 4724 834 4758 868
rect 4814 834 4848 868
rect 4904 834 4938 868
rect 4994 834 5028 868
rect 4454 744 4488 778
rect 4544 744 4578 778
rect 4634 744 4668 778
rect 4724 744 4758 778
rect 4814 744 4848 778
rect 4904 744 4938 778
rect 4994 744 5028 778
rect 4454 654 4488 688
rect 4544 654 4578 688
rect 4634 654 4668 688
rect 4724 654 4758 688
rect 4814 654 4848 688
rect 4904 654 4938 688
rect 4994 654 5028 688
rect 4454 564 4488 598
rect 4544 564 4578 598
rect 4634 564 4668 598
rect 4724 564 4758 598
rect 4814 564 4848 598
rect 4904 564 4938 598
rect 4994 564 5028 598
rect 4454 474 4488 508
rect 4544 474 4578 508
rect 4634 474 4668 508
rect 4724 474 4758 508
rect 4814 474 4848 508
rect 4904 474 4938 508
rect 4994 474 5028 508
rect 4454 384 4488 418
rect 4544 384 4578 418
rect 4634 384 4668 418
rect 4724 384 4758 418
rect 4814 384 4848 418
rect 4904 384 4938 418
rect 4994 384 5028 418
rect 5814 924 5848 958
rect 5904 924 5938 958
rect 5994 924 6028 958
rect 6084 924 6118 958
rect 6174 924 6208 958
rect 6264 924 6298 958
rect 6354 924 6388 958
rect 5814 834 5848 868
rect 5904 834 5938 868
rect 5994 834 6028 868
rect 6084 834 6118 868
rect 6174 834 6208 868
rect 6264 834 6298 868
rect 6354 834 6388 868
rect 5814 744 5848 778
rect 5904 744 5938 778
rect 5994 744 6028 778
rect 6084 744 6118 778
rect 6174 744 6208 778
rect 6264 744 6298 778
rect 6354 744 6388 778
rect 5814 654 5848 688
rect 5904 654 5938 688
rect 5994 654 6028 688
rect 6084 654 6118 688
rect 6174 654 6208 688
rect 6264 654 6298 688
rect 6354 654 6388 688
rect 5814 564 5848 598
rect 5904 564 5938 598
rect 5994 564 6028 598
rect 6084 564 6118 598
rect 6174 564 6208 598
rect 6264 564 6298 598
rect 6354 564 6388 598
rect 5814 474 5848 508
rect 5904 474 5938 508
rect 5994 474 6028 508
rect 6084 474 6118 508
rect 6174 474 6208 508
rect 6264 474 6298 508
rect 6354 474 6388 508
rect 5814 384 5848 418
rect 5904 384 5938 418
rect 5994 384 6028 418
rect 6084 384 6118 418
rect 6174 384 6208 418
rect 6264 384 6298 418
rect 6354 384 6388 418
rect 7174 924 7208 958
rect 7264 924 7298 958
rect 7354 924 7388 958
rect 7444 924 7478 958
rect 7534 924 7568 958
rect 7624 924 7658 958
rect 7714 924 7748 958
rect 7174 834 7208 868
rect 7264 834 7298 868
rect 7354 834 7388 868
rect 7444 834 7478 868
rect 7534 834 7568 868
rect 7624 834 7658 868
rect 7714 834 7748 868
rect 7174 744 7208 778
rect 7264 744 7298 778
rect 7354 744 7388 778
rect 7444 744 7478 778
rect 7534 744 7568 778
rect 7624 744 7658 778
rect 7714 744 7748 778
rect 7174 654 7208 688
rect 7264 654 7298 688
rect 7354 654 7388 688
rect 7444 654 7478 688
rect 7534 654 7568 688
rect 7624 654 7658 688
rect 7714 654 7748 688
rect 7174 564 7208 598
rect 7264 564 7298 598
rect 7354 564 7388 598
rect 7444 564 7478 598
rect 7534 564 7568 598
rect 7624 564 7658 598
rect 7714 564 7748 598
rect 7174 474 7208 508
rect 7264 474 7298 508
rect 7354 474 7388 508
rect 7444 474 7478 508
rect 7534 474 7568 508
rect 7624 474 7658 508
rect 7714 474 7748 508
rect 7174 384 7208 418
rect 7264 384 7298 418
rect 7354 384 7388 418
rect 7444 384 7478 418
rect 7534 384 7568 418
rect 7624 384 7658 418
rect 7714 384 7748 418
rect 8534 924 8568 958
rect 8624 924 8658 958
rect 8714 924 8748 958
rect 8804 924 8838 958
rect 8894 924 8928 958
rect 8984 924 9018 958
rect 9074 924 9108 958
rect 8534 834 8568 868
rect 8624 834 8658 868
rect 8714 834 8748 868
rect 8804 834 8838 868
rect 8894 834 8928 868
rect 8984 834 9018 868
rect 9074 834 9108 868
rect 8534 744 8568 778
rect 8624 744 8658 778
rect 8714 744 8748 778
rect 8804 744 8838 778
rect 8894 744 8928 778
rect 8984 744 9018 778
rect 9074 744 9108 778
rect 8534 654 8568 688
rect 8624 654 8658 688
rect 8714 654 8748 688
rect 8804 654 8838 688
rect 8894 654 8928 688
rect 8984 654 9018 688
rect 9074 654 9108 688
rect 8534 564 8568 598
rect 8624 564 8658 598
rect 8714 564 8748 598
rect 8804 564 8838 598
rect 8894 564 8928 598
rect 8984 564 9018 598
rect 9074 564 9108 598
rect 8534 474 8568 508
rect 8624 474 8658 508
rect 8714 474 8748 508
rect 8804 474 8838 508
rect 8894 474 8928 508
rect 8984 474 9018 508
rect 9074 474 9108 508
rect 8534 384 8568 418
rect 8624 384 8658 418
rect 8714 384 8748 418
rect 8804 384 8838 418
rect 8894 384 8928 418
rect 8984 384 9018 418
rect 9074 384 9108 418
<< psubdiff >>
rect 5060 3290 5140 3320
rect 5060 3250 5080 3290
rect 5120 3250 5140 3290
rect 5060 3190 5140 3250
rect 5060 3150 5080 3190
rect 5120 3150 5140 3190
rect 5060 3120 5140 3150
rect 6420 3290 6500 3320
rect 6420 3250 6440 3290
rect 6480 3250 6500 3290
rect 6420 3190 6500 3250
rect 6420 3150 6440 3190
rect 6480 3150 6500 3190
rect 6420 3120 6500 3150
rect 7780 3290 7860 3320
rect 7780 3250 7800 3290
rect 7840 3250 7860 3290
rect 7780 3190 7860 3250
rect 7780 3150 7800 3190
rect 7840 3150 7860 3190
rect 7780 3120 7860 3150
rect 4580 2740 4660 2770
rect 4580 2700 4600 2740
rect 4640 2700 4660 2740
rect 4580 2640 4660 2700
rect 4580 2600 4600 2640
rect 4640 2600 4660 2640
rect 4580 2540 4660 2600
rect 4580 2500 4600 2540
rect 4640 2500 4660 2540
rect 4580 2440 4660 2500
rect 4580 2400 4600 2440
rect 4640 2400 4660 2440
rect 4580 2340 4660 2400
rect 4580 2300 4600 2340
rect 4640 2300 4660 2340
rect 4580 2240 4660 2300
rect 4580 2200 4600 2240
rect 4640 2200 4660 2240
rect 4580 2140 4660 2200
rect 4580 2100 4600 2140
rect 4640 2100 4660 2140
rect 4580 2040 4660 2100
rect 4580 2000 4600 2040
rect 4640 2000 4660 2040
rect 4580 1970 4660 2000
rect 8260 2740 8340 2770
rect 8260 2700 8280 2740
rect 8320 2700 8340 2740
rect 8260 2640 8340 2700
rect 8260 2600 8280 2640
rect 8320 2600 8340 2640
rect 8260 2540 8340 2600
rect 8260 2500 8280 2540
rect 8320 2500 8340 2540
rect 8260 2440 8340 2500
rect 8260 2400 8280 2440
rect 8320 2400 8340 2440
rect 8260 2340 8340 2400
rect 8260 2300 8280 2340
rect 8320 2300 8340 2340
rect 8260 2240 8340 2300
rect 8260 2200 8280 2240
rect 8320 2200 8340 2240
rect 8260 2140 8340 2200
rect 8260 2100 8280 2140
rect 8320 2100 8340 2140
rect 8260 2040 8340 2100
rect 8260 2000 8280 2040
rect 8320 2000 8340 2040
rect 8260 1970 8340 2000
rect 7520 1680 7600 1710
rect 7520 1640 7540 1680
rect 7580 1640 7600 1680
rect 7520 1580 7600 1640
rect 7520 1540 7540 1580
rect 7580 1540 7600 1580
rect 7520 1510 7600 1540
rect 1376 1279 2664 1314
rect 1376 1256 1506 1279
rect 1376 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2664 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2664 1256
rect 1376 1213 2664 1222
rect 1376 1166 1477 1213
rect 1376 1132 1410 1166
rect 1444 1132 1477 1166
rect 2563 1166 2664 1213
rect 1376 1076 1477 1132
rect 1376 1042 1410 1076
rect 1444 1042 1477 1076
rect 1376 986 1477 1042
rect 1376 952 1410 986
rect 1444 952 1477 986
rect 1376 896 1477 952
rect 1376 862 1410 896
rect 1444 862 1477 896
rect 1376 806 1477 862
rect 1376 772 1410 806
rect 1444 772 1477 806
rect 1376 716 1477 772
rect 1376 682 1410 716
rect 1444 682 1477 716
rect 1376 626 1477 682
rect 1376 592 1410 626
rect 1444 592 1477 626
rect 1376 536 1477 592
rect 1376 502 1410 536
rect 1444 502 1477 536
rect 1376 446 1477 502
rect 1376 412 1410 446
rect 1444 412 1477 446
rect 1376 356 1477 412
rect 1376 322 1410 356
rect 1444 322 1477 356
rect 1376 266 1477 322
rect 1376 232 1410 266
rect 1444 232 1477 266
rect 1376 176 1477 232
rect 2563 1132 2597 1166
rect 2631 1132 2664 1166
rect 2563 1076 2664 1132
rect 2563 1042 2597 1076
rect 2631 1042 2664 1076
rect 2563 986 2664 1042
rect 2563 952 2597 986
rect 2631 952 2664 986
rect 2563 896 2664 952
rect 2563 862 2597 896
rect 2631 862 2664 896
rect 2563 806 2664 862
rect 2563 772 2597 806
rect 2631 772 2664 806
rect 2563 716 2664 772
rect 2563 682 2597 716
rect 2631 682 2664 716
rect 2563 626 2664 682
rect 2563 592 2597 626
rect 2631 592 2664 626
rect 2563 536 2664 592
rect 2563 502 2597 536
rect 2631 502 2664 536
rect 2563 446 2664 502
rect 2563 412 2597 446
rect 2631 412 2664 446
rect 2563 356 2664 412
rect 2563 322 2597 356
rect 2631 322 2664 356
rect 2563 266 2664 322
rect 2563 232 2597 266
rect 2631 232 2664 266
rect 1376 142 1410 176
rect 1444 142 1477 176
rect 1376 127 1477 142
rect 2563 176 2664 232
rect 2563 142 2597 176
rect 2631 142 2664 176
rect 2563 127 2664 142
rect 1376 92 2664 127
rect 40 50 80 90
rect 1376 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 90 2586 92
rect 2530 58 2600 90
rect 2620 58 2664 92
rect 1376 26 2664 58
rect 2736 1279 4024 1314
rect 2736 1256 2866 1279
rect 2736 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4024 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4024 1256
rect 2736 1213 4024 1222
rect 2736 1166 2837 1213
rect 2736 1132 2770 1166
rect 2804 1132 2837 1166
rect 3923 1166 4024 1213
rect 2736 1076 2837 1132
rect 2736 1042 2770 1076
rect 2804 1042 2837 1076
rect 2736 986 2837 1042
rect 2736 952 2770 986
rect 2804 952 2837 986
rect 2736 896 2837 952
rect 2736 862 2770 896
rect 2804 862 2837 896
rect 2736 806 2837 862
rect 2736 772 2770 806
rect 2804 772 2837 806
rect 2736 716 2837 772
rect 2736 682 2770 716
rect 2804 682 2837 716
rect 2736 626 2837 682
rect 2736 592 2770 626
rect 2804 592 2837 626
rect 2736 536 2837 592
rect 2736 502 2770 536
rect 2804 502 2837 536
rect 2736 446 2837 502
rect 2736 412 2770 446
rect 2804 412 2837 446
rect 2736 356 2837 412
rect 2736 322 2770 356
rect 2804 322 2837 356
rect 2736 266 2837 322
rect 2736 232 2770 266
rect 2804 232 2837 266
rect 2736 176 2837 232
rect 3923 1132 3957 1166
rect 3991 1132 4024 1166
rect 3923 1076 4024 1132
rect 3923 1042 3957 1076
rect 3991 1042 4024 1076
rect 3923 986 4024 1042
rect 3923 952 3957 986
rect 3991 952 4024 986
rect 3923 896 4024 952
rect 3923 862 3957 896
rect 3991 862 4024 896
rect 3923 806 4024 862
rect 3923 772 3957 806
rect 3991 772 4024 806
rect 3923 716 4024 772
rect 3923 682 3957 716
rect 3991 682 4024 716
rect 3923 626 4024 682
rect 3923 592 3957 626
rect 3991 592 4024 626
rect 3923 536 4024 592
rect 3923 502 3957 536
rect 3991 502 4024 536
rect 3923 446 4024 502
rect 3923 412 3957 446
rect 3991 412 4024 446
rect 3923 356 4024 412
rect 3923 322 3957 356
rect 3991 322 4024 356
rect 3923 266 4024 322
rect 3923 232 3957 266
rect 3991 232 4024 266
rect 2736 142 2770 176
rect 2804 142 2837 176
rect 2736 127 2837 142
rect 3923 176 4024 232
rect 3923 142 3957 176
rect 3991 142 4024 176
rect 3923 127 4024 142
rect 2736 92 4024 127
rect 4096 1279 5384 1314
rect 4096 1256 4226 1279
rect 4096 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5384 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5384 1256
rect 4096 1213 5384 1222
rect 4096 1166 4197 1213
rect 4096 1132 4130 1166
rect 4164 1132 4197 1166
rect 5283 1166 5384 1213
rect 4096 1076 4197 1132
rect 4096 1042 4130 1076
rect 4164 1042 4197 1076
rect 4096 986 4197 1042
rect 4096 952 4130 986
rect 4164 952 4197 986
rect 4096 896 4197 952
rect 4096 862 4130 896
rect 4164 862 4197 896
rect 4096 806 4197 862
rect 4096 772 4130 806
rect 4164 772 4197 806
rect 4096 716 4197 772
rect 4096 682 4130 716
rect 4164 682 4197 716
rect 4096 626 4197 682
rect 4096 592 4130 626
rect 4164 592 4197 626
rect 4096 536 4197 592
rect 4096 502 4130 536
rect 4164 502 4197 536
rect 4096 446 4197 502
rect 4096 412 4130 446
rect 4164 412 4197 446
rect 4096 356 4197 412
rect 4096 322 4130 356
rect 4164 322 4197 356
rect 4096 266 4197 322
rect 4096 232 4130 266
rect 4164 232 4197 266
rect 4096 176 4197 232
rect 5283 1132 5317 1166
rect 5351 1132 5384 1166
rect 5283 1076 5384 1132
rect 5283 1042 5317 1076
rect 5351 1042 5384 1076
rect 5283 986 5384 1042
rect 5283 952 5317 986
rect 5351 952 5384 986
rect 5283 896 5384 952
rect 5283 862 5317 896
rect 5351 862 5384 896
rect 5283 806 5384 862
rect 5283 772 5317 806
rect 5351 772 5384 806
rect 5283 716 5384 772
rect 5283 682 5317 716
rect 5351 682 5384 716
rect 5283 626 5384 682
rect 5283 592 5317 626
rect 5351 592 5384 626
rect 5283 536 5384 592
rect 5283 502 5317 536
rect 5351 502 5384 536
rect 5283 446 5384 502
rect 5283 412 5317 446
rect 5351 412 5384 446
rect 5283 356 5384 412
rect 5283 322 5317 356
rect 5351 322 5384 356
rect 5283 266 5384 322
rect 5283 232 5317 266
rect 5351 232 5384 266
rect 4096 142 4130 176
rect 4164 142 4197 176
rect 4096 127 4197 142
rect 5283 176 5384 232
rect 5283 142 5317 176
rect 5351 142 5384 176
rect 5283 127 5384 142
rect 4096 92 5384 127
rect 5456 1279 6744 1314
rect 5456 1256 5586 1279
rect 5456 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6744 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6744 1256
rect 5456 1213 6744 1222
rect 5456 1166 5557 1213
rect 5456 1132 5490 1166
rect 5524 1132 5557 1166
rect 6643 1166 6744 1213
rect 5456 1076 5557 1132
rect 5456 1042 5490 1076
rect 5524 1042 5557 1076
rect 5456 986 5557 1042
rect 5456 952 5490 986
rect 5524 952 5557 986
rect 5456 896 5557 952
rect 5456 862 5490 896
rect 5524 862 5557 896
rect 5456 806 5557 862
rect 5456 772 5490 806
rect 5524 772 5557 806
rect 5456 716 5557 772
rect 5456 682 5490 716
rect 5524 682 5557 716
rect 5456 626 5557 682
rect 5456 592 5490 626
rect 5524 592 5557 626
rect 5456 536 5557 592
rect 5456 502 5490 536
rect 5524 502 5557 536
rect 5456 446 5557 502
rect 5456 412 5490 446
rect 5524 412 5557 446
rect 5456 356 5557 412
rect 5456 322 5490 356
rect 5524 322 5557 356
rect 5456 266 5557 322
rect 5456 232 5490 266
rect 5524 232 5557 266
rect 5456 176 5557 232
rect 6643 1132 6677 1166
rect 6711 1132 6744 1166
rect 6643 1076 6744 1132
rect 6643 1042 6677 1076
rect 6711 1042 6744 1076
rect 6643 986 6744 1042
rect 6643 952 6677 986
rect 6711 952 6744 986
rect 6643 896 6744 952
rect 6643 862 6677 896
rect 6711 862 6744 896
rect 6643 806 6744 862
rect 6643 772 6677 806
rect 6711 772 6744 806
rect 6643 716 6744 772
rect 6643 682 6677 716
rect 6711 682 6744 716
rect 6643 626 6744 682
rect 6643 592 6677 626
rect 6711 592 6744 626
rect 6643 536 6744 592
rect 6643 502 6677 536
rect 6711 502 6744 536
rect 6643 446 6744 502
rect 6643 412 6677 446
rect 6711 412 6744 446
rect 6643 356 6744 412
rect 6643 322 6677 356
rect 6711 322 6744 356
rect 6643 266 6744 322
rect 6643 232 6677 266
rect 6711 232 6744 266
rect 5456 142 5490 176
rect 5524 142 5557 176
rect 5456 127 5557 142
rect 6643 176 6744 232
rect 6643 142 6677 176
rect 6711 142 6744 176
rect 6643 127 6744 142
rect 5456 92 6744 127
rect 6816 1279 8104 1314
rect 6816 1256 6946 1279
rect 6816 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8104 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8104 1256
rect 6816 1213 8104 1222
rect 6816 1166 6917 1213
rect 6816 1132 6850 1166
rect 6884 1132 6917 1166
rect 8003 1166 8104 1213
rect 6816 1076 6917 1132
rect 6816 1042 6850 1076
rect 6884 1042 6917 1076
rect 6816 986 6917 1042
rect 6816 952 6850 986
rect 6884 952 6917 986
rect 6816 896 6917 952
rect 6816 862 6850 896
rect 6884 862 6917 896
rect 6816 806 6917 862
rect 6816 772 6850 806
rect 6884 772 6917 806
rect 6816 716 6917 772
rect 6816 682 6850 716
rect 6884 682 6917 716
rect 6816 626 6917 682
rect 6816 592 6850 626
rect 6884 592 6917 626
rect 6816 536 6917 592
rect 6816 502 6850 536
rect 6884 502 6917 536
rect 6816 446 6917 502
rect 6816 412 6850 446
rect 6884 412 6917 446
rect 6816 356 6917 412
rect 6816 322 6850 356
rect 6884 322 6917 356
rect 6816 266 6917 322
rect 6816 232 6850 266
rect 6884 232 6917 266
rect 6816 176 6917 232
rect 8003 1132 8037 1166
rect 8071 1132 8104 1166
rect 8003 1076 8104 1132
rect 8003 1042 8037 1076
rect 8071 1042 8104 1076
rect 8003 986 8104 1042
rect 8003 952 8037 986
rect 8071 952 8104 986
rect 8003 896 8104 952
rect 8003 862 8037 896
rect 8071 862 8104 896
rect 8003 806 8104 862
rect 8003 772 8037 806
rect 8071 772 8104 806
rect 8003 716 8104 772
rect 8003 682 8037 716
rect 8071 682 8104 716
rect 8003 626 8104 682
rect 8003 592 8037 626
rect 8071 592 8104 626
rect 8003 536 8104 592
rect 8003 502 8037 536
rect 8071 502 8104 536
rect 8003 446 8104 502
rect 8003 412 8037 446
rect 8071 412 8104 446
rect 8003 356 8104 412
rect 8003 322 8037 356
rect 8071 322 8104 356
rect 8003 266 8104 322
rect 8003 232 8037 266
rect 8071 232 8104 266
rect 6816 142 6850 176
rect 6884 142 6917 176
rect 6816 127 6917 142
rect 8003 176 8104 232
rect 8003 142 8037 176
rect 8071 142 8104 176
rect 8003 127 8104 142
rect 6816 92 8104 127
rect 8176 1279 9464 1314
rect 8176 1256 8306 1279
rect 8176 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9464 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9464 1256
rect 8176 1213 9464 1222
rect 8176 1166 8277 1213
rect 8176 1132 8210 1166
rect 8244 1132 8277 1166
rect 9363 1166 9464 1213
rect 8176 1076 8277 1132
rect 8176 1042 8210 1076
rect 8244 1042 8277 1076
rect 8176 986 8277 1042
rect 8176 952 8210 986
rect 8244 952 8277 986
rect 8176 896 8277 952
rect 8176 862 8210 896
rect 8244 862 8277 896
rect 8176 806 8277 862
rect 8176 772 8210 806
rect 8244 772 8277 806
rect 8176 716 8277 772
rect 8176 682 8210 716
rect 8244 682 8277 716
rect 8176 626 8277 682
rect 8176 592 8210 626
rect 8244 592 8277 626
rect 8176 536 8277 592
rect 8176 502 8210 536
rect 8244 502 8277 536
rect 8176 446 8277 502
rect 8176 412 8210 446
rect 8244 412 8277 446
rect 8176 356 8277 412
rect 8176 322 8210 356
rect 8244 322 8277 356
rect 8176 266 8277 322
rect 8176 232 8210 266
rect 8244 232 8277 266
rect 8176 176 8277 232
rect 9363 1132 9397 1166
rect 9431 1132 9464 1166
rect 9363 1076 9464 1132
rect 9363 1042 9397 1076
rect 9431 1042 9464 1076
rect 9363 986 9464 1042
rect 9363 952 9397 986
rect 9431 952 9464 986
rect 9363 896 9464 952
rect 9363 862 9397 896
rect 9431 862 9464 896
rect 9363 806 9464 862
rect 9363 772 9397 806
rect 9431 772 9464 806
rect 9363 716 9464 772
rect 9363 682 9397 716
rect 9431 682 9464 716
rect 9363 626 9464 682
rect 9363 592 9397 626
rect 9431 592 9464 626
rect 9363 536 9464 592
rect 9363 502 9397 536
rect 9431 502 9464 536
rect 9363 446 9464 502
rect 9363 412 9397 446
rect 9431 412 9464 446
rect 9363 356 9464 412
rect 9363 322 9397 356
rect 9431 322 9464 356
rect 9363 266 9464 322
rect 9363 232 9397 266
rect 9431 232 9464 266
rect 8176 142 8210 176
rect 8244 142 8277 176
rect 8176 127 8277 142
rect 9363 176 9464 232
rect 9363 142 9397 176
rect 9431 142 9464 176
rect 9363 127 9464 142
rect 8176 92 9464 127
rect 2736 90 2766 92
rect 2736 58 2780 90
rect 2800 58 2866 92
rect 2900 90 2946 92
rect 2900 58 2956 90
rect 2990 58 3046 92
rect 3080 90 3126 92
rect 3080 58 3136 90
rect 3170 58 3226 92
rect 3260 90 3306 92
rect 3260 58 3316 90
rect 3350 58 3406 92
rect 3440 90 3486 92
rect 3440 58 3496 90
rect 3530 58 3586 92
rect 3620 90 3666 92
rect 3620 58 3676 90
rect 3710 58 3766 92
rect 3800 90 3846 92
rect 3800 58 3856 90
rect 3890 58 3970 92
rect 3980 58 4024 92
rect 4096 58 4150 92
rect 4160 90 4206 92
rect 4160 58 4220 90
rect 4260 58 4316 92
rect 4350 90 4386 92
rect 4350 58 4400 90
rect 4440 58 4496 92
rect 4530 90 4566 92
rect 4530 58 4580 90
rect 4620 58 4676 92
rect 4710 90 4746 92
rect 4710 58 4760 90
rect 4800 58 4856 92
rect 4890 90 4926 92
rect 4890 58 4940 90
rect 4980 58 5036 92
rect 5070 90 5106 92
rect 5070 58 5120 90
rect 5160 58 5216 92
rect 5250 90 5286 92
rect 5250 58 5300 90
rect 5330 58 5384 92
rect 5456 90 5466 92
rect 5456 58 5480 90
rect 5510 58 5586 92
rect 5620 90 5646 92
rect 5620 58 5660 90
rect 5710 58 5766 92
rect 5800 90 5826 92
rect 5800 58 5840 90
rect 5890 58 5946 92
rect 5980 90 6006 92
rect 5980 58 6020 90
rect 6070 58 6126 92
rect 6160 90 6186 92
rect 6160 58 6200 90
rect 6250 58 6306 92
rect 6340 90 6366 92
rect 6340 58 6380 90
rect 6430 58 6486 92
rect 6520 90 6546 92
rect 6520 58 6560 90
rect 6610 58 6670 92
rect 6700 90 6726 92
rect 6700 58 6740 90
rect 6816 58 6850 92
rect 6880 90 6906 92
rect 6880 58 6920 90
rect 6980 58 7030 92
rect 7070 90 7086 92
rect 7070 58 7100 90
rect 7160 58 7210 92
rect 7250 90 7266 92
rect 7250 58 7280 90
rect 7340 58 7390 92
rect 7430 90 7446 92
rect 7430 58 7460 90
rect 7520 58 7570 92
rect 7610 90 7626 92
rect 7610 58 7640 90
rect 7700 58 7750 92
rect 7790 90 7806 92
rect 7790 58 7820 90
rect 7880 58 7930 92
rect 7970 90 7986 92
rect 7970 58 8000 90
rect 8030 58 8104 92
rect 8176 58 8180 90
rect 8210 58 8290 92
rect 8340 90 8346 92
rect 8340 58 8360 90
rect 8390 58 8396 92
rect 8430 58 8470 92
rect 8520 90 8526 92
rect 8520 58 8540 90
rect 8570 58 8576 92
rect 8610 58 8650 92
rect 8700 90 8706 92
rect 8700 58 8720 90
rect 8750 58 8756 92
rect 8790 58 8830 92
rect 8880 90 8886 92
rect 8880 58 8900 90
rect 8930 58 8936 92
rect 8970 58 9010 92
rect 9060 90 9066 92
rect 9060 58 9080 90
rect 9110 58 9116 92
rect 9150 58 9190 92
rect 9240 90 9246 92
rect 9240 58 9260 90
rect 9290 58 9296 92
rect 9330 58 9370 92
rect 9420 90 9426 92
rect 9400 58 9440 90
rect 2736 26 4024 58
rect 4096 26 5384 58
rect 5456 26 6744 58
rect 6816 26 8104 58
rect 8176 26 9464 58
<< nsubdiff >>
rect 4340 5410 4420 5440
rect 4340 5370 4360 5410
rect 4400 5370 4420 5410
rect 4340 5310 4420 5370
rect 4340 5270 4360 5310
rect 4400 5270 4420 5310
rect 4340 5210 4420 5270
rect 4340 5170 4360 5210
rect 4400 5170 4420 5210
rect 4340 5110 4420 5170
rect 4340 5070 4360 5110
rect 4400 5070 4420 5110
rect 4340 5010 4420 5070
rect 4340 4970 4360 5010
rect 4400 4970 4420 5010
rect 4340 4910 4420 4970
rect 4340 4870 4360 4910
rect 4400 4870 4420 4910
rect 4340 4810 4420 4870
rect 4340 4770 4360 4810
rect 4400 4770 4420 4810
rect 4340 4710 4420 4770
rect 4340 4670 4360 4710
rect 4400 4670 4420 4710
rect 4340 4640 4420 4670
rect 8500 5410 8580 5440
rect 8500 5370 8520 5410
rect 8560 5370 8580 5410
rect 8500 5310 8580 5370
rect 8500 5270 8520 5310
rect 8560 5270 8580 5310
rect 8500 5210 8580 5270
rect 8500 5170 8520 5210
rect 8560 5170 8580 5210
rect 8500 5110 8580 5170
rect 8500 5070 8520 5110
rect 8560 5070 8580 5110
rect 8500 5010 8580 5070
rect 8500 4970 8520 5010
rect 8560 4970 8580 5010
rect 8500 4910 8580 4970
rect 8500 4870 8520 4910
rect 8560 4870 8580 4910
rect 8500 4810 8580 4870
rect 8500 4770 8520 4810
rect 8560 4770 8580 4810
rect 8500 4710 8580 4770
rect 8500 4670 8520 4710
rect 8560 4670 8580 4710
rect 8500 4640 8580 4670
rect 4380 4100 4460 4130
rect 4380 4060 4400 4100
rect 4440 4060 4460 4100
rect 4380 4000 4460 4060
rect 4380 3960 4400 4000
rect 4440 3960 4460 4000
rect 4380 3900 4460 3960
rect 4380 3860 4400 3900
rect 4440 3860 4460 3900
rect 4380 3800 4460 3860
rect 4380 3760 4400 3800
rect 4440 3760 4460 3800
rect 4380 3730 4460 3760
rect 5740 4100 5820 4130
rect 5740 4060 5760 4100
rect 5800 4060 5820 4100
rect 5740 4000 5820 4060
rect 5740 3960 5760 4000
rect 5800 3960 5820 4000
rect 5740 3900 5820 3960
rect 5740 3860 5760 3900
rect 5800 3860 5820 3900
rect 5740 3800 5820 3860
rect 5740 3760 5760 3800
rect 5800 3760 5820 3800
rect 5740 3730 5820 3760
rect 7100 4100 7180 4130
rect 7100 4060 7120 4100
rect 7160 4060 7180 4100
rect 7100 4000 7180 4060
rect 7100 3960 7120 4000
rect 7160 3960 7180 4000
rect 7100 3900 7180 3960
rect 7100 3860 7120 3900
rect 7160 3860 7180 3900
rect 7100 3800 7180 3860
rect 7100 3760 7120 3800
rect 7160 3760 7180 3800
rect 7100 3730 7180 3760
rect 8460 4100 8540 4130
rect 8460 4060 8480 4100
rect 8520 4060 8540 4100
rect 8460 4000 8540 4060
rect 8460 3960 8480 4000
rect 8520 3960 8540 4000
rect 8460 3900 8540 3960
rect 8460 3860 8480 3900
rect 8520 3860 8540 3900
rect 8460 3800 8540 3860
rect 8460 3760 8480 3800
rect 8520 3760 8540 3800
rect 8460 3730 8540 3760
rect 9190 4100 9270 4130
rect 9190 4060 9210 4100
rect 9250 4060 9270 4100
rect 9190 4000 9270 4060
rect 9190 3960 9210 4000
rect 9250 3960 9270 4000
rect 9190 3900 9270 3960
rect 9190 3860 9210 3900
rect 9250 3860 9270 3900
rect 9190 3800 9270 3860
rect 9190 3760 9210 3800
rect 9250 3760 9270 3800
rect 9190 3730 9270 3760
rect 1539 1132 2501 1151
rect 1539 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 2501 1132
rect 1539 1079 2501 1098
rect 1539 1075 1611 1079
rect 1539 1041 1558 1075
rect 1592 1041 1611 1075
rect 1539 985 1611 1041
rect 2429 1056 2501 1079
rect 2429 1022 2448 1056
rect 2482 1022 2501 1056
rect 1539 951 1558 985
rect 1592 951 1611 985
rect 1539 895 1611 951
rect 1539 861 1558 895
rect 1592 861 1611 895
rect 1539 805 1611 861
rect 1539 771 1558 805
rect 1592 771 1611 805
rect 1539 715 1611 771
rect 1539 681 1558 715
rect 1592 681 1611 715
rect 1539 625 1611 681
rect 1539 591 1558 625
rect 1592 591 1611 625
rect 1539 535 1611 591
rect 1539 501 1558 535
rect 1592 501 1611 535
rect 1539 445 1611 501
rect 1539 411 1558 445
rect 1592 411 1611 445
rect 1539 355 1611 411
rect 1539 321 1558 355
rect 1592 321 1611 355
rect 2429 966 2501 1022
rect 2429 932 2448 966
rect 2482 932 2501 966
rect 2429 876 2501 932
rect 2429 842 2448 876
rect 2482 842 2501 876
rect 2429 786 2501 842
rect 2429 752 2448 786
rect 2482 752 2501 786
rect 2429 696 2501 752
rect 2429 662 2448 696
rect 2482 662 2501 696
rect 2429 606 2501 662
rect 2429 572 2448 606
rect 2482 572 2501 606
rect 2429 516 2501 572
rect 2429 482 2448 516
rect 2482 482 2501 516
rect 2429 426 2501 482
rect 2429 392 2448 426
rect 2482 392 2501 426
rect 2429 336 2501 392
rect 1539 261 1611 321
rect 2429 302 2448 336
rect 2482 302 2501 336
rect 2429 261 2501 302
rect 1539 242 2501 261
rect 1539 208 1636 242
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 208 2501 242
rect 1539 189 2501 208
rect 2899 1132 3861 1151
rect 2899 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 3861 1132
rect 2899 1079 3861 1098
rect 2899 1075 2971 1079
rect 2899 1041 2918 1075
rect 2952 1041 2971 1075
rect 2899 985 2971 1041
rect 3789 1056 3861 1079
rect 3789 1022 3808 1056
rect 3842 1022 3861 1056
rect 2899 951 2918 985
rect 2952 951 2971 985
rect 2899 895 2971 951
rect 2899 861 2918 895
rect 2952 861 2971 895
rect 2899 805 2971 861
rect 2899 771 2918 805
rect 2952 771 2971 805
rect 2899 715 2971 771
rect 2899 681 2918 715
rect 2952 681 2971 715
rect 2899 625 2971 681
rect 2899 591 2918 625
rect 2952 591 2971 625
rect 2899 535 2971 591
rect 2899 501 2918 535
rect 2952 501 2971 535
rect 2899 445 2971 501
rect 2899 411 2918 445
rect 2952 411 2971 445
rect 2899 355 2971 411
rect 2899 321 2918 355
rect 2952 321 2971 355
rect 3789 966 3861 1022
rect 3789 932 3808 966
rect 3842 932 3861 966
rect 3789 876 3861 932
rect 3789 842 3808 876
rect 3842 842 3861 876
rect 3789 786 3861 842
rect 3789 752 3808 786
rect 3842 752 3861 786
rect 3789 696 3861 752
rect 3789 662 3808 696
rect 3842 662 3861 696
rect 3789 606 3861 662
rect 3789 572 3808 606
rect 3842 572 3861 606
rect 3789 516 3861 572
rect 3789 482 3808 516
rect 3842 482 3861 516
rect 3789 426 3861 482
rect 3789 392 3808 426
rect 3842 392 3861 426
rect 3789 336 3861 392
rect 2899 261 2971 321
rect 3789 302 3808 336
rect 3842 302 3861 336
rect 3789 261 3861 302
rect 2899 242 3861 261
rect 2899 208 2996 242
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 208 3861 242
rect 2899 189 3861 208
rect 4259 1132 5221 1151
rect 4259 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5221 1132
rect 4259 1079 5221 1098
rect 4259 1075 4331 1079
rect 4259 1041 4278 1075
rect 4312 1041 4331 1075
rect 4259 985 4331 1041
rect 5149 1056 5221 1079
rect 5149 1022 5168 1056
rect 5202 1022 5221 1056
rect 4259 951 4278 985
rect 4312 951 4331 985
rect 4259 895 4331 951
rect 4259 861 4278 895
rect 4312 861 4331 895
rect 4259 805 4331 861
rect 4259 771 4278 805
rect 4312 771 4331 805
rect 4259 715 4331 771
rect 4259 681 4278 715
rect 4312 681 4331 715
rect 4259 625 4331 681
rect 4259 591 4278 625
rect 4312 591 4331 625
rect 4259 535 4331 591
rect 4259 501 4278 535
rect 4312 501 4331 535
rect 4259 445 4331 501
rect 4259 411 4278 445
rect 4312 411 4331 445
rect 4259 355 4331 411
rect 4259 321 4278 355
rect 4312 321 4331 355
rect 5149 966 5221 1022
rect 5149 932 5168 966
rect 5202 932 5221 966
rect 5149 876 5221 932
rect 5149 842 5168 876
rect 5202 842 5221 876
rect 5149 786 5221 842
rect 5149 752 5168 786
rect 5202 752 5221 786
rect 5149 696 5221 752
rect 5149 662 5168 696
rect 5202 662 5221 696
rect 5149 606 5221 662
rect 5149 572 5168 606
rect 5202 572 5221 606
rect 5149 516 5221 572
rect 5149 482 5168 516
rect 5202 482 5221 516
rect 5149 426 5221 482
rect 5149 392 5168 426
rect 5202 392 5221 426
rect 5149 336 5221 392
rect 4259 261 4331 321
rect 5149 302 5168 336
rect 5202 302 5221 336
rect 5149 261 5221 302
rect 4259 242 5221 261
rect 4259 208 4356 242
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 208 5221 242
rect 4259 189 5221 208
rect 5619 1132 6581 1151
rect 5619 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 6581 1132
rect 5619 1079 6581 1098
rect 5619 1075 5691 1079
rect 5619 1041 5638 1075
rect 5672 1041 5691 1075
rect 5619 985 5691 1041
rect 6509 1056 6581 1079
rect 6509 1022 6528 1056
rect 6562 1022 6581 1056
rect 5619 951 5638 985
rect 5672 951 5691 985
rect 5619 895 5691 951
rect 5619 861 5638 895
rect 5672 861 5691 895
rect 5619 805 5691 861
rect 5619 771 5638 805
rect 5672 771 5691 805
rect 5619 715 5691 771
rect 5619 681 5638 715
rect 5672 681 5691 715
rect 5619 625 5691 681
rect 5619 591 5638 625
rect 5672 591 5691 625
rect 5619 535 5691 591
rect 5619 501 5638 535
rect 5672 501 5691 535
rect 5619 445 5691 501
rect 5619 411 5638 445
rect 5672 411 5691 445
rect 5619 355 5691 411
rect 5619 321 5638 355
rect 5672 321 5691 355
rect 6509 966 6581 1022
rect 6509 932 6528 966
rect 6562 932 6581 966
rect 6509 876 6581 932
rect 6509 842 6528 876
rect 6562 842 6581 876
rect 6509 786 6581 842
rect 6509 752 6528 786
rect 6562 752 6581 786
rect 6509 696 6581 752
rect 6509 662 6528 696
rect 6562 662 6581 696
rect 6509 606 6581 662
rect 6509 572 6528 606
rect 6562 572 6581 606
rect 6509 516 6581 572
rect 6509 482 6528 516
rect 6562 482 6581 516
rect 6509 426 6581 482
rect 6509 392 6528 426
rect 6562 392 6581 426
rect 6509 336 6581 392
rect 5619 261 5691 321
rect 6509 302 6528 336
rect 6562 302 6581 336
rect 6509 261 6581 302
rect 5619 242 6581 261
rect 5619 208 5716 242
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 208 6581 242
rect 5619 189 6581 208
rect 6979 1132 7941 1151
rect 6979 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 7941 1132
rect 6979 1079 7941 1098
rect 6979 1075 7051 1079
rect 6979 1041 6998 1075
rect 7032 1041 7051 1075
rect 6979 985 7051 1041
rect 7869 1056 7941 1079
rect 7869 1022 7888 1056
rect 7922 1022 7941 1056
rect 6979 951 6998 985
rect 7032 951 7051 985
rect 6979 895 7051 951
rect 6979 861 6998 895
rect 7032 861 7051 895
rect 6979 805 7051 861
rect 6979 771 6998 805
rect 7032 771 7051 805
rect 6979 715 7051 771
rect 6979 681 6998 715
rect 7032 681 7051 715
rect 6979 625 7051 681
rect 6979 591 6998 625
rect 7032 591 7051 625
rect 6979 535 7051 591
rect 6979 501 6998 535
rect 7032 501 7051 535
rect 6979 445 7051 501
rect 6979 411 6998 445
rect 7032 411 7051 445
rect 6979 355 7051 411
rect 6979 321 6998 355
rect 7032 321 7051 355
rect 7869 966 7941 1022
rect 7869 932 7888 966
rect 7922 932 7941 966
rect 7869 876 7941 932
rect 7869 842 7888 876
rect 7922 842 7941 876
rect 7869 786 7941 842
rect 7869 752 7888 786
rect 7922 752 7941 786
rect 7869 696 7941 752
rect 7869 662 7888 696
rect 7922 662 7941 696
rect 7869 606 7941 662
rect 7869 572 7888 606
rect 7922 572 7941 606
rect 7869 516 7941 572
rect 7869 482 7888 516
rect 7922 482 7941 516
rect 7869 426 7941 482
rect 7869 392 7888 426
rect 7922 392 7941 426
rect 7869 336 7941 392
rect 6979 261 7051 321
rect 7869 302 7888 336
rect 7922 302 7941 336
rect 7869 261 7941 302
rect 6979 242 7941 261
rect 6979 208 7076 242
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 208 7941 242
rect 6979 189 7941 208
rect 8339 1132 9301 1151
rect 8339 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9301 1132
rect 8339 1079 9301 1098
rect 8339 1075 8411 1079
rect 8339 1041 8358 1075
rect 8392 1041 8411 1075
rect 8339 985 8411 1041
rect 9229 1056 9301 1079
rect 9229 1022 9248 1056
rect 9282 1022 9301 1056
rect 8339 951 8358 985
rect 8392 951 8411 985
rect 8339 895 8411 951
rect 8339 861 8358 895
rect 8392 861 8411 895
rect 8339 805 8411 861
rect 8339 771 8358 805
rect 8392 771 8411 805
rect 8339 715 8411 771
rect 8339 681 8358 715
rect 8392 681 8411 715
rect 8339 625 8411 681
rect 8339 591 8358 625
rect 8392 591 8411 625
rect 8339 535 8411 591
rect 8339 501 8358 535
rect 8392 501 8411 535
rect 8339 445 8411 501
rect 8339 411 8358 445
rect 8392 411 8411 445
rect 8339 355 8411 411
rect 8339 321 8358 355
rect 8392 321 8411 355
rect 9229 966 9301 1022
rect 9229 932 9248 966
rect 9282 932 9301 966
rect 9229 876 9301 932
rect 9229 842 9248 876
rect 9282 842 9301 876
rect 9229 786 9301 842
rect 9229 752 9248 786
rect 9282 752 9301 786
rect 9229 696 9301 752
rect 9229 662 9248 696
rect 9282 662 9301 696
rect 9229 606 9301 662
rect 9229 572 9248 606
rect 9282 572 9301 606
rect 9229 516 9301 572
rect 9229 482 9248 516
rect 9282 482 9301 516
rect 9229 426 9301 482
rect 9229 392 9248 426
rect 9282 392 9301 426
rect 9229 336 9301 392
rect 8339 261 8411 321
rect 9229 302 9248 336
rect 9282 302 9301 336
rect 9229 261 9301 302
rect 8339 242 9301 261
rect 8339 208 8436 242
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 208 9301 242
rect 8339 189 9301 208
<< psubdiffcont >>
rect 5080 3250 5120 3290
rect 5080 3150 5120 3190
rect 6440 3250 6480 3290
rect 6440 3150 6480 3190
rect 7800 3250 7840 3290
rect 7800 3150 7840 3190
rect 4600 2700 4640 2740
rect 4600 2600 4640 2640
rect 4600 2500 4640 2540
rect 4600 2400 4640 2440
rect 4600 2300 4640 2340
rect 4600 2200 4640 2240
rect 4600 2100 4640 2140
rect 4600 2000 4640 2040
rect 8280 2700 8320 2740
rect 8280 2600 8320 2640
rect 8280 2500 8320 2540
rect 8280 2400 8320 2440
rect 8280 2300 8320 2340
rect 8280 2200 8320 2240
rect 8280 2100 8320 2140
rect 8280 2000 8320 2040
rect 7540 1640 7580 1680
rect 7540 1540 7580 1580
rect 1410 1222 1444 1256
rect 1506 1245 1540 1279
rect 1596 1245 1630 1279
rect 1686 1245 1720 1279
rect 1776 1245 1810 1279
rect 1866 1245 1900 1279
rect 1956 1245 1990 1279
rect 2046 1245 2080 1279
rect 2136 1245 2170 1279
rect 2226 1245 2260 1279
rect 2316 1245 2350 1279
rect 2406 1245 2440 1279
rect 2496 1245 2530 1279
rect 2597 1222 2631 1256
rect 1410 1132 1444 1166
rect 1410 1042 1444 1076
rect 1410 952 1444 986
rect 1410 862 1444 896
rect 1410 772 1444 806
rect 1410 682 1444 716
rect 1410 592 1444 626
rect 1410 502 1444 536
rect 1410 412 1444 446
rect 1410 322 1444 356
rect 1410 232 1444 266
rect 2597 1132 2631 1166
rect 2597 1042 2631 1076
rect 2597 952 2631 986
rect 2597 862 2631 896
rect 2597 772 2631 806
rect 2597 682 2631 716
rect 2597 592 2631 626
rect 2597 502 2631 536
rect 2597 412 2631 446
rect 2597 322 2631 356
rect 2597 232 2631 266
rect 1410 142 1444 176
rect 2597 142 2631 176
rect 1506 58 1540 92
rect 1596 58 1630 92
rect 1686 58 1720 92
rect 1776 58 1810 92
rect 1866 58 1900 92
rect 1956 58 1990 92
rect 2046 58 2080 92
rect 2136 58 2170 92
rect 2226 58 2260 92
rect 2316 58 2350 92
rect 2406 58 2440 92
rect 2496 58 2530 92
rect 2586 90 2620 92
rect 2600 58 2620 90
rect 2770 1222 2804 1256
rect 2866 1245 2900 1279
rect 2956 1245 2990 1279
rect 3046 1245 3080 1279
rect 3136 1245 3170 1279
rect 3226 1245 3260 1279
rect 3316 1245 3350 1279
rect 3406 1245 3440 1279
rect 3496 1245 3530 1279
rect 3586 1245 3620 1279
rect 3676 1245 3710 1279
rect 3766 1245 3800 1279
rect 3856 1245 3890 1279
rect 3957 1222 3991 1256
rect 2770 1132 2804 1166
rect 2770 1042 2804 1076
rect 2770 952 2804 986
rect 2770 862 2804 896
rect 2770 772 2804 806
rect 2770 682 2804 716
rect 2770 592 2804 626
rect 2770 502 2804 536
rect 2770 412 2804 446
rect 2770 322 2804 356
rect 2770 232 2804 266
rect 3957 1132 3991 1166
rect 3957 1042 3991 1076
rect 3957 952 3991 986
rect 3957 862 3991 896
rect 3957 772 3991 806
rect 3957 682 3991 716
rect 3957 592 3991 626
rect 3957 502 3991 536
rect 3957 412 3991 446
rect 3957 322 3991 356
rect 3957 232 3991 266
rect 2770 142 2804 176
rect 3957 142 3991 176
rect 4130 1222 4164 1256
rect 4226 1245 4260 1279
rect 4316 1245 4350 1279
rect 4406 1245 4440 1279
rect 4496 1245 4530 1279
rect 4586 1245 4620 1279
rect 4676 1245 4710 1279
rect 4766 1245 4800 1279
rect 4856 1245 4890 1279
rect 4946 1245 4980 1279
rect 5036 1245 5070 1279
rect 5126 1245 5160 1279
rect 5216 1245 5250 1279
rect 5317 1222 5351 1256
rect 4130 1132 4164 1166
rect 4130 1042 4164 1076
rect 4130 952 4164 986
rect 4130 862 4164 896
rect 4130 772 4164 806
rect 4130 682 4164 716
rect 4130 592 4164 626
rect 4130 502 4164 536
rect 4130 412 4164 446
rect 4130 322 4164 356
rect 4130 232 4164 266
rect 5317 1132 5351 1166
rect 5317 1042 5351 1076
rect 5317 952 5351 986
rect 5317 862 5351 896
rect 5317 772 5351 806
rect 5317 682 5351 716
rect 5317 592 5351 626
rect 5317 502 5351 536
rect 5317 412 5351 446
rect 5317 322 5351 356
rect 5317 232 5351 266
rect 4130 142 4164 176
rect 5317 142 5351 176
rect 5490 1222 5524 1256
rect 5586 1245 5620 1279
rect 5676 1245 5710 1279
rect 5766 1245 5800 1279
rect 5856 1245 5890 1279
rect 5946 1245 5980 1279
rect 6036 1245 6070 1279
rect 6126 1245 6160 1279
rect 6216 1245 6250 1279
rect 6306 1245 6340 1279
rect 6396 1245 6430 1279
rect 6486 1245 6520 1279
rect 6576 1245 6610 1279
rect 6677 1222 6711 1256
rect 5490 1132 5524 1166
rect 5490 1042 5524 1076
rect 5490 952 5524 986
rect 5490 862 5524 896
rect 5490 772 5524 806
rect 5490 682 5524 716
rect 5490 592 5524 626
rect 5490 502 5524 536
rect 5490 412 5524 446
rect 5490 322 5524 356
rect 5490 232 5524 266
rect 6677 1132 6711 1166
rect 6677 1042 6711 1076
rect 6677 952 6711 986
rect 6677 862 6711 896
rect 6677 772 6711 806
rect 6677 682 6711 716
rect 6677 592 6711 626
rect 6677 502 6711 536
rect 6677 412 6711 446
rect 6677 322 6711 356
rect 6677 232 6711 266
rect 5490 142 5524 176
rect 6677 142 6711 176
rect 6850 1222 6884 1256
rect 6946 1245 6980 1279
rect 7036 1245 7070 1279
rect 7126 1245 7160 1279
rect 7216 1245 7250 1279
rect 7306 1245 7340 1279
rect 7396 1245 7430 1279
rect 7486 1245 7520 1279
rect 7576 1245 7610 1279
rect 7666 1245 7700 1279
rect 7756 1245 7790 1279
rect 7846 1245 7880 1279
rect 7936 1245 7970 1279
rect 8037 1222 8071 1256
rect 6850 1132 6884 1166
rect 6850 1042 6884 1076
rect 6850 952 6884 986
rect 6850 862 6884 896
rect 6850 772 6884 806
rect 6850 682 6884 716
rect 6850 592 6884 626
rect 6850 502 6884 536
rect 6850 412 6884 446
rect 6850 322 6884 356
rect 6850 232 6884 266
rect 8037 1132 8071 1166
rect 8037 1042 8071 1076
rect 8037 952 8071 986
rect 8037 862 8071 896
rect 8037 772 8071 806
rect 8037 682 8071 716
rect 8037 592 8071 626
rect 8037 502 8071 536
rect 8037 412 8071 446
rect 8037 322 8071 356
rect 8037 232 8071 266
rect 6850 142 6884 176
rect 8037 142 8071 176
rect 8210 1222 8244 1256
rect 8306 1245 8340 1279
rect 8396 1245 8430 1279
rect 8486 1245 8520 1279
rect 8576 1245 8610 1279
rect 8666 1245 8700 1279
rect 8756 1245 8790 1279
rect 8846 1245 8880 1279
rect 8936 1245 8970 1279
rect 9026 1245 9060 1279
rect 9116 1245 9150 1279
rect 9206 1245 9240 1279
rect 9296 1245 9330 1279
rect 9397 1222 9431 1256
rect 8210 1132 8244 1166
rect 8210 1042 8244 1076
rect 8210 952 8244 986
rect 8210 862 8244 896
rect 8210 772 8244 806
rect 8210 682 8244 716
rect 8210 592 8244 626
rect 8210 502 8244 536
rect 8210 412 8244 446
rect 8210 322 8244 356
rect 8210 232 8244 266
rect 9397 1132 9431 1166
rect 9397 1042 9431 1076
rect 9397 952 9431 986
rect 9397 862 9431 896
rect 9397 772 9431 806
rect 9397 682 9431 716
rect 9397 592 9431 626
rect 9397 502 9431 536
rect 9397 412 9431 446
rect 9397 322 9431 356
rect 9397 232 9431 266
rect 8210 142 8244 176
rect 9397 142 9431 176
rect 2766 90 2800 92
rect 2780 58 2800 90
rect 2866 58 2900 92
rect 2946 90 2990 92
rect 2956 58 2990 90
rect 3046 58 3080 92
rect 3126 90 3170 92
rect 3136 58 3170 90
rect 3226 58 3260 92
rect 3306 90 3350 92
rect 3316 58 3350 90
rect 3406 58 3440 92
rect 3486 90 3530 92
rect 3496 58 3530 90
rect 3586 58 3620 92
rect 3666 90 3710 92
rect 3676 58 3710 90
rect 3766 58 3800 92
rect 3846 90 3890 92
rect 3856 58 3890 90
rect 3970 58 3980 92
rect 4026 90 4070 92
rect 4040 58 4070 90
rect 4150 58 4160 92
rect 4206 90 4260 92
rect 4220 58 4260 90
rect 4316 58 4350 92
rect 4386 90 4440 92
rect 4400 58 4440 90
rect 4496 58 4530 92
rect 4566 90 4620 92
rect 4580 58 4620 90
rect 4676 58 4710 92
rect 4746 90 4800 92
rect 4760 58 4800 90
rect 4856 58 4890 92
rect 4926 90 4980 92
rect 4940 58 4980 90
rect 5036 58 5070 92
rect 5106 90 5160 92
rect 5120 58 5160 90
rect 5216 58 5250 92
rect 5286 90 5330 92
rect 5300 58 5330 90
rect 5410 58 5430 92
rect 5466 90 5510 92
rect 5480 58 5510 90
rect 5586 58 5620 92
rect 5646 90 5710 92
rect 5660 58 5710 90
rect 5766 58 5800 92
rect 5826 90 5890 92
rect 5840 58 5890 90
rect 5946 58 5980 92
rect 6006 90 6070 92
rect 6020 58 6070 90
rect 6126 58 6160 92
rect 6186 90 6250 92
rect 6200 58 6250 90
rect 6306 58 6340 92
rect 6366 90 6430 92
rect 6380 58 6430 90
rect 6486 58 6520 92
rect 6546 90 6610 92
rect 6560 58 6610 90
rect 6670 58 6700 92
rect 6726 90 6770 92
rect 6740 58 6770 90
rect 6850 58 6880 92
rect 6906 90 6980 92
rect 6920 58 6980 90
rect 7030 58 7070 92
rect 7086 90 7160 92
rect 7100 58 7160 90
rect 7210 58 7250 92
rect 7266 90 7340 92
rect 7280 58 7340 90
rect 7390 58 7430 92
rect 7446 90 7520 92
rect 7460 58 7520 90
rect 7570 58 7610 92
rect 7626 90 7700 92
rect 7640 58 7700 90
rect 7750 58 7790 92
rect 7806 90 7880 92
rect 7820 58 7880 90
rect 7930 58 7970 92
rect 7986 90 8030 92
rect 8000 58 8030 90
rect 8110 90 8150 92
rect 8166 90 8210 92
rect 8110 58 8140 90
rect 8180 58 8210 90
rect 8290 58 8340 92
rect 8346 90 8390 92
rect 8360 58 8390 90
rect 8396 58 8430 92
rect 8470 58 8520 92
rect 8526 90 8570 92
rect 8540 58 8570 90
rect 8576 58 8610 92
rect 8650 58 8700 92
rect 8706 90 8750 92
rect 8720 58 8750 90
rect 8756 58 8790 92
rect 8830 58 8880 92
rect 8886 90 8930 92
rect 8900 58 8930 90
rect 8936 58 8970 92
rect 9010 58 9060 92
rect 9066 90 9110 92
rect 9080 58 9110 90
rect 9116 58 9150 92
rect 9190 58 9240 92
rect 9246 90 9290 92
rect 9260 58 9290 90
rect 9296 58 9330 92
rect 9370 90 9420 92
rect 9426 90 9470 92
rect 9370 58 9400 90
rect 9440 58 9470 90
<< nsubdiffcont >>
rect 4360 5370 4400 5410
rect 4360 5270 4400 5310
rect 4360 5170 4400 5210
rect 4360 5070 4400 5110
rect 4360 4970 4400 5010
rect 4360 4870 4400 4910
rect 4360 4770 4400 4810
rect 4360 4670 4400 4710
rect 8520 5370 8560 5410
rect 8520 5270 8560 5310
rect 8520 5170 8560 5210
rect 8520 5070 8560 5110
rect 8520 4970 8560 5010
rect 8520 4870 8560 4910
rect 8520 4770 8560 4810
rect 8520 4670 8560 4710
rect 4400 4060 4440 4100
rect 4400 3960 4440 4000
rect 4400 3860 4440 3900
rect 4400 3760 4440 3800
rect 5760 4060 5800 4100
rect 5760 3960 5800 4000
rect 5760 3860 5800 3900
rect 5760 3760 5800 3800
rect 7120 4060 7160 4100
rect 7120 3960 7160 4000
rect 7120 3860 7160 3900
rect 7120 3760 7160 3800
rect 8480 4060 8520 4100
rect 8480 3960 8520 4000
rect 8480 3860 8520 3900
rect 8480 3760 8520 3800
rect 9210 4060 9250 4100
rect 9210 3960 9250 4000
rect 9210 3860 9250 3900
rect 9210 3760 9250 3800
rect 1670 1098 1704 1132
rect 1760 1098 1794 1132
rect 1850 1098 1884 1132
rect 1940 1098 1974 1132
rect 2030 1098 2064 1132
rect 2120 1098 2154 1132
rect 2210 1098 2244 1132
rect 2300 1098 2334 1132
rect 2390 1098 2424 1132
rect 1558 1041 1592 1075
rect 2448 1022 2482 1056
rect 1558 951 1592 985
rect 1558 861 1592 895
rect 1558 771 1592 805
rect 1558 681 1592 715
rect 1558 591 1592 625
rect 1558 501 1592 535
rect 1558 411 1592 445
rect 1558 321 1592 355
rect 2448 932 2482 966
rect 2448 842 2482 876
rect 2448 752 2482 786
rect 2448 662 2482 696
rect 2448 572 2482 606
rect 2448 482 2482 516
rect 2448 392 2482 426
rect 2448 302 2482 336
rect 1636 208 1670 242
rect 1726 208 1760 242
rect 1816 208 1850 242
rect 1906 208 1940 242
rect 1996 208 2030 242
rect 2086 208 2120 242
rect 2176 208 2210 242
rect 2266 208 2300 242
rect 2356 208 2390 242
rect 3030 1098 3064 1132
rect 3120 1098 3154 1132
rect 3210 1098 3244 1132
rect 3300 1098 3334 1132
rect 3390 1098 3424 1132
rect 3480 1098 3514 1132
rect 3570 1098 3604 1132
rect 3660 1098 3694 1132
rect 3750 1098 3784 1132
rect 2918 1041 2952 1075
rect 3808 1022 3842 1056
rect 2918 951 2952 985
rect 2918 861 2952 895
rect 2918 771 2952 805
rect 2918 681 2952 715
rect 2918 591 2952 625
rect 2918 501 2952 535
rect 2918 411 2952 445
rect 2918 321 2952 355
rect 3808 932 3842 966
rect 3808 842 3842 876
rect 3808 752 3842 786
rect 3808 662 3842 696
rect 3808 572 3842 606
rect 3808 482 3842 516
rect 3808 392 3842 426
rect 3808 302 3842 336
rect 2996 208 3030 242
rect 3086 208 3120 242
rect 3176 208 3210 242
rect 3266 208 3300 242
rect 3356 208 3390 242
rect 3446 208 3480 242
rect 3536 208 3570 242
rect 3626 208 3660 242
rect 3716 208 3750 242
rect 4390 1098 4424 1132
rect 4480 1098 4514 1132
rect 4570 1098 4604 1132
rect 4660 1098 4694 1132
rect 4750 1098 4784 1132
rect 4840 1098 4874 1132
rect 4930 1098 4964 1132
rect 5020 1098 5054 1132
rect 5110 1098 5144 1132
rect 4278 1041 4312 1075
rect 5168 1022 5202 1056
rect 4278 951 4312 985
rect 4278 861 4312 895
rect 4278 771 4312 805
rect 4278 681 4312 715
rect 4278 591 4312 625
rect 4278 501 4312 535
rect 4278 411 4312 445
rect 4278 321 4312 355
rect 5168 932 5202 966
rect 5168 842 5202 876
rect 5168 752 5202 786
rect 5168 662 5202 696
rect 5168 572 5202 606
rect 5168 482 5202 516
rect 5168 392 5202 426
rect 5168 302 5202 336
rect 4356 208 4390 242
rect 4446 208 4480 242
rect 4536 208 4570 242
rect 4626 208 4660 242
rect 4716 208 4750 242
rect 4806 208 4840 242
rect 4896 208 4930 242
rect 4986 208 5020 242
rect 5076 208 5110 242
rect 5750 1098 5784 1132
rect 5840 1098 5874 1132
rect 5930 1098 5964 1132
rect 6020 1098 6054 1132
rect 6110 1098 6144 1132
rect 6200 1098 6234 1132
rect 6290 1098 6324 1132
rect 6380 1098 6414 1132
rect 6470 1098 6504 1132
rect 5638 1041 5672 1075
rect 6528 1022 6562 1056
rect 5638 951 5672 985
rect 5638 861 5672 895
rect 5638 771 5672 805
rect 5638 681 5672 715
rect 5638 591 5672 625
rect 5638 501 5672 535
rect 5638 411 5672 445
rect 5638 321 5672 355
rect 6528 932 6562 966
rect 6528 842 6562 876
rect 6528 752 6562 786
rect 6528 662 6562 696
rect 6528 572 6562 606
rect 6528 482 6562 516
rect 6528 392 6562 426
rect 6528 302 6562 336
rect 5716 208 5750 242
rect 5806 208 5840 242
rect 5896 208 5930 242
rect 5986 208 6020 242
rect 6076 208 6110 242
rect 6166 208 6200 242
rect 6256 208 6290 242
rect 6346 208 6380 242
rect 6436 208 6470 242
rect 7110 1098 7144 1132
rect 7200 1098 7234 1132
rect 7290 1098 7324 1132
rect 7380 1098 7414 1132
rect 7470 1098 7504 1132
rect 7560 1098 7594 1132
rect 7650 1098 7684 1132
rect 7740 1098 7774 1132
rect 7830 1098 7864 1132
rect 6998 1041 7032 1075
rect 7888 1022 7922 1056
rect 6998 951 7032 985
rect 6998 861 7032 895
rect 6998 771 7032 805
rect 6998 681 7032 715
rect 6998 591 7032 625
rect 6998 501 7032 535
rect 6998 411 7032 445
rect 6998 321 7032 355
rect 7888 932 7922 966
rect 7888 842 7922 876
rect 7888 752 7922 786
rect 7888 662 7922 696
rect 7888 572 7922 606
rect 7888 482 7922 516
rect 7888 392 7922 426
rect 7888 302 7922 336
rect 7076 208 7110 242
rect 7166 208 7200 242
rect 7256 208 7290 242
rect 7346 208 7380 242
rect 7436 208 7470 242
rect 7526 208 7560 242
rect 7616 208 7650 242
rect 7706 208 7740 242
rect 7796 208 7830 242
rect 8470 1098 8504 1132
rect 8560 1098 8594 1132
rect 8650 1098 8684 1132
rect 8740 1098 8774 1132
rect 8830 1098 8864 1132
rect 8920 1098 8954 1132
rect 9010 1098 9044 1132
rect 9100 1098 9134 1132
rect 9190 1098 9224 1132
rect 8358 1041 8392 1075
rect 9248 1022 9282 1056
rect 8358 951 8392 985
rect 8358 861 8392 895
rect 8358 771 8392 805
rect 8358 681 8392 715
rect 8358 591 8392 625
rect 8358 501 8392 535
rect 8358 411 8392 445
rect 8358 321 8392 355
rect 9248 932 9282 966
rect 9248 842 9282 876
rect 9248 752 9282 786
rect 9248 662 9282 696
rect 9248 572 9282 606
rect 9248 482 9282 516
rect 9248 392 9282 426
rect 9248 302 9282 336
rect 8436 208 8470 242
rect 8526 208 8560 242
rect 8616 208 8650 242
rect 8706 208 8740 242
rect 8796 208 8830 242
rect 8886 208 8920 242
rect 8976 208 9010 242
rect 9066 208 9100 242
rect 9156 208 9190 242
<< poly >>
rect 4500 5440 4620 5470
rect 4700 5440 4820 5470
rect 4900 5440 5020 5470
rect 5100 5440 5220 5470
rect 5300 5440 5420 5470
rect 5500 5440 5620 5470
rect 5700 5440 5820 5470
rect 5900 5440 6020 5470
rect 6100 5440 6220 5470
rect 6300 5440 6420 5470
rect 6500 5440 6620 5470
rect 6700 5440 6820 5470
rect 6900 5440 7020 5470
rect 7100 5440 7220 5470
rect 7300 5440 7420 5470
rect 7500 5440 7620 5470
rect 7700 5440 7820 5470
rect 7900 5440 8020 5470
rect 8100 5440 8220 5470
rect 8300 5440 8420 5470
rect 4500 4610 4620 4640
rect 4700 4620 4820 4640
rect 4900 4620 5020 4640
rect 5100 4620 5220 4640
rect 5300 4620 5420 4640
rect 5500 4620 5620 4640
rect 5700 4620 5820 4640
rect 5900 4620 6020 4640
rect 6100 4620 6220 4640
rect 6300 4620 6420 4640
rect 6500 4620 6620 4640
rect 6700 4620 6820 4640
rect 6900 4620 7020 4640
rect 7100 4620 7220 4640
rect 7300 4620 7420 4640
rect 7500 4620 7620 4640
rect 7700 4620 7820 4640
rect 7900 4620 8020 4640
rect 8100 4620 8220 4640
rect 4700 4590 8220 4620
rect 8300 4610 8420 4640
rect 6220 4550 6240 4590
rect 6280 4550 6300 4590
rect 6220 4530 6300 4550
rect 6620 4550 6640 4590
rect 6680 4550 6700 4590
rect 6620 4530 6700 4550
rect 8140 4550 8160 4590
rect 8200 4550 8220 4590
rect 8140 4530 8220 4550
rect 9030 4300 9110 4320
rect 9030 4260 9050 4300
rect 9090 4260 9110 4300
rect 9030 4240 9110 4260
rect 4540 4130 4660 4160
rect 4740 4130 4860 4160
rect 4940 4130 5060 4160
rect 5140 4130 5260 4160
rect 5340 4130 5460 4160
rect 5540 4130 5660 4160
rect 5900 4130 6020 4160
rect 6100 4130 6220 4160
rect 6300 4130 6420 4160
rect 6500 4130 6620 4160
rect 6700 4130 6820 4160
rect 6900 4130 7020 4160
rect 7260 4130 7380 4160
rect 7460 4130 7580 4160
rect 7660 4130 7780 4160
rect 7860 4130 7980 4160
rect 8060 4130 8180 4160
rect 8260 4130 8380 4160
rect 8830 4130 8860 4160
rect 9080 4130 9110 4240
rect 4540 3700 4660 3730
rect 4740 3710 4860 3730
rect 4940 3710 5060 3730
rect 5140 3710 5260 3730
rect 5340 3710 5460 3730
rect 4740 3680 5460 3710
rect 5540 3700 5660 3730
rect 5900 3700 6020 3730
rect 6100 3710 6220 3730
rect 6300 3710 6420 3730
rect 6500 3710 6620 3730
rect 6700 3710 6820 3730
rect 6100 3680 6820 3710
rect 6900 3700 7020 3730
rect 7260 3700 7380 3730
rect 7460 3710 7580 3730
rect 7660 3710 7780 3730
rect 7860 3710 7980 3730
rect 8060 3710 8180 3730
rect 7460 3680 8180 3710
rect 8260 3700 8380 3730
rect 5260 3640 5280 3680
rect 5320 3640 5340 3680
rect 5260 3620 5340 3640
rect 6140 3610 6180 3680
rect 6740 3610 6780 3680
rect 7580 3640 7600 3680
rect 7640 3640 7660 3680
rect 7580 3620 7660 3640
rect 8830 3650 8860 3730
rect 9080 3700 9110 3730
rect 8970 3650 9050 3670
rect 8830 3610 8990 3650
rect 9030 3610 9050 3650
rect 6120 3590 6200 3610
rect 6120 3550 6140 3590
rect 6180 3550 6200 3590
rect 6120 3530 6200 3550
rect 6720 3590 6800 3610
rect 8970 3590 9050 3610
rect 6720 3550 6740 3590
rect 6780 3550 6800 3590
rect 6720 3530 6800 3550
rect 6060 3410 6140 3430
rect 6060 3370 6080 3410
rect 6120 3370 6140 3410
rect 5220 3320 5340 3350
rect 5420 3320 5540 3350
rect 5620 3320 5740 3350
rect 5820 3340 6140 3370
rect 6780 3410 6860 3430
rect 6780 3370 6800 3410
rect 6840 3370 6860 3410
rect 5820 3320 5940 3340
rect 6020 3320 6140 3340
rect 6220 3320 6340 3350
rect 6580 3320 6700 3350
rect 6780 3340 7100 3370
rect 6780 3320 6900 3340
rect 6980 3320 7100 3340
rect 7180 3320 7300 3350
rect 7380 3320 7500 3350
rect 7580 3320 7700 3350
rect 5220 3090 5340 3120
rect 5420 3100 5540 3120
rect 5620 3100 5740 3120
rect 5420 3070 5740 3100
rect 5820 3090 5940 3120
rect 6020 3090 6140 3120
rect 6220 3090 6340 3120
rect 6580 3090 6700 3120
rect 6780 3090 6900 3120
rect 6980 3090 7100 3120
rect 7180 3100 7300 3120
rect 7380 3100 7500 3120
rect 7180 3070 7500 3100
rect 7580 3090 7700 3120
rect 5540 3030 5560 3070
rect 5600 3030 5620 3070
rect 5540 3010 5620 3030
rect 7300 3030 7320 3070
rect 7360 3030 7380 3070
rect 7300 3010 7380 3030
rect 5620 2860 6420 2880
rect 5620 2820 5640 2860
rect 5680 2820 5720 2860
rect 5760 2820 5800 2860
rect 5840 2820 5880 2860
rect 5920 2820 5960 2860
rect 6000 2820 6040 2860
rect 6080 2820 6120 2860
rect 6160 2820 6200 2860
rect 6240 2820 6280 2860
rect 6320 2820 6360 2860
rect 6400 2820 6420 2860
rect 4740 2770 5540 2800
rect 5620 2770 6420 2820
rect 6500 2860 7300 2880
rect 6500 2820 6520 2860
rect 6560 2820 6600 2860
rect 6640 2820 6680 2860
rect 6720 2820 6760 2860
rect 6800 2820 6840 2860
rect 6880 2820 6920 2860
rect 6960 2820 7000 2860
rect 7040 2820 7080 2860
rect 7120 2820 7160 2860
rect 7200 2820 7240 2860
rect 7280 2820 7300 2860
rect 6500 2770 7300 2820
rect 7380 2770 8180 2800
rect 4740 1940 5540 1970
rect 5620 1940 6420 1970
rect 6500 1940 7300 1970
rect 7380 1940 8180 1970
rect 5440 1800 5520 1820
rect 5440 1760 5460 1800
rect 5500 1760 5520 1800
rect 5440 1740 5520 1760
rect 5600 1800 5680 1820
rect 5600 1760 5620 1800
rect 5660 1760 5680 1800
rect 5600 1740 5680 1760
rect 5760 1800 5840 1820
rect 5760 1760 5780 1800
rect 5820 1760 5840 1800
rect 5760 1740 5840 1760
rect 5920 1800 6000 1820
rect 5920 1760 5940 1800
rect 5980 1760 6000 1800
rect 5920 1740 6000 1760
rect 6080 1800 6160 1820
rect 6080 1760 6100 1800
rect 6140 1760 6160 1800
rect 6080 1740 6160 1760
rect 6240 1800 6320 1820
rect 6240 1760 6260 1800
rect 6300 1760 6320 1800
rect 6240 1740 6320 1760
rect 6400 1800 6480 1820
rect 6400 1760 6420 1800
rect 6460 1760 6480 1800
rect 6400 1740 6480 1760
rect 6560 1800 6640 1820
rect 6560 1760 6580 1800
rect 6620 1760 6640 1800
rect 6560 1740 6640 1760
rect 6720 1800 6800 1820
rect 6720 1760 6740 1800
rect 6780 1760 6800 1800
rect 6720 1740 6800 1760
rect 6880 1800 6960 1820
rect 6880 1760 6900 1800
rect 6940 1760 6960 1800
rect 6880 1740 6960 1760
rect 7040 1800 7120 1820
rect 7040 1760 7060 1800
rect 7100 1760 7120 1800
rect 7040 1740 7120 1760
rect 7200 1800 7280 1820
rect 7200 1760 7220 1800
rect 7260 1760 7280 1800
rect 7200 1740 7280 1760
rect 7360 1800 7440 1820
rect 7360 1760 7380 1800
rect 7420 1760 7440 1800
rect 7360 1740 7440 1760
rect 5440 1710 7440 1740
rect 5440 1480 7440 1510
<< polycont >>
rect 6240 4550 6280 4590
rect 6640 4550 6680 4590
rect 8160 4550 8200 4590
rect 9050 4260 9090 4300
rect 5280 3640 5320 3680
rect 7600 3640 7640 3680
rect 8990 3610 9030 3650
rect 6140 3550 6180 3590
rect 6740 3550 6780 3590
rect 6080 3370 6120 3410
rect 6800 3370 6840 3410
rect 5560 3030 5600 3070
rect 7320 3030 7360 3070
rect 5640 2820 5680 2860
rect 5720 2820 5760 2860
rect 5800 2820 5840 2860
rect 5880 2820 5920 2860
rect 5960 2820 6000 2860
rect 6040 2820 6080 2860
rect 6120 2820 6160 2860
rect 6200 2820 6240 2860
rect 6280 2820 6320 2860
rect 6360 2820 6400 2860
rect 6520 2820 6560 2860
rect 6600 2820 6640 2860
rect 6680 2820 6720 2860
rect 6760 2820 6800 2860
rect 6840 2820 6880 2860
rect 6920 2820 6960 2860
rect 7000 2820 7040 2860
rect 7080 2820 7120 2860
rect 7160 2820 7200 2860
rect 7240 2820 7280 2860
rect 5460 1760 5500 1800
rect 5620 1760 5660 1800
rect 5780 1760 5820 1800
rect 5940 1760 5980 1800
rect 6100 1760 6140 1800
rect 6260 1760 6300 1800
rect 6420 1760 6460 1800
rect 6580 1760 6620 1800
rect 6740 1760 6780 1800
rect 6900 1760 6940 1800
rect 7060 1760 7100 1800
rect 7220 1760 7260 1800
rect 7380 1760 7420 1800
<< xpolycontact >>
rect 2010 4960 2450 5030
rect 3790 4960 4230 5030
rect 2010 4840 2450 4910
rect 3790 4840 4230 4910
rect 2010 4720 2450 4790
rect 3790 4720 4230 4790
rect 2010 4600 2450 4670
rect 3790 4600 4230 4670
rect 2010 4480 2450 4550
rect 3790 4480 4230 4550
rect 2010 3960 2450 4030
rect 3790 3960 4230 4030
rect 2010 3840 2450 3910
rect 3790 3840 4230 3910
rect 2010 3720 2450 3790
rect 3790 3720 4230 3790
rect 2010 3600 2450 3670
rect 3790 3600 4230 3670
rect 2010 3480 2450 3550
rect 3790 3480 4230 3550
rect 2010 3010 2450 3080
rect 3150 3010 3590 3080
rect 2010 2890 2450 2960
rect 3790 2890 4230 2960
rect 2010 2770 2450 2840
rect 3790 2770 4230 2840
rect 2010 2650 2450 2720
rect 3790 2650 4230 2720
rect 2010 2530 2450 2600
rect 3790 2530 4230 2600
rect 2010 2410 2450 2480
rect 3790 2410 4230 2480
<< xpolyres >>
rect 2450 4960 3790 5030
rect 2450 4840 3790 4910
rect 2450 4720 3790 4790
rect 2450 4600 3790 4670
rect 2450 4480 3790 4550
rect 2450 3960 3790 4030
rect 2450 3840 3790 3910
rect 2450 3720 3790 3790
rect 2450 3600 3790 3670
rect 2450 3480 3790 3550
rect 2450 3010 3150 3080
rect 2450 2890 3790 2960
rect 2450 2770 3790 2840
rect 2450 2650 3790 2720
rect 2450 2530 3790 2600
rect 2450 2410 3790 2480
<< locali >>
rect 4620 5530 4700 5550
rect 4620 5490 4640 5530
rect 4680 5490 4700 5530
rect 4620 5470 4700 5490
rect 5020 5530 5100 5550
rect 5020 5490 5040 5530
rect 5080 5490 5100 5530
rect 5020 5470 5100 5490
rect 5420 5530 5500 5550
rect 5420 5490 5440 5530
rect 5480 5490 5500 5530
rect 5420 5470 5500 5490
rect 5820 5530 5900 5550
rect 5820 5490 5840 5530
rect 5880 5490 5900 5530
rect 5820 5470 5900 5490
rect 6220 5530 6300 5550
rect 6220 5490 6240 5530
rect 6280 5490 6300 5530
rect 6220 5470 6300 5490
rect 6620 5530 6700 5550
rect 6620 5490 6640 5530
rect 6680 5490 6700 5530
rect 6620 5470 6700 5490
rect 7020 5530 7100 5550
rect 7020 5490 7040 5530
rect 7080 5490 7100 5530
rect 7020 5470 7100 5490
rect 7420 5530 7500 5550
rect 7420 5490 7440 5530
rect 7480 5490 7500 5530
rect 7420 5470 7500 5490
rect 7820 5530 7900 5550
rect 7820 5490 7840 5530
rect 7880 5490 7900 5530
rect 7820 5470 7900 5490
rect 8220 5530 8300 5550
rect 8220 5490 8240 5530
rect 8280 5490 8300 5530
rect 8220 5470 8300 5490
rect 4640 5430 4680 5470
rect 5040 5430 5080 5470
rect 5440 5430 5480 5470
rect 5840 5430 5880 5470
rect 6240 5430 6280 5470
rect 6640 5430 6680 5470
rect 7040 5430 7080 5470
rect 7440 5430 7480 5470
rect 7840 5430 7880 5470
rect 8240 5430 8280 5470
rect 4350 5410 4490 5430
rect 4350 5370 4360 5410
rect 4400 5370 4440 5410
rect 4480 5370 4490 5410
rect 4350 5310 4490 5370
rect 4350 5270 4360 5310
rect 4400 5270 4440 5310
rect 4480 5270 4490 5310
rect 4350 5210 4490 5270
rect 4350 5170 4360 5210
rect 4400 5170 4440 5210
rect 4480 5170 4490 5210
rect 4350 5110 4490 5170
rect 4350 5070 4360 5110
rect 4400 5070 4440 5110
rect 4480 5070 4490 5110
rect 1890 5010 2010 5030
rect 1890 4970 1910 5010
rect 1950 4970 2010 5010
rect 1890 4960 2010 4970
rect 1890 4950 1970 4960
rect 3790 4910 4230 4960
rect 4350 5010 4490 5070
rect 4350 4970 4360 5010
rect 4400 4970 4440 5010
rect 4480 4970 4490 5010
rect 4350 4910 4490 4970
rect 4350 4870 4360 4910
rect 4400 4870 4440 4910
rect 4480 4870 4490 4910
rect 2010 4790 2450 4840
rect 4350 4810 4490 4870
rect 3790 4670 4230 4720
rect 4350 4770 4360 4810
rect 4400 4770 4440 4810
rect 4480 4770 4490 4810
rect 4350 4710 4490 4770
rect 4350 4670 4360 4710
rect 4400 4670 4440 4710
rect 4480 4670 4490 4710
rect 4350 4650 4490 4670
rect 4630 5410 4690 5430
rect 4630 5370 4640 5410
rect 4680 5370 4690 5410
rect 4630 5310 4690 5370
rect 4630 5270 4640 5310
rect 4680 5270 4690 5310
rect 4630 5210 4690 5270
rect 4630 5170 4640 5210
rect 4680 5170 4690 5210
rect 4630 5110 4690 5170
rect 4630 5070 4640 5110
rect 4680 5070 4690 5110
rect 4630 5010 4690 5070
rect 4630 4970 4640 5010
rect 4680 4970 4690 5010
rect 4630 4910 4690 4970
rect 4630 4870 4640 4910
rect 4680 4870 4690 4910
rect 4630 4810 4690 4870
rect 4630 4770 4640 4810
rect 4680 4770 4690 4810
rect 4630 4710 4690 4770
rect 4630 4670 4640 4710
rect 4680 4670 4690 4710
rect 4630 4650 4690 4670
rect 4830 5410 4890 5430
rect 4830 5370 4840 5410
rect 4880 5370 4890 5410
rect 4830 5310 4890 5370
rect 4830 5270 4840 5310
rect 4880 5270 4890 5310
rect 4830 5210 4890 5270
rect 4830 5170 4840 5210
rect 4880 5170 4890 5210
rect 4830 5110 4890 5170
rect 4830 5070 4840 5110
rect 4880 5070 4890 5110
rect 4830 5010 4890 5070
rect 4830 4970 4840 5010
rect 4880 4970 4890 5010
rect 4830 4910 4890 4970
rect 4830 4870 4840 4910
rect 4880 4870 4890 4910
rect 4830 4810 4890 4870
rect 4830 4770 4840 4810
rect 4880 4770 4890 4810
rect 4830 4710 4890 4770
rect 4830 4670 4840 4710
rect 4880 4670 4890 4710
rect 4830 4650 4890 4670
rect 5030 5410 5090 5430
rect 5030 5370 5040 5410
rect 5080 5370 5090 5410
rect 5030 5310 5090 5370
rect 5030 5270 5040 5310
rect 5080 5270 5090 5310
rect 5030 5210 5090 5270
rect 5030 5170 5040 5210
rect 5080 5170 5090 5210
rect 5030 5110 5090 5170
rect 5030 5070 5040 5110
rect 5080 5070 5090 5110
rect 5030 5010 5090 5070
rect 5030 4970 5040 5010
rect 5080 4970 5090 5010
rect 5030 4910 5090 4970
rect 5030 4870 5040 4910
rect 5080 4870 5090 4910
rect 5030 4810 5090 4870
rect 5030 4770 5040 4810
rect 5080 4770 5090 4810
rect 5030 4710 5090 4770
rect 5030 4670 5040 4710
rect 5080 4670 5090 4710
rect 5030 4650 5090 4670
rect 5230 5410 5290 5430
rect 5230 5370 5240 5410
rect 5280 5370 5290 5410
rect 5230 5310 5290 5370
rect 5230 5270 5240 5310
rect 5280 5270 5290 5310
rect 5230 5210 5290 5270
rect 5230 5170 5240 5210
rect 5280 5170 5290 5210
rect 5230 5110 5290 5170
rect 5230 5070 5240 5110
rect 5280 5070 5290 5110
rect 5230 5010 5290 5070
rect 5230 4970 5240 5010
rect 5280 4970 5290 5010
rect 5230 4910 5290 4970
rect 5230 4870 5240 4910
rect 5280 4870 5290 4910
rect 5230 4810 5290 4870
rect 5230 4770 5240 4810
rect 5280 4770 5290 4810
rect 5230 4710 5290 4770
rect 5230 4670 5240 4710
rect 5280 4670 5290 4710
rect 5230 4650 5290 4670
rect 5430 5410 5490 5430
rect 5430 5370 5440 5410
rect 5480 5370 5490 5410
rect 5430 5310 5490 5370
rect 5430 5270 5440 5310
rect 5480 5270 5490 5310
rect 5430 5210 5490 5270
rect 5430 5170 5440 5210
rect 5480 5170 5490 5210
rect 5430 5110 5490 5170
rect 5430 5070 5440 5110
rect 5480 5070 5490 5110
rect 5430 5010 5490 5070
rect 5430 4970 5440 5010
rect 5480 4970 5490 5010
rect 5430 4910 5490 4970
rect 5430 4870 5440 4910
rect 5480 4870 5490 4910
rect 5430 4810 5490 4870
rect 5430 4770 5440 4810
rect 5480 4770 5490 4810
rect 5430 4710 5490 4770
rect 5430 4670 5440 4710
rect 5480 4670 5490 4710
rect 5430 4650 5490 4670
rect 5630 5410 5690 5430
rect 5630 5370 5640 5410
rect 5680 5370 5690 5410
rect 5630 5310 5690 5370
rect 5630 5270 5640 5310
rect 5680 5270 5690 5310
rect 5630 5210 5690 5270
rect 5630 5170 5640 5210
rect 5680 5170 5690 5210
rect 5630 5110 5690 5170
rect 5630 5070 5640 5110
rect 5680 5070 5690 5110
rect 5630 5010 5690 5070
rect 5630 4970 5640 5010
rect 5680 4970 5690 5010
rect 5630 4910 5690 4970
rect 5630 4870 5640 4910
rect 5680 4870 5690 4910
rect 5630 4810 5690 4870
rect 5630 4770 5640 4810
rect 5680 4770 5690 4810
rect 5630 4710 5690 4770
rect 5630 4670 5640 4710
rect 5680 4670 5690 4710
rect 5630 4650 5690 4670
rect 5830 5410 5890 5430
rect 5830 5370 5840 5410
rect 5880 5370 5890 5410
rect 5830 5310 5890 5370
rect 5830 5270 5840 5310
rect 5880 5270 5890 5310
rect 5830 5210 5890 5270
rect 5830 5170 5840 5210
rect 5880 5170 5890 5210
rect 5830 5110 5890 5170
rect 5830 5070 5840 5110
rect 5880 5070 5890 5110
rect 5830 5010 5890 5070
rect 5830 4970 5840 5010
rect 5880 4970 5890 5010
rect 5830 4910 5890 4970
rect 5830 4870 5840 4910
rect 5880 4870 5890 4910
rect 5830 4810 5890 4870
rect 5830 4770 5840 4810
rect 5880 4770 5890 4810
rect 5830 4710 5890 4770
rect 5830 4670 5840 4710
rect 5880 4670 5890 4710
rect 5830 4650 5890 4670
rect 6030 5410 6090 5430
rect 6030 5370 6040 5410
rect 6080 5370 6090 5410
rect 6030 5310 6090 5370
rect 6030 5270 6040 5310
rect 6080 5270 6090 5310
rect 6030 5210 6090 5270
rect 6030 5170 6040 5210
rect 6080 5170 6090 5210
rect 6030 5110 6090 5170
rect 6030 5070 6040 5110
rect 6080 5070 6090 5110
rect 6030 5010 6090 5070
rect 6030 4970 6040 5010
rect 6080 4970 6090 5010
rect 6030 4910 6090 4970
rect 6030 4870 6040 4910
rect 6080 4870 6090 4910
rect 6030 4810 6090 4870
rect 6030 4770 6040 4810
rect 6080 4770 6090 4810
rect 6030 4710 6090 4770
rect 6030 4670 6040 4710
rect 6080 4670 6090 4710
rect 6030 4650 6090 4670
rect 6230 5410 6290 5430
rect 6230 5370 6240 5410
rect 6280 5370 6290 5410
rect 6230 5310 6290 5370
rect 6230 5270 6240 5310
rect 6280 5270 6290 5310
rect 6230 5210 6290 5270
rect 6230 5170 6240 5210
rect 6280 5170 6290 5210
rect 6230 5110 6290 5170
rect 6230 5070 6240 5110
rect 6280 5070 6290 5110
rect 6230 5010 6290 5070
rect 6230 4970 6240 5010
rect 6280 4970 6290 5010
rect 6230 4910 6290 4970
rect 6230 4870 6240 4910
rect 6280 4870 6290 4910
rect 6230 4810 6290 4870
rect 6230 4770 6240 4810
rect 6280 4770 6290 4810
rect 6230 4710 6290 4770
rect 6230 4670 6240 4710
rect 6280 4670 6290 4710
rect 6230 4650 6290 4670
rect 6430 5410 6490 5430
rect 6430 5370 6440 5410
rect 6480 5370 6490 5410
rect 6430 5310 6490 5370
rect 6430 5270 6440 5310
rect 6480 5270 6490 5310
rect 6430 5210 6490 5270
rect 6430 5170 6440 5210
rect 6480 5170 6490 5210
rect 6430 5110 6490 5170
rect 6430 5070 6440 5110
rect 6480 5070 6490 5110
rect 6430 5010 6490 5070
rect 6430 4970 6440 5010
rect 6480 4970 6490 5010
rect 6430 4910 6490 4970
rect 6430 4870 6440 4910
rect 6480 4870 6490 4910
rect 6430 4810 6490 4870
rect 6430 4770 6440 4810
rect 6480 4770 6490 4810
rect 6430 4710 6490 4770
rect 6430 4670 6440 4710
rect 6480 4670 6490 4710
rect 6430 4650 6490 4670
rect 6630 5410 6690 5430
rect 6630 5370 6640 5410
rect 6680 5370 6690 5410
rect 6630 5310 6690 5370
rect 6630 5270 6640 5310
rect 6680 5270 6690 5310
rect 6630 5210 6690 5270
rect 6630 5170 6640 5210
rect 6680 5170 6690 5210
rect 6630 5110 6690 5170
rect 6630 5070 6640 5110
rect 6680 5070 6690 5110
rect 6630 5010 6690 5070
rect 6630 4970 6640 5010
rect 6680 4970 6690 5010
rect 6630 4910 6690 4970
rect 6630 4870 6640 4910
rect 6680 4870 6690 4910
rect 6630 4810 6690 4870
rect 6630 4770 6640 4810
rect 6680 4770 6690 4810
rect 6630 4710 6690 4770
rect 6630 4670 6640 4710
rect 6680 4670 6690 4710
rect 6630 4650 6690 4670
rect 6830 5410 6890 5430
rect 6830 5370 6840 5410
rect 6880 5370 6890 5410
rect 6830 5310 6890 5370
rect 6830 5270 6840 5310
rect 6880 5270 6890 5310
rect 6830 5210 6890 5270
rect 6830 5170 6840 5210
rect 6880 5170 6890 5210
rect 6830 5110 6890 5170
rect 6830 5070 6840 5110
rect 6880 5070 6890 5110
rect 6830 5010 6890 5070
rect 6830 4970 6840 5010
rect 6880 4970 6890 5010
rect 6830 4910 6890 4970
rect 6830 4870 6840 4910
rect 6880 4870 6890 4910
rect 6830 4810 6890 4870
rect 6830 4770 6840 4810
rect 6880 4770 6890 4810
rect 6830 4710 6890 4770
rect 6830 4670 6840 4710
rect 6880 4670 6890 4710
rect 6830 4650 6890 4670
rect 7030 5410 7090 5430
rect 7030 5370 7040 5410
rect 7080 5370 7090 5410
rect 7030 5310 7090 5370
rect 7030 5270 7040 5310
rect 7080 5270 7090 5310
rect 7030 5210 7090 5270
rect 7030 5170 7040 5210
rect 7080 5170 7090 5210
rect 7030 5110 7090 5170
rect 7030 5070 7040 5110
rect 7080 5070 7090 5110
rect 7030 5010 7090 5070
rect 7030 4970 7040 5010
rect 7080 4970 7090 5010
rect 7030 4910 7090 4970
rect 7030 4870 7040 4910
rect 7080 4870 7090 4910
rect 7030 4810 7090 4870
rect 7030 4770 7040 4810
rect 7080 4770 7090 4810
rect 7030 4710 7090 4770
rect 7030 4670 7040 4710
rect 7080 4670 7090 4710
rect 7030 4650 7090 4670
rect 7230 5410 7290 5430
rect 7230 5370 7240 5410
rect 7280 5370 7290 5410
rect 7230 5310 7290 5370
rect 7230 5270 7240 5310
rect 7280 5270 7290 5310
rect 7230 5210 7290 5270
rect 7230 5170 7240 5210
rect 7280 5170 7290 5210
rect 7230 5110 7290 5170
rect 7230 5070 7240 5110
rect 7280 5070 7290 5110
rect 7230 5010 7290 5070
rect 7230 4970 7240 5010
rect 7280 4970 7290 5010
rect 7230 4910 7290 4970
rect 7230 4870 7240 4910
rect 7280 4870 7290 4910
rect 7230 4810 7290 4870
rect 7230 4770 7240 4810
rect 7280 4770 7290 4810
rect 7230 4710 7290 4770
rect 7230 4670 7240 4710
rect 7280 4670 7290 4710
rect 7230 4650 7290 4670
rect 7430 5410 7490 5430
rect 7430 5370 7440 5410
rect 7480 5370 7490 5410
rect 7430 5310 7490 5370
rect 7430 5270 7440 5310
rect 7480 5270 7490 5310
rect 7430 5210 7490 5270
rect 7430 5170 7440 5210
rect 7480 5170 7490 5210
rect 7430 5110 7490 5170
rect 7430 5070 7440 5110
rect 7480 5070 7490 5110
rect 7430 5010 7490 5070
rect 7430 4970 7440 5010
rect 7480 4970 7490 5010
rect 7430 4910 7490 4970
rect 7430 4870 7440 4910
rect 7480 4870 7490 4910
rect 7430 4810 7490 4870
rect 7430 4770 7440 4810
rect 7480 4770 7490 4810
rect 7430 4710 7490 4770
rect 7430 4670 7440 4710
rect 7480 4670 7490 4710
rect 7430 4650 7490 4670
rect 7630 5410 7690 5430
rect 7630 5370 7640 5410
rect 7680 5370 7690 5410
rect 7630 5310 7690 5370
rect 7630 5270 7640 5310
rect 7680 5270 7690 5310
rect 7630 5210 7690 5270
rect 7630 5170 7640 5210
rect 7680 5170 7690 5210
rect 7630 5110 7690 5170
rect 7630 5070 7640 5110
rect 7680 5070 7690 5110
rect 7630 5010 7690 5070
rect 7630 4970 7640 5010
rect 7680 4970 7690 5010
rect 7630 4910 7690 4970
rect 7630 4870 7640 4910
rect 7680 4870 7690 4910
rect 7630 4810 7690 4870
rect 7630 4770 7640 4810
rect 7680 4770 7690 4810
rect 7630 4710 7690 4770
rect 7630 4670 7640 4710
rect 7680 4670 7690 4710
rect 7630 4650 7690 4670
rect 7830 5410 7890 5430
rect 7830 5370 7840 5410
rect 7880 5370 7890 5410
rect 7830 5310 7890 5370
rect 7830 5270 7840 5310
rect 7880 5270 7890 5310
rect 7830 5210 7890 5270
rect 7830 5170 7840 5210
rect 7880 5170 7890 5210
rect 7830 5110 7890 5170
rect 7830 5070 7840 5110
rect 7880 5070 7890 5110
rect 7830 5010 7890 5070
rect 7830 4970 7840 5010
rect 7880 4970 7890 5010
rect 7830 4910 7890 4970
rect 7830 4870 7840 4910
rect 7880 4870 7890 4910
rect 7830 4810 7890 4870
rect 7830 4770 7840 4810
rect 7880 4770 7890 4810
rect 7830 4710 7890 4770
rect 7830 4670 7840 4710
rect 7880 4670 7890 4710
rect 7830 4650 7890 4670
rect 8030 5410 8090 5430
rect 8030 5370 8040 5410
rect 8080 5370 8090 5410
rect 8030 5310 8090 5370
rect 8030 5270 8040 5310
rect 8080 5270 8090 5310
rect 8030 5210 8090 5270
rect 8030 5170 8040 5210
rect 8080 5170 8090 5210
rect 8030 5110 8090 5170
rect 8030 5070 8040 5110
rect 8080 5070 8090 5110
rect 8030 5010 8090 5070
rect 8030 4970 8040 5010
rect 8080 4970 8090 5010
rect 8030 4910 8090 4970
rect 8030 4870 8040 4910
rect 8080 4870 8090 4910
rect 8030 4810 8090 4870
rect 8030 4770 8040 4810
rect 8080 4770 8090 4810
rect 8030 4710 8090 4770
rect 8030 4670 8040 4710
rect 8080 4670 8090 4710
rect 8030 4650 8090 4670
rect 8230 5410 8290 5430
rect 8230 5370 8240 5410
rect 8280 5370 8290 5410
rect 8230 5310 8290 5370
rect 8230 5270 8240 5310
rect 8280 5270 8290 5310
rect 8230 5210 8290 5270
rect 8230 5170 8240 5210
rect 8280 5170 8290 5210
rect 8230 5110 8290 5170
rect 8230 5070 8240 5110
rect 8280 5070 8290 5110
rect 8230 5010 8290 5070
rect 8230 4970 8240 5010
rect 8280 4970 8290 5010
rect 8230 4910 8290 4970
rect 8230 4870 8240 4910
rect 8280 4870 8290 4910
rect 8230 4810 8290 4870
rect 8230 4770 8240 4810
rect 8280 4770 8290 4810
rect 8230 4710 8290 4770
rect 8230 4670 8240 4710
rect 8280 4670 8290 4710
rect 8230 4650 8290 4670
rect 8430 5410 8570 5430
rect 8430 5370 8440 5410
rect 8480 5370 8520 5410
rect 8560 5370 8570 5410
rect 8430 5310 8570 5370
rect 8430 5270 8440 5310
rect 8480 5270 8520 5310
rect 8560 5270 8570 5310
rect 8430 5210 8570 5270
rect 8430 5170 8440 5210
rect 8480 5170 8520 5210
rect 8560 5170 8570 5210
rect 8430 5110 8570 5170
rect 8430 5070 8440 5110
rect 8480 5070 8520 5110
rect 8560 5070 8570 5110
rect 8430 5010 8570 5070
rect 8430 4970 8440 5010
rect 8480 4970 8520 5010
rect 8560 4970 8570 5010
rect 8430 4910 8570 4970
rect 8430 4870 8440 4910
rect 8480 4870 8520 4910
rect 8560 4870 8570 4910
rect 8430 4810 8570 4870
rect 8430 4770 8440 4810
rect 8480 4770 8520 4810
rect 8560 4770 8570 4810
rect 8430 4710 8570 4770
rect 8430 4670 8440 4710
rect 8480 4670 8520 4710
rect 8560 4670 8570 4710
rect 8430 4650 8570 4670
rect 4840 4610 4880 4650
rect 2010 4550 2450 4600
rect 4820 4590 4900 4610
rect 4820 4550 4840 4590
rect 4880 4550 4900 4590
rect 4820 4530 4900 4550
rect 5240 4520 5280 4650
rect 3790 4420 4230 4480
rect 5220 4500 5300 4520
rect 5220 4460 5240 4500
rect 5280 4460 5300 4500
rect 5220 4440 5300 4460
rect 5640 4430 5680 4650
rect 6040 4520 6080 4650
rect 6220 4590 6300 4610
rect 6220 4550 6240 4590
rect 6280 4550 6300 4590
rect 6220 4530 6300 4550
rect 6020 4500 6100 4520
rect 6020 4460 6040 4500
rect 6080 4460 6100 4500
rect 6020 4440 6100 4460
rect 6440 4430 6480 4650
rect 6840 4610 6880 4650
rect 6620 4590 6700 4610
rect 6620 4550 6640 4590
rect 6680 4550 6700 4590
rect 6620 4530 6700 4550
rect 6820 4590 6900 4610
rect 6820 4550 6840 4590
rect 6880 4550 6900 4590
rect 6820 4530 6900 4550
rect 7240 4430 7280 4650
rect 7640 4610 7680 4650
rect 7620 4590 7700 4610
rect 7620 4550 7640 4590
rect 7680 4550 7700 4590
rect 7620 4530 7700 4550
rect 8040 4520 8080 4650
rect 8140 4590 8220 4610
rect 8140 4550 8160 4590
rect 8200 4550 8220 4590
rect 8140 4530 8220 4550
rect 8020 4500 8100 4520
rect 8020 4460 8040 4500
rect 8080 4460 8100 4500
rect 8020 4440 8100 4460
rect 3790 4380 3810 4420
rect 3850 4380 3900 4420
rect 3940 4380 3990 4420
rect 4030 4380 4080 4420
rect 4120 4380 4170 4420
rect 4210 4380 4230 4420
rect 3790 4360 4230 4380
rect 5620 4410 5700 4430
rect 5620 4370 5640 4410
rect 5680 4370 5700 4410
rect 5620 4350 5700 4370
rect 6420 4410 6500 4430
rect 6420 4370 6440 4410
rect 6480 4370 6500 4410
rect 6420 4350 6500 4370
rect 7220 4410 7300 4430
rect 7220 4370 7240 4410
rect 7280 4370 7300 4410
rect 7220 4350 7300 4370
rect 8750 4320 8830 4340
rect 8750 4280 8770 4320
rect 8810 4300 9110 4320
rect 8810 4280 9050 4300
rect 8750 4260 8830 4280
rect 9030 4260 9050 4280
rect 9090 4260 9110 4300
rect 4460 4220 4540 4240
rect 4460 4180 4480 4220
rect 4520 4180 4540 4220
rect 4460 4160 4540 4180
rect 4660 4220 4740 4240
rect 4660 4180 4680 4220
rect 4720 4180 4740 4220
rect 4660 4160 4740 4180
rect 5060 4220 5140 4240
rect 5060 4180 5080 4220
rect 5120 4180 5140 4220
rect 5060 4160 5140 4180
rect 5460 4220 5540 4240
rect 5460 4180 5480 4220
rect 5520 4180 5540 4220
rect 5460 4160 5540 4180
rect 5660 4220 5740 4240
rect 5660 4180 5680 4220
rect 5720 4180 5740 4220
rect 5660 4160 5740 4180
rect 5820 4220 5900 4240
rect 5820 4180 5840 4220
rect 5880 4180 5900 4220
rect 5820 4160 5900 4180
rect 6020 4220 6100 4240
rect 6020 4180 6040 4220
rect 6080 4180 6100 4220
rect 6020 4160 6100 4180
rect 6220 4220 6300 4240
rect 6220 4180 6240 4220
rect 6280 4180 6300 4220
rect 6220 4160 6300 4180
rect 6420 4220 6500 4240
rect 6420 4180 6440 4220
rect 6480 4180 6500 4220
rect 6420 4160 6500 4180
rect 6620 4220 6700 4240
rect 6620 4180 6640 4220
rect 6680 4180 6700 4220
rect 6620 4160 6700 4180
rect 6820 4220 6900 4240
rect 6820 4180 6840 4220
rect 6880 4180 6900 4220
rect 6820 4160 6900 4180
rect 7020 4220 7100 4240
rect 7020 4180 7040 4220
rect 7080 4180 7100 4220
rect 7020 4160 7100 4180
rect 7180 4220 7260 4240
rect 7180 4180 7200 4220
rect 7240 4180 7260 4220
rect 7180 4160 7260 4180
rect 7380 4220 7460 4240
rect 7380 4180 7400 4220
rect 7440 4180 7460 4220
rect 7380 4160 7460 4180
rect 7780 4220 7860 4240
rect 7780 4180 7800 4220
rect 7840 4180 7860 4220
rect 7780 4160 7860 4180
rect 8180 4220 8260 4240
rect 8180 4180 8200 4220
rect 8240 4180 8260 4220
rect 8180 4160 8260 4180
rect 8380 4220 8460 4240
rect 8380 4180 8400 4220
rect 8440 4180 8460 4220
rect 8380 4160 8460 4180
rect 4480 4120 4520 4160
rect 4680 4120 4720 4160
rect 5080 4120 5120 4160
rect 5480 4120 5520 4160
rect 5680 4120 5720 4160
rect 5840 4120 5880 4160
rect 6040 4120 6080 4160
rect 6240 4120 6280 4160
rect 6440 4120 6480 4160
rect 6640 4120 6680 4160
rect 6840 4120 6880 4160
rect 7040 4120 7080 4160
rect 7200 4120 7240 4160
rect 7400 4120 7440 4160
rect 7800 4120 7840 4160
rect 8200 4120 8240 4160
rect 8400 4120 8440 4160
rect 8770 4120 8810 4260
rect 9030 4240 9110 4260
rect 9150 4220 9230 4240
rect 9150 4180 9170 4220
rect 9210 4180 9230 4220
rect 9150 4160 9230 4180
rect 9170 4120 9210 4160
rect 4390 4100 4530 4120
rect 4390 4060 4400 4100
rect 4440 4060 4480 4100
rect 4520 4060 4530 4100
rect 1890 4010 2010 4030
rect 1890 3970 1910 4010
rect 1950 3970 2010 4010
rect 1890 3960 2010 3970
rect 1890 3950 1970 3960
rect 3790 3910 4230 3960
rect 4390 4000 4530 4060
rect 4390 3960 4400 4000
rect 4440 3960 4480 4000
rect 4520 3960 4530 4000
rect 4390 3900 4530 3960
rect 4390 3860 4400 3900
rect 4440 3860 4480 3900
rect 4520 3860 4530 3900
rect 2010 3790 2450 3840
rect 4390 3800 4530 3860
rect 4390 3760 4400 3800
rect 4440 3760 4480 3800
rect 4520 3760 4530 3800
rect 4390 3740 4530 3760
rect 4670 4100 4730 4120
rect 4670 4060 4680 4100
rect 4720 4060 4730 4100
rect 4670 4000 4730 4060
rect 4670 3960 4680 4000
rect 4720 3960 4730 4000
rect 4670 3900 4730 3960
rect 4670 3860 4680 3900
rect 4720 3860 4730 3900
rect 4670 3800 4730 3860
rect 4670 3760 4680 3800
rect 4720 3760 4730 3800
rect 4670 3740 4730 3760
rect 4870 4100 4930 4120
rect 4870 4060 4880 4100
rect 4920 4060 4930 4100
rect 4870 4000 4930 4060
rect 4870 3960 4880 4000
rect 4920 3960 4930 4000
rect 4870 3900 4930 3960
rect 4870 3860 4880 3900
rect 4920 3860 4930 3900
rect 4870 3800 4930 3860
rect 4870 3760 4880 3800
rect 4920 3760 4930 3800
rect 4870 3740 4930 3760
rect 5070 4100 5130 4120
rect 5070 4060 5080 4100
rect 5120 4060 5130 4100
rect 5070 4000 5130 4060
rect 5070 3960 5080 4000
rect 5120 3960 5130 4000
rect 5070 3900 5130 3960
rect 5070 3860 5080 3900
rect 5120 3860 5130 3900
rect 5070 3800 5130 3860
rect 5070 3760 5080 3800
rect 5120 3760 5130 3800
rect 5070 3740 5130 3760
rect 5270 4100 5330 4120
rect 5270 4060 5280 4100
rect 5320 4060 5330 4100
rect 5270 4000 5330 4060
rect 5270 3960 5280 4000
rect 5320 3960 5330 4000
rect 5270 3900 5330 3960
rect 5270 3860 5280 3900
rect 5320 3860 5330 3900
rect 5270 3800 5330 3860
rect 5270 3760 5280 3800
rect 5320 3760 5330 3800
rect 5270 3740 5330 3760
rect 5470 4100 5530 4120
rect 5470 4060 5480 4100
rect 5520 4060 5530 4100
rect 5470 4000 5530 4060
rect 5470 3960 5480 4000
rect 5520 3960 5530 4000
rect 5470 3900 5530 3960
rect 5470 3860 5480 3900
rect 5520 3860 5530 3900
rect 5470 3800 5530 3860
rect 5470 3760 5480 3800
rect 5520 3760 5530 3800
rect 5470 3740 5530 3760
rect 5670 4100 5890 4120
rect 5670 4060 5680 4100
rect 5720 4060 5760 4100
rect 5800 4060 5840 4100
rect 5880 4060 5890 4100
rect 5670 4000 5890 4060
rect 5670 3960 5680 4000
rect 5720 3960 5760 4000
rect 5800 3960 5840 4000
rect 5880 3960 5890 4000
rect 5670 3900 5890 3960
rect 5670 3860 5680 3900
rect 5720 3860 5760 3900
rect 5800 3860 5840 3900
rect 5880 3860 5890 3900
rect 5670 3800 5890 3860
rect 5670 3760 5680 3800
rect 5720 3760 5760 3800
rect 5800 3760 5840 3800
rect 5880 3760 5890 3800
rect 5670 3740 5890 3760
rect 6030 4100 6090 4120
rect 6030 4060 6040 4100
rect 6080 4060 6090 4100
rect 6030 4000 6090 4060
rect 6030 3960 6040 4000
rect 6080 3960 6090 4000
rect 6030 3900 6090 3960
rect 6030 3860 6040 3900
rect 6080 3860 6090 3900
rect 6030 3800 6090 3860
rect 6030 3760 6040 3800
rect 6080 3760 6090 3800
rect 6030 3740 6090 3760
rect 6230 4100 6290 4120
rect 6230 4060 6240 4100
rect 6280 4060 6290 4100
rect 6230 4000 6290 4060
rect 6230 3960 6240 4000
rect 6280 3960 6290 4000
rect 6230 3900 6290 3960
rect 6230 3860 6240 3900
rect 6280 3860 6290 3900
rect 6230 3800 6290 3860
rect 6230 3760 6240 3800
rect 6280 3760 6290 3800
rect 6230 3740 6290 3760
rect 6430 4100 6490 4120
rect 6430 4060 6440 4100
rect 6480 4060 6490 4100
rect 6430 4000 6490 4060
rect 6430 3960 6440 4000
rect 6480 3960 6490 4000
rect 6430 3900 6490 3960
rect 6430 3860 6440 3900
rect 6480 3860 6490 3900
rect 6430 3800 6490 3860
rect 6430 3760 6440 3800
rect 6480 3760 6490 3800
rect 6430 3740 6490 3760
rect 6630 4100 6690 4120
rect 6630 4060 6640 4100
rect 6680 4060 6690 4100
rect 6630 4000 6690 4060
rect 6630 3960 6640 4000
rect 6680 3960 6690 4000
rect 6630 3900 6690 3960
rect 6630 3860 6640 3900
rect 6680 3860 6690 3900
rect 6630 3800 6690 3860
rect 6630 3760 6640 3800
rect 6680 3760 6690 3800
rect 6630 3740 6690 3760
rect 6830 4100 6890 4120
rect 6830 4060 6840 4100
rect 6880 4060 6890 4100
rect 6830 4000 6890 4060
rect 6830 3960 6840 4000
rect 6880 3960 6890 4000
rect 6830 3900 6890 3960
rect 6830 3860 6840 3900
rect 6880 3860 6890 3900
rect 6830 3800 6890 3860
rect 6830 3760 6840 3800
rect 6880 3760 6890 3800
rect 6830 3740 6890 3760
rect 7030 4100 7250 4120
rect 7030 4060 7040 4100
rect 7080 4060 7120 4100
rect 7160 4060 7200 4100
rect 7240 4060 7250 4100
rect 7030 4000 7250 4060
rect 7030 3960 7040 4000
rect 7080 3960 7120 4000
rect 7160 3960 7200 4000
rect 7240 3960 7250 4000
rect 7030 3900 7250 3960
rect 7030 3860 7040 3900
rect 7080 3860 7120 3900
rect 7160 3860 7200 3900
rect 7240 3860 7250 3900
rect 7030 3800 7250 3860
rect 7030 3760 7040 3800
rect 7080 3760 7120 3800
rect 7160 3760 7200 3800
rect 7240 3760 7250 3800
rect 7030 3740 7250 3760
rect 7390 4100 7450 4120
rect 7390 4060 7400 4100
rect 7440 4060 7450 4100
rect 7390 4000 7450 4060
rect 7390 3960 7400 4000
rect 7440 3960 7450 4000
rect 7390 3900 7450 3960
rect 7390 3860 7400 3900
rect 7440 3860 7450 3900
rect 7390 3800 7450 3860
rect 7390 3760 7400 3800
rect 7440 3760 7450 3800
rect 7390 3740 7450 3760
rect 7590 4100 7650 4120
rect 7590 4060 7600 4100
rect 7640 4060 7650 4100
rect 7590 4000 7650 4060
rect 7590 3960 7600 4000
rect 7640 3960 7650 4000
rect 7590 3900 7650 3960
rect 7590 3860 7600 3900
rect 7640 3860 7650 3900
rect 7590 3800 7650 3860
rect 7590 3760 7600 3800
rect 7640 3760 7650 3800
rect 7590 3740 7650 3760
rect 7790 4100 7850 4120
rect 7790 4060 7800 4100
rect 7840 4060 7850 4100
rect 7790 4000 7850 4060
rect 7790 3960 7800 4000
rect 7840 3960 7850 4000
rect 7790 3900 7850 3960
rect 7790 3860 7800 3900
rect 7840 3860 7850 3900
rect 7790 3800 7850 3860
rect 7790 3760 7800 3800
rect 7840 3760 7850 3800
rect 7790 3740 7850 3760
rect 7990 4100 8050 4120
rect 7990 4060 8000 4100
rect 8040 4060 8050 4100
rect 7990 4000 8050 4060
rect 7990 3960 8000 4000
rect 8040 3960 8050 4000
rect 7990 3900 8050 3960
rect 7990 3860 8000 3900
rect 8040 3860 8050 3900
rect 7990 3800 8050 3860
rect 7990 3760 8000 3800
rect 8040 3760 8050 3800
rect 7990 3740 8050 3760
rect 8190 4100 8250 4120
rect 8190 4060 8200 4100
rect 8240 4060 8250 4100
rect 8190 4000 8250 4060
rect 8190 3960 8200 4000
rect 8240 3960 8250 4000
rect 8190 3900 8250 3960
rect 8190 3860 8200 3900
rect 8240 3860 8250 3900
rect 8190 3800 8250 3860
rect 8190 3760 8200 3800
rect 8240 3760 8250 3800
rect 8190 3740 8250 3760
rect 8390 4100 8530 4120
rect 8390 4060 8400 4100
rect 8440 4060 8480 4100
rect 8520 4060 8530 4100
rect 8390 4000 8530 4060
rect 8390 3960 8400 4000
rect 8440 3960 8480 4000
rect 8520 3960 8530 4000
rect 8390 3900 8530 3960
rect 8390 3860 8400 3900
rect 8440 3860 8480 3900
rect 8520 3860 8530 3900
rect 8390 3800 8530 3860
rect 8390 3760 8400 3800
rect 8440 3760 8480 3800
rect 8520 3760 8530 3800
rect 8390 3740 8530 3760
rect 8760 4100 8820 4120
rect 8760 4060 8770 4100
rect 8810 4060 8820 4100
rect 8760 4000 8820 4060
rect 8760 3960 8770 4000
rect 8810 3960 8820 4000
rect 8760 3900 8820 3960
rect 8760 3860 8770 3900
rect 8810 3860 8820 3900
rect 8760 3800 8820 3860
rect 8760 3760 8770 3800
rect 8810 3760 8820 3800
rect 8760 3740 8820 3760
rect 8870 4100 8930 4120
rect 8870 4060 8880 4100
rect 8920 4060 8930 4100
rect 8870 4000 8930 4060
rect 8870 3960 8880 4000
rect 8920 3960 8930 4000
rect 8870 3900 8930 3960
rect 8870 3860 8880 3900
rect 8920 3860 8930 3900
rect 8870 3800 8930 3860
rect 8870 3760 8880 3800
rect 8920 3760 8930 3800
rect 8870 3740 8930 3760
rect 9010 4100 9070 4120
rect 9010 4060 9020 4100
rect 9060 4060 9070 4100
rect 9010 4000 9070 4060
rect 9010 3960 9020 4000
rect 9060 3960 9070 4000
rect 9010 3900 9070 3960
rect 9010 3860 9020 3900
rect 9060 3860 9070 3900
rect 9010 3800 9070 3860
rect 9010 3760 9020 3800
rect 9060 3760 9070 3800
rect 9010 3740 9070 3760
rect 9120 4100 9260 4120
rect 9120 4060 9130 4100
rect 9170 4060 9210 4100
rect 9250 4060 9260 4100
rect 9120 4000 9260 4060
rect 9120 3960 9130 4000
rect 9170 3960 9210 4000
rect 9250 3960 9260 4000
rect 9120 3900 9260 3960
rect 9120 3860 9130 3900
rect 9170 3860 9210 3900
rect 9250 3860 9260 3900
rect 9120 3800 9260 3860
rect 9120 3760 9130 3800
rect 9170 3760 9210 3800
rect 9250 3760 9260 3800
rect 9120 3740 9260 3760
rect 3790 3670 4230 3720
rect 4880 3610 4920 3740
rect 5280 3700 5320 3740
rect 6240 3700 6280 3740
rect 6640 3700 6680 3740
rect 7600 3700 7640 3740
rect 5260 3680 5340 3700
rect 5260 3640 5280 3680
rect 5320 3640 5340 3680
rect 6240 3680 6680 3700
rect 6240 3660 6440 3680
rect 5260 3620 5340 3640
rect 6420 3640 6440 3660
rect 6480 3660 6680 3680
rect 7580 3680 7660 3700
rect 6480 3640 6500 3660
rect 6420 3620 6500 3640
rect 7580 3640 7600 3680
rect 7640 3640 7660 3680
rect 7580 3620 7660 3640
rect 8000 3610 8040 3740
rect 2010 3550 2450 3600
rect 4860 3590 4940 3610
rect 4860 3550 4880 3590
rect 4920 3550 4940 3590
rect 4860 3530 4940 3550
rect 5540 3530 5620 3610
rect 6120 3590 6200 3610
rect 6120 3550 6140 3590
rect 6180 3550 6200 3590
rect 6120 3530 6200 3550
rect 6720 3590 6800 3610
rect 6720 3550 6740 3590
rect 6780 3550 6800 3590
rect 6720 3530 6800 3550
rect 7300 3530 7380 3610
rect 7980 3590 8060 3610
rect 7980 3550 8000 3590
rect 8040 3550 8060 3590
rect 7980 3530 8060 3550
rect 3790 3420 4230 3480
rect 6420 3500 6500 3520
rect 6420 3460 6440 3500
rect 6480 3460 6500 3500
rect 6420 3440 6500 3460
rect 8880 3430 8920 3740
rect 9010 3670 9050 3740
rect 8970 3650 9050 3670
rect 8970 3610 8990 3650
rect 9030 3610 9050 3650
rect 8970 3590 9050 3610
rect 3790 3380 3810 3420
rect 3850 3380 3900 3420
rect 3940 3380 3990 3420
rect 4030 3380 4080 3420
rect 4120 3380 4170 3420
rect 4210 3380 4230 3420
rect 3790 3360 4230 3380
rect 5540 3410 5620 3430
rect 5540 3370 5560 3410
rect 5600 3370 5620 3410
rect 5540 3350 5620 3370
rect 5940 3410 6020 3430
rect 5940 3370 5960 3410
rect 6000 3370 6020 3410
rect 5940 3350 6020 3370
rect 6060 3410 6140 3430
rect 6060 3370 6080 3410
rect 6120 3370 6140 3410
rect 6060 3350 6140 3370
rect 6780 3410 6860 3430
rect 6780 3370 6800 3410
rect 6840 3370 6860 3410
rect 6780 3350 6860 3370
rect 6900 3410 6980 3430
rect 6900 3370 6920 3410
rect 6960 3370 6980 3410
rect 6900 3350 6980 3370
rect 7300 3410 7380 3430
rect 7300 3370 7320 3410
rect 7360 3370 7380 3410
rect 7300 3350 7380 3370
rect 8860 3410 8940 3430
rect 8860 3370 8880 3410
rect 8920 3370 8940 3410
rect 8860 3350 8940 3370
rect 5560 3310 5600 3350
rect 5960 3310 6000 3350
rect 6920 3310 6960 3350
rect 7320 3310 7360 3350
rect 5060 3290 5210 3310
rect 5060 3250 5080 3290
rect 5120 3250 5160 3290
rect 5200 3250 5210 3290
rect 5060 3190 5210 3250
rect 5060 3150 5080 3190
rect 5120 3150 5160 3190
rect 5200 3150 5210 3190
rect 5060 3130 5210 3150
rect 5350 3290 5410 3310
rect 5350 3250 5360 3290
rect 5400 3250 5410 3290
rect 5350 3190 5410 3250
rect 5350 3150 5360 3190
rect 5400 3150 5410 3190
rect 5350 3130 5410 3150
rect 5550 3290 5610 3310
rect 5550 3250 5560 3290
rect 5600 3250 5610 3290
rect 5550 3190 5610 3250
rect 5550 3150 5560 3190
rect 5600 3150 5610 3190
rect 5550 3130 5610 3150
rect 5750 3290 5810 3310
rect 5750 3250 5760 3290
rect 5800 3250 5810 3290
rect 5750 3190 5810 3250
rect 5750 3150 5760 3190
rect 5800 3150 5810 3190
rect 5750 3130 5810 3150
rect 5950 3290 6010 3310
rect 5950 3250 5960 3290
rect 6000 3250 6010 3290
rect 5950 3190 6010 3250
rect 5950 3150 5960 3190
rect 6000 3150 6010 3190
rect 5950 3130 6010 3150
rect 6150 3290 6210 3310
rect 6150 3250 6160 3290
rect 6200 3250 6210 3290
rect 6150 3190 6210 3250
rect 6150 3150 6160 3190
rect 6200 3150 6210 3190
rect 6150 3130 6210 3150
rect 6350 3290 6570 3310
rect 6350 3250 6360 3290
rect 6400 3250 6440 3290
rect 6480 3250 6520 3290
rect 6560 3250 6570 3290
rect 6350 3190 6570 3250
rect 6350 3150 6360 3190
rect 6400 3150 6440 3190
rect 6480 3150 6520 3190
rect 6560 3150 6570 3190
rect 6350 3130 6570 3150
rect 6710 3290 6770 3310
rect 6710 3250 6720 3290
rect 6760 3250 6770 3290
rect 6710 3190 6770 3250
rect 6710 3150 6720 3190
rect 6760 3150 6770 3190
rect 6710 3130 6770 3150
rect 6910 3290 6970 3310
rect 6910 3250 6920 3290
rect 6960 3250 6970 3290
rect 6910 3190 6970 3250
rect 6910 3150 6920 3190
rect 6960 3150 6970 3190
rect 6910 3130 6970 3150
rect 7110 3290 7170 3310
rect 7110 3250 7120 3290
rect 7160 3250 7170 3290
rect 7110 3190 7170 3250
rect 7110 3150 7120 3190
rect 7160 3150 7170 3190
rect 7110 3130 7170 3150
rect 7310 3290 7370 3310
rect 7310 3250 7320 3290
rect 7360 3250 7370 3290
rect 7310 3190 7370 3250
rect 7310 3150 7320 3190
rect 7360 3150 7370 3190
rect 7310 3130 7370 3150
rect 7510 3290 7570 3310
rect 7510 3250 7520 3290
rect 7560 3250 7570 3290
rect 7510 3190 7570 3250
rect 7510 3150 7520 3190
rect 7560 3150 7570 3190
rect 7510 3130 7570 3150
rect 7710 3290 7850 3310
rect 7710 3250 7720 3290
rect 7760 3250 7800 3290
rect 7840 3250 7850 3290
rect 7710 3190 7850 3250
rect 7710 3150 7720 3190
rect 7760 3150 7800 3190
rect 7840 3150 7850 3190
rect 7710 3130 7850 3150
rect 1890 3060 2010 3080
rect 1890 3020 1910 3060
rect 1950 3020 2010 3060
rect 1890 3010 2010 3020
rect 3590 3060 4230 3080
rect 3590 3020 3810 3060
rect 3850 3020 3900 3060
rect 3940 3020 3990 3060
rect 4030 3020 4080 3060
rect 4120 3020 4170 3060
rect 4210 3020 4230 3060
rect 3590 3010 4230 3020
rect 1890 3000 1970 3010
rect 3790 2960 4230 3010
rect 5160 3000 5200 3130
rect 5360 3000 5400 3130
rect 5540 3070 5620 3090
rect 5540 3030 5560 3070
rect 5600 3030 5620 3070
rect 5540 3010 5620 3030
rect 5760 3000 5800 3130
rect 6160 3000 6200 3130
rect 6360 3000 6400 3130
rect 6520 3000 6560 3130
rect 6720 3000 6760 3130
rect 7120 3000 7160 3130
rect 7300 3070 7380 3090
rect 7300 3030 7320 3070
rect 7360 3030 7380 3070
rect 7300 3010 7380 3030
rect 7520 3000 7560 3130
rect 7720 3000 7760 3130
rect 5140 2980 5220 3000
rect 5140 2940 5160 2980
rect 5200 2940 5220 2980
rect 5140 2920 5220 2940
rect 5340 2980 5420 3000
rect 5340 2940 5360 2980
rect 5400 2940 5420 2980
rect 5340 2920 5420 2940
rect 5740 2980 5820 3000
rect 5740 2940 5760 2980
rect 5800 2940 5820 2980
rect 5740 2920 5820 2940
rect 6140 2980 6220 3000
rect 6140 2940 6160 2980
rect 6200 2940 6220 2980
rect 6140 2920 6220 2940
rect 6340 2980 6420 3000
rect 6340 2940 6360 2980
rect 6400 2940 6420 2980
rect 6340 2920 6420 2940
rect 6500 2980 6580 3000
rect 6500 2940 6520 2980
rect 6560 2940 6580 2980
rect 6500 2920 6580 2940
rect 6700 2980 6780 3000
rect 6700 2940 6720 2980
rect 6760 2940 6780 2980
rect 6700 2920 6780 2940
rect 7100 2980 7180 3000
rect 7100 2940 7120 2980
rect 7160 2940 7180 2980
rect 7100 2920 7180 2940
rect 7500 2980 7580 3000
rect 7500 2940 7520 2980
rect 7560 2940 7580 2980
rect 7500 2920 7580 2940
rect 7700 2980 7780 3000
rect 7700 2940 7720 2980
rect 7760 2940 7780 2980
rect 7700 2920 7780 2940
rect 2010 2840 2450 2890
rect 5760 2880 5800 2920
rect 6160 2880 6200 2920
rect 5560 2860 6420 2880
rect 3790 2720 4230 2770
rect 5560 2820 5640 2860
rect 5680 2820 5720 2860
rect 5760 2820 5800 2860
rect 5840 2820 5880 2860
rect 5920 2820 5960 2860
rect 6000 2820 6040 2860
rect 6080 2820 6120 2860
rect 6160 2820 6200 2860
rect 6240 2820 6280 2860
rect 6320 2820 6360 2860
rect 6400 2820 6420 2860
rect 5560 2800 6420 2820
rect 6500 2860 7380 2880
rect 6500 2820 6520 2860
rect 6560 2820 6600 2860
rect 6640 2820 6680 2860
rect 6720 2820 6760 2860
rect 6800 2820 6840 2860
rect 6880 2820 6920 2860
rect 6960 2820 7000 2860
rect 7040 2820 7080 2860
rect 7120 2820 7160 2860
rect 7200 2820 7240 2860
rect 7280 2820 7320 2860
rect 7360 2820 7380 2860
rect 6500 2800 7380 2820
rect 5560 2760 5600 2800
rect 7320 2760 7360 2800
rect 4590 2740 4730 2760
rect 4590 2700 4600 2740
rect 4640 2700 4680 2740
rect 4720 2700 4730 2740
rect 2010 2600 2450 2650
rect 4590 2640 4730 2700
rect 4590 2600 4600 2640
rect 4640 2600 4680 2640
rect 4720 2600 4730 2640
rect 1890 2480 1970 2490
rect 3790 2480 4230 2530
rect 1890 2470 2010 2480
rect 1890 2430 1910 2470
rect 1950 2430 2010 2470
rect 1890 2410 2010 2430
rect 4590 2540 4730 2600
rect 4590 2500 4600 2540
rect 4640 2500 4680 2540
rect 4720 2500 4730 2540
rect 4590 2440 4730 2500
rect 4590 2400 4600 2440
rect 4640 2400 4680 2440
rect 4720 2400 4730 2440
rect 4590 2340 4730 2400
rect 4590 2300 4600 2340
rect 4640 2300 4680 2340
rect 4720 2300 4730 2340
rect 4590 2240 4730 2300
rect 4590 2200 4600 2240
rect 4640 2200 4680 2240
rect 4720 2200 4730 2240
rect 4590 2140 4730 2200
rect 4590 2100 4600 2140
rect 4640 2100 4680 2140
rect 4720 2100 4730 2140
rect 4590 2040 4730 2100
rect 4590 2000 4600 2040
rect 4640 2000 4680 2040
rect 4720 2000 4730 2040
rect 4590 1980 4730 2000
rect 5550 2740 5610 2760
rect 5550 2700 5560 2740
rect 5600 2700 5610 2740
rect 5550 2640 5610 2700
rect 5550 2600 5560 2640
rect 5600 2600 5610 2640
rect 5550 2540 5610 2600
rect 5550 2500 5560 2540
rect 5600 2500 5610 2540
rect 5550 2440 5610 2500
rect 5550 2400 5560 2440
rect 5600 2400 5610 2440
rect 5550 2340 5610 2400
rect 5550 2300 5560 2340
rect 5600 2300 5610 2340
rect 5550 2240 5610 2300
rect 5550 2200 5560 2240
rect 5600 2200 5610 2240
rect 5550 2140 5610 2200
rect 5550 2100 5560 2140
rect 5600 2100 5610 2140
rect 5550 2040 5610 2100
rect 5550 2000 5560 2040
rect 5600 2000 5610 2040
rect 5550 1980 5610 2000
rect 6430 2740 6490 2760
rect 6430 2700 6440 2740
rect 6480 2700 6490 2740
rect 6430 2640 6490 2700
rect 6430 2600 6440 2640
rect 6480 2600 6490 2640
rect 6430 2540 6490 2600
rect 6430 2500 6440 2540
rect 6480 2500 6490 2540
rect 6430 2440 6490 2500
rect 6430 2400 6440 2440
rect 6480 2400 6490 2440
rect 6430 2340 6490 2400
rect 6430 2300 6440 2340
rect 6480 2300 6490 2340
rect 6430 2240 6490 2300
rect 6430 2200 6440 2240
rect 6480 2200 6490 2240
rect 6430 2140 6490 2200
rect 6430 2100 6440 2140
rect 6480 2100 6490 2140
rect 6430 2040 6490 2100
rect 6430 2000 6440 2040
rect 6480 2000 6490 2040
rect 6430 1980 6490 2000
rect 7310 2740 7370 2760
rect 7310 2700 7320 2740
rect 7360 2700 7370 2740
rect 7310 2640 7370 2700
rect 7310 2600 7320 2640
rect 7360 2600 7370 2640
rect 7310 2540 7370 2600
rect 7310 2500 7320 2540
rect 7360 2500 7370 2540
rect 7310 2440 7370 2500
rect 7310 2400 7320 2440
rect 7360 2400 7370 2440
rect 7310 2340 7370 2400
rect 7310 2300 7320 2340
rect 7360 2300 7370 2340
rect 7310 2240 7370 2300
rect 7310 2200 7320 2240
rect 7360 2200 7370 2240
rect 7310 2140 7370 2200
rect 7310 2100 7320 2140
rect 7360 2100 7370 2140
rect 7310 2040 7370 2100
rect 7310 2000 7320 2040
rect 7360 2000 7370 2040
rect 7310 1980 7370 2000
rect 8190 2740 8330 2760
rect 8190 2700 8200 2740
rect 8240 2700 8280 2740
rect 8320 2700 8330 2740
rect 8190 2640 8330 2700
rect 8190 2600 8200 2640
rect 8240 2600 8280 2640
rect 8320 2600 8330 2640
rect 8190 2540 8330 2600
rect 8190 2500 8200 2540
rect 8240 2500 8280 2540
rect 8320 2500 8330 2540
rect 8190 2440 8330 2500
rect 8190 2400 8200 2440
rect 8240 2400 8280 2440
rect 8320 2400 8330 2440
rect 8190 2340 8330 2400
rect 8190 2300 8200 2340
rect 8240 2300 8280 2340
rect 8320 2300 8330 2340
rect 8190 2240 8330 2300
rect 8190 2200 8200 2240
rect 8240 2200 8280 2240
rect 8320 2200 8330 2240
rect 8190 2140 8330 2200
rect 8190 2100 8200 2140
rect 8240 2100 8280 2140
rect 8320 2100 8330 2140
rect 8190 2040 8330 2100
rect 8190 2000 8200 2040
rect 8240 2000 8280 2040
rect 8320 2000 8330 2040
rect 8190 1980 8330 2000
rect 4680 1940 4720 1980
rect 6440 1940 6480 1980
rect 8200 1940 8240 1980
rect 4660 1920 4740 1940
rect 4660 1880 4680 1920
rect 4720 1880 4740 1920
rect 4660 1860 4740 1880
rect 6420 1920 6500 1940
rect 6420 1880 6440 1920
rect 6480 1880 6500 1920
rect 6420 1860 6500 1880
rect 8180 1920 8260 1940
rect 8180 1880 8200 1920
rect 8240 1880 8260 1920
rect 8180 1860 8260 1880
rect 5380 1800 7520 1820
rect 5380 1760 5460 1800
rect 5500 1760 5620 1800
rect 5660 1760 5780 1800
rect 5820 1760 5940 1800
rect 5980 1760 6100 1800
rect 6140 1760 6260 1800
rect 6300 1760 6420 1800
rect 6460 1760 6580 1800
rect 6620 1760 6740 1800
rect 6780 1760 6900 1800
rect 6940 1760 7060 1800
rect 7100 1760 7220 1800
rect 7260 1760 7380 1800
rect 7420 1760 7460 1800
rect 7500 1760 7520 1800
rect 5380 1740 7520 1760
rect 5380 1700 5420 1740
rect 5370 1680 5430 1700
rect 5370 1640 5380 1680
rect 5420 1640 5430 1680
rect 5370 1580 5430 1640
rect 5370 1540 5380 1580
rect 5420 1540 5430 1580
rect 5370 1520 5430 1540
rect 7450 1680 7590 1700
rect 7450 1640 7460 1680
rect 7500 1640 7540 1680
rect 7580 1640 7590 1680
rect 7450 1580 7590 1640
rect 7450 1540 7460 1580
rect 7500 1540 7540 1580
rect 7580 1540 7590 1580
rect 7450 1520 7590 1540
rect 1190 1410 1270 1430
rect 1190 1370 1210 1410
rect 1250 1370 1270 1410
rect 1190 1320 1270 1370
rect 1410 1410 1490 1430
rect 1410 1370 1430 1410
rect 1470 1370 1490 1410
rect 1410 1320 1490 1370
rect 10 1279 9470 1320
rect 10 1256 1506 1279
rect 10 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2866 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2770 1256
rect 2804 1245 2866 1256
rect 2900 1245 2956 1279
rect 2990 1245 3046 1279
rect 3080 1245 3136 1279
rect 3170 1245 3226 1279
rect 3260 1245 3316 1279
rect 3350 1245 3406 1279
rect 3440 1245 3496 1279
rect 3530 1245 3586 1279
rect 3620 1245 3676 1279
rect 3710 1245 3766 1279
rect 3800 1245 3856 1279
rect 3890 1256 4226 1279
rect 3890 1245 3957 1256
rect 2804 1222 3957 1245
rect 3991 1222 4130 1256
rect 4164 1245 4226 1256
rect 4260 1245 4316 1279
rect 4350 1245 4406 1279
rect 4440 1245 4496 1279
rect 4530 1245 4586 1279
rect 4620 1245 4676 1279
rect 4710 1245 4766 1279
rect 4800 1245 4856 1279
rect 4890 1245 4946 1279
rect 4980 1245 5036 1279
rect 5070 1245 5126 1279
rect 5160 1245 5216 1279
rect 5250 1256 5586 1279
rect 5250 1245 5317 1256
rect 4164 1222 5317 1245
rect 5351 1222 5490 1256
rect 5524 1245 5586 1256
rect 5620 1245 5676 1279
rect 5710 1245 5766 1279
rect 5800 1245 5856 1279
rect 5890 1245 5946 1279
rect 5980 1245 6036 1279
rect 6070 1245 6126 1279
rect 6160 1245 6216 1279
rect 6250 1245 6306 1279
rect 6340 1245 6396 1279
rect 6430 1245 6486 1279
rect 6520 1245 6576 1279
rect 6610 1256 6946 1279
rect 6610 1245 6677 1256
rect 5524 1222 6677 1245
rect 6711 1222 6850 1256
rect 6884 1245 6946 1256
rect 6980 1245 7036 1279
rect 7070 1245 7126 1279
rect 7160 1245 7216 1279
rect 7250 1245 7306 1279
rect 7340 1245 7396 1279
rect 7430 1245 7486 1279
rect 7520 1245 7576 1279
rect 7610 1245 7666 1279
rect 7700 1245 7756 1279
rect 7790 1245 7846 1279
rect 7880 1245 7936 1279
rect 7970 1256 8306 1279
rect 7970 1245 8037 1256
rect 6884 1222 8037 1245
rect 8071 1222 8210 1256
rect 8244 1245 8306 1256
rect 8340 1245 8396 1279
rect 8430 1245 8486 1279
rect 8520 1245 8576 1279
rect 8610 1245 8666 1279
rect 8700 1245 8756 1279
rect 8790 1245 8846 1279
rect 8880 1245 8936 1279
rect 8970 1245 9026 1279
rect 9060 1245 9116 1279
rect 9150 1245 9206 1279
rect 9240 1245 9296 1279
rect 9330 1256 9470 1279
rect 9330 1245 9397 1256
rect 8244 1222 9397 1245
rect 9431 1222 9470 1256
rect 10 1166 9470 1222
rect 10 1132 1410 1166
rect 1444 1132 2597 1166
rect 2631 1132 2770 1166
rect 2804 1132 3957 1166
rect 3991 1132 4130 1166
rect 4164 1132 5317 1166
rect 5351 1132 5490 1166
rect 5524 1132 6677 1166
rect 6711 1132 6850 1166
rect 6884 1132 8037 1166
rect 8071 1132 8210 1166
rect 8244 1132 9397 1166
rect 9431 1132 9470 1166
rect 10 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 3030 1132
rect 3064 1098 3120 1132
rect 3154 1098 3210 1132
rect 3244 1098 3300 1132
rect 3334 1098 3390 1132
rect 3424 1098 3480 1132
rect 3514 1098 3570 1132
rect 3604 1098 3660 1132
rect 3694 1098 3750 1132
rect 3784 1098 4390 1132
rect 4424 1098 4480 1132
rect 4514 1098 4570 1132
rect 4604 1098 4660 1132
rect 4694 1098 4750 1132
rect 4784 1098 4840 1132
rect 4874 1098 4930 1132
rect 4964 1098 5020 1132
rect 5054 1098 5110 1132
rect 5144 1098 5750 1132
rect 5784 1098 5840 1132
rect 5874 1098 5930 1132
rect 5964 1098 6020 1132
rect 6054 1098 6110 1132
rect 6144 1098 6200 1132
rect 6234 1098 6290 1132
rect 6324 1098 6380 1132
rect 6414 1098 6470 1132
rect 6504 1098 7110 1132
rect 7144 1098 7200 1132
rect 7234 1098 7290 1132
rect 7324 1098 7380 1132
rect 7414 1098 7470 1132
rect 7504 1098 7560 1132
rect 7594 1098 7650 1132
rect 7684 1098 7740 1132
rect 7774 1098 7830 1132
rect 7864 1098 8470 1132
rect 8504 1098 8560 1132
rect 8594 1098 8650 1132
rect 8684 1098 8740 1132
rect 8774 1098 8830 1132
rect 8864 1098 8920 1132
rect 8954 1098 9010 1132
rect 9044 1098 9100 1132
rect 9134 1098 9190 1132
rect 9224 1098 9470 1132
rect 10 1079 9470 1098
rect 10 1076 1620 1079
rect 10 1070 1410 1076
rect 10 270 260 1070
rect 1060 1042 1410 1070
rect 1444 1075 1620 1076
rect 1444 1042 1558 1075
rect 1060 1041 1558 1042
rect 1592 1041 1620 1075
rect 1060 986 1620 1041
rect 2420 1076 2980 1079
rect 2420 1056 2597 1076
rect 2420 1022 2448 1056
rect 2482 1042 2597 1056
rect 2631 1042 2770 1076
rect 2804 1075 2980 1076
rect 2804 1042 2918 1075
rect 2482 1041 2918 1042
rect 2952 1041 2980 1075
rect 2482 1022 2980 1041
rect 1060 952 1410 986
rect 1444 985 1620 986
rect 1444 952 1558 985
rect 1060 951 1558 952
rect 1592 951 1620 985
rect 1060 896 1620 951
rect 1060 862 1410 896
rect 1444 895 1620 896
rect 1444 862 1558 895
rect 1060 861 1558 862
rect 1592 861 1620 895
rect 1060 806 1620 861
rect 1060 772 1410 806
rect 1444 805 1620 806
rect 1444 772 1558 805
rect 1060 771 1558 772
rect 1592 771 1620 805
rect 1060 716 1620 771
rect 1060 682 1410 716
rect 1444 715 1620 716
rect 1444 682 1558 715
rect 1060 681 1558 682
rect 1592 681 1620 715
rect 1060 626 1620 681
rect 1060 592 1410 626
rect 1444 625 1620 626
rect 1444 592 1558 625
rect 1060 591 1558 592
rect 1592 591 1620 625
rect 1060 536 1620 591
rect 1060 502 1410 536
rect 1444 535 1620 536
rect 1444 502 1558 535
rect 1060 501 1558 502
rect 1592 501 1620 535
rect 1060 446 1620 501
rect 1060 412 1410 446
rect 1444 445 1620 446
rect 1444 412 1558 445
rect 1060 411 1558 412
rect 1592 411 1620 445
rect 1060 356 1620 411
rect 1060 322 1410 356
rect 1444 355 1620 356
rect 1444 322 1558 355
rect 1060 321 1558 322
rect 1592 321 1620 355
rect 1673 958 2367 1017
rect 1673 924 1734 958
rect 1768 930 1824 958
rect 1858 930 1914 958
rect 1948 930 2004 958
rect 1780 924 1824 930
rect 1880 924 1914 930
rect 1980 924 2004 930
rect 2038 930 2094 958
rect 2038 924 2046 930
rect 1673 896 1746 924
rect 1780 896 1846 924
rect 1880 896 1946 924
rect 1980 896 2046 924
rect 2080 924 2094 930
rect 2128 930 2184 958
rect 2128 924 2146 930
rect 2080 896 2146 924
rect 2180 924 2184 930
rect 2218 930 2274 958
rect 2218 924 2246 930
rect 2308 924 2367 958
rect 2180 896 2246 924
rect 2280 896 2367 924
rect 1673 868 2367 896
rect 1673 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2367 868
rect 1673 830 2367 834
rect 1673 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2367 830
rect 1673 778 2367 796
rect 1673 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2367 778
rect 1673 730 2367 744
rect 1673 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2367 730
rect 1673 688 2367 696
rect 1673 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2367 688
rect 1673 630 2367 654
rect 1673 598 1746 630
rect 1780 598 1846 630
rect 1880 598 1946 630
rect 1980 598 2046 630
rect 1673 564 1734 598
rect 1780 596 1824 598
rect 1880 596 1914 598
rect 1980 596 2004 598
rect 1768 564 1824 596
rect 1858 564 1914 596
rect 1948 564 2004 596
rect 2038 596 2046 598
rect 2080 598 2146 630
rect 2080 596 2094 598
rect 2038 564 2094 596
rect 2128 596 2146 598
rect 2180 598 2246 630
rect 2280 598 2367 630
rect 2180 596 2184 598
rect 2128 564 2184 596
rect 2218 596 2246 598
rect 2218 564 2274 596
rect 2308 564 2367 598
rect 1673 530 2367 564
rect 1673 508 1746 530
rect 1780 508 1846 530
rect 1880 508 1946 530
rect 1980 508 2046 530
rect 1673 474 1734 508
rect 1780 496 1824 508
rect 1880 496 1914 508
rect 1980 496 2004 508
rect 1768 474 1824 496
rect 1858 474 1914 496
rect 1948 474 2004 496
rect 2038 496 2046 508
rect 2080 508 2146 530
rect 2080 496 2094 508
rect 2038 474 2094 496
rect 2128 496 2146 508
rect 2180 508 2246 530
rect 2280 508 2367 530
rect 2180 496 2184 508
rect 2128 474 2184 496
rect 2218 496 2246 508
rect 2218 474 2274 496
rect 2308 474 2367 508
rect 1673 430 2367 474
rect 1673 418 1746 430
rect 1780 418 1846 430
rect 1880 418 1946 430
rect 1980 418 2046 430
rect 1673 384 1734 418
rect 1780 396 1824 418
rect 1880 396 1914 418
rect 1980 396 2004 418
rect 1768 384 1824 396
rect 1858 384 1914 396
rect 1948 384 2004 396
rect 2038 396 2046 418
rect 2080 418 2146 430
rect 2080 396 2094 418
rect 2038 384 2094 396
rect 2128 396 2146 418
rect 2180 418 2246 430
rect 2280 418 2367 430
rect 2180 396 2184 418
rect 2128 384 2184 396
rect 2218 396 2246 418
rect 2218 384 2274 396
rect 2308 384 2367 418
rect 1673 323 2367 384
rect 2420 986 2980 1022
rect 3780 1076 4340 1079
rect 3780 1056 3957 1076
rect 3780 1022 3808 1056
rect 3842 1042 3957 1056
rect 3991 1042 4130 1076
rect 4164 1075 4340 1076
rect 4164 1042 4278 1075
rect 3842 1041 4278 1042
rect 4312 1041 4340 1075
rect 3842 1022 4340 1041
rect 2420 966 2597 986
rect 2420 932 2448 966
rect 2482 952 2597 966
rect 2631 952 2770 986
rect 2804 985 2980 986
rect 2804 952 2918 985
rect 2482 951 2918 952
rect 2952 951 2980 985
rect 2482 932 2980 951
rect 2420 896 2980 932
rect 2420 876 2597 896
rect 2420 842 2448 876
rect 2482 862 2597 876
rect 2631 862 2770 896
rect 2804 895 2980 896
rect 2804 862 2918 895
rect 2482 861 2918 862
rect 2952 861 2980 895
rect 2482 842 2980 861
rect 2420 806 2980 842
rect 2420 786 2597 806
rect 2420 752 2448 786
rect 2482 772 2597 786
rect 2631 772 2770 806
rect 2804 805 2980 806
rect 2804 772 2918 805
rect 2482 771 2918 772
rect 2952 771 2980 805
rect 2482 752 2980 771
rect 2420 716 2980 752
rect 2420 696 2597 716
rect 2420 662 2448 696
rect 2482 682 2597 696
rect 2631 682 2770 716
rect 2804 715 2980 716
rect 2804 682 2918 715
rect 2482 681 2918 682
rect 2952 681 2980 715
rect 2482 662 2980 681
rect 2420 626 2980 662
rect 2420 606 2597 626
rect 2420 572 2448 606
rect 2482 592 2597 606
rect 2631 592 2770 626
rect 2804 625 2980 626
rect 2804 592 2918 625
rect 2482 591 2918 592
rect 2952 591 2980 625
rect 2482 572 2980 591
rect 2420 536 2980 572
rect 2420 516 2597 536
rect 2420 482 2448 516
rect 2482 502 2597 516
rect 2631 502 2770 536
rect 2804 535 2980 536
rect 2804 502 2918 535
rect 2482 501 2918 502
rect 2952 501 2980 535
rect 2482 482 2980 501
rect 2420 446 2980 482
rect 2420 426 2597 446
rect 2420 392 2448 426
rect 2482 412 2597 426
rect 2631 412 2770 446
rect 2804 445 2980 446
rect 2804 412 2918 445
rect 2482 411 2918 412
rect 2952 411 2980 445
rect 2482 392 2980 411
rect 2420 356 2980 392
rect 2420 336 2597 356
rect 1060 270 1620 321
rect 2420 302 2448 336
rect 2482 322 2597 336
rect 2631 322 2770 356
rect 2804 355 2980 356
rect 2804 322 2918 355
rect 2482 321 2918 322
rect 2952 321 2980 355
rect 3033 958 3727 1017
rect 3033 924 3094 958
rect 3128 930 3184 958
rect 3218 930 3274 958
rect 3308 930 3364 958
rect 3140 924 3184 930
rect 3240 924 3274 930
rect 3340 924 3364 930
rect 3398 930 3454 958
rect 3398 924 3406 930
rect 3033 896 3106 924
rect 3140 896 3206 924
rect 3240 896 3306 924
rect 3340 896 3406 924
rect 3440 924 3454 930
rect 3488 930 3544 958
rect 3488 924 3506 930
rect 3440 896 3506 924
rect 3540 924 3544 930
rect 3578 930 3634 958
rect 3578 924 3606 930
rect 3668 924 3727 958
rect 3540 896 3606 924
rect 3640 896 3727 924
rect 3033 868 3727 896
rect 3033 834 3094 868
rect 3128 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3727 868
rect 3033 830 3727 834
rect 3033 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3727 830
rect 3033 778 3727 796
rect 3033 744 3094 778
rect 3128 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3727 778
rect 3033 730 3727 744
rect 3033 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3727 730
rect 3033 688 3727 696
rect 3033 654 3094 688
rect 3128 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3727 688
rect 3033 630 3727 654
rect 3033 598 3106 630
rect 3140 598 3206 630
rect 3240 598 3306 630
rect 3340 598 3406 630
rect 3033 564 3094 598
rect 3140 596 3184 598
rect 3240 596 3274 598
rect 3340 596 3364 598
rect 3128 564 3184 596
rect 3218 564 3274 596
rect 3308 564 3364 596
rect 3398 596 3406 598
rect 3440 598 3506 630
rect 3440 596 3454 598
rect 3398 564 3454 596
rect 3488 596 3506 598
rect 3540 598 3606 630
rect 3640 598 3727 630
rect 3540 596 3544 598
rect 3488 564 3544 596
rect 3578 596 3606 598
rect 3578 564 3634 596
rect 3668 564 3727 598
rect 3033 530 3727 564
rect 3033 508 3106 530
rect 3140 508 3206 530
rect 3240 508 3306 530
rect 3340 508 3406 530
rect 3033 474 3094 508
rect 3140 496 3184 508
rect 3240 496 3274 508
rect 3340 496 3364 508
rect 3128 474 3184 496
rect 3218 474 3274 496
rect 3308 474 3364 496
rect 3398 496 3406 508
rect 3440 508 3506 530
rect 3440 496 3454 508
rect 3398 474 3454 496
rect 3488 496 3506 508
rect 3540 508 3606 530
rect 3640 508 3727 530
rect 3540 496 3544 508
rect 3488 474 3544 496
rect 3578 496 3606 508
rect 3578 474 3634 496
rect 3668 474 3727 508
rect 3033 430 3727 474
rect 3033 418 3106 430
rect 3140 418 3206 430
rect 3240 418 3306 430
rect 3340 418 3406 430
rect 3033 384 3094 418
rect 3140 396 3184 418
rect 3240 396 3274 418
rect 3340 396 3364 418
rect 3128 384 3184 396
rect 3218 384 3274 396
rect 3308 384 3364 396
rect 3398 396 3406 418
rect 3440 418 3506 430
rect 3440 396 3454 418
rect 3398 384 3454 396
rect 3488 396 3506 418
rect 3540 418 3606 430
rect 3640 418 3727 430
rect 3540 396 3544 418
rect 3488 384 3544 396
rect 3578 396 3606 418
rect 3578 384 3634 396
rect 3668 384 3727 418
rect 3033 323 3727 384
rect 3780 986 4340 1022
rect 5140 1076 5700 1079
rect 5140 1056 5317 1076
rect 5140 1022 5168 1056
rect 5202 1042 5317 1056
rect 5351 1042 5490 1076
rect 5524 1075 5700 1076
rect 5524 1042 5638 1075
rect 5202 1041 5638 1042
rect 5672 1041 5700 1075
rect 5202 1022 5700 1041
rect 3780 966 3957 986
rect 3780 932 3808 966
rect 3842 952 3957 966
rect 3991 952 4130 986
rect 4164 985 4340 986
rect 4164 952 4278 985
rect 3842 951 4278 952
rect 4312 951 4340 985
rect 3842 932 4340 951
rect 3780 896 4340 932
rect 3780 876 3957 896
rect 3780 842 3808 876
rect 3842 862 3957 876
rect 3991 862 4130 896
rect 4164 895 4340 896
rect 4164 862 4278 895
rect 3842 861 4278 862
rect 4312 861 4340 895
rect 3842 842 4340 861
rect 3780 806 4340 842
rect 3780 786 3957 806
rect 3780 752 3808 786
rect 3842 772 3957 786
rect 3991 772 4130 806
rect 4164 805 4340 806
rect 4164 772 4278 805
rect 3842 771 4278 772
rect 4312 771 4340 805
rect 3842 752 4340 771
rect 3780 716 4340 752
rect 3780 696 3957 716
rect 3780 662 3808 696
rect 3842 682 3957 696
rect 3991 682 4130 716
rect 4164 715 4340 716
rect 4164 682 4278 715
rect 3842 681 4278 682
rect 4312 681 4340 715
rect 3842 662 4340 681
rect 3780 626 4340 662
rect 3780 606 3957 626
rect 3780 572 3808 606
rect 3842 592 3957 606
rect 3991 592 4130 626
rect 4164 625 4340 626
rect 4164 592 4278 625
rect 3842 591 4278 592
rect 4312 591 4340 625
rect 3842 572 4340 591
rect 3780 536 4340 572
rect 3780 516 3957 536
rect 3780 482 3808 516
rect 3842 502 3957 516
rect 3991 502 4130 536
rect 4164 535 4340 536
rect 4164 502 4278 535
rect 3842 501 4278 502
rect 4312 501 4340 535
rect 3842 482 4340 501
rect 3780 446 4340 482
rect 3780 426 3957 446
rect 3780 392 3808 426
rect 3842 412 3957 426
rect 3991 412 4130 446
rect 4164 445 4340 446
rect 4164 412 4278 445
rect 3842 411 4278 412
rect 4312 411 4340 445
rect 3842 392 4340 411
rect 3780 356 4340 392
rect 3780 336 3957 356
rect 2482 302 2980 321
rect 2420 270 2980 302
rect 3780 302 3808 336
rect 3842 322 3957 336
rect 3991 322 4130 356
rect 4164 355 4340 356
rect 4164 322 4278 355
rect 3842 321 4278 322
rect 4312 321 4340 355
rect 4393 958 5087 1017
rect 4393 924 4454 958
rect 4488 930 4544 958
rect 4578 930 4634 958
rect 4668 930 4724 958
rect 4500 924 4544 930
rect 4600 924 4634 930
rect 4700 924 4724 930
rect 4758 930 4814 958
rect 4758 924 4766 930
rect 4393 896 4466 924
rect 4500 896 4566 924
rect 4600 896 4666 924
rect 4700 896 4766 924
rect 4800 924 4814 930
rect 4848 930 4904 958
rect 4848 924 4866 930
rect 4800 896 4866 924
rect 4900 924 4904 930
rect 4938 930 4994 958
rect 4938 924 4966 930
rect 5028 924 5087 958
rect 4900 896 4966 924
rect 5000 896 5087 924
rect 4393 868 5087 896
rect 4393 834 4454 868
rect 4488 834 4544 868
rect 4578 834 4634 868
rect 4668 834 4724 868
rect 4758 834 4814 868
rect 4848 834 4904 868
rect 4938 834 4994 868
rect 5028 834 5087 868
rect 4393 830 5087 834
rect 4393 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5087 830
rect 4393 778 5087 796
rect 4393 744 4454 778
rect 4488 744 4544 778
rect 4578 744 4634 778
rect 4668 744 4724 778
rect 4758 744 4814 778
rect 4848 744 4904 778
rect 4938 744 4994 778
rect 5028 744 5087 778
rect 4393 730 5087 744
rect 4393 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5087 730
rect 4393 688 5087 696
rect 4393 654 4454 688
rect 4488 654 4544 688
rect 4578 654 4634 688
rect 4668 654 4724 688
rect 4758 654 4814 688
rect 4848 654 4904 688
rect 4938 654 4994 688
rect 5028 654 5087 688
rect 4393 630 5087 654
rect 4393 598 4466 630
rect 4500 598 4566 630
rect 4600 598 4666 630
rect 4700 598 4766 630
rect 4393 564 4454 598
rect 4500 596 4544 598
rect 4600 596 4634 598
rect 4700 596 4724 598
rect 4488 564 4544 596
rect 4578 564 4634 596
rect 4668 564 4724 596
rect 4758 596 4766 598
rect 4800 598 4866 630
rect 4800 596 4814 598
rect 4758 564 4814 596
rect 4848 596 4866 598
rect 4900 598 4966 630
rect 5000 598 5087 630
rect 4900 596 4904 598
rect 4848 564 4904 596
rect 4938 596 4966 598
rect 4938 564 4994 596
rect 5028 564 5087 598
rect 4393 530 5087 564
rect 4393 508 4466 530
rect 4500 508 4566 530
rect 4600 508 4666 530
rect 4700 508 4766 530
rect 4393 474 4454 508
rect 4500 496 4544 508
rect 4600 496 4634 508
rect 4700 496 4724 508
rect 4488 474 4544 496
rect 4578 474 4634 496
rect 4668 474 4724 496
rect 4758 496 4766 508
rect 4800 508 4866 530
rect 4800 496 4814 508
rect 4758 474 4814 496
rect 4848 496 4866 508
rect 4900 508 4966 530
rect 5000 508 5087 530
rect 4900 496 4904 508
rect 4848 474 4904 496
rect 4938 496 4966 508
rect 4938 474 4994 496
rect 5028 474 5087 508
rect 4393 430 5087 474
rect 4393 418 4466 430
rect 4500 418 4566 430
rect 4600 418 4666 430
rect 4700 418 4766 430
rect 4393 384 4454 418
rect 4500 396 4544 418
rect 4600 396 4634 418
rect 4700 396 4724 418
rect 4488 384 4544 396
rect 4578 384 4634 396
rect 4668 384 4724 396
rect 4758 396 4766 418
rect 4800 418 4866 430
rect 4800 396 4814 418
rect 4758 384 4814 396
rect 4848 396 4866 418
rect 4900 418 4966 430
rect 5000 418 5087 430
rect 4900 396 4904 418
rect 4848 384 4904 396
rect 4938 396 4966 418
rect 4938 384 4994 396
rect 5028 384 5087 418
rect 4393 323 5087 384
rect 5140 986 5700 1022
rect 6500 1076 7060 1079
rect 6500 1056 6677 1076
rect 6500 1022 6528 1056
rect 6562 1042 6677 1056
rect 6711 1042 6850 1076
rect 6884 1075 7060 1076
rect 6884 1042 6998 1075
rect 6562 1041 6998 1042
rect 7032 1041 7060 1075
rect 6562 1022 7060 1041
rect 5140 966 5317 986
rect 5140 932 5168 966
rect 5202 952 5317 966
rect 5351 952 5490 986
rect 5524 985 5700 986
rect 5524 952 5638 985
rect 5202 951 5638 952
rect 5672 951 5700 985
rect 5202 932 5700 951
rect 5140 896 5700 932
rect 5140 876 5317 896
rect 5140 842 5168 876
rect 5202 862 5317 876
rect 5351 862 5490 896
rect 5524 895 5700 896
rect 5524 862 5638 895
rect 5202 861 5638 862
rect 5672 861 5700 895
rect 5202 842 5700 861
rect 5140 806 5700 842
rect 5140 786 5317 806
rect 5140 752 5168 786
rect 5202 772 5317 786
rect 5351 772 5490 806
rect 5524 805 5700 806
rect 5524 772 5638 805
rect 5202 771 5638 772
rect 5672 771 5700 805
rect 5202 752 5700 771
rect 5140 716 5700 752
rect 5140 696 5317 716
rect 5140 662 5168 696
rect 5202 682 5317 696
rect 5351 682 5490 716
rect 5524 715 5700 716
rect 5524 682 5638 715
rect 5202 681 5638 682
rect 5672 681 5700 715
rect 5202 662 5700 681
rect 5140 626 5700 662
rect 5140 606 5317 626
rect 5140 572 5168 606
rect 5202 592 5317 606
rect 5351 592 5490 626
rect 5524 625 5700 626
rect 5524 592 5638 625
rect 5202 591 5638 592
rect 5672 591 5700 625
rect 5202 572 5700 591
rect 5140 536 5700 572
rect 5140 516 5317 536
rect 5140 482 5168 516
rect 5202 502 5317 516
rect 5351 502 5490 536
rect 5524 535 5700 536
rect 5524 502 5638 535
rect 5202 501 5638 502
rect 5672 501 5700 535
rect 5202 482 5700 501
rect 5140 446 5700 482
rect 5140 426 5317 446
rect 5140 392 5168 426
rect 5202 412 5317 426
rect 5351 412 5490 446
rect 5524 445 5700 446
rect 5524 412 5638 445
rect 5202 411 5638 412
rect 5672 411 5700 445
rect 5202 392 5700 411
rect 5140 356 5700 392
rect 5140 336 5317 356
rect 3842 302 4340 321
rect 3780 270 4340 302
rect 5140 302 5168 336
rect 5202 322 5317 336
rect 5351 322 5490 356
rect 5524 355 5700 356
rect 5524 322 5638 355
rect 5202 321 5638 322
rect 5672 321 5700 355
rect 5753 958 6447 1017
rect 5753 924 5814 958
rect 5848 930 5904 958
rect 5938 930 5994 958
rect 6028 930 6084 958
rect 5860 924 5904 930
rect 5960 924 5994 930
rect 6060 924 6084 930
rect 6118 930 6174 958
rect 6118 924 6126 930
rect 5753 896 5826 924
rect 5860 896 5926 924
rect 5960 896 6026 924
rect 6060 896 6126 924
rect 6160 924 6174 930
rect 6208 930 6264 958
rect 6208 924 6226 930
rect 6160 896 6226 924
rect 6260 924 6264 930
rect 6298 930 6354 958
rect 6298 924 6326 930
rect 6388 924 6447 958
rect 6260 896 6326 924
rect 6360 896 6447 924
rect 5753 868 6447 896
rect 5753 834 5814 868
rect 5848 834 5904 868
rect 5938 834 5994 868
rect 6028 834 6084 868
rect 6118 834 6174 868
rect 6208 834 6264 868
rect 6298 834 6354 868
rect 6388 834 6447 868
rect 5753 830 6447 834
rect 5753 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6447 830
rect 5753 778 6447 796
rect 5753 744 5814 778
rect 5848 744 5904 778
rect 5938 744 5994 778
rect 6028 744 6084 778
rect 6118 744 6174 778
rect 6208 744 6264 778
rect 6298 744 6354 778
rect 6388 744 6447 778
rect 5753 730 6447 744
rect 5753 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6447 730
rect 5753 688 6447 696
rect 5753 654 5814 688
rect 5848 654 5904 688
rect 5938 654 5994 688
rect 6028 654 6084 688
rect 6118 654 6174 688
rect 6208 654 6264 688
rect 6298 654 6354 688
rect 6388 654 6447 688
rect 5753 630 6447 654
rect 5753 598 5826 630
rect 5860 598 5926 630
rect 5960 598 6026 630
rect 6060 598 6126 630
rect 5753 564 5814 598
rect 5860 596 5904 598
rect 5960 596 5994 598
rect 6060 596 6084 598
rect 5848 564 5904 596
rect 5938 564 5994 596
rect 6028 564 6084 596
rect 6118 596 6126 598
rect 6160 598 6226 630
rect 6160 596 6174 598
rect 6118 564 6174 596
rect 6208 596 6226 598
rect 6260 598 6326 630
rect 6360 598 6447 630
rect 6260 596 6264 598
rect 6208 564 6264 596
rect 6298 596 6326 598
rect 6298 564 6354 596
rect 6388 564 6447 598
rect 5753 530 6447 564
rect 5753 508 5826 530
rect 5860 508 5926 530
rect 5960 508 6026 530
rect 6060 508 6126 530
rect 5753 474 5814 508
rect 5860 496 5904 508
rect 5960 496 5994 508
rect 6060 496 6084 508
rect 5848 474 5904 496
rect 5938 474 5994 496
rect 6028 474 6084 496
rect 6118 496 6126 508
rect 6160 508 6226 530
rect 6160 496 6174 508
rect 6118 474 6174 496
rect 6208 496 6226 508
rect 6260 508 6326 530
rect 6360 508 6447 530
rect 6260 496 6264 508
rect 6208 474 6264 496
rect 6298 496 6326 508
rect 6298 474 6354 496
rect 6388 474 6447 508
rect 5753 430 6447 474
rect 5753 418 5826 430
rect 5860 418 5926 430
rect 5960 418 6026 430
rect 6060 418 6126 430
rect 5753 384 5814 418
rect 5860 396 5904 418
rect 5960 396 5994 418
rect 6060 396 6084 418
rect 5848 384 5904 396
rect 5938 384 5994 396
rect 6028 384 6084 396
rect 6118 396 6126 418
rect 6160 418 6226 430
rect 6160 396 6174 418
rect 6118 384 6174 396
rect 6208 396 6226 418
rect 6260 418 6326 430
rect 6360 418 6447 430
rect 6260 396 6264 418
rect 6208 384 6264 396
rect 6298 396 6326 418
rect 6298 384 6354 396
rect 6388 384 6447 418
rect 5753 323 6447 384
rect 6500 986 7060 1022
rect 7860 1076 8420 1079
rect 7860 1056 8037 1076
rect 7860 1022 7888 1056
rect 7922 1042 8037 1056
rect 8071 1042 8210 1076
rect 8244 1075 8420 1076
rect 8244 1042 8358 1075
rect 7922 1041 8358 1042
rect 8392 1041 8420 1075
rect 7922 1022 8420 1041
rect 6500 966 6677 986
rect 6500 932 6528 966
rect 6562 952 6677 966
rect 6711 952 6850 986
rect 6884 985 7060 986
rect 6884 952 6998 985
rect 6562 951 6998 952
rect 7032 951 7060 985
rect 6562 932 7060 951
rect 6500 896 7060 932
rect 6500 876 6677 896
rect 6500 842 6528 876
rect 6562 862 6677 876
rect 6711 862 6850 896
rect 6884 895 7060 896
rect 6884 862 6998 895
rect 6562 861 6998 862
rect 7032 861 7060 895
rect 6562 842 7060 861
rect 6500 806 7060 842
rect 6500 786 6677 806
rect 6500 752 6528 786
rect 6562 772 6677 786
rect 6711 772 6850 806
rect 6884 805 7060 806
rect 6884 772 6998 805
rect 6562 771 6998 772
rect 7032 771 7060 805
rect 6562 752 7060 771
rect 6500 716 7060 752
rect 6500 696 6677 716
rect 6500 662 6528 696
rect 6562 682 6677 696
rect 6711 682 6850 716
rect 6884 715 7060 716
rect 6884 682 6998 715
rect 6562 681 6998 682
rect 7032 681 7060 715
rect 6562 662 7060 681
rect 6500 626 7060 662
rect 6500 606 6677 626
rect 6500 572 6528 606
rect 6562 592 6677 606
rect 6711 592 6850 626
rect 6884 625 7060 626
rect 6884 592 6998 625
rect 6562 591 6998 592
rect 7032 591 7060 625
rect 6562 572 7060 591
rect 6500 536 7060 572
rect 6500 516 6677 536
rect 6500 482 6528 516
rect 6562 502 6677 516
rect 6711 502 6850 536
rect 6884 535 7060 536
rect 6884 502 6998 535
rect 6562 501 6998 502
rect 7032 501 7060 535
rect 6562 482 7060 501
rect 6500 446 7060 482
rect 6500 426 6677 446
rect 6500 392 6528 426
rect 6562 412 6677 426
rect 6711 412 6850 446
rect 6884 445 7060 446
rect 6884 412 6998 445
rect 6562 411 6998 412
rect 7032 411 7060 445
rect 6562 392 7060 411
rect 6500 356 7060 392
rect 6500 336 6677 356
rect 5202 302 5700 321
rect 5140 270 5700 302
rect 6500 302 6528 336
rect 6562 322 6677 336
rect 6711 322 6850 356
rect 6884 355 7060 356
rect 6884 322 6998 355
rect 6562 321 6998 322
rect 7032 321 7060 355
rect 7113 958 7807 1017
rect 7113 924 7174 958
rect 7208 930 7264 958
rect 7298 930 7354 958
rect 7388 930 7444 958
rect 7220 924 7264 930
rect 7320 924 7354 930
rect 7420 924 7444 930
rect 7478 930 7534 958
rect 7478 924 7486 930
rect 7113 896 7186 924
rect 7220 896 7286 924
rect 7320 896 7386 924
rect 7420 896 7486 924
rect 7520 924 7534 930
rect 7568 930 7624 958
rect 7568 924 7586 930
rect 7520 896 7586 924
rect 7620 924 7624 930
rect 7658 930 7714 958
rect 7658 924 7686 930
rect 7748 924 7807 958
rect 7620 896 7686 924
rect 7720 896 7807 924
rect 7113 868 7807 896
rect 7113 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7807 868
rect 7113 830 7807 834
rect 7113 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7807 830
rect 7113 778 7807 796
rect 7113 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7807 778
rect 7113 730 7807 744
rect 7113 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7807 730
rect 7113 688 7807 696
rect 7113 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7807 688
rect 7113 630 7807 654
rect 7113 598 7186 630
rect 7220 598 7286 630
rect 7320 598 7386 630
rect 7420 598 7486 630
rect 7113 564 7174 598
rect 7220 596 7264 598
rect 7320 596 7354 598
rect 7420 596 7444 598
rect 7208 564 7264 596
rect 7298 564 7354 596
rect 7388 564 7444 596
rect 7478 596 7486 598
rect 7520 598 7586 630
rect 7520 596 7534 598
rect 7478 564 7534 596
rect 7568 596 7586 598
rect 7620 598 7686 630
rect 7720 598 7807 630
rect 7620 596 7624 598
rect 7568 564 7624 596
rect 7658 596 7686 598
rect 7658 564 7714 596
rect 7748 564 7807 598
rect 7113 530 7807 564
rect 7113 508 7186 530
rect 7220 508 7286 530
rect 7320 508 7386 530
rect 7420 508 7486 530
rect 7113 474 7174 508
rect 7220 496 7264 508
rect 7320 496 7354 508
rect 7420 496 7444 508
rect 7208 474 7264 496
rect 7298 474 7354 496
rect 7388 474 7444 496
rect 7478 496 7486 508
rect 7520 508 7586 530
rect 7520 496 7534 508
rect 7478 474 7534 496
rect 7568 496 7586 508
rect 7620 508 7686 530
rect 7720 508 7807 530
rect 7620 496 7624 508
rect 7568 474 7624 496
rect 7658 496 7686 508
rect 7658 474 7714 496
rect 7748 474 7807 508
rect 7113 430 7807 474
rect 7113 418 7186 430
rect 7220 418 7286 430
rect 7320 418 7386 430
rect 7420 418 7486 430
rect 7113 384 7174 418
rect 7220 396 7264 418
rect 7320 396 7354 418
rect 7420 396 7444 418
rect 7208 384 7264 396
rect 7298 384 7354 396
rect 7388 384 7444 396
rect 7478 396 7486 418
rect 7520 418 7586 430
rect 7520 396 7534 418
rect 7478 384 7534 396
rect 7568 396 7586 418
rect 7620 418 7686 430
rect 7720 418 7807 430
rect 7620 396 7624 418
rect 7568 384 7624 396
rect 7658 396 7686 418
rect 7658 384 7714 396
rect 7748 384 7807 418
rect 7113 323 7807 384
rect 7860 986 8420 1022
rect 9220 1076 9470 1079
rect 9220 1056 9397 1076
rect 9220 1022 9248 1056
rect 9282 1042 9397 1056
rect 9431 1042 9470 1076
rect 9282 1022 9470 1042
rect 7860 966 8037 986
rect 7860 932 7888 966
rect 7922 952 8037 966
rect 8071 952 8210 986
rect 8244 985 8420 986
rect 8244 952 8358 985
rect 7922 951 8358 952
rect 8392 951 8420 985
rect 7922 932 8420 951
rect 7860 896 8420 932
rect 7860 876 8037 896
rect 7860 842 7888 876
rect 7922 862 8037 876
rect 8071 862 8210 896
rect 8244 895 8420 896
rect 8244 862 8358 895
rect 7922 861 8358 862
rect 8392 861 8420 895
rect 7922 842 8420 861
rect 7860 806 8420 842
rect 7860 786 8037 806
rect 7860 752 7888 786
rect 7922 772 8037 786
rect 8071 772 8210 806
rect 8244 805 8420 806
rect 8244 772 8358 805
rect 7922 771 8358 772
rect 8392 771 8420 805
rect 7922 752 8420 771
rect 7860 716 8420 752
rect 7860 696 8037 716
rect 7860 662 7888 696
rect 7922 682 8037 696
rect 8071 682 8210 716
rect 8244 715 8420 716
rect 8244 682 8358 715
rect 7922 681 8358 682
rect 8392 681 8420 715
rect 7922 662 8420 681
rect 7860 626 8420 662
rect 7860 606 8037 626
rect 7860 572 7888 606
rect 7922 592 8037 606
rect 8071 592 8210 626
rect 8244 625 8420 626
rect 8244 592 8358 625
rect 7922 591 8358 592
rect 8392 591 8420 625
rect 7922 572 8420 591
rect 7860 536 8420 572
rect 7860 516 8037 536
rect 7860 482 7888 516
rect 7922 502 8037 516
rect 8071 502 8210 536
rect 8244 535 8420 536
rect 8244 502 8358 535
rect 7922 501 8358 502
rect 8392 501 8420 535
rect 7922 482 8420 501
rect 7860 446 8420 482
rect 7860 426 8037 446
rect 7860 392 7888 426
rect 7922 412 8037 426
rect 8071 412 8210 446
rect 8244 445 8420 446
rect 8244 412 8358 445
rect 7922 411 8358 412
rect 8392 411 8420 445
rect 7922 392 8420 411
rect 7860 356 8420 392
rect 7860 336 8037 356
rect 6562 302 7060 321
rect 6500 270 7060 302
rect 7860 302 7888 336
rect 7922 322 8037 336
rect 8071 322 8210 356
rect 8244 355 8420 356
rect 8244 322 8358 355
rect 7922 321 8358 322
rect 8392 321 8420 355
rect 8473 958 9167 1017
rect 8473 924 8534 958
rect 8568 930 8624 958
rect 8658 930 8714 958
rect 8748 930 8804 958
rect 8580 924 8624 930
rect 8680 924 8714 930
rect 8780 924 8804 930
rect 8838 930 8894 958
rect 8838 924 8846 930
rect 8473 896 8546 924
rect 8580 896 8646 924
rect 8680 896 8746 924
rect 8780 896 8846 924
rect 8880 924 8894 930
rect 8928 930 8984 958
rect 8928 924 8946 930
rect 8880 896 8946 924
rect 8980 924 8984 930
rect 9018 930 9074 958
rect 9018 924 9046 930
rect 9108 924 9167 958
rect 8980 896 9046 924
rect 9080 896 9167 924
rect 8473 868 9167 896
rect 8473 834 8534 868
rect 8568 834 8624 868
rect 8658 834 8714 868
rect 8748 834 8804 868
rect 8838 834 8894 868
rect 8928 834 8984 868
rect 9018 834 9074 868
rect 9108 834 9167 868
rect 8473 830 9167 834
rect 8473 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9167 830
rect 8473 778 9167 796
rect 8473 744 8534 778
rect 8568 744 8624 778
rect 8658 744 8714 778
rect 8748 744 8804 778
rect 8838 744 8894 778
rect 8928 744 8984 778
rect 9018 744 9074 778
rect 9108 744 9167 778
rect 8473 730 9167 744
rect 8473 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9167 730
rect 8473 688 9167 696
rect 8473 654 8534 688
rect 8568 654 8624 688
rect 8658 654 8714 688
rect 8748 654 8804 688
rect 8838 654 8894 688
rect 8928 654 8984 688
rect 9018 654 9074 688
rect 9108 654 9167 688
rect 8473 630 9167 654
rect 8473 598 8546 630
rect 8580 598 8646 630
rect 8680 598 8746 630
rect 8780 598 8846 630
rect 8473 564 8534 598
rect 8580 596 8624 598
rect 8680 596 8714 598
rect 8780 596 8804 598
rect 8568 564 8624 596
rect 8658 564 8714 596
rect 8748 564 8804 596
rect 8838 596 8846 598
rect 8880 598 8946 630
rect 8880 596 8894 598
rect 8838 564 8894 596
rect 8928 596 8946 598
rect 8980 598 9046 630
rect 9080 598 9167 630
rect 8980 596 8984 598
rect 8928 564 8984 596
rect 9018 596 9046 598
rect 9018 564 9074 596
rect 9108 564 9167 598
rect 8473 530 9167 564
rect 8473 508 8546 530
rect 8580 508 8646 530
rect 8680 508 8746 530
rect 8780 508 8846 530
rect 8473 474 8534 508
rect 8580 496 8624 508
rect 8680 496 8714 508
rect 8780 496 8804 508
rect 8568 474 8624 496
rect 8658 474 8714 496
rect 8748 474 8804 496
rect 8838 496 8846 508
rect 8880 508 8946 530
rect 8880 496 8894 508
rect 8838 474 8894 496
rect 8928 496 8946 508
rect 8980 508 9046 530
rect 9080 508 9167 530
rect 8980 496 8984 508
rect 8928 474 8984 496
rect 9018 496 9046 508
rect 9018 474 9074 496
rect 9108 474 9167 508
rect 8473 430 9167 474
rect 8473 418 8546 430
rect 8580 418 8646 430
rect 8680 418 8746 430
rect 8780 418 8846 430
rect 8473 384 8534 418
rect 8580 396 8624 418
rect 8680 396 8714 418
rect 8780 396 8804 418
rect 8568 384 8624 396
rect 8658 384 8714 396
rect 8748 384 8804 396
rect 8838 396 8846 418
rect 8880 418 8946 430
rect 8880 396 8894 418
rect 8838 384 8894 396
rect 8928 396 8946 418
rect 8980 418 9046 430
rect 9080 418 9167 430
rect 8980 396 8984 418
rect 8928 384 8984 396
rect 9018 396 9046 418
rect 9018 384 9074 396
rect 9108 384 9167 418
rect 8473 323 9167 384
rect 9220 986 9470 1022
rect 9220 966 9397 986
rect 9220 932 9248 966
rect 9282 952 9397 966
rect 9431 952 9470 986
rect 9282 932 9470 952
rect 9220 896 9470 932
rect 9220 876 9397 896
rect 9220 842 9248 876
rect 9282 862 9397 876
rect 9431 862 9470 896
rect 9282 842 9470 862
rect 9220 806 9470 842
rect 9220 786 9397 806
rect 9220 752 9248 786
rect 9282 772 9397 786
rect 9431 772 9470 806
rect 9282 752 9470 772
rect 9220 716 9470 752
rect 9220 696 9397 716
rect 9220 662 9248 696
rect 9282 682 9397 696
rect 9431 682 9470 716
rect 9282 662 9470 682
rect 9220 626 9470 662
rect 9220 606 9397 626
rect 9220 572 9248 606
rect 9282 592 9397 606
rect 9431 592 9470 626
rect 9282 572 9470 592
rect 9220 536 9470 572
rect 9220 516 9397 536
rect 9220 482 9248 516
rect 9282 502 9397 516
rect 9431 502 9470 536
rect 9282 482 9470 502
rect 9220 446 9470 482
rect 9220 426 9397 446
rect 9220 392 9248 426
rect 9282 412 9397 426
rect 9431 412 9470 446
rect 9282 392 9470 412
rect 9220 356 9470 392
rect 9220 336 9397 356
rect 7922 302 8420 321
rect 7860 270 8420 302
rect 9220 302 9248 336
rect 9282 322 9397 336
rect 9431 322 9470 356
rect 9282 302 9470 322
rect 9220 270 9470 302
rect 10 266 9470 270
rect 10 232 1410 266
rect 1444 242 2597 266
rect 1444 232 1636 242
rect 10 208 1636 232
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 232 2597 242
rect 2631 232 2770 266
rect 2804 242 3957 266
rect 2804 232 2996 242
rect 2390 208 2996 232
rect 3030 208 3086 242
rect 3120 208 3176 242
rect 3210 208 3266 242
rect 3300 208 3356 242
rect 3390 208 3446 242
rect 3480 208 3536 242
rect 3570 208 3626 242
rect 3660 208 3716 242
rect 3750 232 3957 242
rect 3991 232 4130 266
rect 4164 242 5317 266
rect 4164 232 4356 242
rect 3750 208 4356 232
rect 4390 208 4446 242
rect 4480 208 4536 242
rect 4570 208 4626 242
rect 4660 208 4716 242
rect 4750 208 4806 242
rect 4840 208 4896 242
rect 4930 208 4986 242
rect 5020 208 5076 242
rect 5110 232 5317 242
rect 5351 232 5490 266
rect 5524 242 6677 266
rect 5524 232 5716 242
rect 5110 208 5716 232
rect 5750 208 5806 242
rect 5840 208 5896 242
rect 5930 208 5986 242
rect 6020 208 6076 242
rect 6110 208 6166 242
rect 6200 208 6256 242
rect 6290 208 6346 242
rect 6380 208 6436 242
rect 6470 232 6677 242
rect 6711 232 6850 266
rect 6884 242 8037 266
rect 6884 232 7076 242
rect 6470 208 7076 232
rect 7110 208 7166 242
rect 7200 208 7256 242
rect 7290 208 7346 242
rect 7380 208 7436 242
rect 7470 208 7526 242
rect 7560 208 7616 242
rect 7650 208 7706 242
rect 7740 208 7796 242
rect 7830 232 8037 242
rect 8071 232 8210 266
rect 8244 242 9397 266
rect 8244 232 8436 242
rect 7830 208 8436 232
rect 8470 208 8526 242
rect 8560 208 8616 242
rect 8650 208 8706 242
rect 8740 208 8796 242
rect 8830 208 8886 242
rect 8920 208 8976 242
rect 9010 208 9066 242
rect 9100 208 9156 242
rect 9190 232 9397 242
rect 9431 232 9470 266
rect 9190 208 9470 232
rect 10 176 9470 208
rect 10 142 1410 176
rect 1444 142 2597 176
rect 2631 142 2770 176
rect 2804 142 3957 176
rect 3991 142 4130 176
rect 4164 142 5317 176
rect 5351 142 5490 176
rect 5524 142 6677 176
rect 6711 142 6850 176
rect 6884 142 8037 176
rect 8071 142 8210 176
rect 8244 142 9397 176
rect 9431 142 9470 176
rect 10 92 9470 142
rect 10 90 1506 92
rect 10 50 40 90
rect 80 50 220 90
rect 260 50 400 90
rect 440 50 580 90
rect 620 50 760 90
rect 800 50 940 90
rect 980 50 1120 90
rect 1160 50 1300 90
rect 1340 50 1480 90
rect 1540 58 1596 92
rect 1630 90 1686 92
rect 1630 58 1660 90
rect 1720 58 1776 92
rect 1810 90 1866 92
rect 1810 58 1840 90
rect 1900 58 1956 92
rect 1990 90 2046 92
rect 1990 58 2020 90
rect 2080 58 2136 92
rect 2170 90 2226 92
rect 2170 58 2200 90
rect 2260 58 2316 92
rect 2350 90 2406 92
rect 2350 58 2380 90
rect 2440 58 2496 92
rect 2530 90 2586 92
rect 2620 90 2766 92
rect 2530 58 2560 90
rect 1520 50 1660 58
rect 1700 50 1840 58
rect 1880 50 2020 58
rect 2060 50 2200 58
rect 2240 50 2380 58
rect 2420 50 2560 58
rect 2620 58 2740 90
rect 2600 50 2740 58
rect 2800 58 2866 92
rect 2900 90 2946 92
rect 2900 58 2920 90
rect 2990 58 3046 92
rect 3080 90 3126 92
rect 3080 58 3100 90
rect 3170 58 3226 92
rect 3260 90 3306 92
rect 3260 58 3280 90
rect 3350 58 3406 92
rect 3440 90 3486 92
rect 3440 58 3460 90
rect 3530 58 3586 92
rect 3620 90 3666 92
rect 3620 58 3640 90
rect 3710 58 3766 92
rect 3800 90 3846 92
rect 3800 58 3820 90
rect 3890 58 3970 92
rect 3980 90 4026 92
rect 3980 58 4000 90
rect 2780 50 2920 58
rect 2960 50 3100 58
rect 3140 50 3280 58
rect 3320 50 3460 58
rect 3500 50 3640 58
rect 3680 50 3820 58
rect 3860 50 4000 58
rect 4070 58 4150 92
rect 4160 90 4206 92
rect 4160 58 4180 90
rect 4040 50 4180 58
rect 4260 58 4316 92
rect 4350 90 4386 92
rect 4350 58 4360 90
rect 4220 50 4360 58
rect 4440 58 4496 92
rect 4530 90 4566 92
rect 4530 58 4540 90
rect 4400 50 4540 58
rect 4620 58 4676 92
rect 4710 90 4746 92
rect 4710 58 4720 90
rect 4580 50 4720 58
rect 4800 58 4856 92
rect 4890 90 4926 92
rect 4890 58 4900 90
rect 4760 50 4900 58
rect 4980 58 5036 92
rect 5070 90 5106 92
rect 5070 58 5080 90
rect 4940 50 5080 58
rect 5160 58 5216 92
rect 5250 90 5286 92
rect 5250 58 5260 90
rect 5120 50 5260 58
rect 5330 58 5410 92
rect 5430 90 5466 92
rect 5430 58 5440 90
rect 5300 50 5440 58
rect 5510 58 5586 92
rect 5620 90 5646 92
rect 5480 50 5620 58
rect 5710 58 5766 92
rect 5800 90 5826 92
rect 5660 50 5800 58
rect 5890 58 5946 92
rect 5980 90 6006 92
rect 5840 50 5980 58
rect 6070 58 6126 92
rect 6160 90 6186 92
rect 6020 50 6160 58
rect 6250 58 6306 92
rect 6340 90 6366 92
rect 6200 50 6340 58
rect 6430 58 6486 92
rect 6520 90 6546 92
rect 6380 50 6520 58
rect 6610 58 6670 92
rect 6700 90 6726 92
rect 6560 50 6700 58
rect 6770 58 6850 92
rect 6880 90 6906 92
rect 6740 50 6880 58
rect 6980 58 7030 92
rect 7070 90 7086 92
rect 7160 58 7210 92
rect 7250 90 7266 92
rect 7340 58 7390 92
rect 7430 90 7446 92
rect 7520 58 7570 92
rect 7610 90 7626 92
rect 7700 58 7750 92
rect 7790 90 7806 92
rect 7880 58 7930 92
rect 7970 90 7986 92
rect 8030 58 8110 92
rect 8150 90 8166 92
rect 6920 50 7060 58
rect 7100 50 7240 58
rect 7280 50 7420 58
rect 7460 50 7600 58
rect 7640 50 7780 58
rect 7820 50 7960 58
rect 8000 50 8140 58
rect 8210 58 8290 92
rect 8340 90 8346 92
rect 8390 58 8396 92
rect 8430 58 8470 92
rect 8520 90 8526 92
rect 8570 58 8576 92
rect 8610 58 8650 92
rect 8700 90 8706 92
rect 8750 58 8756 92
rect 8790 58 8830 92
rect 8880 90 8886 92
rect 8930 58 8936 92
rect 8970 58 9010 92
rect 9060 90 9066 92
rect 9110 58 9116 92
rect 9150 58 9190 92
rect 9240 90 9246 92
rect 9290 58 9296 92
rect 9330 58 9370 92
rect 9420 90 9426 92
rect 8180 50 8320 58
rect 8360 50 8500 58
rect 8540 50 8680 58
rect 8720 50 8860 58
rect 8900 50 9040 58
rect 9080 50 9220 58
rect 9260 50 9400 58
rect 9440 50 9470 58
rect 10 20 9470 50
<< viali >>
rect 4640 5490 4680 5530
rect 5040 5490 5080 5530
rect 5440 5490 5480 5530
rect 5840 5490 5880 5530
rect 6240 5490 6280 5530
rect 6640 5490 6680 5530
rect 7040 5490 7080 5530
rect 7440 5490 7480 5530
rect 7840 5490 7880 5530
rect 8240 5490 8280 5530
rect 1910 4970 1950 5010
rect 4840 4550 4880 4590
rect 5240 4460 5280 4500
rect 6240 4550 6280 4590
rect 6040 4460 6080 4500
rect 6640 4550 6680 4590
rect 6840 4550 6880 4590
rect 7640 4550 7680 4590
rect 8160 4550 8200 4590
rect 8040 4460 8080 4500
rect 3810 4380 3850 4420
rect 3900 4380 3940 4420
rect 3990 4380 4030 4420
rect 4080 4380 4120 4420
rect 4170 4380 4210 4420
rect 5640 4370 5680 4410
rect 6440 4370 6480 4410
rect 7240 4370 7280 4410
rect 8770 4280 8810 4320
rect 4480 4180 4520 4220
rect 4680 4180 4720 4220
rect 5080 4180 5120 4220
rect 5480 4180 5520 4220
rect 5680 4180 5720 4220
rect 5840 4180 5880 4220
rect 6040 4180 6080 4220
rect 6240 4180 6280 4220
rect 6440 4180 6480 4220
rect 6640 4180 6680 4220
rect 6840 4180 6880 4220
rect 7040 4180 7080 4220
rect 7200 4180 7240 4220
rect 7400 4180 7440 4220
rect 7800 4180 7840 4220
rect 8200 4180 8240 4220
rect 8400 4180 8440 4220
rect 9170 4180 9210 4220
rect 1910 3970 1950 4010
rect 5280 3640 5320 3680
rect 6440 3640 6480 3680
rect 7600 3640 7640 3680
rect 4880 3550 4920 3590
rect 6140 3550 6180 3590
rect 6740 3550 6780 3590
rect 8000 3550 8040 3590
rect 6440 3460 6480 3500
rect 8990 3610 9030 3650
rect 3810 3380 3850 3420
rect 3900 3380 3940 3420
rect 3990 3380 4030 3420
rect 4080 3380 4120 3420
rect 4170 3380 4210 3420
rect 5560 3370 5600 3410
rect 5960 3370 6000 3410
rect 6080 3370 6120 3410
rect 6800 3370 6840 3410
rect 6920 3370 6960 3410
rect 7320 3370 7360 3410
rect 8880 3370 8920 3410
rect 1910 3020 1950 3060
rect 3810 3020 3850 3060
rect 3900 3020 3940 3060
rect 3990 3020 4030 3060
rect 4080 3020 4120 3060
rect 4170 3020 4210 3060
rect 5560 3030 5600 3070
rect 7320 3030 7360 3070
rect 5160 2940 5200 2980
rect 5360 2940 5400 2980
rect 5760 2940 5800 2980
rect 6160 2940 6200 2980
rect 6360 2940 6400 2980
rect 6520 2940 6560 2980
rect 6720 2940 6760 2980
rect 7120 2940 7160 2980
rect 7520 2940 7560 2980
rect 7720 2940 7760 2980
rect 7320 2820 7360 2860
rect 1910 2430 1950 2470
rect 4680 1880 4720 1920
rect 6440 1880 6480 1920
rect 8200 1880 8240 1920
rect 7460 1760 7500 1800
rect 1210 1370 1250 1410
rect 1430 1370 1470 1410
rect 1746 924 1768 930
rect 1768 924 1780 930
rect 1846 924 1858 930
rect 1858 924 1880 930
rect 1946 924 1948 930
rect 1948 924 1980 930
rect 1746 896 1780 924
rect 1846 896 1880 924
rect 1946 896 1980 924
rect 2046 896 2080 930
rect 2146 896 2180 930
rect 2246 924 2274 930
rect 2274 924 2280 930
rect 2246 896 2280 924
rect 1746 796 1780 830
rect 1846 796 1880 830
rect 1946 796 1980 830
rect 2046 796 2080 830
rect 2146 796 2180 830
rect 2246 796 2280 830
rect 1746 696 1780 730
rect 1846 696 1880 730
rect 1946 696 1980 730
rect 2046 696 2080 730
rect 2146 696 2180 730
rect 2246 696 2280 730
rect 1746 598 1780 630
rect 1846 598 1880 630
rect 1946 598 1980 630
rect 1746 596 1768 598
rect 1768 596 1780 598
rect 1846 596 1858 598
rect 1858 596 1880 598
rect 1946 596 1948 598
rect 1948 596 1980 598
rect 2046 596 2080 630
rect 2146 596 2180 630
rect 2246 598 2280 630
rect 2246 596 2274 598
rect 2274 596 2280 598
rect 1746 508 1780 530
rect 1846 508 1880 530
rect 1946 508 1980 530
rect 1746 496 1768 508
rect 1768 496 1780 508
rect 1846 496 1858 508
rect 1858 496 1880 508
rect 1946 496 1948 508
rect 1948 496 1980 508
rect 2046 496 2080 530
rect 2146 496 2180 530
rect 2246 508 2280 530
rect 2246 496 2274 508
rect 2274 496 2280 508
rect 1746 418 1780 430
rect 1846 418 1880 430
rect 1946 418 1980 430
rect 1746 396 1768 418
rect 1768 396 1780 418
rect 1846 396 1858 418
rect 1858 396 1880 418
rect 1946 396 1948 418
rect 1948 396 1980 418
rect 2046 396 2080 430
rect 2146 396 2180 430
rect 2246 418 2280 430
rect 2246 396 2274 418
rect 2274 396 2280 418
rect 3106 924 3128 930
rect 3128 924 3140 930
rect 3206 924 3218 930
rect 3218 924 3240 930
rect 3306 924 3308 930
rect 3308 924 3340 930
rect 3106 896 3140 924
rect 3206 896 3240 924
rect 3306 896 3340 924
rect 3406 896 3440 930
rect 3506 896 3540 930
rect 3606 924 3634 930
rect 3634 924 3640 930
rect 3606 896 3640 924
rect 3106 796 3140 830
rect 3206 796 3240 830
rect 3306 796 3340 830
rect 3406 796 3440 830
rect 3506 796 3540 830
rect 3606 796 3640 830
rect 3106 696 3140 730
rect 3206 696 3240 730
rect 3306 696 3340 730
rect 3406 696 3440 730
rect 3506 696 3540 730
rect 3606 696 3640 730
rect 3106 598 3140 630
rect 3206 598 3240 630
rect 3306 598 3340 630
rect 3106 596 3128 598
rect 3128 596 3140 598
rect 3206 596 3218 598
rect 3218 596 3240 598
rect 3306 596 3308 598
rect 3308 596 3340 598
rect 3406 596 3440 630
rect 3506 596 3540 630
rect 3606 598 3640 630
rect 3606 596 3634 598
rect 3634 596 3640 598
rect 3106 508 3140 530
rect 3206 508 3240 530
rect 3306 508 3340 530
rect 3106 496 3128 508
rect 3128 496 3140 508
rect 3206 496 3218 508
rect 3218 496 3240 508
rect 3306 496 3308 508
rect 3308 496 3340 508
rect 3406 496 3440 530
rect 3506 496 3540 530
rect 3606 508 3640 530
rect 3606 496 3634 508
rect 3634 496 3640 508
rect 3106 418 3140 430
rect 3206 418 3240 430
rect 3306 418 3340 430
rect 3106 396 3128 418
rect 3128 396 3140 418
rect 3206 396 3218 418
rect 3218 396 3240 418
rect 3306 396 3308 418
rect 3308 396 3340 418
rect 3406 396 3440 430
rect 3506 396 3540 430
rect 3606 418 3640 430
rect 3606 396 3634 418
rect 3634 396 3640 418
rect 4466 924 4488 930
rect 4488 924 4500 930
rect 4566 924 4578 930
rect 4578 924 4600 930
rect 4666 924 4668 930
rect 4668 924 4700 930
rect 4466 896 4500 924
rect 4566 896 4600 924
rect 4666 896 4700 924
rect 4766 896 4800 930
rect 4866 896 4900 930
rect 4966 924 4994 930
rect 4994 924 5000 930
rect 4966 896 5000 924
rect 4466 796 4500 830
rect 4566 796 4600 830
rect 4666 796 4700 830
rect 4766 796 4800 830
rect 4866 796 4900 830
rect 4966 796 5000 830
rect 4466 696 4500 730
rect 4566 696 4600 730
rect 4666 696 4700 730
rect 4766 696 4800 730
rect 4866 696 4900 730
rect 4966 696 5000 730
rect 4466 598 4500 630
rect 4566 598 4600 630
rect 4666 598 4700 630
rect 4466 596 4488 598
rect 4488 596 4500 598
rect 4566 596 4578 598
rect 4578 596 4600 598
rect 4666 596 4668 598
rect 4668 596 4700 598
rect 4766 596 4800 630
rect 4866 596 4900 630
rect 4966 598 5000 630
rect 4966 596 4994 598
rect 4994 596 5000 598
rect 4466 508 4500 530
rect 4566 508 4600 530
rect 4666 508 4700 530
rect 4466 496 4488 508
rect 4488 496 4500 508
rect 4566 496 4578 508
rect 4578 496 4600 508
rect 4666 496 4668 508
rect 4668 496 4700 508
rect 4766 496 4800 530
rect 4866 496 4900 530
rect 4966 508 5000 530
rect 4966 496 4994 508
rect 4994 496 5000 508
rect 4466 418 4500 430
rect 4566 418 4600 430
rect 4666 418 4700 430
rect 4466 396 4488 418
rect 4488 396 4500 418
rect 4566 396 4578 418
rect 4578 396 4600 418
rect 4666 396 4668 418
rect 4668 396 4700 418
rect 4766 396 4800 430
rect 4866 396 4900 430
rect 4966 418 5000 430
rect 4966 396 4994 418
rect 4994 396 5000 418
rect 5826 924 5848 930
rect 5848 924 5860 930
rect 5926 924 5938 930
rect 5938 924 5960 930
rect 6026 924 6028 930
rect 6028 924 6060 930
rect 5826 896 5860 924
rect 5926 896 5960 924
rect 6026 896 6060 924
rect 6126 896 6160 930
rect 6226 896 6260 930
rect 6326 924 6354 930
rect 6354 924 6360 930
rect 6326 896 6360 924
rect 5826 796 5860 830
rect 5926 796 5960 830
rect 6026 796 6060 830
rect 6126 796 6160 830
rect 6226 796 6260 830
rect 6326 796 6360 830
rect 5826 696 5860 730
rect 5926 696 5960 730
rect 6026 696 6060 730
rect 6126 696 6160 730
rect 6226 696 6260 730
rect 6326 696 6360 730
rect 5826 598 5860 630
rect 5926 598 5960 630
rect 6026 598 6060 630
rect 5826 596 5848 598
rect 5848 596 5860 598
rect 5926 596 5938 598
rect 5938 596 5960 598
rect 6026 596 6028 598
rect 6028 596 6060 598
rect 6126 596 6160 630
rect 6226 596 6260 630
rect 6326 598 6360 630
rect 6326 596 6354 598
rect 6354 596 6360 598
rect 5826 508 5860 530
rect 5926 508 5960 530
rect 6026 508 6060 530
rect 5826 496 5848 508
rect 5848 496 5860 508
rect 5926 496 5938 508
rect 5938 496 5960 508
rect 6026 496 6028 508
rect 6028 496 6060 508
rect 6126 496 6160 530
rect 6226 496 6260 530
rect 6326 508 6360 530
rect 6326 496 6354 508
rect 6354 496 6360 508
rect 5826 418 5860 430
rect 5926 418 5960 430
rect 6026 418 6060 430
rect 5826 396 5848 418
rect 5848 396 5860 418
rect 5926 396 5938 418
rect 5938 396 5960 418
rect 6026 396 6028 418
rect 6028 396 6060 418
rect 6126 396 6160 430
rect 6226 396 6260 430
rect 6326 418 6360 430
rect 6326 396 6354 418
rect 6354 396 6360 418
rect 7186 924 7208 930
rect 7208 924 7220 930
rect 7286 924 7298 930
rect 7298 924 7320 930
rect 7386 924 7388 930
rect 7388 924 7420 930
rect 7186 896 7220 924
rect 7286 896 7320 924
rect 7386 896 7420 924
rect 7486 896 7520 930
rect 7586 896 7620 930
rect 7686 924 7714 930
rect 7714 924 7720 930
rect 7686 896 7720 924
rect 7186 796 7220 830
rect 7286 796 7320 830
rect 7386 796 7420 830
rect 7486 796 7520 830
rect 7586 796 7620 830
rect 7686 796 7720 830
rect 7186 696 7220 730
rect 7286 696 7320 730
rect 7386 696 7420 730
rect 7486 696 7520 730
rect 7586 696 7620 730
rect 7686 696 7720 730
rect 7186 598 7220 630
rect 7286 598 7320 630
rect 7386 598 7420 630
rect 7186 596 7208 598
rect 7208 596 7220 598
rect 7286 596 7298 598
rect 7298 596 7320 598
rect 7386 596 7388 598
rect 7388 596 7420 598
rect 7486 596 7520 630
rect 7586 596 7620 630
rect 7686 598 7720 630
rect 7686 596 7714 598
rect 7714 596 7720 598
rect 7186 508 7220 530
rect 7286 508 7320 530
rect 7386 508 7420 530
rect 7186 496 7208 508
rect 7208 496 7220 508
rect 7286 496 7298 508
rect 7298 496 7320 508
rect 7386 496 7388 508
rect 7388 496 7420 508
rect 7486 496 7520 530
rect 7586 496 7620 530
rect 7686 508 7720 530
rect 7686 496 7714 508
rect 7714 496 7720 508
rect 7186 418 7220 430
rect 7286 418 7320 430
rect 7386 418 7420 430
rect 7186 396 7208 418
rect 7208 396 7220 418
rect 7286 396 7298 418
rect 7298 396 7320 418
rect 7386 396 7388 418
rect 7388 396 7420 418
rect 7486 396 7520 430
rect 7586 396 7620 430
rect 7686 418 7720 430
rect 7686 396 7714 418
rect 7714 396 7720 418
rect 8546 924 8568 930
rect 8568 924 8580 930
rect 8646 924 8658 930
rect 8658 924 8680 930
rect 8746 924 8748 930
rect 8748 924 8780 930
rect 8546 896 8580 924
rect 8646 896 8680 924
rect 8746 896 8780 924
rect 8846 896 8880 930
rect 8946 896 8980 930
rect 9046 924 9074 930
rect 9074 924 9080 930
rect 9046 896 9080 924
rect 8546 796 8580 830
rect 8646 796 8680 830
rect 8746 796 8780 830
rect 8846 796 8880 830
rect 8946 796 8980 830
rect 9046 796 9080 830
rect 8546 696 8580 730
rect 8646 696 8680 730
rect 8746 696 8780 730
rect 8846 696 8880 730
rect 8946 696 8980 730
rect 9046 696 9080 730
rect 8546 598 8580 630
rect 8646 598 8680 630
rect 8746 598 8780 630
rect 8546 596 8568 598
rect 8568 596 8580 598
rect 8646 596 8658 598
rect 8658 596 8680 598
rect 8746 596 8748 598
rect 8748 596 8780 598
rect 8846 596 8880 630
rect 8946 596 8980 630
rect 9046 598 9080 630
rect 9046 596 9074 598
rect 9074 596 9080 598
rect 8546 508 8580 530
rect 8646 508 8680 530
rect 8746 508 8780 530
rect 8546 496 8568 508
rect 8568 496 8580 508
rect 8646 496 8658 508
rect 8658 496 8680 508
rect 8746 496 8748 508
rect 8748 496 8780 508
rect 8846 496 8880 530
rect 8946 496 8980 530
rect 9046 508 9080 530
rect 9046 496 9074 508
rect 9074 496 9080 508
rect 8546 418 8580 430
rect 8646 418 8680 430
rect 8746 418 8780 430
rect 8546 396 8568 418
rect 8568 396 8580 418
rect 8646 396 8658 418
rect 8658 396 8680 418
rect 8746 396 8748 418
rect 8748 396 8780 418
rect 8846 396 8880 430
rect 8946 396 8980 430
rect 9046 418 9080 430
rect 9046 396 9074 418
rect 9074 396 9080 418
rect 40 50 80 90
rect 220 50 260 90
rect 400 50 440 90
rect 580 50 620 90
rect 760 50 800 90
rect 940 50 980 90
rect 1120 50 1160 90
rect 1300 50 1340 90
rect 1480 58 1506 90
rect 1506 58 1520 90
rect 1660 58 1686 90
rect 1686 58 1700 90
rect 1840 58 1866 90
rect 1866 58 1880 90
rect 2020 58 2046 90
rect 2046 58 2060 90
rect 2200 58 2226 90
rect 2226 58 2240 90
rect 2380 58 2406 90
rect 2406 58 2420 90
rect 1480 50 1520 58
rect 1660 50 1700 58
rect 1840 50 1880 58
rect 2020 50 2060 58
rect 2200 50 2240 58
rect 2380 50 2420 58
rect 2560 50 2600 90
rect 2740 50 2780 90
rect 2920 58 2956 90
rect 2956 58 2960 90
rect 3100 58 3136 90
rect 3136 58 3140 90
rect 3280 58 3316 90
rect 3316 58 3320 90
rect 3460 58 3496 90
rect 3496 58 3500 90
rect 3640 58 3676 90
rect 3676 58 3680 90
rect 3820 58 3856 90
rect 3856 58 3860 90
rect 2920 50 2960 58
rect 3100 50 3140 58
rect 3280 50 3320 58
rect 3460 50 3500 58
rect 3640 50 3680 58
rect 3820 50 3860 58
rect 4000 50 4040 90
rect 4180 50 4220 90
rect 4360 50 4400 90
rect 4540 50 4580 90
rect 4720 50 4760 90
rect 4900 50 4940 90
rect 5080 50 5120 90
rect 5260 50 5300 90
rect 5440 50 5480 90
rect 5620 50 5660 90
rect 5800 50 5840 90
rect 5980 50 6020 90
rect 6160 50 6200 90
rect 6340 50 6380 90
rect 6520 50 6560 90
rect 6700 50 6740 90
rect 6880 50 6920 90
rect 7060 58 7070 90
rect 7070 58 7100 90
rect 7240 58 7250 90
rect 7250 58 7280 90
rect 7420 58 7430 90
rect 7430 58 7460 90
rect 7600 58 7610 90
rect 7610 58 7640 90
rect 7780 58 7790 90
rect 7790 58 7820 90
rect 7960 58 7970 90
rect 7970 58 8000 90
rect 7060 50 7100 58
rect 7240 50 7280 58
rect 7420 50 7460 58
rect 7600 50 7640 58
rect 7780 50 7820 58
rect 7960 50 8000 58
rect 8140 50 8180 90
rect 8320 58 8340 90
rect 8340 58 8360 90
rect 8500 58 8520 90
rect 8520 58 8540 90
rect 8680 58 8700 90
rect 8700 58 8720 90
rect 8860 58 8880 90
rect 8880 58 8900 90
rect 9040 58 9060 90
rect 9060 58 9080 90
rect 9220 58 9240 90
rect 9240 58 9260 90
rect 8320 50 8360 58
rect 8500 50 8540 58
rect 8680 50 8720 58
rect 8860 50 8900 58
rect 9040 50 9080 58
rect 9220 50 9260 58
rect 9400 50 9440 90
<< metal1 >>
rect 4620 5540 4700 5550
rect 4620 5480 4630 5540
rect 4690 5480 4700 5540
rect 4620 5470 4700 5480
rect 5020 5540 5100 5550
rect 5020 5480 5030 5540
rect 5090 5480 5100 5540
rect 5020 5470 5100 5480
rect 5420 5540 5500 5550
rect 5420 5480 5430 5540
rect 5490 5480 5500 5540
rect 5420 5470 5500 5480
rect 5820 5540 5900 5550
rect 5820 5480 5830 5540
rect 5890 5480 5900 5540
rect 5820 5470 5900 5480
rect 6220 5540 6300 5550
rect 6220 5480 6230 5540
rect 6290 5480 6300 5540
rect 6220 5470 6300 5480
rect 6620 5540 6700 5550
rect 6620 5480 6630 5540
rect 6690 5480 6700 5540
rect 6620 5470 6700 5480
rect 7020 5540 7100 5550
rect 7020 5480 7030 5540
rect 7090 5480 7100 5540
rect 7020 5470 7100 5480
rect 7420 5540 7500 5550
rect 7420 5480 7430 5540
rect 7490 5480 7500 5540
rect 7420 5470 7500 5480
rect 7820 5540 7900 5550
rect 7820 5480 7830 5540
rect 7890 5480 7900 5540
rect 7820 5470 7900 5480
rect 8220 5540 8300 5550
rect 8220 5480 8230 5540
rect 8290 5480 8300 5540
rect 8220 5470 8300 5480
rect 1190 5020 1270 5030
rect 1190 4960 1200 5020
rect 1260 4960 1270 5020
rect 1190 4020 1270 4960
rect 1890 5020 1970 5030
rect 1890 4960 1900 5020
rect 1960 4960 1970 5020
rect 1890 4950 1970 4960
rect 4300 4600 4380 4610
rect 4300 4540 4310 4600
rect 4370 4540 4380 4600
rect 4300 4530 4380 4540
rect 4820 4600 4900 4610
rect 4820 4540 4830 4600
rect 4890 4540 4900 4600
rect 4820 4530 4900 4540
rect 6220 4590 6300 4610
rect 6220 4550 6240 4590
rect 6280 4550 6300 4590
rect 6220 4530 6300 4550
rect 6620 4590 6700 4610
rect 6620 4550 6640 4590
rect 6680 4550 6700 4590
rect 6620 4530 6700 4550
rect 6820 4600 6900 4610
rect 6820 4540 6830 4600
rect 6890 4540 6900 4600
rect 6820 4530 6900 4540
rect 7620 4600 7700 4610
rect 7620 4540 7630 4600
rect 7690 4540 7700 4600
rect 7620 4530 7700 4540
rect 8140 4600 8220 4610
rect 8140 4540 8150 4600
rect 8210 4540 8220 4600
rect 8140 4530 8220 4540
rect 8750 4600 8830 4610
rect 8750 4540 8760 4600
rect 8820 4540 8830 4600
rect 8750 4530 8830 4540
rect 3790 4430 4230 4440
rect 3790 4370 3800 4430
rect 4220 4370 4230 4430
rect 3790 4360 4230 4370
rect 1190 3960 1200 4020
rect 1260 3960 1270 4020
rect 880 3430 960 3440
rect 880 3370 890 3430
rect 950 3370 960 3430
rect 880 1450 960 3370
rect 360 370 960 1450
rect 1190 1410 1270 3960
rect 1890 4020 1970 4030
rect 1890 3960 1900 4020
rect 1960 3960 1970 4020
rect 1890 3950 1970 3960
rect 3790 3430 4230 3440
rect 4320 3430 4360 4530
rect 5220 4510 5300 4520
rect 5220 4450 5230 4510
rect 5290 4450 5300 4510
rect 5220 4440 5300 4450
rect 6020 4510 6100 4520
rect 6020 4450 6030 4510
rect 6090 4450 6100 4510
rect 6020 4440 6100 4450
rect 5620 4420 5700 4430
rect 5620 4360 5630 4420
rect 5690 4360 5700 4420
rect 5620 4350 5700 4360
rect 6240 4240 6280 4530
rect 6420 4420 6500 4430
rect 6420 4360 6430 4420
rect 6490 4360 6500 4420
rect 6420 4350 6500 4360
rect 6640 4240 6680 4530
rect 8020 4510 8100 4520
rect 8020 4450 8030 4510
rect 8090 4450 8100 4510
rect 8020 4440 8100 4450
rect 8630 4510 8710 4520
rect 8630 4450 8640 4510
rect 8700 4450 8710 4510
rect 8630 4440 8710 4450
rect 7220 4420 7300 4430
rect 7220 4360 7230 4420
rect 7290 4360 7300 4420
rect 7220 4350 7300 4360
rect 4460 4230 4540 4240
rect 4460 4170 4470 4230
rect 4530 4170 4540 4230
rect 4460 4160 4540 4170
rect 4660 4230 4740 4240
rect 4660 4170 4670 4230
rect 4730 4170 4740 4230
rect 4660 4160 4740 4170
rect 5060 4230 5140 4240
rect 5060 4170 5070 4230
rect 5130 4170 5140 4230
rect 5060 4160 5140 4170
rect 5460 4230 5540 4240
rect 5460 4170 5470 4230
rect 5530 4170 5540 4230
rect 5460 4160 5540 4170
rect 5660 4230 5740 4240
rect 5660 4170 5670 4230
rect 5730 4170 5740 4230
rect 5660 4160 5740 4170
rect 5820 4230 5900 4240
rect 5820 4170 5830 4230
rect 5890 4170 5900 4230
rect 5820 4160 5900 4170
rect 6020 4230 6100 4240
rect 6020 4170 6030 4230
rect 6090 4170 6100 4230
rect 6020 4160 6100 4170
rect 6220 4220 6300 4240
rect 6220 4180 6240 4220
rect 6280 4180 6300 4220
rect 6220 4160 6300 4180
rect 6420 4230 6500 4240
rect 6420 4170 6430 4230
rect 6490 4170 6500 4230
rect 6420 4160 6500 4170
rect 6620 4220 6700 4240
rect 6620 4180 6640 4220
rect 6680 4180 6700 4220
rect 6620 4160 6700 4180
rect 6820 4230 6900 4240
rect 6820 4170 6830 4230
rect 6890 4170 6900 4230
rect 6820 4160 6900 4170
rect 7020 4230 7100 4240
rect 7020 4170 7030 4230
rect 7090 4170 7100 4230
rect 7020 4160 7100 4170
rect 7180 4230 7260 4240
rect 7180 4170 7190 4230
rect 7250 4170 7260 4230
rect 7180 4160 7260 4170
rect 7380 4230 7460 4240
rect 7380 4170 7390 4230
rect 7450 4170 7460 4230
rect 7380 4160 7460 4170
rect 7780 4230 7860 4240
rect 7780 4170 7790 4230
rect 7850 4170 7860 4230
rect 7780 4160 7860 4170
rect 8180 4230 8260 4240
rect 8180 4170 8190 4230
rect 8250 4170 8260 4230
rect 8180 4160 8260 4170
rect 8380 4230 8460 4240
rect 8380 4170 8390 4230
rect 8450 4170 8460 4230
rect 8380 4160 8460 4170
rect 5260 3690 5340 3700
rect 5260 3630 5270 3690
rect 5330 3630 5340 3690
rect 5260 3620 5340 3630
rect 5940 3690 6020 3700
rect 5940 3630 5950 3690
rect 6010 3630 6020 3690
rect 5940 3620 6020 3630
rect 6420 3680 6500 3700
rect 6420 3640 6440 3680
rect 6480 3640 6500 3680
rect 6420 3620 6500 3640
rect 6900 3690 6980 3700
rect 6900 3630 6910 3690
rect 6970 3630 6980 3690
rect 6900 3620 6980 3630
rect 7580 3690 7660 3700
rect 7580 3630 7590 3690
rect 7650 3630 7660 3690
rect 7580 3620 7660 3630
rect 4860 3600 4940 3610
rect 4860 3540 4870 3600
rect 4930 3540 4940 3600
rect 4860 3530 4940 3540
rect 5540 3600 5620 3610
rect 5540 3540 5550 3600
rect 5610 3540 5620 3600
rect 5540 3530 5620 3540
rect 5560 3430 5600 3530
rect 5960 3430 6000 3620
rect 6120 3600 6200 3610
rect 6120 3540 6130 3600
rect 6190 3540 6200 3600
rect 6120 3530 6200 3540
rect 6440 3520 6480 3620
rect 6720 3600 6800 3610
rect 6720 3540 6730 3600
rect 6790 3540 6800 3600
rect 6720 3530 6800 3540
rect 6420 3510 6500 3520
rect 6420 3450 6430 3510
rect 6490 3450 6500 3510
rect 6420 3440 6500 3450
rect 6920 3430 6960 3620
rect 7300 3600 7380 3610
rect 7300 3540 7310 3600
rect 7370 3540 7380 3600
rect 7300 3530 7380 3540
rect 7980 3600 8060 3610
rect 7980 3540 7990 3600
rect 8050 3540 8060 3600
rect 7980 3530 8060 3540
rect 7320 3430 7360 3530
rect 7840 3510 7920 3520
rect 7840 3450 7850 3510
rect 7910 3450 7920 3510
rect 7840 3440 7920 3450
rect 3790 3370 3800 3430
rect 4220 3370 4230 3430
rect 3790 3360 4230 3370
rect 4300 3420 4380 3430
rect 4300 3360 4310 3420
rect 4370 3360 4380 3420
rect 4300 3350 4380 3360
rect 5540 3410 5620 3430
rect 5540 3370 5560 3410
rect 5600 3370 5620 3410
rect 5540 3350 5620 3370
rect 5940 3410 6020 3430
rect 5940 3370 5960 3410
rect 6000 3370 6020 3410
rect 5940 3350 6020 3370
rect 6060 3420 6140 3430
rect 6060 3360 6070 3420
rect 6130 3360 6140 3420
rect 6060 3350 6140 3360
rect 6780 3420 6860 3430
rect 6780 3360 6790 3420
rect 6850 3360 6860 3420
rect 6780 3350 6860 3360
rect 6900 3410 6980 3430
rect 6900 3370 6920 3410
rect 6960 3370 6980 3410
rect 6900 3350 6980 3370
rect 7300 3410 7380 3430
rect 7300 3370 7320 3410
rect 7360 3370 7380 3410
rect 7300 3350 7380 3370
rect 5540 3080 5620 3090
rect 1720 3070 1800 3080
rect 1720 3010 1730 3070
rect 1790 3010 1800 3070
rect 1190 1370 1210 1410
rect 1250 1370 1270 1410
rect 1190 1340 1270 1370
rect 1410 2480 1490 2490
rect 1410 2420 1420 2480
rect 1480 2420 1490 2480
rect 1410 1410 1490 2420
rect 1410 1370 1430 1410
rect 1470 1370 1490 1410
rect 1410 1340 1490 1370
rect 1720 1460 1800 3010
rect 1890 3070 1970 3080
rect 1890 3010 1900 3070
rect 1960 3010 1970 3070
rect 1890 3000 1970 3010
rect 3790 3070 4230 3080
rect 3790 3010 3800 3070
rect 4220 3010 4230 3070
rect 5540 3020 5550 3080
rect 5610 3020 5620 3080
rect 5540 3010 5620 3020
rect 7300 3080 7380 3090
rect 7300 3020 7310 3080
rect 7370 3020 7380 3080
rect 7300 3010 7380 3020
rect 3790 3000 4230 3010
rect 5140 2990 5220 3000
rect 5140 2930 5150 2990
rect 5210 2930 5220 2990
rect 5140 2920 5220 2930
rect 5340 2990 5420 3000
rect 5340 2930 5350 2990
rect 5410 2930 5420 2990
rect 5340 2920 5420 2930
rect 5740 2990 5820 3000
rect 5740 2930 5750 2990
rect 5810 2930 5820 2990
rect 5740 2920 5820 2930
rect 6140 2990 6220 3000
rect 6140 2930 6150 2990
rect 6210 2930 6220 2990
rect 6140 2920 6220 2930
rect 6340 2990 6420 3000
rect 6340 2930 6350 2990
rect 6410 2930 6420 2990
rect 6340 2920 6420 2930
rect 6500 2990 6580 3000
rect 6500 2930 6510 2990
rect 6570 2930 6580 2990
rect 6500 2920 6580 2930
rect 6700 2990 6780 3000
rect 6700 2930 6710 2990
rect 6770 2930 6780 2990
rect 6700 2920 6780 2930
rect 7100 2990 7180 3000
rect 7100 2930 7110 2990
rect 7170 2930 7180 2990
rect 7100 2920 7180 2930
rect 7500 2990 7580 3000
rect 7500 2930 7510 2990
rect 7570 2930 7580 2990
rect 7500 2920 7580 2930
rect 7700 2990 7780 3000
rect 7700 2930 7710 2990
rect 7770 2930 7780 2990
rect 7700 2920 7780 2930
rect 7860 2880 7900 3440
rect 8650 3090 8690 4440
rect 8770 4340 8810 4530
rect 8750 4320 8830 4340
rect 8750 4280 8770 4320
rect 8810 4280 8830 4320
rect 8750 4260 8830 4280
rect 9150 4230 9230 4240
rect 9150 4170 9160 4230
rect 9220 4170 9230 4230
rect 9150 4160 9230 4170
rect 8970 3650 9050 3670
rect 8970 3610 8990 3650
rect 9030 3610 9050 3650
rect 8970 3590 9050 3610
rect 8860 3420 8940 3430
rect 8860 3360 8870 3420
rect 8930 3360 8940 3420
rect 8860 3350 8940 3360
rect 8630 3080 8710 3090
rect 8630 3020 8640 3080
rect 8700 3020 8710 3080
rect 8630 3010 8710 3020
rect 7300 2870 7380 2880
rect 7300 2810 7310 2870
rect 7370 2810 7380 2870
rect 7300 2800 7380 2810
rect 7840 2870 7920 2880
rect 7840 2810 7850 2870
rect 7910 2810 7920 2870
rect 7840 2800 7920 2810
rect 1890 2480 1970 2490
rect 1890 2420 1900 2480
rect 1960 2420 1970 2480
rect 1890 2410 1970 2420
rect 4660 1930 4740 1940
rect 4660 1870 4670 1930
rect 4730 1870 4740 1930
rect 4660 1860 4740 1870
rect 6420 1930 6500 1940
rect 6420 1870 6430 1930
rect 6490 1870 6500 1930
rect 6420 1860 6500 1870
rect 8180 1930 8260 1940
rect 8180 1870 8190 1930
rect 8250 1870 8260 1930
rect 8180 1860 8260 1870
rect 9010 1820 9050 3590
rect 7440 1810 7520 1820
rect 7440 1750 7450 1810
rect 7510 1750 7520 1810
rect 7440 1740 7520 1750
rect 8990 1810 9070 1820
rect 8990 1750 9000 1810
rect 9060 1750 9070 1810
rect 8990 1740 9070 1750
rect 1720 1420 9120 1460
rect 1720 975 2320 1420
rect 3080 975 3680 1420
rect 4440 975 5040 1420
rect 5800 975 6400 1420
rect 7160 975 7760 1420
rect 8520 975 9120 1420
rect 1715 930 2325 975
rect 1715 896 1746 930
rect 1780 896 1846 930
rect 1880 896 1946 930
rect 1980 896 2046 930
rect 2080 896 2146 930
rect 2180 896 2246 930
rect 2280 896 2325 930
rect 1715 830 2325 896
rect 1715 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2325 830
rect 1715 730 2325 796
rect 1715 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2325 730
rect 1715 630 2325 696
rect 1715 596 1746 630
rect 1780 596 1846 630
rect 1880 596 1946 630
rect 1980 596 2046 630
rect 2080 596 2146 630
rect 2180 596 2246 630
rect 2280 596 2325 630
rect 1715 530 2325 596
rect 1715 496 1746 530
rect 1780 496 1846 530
rect 1880 496 1946 530
rect 1980 496 2046 530
rect 2080 496 2146 530
rect 2180 496 2246 530
rect 2280 496 2325 530
rect 1715 430 2325 496
rect 1715 396 1746 430
rect 1780 396 1846 430
rect 1880 396 1946 430
rect 1980 396 2046 430
rect 2080 396 2146 430
rect 2180 396 2246 430
rect 2280 396 2325 430
rect 1715 365 2325 396
rect 3075 930 3685 975
rect 3075 896 3106 930
rect 3140 896 3206 930
rect 3240 896 3306 930
rect 3340 896 3406 930
rect 3440 896 3506 930
rect 3540 896 3606 930
rect 3640 896 3685 930
rect 3075 830 3685 896
rect 3075 796 3106 830
rect 3140 796 3206 830
rect 3240 796 3306 830
rect 3340 796 3406 830
rect 3440 796 3506 830
rect 3540 796 3606 830
rect 3640 796 3685 830
rect 3075 730 3685 796
rect 3075 696 3106 730
rect 3140 696 3206 730
rect 3240 696 3306 730
rect 3340 696 3406 730
rect 3440 696 3506 730
rect 3540 696 3606 730
rect 3640 696 3685 730
rect 3075 630 3685 696
rect 3075 596 3106 630
rect 3140 596 3206 630
rect 3240 596 3306 630
rect 3340 596 3406 630
rect 3440 596 3506 630
rect 3540 596 3606 630
rect 3640 596 3685 630
rect 3075 530 3685 596
rect 3075 496 3106 530
rect 3140 496 3206 530
rect 3240 496 3306 530
rect 3340 496 3406 530
rect 3440 496 3506 530
rect 3540 496 3606 530
rect 3640 496 3685 530
rect 3075 430 3685 496
rect 3075 396 3106 430
rect 3140 396 3206 430
rect 3240 396 3306 430
rect 3340 396 3406 430
rect 3440 396 3506 430
rect 3540 396 3606 430
rect 3640 396 3685 430
rect 3075 365 3685 396
rect 4435 930 5045 975
rect 4435 896 4466 930
rect 4500 896 4566 930
rect 4600 896 4666 930
rect 4700 896 4766 930
rect 4800 896 4866 930
rect 4900 896 4966 930
rect 5000 896 5045 930
rect 4435 830 5045 896
rect 4435 796 4466 830
rect 4500 796 4566 830
rect 4600 796 4666 830
rect 4700 796 4766 830
rect 4800 796 4866 830
rect 4900 796 4966 830
rect 5000 796 5045 830
rect 4435 730 5045 796
rect 4435 696 4466 730
rect 4500 696 4566 730
rect 4600 696 4666 730
rect 4700 696 4766 730
rect 4800 696 4866 730
rect 4900 696 4966 730
rect 5000 696 5045 730
rect 4435 630 5045 696
rect 4435 596 4466 630
rect 4500 596 4566 630
rect 4600 596 4666 630
rect 4700 596 4766 630
rect 4800 596 4866 630
rect 4900 596 4966 630
rect 5000 596 5045 630
rect 4435 530 5045 596
rect 4435 496 4466 530
rect 4500 496 4566 530
rect 4600 496 4666 530
rect 4700 496 4766 530
rect 4800 496 4866 530
rect 4900 496 4966 530
rect 5000 496 5045 530
rect 4435 430 5045 496
rect 4435 396 4466 430
rect 4500 396 4566 430
rect 4600 396 4666 430
rect 4700 396 4766 430
rect 4800 396 4866 430
rect 4900 396 4966 430
rect 5000 396 5045 430
rect 4435 365 5045 396
rect 5795 930 6405 975
rect 5795 896 5826 930
rect 5860 896 5926 930
rect 5960 896 6026 930
rect 6060 896 6126 930
rect 6160 896 6226 930
rect 6260 896 6326 930
rect 6360 896 6405 930
rect 5795 830 6405 896
rect 5795 796 5826 830
rect 5860 796 5926 830
rect 5960 796 6026 830
rect 6060 796 6126 830
rect 6160 796 6226 830
rect 6260 796 6326 830
rect 6360 796 6405 830
rect 5795 730 6405 796
rect 5795 696 5826 730
rect 5860 696 5926 730
rect 5960 696 6026 730
rect 6060 696 6126 730
rect 6160 696 6226 730
rect 6260 696 6326 730
rect 6360 696 6405 730
rect 5795 630 6405 696
rect 5795 596 5826 630
rect 5860 596 5926 630
rect 5960 596 6026 630
rect 6060 596 6126 630
rect 6160 596 6226 630
rect 6260 596 6326 630
rect 6360 596 6405 630
rect 5795 530 6405 596
rect 5795 496 5826 530
rect 5860 496 5926 530
rect 5960 496 6026 530
rect 6060 496 6126 530
rect 6160 496 6226 530
rect 6260 496 6326 530
rect 6360 496 6405 530
rect 5795 430 6405 496
rect 5795 396 5826 430
rect 5860 396 5926 430
rect 5960 396 6026 430
rect 6060 396 6126 430
rect 6160 396 6226 430
rect 6260 396 6326 430
rect 6360 396 6405 430
rect 5795 365 6405 396
rect 7155 930 7765 975
rect 7155 896 7186 930
rect 7220 896 7286 930
rect 7320 896 7386 930
rect 7420 896 7486 930
rect 7520 896 7586 930
rect 7620 896 7686 930
rect 7720 896 7765 930
rect 7155 830 7765 896
rect 7155 796 7186 830
rect 7220 796 7286 830
rect 7320 796 7386 830
rect 7420 796 7486 830
rect 7520 796 7586 830
rect 7620 796 7686 830
rect 7720 796 7765 830
rect 7155 730 7765 796
rect 7155 696 7186 730
rect 7220 696 7286 730
rect 7320 696 7386 730
rect 7420 696 7486 730
rect 7520 696 7586 730
rect 7620 696 7686 730
rect 7720 696 7765 730
rect 7155 630 7765 696
rect 7155 596 7186 630
rect 7220 596 7286 630
rect 7320 596 7386 630
rect 7420 596 7486 630
rect 7520 596 7586 630
rect 7620 596 7686 630
rect 7720 596 7765 630
rect 7155 530 7765 596
rect 7155 496 7186 530
rect 7220 496 7286 530
rect 7320 496 7386 530
rect 7420 496 7486 530
rect 7520 496 7586 530
rect 7620 496 7686 530
rect 7720 496 7765 530
rect 7155 430 7765 496
rect 7155 396 7186 430
rect 7220 396 7286 430
rect 7320 396 7386 430
rect 7420 396 7486 430
rect 7520 396 7586 430
rect 7620 396 7686 430
rect 7720 396 7765 430
rect 7155 365 7765 396
rect 8515 930 9125 975
rect 8515 896 8546 930
rect 8580 896 8646 930
rect 8680 896 8746 930
rect 8780 896 8846 930
rect 8880 896 8946 930
rect 8980 896 9046 930
rect 9080 896 9125 930
rect 8515 830 9125 896
rect 8515 796 8546 830
rect 8580 796 8646 830
rect 8680 796 8746 830
rect 8780 796 8846 830
rect 8880 796 8946 830
rect 8980 796 9046 830
rect 9080 796 9125 830
rect 8515 730 9125 796
rect 8515 696 8546 730
rect 8580 696 8646 730
rect 8680 696 8746 730
rect 8780 696 8846 730
rect 8880 696 8946 730
rect 8980 696 9046 730
rect 9080 696 9125 730
rect 8515 630 9125 696
rect 8515 596 8546 630
rect 8580 596 8646 630
rect 8680 596 8746 630
rect 8780 596 8846 630
rect 8880 596 8946 630
rect 8980 596 9046 630
rect 9080 596 9125 630
rect 8515 530 9125 596
rect 8515 496 8546 530
rect 8580 496 8646 530
rect 8680 496 8746 530
rect 8780 496 8846 530
rect 8880 496 8946 530
rect 8980 496 9046 530
rect 9080 496 9125 530
rect 8515 430 9125 496
rect 8515 396 8546 430
rect 8580 396 8646 430
rect 8680 396 8746 430
rect 8780 396 8846 430
rect 8880 396 8946 430
rect 8980 396 9046 430
rect 9080 396 9125 430
rect 8515 365 9125 396
rect 10 100 110 120
rect 10 40 30 100
rect 90 40 110 100
rect 10 20 110 40
rect 190 100 290 120
rect 190 40 210 100
rect 270 40 290 100
rect 190 20 290 40
rect 370 100 470 120
rect 370 40 390 100
rect 450 40 470 100
rect 370 20 470 40
rect 550 100 650 120
rect 550 40 570 100
rect 630 40 650 100
rect 550 20 650 40
rect 730 100 830 120
rect 730 40 750 100
rect 810 40 830 100
rect 730 20 830 40
rect 910 100 1010 120
rect 910 40 930 100
rect 990 40 1010 100
rect 910 20 1010 40
rect 1090 100 1190 120
rect 1090 40 1110 100
rect 1170 40 1190 100
rect 1090 20 1190 40
rect 1270 100 1370 120
rect 1270 40 1290 100
rect 1350 40 1370 100
rect 1270 20 1370 40
rect 1450 100 1550 120
rect 1450 40 1470 100
rect 1530 40 1550 100
rect 1450 20 1550 40
rect 1630 100 1730 120
rect 1630 40 1650 100
rect 1710 40 1730 100
rect 1630 20 1730 40
rect 1810 100 1910 120
rect 1810 40 1830 100
rect 1890 40 1910 100
rect 1810 20 1910 40
rect 1990 100 2090 120
rect 1990 40 2010 100
rect 2070 40 2090 100
rect 1990 20 2090 40
rect 2170 100 2270 120
rect 2170 40 2190 100
rect 2250 40 2270 100
rect 2170 20 2270 40
rect 2350 100 2450 120
rect 2350 40 2370 100
rect 2430 40 2450 100
rect 2350 20 2450 40
rect 2530 100 2630 120
rect 2530 40 2550 100
rect 2610 40 2630 100
rect 2530 20 2630 40
rect 2710 100 2810 120
rect 2710 40 2730 100
rect 2790 40 2810 100
rect 2710 20 2810 40
rect 2890 100 2990 120
rect 2890 40 2910 100
rect 2970 40 2990 100
rect 2890 20 2990 40
rect 3070 100 3170 120
rect 3070 40 3090 100
rect 3150 40 3170 100
rect 3070 20 3170 40
rect 3250 100 3350 120
rect 3250 40 3270 100
rect 3330 40 3350 100
rect 3250 20 3350 40
rect 3430 100 3530 120
rect 3430 40 3450 100
rect 3510 40 3530 100
rect 3430 20 3530 40
rect 3610 100 3710 120
rect 3610 40 3630 100
rect 3690 40 3710 100
rect 3610 20 3710 40
rect 3790 100 3890 120
rect 3790 40 3810 100
rect 3870 40 3890 100
rect 3790 20 3890 40
rect 3970 100 4070 120
rect 3970 40 3990 100
rect 4050 40 4070 100
rect 3970 20 4070 40
rect 4150 100 4250 120
rect 4150 40 4170 100
rect 4230 40 4250 100
rect 4150 20 4250 40
rect 4330 100 4430 120
rect 4330 40 4350 100
rect 4410 40 4430 100
rect 4330 20 4430 40
rect 4510 100 4610 120
rect 4510 40 4530 100
rect 4590 40 4610 100
rect 4510 20 4610 40
rect 4690 100 4790 120
rect 4690 40 4710 100
rect 4770 40 4790 100
rect 4690 20 4790 40
rect 4870 100 4970 120
rect 4870 40 4890 100
rect 4950 40 4970 100
rect 4870 20 4970 40
rect 5050 100 5150 120
rect 5050 40 5070 100
rect 5130 40 5150 100
rect 5050 20 5150 40
rect 5230 100 5330 120
rect 5230 40 5250 100
rect 5310 40 5330 100
rect 5230 20 5330 40
rect 5410 100 5510 120
rect 5410 40 5430 100
rect 5490 40 5510 100
rect 5410 20 5510 40
rect 5590 100 5690 120
rect 5590 40 5610 100
rect 5670 40 5690 100
rect 5590 20 5690 40
rect 5770 100 5870 120
rect 5770 40 5790 100
rect 5850 40 5870 100
rect 5770 20 5870 40
rect 5950 100 6050 120
rect 5950 40 5970 100
rect 6030 40 6050 100
rect 5950 20 6050 40
rect 6130 100 6230 120
rect 6130 40 6150 100
rect 6210 40 6230 100
rect 6130 20 6230 40
rect 6310 100 6410 120
rect 6310 40 6330 100
rect 6390 40 6410 100
rect 6310 20 6410 40
rect 6490 100 6590 120
rect 6490 40 6510 100
rect 6570 40 6590 100
rect 6490 20 6590 40
rect 6670 100 6770 120
rect 6670 40 6690 100
rect 6750 40 6770 100
rect 6670 20 6770 40
rect 6850 100 6950 120
rect 6850 40 6870 100
rect 6930 40 6950 100
rect 6850 20 6950 40
rect 7030 100 7130 120
rect 7030 40 7050 100
rect 7110 40 7130 100
rect 7030 20 7130 40
rect 7210 100 7310 120
rect 7210 40 7230 100
rect 7290 40 7310 100
rect 7210 20 7310 40
rect 7390 100 7490 120
rect 7390 40 7410 100
rect 7470 40 7490 100
rect 7390 20 7490 40
rect 7570 100 7670 120
rect 7570 40 7590 100
rect 7650 40 7670 100
rect 7570 20 7670 40
rect 7750 100 7850 120
rect 7750 40 7770 100
rect 7830 40 7850 100
rect 7750 20 7850 40
rect 7930 100 8030 120
rect 7930 40 7950 100
rect 8010 40 8030 100
rect 7930 20 8030 40
rect 8110 100 8210 120
rect 8110 40 8130 100
rect 8190 40 8210 100
rect 8110 20 8210 40
rect 8290 100 8390 120
rect 8290 40 8310 100
rect 8370 40 8390 100
rect 8290 20 8390 40
rect 8470 100 8570 120
rect 8470 40 8490 100
rect 8550 40 8570 100
rect 8470 20 8570 40
rect 8650 100 8750 120
rect 8650 40 8670 100
rect 8730 40 8750 100
rect 8650 20 8750 40
rect 8830 100 8930 120
rect 8830 40 8850 100
rect 8910 40 8930 100
rect 8830 20 8930 40
rect 9010 100 9110 120
rect 9010 40 9030 100
rect 9090 40 9110 100
rect 9010 20 9110 40
rect 9190 100 9290 120
rect 9190 40 9210 100
rect 9270 40 9290 100
rect 9190 20 9290 40
rect 9370 100 9470 120
rect 9370 40 9390 100
rect 9450 40 9470 100
rect 9370 20 9470 40
<< via1 >>
rect 4630 5530 4690 5540
rect 4630 5490 4640 5530
rect 4640 5490 4680 5530
rect 4680 5490 4690 5530
rect 4630 5480 4690 5490
rect 5030 5530 5090 5540
rect 5030 5490 5040 5530
rect 5040 5490 5080 5530
rect 5080 5490 5090 5530
rect 5030 5480 5090 5490
rect 5430 5530 5490 5540
rect 5430 5490 5440 5530
rect 5440 5490 5480 5530
rect 5480 5490 5490 5530
rect 5430 5480 5490 5490
rect 5830 5530 5890 5540
rect 5830 5490 5840 5530
rect 5840 5490 5880 5530
rect 5880 5490 5890 5530
rect 5830 5480 5890 5490
rect 6230 5530 6290 5540
rect 6230 5490 6240 5530
rect 6240 5490 6280 5530
rect 6280 5490 6290 5530
rect 6230 5480 6290 5490
rect 6630 5530 6690 5540
rect 6630 5490 6640 5530
rect 6640 5490 6680 5530
rect 6680 5490 6690 5530
rect 6630 5480 6690 5490
rect 7030 5530 7090 5540
rect 7030 5490 7040 5530
rect 7040 5490 7080 5530
rect 7080 5490 7090 5530
rect 7030 5480 7090 5490
rect 7430 5530 7490 5540
rect 7430 5490 7440 5530
rect 7440 5490 7480 5530
rect 7480 5490 7490 5530
rect 7430 5480 7490 5490
rect 7830 5530 7890 5540
rect 7830 5490 7840 5530
rect 7840 5490 7880 5530
rect 7880 5490 7890 5530
rect 7830 5480 7890 5490
rect 8230 5530 8290 5540
rect 8230 5490 8240 5530
rect 8240 5490 8280 5530
rect 8280 5490 8290 5530
rect 8230 5480 8290 5490
rect 1200 4960 1260 5020
rect 1900 5010 1960 5020
rect 1900 4970 1910 5010
rect 1910 4970 1950 5010
rect 1950 4970 1960 5010
rect 1900 4960 1960 4970
rect 4310 4540 4370 4600
rect 4830 4590 4890 4600
rect 4830 4550 4840 4590
rect 4840 4550 4880 4590
rect 4880 4550 4890 4590
rect 4830 4540 4890 4550
rect 6830 4590 6890 4600
rect 6830 4550 6840 4590
rect 6840 4550 6880 4590
rect 6880 4550 6890 4590
rect 6830 4540 6890 4550
rect 7630 4590 7690 4600
rect 7630 4550 7640 4590
rect 7640 4550 7680 4590
rect 7680 4550 7690 4590
rect 7630 4540 7690 4550
rect 8150 4590 8210 4600
rect 8150 4550 8160 4590
rect 8160 4550 8200 4590
rect 8200 4550 8210 4590
rect 8150 4540 8210 4550
rect 8760 4540 8820 4600
rect 3800 4420 4220 4430
rect 3800 4380 3810 4420
rect 3810 4380 3850 4420
rect 3850 4380 3900 4420
rect 3900 4380 3940 4420
rect 3940 4380 3990 4420
rect 3990 4380 4030 4420
rect 4030 4380 4080 4420
rect 4080 4380 4120 4420
rect 4120 4380 4170 4420
rect 4170 4380 4210 4420
rect 4210 4380 4220 4420
rect 3800 4370 4220 4380
rect 1200 3960 1260 4020
rect 890 3370 950 3430
rect 1900 4010 1960 4020
rect 1900 3970 1910 4010
rect 1910 3970 1950 4010
rect 1950 3970 1960 4010
rect 1900 3960 1960 3970
rect 5230 4500 5290 4510
rect 5230 4460 5240 4500
rect 5240 4460 5280 4500
rect 5280 4460 5290 4500
rect 5230 4450 5290 4460
rect 6030 4500 6090 4510
rect 6030 4460 6040 4500
rect 6040 4460 6080 4500
rect 6080 4460 6090 4500
rect 6030 4450 6090 4460
rect 5630 4410 5690 4420
rect 5630 4370 5640 4410
rect 5640 4370 5680 4410
rect 5680 4370 5690 4410
rect 5630 4360 5690 4370
rect 6430 4410 6490 4420
rect 6430 4370 6440 4410
rect 6440 4370 6480 4410
rect 6480 4370 6490 4410
rect 6430 4360 6490 4370
rect 8030 4500 8090 4510
rect 8030 4460 8040 4500
rect 8040 4460 8080 4500
rect 8080 4460 8090 4500
rect 8030 4450 8090 4460
rect 8640 4450 8700 4510
rect 7230 4410 7290 4420
rect 7230 4370 7240 4410
rect 7240 4370 7280 4410
rect 7280 4370 7290 4410
rect 7230 4360 7290 4370
rect 4470 4220 4530 4230
rect 4470 4180 4480 4220
rect 4480 4180 4520 4220
rect 4520 4180 4530 4220
rect 4470 4170 4530 4180
rect 4670 4220 4730 4230
rect 4670 4180 4680 4220
rect 4680 4180 4720 4220
rect 4720 4180 4730 4220
rect 4670 4170 4730 4180
rect 5070 4220 5130 4230
rect 5070 4180 5080 4220
rect 5080 4180 5120 4220
rect 5120 4180 5130 4220
rect 5070 4170 5130 4180
rect 5470 4220 5530 4230
rect 5470 4180 5480 4220
rect 5480 4180 5520 4220
rect 5520 4180 5530 4220
rect 5470 4170 5530 4180
rect 5670 4220 5730 4230
rect 5670 4180 5680 4220
rect 5680 4180 5720 4220
rect 5720 4180 5730 4220
rect 5670 4170 5730 4180
rect 5830 4220 5890 4230
rect 5830 4180 5840 4220
rect 5840 4180 5880 4220
rect 5880 4180 5890 4220
rect 5830 4170 5890 4180
rect 6030 4220 6090 4230
rect 6030 4180 6040 4220
rect 6040 4180 6080 4220
rect 6080 4180 6090 4220
rect 6030 4170 6090 4180
rect 6430 4220 6490 4230
rect 6430 4180 6440 4220
rect 6440 4180 6480 4220
rect 6480 4180 6490 4220
rect 6430 4170 6490 4180
rect 6830 4220 6890 4230
rect 6830 4180 6840 4220
rect 6840 4180 6880 4220
rect 6880 4180 6890 4220
rect 6830 4170 6890 4180
rect 7030 4220 7090 4230
rect 7030 4180 7040 4220
rect 7040 4180 7080 4220
rect 7080 4180 7090 4220
rect 7030 4170 7090 4180
rect 7190 4220 7250 4230
rect 7190 4180 7200 4220
rect 7200 4180 7240 4220
rect 7240 4180 7250 4220
rect 7190 4170 7250 4180
rect 7390 4220 7450 4230
rect 7390 4180 7400 4220
rect 7400 4180 7440 4220
rect 7440 4180 7450 4220
rect 7390 4170 7450 4180
rect 7790 4220 7850 4230
rect 7790 4180 7800 4220
rect 7800 4180 7840 4220
rect 7840 4180 7850 4220
rect 7790 4170 7850 4180
rect 8190 4220 8250 4230
rect 8190 4180 8200 4220
rect 8200 4180 8240 4220
rect 8240 4180 8250 4220
rect 8190 4170 8250 4180
rect 8390 4220 8450 4230
rect 8390 4180 8400 4220
rect 8400 4180 8440 4220
rect 8440 4180 8450 4220
rect 8390 4170 8450 4180
rect 5270 3680 5330 3690
rect 5270 3640 5280 3680
rect 5280 3640 5320 3680
rect 5320 3640 5330 3680
rect 5270 3630 5330 3640
rect 5950 3630 6010 3690
rect 6910 3630 6970 3690
rect 7590 3680 7650 3690
rect 7590 3640 7600 3680
rect 7600 3640 7640 3680
rect 7640 3640 7650 3680
rect 7590 3630 7650 3640
rect 4870 3590 4930 3600
rect 4870 3550 4880 3590
rect 4880 3550 4920 3590
rect 4920 3550 4930 3590
rect 4870 3540 4930 3550
rect 5550 3540 5610 3600
rect 6130 3590 6190 3600
rect 6130 3550 6140 3590
rect 6140 3550 6180 3590
rect 6180 3550 6190 3590
rect 6130 3540 6190 3550
rect 6730 3590 6790 3600
rect 6730 3550 6740 3590
rect 6740 3550 6780 3590
rect 6780 3550 6790 3590
rect 6730 3540 6790 3550
rect 6430 3500 6490 3510
rect 6430 3460 6440 3500
rect 6440 3460 6480 3500
rect 6480 3460 6490 3500
rect 6430 3450 6490 3460
rect 7310 3540 7370 3600
rect 7990 3590 8050 3600
rect 7990 3550 8000 3590
rect 8000 3550 8040 3590
rect 8040 3550 8050 3590
rect 7990 3540 8050 3550
rect 7850 3450 7910 3510
rect 3800 3420 4220 3430
rect 3800 3380 3810 3420
rect 3810 3380 3850 3420
rect 3850 3380 3900 3420
rect 3900 3380 3940 3420
rect 3940 3380 3990 3420
rect 3990 3380 4030 3420
rect 4030 3380 4080 3420
rect 4080 3380 4120 3420
rect 4120 3380 4170 3420
rect 4170 3380 4210 3420
rect 4210 3380 4220 3420
rect 3800 3370 4220 3380
rect 4310 3360 4370 3420
rect 6070 3410 6130 3420
rect 6070 3370 6080 3410
rect 6080 3370 6120 3410
rect 6120 3370 6130 3410
rect 6070 3360 6130 3370
rect 6790 3410 6850 3420
rect 6790 3370 6800 3410
rect 6800 3370 6840 3410
rect 6840 3370 6850 3410
rect 6790 3360 6850 3370
rect 1730 3010 1790 3070
rect 1420 2420 1480 2480
rect 1900 3060 1960 3070
rect 1900 3020 1910 3060
rect 1910 3020 1950 3060
rect 1950 3020 1960 3060
rect 1900 3010 1960 3020
rect 3800 3060 4220 3070
rect 3800 3020 3810 3060
rect 3810 3020 3850 3060
rect 3850 3020 3900 3060
rect 3900 3020 3940 3060
rect 3940 3020 3990 3060
rect 3990 3020 4030 3060
rect 4030 3020 4080 3060
rect 4080 3020 4120 3060
rect 4120 3020 4170 3060
rect 4170 3020 4210 3060
rect 4210 3020 4220 3060
rect 3800 3010 4220 3020
rect 5550 3070 5610 3080
rect 5550 3030 5560 3070
rect 5560 3030 5600 3070
rect 5600 3030 5610 3070
rect 5550 3020 5610 3030
rect 7310 3070 7370 3080
rect 7310 3030 7320 3070
rect 7320 3030 7360 3070
rect 7360 3030 7370 3070
rect 7310 3020 7370 3030
rect 5150 2980 5210 2990
rect 5150 2940 5160 2980
rect 5160 2940 5200 2980
rect 5200 2940 5210 2980
rect 5150 2930 5210 2940
rect 5350 2980 5410 2990
rect 5350 2940 5360 2980
rect 5360 2940 5400 2980
rect 5400 2940 5410 2980
rect 5350 2930 5410 2940
rect 5750 2980 5810 2990
rect 5750 2940 5760 2980
rect 5760 2940 5800 2980
rect 5800 2940 5810 2980
rect 5750 2930 5810 2940
rect 6150 2980 6210 2990
rect 6150 2940 6160 2980
rect 6160 2940 6200 2980
rect 6200 2940 6210 2980
rect 6150 2930 6210 2940
rect 6350 2980 6410 2990
rect 6350 2940 6360 2980
rect 6360 2940 6400 2980
rect 6400 2940 6410 2980
rect 6350 2930 6410 2940
rect 6510 2980 6570 2990
rect 6510 2940 6520 2980
rect 6520 2940 6560 2980
rect 6560 2940 6570 2980
rect 6510 2930 6570 2940
rect 6710 2980 6770 2990
rect 6710 2940 6720 2980
rect 6720 2940 6760 2980
rect 6760 2940 6770 2980
rect 6710 2930 6770 2940
rect 7110 2980 7170 2990
rect 7110 2940 7120 2980
rect 7120 2940 7160 2980
rect 7160 2940 7170 2980
rect 7110 2930 7170 2940
rect 7510 2980 7570 2990
rect 7510 2940 7520 2980
rect 7520 2940 7560 2980
rect 7560 2940 7570 2980
rect 7510 2930 7570 2940
rect 7710 2980 7770 2990
rect 7710 2940 7720 2980
rect 7720 2940 7760 2980
rect 7760 2940 7770 2980
rect 7710 2930 7770 2940
rect 9160 4220 9220 4230
rect 9160 4180 9170 4220
rect 9170 4180 9210 4220
rect 9210 4180 9220 4220
rect 9160 4170 9220 4180
rect 8870 3410 8930 3420
rect 8870 3370 8880 3410
rect 8880 3370 8920 3410
rect 8920 3370 8930 3410
rect 8870 3360 8930 3370
rect 8640 3020 8700 3080
rect 7310 2860 7370 2870
rect 7310 2820 7320 2860
rect 7320 2820 7360 2860
rect 7360 2820 7370 2860
rect 7310 2810 7370 2820
rect 7850 2810 7910 2870
rect 1900 2470 1960 2480
rect 1900 2430 1910 2470
rect 1910 2430 1950 2470
rect 1950 2430 1960 2470
rect 1900 2420 1960 2430
rect 4670 1920 4730 1930
rect 4670 1880 4680 1920
rect 4680 1880 4720 1920
rect 4720 1880 4730 1920
rect 4670 1870 4730 1880
rect 6430 1920 6490 1930
rect 6430 1880 6440 1920
rect 6440 1880 6480 1920
rect 6480 1880 6490 1920
rect 6430 1870 6490 1880
rect 8190 1920 8250 1930
rect 8190 1880 8200 1920
rect 8200 1880 8240 1920
rect 8240 1880 8250 1920
rect 8190 1870 8250 1880
rect 7450 1800 7510 1810
rect 7450 1760 7460 1800
rect 7460 1760 7500 1800
rect 7500 1760 7510 1800
rect 7450 1750 7510 1760
rect 9000 1750 9060 1810
rect 30 90 90 100
rect 30 50 40 90
rect 40 50 80 90
rect 80 50 90 90
rect 30 40 90 50
rect 210 90 270 100
rect 210 50 220 90
rect 220 50 260 90
rect 260 50 270 90
rect 210 40 270 50
rect 390 90 450 100
rect 390 50 400 90
rect 400 50 440 90
rect 440 50 450 90
rect 390 40 450 50
rect 570 90 630 100
rect 570 50 580 90
rect 580 50 620 90
rect 620 50 630 90
rect 570 40 630 50
rect 750 90 810 100
rect 750 50 760 90
rect 760 50 800 90
rect 800 50 810 90
rect 750 40 810 50
rect 930 90 990 100
rect 930 50 940 90
rect 940 50 980 90
rect 980 50 990 90
rect 930 40 990 50
rect 1110 90 1170 100
rect 1110 50 1120 90
rect 1120 50 1160 90
rect 1160 50 1170 90
rect 1110 40 1170 50
rect 1290 90 1350 100
rect 1290 50 1300 90
rect 1300 50 1340 90
rect 1340 50 1350 90
rect 1290 40 1350 50
rect 1470 90 1530 100
rect 1470 50 1480 90
rect 1480 50 1520 90
rect 1520 50 1530 90
rect 1470 40 1530 50
rect 1650 90 1710 100
rect 1650 50 1660 90
rect 1660 50 1700 90
rect 1700 50 1710 90
rect 1650 40 1710 50
rect 1830 90 1890 100
rect 1830 50 1840 90
rect 1840 50 1880 90
rect 1880 50 1890 90
rect 1830 40 1890 50
rect 2010 90 2070 100
rect 2010 50 2020 90
rect 2020 50 2060 90
rect 2060 50 2070 90
rect 2010 40 2070 50
rect 2190 90 2250 100
rect 2190 50 2200 90
rect 2200 50 2240 90
rect 2240 50 2250 90
rect 2190 40 2250 50
rect 2370 90 2430 100
rect 2370 50 2380 90
rect 2380 50 2420 90
rect 2420 50 2430 90
rect 2370 40 2430 50
rect 2550 90 2610 100
rect 2550 50 2560 90
rect 2560 50 2600 90
rect 2600 50 2610 90
rect 2550 40 2610 50
rect 2730 90 2790 100
rect 2730 50 2740 90
rect 2740 50 2780 90
rect 2780 50 2790 90
rect 2730 40 2790 50
rect 2910 90 2970 100
rect 2910 50 2920 90
rect 2920 50 2960 90
rect 2960 50 2970 90
rect 2910 40 2970 50
rect 3090 90 3150 100
rect 3090 50 3100 90
rect 3100 50 3140 90
rect 3140 50 3150 90
rect 3090 40 3150 50
rect 3270 90 3330 100
rect 3270 50 3280 90
rect 3280 50 3320 90
rect 3320 50 3330 90
rect 3270 40 3330 50
rect 3450 90 3510 100
rect 3450 50 3460 90
rect 3460 50 3500 90
rect 3500 50 3510 90
rect 3450 40 3510 50
rect 3630 90 3690 100
rect 3630 50 3640 90
rect 3640 50 3680 90
rect 3680 50 3690 90
rect 3630 40 3690 50
rect 3810 90 3870 100
rect 3810 50 3820 90
rect 3820 50 3860 90
rect 3860 50 3870 90
rect 3810 40 3870 50
rect 3990 90 4050 100
rect 3990 50 4000 90
rect 4000 50 4040 90
rect 4040 50 4050 90
rect 3990 40 4050 50
rect 4170 90 4230 100
rect 4170 50 4180 90
rect 4180 50 4220 90
rect 4220 50 4230 90
rect 4170 40 4230 50
rect 4350 90 4410 100
rect 4350 50 4360 90
rect 4360 50 4400 90
rect 4400 50 4410 90
rect 4350 40 4410 50
rect 4530 90 4590 100
rect 4530 50 4540 90
rect 4540 50 4580 90
rect 4580 50 4590 90
rect 4530 40 4590 50
rect 4710 90 4770 100
rect 4710 50 4720 90
rect 4720 50 4760 90
rect 4760 50 4770 90
rect 4710 40 4770 50
rect 4890 90 4950 100
rect 4890 50 4900 90
rect 4900 50 4940 90
rect 4940 50 4950 90
rect 4890 40 4950 50
rect 5070 90 5130 100
rect 5070 50 5080 90
rect 5080 50 5120 90
rect 5120 50 5130 90
rect 5070 40 5130 50
rect 5250 90 5310 100
rect 5250 50 5260 90
rect 5260 50 5300 90
rect 5300 50 5310 90
rect 5250 40 5310 50
rect 5430 90 5490 100
rect 5430 50 5440 90
rect 5440 50 5480 90
rect 5480 50 5490 90
rect 5430 40 5490 50
rect 5610 90 5670 100
rect 5610 50 5620 90
rect 5620 50 5660 90
rect 5660 50 5670 90
rect 5610 40 5670 50
rect 5790 90 5850 100
rect 5790 50 5800 90
rect 5800 50 5840 90
rect 5840 50 5850 90
rect 5790 40 5850 50
rect 5970 90 6030 100
rect 5970 50 5980 90
rect 5980 50 6020 90
rect 6020 50 6030 90
rect 5970 40 6030 50
rect 6150 90 6210 100
rect 6150 50 6160 90
rect 6160 50 6200 90
rect 6200 50 6210 90
rect 6150 40 6210 50
rect 6330 90 6390 100
rect 6330 50 6340 90
rect 6340 50 6380 90
rect 6380 50 6390 90
rect 6330 40 6390 50
rect 6510 90 6570 100
rect 6510 50 6520 90
rect 6520 50 6560 90
rect 6560 50 6570 90
rect 6510 40 6570 50
rect 6690 90 6750 100
rect 6690 50 6700 90
rect 6700 50 6740 90
rect 6740 50 6750 90
rect 6690 40 6750 50
rect 6870 90 6930 100
rect 6870 50 6880 90
rect 6880 50 6920 90
rect 6920 50 6930 90
rect 6870 40 6930 50
rect 7050 90 7110 100
rect 7050 50 7060 90
rect 7060 50 7100 90
rect 7100 50 7110 90
rect 7050 40 7110 50
rect 7230 90 7290 100
rect 7230 50 7240 90
rect 7240 50 7280 90
rect 7280 50 7290 90
rect 7230 40 7290 50
rect 7410 90 7470 100
rect 7410 50 7420 90
rect 7420 50 7460 90
rect 7460 50 7470 90
rect 7410 40 7470 50
rect 7590 90 7650 100
rect 7590 50 7600 90
rect 7600 50 7640 90
rect 7640 50 7650 90
rect 7590 40 7650 50
rect 7770 90 7830 100
rect 7770 50 7780 90
rect 7780 50 7820 90
rect 7820 50 7830 90
rect 7770 40 7830 50
rect 7950 90 8010 100
rect 7950 50 7960 90
rect 7960 50 8000 90
rect 8000 50 8010 90
rect 7950 40 8010 50
rect 8130 90 8190 100
rect 8130 50 8140 90
rect 8140 50 8180 90
rect 8180 50 8190 90
rect 8130 40 8190 50
rect 8310 90 8370 100
rect 8310 50 8320 90
rect 8320 50 8360 90
rect 8360 50 8370 90
rect 8310 40 8370 50
rect 8490 90 8550 100
rect 8490 50 8500 90
rect 8500 50 8540 90
rect 8540 50 8550 90
rect 8490 40 8550 50
rect 8670 90 8730 100
rect 8670 50 8680 90
rect 8680 50 8720 90
rect 8720 50 8730 90
rect 8670 40 8730 50
rect 8850 90 8910 100
rect 8850 50 8860 90
rect 8860 50 8900 90
rect 8900 50 8910 90
rect 8850 40 8910 50
rect 9030 90 9090 100
rect 9030 50 9040 90
rect 9040 50 9080 90
rect 9080 50 9090 90
rect 9030 40 9090 50
rect 9210 90 9270 100
rect 9210 50 9220 90
rect 9220 50 9260 90
rect 9260 50 9270 90
rect 9210 40 9270 50
rect 9390 90 9450 100
rect 9390 50 9400 90
rect 9400 50 9440 90
rect 9440 50 9450 90
rect 9390 40 9450 50
<< metal2 >>
rect -1940 6960 -1860 6970
rect -1940 6900 -1930 6960
rect -1870 6900 -1860 6960
rect -1940 6890 -1860 6900
rect 11810 6960 11890 6970
rect 11810 6900 11820 6960
rect 11880 6900 11890 6960
rect 11810 6890 11890 6900
rect -1940 5540 -1860 5550
rect -1940 5530 -1930 5540
rect -3290 5490 -1930 5530
rect -1940 5480 -1930 5490
rect -1870 5530 -1860 5540
rect 4620 5540 4700 5550
rect 4620 5530 4630 5540
rect -1870 5490 4630 5530
rect -1870 5480 -1860 5490
rect -1940 5470 -1860 5480
rect 4620 5480 4630 5490
rect 4690 5530 4700 5540
rect 5020 5540 5100 5550
rect 5020 5530 5030 5540
rect 4690 5490 5030 5530
rect 4690 5480 4700 5490
rect 4620 5470 4700 5480
rect 5020 5480 5030 5490
rect 5090 5530 5100 5540
rect 5420 5540 5500 5550
rect 5420 5530 5430 5540
rect 5090 5490 5430 5530
rect 5090 5480 5100 5490
rect 5020 5470 5100 5480
rect 5420 5480 5430 5490
rect 5490 5530 5500 5540
rect 5820 5540 5900 5550
rect 5820 5530 5830 5540
rect 5490 5490 5830 5530
rect 5490 5480 5500 5490
rect 5420 5470 5500 5480
rect 5820 5480 5830 5490
rect 5890 5530 5900 5540
rect 6220 5540 6300 5550
rect 6220 5530 6230 5540
rect 5890 5490 6230 5530
rect 5890 5480 5900 5490
rect 5820 5470 5900 5480
rect 6220 5480 6230 5490
rect 6290 5530 6300 5540
rect 6620 5540 6700 5550
rect 6620 5530 6630 5540
rect 6290 5490 6630 5530
rect 6290 5480 6300 5490
rect 6220 5470 6300 5480
rect 6620 5480 6630 5490
rect 6690 5530 6700 5540
rect 7020 5540 7100 5550
rect 7020 5530 7030 5540
rect 6690 5490 7030 5530
rect 6690 5480 6700 5490
rect 6620 5470 6700 5480
rect 7020 5480 7030 5490
rect 7090 5530 7100 5540
rect 7420 5540 7500 5550
rect 7420 5530 7430 5540
rect 7090 5490 7430 5530
rect 7090 5480 7100 5490
rect 7020 5470 7100 5480
rect 7420 5480 7430 5490
rect 7490 5530 7500 5540
rect 7820 5540 7900 5550
rect 7820 5530 7830 5540
rect 7490 5490 7830 5530
rect 7490 5480 7500 5490
rect 7420 5470 7500 5480
rect 7820 5480 7830 5490
rect 7890 5530 7900 5540
rect 8220 5540 8300 5550
rect 8220 5530 8230 5540
rect 7890 5490 8230 5530
rect 7890 5480 7900 5490
rect 7820 5470 7900 5480
rect 8220 5480 8230 5490
rect 8290 5530 8300 5540
rect 11810 5540 11890 5550
rect 11810 5530 11820 5540
rect 8290 5490 11820 5530
rect 8290 5480 8300 5490
rect 8220 5470 8300 5480
rect 11810 5480 11820 5490
rect 11880 5530 11890 5540
rect 11880 5490 13010 5530
rect 11880 5480 11890 5490
rect 11810 5470 11890 5480
rect 1190 5020 1970 5030
rect 1190 4960 1200 5020
rect 1260 4960 1900 5020
rect 1960 4960 1970 5020
rect 1190 4950 1970 4960
rect 4300 4600 4380 4610
rect 4300 4540 4310 4600
rect 4370 4590 4380 4600
rect 4820 4600 4900 4610
rect 4820 4590 4830 4600
rect 4370 4550 4830 4590
rect 4370 4540 4380 4550
rect 4300 4530 4380 4540
rect 4820 4540 4830 4550
rect 4890 4590 4900 4600
rect 6820 4600 6900 4610
rect 6820 4590 6830 4600
rect 4890 4550 6830 4590
rect 4890 4540 4900 4550
rect 4820 4530 4900 4540
rect 6820 4540 6830 4550
rect 6890 4590 6900 4600
rect 7620 4600 7700 4610
rect 7620 4590 7630 4600
rect 6890 4550 7630 4590
rect 6890 4540 6900 4550
rect 6820 4530 6900 4540
rect 7620 4540 7630 4550
rect 7690 4540 7700 4600
rect 7620 4530 7700 4540
rect 8140 4600 8220 4610
rect 8140 4540 8150 4600
rect 8210 4590 8220 4600
rect 8750 4600 8830 4610
rect 8750 4590 8760 4600
rect 8210 4550 8760 4590
rect 8210 4540 8220 4550
rect 8140 4530 8220 4540
rect 8750 4540 8760 4550
rect 8820 4540 8830 4600
rect 8750 4530 8830 4540
rect 5220 4510 5300 4520
rect 5220 4450 5230 4510
rect 5290 4500 5300 4510
rect 6020 4510 6100 4520
rect 6020 4500 6030 4510
rect 5290 4460 6030 4500
rect 5290 4450 5300 4460
rect 5220 4440 5300 4450
rect 6020 4450 6030 4460
rect 6090 4500 6100 4510
rect 8020 4510 8100 4520
rect 8020 4500 8030 4510
rect 6090 4460 8030 4500
rect 6090 4450 6100 4460
rect 6020 4440 6100 4450
rect 8020 4450 8030 4460
rect 8090 4500 8100 4510
rect 8630 4510 8710 4520
rect 8630 4500 8640 4510
rect 8090 4460 8640 4500
rect 8090 4450 8100 4460
rect 8020 4440 8100 4450
rect 8630 4450 8640 4460
rect 8700 4450 8710 4510
rect 8630 4440 8710 4450
rect 3790 4430 4230 4440
rect 3790 4370 3800 4430
rect 4220 4410 4230 4430
rect 5620 4420 5700 4430
rect 5620 4410 5630 4420
rect 4220 4370 5630 4410
rect 3790 4360 4230 4370
rect 5620 4360 5630 4370
rect 5690 4410 5700 4420
rect 6420 4420 6500 4430
rect 6420 4410 6430 4420
rect 5690 4370 6430 4410
rect 5690 4360 5700 4370
rect 5620 4350 5700 4360
rect 6420 4360 6430 4370
rect 6490 4410 6500 4420
rect 7220 4420 7300 4430
rect 7220 4410 7230 4420
rect 6490 4370 7230 4410
rect 6490 4360 6500 4370
rect 6420 4350 6500 4360
rect 7220 4360 7230 4370
rect 7290 4360 7300 4420
rect 7220 4350 7300 4360
rect 4460 4230 4540 4240
rect 4460 4170 4470 4230
rect 4530 4220 4540 4230
rect 4660 4230 4740 4240
rect 4660 4220 4670 4230
rect 4530 4180 4670 4220
rect 4530 4170 4540 4180
rect 4460 4160 4540 4170
rect 4660 4170 4670 4180
rect 4730 4220 4740 4230
rect 5060 4230 5140 4240
rect 5060 4220 5070 4230
rect 4730 4180 5070 4220
rect 4730 4170 4740 4180
rect 4660 4160 4740 4170
rect 5060 4170 5070 4180
rect 5130 4220 5140 4230
rect 5460 4230 5540 4240
rect 5460 4220 5470 4230
rect 5130 4180 5470 4220
rect 5130 4170 5140 4180
rect 5060 4160 5140 4170
rect 5460 4170 5470 4180
rect 5530 4220 5540 4230
rect 5660 4230 5740 4240
rect 5660 4220 5670 4230
rect 5530 4180 5670 4220
rect 5530 4170 5540 4180
rect 5460 4160 5540 4170
rect 5660 4170 5670 4180
rect 5730 4220 5740 4230
rect 5820 4230 5900 4240
rect 5820 4220 5830 4230
rect 5730 4180 5830 4220
rect 5730 4170 5740 4180
rect 5660 4160 5740 4170
rect 5820 4170 5830 4180
rect 5890 4220 5900 4230
rect 6020 4230 6100 4240
rect 6020 4220 6030 4230
rect 5890 4180 6030 4220
rect 5890 4170 5900 4180
rect 5820 4160 5900 4170
rect 6020 4170 6030 4180
rect 6090 4220 6100 4230
rect 6420 4230 6500 4240
rect 6420 4220 6430 4230
rect 6090 4180 6430 4220
rect 6090 4170 6100 4180
rect 6020 4160 6100 4170
rect 6420 4170 6430 4180
rect 6490 4220 6500 4230
rect 6820 4230 6900 4240
rect 6820 4220 6830 4230
rect 6490 4180 6830 4220
rect 6490 4170 6500 4180
rect 6420 4160 6500 4170
rect 6820 4170 6830 4180
rect 6890 4220 6900 4230
rect 7020 4230 7100 4240
rect 7020 4220 7030 4230
rect 6890 4180 7030 4220
rect 6890 4170 6900 4180
rect 6820 4160 6900 4170
rect 7020 4170 7030 4180
rect 7090 4220 7100 4230
rect 7180 4230 7260 4240
rect 7180 4220 7190 4230
rect 7090 4180 7190 4220
rect 7090 4170 7100 4180
rect 7020 4160 7100 4170
rect 7180 4170 7190 4180
rect 7250 4220 7260 4230
rect 7380 4230 7460 4240
rect 7380 4220 7390 4230
rect 7250 4180 7390 4220
rect 7250 4170 7260 4180
rect 7180 4160 7260 4170
rect 7380 4170 7390 4180
rect 7450 4220 7460 4230
rect 7780 4230 7860 4240
rect 7780 4220 7790 4230
rect 7450 4180 7790 4220
rect 7450 4170 7460 4180
rect 7380 4160 7460 4170
rect 7780 4170 7790 4180
rect 7850 4220 7860 4230
rect 8180 4230 8260 4240
rect 8180 4220 8190 4230
rect 7850 4180 8190 4220
rect 7850 4170 7860 4180
rect 7780 4160 7860 4170
rect 8180 4170 8190 4180
rect 8250 4220 8260 4230
rect 8380 4230 8460 4240
rect 8380 4220 8390 4230
rect 8250 4180 8390 4220
rect 8250 4170 8260 4180
rect 8180 4160 8260 4170
rect 8380 4170 8390 4180
rect 8450 4220 8460 4230
rect 9150 4230 9230 4240
rect 9150 4220 9160 4230
rect 8450 4180 9160 4220
rect 8450 4170 8460 4180
rect 8380 4160 8460 4170
rect 9150 4170 9160 4180
rect 9220 4220 9230 4230
rect 11810 4230 11890 4240
rect 11810 4220 11820 4230
rect 9220 4180 11820 4220
rect 9220 4170 9230 4180
rect 9150 4160 9230 4170
rect 11810 4170 11820 4180
rect 11880 4220 11890 4230
rect 11880 4180 13050 4220
rect 11880 4170 11890 4180
rect 11810 4160 11890 4170
rect 1190 4020 1970 4030
rect 1190 3960 1200 4020
rect 1260 3960 1900 4020
rect 1960 3960 1970 4020
rect 1190 3950 1970 3960
rect 5260 3690 5340 3700
rect 5260 3630 5270 3690
rect 5330 3680 5340 3690
rect 5940 3690 6020 3700
rect 5940 3680 5950 3690
rect 5330 3640 5950 3680
rect 5330 3630 5340 3640
rect 5260 3620 5340 3630
rect 5940 3630 5950 3640
rect 6010 3680 6020 3690
rect 6900 3690 6980 3700
rect 6900 3680 6910 3690
rect 6010 3640 6910 3680
rect 6010 3630 6020 3640
rect 5940 3620 6020 3630
rect 6900 3630 6910 3640
rect 6970 3680 6980 3690
rect 7580 3690 7660 3700
rect 7580 3680 7590 3690
rect 6970 3640 7590 3680
rect 6970 3630 6980 3640
rect 6900 3620 6980 3630
rect 7580 3630 7590 3640
rect 7650 3630 7660 3690
rect 7580 3620 7660 3630
rect 4860 3600 4940 3610
rect 4860 3540 4870 3600
rect 4930 3590 4940 3600
rect 5540 3600 5620 3610
rect 5540 3590 5550 3600
rect 4930 3550 5550 3590
rect 4930 3540 4940 3550
rect 4860 3530 4940 3540
rect 5540 3540 5550 3550
rect 5610 3590 5620 3600
rect 6120 3600 6200 3610
rect 6120 3590 6130 3600
rect 5610 3550 6130 3590
rect 5610 3540 5620 3550
rect 5540 3530 5620 3540
rect 6120 3540 6130 3550
rect 6190 3590 6200 3600
rect 6720 3600 6800 3610
rect 6720 3590 6730 3600
rect 6190 3550 6730 3590
rect 6190 3540 6200 3550
rect 6120 3530 6200 3540
rect 6720 3540 6730 3550
rect 6790 3590 6800 3600
rect 7300 3600 7380 3610
rect 7300 3590 7310 3600
rect 6790 3550 7310 3590
rect 6790 3540 6800 3550
rect 6720 3530 6800 3540
rect 7300 3540 7310 3550
rect 7370 3590 7380 3600
rect 7980 3600 8060 3610
rect 7980 3590 7990 3600
rect 7370 3550 7990 3590
rect 7370 3540 7380 3550
rect 7300 3530 7380 3540
rect 7980 3540 7990 3550
rect 8050 3540 8060 3600
rect 7980 3530 8060 3540
rect 6420 3510 6500 3520
rect 6420 3450 6430 3510
rect 6490 3500 6500 3510
rect 7840 3510 7920 3520
rect 7840 3500 7850 3510
rect 6490 3460 7850 3500
rect 6490 3450 6500 3460
rect 6420 3440 6500 3450
rect 7840 3450 7850 3460
rect 7910 3450 7920 3510
rect 7840 3440 7920 3450
rect 880 3430 4230 3440
rect 880 3370 890 3430
rect 950 3370 3800 3430
rect 4220 3410 4230 3430
rect 4300 3420 4380 3430
rect 4300 3410 4310 3420
rect 4220 3370 4310 3410
rect 880 3360 4230 3370
rect 4300 3360 4310 3370
rect 4370 3410 4380 3420
rect 6060 3420 6140 3430
rect 6060 3410 6070 3420
rect 4370 3370 6070 3410
rect 4370 3360 4380 3370
rect 4300 3350 4380 3360
rect 6060 3360 6070 3370
rect 6130 3410 6140 3420
rect 6780 3420 6860 3430
rect 6780 3410 6790 3420
rect 6130 3370 6790 3410
rect 6130 3360 6140 3370
rect 6060 3350 6140 3360
rect 6780 3360 6790 3370
rect 6850 3410 6860 3420
rect 8860 3420 8940 3430
rect 8860 3410 8870 3420
rect 6850 3370 8870 3410
rect 6850 3360 6860 3370
rect 6780 3350 6860 3360
rect 8860 3360 8870 3370
rect 8930 3360 8940 3420
rect 8860 3350 8940 3360
rect 5540 3080 5620 3090
rect 1720 3070 1970 3080
rect 1720 3010 1730 3070
rect 1790 3010 1900 3070
rect 1960 3010 1970 3070
rect 1720 3000 1970 3010
rect 3790 3070 4230 3080
rect 5540 3070 5550 3080
rect 3790 3010 3800 3070
rect 4220 3030 5550 3070
rect 4220 3010 4230 3030
rect 5540 3020 5550 3030
rect 5610 3070 5620 3080
rect 7300 3080 7380 3090
rect 7300 3070 7310 3080
rect 5610 3030 7310 3070
rect 5610 3020 5620 3030
rect 5540 3010 5620 3020
rect 7300 3020 7310 3030
rect 7370 3070 7380 3080
rect 8630 3080 8710 3090
rect 8630 3070 8640 3080
rect 7370 3030 8640 3070
rect 7370 3020 7380 3030
rect 7300 3010 7380 3020
rect 8630 3020 8640 3030
rect 8700 3020 8710 3080
rect 8630 3010 8710 3020
rect 3790 3000 4230 3010
rect 5140 2990 5220 3000
rect 5140 2930 5150 2990
rect 5210 2980 5220 2990
rect 5340 2990 5420 3000
rect 5340 2980 5350 2990
rect 5210 2940 5350 2980
rect 5210 2930 5220 2940
rect 5140 2920 5220 2930
rect 5340 2930 5350 2940
rect 5410 2980 5420 2990
rect 5740 2990 5820 3000
rect 5740 2980 5750 2990
rect 5410 2940 5750 2980
rect 5410 2930 5420 2940
rect 5340 2920 5420 2930
rect 5740 2930 5750 2940
rect 5810 2980 5820 2990
rect 6140 2990 6220 3000
rect 6140 2980 6150 2990
rect 5810 2940 6150 2980
rect 5810 2930 5820 2940
rect 5740 2920 5820 2930
rect 6140 2930 6150 2940
rect 6210 2980 6220 2990
rect 6340 2990 6420 3000
rect 6340 2980 6350 2990
rect 6210 2940 6350 2980
rect 6210 2930 6220 2940
rect 6140 2920 6220 2930
rect 6340 2930 6350 2940
rect 6410 2980 6420 2990
rect 6500 2990 6580 3000
rect 6500 2980 6510 2990
rect 6410 2940 6510 2980
rect 6410 2930 6420 2940
rect 6340 2920 6420 2930
rect 6500 2930 6510 2940
rect 6570 2980 6580 2990
rect 6700 2990 6780 3000
rect 6700 2980 6710 2990
rect 6570 2940 6710 2980
rect 6570 2930 6580 2940
rect 6500 2920 6580 2930
rect 6700 2930 6710 2940
rect 6770 2980 6780 2990
rect 7100 2990 7180 3000
rect 7100 2980 7110 2990
rect 6770 2940 7110 2980
rect 6770 2930 6780 2940
rect 6700 2920 6780 2930
rect 7100 2930 7110 2940
rect 7170 2980 7180 2990
rect 7500 2990 7580 3000
rect 7500 2980 7510 2990
rect 7170 2940 7510 2980
rect 7170 2930 7180 2940
rect 7100 2920 7180 2930
rect 7500 2930 7510 2940
rect 7570 2980 7580 2990
rect 7700 2990 7780 3000
rect 7700 2980 7710 2990
rect 7570 2940 7710 2980
rect 7570 2930 7580 2940
rect 7500 2920 7580 2930
rect 7700 2930 7710 2940
rect 7770 2930 7780 2990
rect 7700 2920 7780 2930
rect 7300 2870 7380 2880
rect 7300 2810 7310 2870
rect 7370 2860 7380 2870
rect 7840 2870 7920 2880
rect 7840 2860 7850 2870
rect 7370 2820 7850 2860
rect 7370 2810 7380 2820
rect 7300 2800 7380 2810
rect 7840 2810 7850 2820
rect 7910 2810 7920 2870
rect 7840 2800 7920 2810
rect 1410 2480 1970 2490
rect 1410 2420 1420 2480
rect 1480 2420 1900 2480
rect 1960 2420 1970 2480
rect 1410 2410 1970 2420
rect 4660 1930 4740 1940
rect 4660 1870 4670 1930
rect 4730 1920 4740 1930
rect 6420 1930 6500 1940
rect 6420 1920 6430 1930
rect 4730 1880 6430 1920
rect 4730 1870 4740 1880
rect 4660 1860 4740 1870
rect 6420 1870 6430 1880
rect 6490 1920 6500 1930
rect 8180 1930 8260 1940
rect 8180 1920 8190 1930
rect 6490 1880 8190 1920
rect 6490 1870 6500 1880
rect 6420 1860 6500 1870
rect 8180 1870 8190 1880
rect 8250 1920 8260 1930
rect 9920 1930 10000 1940
rect 9920 1920 9930 1930
rect 8250 1880 9930 1920
rect 8250 1870 8260 1880
rect 8180 1860 8260 1870
rect 9920 1870 9930 1880
rect 9990 1920 10000 1930
rect 9990 1880 10770 1920
rect 9990 1870 10000 1880
rect 9920 1860 10000 1870
rect 7440 1810 7520 1820
rect 7440 1750 7450 1810
rect 7510 1800 7520 1810
rect 8990 1810 9070 1820
rect 8990 1800 9000 1810
rect 7510 1760 9000 1800
rect 7510 1750 7520 1760
rect 7440 1740 7520 1750
rect 8990 1750 9000 1760
rect 9060 1750 9070 1810
rect 8990 1740 9070 1750
rect 9920 1630 10000 1640
rect 9920 1620 9930 1630
rect 7600 1580 9930 1620
rect 9920 1570 9930 1580
rect 9990 1620 10000 1630
rect 9990 1580 10770 1620
rect 9990 1570 10000 1580
rect 9920 1560 10000 1570
rect -940 100 11060 110
rect -940 40 -470 100
rect -410 40 30 100
rect 90 40 210 100
rect 270 40 390 100
rect 450 40 570 100
rect 630 40 750 100
rect 810 40 930 100
rect 990 40 1110 100
rect 1170 40 1290 100
rect 1350 40 1470 100
rect 1530 40 1650 100
rect 1710 40 1830 100
rect 1890 40 2010 100
rect 2070 40 2190 100
rect 2250 40 2370 100
rect 2430 40 2550 100
rect 2610 40 2730 100
rect 2790 40 2910 100
rect 2970 40 3090 100
rect 3150 40 3270 100
rect 3330 40 3450 100
rect 3510 40 3630 100
rect 3690 40 3810 100
rect 3870 40 3990 100
rect 4050 40 4170 100
rect 4230 40 4350 100
rect 4410 40 4530 100
rect 4590 40 4710 100
rect 4770 40 4890 100
rect 4950 40 5070 100
rect 5130 40 5250 100
rect 5310 40 5430 100
rect 5490 40 5610 100
rect 5670 40 5790 100
rect 5850 40 5970 100
rect 6030 40 6150 100
rect 6210 40 6330 100
rect 6390 40 6510 100
rect 6570 40 6690 100
rect 6750 40 6870 100
rect 6930 40 7050 100
rect 7110 40 7230 100
rect 7290 40 7410 100
rect 7470 40 7590 100
rect 7650 40 7770 100
rect 7830 40 7950 100
rect 8010 40 8130 100
rect 8190 40 8310 100
rect 8370 40 8490 100
rect 8550 40 8670 100
rect 8730 40 8850 100
rect 8910 40 9030 100
rect 9090 40 9210 100
rect 9270 40 9390 100
rect 9450 40 9930 100
rect 9990 40 11060 100
rect -940 30 11060 40
rect -1940 -1240 -1860 -1230
rect -1940 -1300 -1930 -1240
rect -1870 -1300 -1860 -1240
rect -1940 -1310 -1860 -1300
<< via2 >>
rect -1930 6900 -1870 6960
rect 11820 6900 11880 6960
rect -1930 5480 -1870 5540
rect 11820 5480 11880 5540
rect 11820 4170 11880 4230
rect 9930 1870 9990 1930
rect 9930 1570 9990 1630
rect -470 40 -410 100
rect 9930 40 9990 100
rect -1930 -1300 -1870 -1240
<< metal3 >>
rect -1940 6980 -1860 7500
rect 11810 6980 11890 7520
rect -1950 6970 -1850 6980
rect -1950 6890 -1940 6970
rect -1860 6890 -1850 6970
rect -1950 6880 -1850 6890
rect 11800 6970 11900 6980
rect 11800 6890 11810 6970
rect 11890 6890 11900 6970
rect 11800 6880 11900 6890
rect -1940 5540 -1860 6880
rect -480 6080 -400 6370
rect 9920 6080 10000 6370
rect -490 6070 -390 6080
rect -490 5990 -480 6070
rect -400 5990 -390 6070
rect -490 5980 -390 5990
rect 9910 6070 10010 6080
rect 9910 5990 9920 6070
rect 10000 5990 10010 6070
rect 9910 5980 10010 5990
rect -1940 5480 -1930 5540
rect -1870 5480 -1860 5540
rect -1940 -1220 -1860 5480
rect -480 100 -400 5980
rect -480 40 -470 100
rect -410 40 -400 100
rect -480 -220 -400 40
rect 9920 1930 10000 5980
rect 9920 1870 9930 1930
rect 9990 1870 10000 1930
rect 9920 1630 10000 1870
rect 9920 1570 9930 1630
rect 9990 1570 10000 1630
rect 9920 100 10000 1570
rect 9920 40 9930 100
rect 9990 40 10000 100
rect 9920 -220 10000 40
rect 11810 5540 11890 6880
rect 11810 5480 11820 5540
rect 11880 5480 11890 5540
rect 11810 4230 11890 5480
rect 11810 4170 11820 4230
rect 11880 4170 11890 4230
rect -490 -230 -390 -220
rect -490 -310 -480 -230
rect -400 -310 -390 -230
rect -490 -320 -390 -310
rect 9910 -230 10010 -220
rect 9910 -310 9920 -230
rect 10000 -310 10010 -230
rect 9910 -320 10010 -310
rect -480 -900 -400 -320
rect 9920 -810 10000 -320
rect 11810 -1220 11890 4170
rect -1950 -1230 -1850 -1220
rect -1950 -1310 -1940 -1230
rect -1860 -1310 -1850 -1230
rect -1950 -1320 -1850 -1310
rect 11800 -1230 11900 -1220
rect 11800 -1310 11810 -1230
rect 11890 -1310 11900 -1230
rect 11800 -1320 11900 -1310
rect -1940 -1820 -1860 -1320
rect 11810 -1800 11890 -1320
<< via3 >>
rect -1940 6960 -1860 6970
rect -1940 6900 -1930 6960
rect -1930 6900 -1870 6960
rect -1870 6900 -1860 6960
rect -1940 6890 -1860 6900
rect 11810 6960 11890 6970
rect 11810 6900 11820 6960
rect 11820 6900 11880 6960
rect 11880 6900 11890 6960
rect 11810 6890 11890 6900
rect -480 5990 -400 6070
rect 9920 5990 10000 6070
rect -480 -310 -400 -230
rect 9920 -310 10000 -230
rect -1940 -1240 -1860 -1230
rect -1940 -1300 -1930 -1240
rect -1930 -1300 -1870 -1240
rect -1870 -1300 -1860 -1240
rect -1940 -1310 -1860 -1300
rect 11810 -1310 11890 -1230
<< metal4 >>
rect -1950 6970 -1850 6980
rect 11800 6970 11900 6980
rect -2830 6890 -1940 6970
rect -1860 6890 11810 6970
rect 11890 6890 12840 6970
rect -1950 6880 -1850 6890
rect 11800 6880 11900 6890
rect -490 6070 -390 6080
rect 9910 6070 10010 6080
rect -940 5990 -480 6070
rect -400 5990 9920 6070
rect 10000 5990 11060 6070
rect -490 5980 -390 5990
rect 9910 5980 10010 5990
rect -490 -230 -390 -220
rect 9910 -230 10010 -220
rect -940 -310 -480 -230
rect -400 -310 9920 -230
rect 10000 -310 11060 -230
rect -490 -320 -390 -310
rect 9910 -320 10010 -310
rect -1950 -1230 -1850 -1220
rect 11800 -1230 11900 -1220
rect -2830 -1310 -1940 -1230
rect -1860 -1310 11810 -1230
rect 11890 -1310 12840 -1230
rect -1950 -1320 -1850 -1310
rect 11800 -1320 11900 -1310
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 -10 0 1 0
box 0 0 1340 1340
<< labels >>
flabel locali s 4660 1102 4778 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 4683 1252 4784 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 4624 626 4872 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 6020 1102 6138 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 6043 1252 6144 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 5984 626 6232 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 7380 1102 7498 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 7403 1252 7504 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 7344 626 7592 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 8740 1102 8858 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 8763 1252 8864 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 8704 626 8952 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 3264 626 3512 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 3323 1252 3424 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 3300 1102 3418 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 1940 1102 2058 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 1963 1252 2064 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 1904 626 2152 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
<< end >>
