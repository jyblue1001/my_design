magic
tech sky130A
timestamp 1739803560
<< psubdiff >>
rect 2600 -6165 2650 -6150
rect 2600 -6185 2615 -6165
rect 2635 -6185 2650 -6165
rect 2600 -6200 2650 -6185
<< psubdiffcont >>
rect 2615 -6185 2635 -6165
<< xpolycontact >>
rect 5520 195 5740 230
rect 6476 195 6696 230
<< xpolyres >>
rect 5740 195 6476 230
<< locali >>
rect 1135 220 1185 230
rect 1135 190 1145 220
rect 1175 190 1185 220
rect 5480 225 5520 230
rect 5480 200 5485 225
rect 5510 200 5520 225
rect 5480 195 5520 200
rect 6696 225 6736 230
rect 6696 200 6706 225
rect 6731 200 6736 225
rect 6696 195 6736 200
rect 1135 180 1185 190
rect 2475 -6105 2530 -6095
rect 2475 -6140 2485 -6105
rect 2520 -6130 2530 -6105
rect 2725 -6105 2780 -6095
rect 2725 -6130 2735 -6105
rect 2520 -6140 2735 -6130
rect 2770 -6140 2780 -6105
rect 2475 -6150 2780 -6140
rect 2600 -6165 2650 -6150
rect 2600 -6185 2615 -6165
rect 2635 -6185 2650 -6165
rect 2600 -6200 2650 -6185
<< viali >>
rect 1145 190 1175 220
rect 5485 200 5510 225
rect 6706 200 6731 225
rect 2485 -6140 2520 -6105
rect 2735 -6140 2770 -6105
<< metal1 >>
rect 1135 225 5520 230
rect 1135 220 5485 225
rect 1135 190 1145 220
rect 1175 200 5485 220
rect 5510 200 5520 225
rect 1175 195 5520 200
rect 6695 225 9720 230
rect 6695 200 6706 225
rect 6731 220 9720 225
rect 6731 200 9680 220
rect 6695 195 9680 200
rect 1175 190 1185 195
rect 1135 180 1185 190
rect 9670 190 9680 195
rect 9710 190 9720 220
rect 9670 180 9720 190
rect 2475 -6105 2530 -6095
rect 2475 -6140 2485 -6105
rect 2520 -6140 2530 -6105
rect 2475 -6150 2530 -6140
rect 2725 -6105 2780 -6095
rect 2725 -6140 2735 -6105
rect 2770 -6140 2780 -6105
rect 2725 -6150 2780 -6140
<< via1 >>
rect 1145 190 1175 220
rect 9680 190 9710 220
rect 2485 -6140 2520 -6105
rect 2735 -6140 2770 -6105
<< metal2 >>
rect 1135 220 1185 230
rect 1135 190 1145 220
rect 1175 190 1185 220
rect 1135 180 1185 190
rect 9670 220 9720 230
rect 9670 190 9680 220
rect 9710 190 9720 220
rect 9670 180 9720 190
rect 2475 -6105 2530 -6095
rect 2475 -6140 2485 -6105
rect 2520 -6140 2530 -6105
rect 2475 -6150 2530 -6140
rect 2725 -6105 2780 -6095
rect 2725 -6140 2735 -6105
rect 2770 -6140 2780 -6105
rect 2725 -6150 2780 -6140
<< via2 >>
rect 1145 190 1175 220
rect 9680 190 9710 220
rect 2485 -6140 2520 -6105
rect 2735 -6140 2770 -6105
<< metal3 >>
rect 1135 220 1185 230
rect 1135 190 1145 220
rect 1175 190 1185 220
rect 1135 55 1185 190
rect 9670 220 9720 230
rect 9670 190 9680 220
rect 9710 190 9720 220
rect 9670 55 9720 190
rect 1135 -5975 2545 55
rect 2710 -5975 9720 55
rect 2475 -6105 2530 -6095
rect 2475 -6140 2485 -6105
rect 2520 -6140 2530 -6105
rect 2475 -6150 2530 -6140
rect 2725 -6105 2780 -6095
rect 2725 -6140 2735 -6105
rect 2770 -6140 2780 -6105
rect 2725 -6150 2780 -6140
<< via3 >>
rect 2485 -6140 2520 -6105
rect 2735 -6140 2770 -6105
<< mimcap >>
rect 1150 -5915 2530 40
rect 1150 -5950 2485 -5915
rect 2520 -5950 2530 -5915
rect 1150 -5960 2530 -5950
rect 2725 -5915 9705 40
rect 2725 -5950 2735 -5915
rect 2770 -5950 9705 -5915
rect 2725 -5960 9705 -5950
<< mimcapcontact >>
rect 2485 -5950 2520 -5915
rect 2735 -5950 2770 -5915
<< metal4 >>
rect 2475 -5915 2530 -5910
rect 2475 -5950 2485 -5915
rect 2520 -5950 2530 -5915
rect 2475 -6105 2530 -5950
rect 2475 -6140 2485 -6105
rect 2520 -6140 2530 -6105
rect 2475 -6150 2530 -6140
rect 2725 -5915 2780 -5910
rect 2725 -5950 2735 -5915
rect 2770 -5950 2780 -5915
rect 2725 -6105 2780 -5950
rect 2725 -6140 2735 -6105
rect 2770 -6140 2780 -6105
rect 2725 -6150 2780 -6140
<< labels >>
flabel locali 2625 -6150 2625 -6150 5 FreeSans 800 0 0 -400 GNDA
port 2 s
flabel metal1 2620 230 2620 230 1 FreeSans 800 0 0 400 V_OUT
port 1 n
flabel metal1 8230 230 8230 230 1 FreeSans 800 0 0 400 R1_C1
<< end >>
